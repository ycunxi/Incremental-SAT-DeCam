module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);

input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;//RE__PI;

input s_0,s_1;//RE__ALLOW(00,01,10,11);
input s_2,s_3;//RE__ALLOW(00,01,10,11);
input s_4,s_5;//RE__ALLOW(00,01,10,11);
input s_6,s_7;//RE__ALLOW(00,01,10,11);
input s_8,s_9;//RE__ALLOW(00,01,10,11);
input s_10,s_11;//RE__ALLOW(00,01,10,11);
input s_12,s_13;//RE__ALLOW(00,01,10,11);
input s_14,s_15;//RE__ALLOW(00,01,10,11);
input s_16,s_17;//RE__ALLOW(00,01,10,11);
input s_18,s_19;//RE__ALLOW(00,01,10,11);
input s_20,s_21;//RE__ALLOW(00,01,10,11);
input s_22,s_23;//RE__ALLOW(00,01,10,11);
input s_24,s_25;//RE__ALLOW(00,01,10,11);
input s_26,s_27;//RE__ALLOW(00,01,10,11);
input s_28,s_29;//RE__ALLOW(00,01,10,11);
input s_30,s_31;//RE__ALLOW(00,01,10,11);
input s_32,s_33;//RE__ALLOW(00,01,10,11);
input s_34,s_35;//RE__ALLOW(00,01,10,11);
input s_36,s_37;//RE__ALLOW(00,01,10,11);
input s_38,s_39;//RE__ALLOW(00,01,10,11);
input s_40,s_41;//RE__ALLOW(00,01,10,11);
input s_42,s_43;//RE__ALLOW(00,01,10,11);
input s_44,s_45;//RE__ALLOW(00,01,10,11);
input s_46,s_47;//RE__ALLOW(00,01,10,11);
input s_48,s_49;//RE__ALLOW(00,01,10,11);
input s_50,s_51;//RE__ALLOW(00,01,10,11);
input s_52,s_53;//RE__ALLOW(00,01,10,11);
input s_54,s_55;//RE__ALLOW(00,01,10,11);
input s_56,s_57;//RE__ALLOW(00,01,10,11);
input s_58,s_59;//RE__ALLOW(00,01,10,11);
input s_60,s_61;//RE__ALLOW(00,01,10,11);
input s_62,s_63;//RE__ALLOW(00,01,10,11);
input s_64,s_65;//RE__ALLOW(00,01,10,11);
input s_66,s_67;//RE__ALLOW(00,01,10,11);
input s_68,s_69;//RE__ALLOW(00,01,10,11);
input s_70,s_71;//RE__ALLOW(00,01,10,11);
input s_72,s_73;//RE__ALLOW(00,01,10,11);
input s_74,s_75;//RE__ALLOW(00,01,10,11);
input s_76,s_77;//RE__ALLOW(00,01,10,11);
input s_78,s_79;//RE__ALLOW(00,01,10,11);
input s_80,s_81;//RE__ALLOW(00,01,10,11);
input s_82,s_83;//RE__ALLOW(00,01,10,11);
input s_84,s_85;//RE__ALLOW(00,01,10,11);
input s_86,s_87;//RE__ALLOW(00,01,10,11);
input s_88,s_89;//RE__ALLOW(00,01,10,11);
input s_90,s_91;//RE__ALLOW(00,01,10,11);
input s_92,s_93;//RE__ALLOW(00,01,10,11);
input s_94,s_95;//RE__ALLOW(00,01,10,11);
input s_96,s_97;//RE__ALLOW(00,01,10,11);
input s_98,s_99;//RE__ALLOW(00,01,10,11);
input s_100,s_101;//RE__ALLOW(00,01,10,11);
input s_102,s_103;//RE__ALLOW(00,01,10,11);
input s_104,s_105;//RE__ALLOW(00,01,10,11);
input s_106,s_107;//RE__ALLOW(00,01,10,11);
input s_108,s_109;//RE__ALLOW(00,01,10,11);
input s_110,s_111;//RE__ALLOW(00,01,10,11);
input s_112,s_113;//RE__ALLOW(00,01,10,11);
input s_114,s_115;//RE__ALLOW(00,01,10,11);
input s_116,s_117;//RE__ALLOW(00,01,10,11);
input s_118,s_119;//RE__ALLOW(00,01,10,11);
input s_120,s_121;//RE__ALLOW(00,01,10,11);
input s_122,s_123;//RE__ALLOW(00,01,10,11);
input s_124,s_125;//RE__ALLOW(00,01,10,11);
input s_126,s_127;//RE__ALLOW(00,01,10,11);
input s_128,s_129;//RE__ALLOW(00,01,10,11);
input s_130,s_131;//RE__ALLOW(00,01,10,11);
input s_132,s_133;//RE__ALLOW(00,01,10,11);
input s_134,s_135;//RE__ALLOW(00,01,10,11);
input s_136,s_137;//RE__ALLOW(00,01,10,11);
input s_138,s_139;//RE__ALLOW(00,01,10,11);
input s_140,s_141;//RE__ALLOW(00,01,10,11);
input s_142,s_143;//RE__ALLOW(00,01,10,11);
input s_144,s_145;//RE__ALLOW(00,01,10,11);
input s_146,s_147;//RE__ALLOW(00,01,10,11);
input s_148,s_149;//RE__ALLOW(00,01,10,11);
input s_150,s_151;//RE__ALLOW(00,01,10,11);
input s_152,s_153;//RE__ALLOW(00,01,10,11);
input s_154,s_155;//RE__ALLOW(00,01,10,11);
input s_156,s_157;//RE__ALLOW(00,01,10,11);
input s_158,s_159;//RE__ALLOW(00,01,10,11);
input s_160,s_161;//RE__ALLOW(00,01,10,11);
input s_162,s_163;//RE__ALLOW(00,01,10,11);
input s_164,s_165;//RE__ALLOW(00,01,10,11);
input s_166,s_167;//RE__ALLOW(00,01,10,11);
input s_168,s_169;//RE__ALLOW(00,01,10,11);
input s_170,s_171;//RE__ALLOW(00,01,10,11);
input s_172,s_173;//RE__ALLOW(00,01,10,11);
input s_174,s_175;//RE__ALLOW(00,01,10,11);
input s_176,s_177;//RE__ALLOW(00,01,10,11);
input s_178,s_179;//RE__ALLOW(00,01,10,11);
input s_180,s_181;//RE__ALLOW(00,01,10,11);
input s_182,s_183;//RE__ALLOW(00,01,10,11);
input s_184,s_185;//RE__ALLOW(00,01,10,11);
input s_186,s_187;//RE__ALLOW(00,01,10,11);
input s_188,s_189;//RE__ALLOW(00,01,10,11);
input s_190,s_191;//RE__ALLOW(00,01,10,11);
input s_192,s_193;//RE__ALLOW(00,01,10,11);
input s_194,s_195;//RE__ALLOW(00,01,10,11);
input s_196,s_197;//RE__ALLOW(00,01,10,11);
input s_198,s_199;//RE__ALLOW(00,01,10,11);
input s_200,s_201;//RE__ALLOW(00,01,10,11);
input s_202,s_203;//RE__ALLOW(00,01,10,11);
input s_204,s_205;//RE__ALLOW(00,01,10,11);
input s_206,s_207;//RE__ALLOW(00,01,10,11);
input s_208,s_209;//RE__ALLOW(00,01,10,11);
input s_210,s_211;//RE__ALLOW(00,01,10,11);
input s_212,s_213;//RE__ALLOW(00,01,10,11);
input s_214,s_215;//RE__ALLOW(00,01,10,11);
input s_216,s_217;//RE__ALLOW(00,01,10,11);
input s_218,s_219;//RE__ALLOW(00,01,10,11);
input s_220,s_221;//RE__ALLOW(00,01,10,11);
input s_222,s_223;//RE__ALLOW(00,01,10,11);
input s_224,s_225;//RE__ALLOW(00,01,10,11);
input s_226,s_227;//RE__ALLOW(00,01,10,11);
input s_228,s_229;//RE__ALLOW(00,01,10,11);
input s_230,s_231;//RE__ALLOW(00,01,10,11);
input s_232,s_233;//RE__ALLOW(00,01,10,11);
input s_234,s_235;//RE__ALLOW(00,01,10,11);
input s_236,s_237;//RE__ALLOW(00,01,10,11);
input s_238,s_239;//RE__ALLOW(00,01,10,11);
input s_240,s_241;//RE__ALLOW(00,01,10,11);
input s_242,s_243;//RE__ALLOW(00,01,10,11);
input s_244,s_245;//RE__ALLOW(00,01,10,11);
input s_246,s_247;//RE__ALLOW(00,01,10,11);
input s_248,s_249;//RE__ALLOW(00,01,10,11);
input s_250,s_251;//RE__ALLOW(00,01,10,11);
input s_252,s_253;//RE__ALLOW(00,01,10,11);
input s_254,s_255;//RE__ALLOW(00,01,10,11);
input s_256,s_257;//RE__ALLOW(00,01,10,11);
input s_258,s_259;//RE__ALLOW(00,01,10,11);
input s_260,s_261;//RE__ALLOW(00,01,10,11);
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;

  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate235inter0, gate235inter1, gate235inter2, gate235inter3, gate235inter4, gate235inter5, gate235inter6, gate235inter7, gate235inter8, gate235inter9, gate235inter10, gate235inter11, gate235inter12, gate244inter0, gate244inter1, gate244inter2, gate244inter3, gate244inter4, gate244inter5, gate244inter6, gate244inter7, gate244inter8, gate244inter9, gate244inter10, gate244inter11, gate244inter12, gate179inter0, gate179inter1, gate179inter2, gate179inter3, gate179inter4, gate179inter5, gate179inter6, gate179inter7, gate179inter8, gate179inter9, gate179inter10, gate179inter11, gate179inter12, gate128inter0, gate128inter1, gate128inter2, gate128inter3, gate128inter4, gate128inter5, gate128inter6, gate128inter7, gate128inter8, gate128inter9, gate128inter10, gate128inter11, gate128inter12, gate63inter0, gate63inter1, gate63inter2, gate63inter3, gate63inter4, gate63inter5, gate63inter6, gate63inter7, gate63inter8, gate63inter9, gate63inter10, gate63inter11, gate63inter12, gate495inter0, gate495inter1, gate495inter2, gate495inter3, gate495inter4, gate495inter5, gate495inter6, gate495inter7, gate495inter8, gate495inter9, gate495inter10, gate495inter11, gate495inter12, gate489inter0, gate489inter1, gate489inter2, gate489inter3, gate489inter4, gate489inter5, gate489inter6, gate489inter7, gate489inter8, gate489inter9, gate489inter10, gate489inter11, gate489inter12, gate438inter0, gate438inter1, gate438inter2, gate438inter3, gate438inter4, gate438inter5, gate438inter6, gate438inter7, gate438inter8, gate438inter9, gate438inter10, gate438inter11, gate438inter12, gate54inter0, gate54inter1, gate54inter2, gate54inter3, gate54inter4, gate54inter5, gate54inter6, gate54inter7, gate54inter8, gate54inter9, gate54inter10, gate54inter11, gate54inter12, gate263inter0, gate263inter1, gate263inter2, gate263inter3, gate263inter4, gate263inter5, gate263inter6, gate263inter7, gate263inter8, gate263inter9, gate263inter10, gate263inter11, gate263inter12, gate406inter0, gate406inter1, gate406inter2, gate406inter3, gate406inter4, gate406inter5, gate406inter6, gate406inter7, gate406inter8, gate406inter9, gate406inter10, gate406inter11, gate406inter12, gate290inter0, gate290inter1, gate290inter2, gate290inter3, gate290inter4, gate290inter5, gate290inter6, gate290inter7, gate290inter8, gate290inter9, gate290inter10, gate290inter11, gate290inter12, gate223inter0, gate223inter1, gate223inter2, gate223inter3, gate223inter4, gate223inter5, gate223inter6, gate223inter7, gate223inter8, gate223inter9, gate223inter10, gate223inter11, gate223inter12, gate131inter0, gate131inter1, gate131inter2, gate131inter3, gate131inter4, gate131inter5, gate131inter6, gate131inter7, gate131inter8, gate131inter9, gate131inter10, gate131inter11, gate131inter12, gate194inter0, gate194inter1, gate194inter2, gate194inter3, gate194inter4, gate194inter5, gate194inter6, gate194inter7, gate194inter8, gate194inter9, gate194inter10, gate194inter11, gate194inter12, gate472inter0, gate472inter1, gate472inter2, gate472inter3, gate472inter4, gate472inter5, gate472inter6, gate472inter7, gate472inter8, gate472inter9, gate472inter10, gate472inter11, gate472inter12, gate512inter0, gate512inter1, gate512inter2, gate512inter3, gate512inter4, gate512inter5, gate512inter6, gate512inter7, gate512inter8, gate512inter9, gate512inter10, gate512inter11, gate512inter12, gate473inter0, gate473inter1, gate473inter2, gate473inter3, gate473inter4, gate473inter5, gate473inter6, gate473inter7, gate473inter8, gate473inter9, gate473inter10, gate473inter11, gate473inter12, gate216inter0, gate216inter1, gate216inter2, gate216inter3, gate216inter4, gate216inter5, gate216inter6, gate216inter7, gate216inter8, gate216inter9, gate216inter10, gate216inter11, gate216inter12, gate31inter0, gate31inter1, gate31inter2, gate31inter3, gate31inter4, gate31inter5, gate31inter6, gate31inter7, gate31inter8, gate31inter9, gate31inter10, gate31inter11, gate31inter12, gate504inter0, gate504inter1, gate504inter2, gate504inter3, gate504inter4, gate504inter5, gate504inter6, gate504inter7, gate504inter8, gate504inter9, gate504inter10, gate504inter11, gate504inter12, gate85inter0, gate85inter1, gate85inter2, gate85inter3, gate85inter4, gate85inter5, gate85inter6, gate85inter7, gate85inter8, gate85inter9, gate85inter10, gate85inter11, gate85inter12, gate393inter0, gate393inter1, gate393inter2, gate393inter3, gate393inter4, gate393inter5, gate393inter6, gate393inter7, gate393inter8, gate393inter9, gate393inter10, gate393inter11, gate393inter12, gate38inter0, gate38inter1, gate38inter2, gate38inter3, gate38inter4, gate38inter5, gate38inter6, gate38inter7, gate38inter8, gate38inter9, gate38inter10, gate38inter11, gate38inter12, gate414inter0, gate414inter1, gate414inter2, gate414inter3, gate414inter4, gate414inter5, gate414inter6, gate414inter7, gate414inter8, gate414inter9, gate414inter10, gate414inter11, gate414inter12, gate109inter0, gate109inter1, gate109inter2, gate109inter3, gate109inter4, gate109inter5, gate109inter6, gate109inter7, gate109inter8, gate109inter9, gate109inter10, gate109inter11, gate109inter12, gate165inter0, gate165inter1, gate165inter2, gate165inter3, gate165inter4, gate165inter5, gate165inter6, gate165inter7, gate165inter8, gate165inter9, gate165inter10, gate165inter11, gate165inter12, gate460inter0, gate460inter1, gate460inter2, gate460inter3, gate460inter4, gate460inter5, gate460inter6, gate460inter7, gate460inter8, gate460inter9, gate460inter10, gate460inter11, gate460inter12, gate494inter0, gate494inter1, gate494inter2, gate494inter3, gate494inter4, gate494inter5, gate494inter6, gate494inter7, gate494inter8, gate494inter9, gate494inter10, gate494inter11, gate494inter12, gate14inter0, gate14inter1, gate14inter2, gate14inter3, gate14inter4, gate14inter5, gate14inter6, gate14inter7, gate14inter8, gate14inter9, gate14inter10, gate14inter11, gate14inter12, gate87inter0, gate87inter1, gate87inter2, gate87inter3, gate87inter4, gate87inter5, gate87inter6, gate87inter7, gate87inter8, gate87inter9, gate87inter10, gate87inter11, gate87inter12, gate409inter0, gate409inter1, gate409inter2, gate409inter3, gate409inter4, gate409inter5, gate409inter6, gate409inter7, gate409inter8, gate409inter9, gate409inter10, gate409inter11, gate409inter12, gate420inter0, gate420inter1, gate420inter2, gate420inter3, gate420inter4, gate420inter5, gate420inter6, gate420inter7, gate420inter8, gate420inter9, gate420inter10, gate420inter11, gate420inter12, gate49inter0, gate49inter1, gate49inter2, gate49inter3, gate49inter4, gate49inter5, gate49inter6, gate49inter7, gate49inter8, gate49inter9, gate49inter10, gate49inter11, gate49inter12, gate52inter0, gate52inter1, gate52inter2, gate52inter3, gate52inter4, gate52inter5, gate52inter6, gate52inter7, gate52inter8, gate52inter9, gate52inter10, gate52inter11, gate52inter12, gate261inter0, gate261inter1, gate261inter2, gate261inter3, gate261inter4, gate261inter5, gate261inter6, gate261inter7, gate261inter8, gate261inter9, gate261inter10, gate261inter11, gate261inter12, gate18inter0, gate18inter1, gate18inter2, gate18inter3, gate18inter4, gate18inter5, gate18inter6, gate18inter7, gate18inter8, gate18inter9, gate18inter10, gate18inter11, gate18inter12, gate514inter0, gate514inter1, gate514inter2, gate514inter3, gate514inter4, gate514inter5, gate514inter6, gate514inter7, gate514inter8, gate514inter9, gate514inter10, gate514inter11, gate514inter12, gate278inter0, gate278inter1, gate278inter2, gate278inter3, gate278inter4, gate278inter5, gate278inter6, gate278inter7, gate278inter8, gate278inter9, gate278inter10, gate278inter11, gate278inter12, gate488inter0, gate488inter1, gate488inter2, gate488inter3, gate488inter4, gate488inter5, gate488inter6, gate488inter7, gate488inter8, gate488inter9, gate488inter10, gate488inter11, gate488inter12, gate390inter0, gate390inter1, gate390inter2, gate390inter3, gate390inter4, gate390inter5, gate390inter6, gate390inter7, gate390inter8, gate390inter9, gate390inter10, gate390inter11, gate390inter12, gate105inter0, gate105inter1, gate105inter2, gate105inter3, gate105inter4, gate105inter5, gate105inter6, gate105inter7, gate105inter8, gate105inter9, gate105inter10, gate105inter11, gate105inter12, gate466inter0, gate466inter1, gate466inter2, gate466inter3, gate466inter4, gate466inter5, gate466inter6, gate466inter7, gate466inter8, gate466inter9, gate466inter10, gate466inter11, gate466inter12, gate29inter0, gate29inter1, gate29inter2, gate29inter3, gate29inter4, gate29inter5, gate29inter6, gate29inter7, gate29inter8, gate29inter9, gate29inter10, gate29inter11, gate29inter12, gate78inter0, gate78inter1, gate78inter2, gate78inter3, gate78inter4, gate78inter5, gate78inter6, gate78inter7, gate78inter8, gate78inter9, gate78inter10, gate78inter11, gate78inter12, gate62inter0, gate62inter1, gate62inter2, gate62inter3, gate62inter4, gate62inter5, gate62inter6, gate62inter7, gate62inter8, gate62inter9, gate62inter10, gate62inter11, gate62inter12, gate454inter0, gate454inter1, gate454inter2, gate454inter3, gate454inter4, gate454inter5, gate454inter6, gate454inter7, gate454inter8, gate454inter9, gate454inter10, gate454inter11, gate454inter12, gate187inter0, gate187inter1, gate187inter2, gate187inter3, gate187inter4, gate187inter5, gate187inter6, gate187inter7, gate187inter8, gate187inter9, gate187inter10, gate187inter11, gate187inter12, gate441inter0, gate441inter1, gate441inter2, gate441inter3, gate441inter4, gate441inter5, gate441inter6, gate441inter7, gate441inter8, gate441inter9, gate441inter10, gate441inter11, gate441inter12, gate426inter0, gate426inter1, gate426inter2, gate426inter3, gate426inter4, gate426inter5, gate426inter6, gate426inter7, gate426inter8, gate426inter9, gate426inter10, gate426inter11, gate426inter12, gate401inter0, gate401inter1, gate401inter2, gate401inter3, gate401inter4, gate401inter5, gate401inter6, gate401inter7, gate401inter8, gate401inter9, gate401inter10, gate401inter11, gate401inter12, gate37inter0, gate37inter1, gate37inter2, gate37inter3, gate37inter4, gate37inter5, gate37inter6, gate37inter7, gate37inter8, gate37inter9, gate37inter10, gate37inter11, gate37inter12, gate205inter0, gate205inter1, gate205inter2, gate205inter3, gate205inter4, gate205inter5, gate205inter6, gate205inter7, gate205inter8, gate205inter9, gate205inter10, gate205inter11, gate205inter12, gate161inter0, gate161inter1, gate161inter2, gate161inter3, gate161inter4, gate161inter5, gate161inter6, gate161inter7, gate161inter8, gate161inter9, gate161inter10, gate161inter11, gate161inter12, gate293inter0, gate293inter1, gate293inter2, gate293inter3, gate293inter4, gate293inter5, gate293inter6, gate293inter7, gate293inter8, gate293inter9, gate293inter10, gate293inter11, gate293inter12, gate243inter0, gate243inter1, gate243inter2, gate243inter3, gate243inter4, gate243inter5, gate243inter6, gate243inter7, gate243inter8, gate243inter9, gate243inter10, gate243inter11, gate243inter12, gate248inter0, gate248inter1, gate248inter2, gate248inter3, gate248inter4, gate248inter5, gate248inter6, gate248inter7, gate248inter8, gate248inter9, gate248inter10, gate248inter11, gate248inter12, gate189inter0, gate189inter1, gate189inter2, gate189inter3, gate189inter4, gate189inter5, gate189inter6, gate189inter7, gate189inter8, gate189inter9, gate189inter10, gate189inter11, gate189inter12, gate141inter0, gate141inter1, gate141inter2, gate141inter3, gate141inter4, gate141inter5, gate141inter6, gate141inter7, gate141inter8, gate141inter9, gate141inter10, gate141inter11, gate141inter12, gate91inter0, gate91inter1, gate91inter2, gate91inter3, gate91inter4, gate91inter5, gate91inter6, gate91inter7, gate91inter8, gate91inter9, gate91inter10, gate91inter11, gate91inter12, gate180inter0, gate180inter1, gate180inter2, gate180inter3, gate180inter4, gate180inter5, gate180inter6, gate180inter7, gate180inter8, gate180inter9, gate180inter10, gate180inter11, gate180inter12, gate213inter0, gate213inter1, gate213inter2, gate213inter3, gate213inter4, gate213inter5, gate213inter6, gate213inter7, gate213inter8, gate213inter9, gate213inter10, gate213inter11, gate213inter12, gate186inter0, gate186inter1, gate186inter2, gate186inter3, gate186inter4, gate186inter5, gate186inter6, gate186inter7, gate186inter8, gate186inter9, gate186inter10, gate186inter11, gate186inter12, gate285inter0, gate285inter1, gate285inter2, gate285inter3, gate285inter4, gate285inter5, gate285inter6, gate285inter7, gate285inter8, gate285inter9, gate285inter10, gate285inter11, gate285inter12, gate191inter0, gate191inter1, gate191inter2, gate191inter3, gate191inter4, gate191inter5, gate191inter6, gate191inter7, gate191inter8, gate191inter9, gate191inter10, gate191inter11, gate191inter12, gate166inter0, gate166inter1, gate166inter2, gate166inter3, gate166inter4, gate166inter5, gate166inter6, gate166inter7, gate166inter8, gate166inter9, gate166inter10, gate166inter11, gate166inter12, gate174inter0, gate174inter1, gate174inter2, gate174inter3, gate174inter4, gate174inter5, gate174inter6, gate174inter7, gate174inter8, gate174inter9, gate174inter10, gate174inter11, gate174inter12, gate56inter0, gate56inter1, gate56inter2, gate56inter3, gate56inter4, gate56inter5, gate56inter6, gate56inter7, gate56inter8, gate56inter9, gate56inter10, gate56inter11, gate56inter12, gate465inter0, gate465inter1, gate465inter2, gate465inter3, gate465inter4, gate465inter5, gate465inter6, gate465inter7, gate465inter8, gate465inter9, gate465inter10, gate465inter11, gate465inter12, gate136inter0, gate136inter1, gate136inter2, gate136inter3, gate136inter4, gate136inter5, gate136inter6, gate136inter7, gate136inter8, gate136inter9, gate136inter10, gate136inter11, gate136inter12, gate492inter0, gate492inter1, gate492inter2, gate492inter3, gate492inter4, gate492inter5, gate492inter6, gate492inter7, gate492inter8, gate492inter9, gate492inter10, gate492inter11, gate492inter12, gate28inter0, gate28inter1, gate28inter2, gate28inter3, gate28inter4, gate28inter5, gate28inter6, gate28inter7, gate28inter8, gate28inter9, gate28inter10, gate28inter11, gate28inter12, gate397inter0, gate397inter1, gate397inter2, gate397inter3, gate397inter4, gate397inter5, gate397inter6, gate397inter7, gate397inter8, gate397inter9, gate397inter10, gate397inter11, gate397inter12, gate267inter0, gate267inter1, gate267inter2, gate267inter3, gate267inter4, gate267inter5, gate267inter6, gate267inter7, gate267inter8, gate267inter9, gate267inter10, gate267inter11, gate267inter12, gate119inter0, gate119inter1, gate119inter2, gate119inter3, gate119inter4, gate119inter5, gate119inter6, gate119inter7, gate119inter8, gate119inter9, gate119inter10, gate119inter11, gate119inter12, gate160inter0, gate160inter1, gate160inter2, gate160inter3, gate160inter4, gate160inter5, gate160inter6, gate160inter7, gate160inter8, gate160inter9, gate160inter10, gate160inter11, gate160inter12, gate132inter0, gate132inter1, gate132inter2, gate132inter3, gate132inter4, gate132inter5, gate132inter6, gate132inter7, gate132inter8, gate132inter9, gate132inter10, gate132inter11, gate132inter12, gate169inter0, gate169inter1, gate169inter2, gate169inter3, gate169inter4, gate169inter5, gate169inter6, gate169inter7, gate169inter8, gate169inter9, gate169inter10, gate169inter11, gate169inter12, gate25inter0, gate25inter1, gate25inter2, gate25inter3, gate25inter4, gate25inter5, gate25inter6, gate25inter7, gate25inter8, gate25inter9, gate25inter10, gate25inter11, gate25inter12, gate92inter0, gate92inter1, gate92inter2, gate92inter3, gate92inter4, gate92inter5, gate92inter6, gate92inter7, gate92inter8, gate92inter9, gate92inter10, gate92inter11, gate92inter12, gate148inter0, gate148inter1, gate148inter2, gate148inter3, gate148inter4, gate148inter5, gate148inter6, gate148inter7, gate148inter8, gate148inter9, gate148inter10, gate148inter11, gate148inter12, gate158inter0, gate158inter1, gate158inter2, gate158inter3, gate158inter4, gate158inter5, gate158inter6, gate158inter7, gate158inter8, gate158inter9, gate158inter10, gate158inter11, gate158inter12, gate500inter0, gate500inter1, gate500inter2, gate500inter3, gate500inter4, gate500inter5, gate500inter6, gate500inter7, gate500inter8, gate500inter9, gate500inter10, gate500inter11, gate500inter12, gate118inter0, gate118inter1, gate118inter2, gate118inter3, gate118inter4, gate118inter5, gate118inter6, gate118inter7, gate118inter8, gate118inter9, gate118inter10, gate118inter11, gate118inter12, gate21inter0, gate21inter1, gate21inter2, gate21inter3, gate21inter4, gate21inter5, gate21inter6, gate21inter7, gate21inter8, gate21inter9, gate21inter10, gate21inter11, gate21inter12, gate455inter0, gate455inter1, gate455inter2, gate455inter3, gate455inter4, gate455inter5, gate455inter6, gate455inter7, gate455inter8, gate455inter9, gate455inter10, gate455inter11, gate455inter12, gate266inter0, gate266inter1, gate266inter2, gate266inter3, gate266inter4, gate266inter5, gate266inter6, gate266inter7, gate266inter8, gate266inter9, gate266inter10, gate266inter11, gate266inter12, gate9inter0, gate9inter1, gate9inter2, gate9inter3, gate9inter4, gate9inter5, gate9inter6, gate9inter7, gate9inter8, gate9inter9, gate9inter10, gate9inter11, gate9inter12, gate416inter0, gate416inter1, gate416inter2, gate416inter3, gate416inter4, gate416inter5, gate416inter6, gate416inter7, gate416inter8, gate416inter9, gate416inter10, gate416inter11, gate416inter12, gate237inter0, gate237inter1, gate237inter2, gate237inter3, gate237inter4, gate237inter5, gate237inter6, gate237inter7, gate237inter8, gate237inter9, gate237inter10, gate237inter11, gate237inter12, gate96inter0, gate96inter1, gate96inter2, gate96inter3, gate96inter4, gate96inter5, gate96inter6, gate96inter7, gate96inter8, gate96inter9, gate96inter10, gate96inter11, gate96inter12, gate172inter0, gate172inter1, gate172inter2, gate172inter3, gate172inter4, gate172inter5, gate172inter6, gate172inter7, gate172inter8, gate172inter9, gate172inter10, gate172inter11, gate172inter12, gate392inter0, gate392inter1, gate392inter2, gate392inter3, gate392inter4, gate392inter5, gate392inter6, gate392inter7, gate392inter8, gate392inter9, gate392inter10, gate392inter11, gate392inter12, gate487inter0, gate487inter1, gate487inter2, gate487inter3, gate487inter4, gate487inter5, gate487inter6, gate487inter7, gate487inter8, gate487inter9, gate487inter10, gate487inter11, gate487inter12, gate238inter0, gate238inter1, gate238inter2, gate238inter3, gate238inter4, gate238inter5, gate238inter6, gate238inter7, gate238inter8, gate238inter9, gate238inter10, gate238inter11, gate238inter12, gate19inter0, gate19inter1, gate19inter2, gate19inter3, gate19inter4, gate19inter5, gate19inter6, gate19inter7, gate19inter8, gate19inter9, gate19inter10, gate19inter11, gate19inter12, gate102inter0, gate102inter1, gate102inter2, gate102inter3, gate102inter4, gate102inter5, gate102inter6, gate102inter7, gate102inter8, gate102inter9, gate102inter10, gate102inter11, gate102inter12, gate188inter0, gate188inter1, gate188inter2, gate188inter3, gate188inter4, gate188inter5, gate188inter6, gate188inter7, gate188inter8, gate188inter9, gate188inter10, gate188inter11, gate188inter12, gate258inter0, gate258inter1, gate258inter2, gate258inter3, gate258inter4, gate258inter5, gate258inter6, gate258inter7, gate258inter8, gate258inter9, gate258inter10, gate258inter11, gate258inter12, gate61inter0, gate61inter1, gate61inter2, gate61inter3, gate61inter4, gate61inter5, gate61inter6, gate61inter7, gate61inter8, gate61inter9, gate61inter10, gate61inter11, gate61inter12, gate222inter0, gate222inter1, gate222inter2, gate222inter3, gate222inter4, gate222inter5, gate222inter6, gate222inter7, gate222inter8, gate222inter9, gate222inter10, gate222inter11, gate222inter12, gate120inter0, gate120inter1, gate120inter2, gate120inter3, gate120inter4, gate120inter5, gate120inter6, gate120inter7, gate120inter8, gate120inter9, gate120inter10, gate120inter11, gate120inter12, gate80inter0, gate80inter1, gate80inter2, gate80inter3, gate80inter4, gate80inter5, gate80inter6, gate80inter7, gate80inter8, gate80inter9, gate80inter10, gate80inter11, gate80inter12, gate51inter0, gate51inter1, gate51inter2, gate51inter3, gate51inter4, gate51inter5, gate51inter6, gate51inter7, gate51inter8, gate51inter9, gate51inter10, gate51inter11, gate51inter12, gate405inter0, gate405inter1, gate405inter2, gate405inter3, gate405inter4, gate405inter5, gate405inter6, gate405inter7, gate405inter8, gate405inter9, gate405inter10, gate405inter11, gate405inter12, gate499inter0, gate499inter1, gate499inter2, gate499inter3, gate499inter4, gate499inter5, gate499inter6, gate499inter7, gate499inter8, gate499inter9, gate499inter10, gate499inter11, gate499inter12, gate275inter0, gate275inter1, gate275inter2, gate275inter3, gate275inter4, gate275inter5, gate275inter6, gate275inter7, gate275inter8, gate275inter9, gate275inter10, gate275inter11, gate275inter12, gate402inter0, gate402inter1, gate402inter2, gate402inter3, gate402inter4, gate402inter5, gate402inter6, gate402inter7, gate402inter8, gate402inter9, gate402inter10, gate402inter11, gate402inter12, gate467inter0, gate467inter1, gate467inter2, gate467inter3, gate467inter4, gate467inter5, gate467inter6, gate467inter7, gate467inter8, gate467inter9, gate467inter10, gate467inter11, gate467inter12, gate506inter0, gate506inter1, gate506inter2, gate506inter3, gate506inter4, gate506inter5, gate506inter6, gate506inter7, gate506inter8, gate506inter9, gate506inter10, gate506inter11, gate506inter12, gate177inter0, gate177inter1, gate177inter2, gate177inter3, gate177inter4, gate177inter5, gate177inter6, gate177inter7, gate177inter8, gate177inter9, gate177inter10, gate177inter11, gate177inter12, gate196inter0, gate196inter1, gate196inter2, gate196inter3, gate196inter4, gate196inter5, gate196inter6, gate196inter7, gate196inter8, gate196inter9, gate196inter10, gate196inter11, gate196inter12, gate398inter0, gate398inter1, gate398inter2, gate398inter3, gate398inter4, gate398inter5, gate398inter6, gate398inter7, gate398inter8, gate398inter9, gate398inter10, gate398inter11, gate398inter12, gate291inter0, gate291inter1, gate291inter2, gate291inter3, gate291inter4, gate291inter5, gate291inter6, gate291inter7, gate291inter8, gate291inter9, gate291inter10, gate291inter11, gate291inter12, gate232inter0, gate232inter1, gate232inter2, gate232inter3, gate232inter4, gate232inter5, gate232inter6, gate232inter7, gate232inter8, gate232inter9, gate232inter10, gate232inter11, gate232inter12, gate430inter0, gate430inter1, gate430inter2, gate430inter3, gate430inter4, gate430inter5, gate430inter6, gate430inter7, gate430inter8, gate430inter9, gate430inter10, gate430inter11, gate430inter12, gate273inter0, gate273inter1, gate273inter2, gate273inter3, gate273inter4, gate273inter5, gate273inter6, gate273inter7, gate273inter8, gate273inter9, gate273inter10, gate273inter11, gate273inter12, gate207inter0, gate207inter1, gate207inter2, gate207inter3, gate207inter4, gate207inter5, gate207inter6, gate207inter7, gate207inter8, gate207inter9, gate207inter10, gate207inter11, gate207inter12, gate431inter0, gate431inter1, gate431inter2, gate431inter3, gate431inter4, gate431inter5, gate431inter6, gate431inter7, gate431inter8, gate431inter9, gate431inter10, gate431inter11, gate431inter12, gate27inter0, gate27inter1, gate27inter2, gate27inter3, gate27inter4, gate27inter5, gate27inter6, gate27inter7, gate27inter8, gate27inter9, gate27inter10, gate27inter11, gate27inter12, gate185inter0, gate185inter1, gate185inter2, gate185inter3, gate185inter4, gate185inter5, gate185inter6, gate185inter7, gate185inter8, gate185inter9, gate185inter10, gate185inter11, gate185inter12, gate427inter0, gate427inter1, gate427inter2, gate427inter3, gate427inter4, gate427inter5, gate427inter6, gate427inter7, gate427inter8, gate427inter9, gate427inter10, gate427inter11, gate427inter12, gate433inter0, gate433inter1, gate433inter2, gate433inter3, gate433inter4, gate433inter5, gate433inter6, gate433inter7, gate433inter8, gate433inter9, gate433inter10, gate433inter11, gate433inter12, gate264inter0, gate264inter1, gate264inter2, gate264inter3, gate264inter4, gate264inter5, gate264inter6, gate264inter7, gate264inter8, gate264inter9, gate264inter10, gate264inter11, gate264inter12, gate413inter0, gate413inter1, gate413inter2, gate413inter3, gate413inter4, gate413inter5, gate413inter6, gate413inter7, gate413inter8, gate413inter9, gate413inter10, gate413inter11, gate413inter12, gate47inter0, gate47inter1, gate47inter2, gate47inter3, gate47inter4, gate47inter5, gate47inter6, gate47inter7, gate47inter8, gate47inter9, gate47inter10, gate47inter11, gate47inter12, gate240inter0, gate240inter1, gate240inter2, gate240inter3, gate240inter4, gate240inter5, gate240inter6, gate240inter7, gate240inter8, gate240inter9, gate240inter10, gate240inter11, gate240inter12, gate15inter0, gate15inter1, gate15inter2, gate15inter3, gate15inter4, gate15inter5, gate15inter6, gate15inter7, gate15inter8, gate15inter9, gate15inter10, gate15inter11, gate15inter12, gate24inter0, gate24inter1, gate24inter2, gate24inter3, gate24inter4, gate24inter5, gate24inter6, gate24inter7, gate24inter8, gate24inter9, gate24inter10, gate24inter11, gate24inter12, gate39inter0, gate39inter1, gate39inter2, gate39inter3, gate39inter4, gate39inter5, gate39inter6, gate39inter7, gate39inter8, gate39inter9, gate39inter10, gate39inter11, gate39inter12, gate282inter0, gate282inter1, gate282inter2, gate282inter3, gate282inter4, gate282inter5, gate282inter6, gate282inter7, gate282inter8, gate282inter9, gate282inter10, gate282inter11, gate282inter12;



and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );

  xor2  gate1765(.a(G2), .b(G1), .O(gate9inter0));
  nand2 gate1766(.a(gate9inter0), .b(s_174), .O(gate9inter1));
  and2  gate1767(.a(G2), .b(G1), .O(gate9inter2));
  inv1  gate1768(.a(s_174), .O(gate9inter3));
  inv1  gate1769(.a(s_175), .O(gate9inter4));
  nand2 gate1770(.a(gate9inter4), .b(gate9inter3), .O(gate9inter5));
  nor2  gate1771(.a(gate9inter5), .b(gate9inter2), .O(gate9inter6));
  inv1  gate1772(.a(G1), .O(gate9inter7));
  inv1  gate1773(.a(G2), .O(gate9inter8));
  nand2 gate1774(.a(gate9inter8), .b(gate9inter7), .O(gate9inter9));
  nand2 gate1775(.a(s_175), .b(gate9inter3), .O(gate9inter10));
  nor2  gate1776(.a(gate9inter10), .b(gate9inter9), .O(gate9inter11));
  nor2  gate1777(.a(gate9inter11), .b(gate9inter6), .O(gate9inter12));
  nand2 gate1778(.a(gate9inter12), .b(gate9inter1), .O(G266));
nand2 gate10( .a(G3), .b(G4), .O(G269) );
nand2 gate11( .a(G5), .b(G6), .O(G272) );
nand2 gate12( .a(G7), .b(G8), .O(G275) );
nand2 gate13( .a(G9), .b(G10), .O(G278) );

  xor2  gate953(.a(G12), .b(G11), .O(gate14inter0));
  nand2 gate954(.a(gate14inter0), .b(s_58), .O(gate14inter1));
  and2  gate955(.a(G12), .b(G11), .O(gate14inter2));
  inv1  gate956(.a(s_58), .O(gate14inter3));
  inv1  gate957(.a(s_59), .O(gate14inter4));
  nand2 gate958(.a(gate14inter4), .b(gate14inter3), .O(gate14inter5));
  nor2  gate959(.a(gate14inter5), .b(gate14inter2), .O(gate14inter6));
  inv1  gate960(.a(G11), .O(gate14inter7));
  inv1  gate961(.a(G12), .O(gate14inter8));
  nand2 gate962(.a(gate14inter8), .b(gate14inter7), .O(gate14inter9));
  nand2 gate963(.a(s_59), .b(gate14inter3), .O(gate14inter10));
  nor2  gate964(.a(gate14inter10), .b(gate14inter9), .O(gate14inter11));
  nor2  gate965(.a(gate14inter11), .b(gate14inter6), .O(gate14inter12));
  nand2 gate966(.a(gate14inter12), .b(gate14inter1), .O(G281));

  xor2  gate2325(.a(G14), .b(G13), .O(gate15inter0));
  nand2 gate2326(.a(gate15inter0), .b(s_254), .O(gate15inter1));
  and2  gate2327(.a(G14), .b(G13), .O(gate15inter2));
  inv1  gate2328(.a(s_254), .O(gate15inter3));
  inv1  gate2329(.a(s_255), .O(gate15inter4));
  nand2 gate2330(.a(gate15inter4), .b(gate15inter3), .O(gate15inter5));
  nor2  gate2331(.a(gate15inter5), .b(gate15inter2), .O(gate15inter6));
  inv1  gate2332(.a(G13), .O(gate15inter7));
  inv1  gate2333(.a(G14), .O(gate15inter8));
  nand2 gate2334(.a(gate15inter8), .b(gate15inter7), .O(gate15inter9));
  nand2 gate2335(.a(s_255), .b(gate15inter3), .O(gate15inter10));
  nor2  gate2336(.a(gate15inter10), .b(gate15inter9), .O(gate15inter11));
  nor2  gate2337(.a(gate15inter11), .b(gate15inter6), .O(gate15inter12));
  nand2 gate2338(.a(gate15inter12), .b(gate15inter1), .O(G284));
nand2 gate16( .a(G15), .b(G16), .O(G287) );
nand2 gate17( .a(G17), .b(G18), .O(G290) );

  xor2  gate1051(.a(G20), .b(G19), .O(gate18inter0));
  nand2 gate1052(.a(gate18inter0), .b(s_72), .O(gate18inter1));
  and2  gate1053(.a(G20), .b(G19), .O(gate18inter2));
  inv1  gate1054(.a(s_72), .O(gate18inter3));
  inv1  gate1055(.a(s_73), .O(gate18inter4));
  nand2 gate1056(.a(gate18inter4), .b(gate18inter3), .O(gate18inter5));
  nor2  gate1057(.a(gate18inter5), .b(gate18inter2), .O(gate18inter6));
  inv1  gate1058(.a(G19), .O(gate18inter7));
  inv1  gate1059(.a(G20), .O(gate18inter8));
  nand2 gate1060(.a(gate18inter8), .b(gate18inter7), .O(gate18inter9));
  nand2 gate1061(.a(s_73), .b(gate18inter3), .O(gate18inter10));
  nor2  gate1062(.a(gate18inter10), .b(gate18inter9), .O(gate18inter11));
  nor2  gate1063(.a(gate18inter11), .b(gate18inter6), .O(gate18inter12));
  nand2 gate1064(.a(gate18inter12), .b(gate18inter1), .O(G293));

  xor2  gate1877(.a(G22), .b(G21), .O(gate19inter0));
  nand2 gate1878(.a(gate19inter0), .b(s_190), .O(gate19inter1));
  and2  gate1879(.a(G22), .b(G21), .O(gate19inter2));
  inv1  gate1880(.a(s_190), .O(gate19inter3));
  inv1  gate1881(.a(s_191), .O(gate19inter4));
  nand2 gate1882(.a(gate19inter4), .b(gate19inter3), .O(gate19inter5));
  nor2  gate1883(.a(gate19inter5), .b(gate19inter2), .O(gate19inter6));
  inv1  gate1884(.a(G21), .O(gate19inter7));
  inv1  gate1885(.a(G22), .O(gate19inter8));
  nand2 gate1886(.a(gate19inter8), .b(gate19inter7), .O(gate19inter9));
  nand2 gate1887(.a(s_191), .b(gate19inter3), .O(gate19inter10));
  nor2  gate1888(.a(gate19inter10), .b(gate19inter9), .O(gate19inter11));
  nor2  gate1889(.a(gate19inter11), .b(gate19inter6), .O(gate19inter12));
  nand2 gate1890(.a(gate19inter12), .b(gate19inter1), .O(G296));
nand2 gate20( .a(G23), .b(G24), .O(G299) );

  xor2  gate1723(.a(G26), .b(G25), .O(gate21inter0));
  nand2 gate1724(.a(gate21inter0), .b(s_168), .O(gate21inter1));
  and2  gate1725(.a(G26), .b(G25), .O(gate21inter2));
  inv1  gate1726(.a(s_168), .O(gate21inter3));
  inv1  gate1727(.a(s_169), .O(gate21inter4));
  nand2 gate1728(.a(gate21inter4), .b(gate21inter3), .O(gate21inter5));
  nor2  gate1729(.a(gate21inter5), .b(gate21inter2), .O(gate21inter6));
  inv1  gate1730(.a(G25), .O(gate21inter7));
  inv1  gate1731(.a(G26), .O(gate21inter8));
  nand2 gate1732(.a(gate21inter8), .b(gate21inter7), .O(gate21inter9));
  nand2 gate1733(.a(s_169), .b(gate21inter3), .O(gate21inter10));
  nor2  gate1734(.a(gate21inter10), .b(gate21inter9), .O(gate21inter11));
  nor2  gate1735(.a(gate21inter11), .b(gate21inter6), .O(gate21inter12));
  nand2 gate1736(.a(gate21inter12), .b(gate21inter1), .O(G302));
nand2 gate22( .a(G27), .b(G28), .O(G305) );
nand2 gate23( .a(G29), .b(G30), .O(G308) );

  xor2  gate2339(.a(G32), .b(G31), .O(gate24inter0));
  nand2 gate2340(.a(gate24inter0), .b(s_256), .O(gate24inter1));
  and2  gate2341(.a(G32), .b(G31), .O(gate24inter2));
  inv1  gate2342(.a(s_256), .O(gate24inter3));
  inv1  gate2343(.a(s_257), .O(gate24inter4));
  nand2 gate2344(.a(gate24inter4), .b(gate24inter3), .O(gate24inter5));
  nor2  gate2345(.a(gate24inter5), .b(gate24inter2), .O(gate24inter6));
  inv1  gate2346(.a(G31), .O(gate24inter7));
  inv1  gate2347(.a(G32), .O(gate24inter8));
  nand2 gate2348(.a(gate24inter8), .b(gate24inter7), .O(gate24inter9));
  nand2 gate2349(.a(s_257), .b(gate24inter3), .O(gate24inter10));
  nor2  gate2350(.a(gate24inter10), .b(gate24inter9), .O(gate24inter11));
  nor2  gate2351(.a(gate24inter11), .b(gate24inter6), .O(gate24inter12));
  nand2 gate2352(.a(gate24inter12), .b(gate24inter1), .O(G311));

  xor2  gate1639(.a(G5), .b(G1), .O(gate25inter0));
  nand2 gate1640(.a(gate25inter0), .b(s_156), .O(gate25inter1));
  and2  gate1641(.a(G5), .b(G1), .O(gate25inter2));
  inv1  gate1642(.a(s_156), .O(gate25inter3));
  inv1  gate1643(.a(s_157), .O(gate25inter4));
  nand2 gate1644(.a(gate25inter4), .b(gate25inter3), .O(gate25inter5));
  nor2  gate1645(.a(gate25inter5), .b(gate25inter2), .O(gate25inter6));
  inv1  gate1646(.a(G1), .O(gate25inter7));
  inv1  gate1647(.a(G5), .O(gate25inter8));
  nand2 gate1648(.a(gate25inter8), .b(gate25inter7), .O(gate25inter9));
  nand2 gate1649(.a(s_157), .b(gate25inter3), .O(gate25inter10));
  nor2  gate1650(.a(gate25inter10), .b(gate25inter9), .O(gate25inter11));
  nor2  gate1651(.a(gate25inter11), .b(gate25inter6), .O(gate25inter12));
  nand2 gate1652(.a(gate25inter12), .b(gate25inter1), .O(G314));
nand2 gate26( .a(G9), .b(G13), .O(G317) );

  xor2  gate2213(.a(G6), .b(G2), .O(gate27inter0));
  nand2 gate2214(.a(gate27inter0), .b(s_238), .O(gate27inter1));
  and2  gate2215(.a(G6), .b(G2), .O(gate27inter2));
  inv1  gate2216(.a(s_238), .O(gate27inter3));
  inv1  gate2217(.a(s_239), .O(gate27inter4));
  nand2 gate2218(.a(gate27inter4), .b(gate27inter3), .O(gate27inter5));
  nor2  gate2219(.a(gate27inter5), .b(gate27inter2), .O(gate27inter6));
  inv1  gate2220(.a(G2), .O(gate27inter7));
  inv1  gate2221(.a(G6), .O(gate27inter8));
  nand2 gate2222(.a(gate27inter8), .b(gate27inter7), .O(gate27inter9));
  nand2 gate2223(.a(s_239), .b(gate27inter3), .O(gate27inter10));
  nor2  gate2224(.a(gate27inter10), .b(gate27inter9), .O(gate27inter11));
  nor2  gate2225(.a(gate27inter11), .b(gate27inter6), .O(gate27inter12));
  nand2 gate2226(.a(gate27inter12), .b(gate27inter1), .O(G320));

  xor2  gate1541(.a(G14), .b(G10), .O(gate28inter0));
  nand2 gate1542(.a(gate28inter0), .b(s_142), .O(gate28inter1));
  and2  gate1543(.a(G14), .b(G10), .O(gate28inter2));
  inv1  gate1544(.a(s_142), .O(gate28inter3));
  inv1  gate1545(.a(s_143), .O(gate28inter4));
  nand2 gate1546(.a(gate28inter4), .b(gate28inter3), .O(gate28inter5));
  nor2  gate1547(.a(gate28inter5), .b(gate28inter2), .O(gate28inter6));
  inv1  gate1548(.a(G10), .O(gate28inter7));
  inv1  gate1549(.a(G14), .O(gate28inter8));
  nand2 gate1550(.a(gate28inter8), .b(gate28inter7), .O(gate28inter9));
  nand2 gate1551(.a(s_143), .b(gate28inter3), .O(gate28inter10));
  nor2  gate1552(.a(gate28inter10), .b(gate28inter9), .O(gate28inter11));
  nor2  gate1553(.a(gate28inter11), .b(gate28inter6), .O(gate28inter12));
  nand2 gate1554(.a(gate28inter12), .b(gate28inter1), .O(G323));

  xor2  gate1149(.a(G7), .b(G3), .O(gate29inter0));
  nand2 gate1150(.a(gate29inter0), .b(s_86), .O(gate29inter1));
  and2  gate1151(.a(G7), .b(G3), .O(gate29inter2));
  inv1  gate1152(.a(s_86), .O(gate29inter3));
  inv1  gate1153(.a(s_87), .O(gate29inter4));
  nand2 gate1154(.a(gate29inter4), .b(gate29inter3), .O(gate29inter5));
  nor2  gate1155(.a(gate29inter5), .b(gate29inter2), .O(gate29inter6));
  inv1  gate1156(.a(G3), .O(gate29inter7));
  inv1  gate1157(.a(G7), .O(gate29inter8));
  nand2 gate1158(.a(gate29inter8), .b(gate29inter7), .O(gate29inter9));
  nand2 gate1159(.a(s_87), .b(gate29inter3), .O(gate29inter10));
  nor2  gate1160(.a(gate29inter10), .b(gate29inter9), .O(gate29inter11));
  nor2  gate1161(.a(gate29inter11), .b(gate29inter6), .O(gate29inter12));
  nand2 gate1162(.a(gate29inter12), .b(gate29inter1), .O(G326));
nand2 gate30( .a(G11), .b(G15), .O(G329) );

  xor2  gate813(.a(G8), .b(G4), .O(gate31inter0));
  nand2 gate814(.a(gate31inter0), .b(s_38), .O(gate31inter1));
  and2  gate815(.a(G8), .b(G4), .O(gate31inter2));
  inv1  gate816(.a(s_38), .O(gate31inter3));
  inv1  gate817(.a(s_39), .O(gate31inter4));
  nand2 gate818(.a(gate31inter4), .b(gate31inter3), .O(gate31inter5));
  nor2  gate819(.a(gate31inter5), .b(gate31inter2), .O(gate31inter6));
  inv1  gate820(.a(G4), .O(gate31inter7));
  inv1  gate821(.a(G8), .O(gate31inter8));
  nand2 gate822(.a(gate31inter8), .b(gate31inter7), .O(gate31inter9));
  nand2 gate823(.a(s_39), .b(gate31inter3), .O(gate31inter10));
  nor2  gate824(.a(gate31inter10), .b(gate31inter9), .O(gate31inter11));
  nor2  gate825(.a(gate31inter11), .b(gate31inter6), .O(gate31inter12));
  nand2 gate826(.a(gate31inter12), .b(gate31inter1), .O(G332));
nand2 gate32( .a(G12), .b(G16), .O(G335) );
nand2 gate33( .a(G17), .b(G21), .O(G338) );
nand2 gate34( .a(G25), .b(G29), .O(G341) );
nand2 gate35( .a(G18), .b(G22), .O(G344) );
nand2 gate36( .a(G26), .b(G30), .O(G347) );

  xor2  gate1261(.a(G23), .b(G19), .O(gate37inter0));
  nand2 gate1262(.a(gate37inter0), .b(s_102), .O(gate37inter1));
  and2  gate1263(.a(G23), .b(G19), .O(gate37inter2));
  inv1  gate1264(.a(s_102), .O(gate37inter3));
  inv1  gate1265(.a(s_103), .O(gate37inter4));
  nand2 gate1266(.a(gate37inter4), .b(gate37inter3), .O(gate37inter5));
  nor2  gate1267(.a(gate37inter5), .b(gate37inter2), .O(gate37inter6));
  inv1  gate1268(.a(G19), .O(gate37inter7));
  inv1  gate1269(.a(G23), .O(gate37inter8));
  nand2 gate1270(.a(gate37inter8), .b(gate37inter7), .O(gate37inter9));
  nand2 gate1271(.a(s_103), .b(gate37inter3), .O(gate37inter10));
  nor2  gate1272(.a(gate37inter10), .b(gate37inter9), .O(gate37inter11));
  nor2  gate1273(.a(gate37inter11), .b(gate37inter6), .O(gate37inter12));
  nand2 gate1274(.a(gate37inter12), .b(gate37inter1), .O(G350));

  xor2  gate869(.a(G31), .b(G27), .O(gate38inter0));
  nand2 gate870(.a(gate38inter0), .b(s_46), .O(gate38inter1));
  and2  gate871(.a(G31), .b(G27), .O(gate38inter2));
  inv1  gate872(.a(s_46), .O(gate38inter3));
  inv1  gate873(.a(s_47), .O(gate38inter4));
  nand2 gate874(.a(gate38inter4), .b(gate38inter3), .O(gate38inter5));
  nor2  gate875(.a(gate38inter5), .b(gate38inter2), .O(gate38inter6));
  inv1  gate876(.a(G27), .O(gate38inter7));
  inv1  gate877(.a(G31), .O(gate38inter8));
  nand2 gate878(.a(gate38inter8), .b(gate38inter7), .O(gate38inter9));
  nand2 gate879(.a(s_47), .b(gate38inter3), .O(gate38inter10));
  nor2  gate880(.a(gate38inter10), .b(gate38inter9), .O(gate38inter11));
  nor2  gate881(.a(gate38inter11), .b(gate38inter6), .O(gate38inter12));
  nand2 gate882(.a(gate38inter12), .b(gate38inter1), .O(G353));

  xor2  gate2353(.a(G24), .b(G20), .O(gate39inter0));
  nand2 gate2354(.a(gate39inter0), .b(s_258), .O(gate39inter1));
  and2  gate2355(.a(G24), .b(G20), .O(gate39inter2));
  inv1  gate2356(.a(s_258), .O(gate39inter3));
  inv1  gate2357(.a(s_259), .O(gate39inter4));
  nand2 gate2358(.a(gate39inter4), .b(gate39inter3), .O(gate39inter5));
  nor2  gate2359(.a(gate39inter5), .b(gate39inter2), .O(gate39inter6));
  inv1  gate2360(.a(G20), .O(gate39inter7));
  inv1  gate2361(.a(G24), .O(gate39inter8));
  nand2 gate2362(.a(gate39inter8), .b(gate39inter7), .O(gate39inter9));
  nand2 gate2363(.a(s_259), .b(gate39inter3), .O(gate39inter10));
  nor2  gate2364(.a(gate39inter10), .b(gate39inter9), .O(gate39inter11));
  nor2  gate2365(.a(gate39inter11), .b(gate39inter6), .O(gate39inter12));
  nand2 gate2366(.a(gate39inter12), .b(gate39inter1), .O(G356));
nand2 gate40( .a(G28), .b(G32), .O(G359) );
nand2 gate41( .a(G1), .b(G266), .O(G362) );
nand2 gate42( .a(G2), .b(G266), .O(G363) );
nand2 gate43( .a(G3), .b(G269), .O(G364) );
nand2 gate44( .a(G4), .b(G269), .O(G365) );
nand2 gate45( .a(G5), .b(G272), .O(G366) );
nand2 gate46( .a(G6), .b(G272), .O(G367) );

  xor2  gate2297(.a(G275), .b(G7), .O(gate47inter0));
  nand2 gate2298(.a(gate47inter0), .b(s_250), .O(gate47inter1));
  and2  gate2299(.a(G275), .b(G7), .O(gate47inter2));
  inv1  gate2300(.a(s_250), .O(gate47inter3));
  inv1  gate2301(.a(s_251), .O(gate47inter4));
  nand2 gate2302(.a(gate47inter4), .b(gate47inter3), .O(gate47inter5));
  nor2  gate2303(.a(gate47inter5), .b(gate47inter2), .O(gate47inter6));
  inv1  gate2304(.a(G7), .O(gate47inter7));
  inv1  gate2305(.a(G275), .O(gate47inter8));
  nand2 gate2306(.a(gate47inter8), .b(gate47inter7), .O(gate47inter9));
  nand2 gate2307(.a(s_251), .b(gate47inter3), .O(gate47inter10));
  nor2  gate2308(.a(gate47inter10), .b(gate47inter9), .O(gate47inter11));
  nor2  gate2309(.a(gate47inter11), .b(gate47inter6), .O(gate47inter12));
  nand2 gate2310(.a(gate47inter12), .b(gate47inter1), .O(G368));
nand2 gate48( .a(G8), .b(G275), .O(G369) );

  xor2  gate1009(.a(G278), .b(G9), .O(gate49inter0));
  nand2 gate1010(.a(gate49inter0), .b(s_66), .O(gate49inter1));
  and2  gate1011(.a(G278), .b(G9), .O(gate49inter2));
  inv1  gate1012(.a(s_66), .O(gate49inter3));
  inv1  gate1013(.a(s_67), .O(gate49inter4));
  nand2 gate1014(.a(gate49inter4), .b(gate49inter3), .O(gate49inter5));
  nor2  gate1015(.a(gate49inter5), .b(gate49inter2), .O(gate49inter6));
  inv1  gate1016(.a(G9), .O(gate49inter7));
  inv1  gate1017(.a(G278), .O(gate49inter8));
  nand2 gate1018(.a(gate49inter8), .b(gate49inter7), .O(gate49inter9));
  nand2 gate1019(.a(s_67), .b(gate49inter3), .O(gate49inter10));
  nor2  gate1020(.a(gate49inter10), .b(gate49inter9), .O(gate49inter11));
  nor2  gate1021(.a(gate49inter11), .b(gate49inter6), .O(gate49inter12));
  nand2 gate1022(.a(gate49inter12), .b(gate49inter1), .O(G370));
nand2 gate50( .a(G10), .b(G278), .O(G371) );

  xor2  gate1989(.a(G281), .b(G11), .O(gate51inter0));
  nand2 gate1990(.a(gate51inter0), .b(s_206), .O(gate51inter1));
  and2  gate1991(.a(G281), .b(G11), .O(gate51inter2));
  inv1  gate1992(.a(s_206), .O(gate51inter3));
  inv1  gate1993(.a(s_207), .O(gate51inter4));
  nand2 gate1994(.a(gate51inter4), .b(gate51inter3), .O(gate51inter5));
  nor2  gate1995(.a(gate51inter5), .b(gate51inter2), .O(gate51inter6));
  inv1  gate1996(.a(G11), .O(gate51inter7));
  inv1  gate1997(.a(G281), .O(gate51inter8));
  nand2 gate1998(.a(gate51inter8), .b(gate51inter7), .O(gate51inter9));
  nand2 gate1999(.a(s_207), .b(gate51inter3), .O(gate51inter10));
  nor2  gate2000(.a(gate51inter10), .b(gate51inter9), .O(gate51inter11));
  nor2  gate2001(.a(gate51inter11), .b(gate51inter6), .O(gate51inter12));
  nand2 gate2002(.a(gate51inter12), .b(gate51inter1), .O(G372));

  xor2  gate1023(.a(G281), .b(G12), .O(gate52inter0));
  nand2 gate1024(.a(gate52inter0), .b(s_68), .O(gate52inter1));
  and2  gate1025(.a(G281), .b(G12), .O(gate52inter2));
  inv1  gate1026(.a(s_68), .O(gate52inter3));
  inv1  gate1027(.a(s_69), .O(gate52inter4));
  nand2 gate1028(.a(gate52inter4), .b(gate52inter3), .O(gate52inter5));
  nor2  gate1029(.a(gate52inter5), .b(gate52inter2), .O(gate52inter6));
  inv1  gate1030(.a(G12), .O(gate52inter7));
  inv1  gate1031(.a(G281), .O(gate52inter8));
  nand2 gate1032(.a(gate52inter8), .b(gate52inter7), .O(gate52inter9));
  nand2 gate1033(.a(s_69), .b(gate52inter3), .O(gate52inter10));
  nor2  gate1034(.a(gate52inter10), .b(gate52inter9), .O(gate52inter11));
  nor2  gate1035(.a(gate52inter11), .b(gate52inter6), .O(gate52inter12));
  nand2 gate1036(.a(gate52inter12), .b(gate52inter1), .O(G373));
nand2 gate53( .a(G13), .b(G284), .O(G374) );

  xor2  gate659(.a(G284), .b(G14), .O(gate54inter0));
  nand2 gate660(.a(gate54inter0), .b(s_16), .O(gate54inter1));
  and2  gate661(.a(G284), .b(G14), .O(gate54inter2));
  inv1  gate662(.a(s_16), .O(gate54inter3));
  inv1  gate663(.a(s_17), .O(gate54inter4));
  nand2 gate664(.a(gate54inter4), .b(gate54inter3), .O(gate54inter5));
  nor2  gate665(.a(gate54inter5), .b(gate54inter2), .O(gate54inter6));
  inv1  gate666(.a(G14), .O(gate54inter7));
  inv1  gate667(.a(G284), .O(gate54inter8));
  nand2 gate668(.a(gate54inter8), .b(gate54inter7), .O(gate54inter9));
  nand2 gate669(.a(s_17), .b(gate54inter3), .O(gate54inter10));
  nor2  gate670(.a(gate54inter10), .b(gate54inter9), .O(gate54inter11));
  nor2  gate671(.a(gate54inter11), .b(gate54inter6), .O(gate54inter12));
  nand2 gate672(.a(gate54inter12), .b(gate54inter1), .O(G375));
nand2 gate55( .a(G15), .b(G287), .O(G376) );

  xor2  gate1485(.a(G287), .b(G16), .O(gate56inter0));
  nand2 gate1486(.a(gate56inter0), .b(s_134), .O(gate56inter1));
  and2  gate1487(.a(G287), .b(G16), .O(gate56inter2));
  inv1  gate1488(.a(s_134), .O(gate56inter3));
  inv1  gate1489(.a(s_135), .O(gate56inter4));
  nand2 gate1490(.a(gate56inter4), .b(gate56inter3), .O(gate56inter5));
  nor2  gate1491(.a(gate56inter5), .b(gate56inter2), .O(gate56inter6));
  inv1  gate1492(.a(G16), .O(gate56inter7));
  inv1  gate1493(.a(G287), .O(gate56inter8));
  nand2 gate1494(.a(gate56inter8), .b(gate56inter7), .O(gate56inter9));
  nand2 gate1495(.a(s_135), .b(gate56inter3), .O(gate56inter10));
  nor2  gate1496(.a(gate56inter10), .b(gate56inter9), .O(gate56inter11));
  nor2  gate1497(.a(gate56inter11), .b(gate56inter6), .O(gate56inter12));
  nand2 gate1498(.a(gate56inter12), .b(gate56inter1), .O(G377));
nand2 gate57( .a(G17), .b(G290), .O(G378) );
nand2 gate58( .a(G18), .b(G290), .O(G379) );
nand2 gate59( .a(G19), .b(G293), .O(G380) );
nand2 gate60( .a(G20), .b(G293), .O(G381) );

  xor2  gate1933(.a(G296), .b(G21), .O(gate61inter0));
  nand2 gate1934(.a(gate61inter0), .b(s_198), .O(gate61inter1));
  and2  gate1935(.a(G296), .b(G21), .O(gate61inter2));
  inv1  gate1936(.a(s_198), .O(gate61inter3));
  inv1  gate1937(.a(s_199), .O(gate61inter4));
  nand2 gate1938(.a(gate61inter4), .b(gate61inter3), .O(gate61inter5));
  nor2  gate1939(.a(gate61inter5), .b(gate61inter2), .O(gate61inter6));
  inv1  gate1940(.a(G21), .O(gate61inter7));
  inv1  gate1941(.a(G296), .O(gate61inter8));
  nand2 gate1942(.a(gate61inter8), .b(gate61inter7), .O(gate61inter9));
  nand2 gate1943(.a(s_199), .b(gate61inter3), .O(gate61inter10));
  nor2  gate1944(.a(gate61inter10), .b(gate61inter9), .O(gate61inter11));
  nor2  gate1945(.a(gate61inter11), .b(gate61inter6), .O(gate61inter12));
  nand2 gate1946(.a(gate61inter12), .b(gate61inter1), .O(G382));

  xor2  gate1177(.a(G296), .b(G22), .O(gate62inter0));
  nand2 gate1178(.a(gate62inter0), .b(s_90), .O(gate62inter1));
  and2  gate1179(.a(G296), .b(G22), .O(gate62inter2));
  inv1  gate1180(.a(s_90), .O(gate62inter3));
  inv1  gate1181(.a(s_91), .O(gate62inter4));
  nand2 gate1182(.a(gate62inter4), .b(gate62inter3), .O(gate62inter5));
  nor2  gate1183(.a(gate62inter5), .b(gate62inter2), .O(gate62inter6));
  inv1  gate1184(.a(G22), .O(gate62inter7));
  inv1  gate1185(.a(G296), .O(gate62inter8));
  nand2 gate1186(.a(gate62inter8), .b(gate62inter7), .O(gate62inter9));
  nand2 gate1187(.a(s_91), .b(gate62inter3), .O(gate62inter10));
  nor2  gate1188(.a(gate62inter10), .b(gate62inter9), .O(gate62inter11));
  nor2  gate1189(.a(gate62inter11), .b(gate62inter6), .O(gate62inter12));
  nand2 gate1190(.a(gate62inter12), .b(gate62inter1), .O(G383));

  xor2  gate603(.a(G299), .b(G23), .O(gate63inter0));
  nand2 gate604(.a(gate63inter0), .b(s_8), .O(gate63inter1));
  and2  gate605(.a(G299), .b(G23), .O(gate63inter2));
  inv1  gate606(.a(s_8), .O(gate63inter3));
  inv1  gate607(.a(s_9), .O(gate63inter4));
  nand2 gate608(.a(gate63inter4), .b(gate63inter3), .O(gate63inter5));
  nor2  gate609(.a(gate63inter5), .b(gate63inter2), .O(gate63inter6));
  inv1  gate610(.a(G23), .O(gate63inter7));
  inv1  gate611(.a(G299), .O(gate63inter8));
  nand2 gate612(.a(gate63inter8), .b(gate63inter7), .O(gate63inter9));
  nand2 gate613(.a(s_9), .b(gate63inter3), .O(gate63inter10));
  nor2  gate614(.a(gate63inter10), .b(gate63inter9), .O(gate63inter11));
  nor2  gate615(.a(gate63inter11), .b(gate63inter6), .O(gate63inter12));
  nand2 gate616(.a(gate63inter12), .b(gate63inter1), .O(G384));
nand2 gate64( .a(G24), .b(G299), .O(G385) );
nand2 gate65( .a(G25), .b(G302), .O(G386) );
nand2 gate66( .a(G26), .b(G302), .O(G387) );
nand2 gate67( .a(G27), .b(G305), .O(G388) );
nand2 gate68( .a(G28), .b(G305), .O(G389) );
nand2 gate69( .a(G29), .b(G308), .O(G390) );
nand2 gate70( .a(G30), .b(G308), .O(G391) );
nand2 gate71( .a(G31), .b(G311), .O(G392) );
nand2 gate72( .a(G32), .b(G311), .O(G393) );
nand2 gate73( .a(G1), .b(G314), .O(G394) );
nand2 gate74( .a(G5), .b(G314), .O(G395) );
nand2 gate75( .a(G9), .b(G317), .O(G396) );
nand2 gate76( .a(G13), .b(G317), .O(G397) );
nand2 gate77( .a(G2), .b(G320), .O(G398) );

  xor2  gate1163(.a(G320), .b(G6), .O(gate78inter0));
  nand2 gate1164(.a(gate78inter0), .b(s_88), .O(gate78inter1));
  and2  gate1165(.a(G320), .b(G6), .O(gate78inter2));
  inv1  gate1166(.a(s_88), .O(gate78inter3));
  inv1  gate1167(.a(s_89), .O(gate78inter4));
  nand2 gate1168(.a(gate78inter4), .b(gate78inter3), .O(gate78inter5));
  nor2  gate1169(.a(gate78inter5), .b(gate78inter2), .O(gate78inter6));
  inv1  gate1170(.a(G6), .O(gate78inter7));
  inv1  gate1171(.a(G320), .O(gate78inter8));
  nand2 gate1172(.a(gate78inter8), .b(gate78inter7), .O(gate78inter9));
  nand2 gate1173(.a(s_89), .b(gate78inter3), .O(gate78inter10));
  nor2  gate1174(.a(gate78inter10), .b(gate78inter9), .O(gate78inter11));
  nor2  gate1175(.a(gate78inter11), .b(gate78inter6), .O(gate78inter12));
  nand2 gate1176(.a(gate78inter12), .b(gate78inter1), .O(G399));
nand2 gate79( .a(G10), .b(G323), .O(G400) );

  xor2  gate1975(.a(G323), .b(G14), .O(gate80inter0));
  nand2 gate1976(.a(gate80inter0), .b(s_204), .O(gate80inter1));
  and2  gate1977(.a(G323), .b(G14), .O(gate80inter2));
  inv1  gate1978(.a(s_204), .O(gate80inter3));
  inv1  gate1979(.a(s_205), .O(gate80inter4));
  nand2 gate1980(.a(gate80inter4), .b(gate80inter3), .O(gate80inter5));
  nor2  gate1981(.a(gate80inter5), .b(gate80inter2), .O(gate80inter6));
  inv1  gate1982(.a(G14), .O(gate80inter7));
  inv1  gate1983(.a(G323), .O(gate80inter8));
  nand2 gate1984(.a(gate80inter8), .b(gate80inter7), .O(gate80inter9));
  nand2 gate1985(.a(s_205), .b(gate80inter3), .O(gate80inter10));
  nor2  gate1986(.a(gate80inter10), .b(gate80inter9), .O(gate80inter11));
  nor2  gate1987(.a(gate80inter11), .b(gate80inter6), .O(gate80inter12));
  nand2 gate1988(.a(gate80inter12), .b(gate80inter1), .O(G401));
nand2 gate81( .a(G3), .b(G326), .O(G402) );
nand2 gate82( .a(G7), .b(G326), .O(G403) );
nand2 gate83( .a(G11), .b(G329), .O(G404) );
nand2 gate84( .a(G15), .b(G329), .O(G405) );

  xor2  gate841(.a(G332), .b(G4), .O(gate85inter0));
  nand2 gate842(.a(gate85inter0), .b(s_42), .O(gate85inter1));
  and2  gate843(.a(G332), .b(G4), .O(gate85inter2));
  inv1  gate844(.a(s_42), .O(gate85inter3));
  inv1  gate845(.a(s_43), .O(gate85inter4));
  nand2 gate846(.a(gate85inter4), .b(gate85inter3), .O(gate85inter5));
  nor2  gate847(.a(gate85inter5), .b(gate85inter2), .O(gate85inter6));
  inv1  gate848(.a(G4), .O(gate85inter7));
  inv1  gate849(.a(G332), .O(gate85inter8));
  nand2 gate850(.a(gate85inter8), .b(gate85inter7), .O(gate85inter9));
  nand2 gate851(.a(s_43), .b(gate85inter3), .O(gate85inter10));
  nor2  gate852(.a(gate85inter10), .b(gate85inter9), .O(gate85inter11));
  nor2  gate853(.a(gate85inter11), .b(gate85inter6), .O(gate85inter12));
  nand2 gate854(.a(gate85inter12), .b(gate85inter1), .O(G406));
nand2 gate86( .a(G8), .b(G332), .O(G407) );

  xor2  gate967(.a(G335), .b(G12), .O(gate87inter0));
  nand2 gate968(.a(gate87inter0), .b(s_60), .O(gate87inter1));
  and2  gate969(.a(G335), .b(G12), .O(gate87inter2));
  inv1  gate970(.a(s_60), .O(gate87inter3));
  inv1  gate971(.a(s_61), .O(gate87inter4));
  nand2 gate972(.a(gate87inter4), .b(gate87inter3), .O(gate87inter5));
  nor2  gate973(.a(gate87inter5), .b(gate87inter2), .O(gate87inter6));
  inv1  gate974(.a(G12), .O(gate87inter7));
  inv1  gate975(.a(G335), .O(gate87inter8));
  nand2 gate976(.a(gate87inter8), .b(gate87inter7), .O(gate87inter9));
  nand2 gate977(.a(s_61), .b(gate87inter3), .O(gate87inter10));
  nor2  gate978(.a(gate87inter10), .b(gate87inter9), .O(gate87inter11));
  nor2  gate979(.a(gate87inter11), .b(gate87inter6), .O(gate87inter12));
  nand2 gate980(.a(gate87inter12), .b(gate87inter1), .O(G408));
nand2 gate88( .a(G16), .b(G335), .O(G409) );
nand2 gate89( .a(G17), .b(G338), .O(G410) );
nand2 gate90( .a(G21), .b(G338), .O(G411) );

  xor2  gate1373(.a(G341), .b(G25), .O(gate91inter0));
  nand2 gate1374(.a(gate91inter0), .b(s_118), .O(gate91inter1));
  and2  gate1375(.a(G341), .b(G25), .O(gate91inter2));
  inv1  gate1376(.a(s_118), .O(gate91inter3));
  inv1  gate1377(.a(s_119), .O(gate91inter4));
  nand2 gate1378(.a(gate91inter4), .b(gate91inter3), .O(gate91inter5));
  nor2  gate1379(.a(gate91inter5), .b(gate91inter2), .O(gate91inter6));
  inv1  gate1380(.a(G25), .O(gate91inter7));
  inv1  gate1381(.a(G341), .O(gate91inter8));
  nand2 gate1382(.a(gate91inter8), .b(gate91inter7), .O(gate91inter9));
  nand2 gate1383(.a(s_119), .b(gate91inter3), .O(gate91inter10));
  nor2  gate1384(.a(gate91inter10), .b(gate91inter9), .O(gate91inter11));
  nor2  gate1385(.a(gate91inter11), .b(gate91inter6), .O(gate91inter12));
  nand2 gate1386(.a(gate91inter12), .b(gate91inter1), .O(G412));

  xor2  gate1653(.a(G341), .b(G29), .O(gate92inter0));
  nand2 gate1654(.a(gate92inter0), .b(s_158), .O(gate92inter1));
  and2  gate1655(.a(G341), .b(G29), .O(gate92inter2));
  inv1  gate1656(.a(s_158), .O(gate92inter3));
  inv1  gate1657(.a(s_159), .O(gate92inter4));
  nand2 gate1658(.a(gate92inter4), .b(gate92inter3), .O(gate92inter5));
  nor2  gate1659(.a(gate92inter5), .b(gate92inter2), .O(gate92inter6));
  inv1  gate1660(.a(G29), .O(gate92inter7));
  inv1  gate1661(.a(G341), .O(gate92inter8));
  nand2 gate1662(.a(gate92inter8), .b(gate92inter7), .O(gate92inter9));
  nand2 gate1663(.a(s_159), .b(gate92inter3), .O(gate92inter10));
  nor2  gate1664(.a(gate92inter10), .b(gate92inter9), .O(gate92inter11));
  nor2  gate1665(.a(gate92inter11), .b(gate92inter6), .O(gate92inter12));
  nand2 gate1666(.a(gate92inter12), .b(gate92inter1), .O(G413));
nand2 gate93( .a(G18), .b(G344), .O(G414) );
nand2 gate94( .a(G22), .b(G344), .O(G415) );
nand2 gate95( .a(G26), .b(G347), .O(G416) );

  xor2  gate1807(.a(G347), .b(G30), .O(gate96inter0));
  nand2 gate1808(.a(gate96inter0), .b(s_180), .O(gate96inter1));
  and2  gate1809(.a(G347), .b(G30), .O(gate96inter2));
  inv1  gate1810(.a(s_180), .O(gate96inter3));
  inv1  gate1811(.a(s_181), .O(gate96inter4));
  nand2 gate1812(.a(gate96inter4), .b(gate96inter3), .O(gate96inter5));
  nor2  gate1813(.a(gate96inter5), .b(gate96inter2), .O(gate96inter6));
  inv1  gate1814(.a(G30), .O(gate96inter7));
  inv1  gate1815(.a(G347), .O(gate96inter8));
  nand2 gate1816(.a(gate96inter8), .b(gate96inter7), .O(gate96inter9));
  nand2 gate1817(.a(s_181), .b(gate96inter3), .O(gate96inter10));
  nor2  gate1818(.a(gate96inter10), .b(gate96inter9), .O(gate96inter11));
  nor2  gate1819(.a(gate96inter11), .b(gate96inter6), .O(gate96inter12));
  nand2 gate1820(.a(gate96inter12), .b(gate96inter1), .O(G417));
nand2 gate97( .a(G19), .b(G350), .O(G418) );
nand2 gate98( .a(G23), .b(G350), .O(G419) );
nand2 gate99( .a(G27), .b(G353), .O(G420) );
nand2 gate100( .a(G31), .b(G353), .O(G421) );
nand2 gate101( .a(G20), .b(G356), .O(G422) );

  xor2  gate1891(.a(G356), .b(G24), .O(gate102inter0));
  nand2 gate1892(.a(gate102inter0), .b(s_192), .O(gate102inter1));
  and2  gate1893(.a(G356), .b(G24), .O(gate102inter2));
  inv1  gate1894(.a(s_192), .O(gate102inter3));
  inv1  gate1895(.a(s_193), .O(gate102inter4));
  nand2 gate1896(.a(gate102inter4), .b(gate102inter3), .O(gate102inter5));
  nor2  gate1897(.a(gate102inter5), .b(gate102inter2), .O(gate102inter6));
  inv1  gate1898(.a(G24), .O(gate102inter7));
  inv1  gate1899(.a(G356), .O(gate102inter8));
  nand2 gate1900(.a(gate102inter8), .b(gate102inter7), .O(gate102inter9));
  nand2 gate1901(.a(s_193), .b(gate102inter3), .O(gate102inter10));
  nor2  gate1902(.a(gate102inter10), .b(gate102inter9), .O(gate102inter11));
  nor2  gate1903(.a(gate102inter11), .b(gate102inter6), .O(gate102inter12));
  nand2 gate1904(.a(gate102inter12), .b(gate102inter1), .O(G423));
nand2 gate103( .a(G28), .b(G359), .O(G424) );
nand2 gate104( .a(G32), .b(G359), .O(G425) );

  xor2  gate1121(.a(G363), .b(G362), .O(gate105inter0));
  nand2 gate1122(.a(gate105inter0), .b(s_82), .O(gate105inter1));
  and2  gate1123(.a(G363), .b(G362), .O(gate105inter2));
  inv1  gate1124(.a(s_82), .O(gate105inter3));
  inv1  gate1125(.a(s_83), .O(gate105inter4));
  nand2 gate1126(.a(gate105inter4), .b(gate105inter3), .O(gate105inter5));
  nor2  gate1127(.a(gate105inter5), .b(gate105inter2), .O(gate105inter6));
  inv1  gate1128(.a(G362), .O(gate105inter7));
  inv1  gate1129(.a(G363), .O(gate105inter8));
  nand2 gate1130(.a(gate105inter8), .b(gate105inter7), .O(gate105inter9));
  nand2 gate1131(.a(s_83), .b(gate105inter3), .O(gate105inter10));
  nor2  gate1132(.a(gate105inter10), .b(gate105inter9), .O(gate105inter11));
  nor2  gate1133(.a(gate105inter11), .b(gate105inter6), .O(gate105inter12));
  nand2 gate1134(.a(gate105inter12), .b(gate105inter1), .O(G426));
nand2 gate106( .a(G364), .b(G365), .O(G429) );
nand2 gate107( .a(G366), .b(G367), .O(G432) );
nand2 gate108( .a(G368), .b(G369), .O(G435) );

  xor2  gate897(.a(G371), .b(G370), .O(gate109inter0));
  nand2 gate898(.a(gate109inter0), .b(s_50), .O(gate109inter1));
  and2  gate899(.a(G371), .b(G370), .O(gate109inter2));
  inv1  gate900(.a(s_50), .O(gate109inter3));
  inv1  gate901(.a(s_51), .O(gate109inter4));
  nand2 gate902(.a(gate109inter4), .b(gate109inter3), .O(gate109inter5));
  nor2  gate903(.a(gate109inter5), .b(gate109inter2), .O(gate109inter6));
  inv1  gate904(.a(G370), .O(gate109inter7));
  inv1  gate905(.a(G371), .O(gate109inter8));
  nand2 gate906(.a(gate109inter8), .b(gate109inter7), .O(gate109inter9));
  nand2 gate907(.a(s_51), .b(gate109inter3), .O(gate109inter10));
  nor2  gate908(.a(gate109inter10), .b(gate109inter9), .O(gate109inter11));
  nor2  gate909(.a(gate109inter11), .b(gate109inter6), .O(gate109inter12));
  nand2 gate910(.a(gate109inter12), .b(gate109inter1), .O(G438));
nand2 gate110( .a(G372), .b(G373), .O(G441) );
nand2 gate111( .a(G374), .b(G375), .O(G444) );
nand2 gate112( .a(G376), .b(G377), .O(G447) );
nand2 gate113( .a(G378), .b(G379), .O(G450) );
nand2 gate114( .a(G380), .b(G381), .O(G453) );
nand2 gate115( .a(G382), .b(G383), .O(G456) );
nand2 gate116( .a(G384), .b(G385), .O(G459) );
nand2 gate117( .a(G386), .b(G387), .O(G462) );

  xor2  gate1709(.a(G389), .b(G388), .O(gate118inter0));
  nand2 gate1710(.a(gate118inter0), .b(s_166), .O(gate118inter1));
  and2  gate1711(.a(G389), .b(G388), .O(gate118inter2));
  inv1  gate1712(.a(s_166), .O(gate118inter3));
  inv1  gate1713(.a(s_167), .O(gate118inter4));
  nand2 gate1714(.a(gate118inter4), .b(gate118inter3), .O(gate118inter5));
  nor2  gate1715(.a(gate118inter5), .b(gate118inter2), .O(gate118inter6));
  inv1  gate1716(.a(G388), .O(gate118inter7));
  inv1  gate1717(.a(G389), .O(gate118inter8));
  nand2 gate1718(.a(gate118inter8), .b(gate118inter7), .O(gate118inter9));
  nand2 gate1719(.a(s_167), .b(gate118inter3), .O(gate118inter10));
  nor2  gate1720(.a(gate118inter10), .b(gate118inter9), .O(gate118inter11));
  nor2  gate1721(.a(gate118inter11), .b(gate118inter6), .O(gate118inter12));
  nand2 gate1722(.a(gate118inter12), .b(gate118inter1), .O(G465));

  xor2  gate1583(.a(G391), .b(G390), .O(gate119inter0));
  nand2 gate1584(.a(gate119inter0), .b(s_148), .O(gate119inter1));
  and2  gate1585(.a(G391), .b(G390), .O(gate119inter2));
  inv1  gate1586(.a(s_148), .O(gate119inter3));
  inv1  gate1587(.a(s_149), .O(gate119inter4));
  nand2 gate1588(.a(gate119inter4), .b(gate119inter3), .O(gate119inter5));
  nor2  gate1589(.a(gate119inter5), .b(gate119inter2), .O(gate119inter6));
  inv1  gate1590(.a(G390), .O(gate119inter7));
  inv1  gate1591(.a(G391), .O(gate119inter8));
  nand2 gate1592(.a(gate119inter8), .b(gate119inter7), .O(gate119inter9));
  nand2 gate1593(.a(s_149), .b(gate119inter3), .O(gate119inter10));
  nor2  gate1594(.a(gate119inter10), .b(gate119inter9), .O(gate119inter11));
  nor2  gate1595(.a(gate119inter11), .b(gate119inter6), .O(gate119inter12));
  nand2 gate1596(.a(gate119inter12), .b(gate119inter1), .O(G468));

  xor2  gate1961(.a(G393), .b(G392), .O(gate120inter0));
  nand2 gate1962(.a(gate120inter0), .b(s_202), .O(gate120inter1));
  and2  gate1963(.a(G393), .b(G392), .O(gate120inter2));
  inv1  gate1964(.a(s_202), .O(gate120inter3));
  inv1  gate1965(.a(s_203), .O(gate120inter4));
  nand2 gate1966(.a(gate120inter4), .b(gate120inter3), .O(gate120inter5));
  nor2  gate1967(.a(gate120inter5), .b(gate120inter2), .O(gate120inter6));
  inv1  gate1968(.a(G392), .O(gate120inter7));
  inv1  gate1969(.a(G393), .O(gate120inter8));
  nand2 gate1970(.a(gate120inter8), .b(gate120inter7), .O(gate120inter9));
  nand2 gate1971(.a(s_203), .b(gate120inter3), .O(gate120inter10));
  nor2  gate1972(.a(gate120inter10), .b(gate120inter9), .O(gate120inter11));
  nor2  gate1973(.a(gate120inter11), .b(gate120inter6), .O(gate120inter12));
  nand2 gate1974(.a(gate120inter12), .b(gate120inter1), .O(G471));
nand2 gate121( .a(G394), .b(G395), .O(G474) );
nand2 gate122( .a(G396), .b(G397), .O(G477) );
nand2 gate123( .a(G398), .b(G399), .O(G480) );
nand2 gate124( .a(G400), .b(G401), .O(G483) );
nand2 gate125( .a(G402), .b(G403), .O(G486) );
nand2 gate126( .a(G404), .b(G405), .O(G489) );
nand2 gate127( .a(G406), .b(G407), .O(G492) );

  xor2  gate589(.a(G409), .b(G408), .O(gate128inter0));
  nand2 gate590(.a(gate128inter0), .b(s_6), .O(gate128inter1));
  and2  gate591(.a(G409), .b(G408), .O(gate128inter2));
  inv1  gate592(.a(s_6), .O(gate128inter3));
  inv1  gate593(.a(s_7), .O(gate128inter4));
  nand2 gate594(.a(gate128inter4), .b(gate128inter3), .O(gate128inter5));
  nor2  gate595(.a(gate128inter5), .b(gate128inter2), .O(gate128inter6));
  inv1  gate596(.a(G408), .O(gate128inter7));
  inv1  gate597(.a(G409), .O(gate128inter8));
  nand2 gate598(.a(gate128inter8), .b(gate128inter7), .O(gate128inter9));
  nand2 gate599(.a(s_7), .b(gate128inter3), .O(gate128inter10));
  nor2  gate600(.a(gate128inter10), .b(gate128inter9), .O(gate128inter11));
  nor2  gate601(.a(gate128inter11), .b(gate128inter6), .O(gate128inter12));
  nand2 gate602(.a(gate128inter12), .b(gate128inter1), .O(G495));
nand2 gate129( .a(G410), .b(G411), .O(G498) );
nand2 gate130( .a(G412), .b(G413), .O(G501) );

  xor2  gate729(.a(G415), .b(G414), .O(gate131inter0));
  nand2 gate730(.a(gate131inter0), .b(s_26), .O(gate131inter1));
  and2  gate731(.a(G415), .b(G414), .O(gate131inter2));
  inv1  gate732(.a(s_26), .O(gate131inter3));
  inv1  gate733(.a(s_27), .O(gate131inter4));
  nand2 gate734(.a(gate131inter4), .b(gate131inter3), .O(gate131inter5));
  nor2  gate735(.a(gate131inter5), .b(gate131inter2), .O(gate131inter6));
  inv1  gate736(.a(G414), .O(gate131inter7));
  inv1  gate737(.a(G415), .O(gate131inter8));
  nand2 gate738(.a(gate131inter8), .b(gate131inter7), .O(gate131inter9));
  nand2 gate739(.a(s_27), .b(gate131inter3), .O(gate131inter10));
  nor2  gate740(.a(gate131inter10), .b(gate131inter9), .O(gate131inter11));
  nor2  gate741(.a(gate131inter11), .b(gate131inter6), .O(gate131inter12));
  nand2 gate742(.a(gate131inter12), .b(gate131inter1), .O(G504));

  xor2  gate1611(.a(G417), .b(G416), .O(gate132inter0));
  nand2 gate1612(.a(gate132inter0), .b(s_152), .O(gate132inter1));
  and2  gate1613(.a(G417), .b(G416), .O(gate132inter2));
  inv1  gate1614(.a(s_152), .O(gate132inter3));
  inv1  gate1615(.a(s_153), .O(gate132inter4));
  nand2 gate1616(.a(gate132inter4), .b(gate132inter3), .O(gate132inter5));
  nor2  gate1617(.a(gate132inter5), .b(gate132inter2), .O(gate132inter6));
  inv1  gate1618(.a(G416), .O(gate132inter7));
  inv1  gate1619(.a(G417), .O(gate132inter8));
  nand2 gate1620(.a(gate132inter8), .b(gate132inter7), .O(gate132inter9));
  nand2 gate1621(.a(s_153), .b(gate132inter3), .O(gate132inter10));
  nor2  gate1622(.a(gate132inter10), .b(gate132inter9), .O(gate132inter11));
  nor2  gate1623(.a(gate132inter11), .b(gate132inter6), .O(gate132inter12));
  nand2 gate1624(.a(gate132inter12), .b(gate132inter1), .O(G507));
nand2 gate133( .a(G418), .b(G419), .O(G510) );
nand2 gate134( .a(G420), .b(G421), .O(G513) );
nand2 gate135( .a(G422), .b(G423), .O(G516) );

  xor2  gate1513(.a(G425), .b(G424), .O(gate136inter0));
  nand2 gate1514(.a(gate136inter0), .b(s_138), .O(gate136inter1));
  and2  gate1515(.a(G425), .b(G424), .O(gate136inter2));
  inv1  gate1516(.a(s_138), .O(gate136inter3));
  inv1  gate1517(.a(s_139), .O(gate136inter4));
  nand2 gate1518(.a(gate136inter4), .b(gate136inter3), .O(gate136inter5));
  nor2  gate1519(.a(gate136inter5), .b(gate136inter2), .O(gate136inter6));
  inv1  gate1520(.a(G424), .O(gate136inter7));
  inv1  gate1521(.a(G425), .O(gate136inter8));
  nand2 gate1522(.a(gate136inter8), .b(gate136inter7), .O(gate136inter9));
  nand2 gate1523(.a(s_139), .b(gate136inter3), .O(gate136inter10));
  nor2  gate1524(.a(gate136inter10), .b(gate136inter9), .O(gate136inter11));
  nor2  gate1525(.a(gate136inter11), .b(gate136inter6), .O(gate136inter12));
  nand2 gate1526(.a(gate136inter12), .b(gate136inter1), .O(G519));
nand2 gate137( .a(G426), .b(G429), .O(G522) );
nand2 gate138( .a(G432), .b(G435), .O(G525) );
nand2 gate139( .a(G438), .b(G441), .O(G528) );
nand2 gate140( .a(G444), .b(G447), .O(G531) );

  xor2  gate1359(.a(G453), .b(G450), .O(gate141inter0));
  nand2 gate1360(.a(gate141inter0), .b(s_116), .O(gate141inter1));
  and2  gate1361(.a(G453), .b(G450), .O(gate141inter2));
  inv1  gate1362(.a(s_116), .O(gate141inter3));
  inv1  gate1363(.a(s_117), .O(gate141inter4));
  nand2 gate1364(.a(gate141inter4), .b(gate141inter3), .O(gate141inter5));
  nor2  gate1365(.a(gate141inter5), .b(gate141inter2), .O(gate141inter6));
  inv1  gate1366(.a(G450), .O(gate141inter7));
  inv1  gate1367(.a(G453), .O(gate141inter8));
  nand2 gate1368(.a(gate141inter8), .b(gate141inter7), .O(gate141inter9));
  nand2 gate1369(.a(s_117), .b(gate141inter3), .O(gate141inter10));
  nor2  gate1370(.a(gate141inter10), .b(gate141inter9), .O(gate141inter11));
  nor2  gate1371(.a(gate141inter11), .b(gate141inter6), .O(gate141inter12));
  nand2 gate1372(.a(gate141inter12), .b(gate141inter1), .O(G534));
nand2 gate142( .a(G456), .b(G459), .O(G537) );
nand2 gate143( .a(G462), .b(G465), .O(G540) );
nand2 gate144( .a(G468), .b(G471), .O(G543) );
nand2 gate145( .a(G474), .b(G477), .O(G546) );
nand2 gate146( .a(G480), .b(G483), .O(G549) );
nand2 gate147( .a(G486), .b(G489), .O(G552) );

  xor2  gate1667(.a(G495), .b(G492), .O(gate148inter0));
  nand2 gate1668(.a(gate148inter0), .b(s_160), .O(gate148inter1));
  and2  gate1669(.a(G495), .b(G492), .O(gate148inter2));
  inv1  gate1670(.a(s_160), .O(gate148inter3));
  inv1  gate1671(.a(s_161), .O(gate148inter4));
  nand2 gate1672(.a(gate148inter4), .b(gate148inter3), .O(gate148inter5));
  nor2  gate1673(.a(gate148inter5), .b(gate148inter2), .O(gate148inter6));
  inv1  gate1674(.a(G492), .O(gate148inter7));
  inv1  gate1675(.a(G495), .O(gate148inter8));
  nand2 gate1676(.a(gate148inter8), .b(gate148inter7), .O(gate148inter9));
  nand2 gate1677(.a(s_161), .b(gate148inter3), .O(gate148inter10));
  nor2  gate1678(.a(gate148inter10), .b(gate148inter9), .O(gate148inter11));
  nor2  gate1679(.a(gate148inter11), .b(gate148inter6), .O(gate148inter12));
  nand2 gate1680(.a(gate148inter12), .b(gate148inter1), .O(G555));
nand2 gate149( .a(G498), .b(G501), .O(G558) );
nand2 gate150( .a(G504), .b(G507), .O(G561) );
nand2 gate151( .a(G510), .b(G513), .O(G564) );
nand2 gate152( .a(G516), .b(G519), .O(G567) );
nand2 gate153( .a(G426), .b(G522), .O(G570) );
nand2 gate154( .a(G429), .b(G522), .O(G571) );
nand2 gate155( .a(G432), .b(G525), .O(G572) );
nand2 gate156( .a(G435), .b(G525), .O(G573) );
nand2 gate157( .a(G438), .b(G528), .O(G574) );

  xor2  gate1681(.a(G528), .b(G441), .O(gate158inter0));
  nand2 gate1682(.a(gate158inter0), .b(s_162), .O(gate158inter1));
  and2  gate1683(.a(G528), .b(G441), .O(gate158inter2));
  inv1  gate1684(.a(s_162), .O(gate158inter3));
  inv1  gate1685(.a(s_163), .O(gate158inter4));
  nand2 gate1686(.a(gate158inter4), .b(gate158inter3), .O(gate158inter5));
  nor2  gate1687(.a(gate158inter5), .b(gate158inter2), .O(gate158inter6));
  inv1  gate1688(.a(G441), .O(gate158inter7));
  inv1  gate1689(.a(G528), .O(gate158inter8));
  nand2 gate1690(.a(gate158inter8), .b(gate158inter7), .O(gate158inter9));
  nand2 gate1691(.a(s_163), .b(gate158inter3), .O(gate158inter10));
  nor2  gate1692(.a(gate158inter10), .b(gate158inter9), .O(gate158inter11));
  nor2  gate1693(.a(gate158inter11), .b(gate158inter6), .O(gate158inter12));
  nand2 gate1694(.a(gate158inter12), .b(gate158inter1), .O(G575));
nand2 gate159( .a(G444), .b(G531), .O(G576) );

  xor2  gate1597(.a(G531), .b(G447), .O(gate160inter0));
  nand2 gate1598(.a(gate160inter0), .b(s_150), .O(gate160inter1));
  and2  gate1599(.a(G531), .b(G447), .O(gate160inter2));
  inv1  gate1600(.a(s_150), .O(gate160inter3));
  inv1  gate1601(.a(s_151), .O(gate160inter4));
  nand2 gate1602(.a(gate160inter4), .b(gate160inter3), .O(gate160inter5));
  nor2  gate1603(.a(gate160inter5), .b(gate160inter2), .O(gate160inter6));
  inv1  gate1604(.a(G447), .O(gate160inter7));
  inv1  gate1605(.a(G531), .O(gate160inter8));
  nand2 gate1606(.a(gate160inter8), .b(gate160inter7), .O(gate160inter9));
  nand2 gate1607(.a(s_151), .b(gate160inter3), .O(gate160inter10));
  nor2  gate1608(.a(gate160inter10), .b(gate160inter9), .O(gate160inter11));
  nor2  gate1609(.a(gate160inter11), .b(gate160inter6), .O(gate160inter12));
  nand2 gate1610(.a(gate160inter12), .b(gate160inter1), .O(G577));

  xor2  gate1289(.a(G534), .b(G450), .O(gate161inter0));
  nand2 gate1290(.a(gate161inter0), .b(s_106), .O(gate161inter1));
  and2  gate1291(.a(G534), .b(G450), .O(gate161inter2));
  inv1  gate1292(.a(s_106), .O(gate161inter3));
  inv1  gate1293(.a(s_107), .O(gate161inter4));
  nand2 gate1294(.a(gate161inter4), .b(gate161inter3), .O(gate161inter5));
  nor2  gate1295(.a(gate161inter5), .b(gate161inter2), .O(gate161inter6));
  inv1  gate1296(.a(G450), .O(gate161inter7));
  inv1  gate1297(.a(G534), .O(gate161inter8));
  nand2 gate1298(.a(gate161inter8), .b(gate161inter7), .O(gate161inter9));
  nand2 gate1299(.a(s_107), .b(gate161inter3), .O(gate161inter10));
  nor2  gate1300(.a(gate161inter10), .b(gate161inter9), .O(gate161inter11));
  nor2  gate1301(.a(gate161inter11), .b(gate161inter6), .O(gate161inter12));
  nand2 gate1302(.a(gate161inter12), .b(gate161inter1), .O(G578));
nand2 gate162( .a(G453), .b(G534), .O(G579) );
nand2 gate163( .a(G456), .b(G537), .O(G580) );
nand2 gate164( .a(G459), .b(G537), .O(G581) );

  xor2  gate911(.a(G540), .b(G462), .O(gate165inter0));
  nand2 gate912(.a(gate165inter0), .b(s_52), .O(gate165inter1));
  and2  gate913(.a(G540), .b(G462), .O(gate165inter2));
  inv1  gate914(.a(s_52), .O(gate165inter3));
  inv1  gate915(.a(s_53), .O(gate165inter4));
  nand2 gate916(.a(gate165inter4), .b(gate165inter3), .O(gate165inter5));
  nor2  gate917(.a(gate165inter5), .b(gate165inter2), .O(gate165inter6));
  inv1  gate918(.a(G462), .O(gate165inter7));
  inv1  gate919(.a(G540), .O(gate165inter8));
  nand2 gate920(.a(gate165inter8), .b(gate165inter7), .O(gate165inter9));
  nand2 gate921(.a(s_53), .b(gate165inter3), .O(gate165inter10));
  nor2  gate922(.a(gate165inter10), .b(gate165inter9), .O(gate165inter11));
  nor2  gate923(.a(gate165inter11), .b(gate165inter6), .O(gate165inter12));
  nand2 gate924(.a(gate165inter12), .b(gate165inter1), .O(G582));

  xor2  gate1457(.a(G540), .b(G465), .O(gate166inter0));
  nand2 gate1458(.a(gate166inter0), .b(s_130), .O(gate166inter1));
  and2  gate1459(.a(G540), .b(G465), .O(gate166inter2));
  inv1  gate1460(.a(s_130), .O(gate166inter3));
  inv1  gate1461(.a(s_131), .O(gate166inter4));
  nand2 gate1462(.a(gate166inter4), .b(gate166inter3), .O(gate166inter5));
  nor2  gate1463(.a(gate166inter5), .b(gate166inter2), .O(gate166inter6));
  inv1  gate1464(.a(G465), .O(gate166inter7));
  inv1  gate1465(.a(G540), .O(gate166inter8));
  nand2 gate1466(.a(gate166inter8), .b(gate166inter7), .O(gate166inter9));
  nand2 gate1467(.a(s_131), .b(gate166inter3), .O(gate166inter10));
  nor2  gate1468(.a(gate166inter10), .b(gate166inter9), .O(gate166inter11));
  nor2  gate1469(.a(gate166inter11), .b(gate166inter6), .O(gate166inter12));
  nand2 gate1470(.a(gate166inter12), .b(gate166inter1), .O(G583));
nand2 gate167( .a(G468), .b(G543), .O(G584) );
nand2 gate168( .a(G471), .b(G543), .O(G585) );

  xor2  gate1625(.a(G546), .b(G474), .O(gate169inter0));
  nand2 gate1626(.a(gate169inter0), .b(s_154), .O(gate169inter1));
  and2  gate1627(.a(G546), .b(G474), .O(gate169inter2));
  inv1  gate1628(.a(s_154), .O(gate169inter3));
  inv1  gate1629(.a(s_155), .O(gate169inter4));
  nand2 gate1630(.a(gate169inter4), .b(gate169inter3), .O(gate169inter5));
  nor2  gate1631(.a(gate169inter5), .b(gate169inter2), .O(gate169inter6));
  inv1  gate1632(.a(G474), .O(gate169inter7));
  inv1  gate1633(.a(G546), .O(gate169inter8));
  nand2 gate1634(.a(gate169inter8), .b(gate169inter7), .O(gate169inter9));
  nand2 gate1635(.a(s_155), .b(gate169inter3), .O(gate169inter10));
  nor2  gate1636(.a(gate169inter10), .b(gate169inter9), .O(gate169inter11));
  nor2  gate1637(.a(gate169inter11), .b(gate169inter6), .O(gate169inter12));
  nand2 gate1638(.a(gate169inter12), .b(gate169inter1), .O(G586));
nand2 gate170( .a(G477), .b(G546), .O(G587) );
nand2 gate171( .a(G480), .b(G549), .O(G588) );

  xor2  gate1821(.a(G549), .b(G483), .O(gate172inter0));
  nand2 gate1822(.a(gate172inter0), .b(s_182), .O(gate172inter1));
  and2  gate1823(.a(G549), .b(G483), .O(gate172inter2));
  inv1  gate1824(.a(s_182), .O(gate172inter3));
  inv1  gate1825(.a(s_183), .O(gate172inter4));
  nand2 gate1826(.a(gate172inter4), .b(gate172inter3), .O(gate172inter5));
  nor2  gate1827(.a(gate172inter5), .b(gate172inter2), .O(gate172inter6));
  inv1  gate1828(.a(G483), .O(gate172inter7));
  inv1  gate1829(.a(G549), .O(gate172inter8));
  nand2 gate1830(.a(gate172inter8), .b(gate172inter7), .O(gate172inter9));
  nand2 gate1831(.a(s_183), .b(gate172inter3), .O(gate172inter10));
  nor2  gate1832(.a(gate172inter10), .b(gate172inter9), .O(gate172inter11));
  nor2  gate1833(.a(gate172inter11), .b(gate172inter6), .O(gate172inter12));
  nand2 gate1834(.a(gate172inter12), .b(gate172inter1), .O(G589));
nand2 gate173( .a(G486), .b(G552), .O(G590) );

  xor2  gate1471(.a(G552), .b(G489), .O(gate174inter0));
  nand2 gate1472(.a(gate174inter0), .b(s_132), .O(gate174inter1));
  and2  gate1473(.a(G552), .b(G489), .O(gate174inter2));
  inv1  gate1474(.a(s_132), .O(gate174inter3));
  inv1  gate1475(.a(s_133), .O(gate174inter4));
  nand2 gate1476(.a(gate174inter4), .b(gate174inter3), .O(gate174inter5));
  nor2  gate1477(.a(gate174inter5), .b(gate174inter2), .O(gate174inter6));
  inv1  gate1478(.a(G489), .O(gate174inter7));
  inv1  gate1479(.a(G552), .O(gate174inter8));
  nand2 gate1480(.a(gate174inter8), .b(gate174inter7), .O(gate174inter9));
  nand2 gate1481(.a(s_133), .b(gate174inter3), .O(gate174inter10));
  nor2  gate1482(.a(gate174inter10), .b(gate174inter9), .O(gate174inter11));
  nor2  gate1483(.a(gate174inter11), .b(gate174inter6), .O(gate174inter12));
  nand2 gate1484(.a(gate174inter12), .b(gate174inter1), .O(G591));
nand2 gate175( .a(G492), .b(G555), .O(G592) );
nand2 gate176( .a(G495), .b(G555), .O(G593) );

  xor2  gate2087(.a(G558), .b(G498), .O(gate177inter0));
  nand2 gate2088(.a(gate177inter0), .b(s_220), .O(gate177inter1));
  and2  gate2089(.a(G558), .b(G498), .O(gate177inter2));
  inv1  gate2090(.a(s_220), .O(gate177inter3));
  inv1  gate2091(.a(s_221), .O(gate177inter4));
  nand2 gate2092(.a(gate177inter4), .b(gate177inter3), .O(gate177inter5));
  nor2  gate2093(.a(gate177inter5), .b(gate177inter2), .O(gate177inter6));
  inv1  gate2094(.a(G498), .O(gate177inter7));
  inv1  gate2095(.a(G558), .O(gate177inter8));
  nand2 gate2096(.a(gate177inter8), .b(gate177inter7), .O(gate177inter9));
  nand2 gate2097(.a(s_221), .b(gate177inter3), .O(gate177inter10));
  nor2  gate2098(.a(gate177inter10), .b(gate177inter9), .O(gate177inter11));
  nor2  gate2099(.a(gate177inter11), .b(gate177inter6), .O(gate177inter12));
  nand2 gate2100(.a(gate177inter12), .b(gate177inter1), .O(G594));
nand2 gate178( .a(G501), .b(G558), .O(G595) );

  xor2  gate575(.a(G561), .b(G504), .O(gate179inter0));
  nand2 gate576(.a(gate179inter0), .b(s_4), .O(gate179inter1));
  and2  gate577(.a(G561), .b(G504), .O(gate179inter2));
  inv1  gate578(.a(s_4), .O(gate179inter3));
  inv1  gate579(.a(s_5), .O(gate179inter4));
  nand2 gate580(.a(gate179inter4), .b(gate179inter3), .O(gate179inter5));
  nor2  gate581(.a(gate179inter5), .b(gate179inter2), .O(gate179inter6));
  inv1  gate582(.a(G504), .O(gate179inter7));
  inv1  gate583(.a(G561), .O(gate179inter8));
  nand2 gate584(.a(gate179inter8), .b(gate179inter7), .O(gate179inter9));
  nand2 gate585(.a(s_5), .b(gate179inter3), .O(gate179inter10));
  nor2  gate586(.a(gate179inter10), .b(gate179inter9), .O(gate179inter11));
  nor2  gate587(.a(gate179inter11), .b(gate179inter6), .O(gate179inter12));
  nand2 gate588(.a(gate179inter12), .b(gate179inter1), .O(G596));

  xor2  gate1387(.a(G561), .b(G507), .O(gate180inter0));
  nand2 gate1388(.a(gate180inter0), .b(s_120), .O(gate180inter1));
  and2  gate1389(.a(G561), .b(G507), .O(gate180inter2));
  inv1  gate1390(.a(s_120), .O(gate180inter3));
  inv1  gate1391(.a(s_121), .O(gate180inter4));
  nand2 gate1392(.a(gate180inter4), .b(gate180inter3), .O(gate180inter5));
  nor2  gate1393(.a(gate180inter5), .b(gate180inter2), .O(gate180inter6));
  inv1  gate1394(.a(G507), .O(gate180inter7));
  inv1  gate1395(.a(G561), .O(gate180inter8));
  nand2 gate1396(.a(gate180inter8), .b(gate180inter7), .O(gate180inter9));
  nand2 gate1397(.a(s_121), .b(gate180inter3), .O(gate180inter10));
  nor2  gate1398(.a(gate180inter10), .b(gate180inter9), .O(gate180inter11));
  nor2  gate1399(.a(gate180inter11), .b(gate180inter6), .O(gate180inter12));
  nand2 gate1400(.a(gate180inter12), .b(gate180inter1), .O(G597));
nand2 gate181( .a(G510), .b(G564), .O(G598) );
nand2 gate182( .a(G513), .b(G564), .O(G599) );
nand2 gate183( .a(G516), .b(G567), .O(G600) );
nand2 gate184( .a(G519), .b(G567), .O(G601) );

  xor2  gate2227(.a(G571), .b(G570), .O(gate185inter0));
  nand2 gate2228(.a(gate185inter0), .b(s_240), .O(gate185inter1));
  and2  gate2229(.a(G571), .b(G570), .O(gate185inter2));
  inv1  gate2230(.a(s_240), .O(gate185inter3));
  inv1  gate2231(.a(s_241), .O(gate185inter4));
  nand2 gate2232(.a(gate185inter4), .b(gate185inter3), .O(gate185inter5));
  nor2  gate2233(.a(gate185inter5), .b(gate185inter2), .O(gate185inter6));
  inv1  gate2234(.a(G570), .O(gate185inter7));
  inv1  gate2235(.a(G571), .O(gate185inter8));
  nand2 gate2236(.a(gate185inter8), .b(gate185inter7), .O(gate185inter9));
  nand2 gate2237(.a(s_241), .b(gate185inter3), .O(gate185inter10));
  nor2  gate2238(.a(gate185inter10), .b(gate185inter9), .O(gate185inter11));
  nor2  gate2239(.a(gate185inter11), .b(gate185inter6), .O(gate185inter12));
  nand2 gate2240(.a(gate185inter12), .b(gate185inter1), .O(G602));

  xor2  gate1415(.a(G573), .b(G572), .O(gate186inter0));
  nand2 gate1416(.a(gate186inter0), .b(s_124), .O(gate186inter1));
  and2  gate1417(.a(G573), .b(G572), .O(gate186inter2));
  inv1  gate1418(.a(s_124), .O(gate186inter3));
  inv1  gate1419(.a(s_125), .O(gate186inter4));
  nand2 gate1420(.a(gate186inter4), .b(gate186inter3), .O(gate186inter5));
  nor2  gate1421(.a(gate186inter5), .b(gate186inter2), .O(gate186inter6));
  inv1  gate1422(.a(G572), .O(gate186inter7));
  inv1  gate1423(.a(G573), .O(gate186inter8));
  nand2 gate1424(.a(gate186inter8), .b(gate186inter7), .O(gate186inter9));
  nand2 gate1425(.a(s_125), .b(gate186inter3), .O(gate186inter10));
  nor2  gate1426(.a(gate186inter10), .b(gate186inter9), .O(gate186inter11));
  nor2  gate1427(.a(gate186inter11), .b(gate186inter6), .O(gate186inter12));
  nand2 gate1428(.a(gate186inter12), .b(gate186inter1), .O(G607));

  xor2  gate1205(.a(G575), .b(G574), .O(gate187inter0));
  nand2 gate1206(.a(gate187inter0), .b(s_94), .O(gate187inter1));
  and2  gate1207(.a(G575), .b(G574), .O(gate187inter2));
  inv1  gate1208(.a(s_94), .O(gate187inter3));
  inv1  gate1209(.a(s_95), .O(gate187inter4));
  nand2 gate1210(.a(gate187inter4), .b(gate187inter3), .O(gate187inter5));
  nor2  gate1211(.a(gate187inter5), .b(gate187inter2), .O(gate187inter6));
  inv1  gate1212(.a(G574), .O(gate187inter7));
  inv1  gate1213(.a(G575), .O(gate187inter8));
  nand2 gate1214(.a(gate187inter8), .b(gate187inter7), .O(gate187inter9));
  nand2 gate1215(.a(s_95), .b(gate187inter3), .O(gate187inter10));
  nor2  gate1216(.a(gate187inter10), .b(gate187inter9), .O(gate187inter11));
  nor2  gate1217(.a(gate187inter11), .b(gate187inter6), .O(gate187inter12));
  nand2 gate1218(.a(gate187inter12), .b(gate187inter1), .O(G612));

  xor2  gate1905(.a(G577), .b(G576), .O(gate188inter0));
  nand2 gate1906(.a(gate188inter0), .b(s_194), .O(gate188inter1));
  and2  gate1907(.a(G577), .b(G576), .O(gate188inter2));
  inv1  gate1908(.a(s_194), .O(gate188inter3));
  inv1  gate1909(.a(s_195), .O(gate188inter4));
  nand2 gate1910(.a(gate188inter4), .b(gate188inter3), .O(gate188inter5));
  nor2  gate1911(.a(gate188inter5), .b(gate188inter2), .O(gate188inter6));
  inv1  gate1912(.a(G576), .O(gate188inter7));
  inv1  gate1913(.a(G577), .O(gate188inter8));
  nand2 gate1914(.a(gate188inter8), .b(gate188inter7), .O(gate188inter9));
  nand2 gate1915(.a(s_195), .b(gate188inter3), .O(gate188inter10));
  nor2  gate1916(.a(gate188inter10), .b(gate188inter9), .O(gate188inter11));
  nor2  gate1917(.a(gate188inter11), .b(gate188inter6), .O(gate188inter12));
  nand2 gate1918(.a(gate188inter12), .b(gate188inter1), .O(G617));

  xor2  gate1345(.a(G579), .b(G578), .O(gate189inter0));
  nand2 gate1346(.a(gate189inter0), .b(s_114), .O(gate189inter1));
  and2  gate1347(.a(G579), .b(G578), .O(gate189inter2));
  inv1  gate1348(.a(s_114), .O(gate189inter3));
  inv1  gate1349(.a(s_115), .O(gate189inter4));
  nand2 gate1350(.a(gate189inter4), .b(gate189inter3), .O(gate189inter5));
  nor2  gate1351(.a(gate189inter5), .b(gate189inter2), .O(gate189inter6));
  inv1  gate1352(.a(G578), .O(gate189inter7));
  inv1  gate1353(.a(G579), .O(gate189inter8));
  nand2 gate1354(.a(gate189inter8), .b(gate189inter7), .O(gate189inter9));
  nand2 gate1355(.a(s_115), .b(gate189inter3), .O(gate189inter10));
  nor2  gate1356(.a(gate189inter10), .b(gate189inter9), .O(gate189inter11));
  nor2  gate1357(.a(gate189inter11), .b(gate189inter6), .O(gate189inter12));
  nand2 gate1358(.a(gate189inter12), .b(gate189inter1), .O(G622));
nand2 gate190( .a(G580), .b(G581), .O(G627) );

  xor2  gate1443(.a(G583), .b(G582), .O(gate191inter0));
  nand2 gate1444(.a(gate191inter0), .b(s_128), .O(gate191inter1));
  and2  gate1445(.a(G583), .b(G582), .O(gate191inter2));
  inv1  gate1446(.a(s_128), .O(gate191inter3));
  inv1  gate1447(.a(s_129), .O(gate191inter4));
  nand2 gate1448(.a(gate191inter4), .b(gate191inter3), .O(gate191inter5));
  nor2  gate1449(.a(gate191inter5), .b(gate191inter2), .O(gate191inter6));
  inv1  gate1450(.a(G582), .O(gate191inter7));
  inv1  gate1451(.a(G583), .O(gate191inter8));
  nand2 gate1452(.a(gate191inter8), .b(gate191inter7), .O(gate191inter9));
  nand2 gate1453(.a(s_129), .b(gate191inter3), .O(gate191inter10));
  nor2  gate1454(.a(gate191inter10), .b(gate191inter9), .O(gate191inter11));
  nor2  gate1455(.a(gate191inter11), .b(gate191inter6), .O(gate191inter12));
  nand2 gate1456(.a(gate191inter12), .b(gate191inter1), .O(G632));
nand2 gate192( .a(G584), .b(G585), .O(G637) );
nand2 gate193( .a(G586), .b(G587), .O(G642) );

  xor2  gate743(.a(G589), .b(G588), .O(gate194inter0));
  nand2 gate744(.a(gate194inter0), .b(s_28), .O(gate194inter1));
  and2  gate745(.a(G589), .b(G588), .O(gate194inter2));
  inv1  gate746(.a(s_28), .O(gate194inter3));
  inv1  gate747(.a(s_29), .O(gate194inter4));
  nand2 gate748(.a(gate194inter4), .b(gate194inter3), .O(gate194inter5));
  nor2  gate749(.a(gate194inter5), .b(gate194inter2), .O(gate194inter6));
  inv1  gate750(.a(G588), .O(gate194inter7));
  inv1  gate751(.a(G589), .O(gate194inter8));
  nand2 gate752(.a(gate194inter8), .b(gate194inter7), .O(gate194inter9));
  nand2 gate753(.a(s_29), .b(gate194inter3), .O(gate194inter10));
  nor2  gate754(.a(gate194inter10), .b(gate194inter9), .O(gate194inter11));
  nor2  gate755(.a(gate194inter11), .b(gate194inter6), .O(gate194inter12));
  nand2 gate756(.a(gate194inter12), .b(gate194inter1), .O(G645));
nand2 gate195( .a(G590), .b(G591), .O(G648) );

  xor2  gate2101(.a(G593), .b(G592), .O(gate196inter0));
  nand2 gate2102(.a(gate196inter0), .b(s_222), .O(gate196inter1));
  and2  gate2103(.a(G593), .b(G592), .O(gate196inter2));
  inv1  gate2104(.a(s_222), .O(gate196inter3));
  inv1  gate2105(.a(s_223), .O(gate196inter4));
  nand2 gate2106(.a(gate196inter4), .b(gate196inter3), .O(gate196inter5));
  nor2  gate2107(.a(gate196inter5), .b(gate196inter2), .O(gate196inter6));
  inv1  gate2108(.a(G592), .O(gate196inter7));
  inv1  gate2109(.a(G593), .O(gate196inter8));
  nand2 gate2110(.a(gate196inter8), .b(gate196inter7), .O(gate196inter9));
  nand2 gate2111(.a(s_223), .b(gate196inter3), .O(gate196inter10));
  nor2  gate2112(.a(gate196inter10), .b(gate196inter9), .O(gate196inter11));
  nor2  gate2113(.a(gate196inter11), .b(gate196inter6), .O(gate196inter12));
  nand2 gate2114(.a(gate196inter12), .b(gate196inter1), .O(G651));
nand2 gate197( .a(G594), .b(G595), .O(G654) );
nand2 gate198( .a(G596), .b(G597), .O(G657) );
nand2 gate199( .a(G598), .b(G599), .O(G660) );
nand2 gate200( .a(G600), .b(G601), .O(G663) );
nand2 gate201( .a(G602), .b(G607), .O(G666) );
nand2 gate202( .a(G612), .b(G617), .O(G669) );
nand2 gate203( .a(G602), .b(G612), .O(G672) );
nand2 gate204( .a(G607), .b(G617), .O(G675) );

  xor2  gate1275(.a(G627), .b(G622), .O(gate205inter0));
  nand2 gate1276(.a(gate205inter0), .b(s_104), .O(gate205inter1));
  and2  gate1277(.a(G627), .b(G622), .O(gate205inter2));
  inv1  gate1278(.a(s_104), .O(gate205inter3));
  inv1  gate1279(.a(s_105), .O(gate205inter4));
  nand2 gate1280(.a(gate205inter4), .b(gate205inter3), .O(gate205inter5));
  nor2  gate1281(.a(gate205inter5), .b(gate205inter2), .O(gate205inter6));
  inv1  gate1282(.a(G622), .O(gate205inter7));
  inv1  gate1283(.a(G627), .O(gate205inter8));
  nand2 gate1284(.a(gate205inter8), .b(gate205inter7), .O(gate205inter9));
  nand2 gate1285(.a(s_105), .b(gate205inter3), .O(gate205inter10));
  nor2  gate1286(.a(gate205inter10), .b(gate205inter9), .O(gate205inter11));
  nor2  gate1287(.a(gate205inter11), .b(gate205inter6), .O(gate205inter12));
  nand2 gate1288(.a(gate205inter12), .b(gate205inter1), .O(G678));
nand2 gate206( .a(G632), .b(G637), .O(G681) );

  xor2  gate2185(.a(G632), .b(G622), .O(gate207inter0));
  nand2 gate2186(.a(gate207inter0), .b(s_234), .O(gate207inter1));
  and2  gate2187(.a(G632), .b(G622), .O(gate207inter2));
  inv1  gate2188(.a(s_234), .O(gate207inter3));
  inv1  gate2189(.a(s_235), .O(gate207inter4));
  nand2 gate2190(.a(gate207inter4), .b(gate207inter3), .O(gate207inter5));
  nor2  gate2191(.a(gate207inter5), .b(gate207inter2), .O(gate207inter6));
  inv1  gate2192(.a(G622), .O(gate207inter7));
  inv1  gate2193(.a(G632), .O(gate207inter8));
  nand2 gate2194(.a(gate207inter8), .b(gate207inter7), .O(gate207inter9));
  nand2 gate2195(.a(s_235), .b(gate207inter3), .O(gate207inter10));
  nor2  gate2196(.a(gate207inter10), .b(gate207inter9), .O(gate207inter11));
  nor2  gate2197(.a(gate207inter11), .b(gate207inter6), .O(gate207inter12));
  nand2 gate2198(.a(gate207inter12), .b(gate207inter1), .O(G684));
nand2 gate208( .a(G627), .b(G637), .O(G687) );
nand2 gate209( .a(G602), .b(G666), .O(G690) );
nand2 gate210( .a(G607), .b(G666), .O(G691) );
nand2 gate211( .a(G612), .b(G669), .O(G692) );
nand2 gate212( .a(G617), .b(G669), .O(G693) );

  xor2  gate1401(.a(G672), .b(G602), .O(gate213inter0));
  nand2 gate1402(.a(gate213inter0), .b(s_122), .O(gate213inter1));
  and2  gate1403(.a(G672), .b(G602), .O(gate213inter2));
  inv1  gate1404(.a(s_122), .O(gate213inter3));
  inv1  gate1405(.a(s_123), .O(gate213inter4));
  nand2 gate1406(.a(gate213inter4), .b(gate213inter3), .O(gate213inter5));
  nor2  gate1407(.a(gate213inter5), .b(gate213inter2), .O(gate213inter6));
  inv1  gate1408(.a(G602), .O(gate213inter7));
  inv1  gate1409(.a(G672), .O(gate213inter8));
  nand2 gate1410(.a(gate213inter8), .b(gate213inter7), .O(gate213inter9));
  nand2 gate1411(.a(s_123), .b(gate213inter3), .O(gate213inter10));
  nor2  gate1412(.a(gate213inter10), .b(gate213inter9), .O(gate213inter11));
  nor2  gate1413(.a(gate213inter11), .b(gate213inter6), .O(gate213inter12));
  nand2 gate1414(.a(gate213inter12), .b(gate213inter1), .O(G694));
nand2 gate214( .a(G612), .b(G672), .O(G695) );
nand2 gate215( .a(G607), .b(G675), .O(G696) );

  xor2  gate799(.a(G675), .b(G617), .O(gate216inter0));
  nand2 gate800(.a(gate216inter0), .b(s_36), .O(gate216inter1));
  and2  gate801(.a(G675), .b(G617), .O(gate216inter2));
  inv1  gate802(.a(s_36), .O(gate216inter3));
  inv1  gate803(.a(s_37), .O(gate216inter4));
  nand2 gate804(.a(gate216inter4), .b(gate216inter3), .O(gate216inter5));
  nor2  gate805(.a(gate216inter5), .b(gate216inter2), .O(gate216inter6));
  inv1  gate806(.a(G617), .O(gate216inter7));
  inv1  gate807(.a(G675), .O(gate216inter8));
  nand2 gate808(.a(gate216inter8), .b(gate216inter7), .O(gate216inter9));
  nand2 gate809(.a(s_37), .b(gate216inter3), .O(gate216inter10));
  nor2  gate810(.a(gate216inter10), .b(gate216inter9), .O(gate216inter11));
  nor2  gate811(.a(gate216inter11), .b(gate216inter6), .O(gate216inter12));
  nand2 gate812(.a(gate216inter12), .b(gate216inter1), .O(G697));
nand2 gate217( .a(G622), .b(G678), .O(G698) );
nand2 gate218( .a(G627), .b(G678), .O(G699) );
nand2 gate219( .a(G632), .b(G681), .O(G700) );
nand2 gate220( .a(G637), .b(G681), .O(G701) );
nand2 gate221( .a(G622), .b(G684), .O(G702) );

  xor2  gate1947(.a(G684), .b(G632), .O(gate222inter0));
  nand2 gate1948(.a(gate222inter0), .b(s_200), .O(gate222inter1));
  and2  gate1949(.a(G684), .b(G632), .O(gate222inter2));
  inv1  gate1950(.a(s_200), .O(gate222inter3));
  inv1  gate1951(.a(s_201), .O(gate222inter4));
  nand2 gate1952(.a(gate222inter4), .b(gate222inter3), .O(gate222inter5));
  nor2  gate1953(.a(gate222inter5), .b(gate222inter2), .O(gate222inter6));
  inv1  gate1954(.a(G632), .O(gate222inter7));
  inv1  gate1955(.a(G684), .O(gate222inter8));
  nand2 gate1956(.a(gate222inter8), .b(gate222inter7), .O(gate222inter9));
  nand2 gate1957(.a(s_201), .b(gate222inter3), .O(gate222inter10));
  nor2  gate1958(.a(gate222inter10), .b(gate222inter9), .O(gate222inter11));
  nor2  gate1959(.a(gate222inter11), .b(gate222inter6), .O(gate222inter12));
  nand2 gate1960(.a(gate222inter12), .b(gate222inter1), .O(G703));

  xor2  gate715(.a(G687), .b(G627), .O(gate223inter0));
  nand2 gate716(.a(gate223inter0), .b(s_24), .O(gate223inter1));
  and2  gate717(.a(G687), .b(G627), .O(gate223inter2));
  inv1  gate718(.a(s_24), .O(gate223inter3));
  inv1  gate719(.a(s_25), .O(gate223inter4));
  nand2 gate720(.a(gate223inter4), .b(gate223inter3), .O(gate223inter5));
  nor2  gate721(.a(gate223inter5), .b(gate223inter2), .O(gate223inter6));
  inv1  gate722(.a(G627), .O(gate223inter7));
  inv1  gate723(.a(G687), .O(gate223inter8));
  nand2 gate724(.a(gate223inter8), .b(gate223inter7), .O(gate223inter9));
  nand2 gate725(.a(s_25), .b(gate223inter3), .O(gate223inter10));
  nor2  gate726(.a(gate223inter10), .b(gate223inter9), .O(gate223inter11));
  nor2  gate727(.a(gate223inter11), .b(gate223inter6), .O(gate223inter12));
  nand2 gate728(.a(gate223inter12), .b(gate223inter1), .O(G704));
nand2 gate224( .a(G637), .b(G687), .O(G705) );
nand2 gate225( .a(G690), .b(G691), .O(G706) );
nand2 gate226( .a(G692), .b(G693), .O(G709) );
nand2 gate227( .a(G694), .b(G695), .O(G712) );
nand2 gate228( .a(G696), .b(G697), .O(G715) );
nand2 gate229( .a(G698), .b(G699), .O(G718) );
nand2 gate230( .a(G700), .b(G701), .O(G721) );
nand2 gate231( .a(G702), .b(G703), .O(G724) );

  xor2  gate2143(.a(G705), .b(G704), .O(gate232inter0));
  nand2 gate2144(.a(gate232inter0), .b(s_228), .O(gate232inter1));
  and2  gate2145(.a(G705), .b(G704), .O(gate232inter2));
  inv1  gate2146(.a(s_228), .O(gate232inter3));
  inv1  gate2147(.a(s_229), .O(gate232inter4));
  nand2 gate2148(.a(gate232inter4), .b(gate232inter3), .O(gate232inter5));
  nor2  gate2149(.a(gate232inter5), .b(gate232inter2), .O(gate232inter6));
  inv1  gate2150(.a(G704), .O(gate232inter7));
  inv1  gate2151(.a(G705), .O(gate232inter8));
  nand2 gate2152(.a(gate232inter8), .b(gate232inter7), .O(gate232inter9));
  nand2 gate2153(.a(s_229), .b(gate232inter3), .O(gate232inter10));
  nor2  gate2154(.a(gate232inter10), .b(gate232inter9), .O(gate232inter11));
  nor2  gate2155(.a(gate232inter11), .b(gate232inter6), .O(gate232inter12));
  nand2 gate2156(.a(gate232inter12), .b(gate232inter1), .O(G727));
nand2 gate233( .a(G242), .b(G718), .O(G730) );
nand2 gate234( .a(G245), .b(G721), .O(G733) );

  xor2  gate547(.a(G724), .b(G248), .O(gate235inter0));
  nand2 gate548(.a(gate235inter0), .b(s_0), .O(gate235inter1));
  and2  gate549(.a(G724), .b(G248), .O(gate235inter2));
  inv1  gate550(.a(s_0), .O(gate235inter3));
  inv1  gate551(.a(s_1), .O(gate235inter4));
  nand2 gate552(.a(gate235inter4), .b(gate235inter3), .O(gate235inter5));
  nor2  gate553(.a(gate235inter5), .b(gate235inter2), .O(gate235inter6));
  inv1  gate554(.a(G248), .O(gate235inter7));
  inv1  gate555(.a(G724), .O(gate235inter8));
  nand2 gate556(.a(gate235inter8), .b(gate235inter7), .O(gate235inter9));
  nand2 gate557(.a(s_1), .b(gate235inter3), .O(gate235inter10));
  nor2  gate558(.a(gate235inter10), .b(gate235inter9), .O(gate235inter11));
  nor2  gate559(.a(gate235inter11), .b(gate235inter6), .O(gate235inter12));
  nand2 gate560(.a(gate235inter12), .b(gate235inter1), .O(G736));
nand2 gate236( .a(G251), .b(G727), .O(G739) );

  xor2  gate1793(.a(G706), .b(G254), .O(gate237inter0));
  nand2 gate1794(.a(gate237inter0), .b(s_178), .O(gate237inter1));
  and2  gate1795(.a(G706), .b(G254), .O(gate237inter2));
  inv1  gate1796(.a(s_178), .O(gate237inter3));
  inv1  gate1797(.a(s_179), .O(gate237inter4));
  nand2 gate1798(.a(gate237inter4), .b(gate237inter3), .O(gate237inter5));
  nor2  gate1799(.a(gate237inter5), .b(gate237inter2), .O(gate237inter6));
  inv1  gate1800(.a(G254), .O(gate237inter7));
  inv1  gate1801(.a(G706), .O(gate237inter8));
  nand2 gate1802(.a(gate237inter8), .b(gate237inter7), .O(gate237inter9));
  nand2 gate1803(.a(s_179), .b(gate237inter3), .O(gate237inter10));
  nor2  gate1804(.a(gate237inter10), .b(gate237inter9), .O(gate237inter11));
  nor2  gate1805(.a(gate237inter11), .b(gate237inter6), .O(gate237inter12));
  nand2 gate1806(.a(gate237inter12), .b(gate237inter1), .O(G742));

  xor2  gate1863(.a(G709), .b(G257), .O(gate238inter0));
  nand2 gate1864(.a(gate238inter0), .b(s_188), .O(gate238inter1));
  and2  gate1865(.a(G709), .b(G257), .O(gate238inter2));
  inv1  gate1866(.a(s_188), .O(gate238inter3));
  inv1  gate1867(.a(s_189), .O(gate238inter4));
  nand2 gate1868(.a(gate238inter4), .b(gate238inter3), .O(gate238inter5));
  nor2  gate1869(.a(gate238inter5), .b(gate238inter2), .O(gate238inter6));
  inv1  gate1870(.a(G257), .O(gate238inter7));
  inv1  gate1871(.a(G709), .O(gate238inter8));
  nand2 gate1872(.a(gate238inter8), .b(gate238inter7), .O(gate238inter9));
  nand2 gate1873(.a(s_189), .b(gate238inter3), .O(gate238inter10));
  nor2  gate1874(.a(gate238inter10), .b(gate238inter9), .O(gate238inter11));
  nor2  gate1875(.a(gate238inter11), .b(gate238inter6), .O(gate238inter12));
  nand2 gate1876(.a(gate238inter12), .b(gate238inter1), .O(G745));
nand2 gate239( .a(G260), .b(G712), .O(G748) );

  xor2  gate2311(.a(G715), .b(G263), .O(gate240inter0));
  nand2 gate2312(.a(gate240inter0), .b(s_252), .O(gate240inter1));
  and2  gate2313(.a(G715), .b(G263), .O(gate240inter2));
  inv1  gate2314(.a(s_252), .O(gate240inter3));
  inv1  gate2315(.a(s_253), .O(gate240inter4));
  nand2 gate2316(.a(gate240inter4), .b(gate240inter3), .O(gate240inter5));
  nor2  gate2317(.a(gate240inter5), .b(gate240inter2), .O(gate240inter6));
  inv1  gate2318(.a(G263), .O(gate240inter7));
  inv1  gate2319(.a(G715), .O(gate240inter8));
  nand2 gate2320(.a(gate240inter8), .b(gate240inter7), .O(gate240inter9));
  nand2 gate2321(.a(s_253), .b(gate240inter3), .O(gate240inter10));
  nor2  gate2322(.a(gate240inter10), .b(gate240inter9), .O(gate240inter11));
  nor2  gate2323(.a(gate240inter11), .b(gate240inter6), .O(gate240inter12));
  nand2 gate2324(.a(gate240inter12), .b(gate240inter1), .O(G751));
nand2 gate241( .a(G242), .b(G730), .O(G754) );
nand2 gate242( .a(G718), .b(G730), .O(G755) );

  xor2  gate1317(.a(G733), .b(G245), .O(gate243inter0));
  nand2 gate1318(.a(gate243inter0), .b(s_110), .O(gate243inter1));
  and2  gate1319(.a(G733), .b(G245), .O(gate243inter2));
  inv1  gate1320(.a(s_110), .O(gate243inter3));
  inv1  gate1321(.a(s_111), .O(gate243inter4));
  nand2 gate1322(.a(gate243inter4), .b(gate243inter3), .O(gate243inter5));
  nor2  gate1323(.a(gate243inter5), .b(gate243inter2), .O(gate243inter6));
  inv1  gate1324(.a(G245), .O(gate243inter7));
  inv1  gate1325(.a(G733), .O(gate243inter8));
  nand2 gate1326(.a(gate243inter8), .b(gate243inter7), .O(gate243inter9));
  nand2 gate1327(.a(s_111), .b(gate243inter3), .O(gate243inter10));
  nor2  gate1328(.a(gate243inter10), .b(gate243inter9), .O(gate243inter11));
  nor2  gate1329(.a(gate243inter11), .b(gate243inter6), .O(gate243inter12));
  nand2 gate1330(.a(gate243inter12), .b(gate243inter1), .O(G756));

  xor2  gate561(.a(G733), .b(G721), .O(gate244inter0));
  nand2 gate562(.a(gate244inter0), .b(s_2), .O(gate244inter1));
  and2  gate563(.a(G733), .b(G721), .O(gate244inter2));
  inv1  gate564(.a(s_2), .O(gate244inter3));
  inv1  gate565(.a(s_3), .O(gate244inter4));
  nand2 gate566(.a(gate244inter4), .b(gate244inter3), .O(gate244inter5));
  nor2  gate567(.a(gate244inter5), .b(gate244inter2), .O(gate244inter6));
  inv1  gate568(.a(G721), .O(gate244inter7));
  inv1  gate569(.a(G733), .O(gate244inter8));
  nand2 gate570(.a(gate244inter8), .b(gate244inter7), .O(gate244inter9));
  nand2 gate571(.a(s_3), .b(gate244inter3), .O(gate244inter10));
  nor2  gate572(.a(gate244inter10), .b(gate244inter9), .O(gate244inter11));
  nor2  gate573(.a(gate244inter11), .b(gate244inter6), .O(gate244inter12));
  nand2 gate574(.a(gate244inter12), .b(gate244inter1), .O(G757));
nand2 gate245( .a(G248), .b(G736), .O(G758) );
nand2 gate246( .a(G724), .b(G736), .O(G759) );
nand2 gate247( .a(G251), .b(G739), .O(G760) );

  xor2  gate1331(.a(G739), .b(G727), .O(gate248inter0));
  nand2 gate1332(.a(gate248inter0), .b(s_112), .O(gate248inter1));
  and2  gate1333(.a(G739), .b(G727), .O(gate248inter2));
  inv1  gate1334(.a(s_112), .O(gate248inter3));
  inv1  gate1335(.a(s_113), .O(gate248inter4));
  nand2 gate1336(.a(gate248inter4), .b(gate248inter3), .O(gate248inter5));
  nor2  gate1337(.a(gate248inter5), .b(gate248inter2), .O(gate248inter6));
  inv1  gate1338(.a(G727), .O(gate248inter7));
  inv1  gate1339(.a(G739), .O(gate248inter8));
  nand2 gate1340(.a(gate248inter8), .b(gate248inter7), .O(gate248inter9));
  nand2 gate1341(.a(s_113), .b(gate248inter3), .O(gate248inter10));
  nor2  gate1342(.a(gate248inter10), .b(gate248inter9), .O(gate248inter11));
  nor2  gate1343(.a(gate248inter11), .b(gate248inter6), .O(gate248inter12));
  nand2 gate1344(.a(gate248inter12), .b(gate248inter1), .O(G761));
nand2 gate249( .a(G254), .b(G742), .O(G762) );
nand2 gate250( .a(G706), .b(G742), .O(G763) );
nand2 gate251( .a(G257), .b(G745), .O(G764) );
nand2 gate252( .a(G709), .b(G745), .O(G765) );
nand2 gate253( .a(G260), .b(G748), .O(G766) );
nand2 gate254( .a(G712), .b(G748), .O(G767) );
nand2 gate255( .a(G263), .b(G751), .O(G768) );
nand2 gate256( .a(G715), .b(G751), .O(G769) );
nand2 gate257( .a(G754), .b(G755), .O(G770) );

  xor2  gate1919(.a(G757), .b(G756), .O(gate258inter0));
  nand2 gate1920(.a(gate258inter0), .b(s_196), .O(gate258inter1));
  and2  gate1921(.a(G757), .b(G756), .O(gate258inter2));
  inv1  gate1922(.a(s_196), .O(gate258inter3));
  inv1  gate1923(.a(s_197), .O(gate258inter4));
  nand2 gate1924(.a(gate258inter4), .b(gate258inter3), .O(gate258inter5));
  nor2  gate1925(.a(gate258inter5), .b(gate258inter2), .O(gate258inter6));
  inv1  gate1926(.a(G756), .O(gate258inter7));
  inv1  gate1927(.a(G757), .O(gate258inter8));
  nand2 gate1928(.a(gate258inter8), .b(gate258inter7), .O(gate258inter9));
  nand2 gate1929(.a(s_197), .b(gate258inter3), .O(gate258inter10));
  nor2  gate1930(.a(gate258inter10), .b(gate258inter9), .O(gate258inter11));
  nor2  gate1931(.a(gate258inter11), .b(gate258inter6), .O(gate258inter12));
  nand2 gate1932(.a(gate258inter12), .b(gate258inter1), .O(G773));
nand2 gate259( .a(G758), .b(G759), .O(G776) );
nand2 gate260( .a(G760), .b(G761), .O(G779) );

  xor2  gate1037(.a(G763), .b(G762), .O(gate261inter0));
  nand2 gate1038(.a(gate261inter0), .b(s_70), .O(gate261inter1));
  and2  gate1039(.a(G763), .b(G762), .O(gate261inter2));
  inv1  gate1040(.a(s_70), .O(gate261inter3));
  inv1  gate1041(.a(s_71), .O(gate261inter4));
  nand2 gate1042(.a(gate261inter4), .b(gate261inter3), .O(gate261inter5));
  nor2  gate1043(.a(gate261inter5), .b(gate261inter2), .O(gate261inter6));
  inv1  gate1044(.a(G762), .O(gate261inter7));
  inv1  gate1045(.a(G763), .O(gate261inter8));
  nand2 gate1046(.a(gate261inter8), .b(gate261inter7), .O(gate261inter9));
  nand2 gate1047(.a(s_71), .b(gate261inter3), .O(gate261inter10));
  nor2  gate1048(.a(gate261inter10), .b(gate261inter9), .O(gate261inter11));
  nor2  gate1049(.a(gate261inter11), .b(gate261inter6), .O(gate261inter12));
  nand2 gate1050(.a(gate261inter12), .b(gate261inter1), .O(G782));
nand2 gate262( .a(G764), .b(G765), .O(G785) );

  xor2  gate673(.a(G767), .b(G766), .O(gate263inter0));
  nand2 gate674(.a(gate263inter0), .b(s_18), .O(gate263inter1));
  and2  gate675(.a(G767), .b(G766), .O(gate263inter2));
  inv1  gate676(.a(s_18), .O(gate263inter3));
  inv1  gate677(.a(s_19), .O(gate263inter4));
  nand2 gate678(.a(gate263inter4), .b(gate263inter3), .O(gate263inter5));
  nor2  gate679(.a(gate263inter5), .b(gate263inter2), .O(gate263inter6));
  inv1  gate680(.a(G766), .O(gate263inter7));
  inv1  gate681(.a(G767), .O(gate263inter8));
  nand2 gate682(.a(gate263inter8), .b(gate263inter7), .O(gate263inter9));
  nand2 gate683(.a(s_19), .b(gate263inter3), .O(gate263inter10));
  nor2  gate684(.a(gate263inter10), .b(gate263inter9), .O(gate263inter11));
  nor2  gate685(.a(gate263inter11), .b(gate263inter6), .O(gate263inter12));
  nand2 gate686(.a(gate263inter12), .b(gate263inter1), .O(G788));

  xor2  gate2269(.a(G769), .b(G768), .O(gate264inter0));
  nand2 gate2270(.a(gate264inter0), .b(s_246), .O(gate264inter1));
  and2  gate2271(.a(G769), .b(G768), .O(gate264inter2));
  inv1  gate2272(.a(s_246), .O(gate264inter3));
  inv1  gate2273(.a(s_247), .O(gate264inter4));
  nand2 gate2274(.a(gate264inter4), .b(gate264inter3), .O(gate264inter5));
  nor2  gate2275(.a(gate264inter5), .b(gate264inter2), .O(gate264inter6));
  inv1  gate2276(.a(G768), .O(gate264inter7));
  inv1  gate2277(.a(G769), .O(gate264inter8));
  nand2 gate2278(.a(gate264inter8), .b(gate264inter7), .O(gate264inter9));
  nand2 gate2279(.a(s_247), .b(gate264inter3), .O(gate264inter10));
  nor2  gate2280(.a(gate264inter10), .b(gate264inter9), .O(gate264inter11));
  nor2  gate2281(.a(gate264inter11), .b(gate264inter6), .O(gate264inter12));
  nand2 gate2282(.a(gate264inter12), .b(gate264inter1), .O(G791));
nand2 gate265( .a(G642), .b(G770), .O(G794) );

  xor2  gate1751(.a(G773), .b(G645), .O(gate266inter0));
  nand2 gate1752(.a(gate266inter0), .b(s_172), .O(gate266inter1));
  and2  gate1753(.a(G773), .b(G645), .O(gate266inter2));
  inv1  gate1754(.a(s_172), .O(gate266inter3));
  inv1  gate1755(.a(s_173), .O(gate266inter4));
  nand2 gate1756(.a(gate266inter4), .b(gate266inter3), .O(gate266inter5));
  nor2  gate1757(.a(gate266inter5), .b(gate266inter2), .O(gate266inter6));
  inv1  gate1758(.a(G645), .O(gate266inter7));
  inv1  gate1759(.a(G773), .O(gate266inter8));
  nand2 gate1760(.a(gate266inter8), .b(gate266inter7), .O(gate266inter9));
  nand2 gate1761(.a(s_173), .b(gate266inter3), .O(gate266inter10));
  nor2  gate1762(.a(gate266inter10), .b(gate266inter9), .O(gate266inter11));
  nor2  gate1763(.a(gate266inter11), .b(gate266inter6), .O(gate266inter12));
  nand2 gate1764(.a(gate266inter12), .b(gate266inter1), .O(G797));

  xor2  gate1569(.a(G776), .b(G648), .O(gate267inter0));
  nand2 gate1570(.a(gate267inter0), .b(s_146), .O(gate267inter1));
  and2  gate1571(.a(G776), .b(G648), .O(gate267inter2));
  inv1  gate1572(.a(s_146), .O(gate267inter3));
  inv1  gate1573(.a(s_147), .O(gate267inter4));
  nand2 gate1574(.a(gate267inter4), .b(gate267inter3), .O(gate267inter5));
  nor2  gate1575(.a(gate267inter5), .b(gate267inter2), .O(gate267inter6));
  inv1  gate1576(.a(G648), .O(gate267inter7));
  inv1  gate1577(.a(G776), .O(gate267inter8));
  nand2 gate1578(.a(gate267inter8), .b(gate267inter7), .O(gate267inter9));
  nand2 gate1579(.a(s_147), .b(gate267inter3), .O(gate267inter10));
  nor2  gate1580(.a(gate267inter10), .b(gate267inter9), .O(gate267inter11));
  nor2  gate1581(.a(gate267inter11), .b(gate267inter6), .O(gate267inter12));
  nand2 gate1582(.a(gate267inter12), .b(gate267inter1), .O(G800));
nand2 gate268( .a(G651), .b(G779), .O(G803) );
nand2 gate269( .a(G654), .b(G782), .O(G806) );
nand2 gate270( .a(G657), .b(G785), .O(G809) );
nand2 gate271( .a(G660), .b(G788), .O(G812) );
nand2 gate272( .a(G663), .b(G791), .O(G815) );

  xor2  gate2171(.a(G794), .b(G642), .O(gate273inter0));
  nand2 gate2172(.a(gate273inter0), .b(s_232), .O(gate273inter1));
  and2  gate2173(.a(G794), .b(G642), .O(gate273inter2));
  inv1  gate2174(.a(s_232), .O(gate273inter3));
  inv1  gate2175(.a(s_233), .O(gate273inter4));
  nand2 gate2176(.a(gate273inter4), .b(gate273inter3), .O(gate273inter5));
  nor2  gate2177(.a(gate273inter5), .b(gate273inter2), .O(gate273inter6));
  inv1  gate2178(.a(G642), .O(gate273inter7));
  inv1  gate2179(.a(G794), .O(gate273inter8));
  nand2 gate2180(.a(gate273inter8), .b(gate273inter7), .O(gate273inter9));
  nand2 gate2181(.a(s_233), .b(gate273inter3), .O(gate273inter10));
  nor2  gate2182(.a(gate273inter10), .b(gate273inter9), .O(gate273inter11));
  nor2  gate2183(.a(gate273inter11), .b(gate273inter6), .O(gate273inter12));
  nand2 gate2184(.a(gate273inter12), .b(gate273inter1), .O(G818));
nand2 gate274( .a(G770), .b(G794), .O(G819) );

  xor2  gate2031(.a(G797), .b(G645), .O(gate275inter0));
  nand2 gate2032(.a(gate275inter0), .b(s_212), .O(gate275inter1));
  and2  gate2033(.a(G797), .b(G645), .O(gate275inter2));
  inv1  gate2034(.a(s_212), .O(gate275inter3));
  inv1  gate2035(.a(s_213), .O(gate275inter4));
  nand2 gate2036(.a(gate275inter4), .b(gate275inter3), .O(gate275inter5));
  nor2  gate2037(.a(gate275inter5), .b(gate275inter2), .O(gate275inter6));
  inv1  gate2038(.a(G645), .O(gate275inter7));
  inv1  gate2039(.a(G797), .O(gate275inter8));
  nand2 gate2040(.a(gate275inter8), .b(gate275inter7), .O(gate275inter9));
  nand2 gate2041(.a(s_213), .b(gate275inter3), .O(gate275inter10));
  nor2  gate2042(.a(gate275inter10), .b(gate275inter9), .O(gate275inter11));
  nor2  gate2043(.a(gate275inter11), .b(gate275inter6), .O(gate275inter12));
  nand2 gate2044(.a(gate275inter12), .b(gate275inter1), .O(G820));
nand2 gate276( .a(G773), .b(G797), .O(G821) );
nand2 gate277( .a(G648), .b(G800), .O(G822) );

  xor2  gate1079(.a(G800), .b(G776), .O(gate278inter0));
  nand2 gate1080(.a(gate278inter0), .b(s_76), .O(gate278inter1));
  and2  gate1081(.a(G800), .b(G776), .O(gate278inter2));
  inv1  gate1082(.a(s_76), .O(gate278inter3));
  inv1  gate1083(.a(s_77), .O(gate278inter4));
  nand2 gate1084(.a(gate278inter4), .b(gate278inter3), .O(gate278inter5));
  nor2  gate1085(.a(gate278inter5), .b(gate278inter2), .O(gate278inter6));
  inv1  gate1086(.a(G776), .O(gate278inter7));
  inv1  gate1087(.a(G800), .O(gate278inter8));
  nand2 gate1088(.a(gate278inter8), .b(gate278inter7), .O(gate278inter9));
  nand2 gate1089(.a(s_77), .b(gate278inter3), .O(gate278inter10));
  nor2  gate1090(.a(gate278inter10), .b(gate278inter9), .O(gate278inter11));
  nor2  gate1091(.a(gate278inter11), .b(gate278inter6), .O(gate278inter12));
  nand2 gate1092(.a(gate278inter12), .b(gate278inter1), .O(G823));
nand2 gate279( .a(G651), .b(G803), .O(G824) );
nand2 gate280( .a(G779), .b(G803), .O(G825) );
nand2 gate281( .a(G654), .b(G806), .O(G826) );

  xor2  gate2367(.a(G806), .b(G782), .O(gate282inter0));
  nand2 gate2368(.a(gate282inter0), .b(s_260), .O(gate282inter1));
  and2  gate2369(.a(G806), .b(G782), .O(gate282inter2));
  inv1  gate2370(.a(s_260), .O(gate282inter3));
  inv1  gate2371(.a(s_261), .O(gate282inter4));
  nand2 gate2372(.a(gate282inter4), .b(gate282inter3), .O(gate282inter5));
  nor2  gate2373(.a(gate282inter5), .b(gate282inter2), .O(gate282inter6));
  inv1  gate2374(.a(G782), .O(gate282inter7));
  inv1  gate2375(.a(G806), .O(gate282inter8));
  nand2 gate2376(.a(gate282inter8), .b(gate282inter7), .O(gate282inter9));
  nand2 gate2377(.a(s_261), .b(gate282inter3), .O(gate282inter10));
  nor2  gate2378(.a(gate282inter10), .b(gate282inter9), .O(gate282inter11));
  nor2  gate2379(.a(gate282inter11), .b(gate282inter6), .O(gate282inter12));
  nand2 gate2380(.a(gate282inter12), .b(gate282inter1), .O(G827));
nand2 gate283( .a(G657), .b(G809), .O(G828) );
nand2 gate284( .a(G785), .b(G809), .O(G829) );

  xor2  gate1429(.a(G812), .b(G660), .O(gate285inter0));
  nand2 gate1430(.a(gate285inter0), .b(s_126), .O(gate285inter1));
  and2  gate1431(.a(G812), .b(G660), .O(gate285inter2));
  inv1  gate1432(.a(s_126), .O(gate285inter3));
  inv1  gate1433(.a(s_127), .O(gate285inter4));
  nand2 gate1434(.a(gate285inter4), .b(gate285inter3), .O(gate285inter5));
  nor2  gate1435(.a(gate285inter5), .b(gate285inter2), .O(gate285inter6));
  inv1  gate1436(.a(G660), .O(gate285inter7));
  inv1  gate1437(.a(G812), .O(gate285inter8));
  nand2 gate1438(.a(gate285inter8), .b(gate285inter7), .O(gate285inter9));
  nand2 gate1439(.a(s_127), .b(gate285inter3), .O(gate285inter10));
  nor2  gate1440(.a(gate285inter10), .b(gate285inter9), .O(gate285inter11));
  nor2  gate1441(.a(gate285inter11), .b(gate285inter6), .O(gate285inter12));
  nand2 gate1442(.a(gate285inter12), .b(gate285inter1), .O(G830));
nand2 gate286( .a(G788), .b(G812), .O(G831) );
nand2 gate287( .a(G663), .b(G815), .O(G832) );
nand2 gate288( .a(G791), .b(G815), .O(G833) );
nand2 gate289( .a(G818), .b(G819), .O(G834) );

  xor2  gate701(.a(G821), .b(G820), .O(gate290inter0));
  nand2 gate702(.a(gate290inter0), .b(s_22), .O(gate290inter1));
  and2  gate703(.a(G821), .b(G820), .O(gate290inter2));
  inv1  gate704(.a(s_22), .O(gate290inter3));
  inv1  gate705(.a(s_23), .O(gate290inter4));
  nand2 gate706(.a(gate290inter4), .b(gate290inter3), .O(gate290inter5));
  nor2  gate707(.a(gate290inter5), .b(gate290inter2), .O(gate290inter6));
  inv1  gate708(.a(G820), .O(gate290inter7));
  inv1  gate709(.a(G821), .O(gate290inter8));
  nand2 gate710(.a(gate290inter8), .b(gate290inter7), .O(gate290inter9));
  nand2 gate711(.a(s_23), .b(gate290inter3), .O(gate290inter10));
  nor2  gate712(.a(gate290inter10), .b(gate290inter9), .O(gate290inter11));
  nor2  gate713(.a(gate290inter11), .b(gate290inter6), .O(gate290inter12));
  nand2 gate714(.a(gate290inter12), .b(gate290inter1), .O(G847));

  xor2  gate2129(.a(G823), .b(G822), .O(gate291inter0));
  nand2 gate2130(.a(gate291inter0), .b(s_226), .O(gate291inter1));
  and2  gate2131(.a(G823), .b(G822), .O(gate291inter2));
  inv1  gate2132(.a(s_226), .O(gate291inter3));
  inv1  gate2133(.a(s_227), .O(gate291inter4));
  nand2 gate2134(.a(gate291inter4), .b(gate291inter3), .O(gate291inter5));
  nor2  gate2135(.a(gate291inter5), .b(gate291inter2), .O(gate291inter6));
  inv1  gate2136(.a(G822), .O(gate291inter7));
  inv1  gate2137(.a(G823), .O(gate291inter8));
  nand2 gate2138(.a(gate291inter8), .b(gate291inter7), .O(gate291inter9));
  nand2 gate2139(.a(s_227), .b(gate291inter3), .O(gate291inter10));
  nor2  gate2140(.a(gate291inter10), .b(gate291inter9), .O(gate291inter11));
  nor2  gate2141(.a(gate291inter11), .b(gate291inter6), .O(gate291inter12));
  nand2 gate2142(.a(gate291inter12), .b(gate291inter1), .O(G860));
nand2 gate292( .a(G824), .b(G825), .O(G873) );

  xor2  gate1303(.a(G829), .b(G828), .O(gate293inter0));
  nand2 gate1304(.a(gate293inter0), .b(s_108), .O(gate293inter1));
  and2  gate1305(.a(G829), .b(G828), .O(gate293inter2));
  inv1  gate1306(.a(s_108), .O(gate293inter3));
  inv1  gate1307(.a(s_109), .O(gate293inter4));
  nand2 gate1308(.a(gate293inter4), .b(gate293inter3), .O(gate293inter5));
  nor2  gate1309(.a(gate293inter5), .b(gate293inter2), .O(gate293inter6));
  inv1  gate1310(.a(G828), .O(gate293inter7));
  inv1  gate1311(.a(G829), .O(gate293inter8));
  nand2 gate1312(.a(gate293inter8), .b(gate293inter7), .O(gate293inter9));
  nand2 gate1313(.a(s_109), .b(gate293inter3), .O(gate293inter10));
  nor2  gate1314(.a(gate293inter10), .b(gate293inter9), .O(gate293inter11));
  nor2  gate1315(.a(gate293inter11), .b(gate293inter6), .O(gate293inter12));
  nand2 gate1316(.a(gate293inter12), .b(gate293inter1), .O(G886));
nand2 gate294( .a(G832), .b(G833), .O(G899) );
nand2 gate295( .a(G830), .b(G831), .O(G912) );
nand2 gate296( .a(G826), .b(G827), .O(G925) );
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );
nand2 gate387( .a(G1), .b(G1036), .O(G1132) );
nand2 gate388( .a(G2), .b(G1039), .O(G1135) );
nand2 gate389( .a(G3), .b(G1042), .O(G1138) );

  xor2  gate1107(.a(G1045), .b(G4), .O(gate390inter0));
  nand2 gate1108(.a(gate390inter0), .b(s_80), .O(gate390inter1));
  and2  gate1109(.a(G1045), .b(G4), .O(gate390inter2));
  inv1  gate1110(.a(s_80), .O(gate390inter3));
  inv1  gate1111(.a(s_81), .O(gate390inter4));
  nand2 gate1112(.a(gate390inter4), .b(gate390inter3), .O(gate390inter5));
  nor2  gate1113(.a(gate390inter5), .b(gate390inter2), .O(gate390inter6));
  inv1  gate1114(.a(G4), .O(gate390inter7));
  inv1  gate1115(.a(G1045), .O(gate390inter8));
  nand2 gate1116(.a(gate390inter8), .b(gate390inter7), .O(gate390inter9));
  nand2 gate1117(.a(s_81), .b(gate390inter3), .O(gate390inter10));
  nor2  gate1118(.a(gate390inter10), .b(gate390inter9), .O(gate390inter11));
  nor2  gate1119(.a(gate390inter11), .b(gate390inter6), .O(gate390inter12));
  nand2 gate1120(.a(gate390inter12), .b(gate390inter1), .O(G1141));
nand2 gate391( .a(G5), .b(G1048), .O(G1144) );

  xor2  gate1835(.a(G1051), .b(G6), .O(gate392inter0));
  nand2 gate1836(.a(gate392inter0), .b(s_184), .O(gate392inter1));
  and2  gate1837(.a(G1051), .b(G6), .O(gate392inter2));
  inv1  gate1838(.a(s_184), .O(gate392inter3));
  inv1  gate1839(.a(s_185), .O(gate392inter4));
  nand2 gate1840(.a(gate392inter4), .b(gate392inter3), .O(gate392inter5));
  nor2  gate1841(.a(gate392inter5), .b(gate392inter2), .O(gate392inter6));
  inv1  gate1842(.a(G6), .O(gate392inter7));
  inv1  gate1843(.a(G1051), .O(gate392inter8));
  nand2 gate1844(.a(gate392inter8), .b(gate392inter7), .O(gate392inter9));
  nand2 gate1845(.a(s_185), .b(gate392inter3), .O(gate392inter10));
  nor2  gate1846(.a(gate392inter10), .b(gate392inter9), .O(gate392inter11));
  nor2  gate1847(.a(gate392inter11), .b(gate392inter6), .O(gate392inter12));
  nand2 gate1848(.a(gate392inter12), .b(gate392inter1), .O(G1147));

  xor2  gate855(.a(G1054), .b(G7), .O(gate393inter0));
  nand2 gate856(.a(gate393inter0), .b(s_44), .O(gate393inter1));
  and2  gate857(.a(G1054), .b(G7), .O(gate393inter2));
  inv1  gate858(.a(s_44), .O(gate393inter3));
  inv1  gate859(.a(s_45), .O(gate393inter4));
  nand2 gate860(.a(gate393inter4), .b(gate393inter3), .O(gate393inter5));
  nor2  gate861(.a(gate393inter5), .b(gate393inter2), .O(gate393inter6));
  inv1  gate862(.a(G7), .O(gate393inter7));
  inv1  gate863(.a(G1054), .O(gate393inter8));
  nand2 gate864(.a(gate393inter8), .b(gate393inter7), .O(gate393inter9));
  nand2 gate865(.a(s_45), .b(gate393inter3), .O(gate393inter10));
  nor2  gate866(.a(gate393inter10), .b(gate393inter9), .O(gate393inter11));
  nor2  gate867(.a(gate393inter11), .b(gate393inter6), .O(gate393inter12));
  nand2 gate868(.a(gate393inter12), .b(gate393inter1), .O(G1150));
nand2 gate394( .a(G8), .b(G1057), .O(G1153) );
nand2 gate395( .a(G9), .b(G1060), .O(G1156) );
nand2 gate396( .a(G10), .b(G1063), .O(G1159) );

  xor2  gate1555(.a(G1066), .b(G11), .O(gate397inter0));
  nand2 gate1556(.a(gate397inter0), .b(s_144), .O(gate397inter1));
  and2  gate1557(.a(G1066), .b(G11), .O(gate397inter2));
  inv1  gate1558(.a(s_144), .O(gate397inter3));
  inv1  gate1559(.a(s_145), .O(gate397inter4));
  nand2 gate1560(.a(gate397inter4), .b(gate397inter3), .O(gate397inter5));
  nor2  gate1561(.a(gate397inter5), .b(gate397inter2), .O(gate397inter6));
  inv1  gate1562(.a(G11), .O(gate397inter7));
  inv1  gate1563(.a(G1066), .O(gate397inter8));
  nand2 gate1564(.a(gate397inter8), .b(gate397inter7), .O(gate397inter9));
  nand2 gate1565(.a(s_145), .b(gate397inter3), .O(gate397inter10));
  nor2  gate1566(.a(gate397inter10), .b(gate397inter9), .O(gate397inter11));
  nor2  gate1567(.a(gate397inter11), .b(gate397inter6), .O(gate397inter12));
  nand2 gate1568(.a(gate397inter12), .b(gate397inter1), .O(G1162));

  xor2  gate2115(.a(G1069), .b(G12), .O(gate398inter0));
  nand2 gate2116(.a(gate398inter0), .b(s_224), .O(gate398inter1));
  and2  gate2117(.a(G1069), .b(G12), .O(gate398inter2));
  inv1  gate2118(.a(s_224), .O(gate398inter3));
  inv1  gate2119(.a(s_225), .O(gate398inter4));
  nand2 gate2120(.a(gate398inter4), .b(gate398inter3), .O(gate398inter5));
  nor2  gate2121(.a(gate398inter5), .b(gate398inter2), .O(gate398inter6));
  inv1  gate2122(.a(G12), .O(gate398inter7));
  inv1  gate2123(.a(G1069), .O(gate398inter8));
  nand2 gate2124(.a(gate398inter8), .b(gate398inter7), .O(gate398inter9));
  nand2 gate2125(.a(s_225), .b(gate398inter3), .O(gate398inter10));
  nor2  gate2126(.a(gate398inter10), .b(gate398inter9), .O(gate398inter11));
  nor2  gate2127(.a(gate398inter11), .b(gate398inter6), .O(gate398inter12));
  nand2 gate2128(.a(gate398inter12), .b(gate398inter1), .O(G1165));
nand2 gate399( .a(G13), .b(G1072), .O(G1168) );
nand2 gate400( .a(G14), .b(G1075), .O(G1171) );

  xor2  gate1247(.a(G1078), .b(G15), .O(gate401inter0));
  nand2 gate1248(.a(gate401inter0), .b(s_100), .O(gate401inter1));
  and2  gate1249(.a(G1078), .b(G15), .O(gate401inter2));
  inv1  gate1250(.a(s_100), .O(gate401inter3));
  inv1  gate1251(.a(s_101), .O(gate401inter4));
  nand2 gate1252(.a(gate401inter4), .b(gate401inter3), .O(gate401inter5));
  nor2  gate1253(.a(gate401inter5), .b(gate401inter2), .O(gate401inter6));
  inv1  gate1254(.a(G15), .O(gate401inter7));
  inv1  gate1255(.a(G1078), .O(gate401inter8));
  nand2 gate1256(.a(gate401inter8), .b(gate401inter7), .O(gate401inter9));
  nand2 gate1257(.a(s_101), .b(gate401inter3), .O(gate401inter10));
  nor2  gate1258(.a(gate401inter10), .b(gate401inter9), .O(gate401inter11));
  nor2  gate1259(.a(gate401inter11), .b(gate401inter6), .O(gate401inter12));
  nand2 gate1260(.a(gate401inter12), .b(gate401inter1), .O(G1174));

  xor2  gate2045(.a(G1081), .b(G16), .O(gate402inter0));
  nand2 gate2046(.a(gate402inter0), .b(s_214), .O(gate402inter1));
  and2  gate2047(.a(G1081), .b(G16), .O(gate402inter2));
  inv1  gate2048(.a(s_214), .O(gate402inter3));
  inv1  gate2049(.a(s_215), .O(gate402inter4));
  nand2 gate2050(.a(gate402inter4), .b(gate402inter3), .O(gate402inter5));
  nor2  gate2051(.a(gate402inter5), .b(gate402inter2), .O(gate402inter6));
  inv1  gate2052(.a(G16), .O(gate402inter7));
  inv1  gate2053(.a(G1081), .O(gate402inter8));
  nand2 gate2054(.a(gate402inter8), .b(gate402inter7), .O(gate402inter9));
  nand2 gate2055(.a(s_215), .b(gate402inter3), .O(gate402inter10));
  nor2  gate2056(.a(gate402inter10), .b(gate402inter9), .O(gate402inter11));
  nor2  gate2057(.a(gate402inter11), .b(gate402inter6), .O(gate402inter12));
  nand2 gate2058(.a(gate402inter12), .b(gate402inter1), .O(G1177));
nand2 gate403( .a(G17), .b(G1084), .O(G1180) );
nand2 gate404( .a(G18), .b(G1087), .O(G1183) );

  xor2  gate2003(.a(G1090), .b(G19), .O(gate405inter0));
  nand2 gate2004(.a(gate405inter0), .b(s_208), .O(gate405inter1));
  and2  gate2005(.a(G1090), .b(G19), .O(gate405inter2));
  inv1  gate2006(.a(s_208), .O(gate405inter3));
  inv1  gate2007(.a(s_209), .O(gate405inter4));
  nand2 gate2008(.a(gate405inter4), .b(gate405inter3), .O(gate405inter5));
  nor2  gate2009(.a(gate405inter5), .b(gate405inter2), .O(gate405inter6));
  inv1  gate2010(.a(G19), .O(gate405inter7));
  inv1  gate2011(.a(G1090), .O(gate405inter8));
  nand2 gate2012(.a(gate405inter8), .b(gate405inter7), .O(gate405inter9));
  nand2 gate2013(.a(s_209), .b(gate405inter3), .O(gate405inter10));
  nor2  gate2014(.a(gate405inter10), .b(gate405inter9), .O(gate405inter11));
  nor2  gate2015(.a(gate405inter11), .b(gate405inter6), .O(gate405inter12));
  nand2 gate2016(.a(gate405inter12), .b(gate405inter1), .O(G1186));

  xor2  gate687(.a(G1093), .b(G20), .O(gate406inter0));
  nand2 gate688(.a(gate406inter0), .b(s_20), .O(gate406inter1));
  and2  gate689(.a(G1093), .b(G20), .O(gate406inter2));
  inv1  gate690(.a(s_20), .O(gate406inter3));
  inv1  gate691(.a(s_21), .O(gate406inter4));
  nand2 gate692(.a(gate406inter4), .b(gate406inter3), .O(gate406inter5));
  nor2  gate693(.a(gate406inter5), .b(gate406inter2), .O(gate406inter6));
  inv1  gate694(.a(G20), .O(gate406inter7));
  inv1  gate695(.a(G1093), .O(gate406inter8));
  nand2 gate696(.a(gate406inter8), .b(gate406inter7), .O(gate406inter9));
  nand2 gate697(.a(s_21), .b(gate406inter3), .O(gate406inter10));
  nor2  gate698(.a(gate406inter10), .b(gate406inter9), .O(gate406inter11));
  nor2  gate699(.a(gate406inter11), .b(gate406inter6), .O(gate406inter12));
  nand2 gate700(.a(gate406inter12), .b(gate406inter1), .O(G1189));
nand2 gate407( .a(G21), .b(G1096), .O(G1192) );
nand2 gate408( .a(G22), .b(G1099), .O(G1195) );

  xor2  gate981(.a(G1102), .b(G23), .O(gate409inter0));
  nand2 gate982(.a(gate409inter0), .b(s_62), .O(gate409inter1));
  and2  gate983(.a(G1102), .b(G23), .O(gate409inter2));
  inv1  gate984(.a(s_62), .O(gate409inter3));
  inv1  gate985(.a(s_63), .O(gate409inter4));
  nand2 gate986(.a(gate409inter4), .b(gate409inter3), .O(gate409inter5));
  nor2  gate987(.a(gate409inter5), .b(gate409inter2), .O(gate409inter6));
  inv1  gate988(.a(G23), .O(gate409inter7));
  inv1  gate989(.a(G1102), .O(gate409inter8));
  nand2 gate990(.a(gate409inter8), .b(gate409inter7), .O(gate409inter9));
  nand2 gate991(.a(s_63), .b(gate409inter3), .O(gate409inter10));
  nor2  gate992(.a(gate409inter10), .b(gate409inter9), .O(gate409inter11));
  nor2  gate993(.a(gate409inter11), .b(gate409inter6), .O(gate409inter12));
  nand2 gate994(.a(gate409inter12), .b(gate409inter1), .O(G1198));
nand2 gate410( .a(G24), .b(G1105), .O(G1201) );
nand2 gate411( .a(G25), .b(G1108), .O(G1204) );
nand2 gate412( .a(G26), .b(G1111), .O(G1207) );

  xor2  gate2283(.a(G1114), .b(G27), .O(gate413inter0));
  nand2 gate2284(.a(gate413inter0), .b(s_248), .O(gate413inter1));
  and2  gate2285(.a(G1114), .b(G27), .O(gate413inter2));
  inv1  gate2286(.a(s_248), .O(gate413inter3));
  inv1  gate2287(.a(s_249), .O(gate413inter4));
  nand2 gate2288(.a(gate413inter4), .b(gate413inter3), .O(gate413inter5));
  nor2  gate2289(.a(gate413inter5), .b(gate413inter2), .O(gate413inter6));
  inv1  gate2290(.a(G27), .O(gate413inter7));
  inv1  gate2291(.a(G1114), .O(gate413inter8));
  nand2 gate2292(.a(gate413inter8), .b(gate413inter7), .O(gate413inter9));
  nand2 gate2293(.a(s_249), .b(gate413inter3), .O(gate413inter10));
  nor2  gate2294(.a(gate413inter10), .b(gate413inter9), .O(gate413inter11));
  nor2  gate2295(.a(gate413inter11), .b(gate413inter6), .O(gate413inter12));
  nand2 gate2296(.a(gate413inter12), .b(gate413inter1), .O(G1210));

  xor2  gate883(.a(G1117), .b(G28), .O(gate414inter0));
  nand2 gate884(.a(gate414inter0), .b(s_48), .O(gate414inter1));
  and2  gate885(.a(G1117), .b(G28), .O(gate414inter2));
  inv1  gate886(.a(s_48), .O(gate414inter3));
  inv1  gate887(.a(s_49), .O(gate414inter4));
  nand2 gate888(.a(gate414inter4), .b(gate414inter3), .O(gate414inter5));
  nor2  gate889(.a(gate414inter5), .b(gate414inter2), .O(gate414inter6));
  inv1  gate890(.a(G28), .O(gate414inter7));
  inv1  gate891(.a(G1117), .O(gate414inter8));
  nand2 gate892(.a(gate414inter8), .b(gate414inter7), .O(gate414inter9));
  nand2 gate893(.a(s_49), .b(gate414inter3), .O(gate414inter10));
  nor2  gate894(.a(gate414inter10), .b(gate414inter9), .O(gate414inter11));
  nor2  gate895(.a(gate414inter11), .b(gate414inter6), .O(gate414inter12));
  nand2 gate896(.a(gate414inter12), .b(gate414inter1), .O(G1213));
nand2 gate415( .a(G29), .b(G1120), .O(G1216) );

  xor2  gate1779(.a(G1123), .b(G30), .O(gate416inter0));
  nand2 gate1780(.a(gate416inter0), .b(s_176), .O(gate416inter1));
  and2  gate1781(.a(G1123), .b(G30), .O(gate416inter2));
  inv1  gate1782(.a(s_176), .O(gate416inter3));
  inv1  gate1783(.a(s_177), .O(gate416inter4));
  nand2 gate1784(.a(gate416inter4), .b(gate416inter3), .O(gate416inter5));
  nor2  gate1785(.a(gate416inter5), .b(gate416inter2), .O(gate416inter6));
  inv1  gate1786(.a(G30), .O(gate416inter7));
  inv1  gate1787(.a(G1123), .O(gate416inter8));
  nand2 gate1788(.a(gate416inter8), .b(gate416inter7), .O(gate416inter9));
  nand2 gate1789(.a(s_177), .b(gate416inter3), .O(gate416inter10));
  nor2  gate1790(.a(gate416inter10), .b(gate416inter9), .O(gate416inter11));
  nor2  gate1791(.a(gate416inter11), .b(gate416inter6), .O(gate416inter12));
  nand2 gate1792(.a(gate416inter12), .b(gate416inter1), .O(G1219));
nand2 gate417( .a(G31), .b(G1126), .O(G1222) );
nand2 gate418( .a(G32), .b(G1129), .O(G1225) );
nand2 gate419( .a(G1), .b(G1132), .O(G1228) );

  xor2  gate995(.a(G1132), .b(G1036), .O(gate420inter0));
  nand2 gate996(.a(gate420inter0), .b(s_64), .O(gate420inter1));
  and2  gate997(.a(G1132), .b(G1036), .O(gate420inter2));
  inv1  gate998(.a(s_64), .O(gate420inter3));
  inv1  gate999(.a(s_65), .O(gate420inter4));
  nand2 gate1000(.a(gate420inter4), .b(gate420inter3), .O(gate420inter5));
  nor2  gate1001(.a(gate420inter5), .b(gate420inter2), .O(gate420inter6));
  inv1  gate1002(.a(G1036), .O(gate420inter7));
  inv1  gate1003(.a(G1132), .O(gate420inter8));
  nand2 gate1004(.a(gate420inter8), .b(gate420inter7), .O(gate420inter9));
  nand2 gate1005(.a(s_65), .b(gate420inter3), .O(gate420inter10));
  nor2  gate1006(.a(gate420inter10), .b(gate420inter9), .O(gate420inter11));
  nor2  gate1007(.a(gate420inter11), .b(gate420inter6), .O(gate420inter12));
  nand2 gate1008(.a(gate420inter12), .b(gate420inter1), .O(G1229));
nand2 gate421( .a(G2), .b(G1135), .O(G1230) );
nand2 gate422( .a(G1039), .b(G1135), .O(G1231) );
nand2 gate423( .a(G3), .b(G1138), .O(G1232) );
nand2 gate424( .a(G1042), .b(G1138), .O(G1233) );
nand2 gate425( .a(G4), .b(G1141), .O(G1234) );

  xor2  gate1233(.a(G1141), .b(G1045), .O(gate426inter0));
  nand2 gate1234(.a(gate426inter0), .b(s_98), .O(gate426inter1));
  and2  gate1235(.a(G1141), .b(G1045), .O(gate426inter2));
  inv1  gate1236(.a(s_98), .O(gate426inter3));
  inv1  gate1237(.a(s_99), .O(gate426inter4));
  nand2 gate1238(.a(gate426inter4), .b(gate426inter3), .O(gate426inter5));
  nor2  gate1239(.a(gate426inter5), .b(gate426inter2), .O(gate426inter6));
  inv1  gate1240(.a(G1045), .O(gate426inter7));
  inv1  gate1241(.a(G1141), .O(gate426inter8));
  nand2 gate1242(.a(gate426inter8), .b(gate426inter7), .O(gate426inter9));
  nand2 gate1243(.a(s_99), .b(gate426inter3), .O(gate426inter10));
  nor2  gate1244(.a(gate426inter10), .b(gate426inter9), .O(gate426inter11));
  nor2  gate1245(.a(gate426inter11), .b(gate426inter6), .O(gate426inter12));
  nand2 gate1246(.a(gate426inter12), .b(gate426inter1), .O(G1235));

  xor2  gate2241(.a(G1144), .b(G5), .O(gate427inter0));
  nand2 gate2242(.a(gate427inter0), .b(s_242), .O(gate427inter1));
  and2  gate2243(.a(G1144), .b(G5), .O(gate427inter2));
  inv1  gate2244(.a(s_242), .O(gate427inter3));
  inv1  gate2245(.a(s_243), .O(gate427inter4));
  nand2 gate2246(.a(gate427inter4), .b(gate427inter3), .O(gate427inter5));
  nor2  gate2247(.a(gate427inter5), .b(gate427inter2), .O(gate427inter6));
  inv1  gate2248(.a(G5), .O(gate427inter7));
  inv1  gate2249(.a(G1144), .O(gate427inter8));
  nand2 gate2250(.a(gate427inter8), .b(gate427inter7), .O(gate427inter9));
  nand2 gate2251(.a(s_243), .b(gate427inter3), .O(gate427inter10));
  nor2  gate2252(.a(gate427inter10), .b(gate427inter9), .O(gate427inter11));
  nor2  gate2253(.a(gate427inter11), .b(gate427inter6), .O(gate427inter12));
  nand2 gate2254(.a(gate427inter12), .b(gate427inter1), .O(G1236));
nand2 gate428( .a(G1048), .b(G1144), .O(G1237) );
nand2 gate429( .a(G6), .b(G1147), .O(G1238) );

  xor2  gate2157(.a(G1147), .b(G1051), .O(gate430inter0));
  nand2 gate2158(.a(gate430inter0), .b(s_230), .O(gate430inter1));
  and2  gate2159(.a(G1147), .b(G1051), .O(gate430inter2));
  inv1  gate2160(.a(s_230), .O(gate430inter3));
  inv1  gate2161(.a(s_231), .O(gate430inter4));
  nand2 gate2162(.a(gate430inter4), .b(gate430inter3), .O(gate430inter5));
  nor2  gate2163(.a(gate430inter5), .b(gate430inter2), .O(gate430inter6));
  inv1  gate2164(.a(G1051), .O(gate430inter7));
  inv1  gate2165(.a(G1147), .O(gate430inter8));
  nand2 gate2166(.a(gate430inter8), .b(gate430inter7), .O(gate430inter9));
  nand2 gate2167(.a(s_231), .b(gate430inter3), .O(gate430inter10));
  nor2  gate2168(.a(gate430inter10), .b(gate430inter9), .O(gate430inter11));
  nor2  gate2169(.a(gate430inter11), .b(gate430inter6), .O(gate430inter12));
  nand2 gate2170(.a(gate430inter12), .b(gate430inter1), .O(G1239));

  xor2  gate2199(.a(G1150), .b(G7), .O(gate431inter0));
  nand2 gate2200(.a(gate431inter0), .b(s_236), .O(gate431inter1));
  and2  gate2201(.a(G1150), .b(G7), .O(gate431inter2));
  inv1  gate2202(.a(s_236), .O(gate431inter3));
  inv1  gate2203(.a(s_237), .O(gate431inter4));
  nand2 gate2204(.a(gate431inter4), .b(gate431inter3), .O(gate431inter5));
  nor2  gate2205(.a(gate431inter5), .b(gate431inter2), .O(gate431inter6));
  inv1  gate2206(.a(G7), .O(gate431inter7));
  inv1  gate2207(.a(G1150), .O(gate431inter8));
  nand2 gate2208(.a(gate431inter8), .b(gate431inter7), .O(gate431inter9));
  nand2 gate2209(.a(s_237), .b(gate431inter3), .O(gate431inter10));
  nor2  gate2210(.a(gate431inter10), .b(gate431inter9), .O(gate431inter11));
  nor2  gate2211(.a(gate431inter11), .b(gate431inter6), .O(gate431inter12));
  nand2 gate2212(.a(gate431inter12), .b(gate431inter1), .O(G1240));
nand2 gate432( .a(G1054), .b(G1150), .O(G1241) );

  xor2  gate2255(.a(G1153), .b(G8), .O(gate433inter0));
  nand2 gate2256(.a(gate433inter0), .b(s_244), .O(gate433inter1));
  and2  gate2257(.a(G1153), .b(G8), .O(gate433inter2));
  inv1  gate2258(.a(s_244), .O(gate433inter3));
  inv1  gate2259(.a(s_245), .O(gate433inter4));
  nand2 gate2260(.a(gate433inter4), .b(gate433inter3), .O(gate433inter5));
  nor2  gate2261(.a(gate433inter5), .b(gate433inter2), .O(gate433inter6));
  inv1  gate2262(.a(G8), .O(gate433inter7));
  inv1  gate2263(.a(G1153), .O(gate433inter8));
  nand2 gate2264(.a(gate433inter8), .b(gate433inter7), .O(gate433inter9));
  nand2 gate2265(.a(s_245), .b(gate433inter3), .O(gate433inter10));
  nor2  gate2266(.a(gate433inter10), .b(gate433inter9), .O(gate433inter11));
  nor2  gate2267(.a(gate433inter11), .b(gate433inter6), .O(gate433inter12));
  nand2 gate2268(.a(gate433inter12), .b(gate433inter1), .O(G1242));
nand2 gate434( .a(G1057), .b(G1153), .O(G1243) );
nand2 gate435( .a(G9), .b(G1156), .O(G1244) );
nand2 gate436( .a(G1060), .b(G1156), .O(G1245) );
nand2 gate437( .a(G10), .b(G1159), .O(G1246) );

  xor2  gate645(.a(G1159), .b(G1063), .O(gate438inter0));
  nand2 gate646(.a(gate438inter0), .b(s_14), .O(gate438inter1));
  and2  gate647(.a(G1159), .b(G1063), .O(gate438inter2));
  inv1  gate648(.a(s_14), .O(gate438inter3));
  inv1  gate649(.a(s_15), .O(gate438inter4));
  nand2 gate650(.a(gate438inter4), .b(gate438inter3), .O(gate438inter5));
  nor2  gate651(.a(gate438inter5), .b(gate438inter2), .O(gate438inter6));
  inv1  gate652(.a(G1063), .O(gate438inter7));
  inv1  gate653(.a(G1159), .O(gate438inter8));
  nand2 gate654(.a(gate438inter8), .b(gate438inter7), .O(gate438inter9));
  nand2 gate655(.a(s_15), .b(gate438inter3), .O(gate438inter10));
  nor2  gate656(.a(gate438inter10), .b(gate438inter9), .O(gate438inter11));
  nor2  gate657(.a(gate438inter11), .b(gate438inter6), .O(gate438inter12));
  nand2 gate658(.a(gate438inter12), .b(gate438inter1), .O(G1247));
nand2 gate439( .a(G11), .b(G1162), .O(G1248) );
nand2 gate440( .a(G1066), .b(G1162), .O(G1249) );

  xor2  gate1219(.a(G1165), .b(G12), .O(gate441inter0));
  nand2 gate1220(.a(gate441inter0), .b(s_96), .O(gate441inter1));
  and2  gate1221(.a(G1165), .b(G12), .O(gate441inter2));
  inv1  gate1222(.a(s_96), .O(gate441inter3));
  inv1  gate1223(.a(s_97), .O(gate441inter4));
  nand2 gate1224(.a(gate441inter4), .b(gate441inter3), .O(gate441inter5));
  nor2  gate1225(.a(gate441inter5), .b(gate441inter2), .O(gate441inter6));
  inv1  gate1226(.a(G12), .O(gate441inter7));
  inv1  gate1227(.a(G1165), .O(gate441inter8));
  nand2 gate1228(.a(gate441inter8), .b(gate441inter7), .O(gate441inter9));
  nand2 gate1229(.a(s_97), .b(gate441inter3), .O(gate441inter10));
  nor2  gate1230(.a(gate441inter10), .b(gate441inter9), .O(gate441inter11));
  nor2  gate1231(.a(gate441inter11), .b(gate441inter6), .O(gate441inter12));
  nand2 gate1232(.a(gate441inter12), .b(gate441inter1), .O(G1250));
nand2 gate442( .a(G1069), .b(G1165), .O(G1251) );
nand2 gate443( .a(G13), .b(G1168), .O(G1252) );
nand2 gate444( .a(G1072), .b(G1168), .O(G1253) );
nand2 gate445( .a(G14), .b(G1171), .O(G1254) );
nand2 gate446( .a(G1075), .b(G1171), .O(G1255) );
nand2 gate447( .a(G15), .b(G1174), .O(G1256) );
nand2 gate448( .a(G1078), .b(G1174), .O(G1257) );
nand2 gate449( .a(G16), .b(G1177), .O(G1258) );
nand2 gate450( .a(G1081), .b(G1177), .O(G1259) );
nand2 gate451( .a(G17), .b(G1180), .O(G1260) );
nand2 gate452( .a(G1084), .b(G1180), .O(G1261) );
nand2 gate453( .a(G18), .b(G1183), .O(G1262) );

  xor2  gate1191(.a(G1183), .b(G1087), .O(gate454inter0));
  nand2 gate1192(.a(gate454inter0), .b(s_92), .O(gate454inter1));
  and2  gate1193(.a(G1183), .b(G1087), .O(gate454inter2));
  inv1  gate1194(.a(s_92), .O(gate454inter3));
  inv1  gate1195(.a(s_93), .O(gate454inter4));
  nand2 gate1196(.a(gate454inter4), .b(gate454inter3), .O(gate454inter5));
  nor2  gate1197(.a(gate454inter5), .b(gate454inter2), .O(gate454inter6));
  inv1  gate1198(.a(G1087), .O(gate454inter7));
  inv1  gate1199(.a(G1183), .O(gate454inter8));
  nand2 gate1200(.a(gate454inter8), .b(gate454inter7), .O(gate454inter9));
  nand2 gate1201(.a(s_93), .b(gate454inter3), .O(gate454inter10));
  nor2  gate1202(.a(gate454inter10), .b(gate454inter9), .O(gate454inter11));
  nor2  gate1203(.a(gate454inter11), .b(gate454inter6), .O(gate454inter12));
  nand2 gate1204(.a(gate454inter12), .b(gate454inter1), .O(G1263));

  xor2  gate1737(.a(G1186), .b(G19), .O(gate455inter0));
  nand2 gate1738(.a(gate455inter0), .b(s_170), .O(gate455inter1));
  and2  gate1739(.a(G1186), .b(G19), .O(gate455inter2));
  inv1  gate1740(.a(s_170), .O(gate455inter3));
  inv1  gate1741(.a(s_171), .O(gate455inter4));
  nand2 gate1742(.a(gate455inter4), .b(gate455inter3), .O(gate455inter5));
  nor2  gate1743(.a(gate455inter5), .b(gate455inter2), .O(gate455inter6));
  inv1  gate1744(.a(G19), .O(gate455inter7));
  inv1  gate1745(.a(G1186), .O(gate455inter8));
  nand2 gate1746(.a(gate455inter8), .b(gate455inter7), .O(gate455inter9));
  nand2 gate1747(.a(s_171), .b(gate455inter3), .O(gate455inter10));
  nor2  gate1748(.a(gate455inter10), .b(gate455inter9), .O(gate455inter11));
  nor2  gate1749(.a(gate455inter11), .b(gate455inter6), .O(gate455inter12));
  nand2 gate1750(.a(gate455inter12), .b(gate455inter1), .O(G1264));
nand2 gate456( .a(G1090), .b(G1186), .O(G1265) );
nand2 gate457( .a(G20), .b(G1189), .O(G1266) );
nand2 gate458( .a(G1093), .b(G1189), .O(G1267) );
nand2 gate459( .a(G21), .b(G1192), .O(G1268) );

  xor2  gate925(.a(G1192), .b(G1096), .O(gate460inter0));
  nand2 gate926(.a(gate460inter0), .b(s_54), .O(gate460inter1));
  and2  gate927(.a(G1192), .b(G1096), .O(gate460inter2));
  inv1  gate928(.a(s_54), .O(gate460inter3));
  inv1  gate929(.a(s_55), .O(gate460inter4));
  nand2 gate930(.a(gate460inter4), .b(gate460inter3), .O(gate460inter5));
  nor2  gate931(.a(gate460inter5), .b(gate460inter2), .O(gate460inter6));
  inv1  gate932(.a(G1096), .O(gate460inter7));
  inv1  gate933(.a(G1192), .O(gate460inter8));
  nand2 gate934(.a(gate460inter8), .b(gate460inter7), .O(gate460inter9));
  nand2 gate935(.a(s_55), .b(gate460inter3), .O(gate460inter10));
  nor2  gate936(.a(gate460inter10), .b(gate460inter9), .O(gate460inter11));
  nor2  gate937(.a(gate460inter11), .b(gate460inter6), .O(gate460inter12));
  nand2 gate938(.a(gate460inter12), .b(gate460inter1), .O(G1269));
nand2 gate461( .a(G22), .b(G1195), .O(G1270) );
nand2 gate462( .a(G1099), .b(G1195), .O(G1271) );
nand2 gate463( .a(G23), .b(G1198), .O(G1272) );
nand2 gate464( .a(G1102), .b(G1198), .O(G1273) );

  xor2  gate1499(.a(G1201), .b(G24), .O(gate465inter0));
  nand2 gate1500(.a(gate465inter0), .b(s_136), .O(gate465inter1));
  and2  gate1501(.a(G1201), .b(G24), .O(gate465inter2));
  inv1  gate1502(.a(s_136), .O(gate465inter3));
  inv1  gate1503(.a(s_137), .O(gate465inter4));
  nand2 gate1504(.a(gate465inter4), .b(gate465inter3), .O(gate465inter5));
  nor2  gate1505(.a(gate465inter5), .b(gate465inter2), .O(gate465inter6));
  inv1  gate1506(.a(G24), .O(gate465inter7));
  inv1  gate1507(.a(G1201), .O(gate465inter8));
  nand2 gate1508(.a(gate465inter8), .b(gate465inter7), .O(gate465inter9));
  nand2 gate1509(.a(s_137), .b(gate465inter3), .O(gate465inter10));
  nor2  gate1510(.a(gate465inter10), .b(gate465inter9), .O(gate465inter11));
  nor2  gate1511(.a(gate465inter11), .b(gate465inter6), .O(gate465inter12));
  nand2 gate1512(.a(gate465inter12), .b(gate465inter1), .O(G1274));

  xor2  gate1135(.a(G1201), .b(G1105), .O(gate466inter0));
  nand2 gate1136(.a(gate466inter0), .b(s_84), .O(gate466inter1));
  and2  gate1137(.a(G1201), .b(G1105), .O(gate466inter2));
  inv1  gate1138(.a(s_84), .O(gate466inter3));
  inv1  gate1139(.a(s_85), .O(gate466inter4));
  nand2 gate1140(.a(gate466inter4), .b(gate466inter3), .O(gate466inter5));
  nor2  gate1141(.a(gate466inter5), .b(gate466inter2), .O(gate466inter6));
  inv1  gate1142(.a(G1105), .O(gate466inter7));
  inv1  gate1143(.a(G1201), .O(gate466inter8));
  nand2 gate1144(.a(gate466inter8), .b(gate466inter7), .O(gate466inter9));
  nand2 gate1145(.a(s_85), .b(gate466inter3), .O(gate466inter10));
  nor2  gate1146(.a(gate466inter10), .b(gate466inter9), .O(gate466inter11));
  nor2  gate1147(.a(gate466inter11), .b(gate466inter6), .O(gate466inter12));
  nand2 gate1148(.a(gate466inter12), .b(gate466inter1), .O(G1275));

  xor2  gate2059(.a(G1204), .b(G25), .O(gate467inter0));
  nand2 gate2060(.a(gate467inter0), .b(s_216), .O(gate467inter1));
  and2  gate2061(.a(G1204), .b(G25), .O(gate467inter2));
  inv1  gate2062(.a(s_216), .O(gate467inter3));
  inv1  gate2063(.a(s_217), .O(gate467inter4));
  nand2 gate2064(.a(gate467inter4), .b(gate467inter3), .O(gate467inter5));
  nor2  gate2065(.a(gate467inter5), .b(gate467inter2), .O(gate467inter6));
  inv1  gate2066(.a(G25), .O(gate467inter7));
  inv1  gate2067(.a(G1204), .O(gate467inter8));
  nand2 gate2068(.a(gate467inter8), .b(gate467inter7), .O(gate467inter9));
  nand2 gate2069(.a(s_217), .b(gate467inter3), .O(gate467inter10));
  nor2  gate2070(.a(gate467inter10), .b(gate467inter9), .O(gate467inter11));
  nor2  gate2071(.a(gate467inter11), .b(gate467inter6), .O(gate467inter12));
  nand2 gate2072(.a(gate467inter12), .b(gate467inter1), .O(G1276));
nand2 gate468( .a(G1108), .b(G1204), .O(G1277) );
nand2 gate469( .a(G26), .b(G1207), .O(G1278) );
nand2 gate470( .a(G1111), .b(G1207), .O(G1279) );
nand2 gate471( .a(G27), .b(G1210), .O(G1280) );

  xor2  gate757(.a(G1210), .b(G1114), .O(gate472inter0));
  nand2 gate758(.a(gate472inter0), .b(s_30), .O(gate472inter1));
  and2  gate759(.a(G1210), .b(G1114), .O(gate472inter2));
  inv1  gate760(.a(s_30), .O(gate472inter3));
  inv1  gate761(.a(s_31), .O(gate472inter4));
  nand2 gate762(.a(gate472inter4), .b(gate472inter3), .O(gate472inter5));
  nor2  gate763(.a(gate472inter5), .b(gate472inter2), .O(gate472inter6));
  inv1  gate764(.a(G1114), .O(gate472inter7));
  inv1  gate765(.a(G1210), .O(gate472inter8));
  nand2 gate766(.a(gate472inter8), .b(gate472inter7), .O(gate472inter9));
  nand2 gate767(.a(s_31), .b(gate472inter3), .O(gate472inter10));
  nor2  gate768(.a(gate472inter10), .b(gate472inter9), .O(gate472inter11));
  nor2  gate769(.a(gate472inter11), .b(gate472inter6), .O(gate472inter12));
  nand2 gate770(.a(gate472inter12), .b(gate472inter1), .O(G1281));

  xor2  gate785(.a(G1213), .b(G28), .O(gate473inter0));
  nand2 gate786(.a(gate473inter0), .b(s_34), .O(gate473inter1));
  and2  gate787(.a(G1213), .b(G28), .O(gate473inter2));
  inv1  gate788(.a(s_34), .O(gate473inter3));
  inv1  gate789(.a(s_35), .O(gate473inter4));
  nand2 gate790(.a(gate473inter4), .b(gate473inter3), .O(gate473inter5));
  nor2  gate791(.a(gate473inter5), .b(gate473inter2), .O(gate473inter6));
  inv1  gate792(.a(G28), .O(gate473inter7));
  inv1  gate793(.a(G1213), .O(gate473inter8));
  nand2 gate794(.a(gate473inter8), .b(gate473inter7), .O(gate473inter9));
  nand2 gate795(.a(s_35), .b(gate473inter3), .O(gate473inter10));
  nor2  gate796(.a(gate473inter10), .b(gate473inter9), .O(gate473inter11));
  nor2  gate797(.a(gate473inter11), .b(gate473inter6), .O(gate473inter12));
  nand2 gate798(.a(gate473inter12), .b(gate473inter1), .O(G1282));
nand2 gate474( .a(G1117), .b(G1213), .O(G1283) );
nand2 gate475( .a(G29), .b(G1216), .O(G1284) );
nand2 gate476( .a(G1120), .b(G1216), .O(G1285) );
nand2 gate477( .a(G30), .b(G1219), .O(G1286) );
nand2 gate478( .a(G1123), .b(G1219), .O(G1287) );
nand2 gate479( .a(G31), .b(G1222), .O(G1288) );
nand2 gate480( .a(G1126), .b(G1222), .O(G1289) );
nand2 gate481( .a(G32), .b(G1225), .O(G1290) );
nand2 gate482( .a(G1129), .b(G1225), .O(G1291) );
nand2 gate483( .a(G1228), .b(G1229), .O(G1292) );
nand2 gate484( .a(G1230), .b(G1231), .O(G1293) );
nand2 gate485( .a(G1232), .b(G1233), .O(G1294) );
nand2 gate486( .a(G1234), .b(G1235), .O(G1295) );

  xor2  gate1849(.a(G1237), .b(G1236), .O(gate487inter0));
  nand2 gate1850(.a(gate487inter0), .b(s_186), .O(gate487inter1));
  and2  gate1851(.a(G1237), .b(G1236), .O(gate487inter2));
  inv1  gate1852(.a(s_186), .O(gate487inter3));
  inv1  gate1853(.a(s_187), .O(gate487inter4));
  nand2 gate1854(.a(gate487inter4), .b(gate487inter3), .O(gate487inter5));
  nor2  gate1855(.a(gate487inter5), .b(gate487inter2), .O(gate487inter6));
  inv1  gate1856(.a(G1236), .O(gate487inter7));
  inv1  gate1857(.a(G1237), .O(gate487inter8));
  nand2 gate1858(.a(gate487inter8), .b(gate487inter7), .O(gate487inter9));
  nand2 gate1859(.a(s_187), .b(gate487inter3), .O(gate487inter10));
  nor2  gate1860(.a(gate487inter10), .b(gate487inter9), .O(gate487inter11));
  nor2  gate1861(.a(gate487inter11), .b(gate487inter6), .O(gate487inter12));
  nand2 gate1862(.a(gate487inter12), .b(gate487inter1), .O(G1296));

  xor2  gate1093(.a(G1239), .b(G1238), .O(gate488inter0));
  nand2 gate1094(.a(gate488inter0), .b(s_78), .O(gate488inter1));
  and2  gate1095(.a(G1239), .b(G1238), .O(gate488inter2));
  inv1  gate1096(.a(s_78), .O(gate488inter3));
  inv1  gate1097(.a(s_79), .O(gate488inter4));
  nand2 gate1098(.a(gate488inter4), .b(gate488inter3), .O(gate488inter5));
  nor2  gate1099(.a(gate488inter5), .b(gate488inter2), .O(gate488inter6));
  inv1  gate1100(.a(G1238), .O(gate488inter7));
  inv1  gate1101(.a(G1239), .O(gate488inter8));
  nand2 gate1102(.a(gate488inter8), .b(gate488inter7), .O(gate488inter9));
  nand2 gate1103(.a(s_79), .b(gate488inter3), .O(gate488inter10));
  nor2  gate1104(.a(gate488inter10), .b(gate488inter9), .O(gate488inter11));
  nor2  gate1105(.a(gate488inter11), .b(gate488inter6), .O(gate488inter12));
  nand2 gate1106(.a(gate488inter12), .b(gate488inter1), .O(G1297));

  xor2  gate631(.a(G1241), .b(G1240), .O(gate489inter0));
  nand2 gate632(.a(gate489inter0), .b(s_12), .O(gate489inter1));
  and2  gate633(.a(G1241), .b(G1240), .O(gate489inter2));
  inv1  gate634(.a(s_12), .O(gate489inter3));
  inv1  gate635(.a(s_13), .O(gate489inter4));
  nand2 gate636(.a(gate489inter4), .b(gate489inter3), .O(gate489inter5));
  nor2  gate637(.a(gate489inter5), .b(gate489inter2), .O(gate489inter6));
  inv1  gate638(.a(G1240), .O(gate489inter7));
  inv1  gate639(.a(G1241), .O(gate489inter8));
  nand2 gate640(.a(gate489inter8), .b(gate489inter7), .O(gate489inter9));
  nand2 gate641(.a(s_13), .b(gate489inter3), .O(gate489inter10));
  nor2  gate642(.a(gate489inter10), .b(gate489inter9), .O(gate489inter11));
  nor2  gate643(.a(gate489inter11), .b(gate489inter6), .O(gate489inter12));
  nand2 gate644(.a(gate489inter12), .b(gate489inter1), .O(G1298));
nand2 gate490( .a(G1242), .b(G1243), .O(G1299) );
nand2 gate491( .a(G1244), .b(G1245), .O(G1300) );

  xor2  gate1527(.a(G1247), .b(G1246), .O(gate492inter0));
  nand2 gate1528(.a(gate492inter0), .b(s_140), .O(gate492inter1));
  and2  gate1529(.a(G1247), .b(G1246), .O(gate492inter2));
  inv1  gate1530(.a(s_140), .O(gate492inter3));
  inv1  gate1531(.a(s_141), .O(gate492inter4));
  nand2 gate1532(.a(gate492inter4), .b(gate492inter3), .O(gate492inter5));
  nor2  gate1533(.a(gate492inter5), .b(gate492inter2), .O(gate492inter6));
  inv1  gate1534(.a(G1246), .O(gate492inter7));
  inv1  gate1535(.a(G1247), .O(gate492inter8));
  nand2 gate1536(.a(gate492inter8), .b(gate492inter7), .O(gate492inter9));
  nand2 gate1537(.a(s_141), .b(gate492inter3), .O(gate492inter10));
  nor2  gate1538(.a(gate492inter10), .b(gate492inter9), .O(gate492inter11));
  nor2  gate1539(.a(gate492inter11), .b(gate492inter6), .O(gate492inter12));
  nand2 gate1540(.a(gate492inter12), .b(gate492inter1), .O(G1301));
nand2 gate493( .a(G1248), .b(G1249), .O(G1302) );

  xor2  gate939(.a(G1251), .b(G1250), .O(gate494inter0));
  nand2 gate940(.a(gate494inter0), .b(s_56), .O(gate494inter1));
  and2  gate941(.a(G1251), .b(G1250), .O(gate494inter2));
  inv1  gate942(.a(s_56), .O(gate494inter3));
  inv1  gate943(.a(s_57), .O(gate494inter4));
  nand2 gate944(.a(gate494inter4), .b(gate494inter3), .O(gate494inter5));
  nor2  gate945(.a(gate494inter5), .b(gate494inter2), .O(gate494inter6));
  inv1  gate946(.a(G1250), .O(gate494inter7));
  inv1  gate947(.a(G1251), .O(gate494inter8));
  nand2 gate948(.a(gate494inter8), .b(gate494inter7), .O(gate494inter9));
  nand2 gate949(.a(s_57), .b(gate494inter3), .O(gate494inter10));
  nor2  gate950(.a(gate494inter10), .b(gate494inter9), .O(gate494inter11));
  nor2  gate951(.a(gate494inter11), .b(gate494inter6), .O(gate494inter12));
  nand2 gate952(.a(gate494inter12), .b(gate494inter1), .O(G1303));

  xor2  gate617(.a(G1253), .b(G1252), .O(gate495inter0));
  nand2 gate618(.a(gate495inter0), .b(s_10), .O(gate495inter1));
  and2  gate619(.a(G1253), .b(G1252), .O(gate495inter2));
  inv1  gate620(.a(s_10), .O(gate495inter3));
  inv1  gate621(.a(s_11), .O(gate495inter4));
  nand2 gate622(.a(gate495inter4), .b(gate495inter3), .O(gate495inter5));
  nor2  gate623(.a(gate495inter5), .b(gate495inter2), .O(gate495inter6));
  inv1  gate624(.a(G1252), .O(gate495inter7));
  inv1  gate625(.a(G1253), .O(gate495inter8));
  nand2 gate626(.a(gate495inter8), .b(gate495inter7), .O(gate495inter9));
  nand2 gate627(.a(s_11), .b(gate495inter3), .O(gate495inter10));
  nor2  gate628(.a(gate495inter10), .b(gate495inter9), .O(gate495inter11));
  nor2  gate629(.a(gate495inter11), .b(gate495inter6), .O(gate495inter12));
  nand2 gate630(.a(gate495inter12), .b(gate495inter1), .O(G1304));
nand2 gate496( .a(G1254), .b(G1255), .O(G1305) );
nand2 gate497( .a(G1256), .b(G1257), .O(G1306) );
nand2 gate498( .a(G1258), .b(G1259), .O(G1307) );

  xor2  gate2017(.a(G1261), .b(G1260), .O(gate499inter0));
  nand2 gate2018(.a(gate499inter0), .b(s_210), .O(gate499inter1));
  and2  gate2019(.a(G1261), .b(G1260), .O(gate499inter2));
  inv1  gate2020(.a(s_210), .O(gate499inter3));
  inv1  gate2021(.a(s_211), .O(gate499inter4));
  nand2 gate2022(.a(gate499inter4), .b(gate499inter3), .O(gate499inter5));
  nor2  gate2023(.a(gate499inter5), .b(gate499inter2), .O(gate499inter6));
  inv1  gate2024(.a(G1260), .O(gate499inter7));
  inv1  gate2025(.a(G1261), .O(gate499inter8));
  nand2 gate2026(.a(gate499inter8), .b(gate499inter7), .O(gate499inter9));
  nand2 gate2027(.a(s_211), .b(gate499inter3), .O(gate499inter10));
  nor2  gate2028(.a(gate499inter10), .b(gate499inter9), .O(gate499inter11));
  nor2  gate2029(.a(gate499inter11), .b(gate499inter6), .O(gate499inter12));
  nand2 gate2030(.a(gate499inter12), .b(gate499inter1), .O(G1308));

  xor2  gate1695(.a(G1263), .b(G1262), .O(gate500inter0));
  nand2 gate1696(.a(gate500inter0), .b(s_164), .O(gate500inter1));
  and2  gate1697(.a(G1263), .b(G1262), .O(gate500inter2));
  inv1  gate1698(.a(s_164), .O(gate500inter3));
  inv1  gate1699(.a(s_165), .O(gate500inter4));
  nand2 gate1700(.a(gate500inter4), .b(gate500inter3), .O(gate500inter5));
  nor2  gate1701(.a(gate500inter5), .b(gate500inter2), .O(gate500inter6));
  inv1  gate1702(.a(G1262), .O(gate500inter7));
  inv1  gate1703(.a(G1263), .O(gate500inter8));
  nand2 gate1704(.a(gate500inter8), .b(gate500inter7), .O(gate500inter9));
  nand2 gate1705(.a(s_165), .b(gate500inter3), .O(gate500inter10));
  nor2  gate1706(.a(gate500inter10), .b(gate500inter9), .O(gate500inter11));
  nor2  gate1707(.a(gate500inter11), .b(gate500inter6), .O(gate500inter12));
  nand2 gate1708(.a(gate500inter12), .b(gate500inter1), .O(G1309));
nand2 gate501( .a(G1264), .b(G1265), .O(G1310) );
nand2 gate502( .a(G1266), .b(G1267), .O(G1311) );
nand2 gate503( .a(G1268), .b(G1269), .O(G1312) );

  xor2  gate827(.a(G1271), .b(G1270), .O(gate504inter0));
  nand2 gate828(.a(gate504inter0), .b(s_40), .O(gate504inter1));
  and2  gate829(.a(G1271), .b(G1270), .O(gate504inter2));
  inv1  gate830(.a(s_40), .O(gate504inter3));
  inv1  gate831(.a(s_41), .O(gate504inter4));
  nand2 gate832(.a(gate504inter4), .b(gate504inter3), .O(gate504inter5));
  nor2  gate833(.a(gate504inter5), .b(gate504inter2), .O(gate504inter6));
  inv1  gate834(.a(G1270), .O(gate504inter7));
  inv1  gate835(.a(G1271), .O(gate504inter8));
  nand2 gate836(.a(gate504inter8), .b(gate504inter7), .O(gate504inter9));
  nand2 gate837(.a(s_41), .b(gate504inter3), .O(gate504inter10));
  nor2  gate838(.a(gate504inter10), .b(gate504inter9), .O(gate504inter11));
  nor2  gate839(.a(gate504inter11), .b(gate504inter6), .O(gate504inter12));
  nand2 gate840(.a(gate504inter12), .b(gate504inter1), .O(G1313));
nand2 gate505( .a(G1272), .b(G1273), .O(G1314) );

  xor2  gate2073(.a(G1275), .b(G1274), .O(gate506inter0));
  nand2 gate2074(.a(gate506inter0), .b(s_218), .O(gate506inter1));
  and2  gate2075(.a(G1275), .b(G1274), .O(gate506inter2));
  inv1  gate2076(.a(s_218), .O(gate506inter3));
  inv1  gate2077(.a(s_219), .O(gate506inter4));
  nand2 gate2078(.a(gate506inter4), .b(gate506inter3), .O(gate506inter5));
  nor2  gate2079(.a(gate506inter5), .b(gate506inter2), .O(gate506inter6));
  inv1  gate2080(.a(G1274), .O(gate506inter7));
  inv1  gate2081(.a(G1275), .O(gate506inter8));
  nand2 gate2082(.a(gate506inter8), .b(gate506inter7), .O(gate506inter9));
  nand2 gate2083(.a(s_219), .b(gate506inter3), .O(gate506inter10));
  nor2  gate2084(.a(gate506inter10), .b(gate506inter9), .O(gate506inter11));
  nor2  gate2085(.a(gate506inter11), .b(gate506inter6), .O(gate506inter12));
  nand2 gate2086(.a(gate506inter12), .b(gate506inter1), .O(G1315));
nand2 gate507( .a(G1276), .b(G1277), .O(G1316) );
nand2 gate508( .a(G1278), .b(G1279), .O(G1317) );
nand2 gate509( .a(G1280), .b(G1281), .O(G1318) );
nand2 gate510( .a(G1282), .b(G1283), .O(G1319) );
nand2 gate511( .a(G1284), .b(G1285), .O(G1320) );

  xor2  gate771(.a(G1287), .b(G1286), .O(gate512inter0));
  nand2 gate772(.a(gate512inter0), .b(s_32), .O(gate512inter1));
  and2  gate773(.a(G1287), .b(G1286), .O(gate512inter2));
  inv1  gate774(.a(s_32), .O(gate512inter3));
  inv1  gate775(.a(s_33), .O(gate512inter4));
  nand2 gate776(.a(gate512inter4), .b(gate512inter3), .O(gate512inter5));
  nor2  gate777(.a(gate512inter5), .b(gate512inter2), .O(gate512inter6));
  inv1  gate778(.a(G1286), .O(gate512inter7));
  inv1  gate779(.a(G1287), .O(gate512inter8));
  nand2 gate780(.a(gate512inter8), .b(gate512inter7), .O(gate512inter9));
  nand2 gate781(.a(s_33), .b(gate512inter3), .O(gate512inter10));
  nor2  gate782(.a(gate512inter10), .b(gate512inter9), .O(gate512inter11));
  nor2  gate783(.a(gate512inter11), .b(gate512inter6), .O(gate512inter12));
  nand2 gate784(.a(gate512inter12), .b(gate512inter1), .O(G1321));
nand2 gate513( .a(G1288), .b(G1289), .O(G1322) );

  xor2  gate1065(.a(G1291), .b(G1290), .O(gate514inter0));
  nand2 gate1066(.a(gate514inter0), .b(s_74), .O(gate514inter1));
  and2  gate1067(.a(G1291), .b(G1290), .O(gate514inter2));
  inv1  gate1068(.a(s_74), .O(gate514inter3));
  inv1  gate1069(.a(s_75), .O(gate514inter4));
  nand2 gate1070(.a(gate514inter4), .b(gate514inter3), .O(gate514inter5));
  nor2  gate1071(.a(gate514inter5), .b(gate514inter2), .O(gate514inter6));
  inv1  gate1072(.a(G1290), .O(gate514inter7));
  inv1  gate1073(.a(G1291), .O(gate514inter8));
  nand2 gate1074(.a(gate514inter8), .b(gate514inter7), .O(gate514inter9));
  nand2 gate1075(.a(s_75), .b(gate514inter3), .O(gate514inter10));
  nor2  gate1076(.a(gate514inter10), .b(gate514inter9), .O(gate514inter11));
  nor2  gate1077(.a(gate514inter11), .b(gate514inter6), .O(gate514inter12));
  nand2 gate1078(.a(gate514inter12), .b(gate514inter1), .O(G1323));
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule