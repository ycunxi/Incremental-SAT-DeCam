module c432 (N1,N4,N8,N11,N14,N17,N21,N24,N27,N30,
             N34,N37,N40,N43,N47,N50,N53,N56,N60,N63,
             N66,N69,N73,N76,N79,N82,N86,N89,N92,N95,
             N99,N102,N105,N108,N112,N115,N223,N329,N370,N421,
             N430,N431,N432);

input N1,N4,N8,N11,N14,N17,N21,N24,N27,N30,
      N34,N37,N40,N43,N47,N50,N53,N56,N60,N63,
      N66,N69,N73,N76,N79,N82,N86,N89,N92,N95,
      N99,N102,N105,N108,N112,N115;//RE__PI;

input s_0,s_1;//RE__ALLOW(00,01,10,11);
input s_2,s_3;//RE__ALLOW(00,01,10,11);
input s_4,s_5;//RE__ALLOW(00,01,10,11);
input s_6,s_7;//RE__ALLOW(00,01,10,11);
input s_8,s_9;//RE__ALLOW(00,01,10,11);
input s_10,s_11;//RE__ALLOW(00,01,10,11);
input s_12,s_13;//RE__ALLOW(00,01,10,11);
input s_14,s_15;//RE__ALLOW(00,01,10,11);
input s_16,s_17;//RE__ALLOW(00,01,10,11);
input s_18,s_19;//RE__ALLOW(00,01,10,11);
input s_20,s_21;//RE__ALLOW(00,01,10,11);
input s_22,s_23;//RE__ALLOW(00,01,10,11);
input s_24,s_25;//RE__ALLOW(00,01,10,11);
input s_26,s_27;//RE__ALLOW(00,01,10,11);
input s_28,s_29;//RE__ALLOW(00,01,10,11);
input s_30,s_31;//RE__ALLOW(00,01,10,11);
input s_32,s_33;//RE__ALLOW(00,01,10,11);
input s_34,s_35;//RE__ALLOW(00,01,10,11);
input s_36,s_37;//RE__ALLOW(00,01,10,11);
input s_38,s_39;//RE__ALLOW(00,01,10,11);
input s_40,s_41;//RE__ALLOW(00,01,10,11);
input s_42,s_43;//RE__ALLOW(00,01,10,11);
input s_44,s_45;//RE__ALLOW(00,01,10,11);
input s_46,s_47;//RE__ALLOW(00,01,10,11);
input s_48,s_49;//RE__ALLOW(00,01,10,11);
input s_50,s_51;//RE__ALLOW(00,01,10,11);
input s_52,s_53;//RE__ALLOW(00,01,10,11);
input s_54,s_55;//RE__ALLOW(00,01,10,11);
input s_56,s_57;//RE__ALLOW(00,01,10,11);
input s_58,s_59;//RE__ALLOW(00,01,10,11);
input s_60,s_61;//RE__ALLOW(00,01,10,11);
input s_62,s_63;//RE__ALLOW(00,01,10,11);
input s_64,s_65;//RE__ALLOW(00,01,10,11);
input s_66,s_67;//RE__ALLOW(00,01,10,11);
input s_68,s_69;//RE__ALLOW(00,01,10,11);
input s_70,s_71;//RE__ALLOW(00,01,10,11);
output N223,N329,N370,N421,N430,N431,N432;

wire N118,N119,N122,N123,N126,N127,N130,N131,N134,N135,
     N138,N139,N142,N143,N146,N147,N150,N151,N154,N157,
     N158,N159,N162,N165,N168,N171,N174,N177,N180,N183,
     N184,N185,N186,N187,N188,N189,N190,N191,N192,N193,
     N194,N195,N196,N197,N198,N199,N203,N213,N224,N227,
     N230,N233,N236,N239,N242,N243,N246,N247,N250,N251,
     N254,N255,N256,N257,N258,N259,N260,N263,N264,N267,
     N270,N273,N276,N279,N282,N285,N288,N289,N290,N291,
     N292,N293,N294,N295,N296,N300,N301,N302,N303,N304,
     N305,N306,N307,N308,N309,N319,N330,N331,N332,N333,
     N334,N335,N336,N337,N338,N339,N340,N341,N342,N343,
     N344,N345,N346,N347,N348,N349,N350,N351,N352,N353,
     N354,N355,N356,N357,N360,N371,N372,N373,N374,N375,
     N376,N377,N378,N379,N380,N381,N386,N393,N399,N404,
     N407,N411,N414,N415,N416,N417,N418,N419,N420,N422,
     N425,N428,N429, gate71inter0, gate71inter1, gate71inter2, gate71inter3, gate71inter4, gate71inter5, gate71inter6, gate71inter7, gate71inter8, gate71inter9, gate71inter10, gate71inter11, gate71inter12, gate83inter0, gate83inter1, gate83inter2, gate83inter3, gate83inter4, gate83inter5, gate83inter6, gate83inter7, gate83inter8, gate83inter9, gate83inter10, gate83inter11, gate83inter12, gate132inter0, gate132inter1, gate132inter2, gate132inter3, gate132inter4, gate132inter5, gate132inter6, gate132inter7, gate132inter8, gate132inter9, gate132inter10, gate132inter11, gate132inter12, gate72inter0, gate72inter1, gate72inter2, gate72inter3, gate72inter4, gate72inter5, gate72inter6, gate72inter7, gate72inter8, gate72inter9, gate72inter10, gate72inter11, gate72inter12, gate117inter0, gate117inter1, gate117inter2, gate117inter3, gate117inter4, gate117inter5, gate117inter6, gate117inter7, gate117inter8, gate117inter9, gate117inter10, gate117inter11, gate117inter12, gate42inter0, gate42inter1, gate42inter2, gate42inter3, gate42inter4, gate42inter5, gate42inter6, gate42inter7, gate42inter8, gate42inter9, gate42inter10, gate42inter11, gate42inter12, gate130inter0, gate130inter1, gate130inter2, gate130inter3, gate130inter4, gate130inter5, gate130inter6, gate130inter7, gate130inter8, gate130inter9, gate130inter10, gate130inter11, gate130inter12, gate70inter0, gate70inter1, gate70inter2, gate70inter3, gate70inter4, gate70inter5, gate70inter6, gate70inter7, gate70inter8, gate70inter9, gate70inter10, gate70inter11, gate70inter12, gate60inter0, gate60inter1, gate60inter2, gate60inter3, gate60inter4, gate60inter5, gate60inter6, gate60inter7, gate60inter8, gate60inter9, gate60inter10, gate60inter11, gate60inter12, gate24inter0, gate24inter1, gate24inter2, gate24inter3, gate24inter4, gate24inter5, gate24inter6, gate24inter7, gate24inter8, gate24inter9, gate24inter10, gate24inter11, gate24inter12, gate52inter0, gate52inter1, gate52inter2, gate52inter3, gate52inter4, gate52inter5, gate52inter6, gate52inter7, gate52inter8, gate52inter9, gate52inter10, gate52inter11, gate52inter12, gate107inter0, gate107inter1, gate107inter2, gate107inter3, gate107inter4, gate107inter5, gate107inter6, gate107inter7, gate107inter8, gate107inter9, gate107inter10, gate107inter11, gate107inter12, gate115inter0, gate115inter1, gate115inter2, gate115inter3, gate115inter4, gate115inter5, gate115inter6, gate115inter7, gate115inter8, gate115inter9, gate115inter10, gate115inter11, gate115inter12, gate77inter0, gate77inter1, gate77inter2, gate77inter3, gate77inter4, gate77inter5, gate77inter6, gate77inter7, gate77inter8, gate77inter9, gate77inter10, gate77inter11, gate77inter12, gate22inter0, gate22inter1, gate22inter2, gate22inter3, gate22inter4, gate22inter5, gate22inter6, gate22inter7, gate22inter8, gate22inter9, gate22inter10, gate22inter11, gate22inter12, gate121inter0, gate121inter1, gate121inter2, gate121inter3, gate121inter4, gate121inter5, gate121inter6, gate121inter7, gate121inter8, gate121inter9, gate121inter10, gate121inter11, gate121inter12, gate69inter0, gate69inter1, gate69inter2, gate69inter3, gate69inter4, gate69inter5, gate69inter6, gate69inter7, gate69inter8, gate69inter9, gate69inter10, gate69inter11, gate69inter12, gate29inter0, gate29inter1, gate29inter2, gate29inter3, gate29inter4, gate29inter5, gate29inter6, gate29inter7, gate29inter8, gate29inter9, gate29inter10, gate29inter11, gate29inter12, gate30inter0, gate30inter1, gate30inter2, gate30inter3, gate30inter4, gate30inter5, gate30inter6, gate30inter7, gate30inter8, gate30inter9, gate30inter10, gate30inter11, gate30inter12, gate57inter0, gate57inter1, gate57inter2, gate57inter3, gate57inter4, gate57inter5, gate57inter6, gate57inter7, gate57inter8, gate57inter9, gate57inter10, gate57inter11, gate57inter12, gate112inter0, gate112inter1, gate112inter2, gate112inter3, gate112inter4, gate112inter5, gate112inter6, gate112inter7, gate112inter8, gate112inter9, gate112inter10, gate112inter11, gate112inter12, gate41inter0, gate41inter1, gate41inter2, gate41inter3, gate41inter4, gate41inter5, gate41inter6, gate41inter7, gate41inter8, gate41inter9, gate41inter10, gate41inter11, gate41inter12, gate65inter0, gate65inter1, gate65inter2, gate65inter3, gate65inter4, gate65inter5, gate65inter6, gate65inter7, gate65inter8, gate65inter9, gate65inter10, gate65inter11, gate65inter12, gate74inter0, gate74inter1, gate74inter2, gate74inter3, gate74inter4, gate74inter5, gate74inter6, gate74inter7, gate74inter8, gate74inter9, gate74inter10, gate74inter11, gate74inter12, gate35inter0, gate35inter1, gate35inter2, gate35inter3, gate35inter4, gate35inter5, gate35inter6, gate35inter7, gate35inter8, gate35inter9, gate35inter10, gate35inter11, gate35inter12, gate100inter0, gate100inter1, gate100inter2, gate100inter3, gate100inter4, gate100inter5, gate100inter6, gate100inter7, gate100inter8, gate100inter9, gate100inter10, gate100inter11, gate100inter12, gate63inter0, gate63inter1, gate63inter2, gate63inter3, gate63inter4, gate63inter5, gate63inter6, gate63inter7, gate63inter8, gate63inter9, gate63inter10, gate63inter11, gate63inter12, gate79inter0, gate79inter1, gate79inter2, gate79inter3, gate79inter4, gate79inter5, gate79inter6, gate79inter7, gate79inter8, gate79inter9, gate79inter10, gate79inter11, gate79inter12, gate103inter0, gate103inter1, gate103inter2, gate103inter3, gate103inter4, gate103inter5, gate103inter6, gate103inter7, gate103inter8, gate103inter9, gate103inter10, gate103inter11, gate103inter12, gate122inter0, gate122inter1, gate122inter2, gate122inter3, gate122inter4, gate122inter5, gate122inter6, gate122inter7, gate122inter8, gate122inter9, gate122inter10, gate122inter11, gate122inter12, gate50inter0, gate50inter1, gate50inter2, gate50inter3, gate50inter4, gate50inter5, gate50inter6, gate50inter7, gate50inter8, gate50inter9, gate50inter10, gate50inter11, gate50inter12, gate25inter0, gate25inter1, gate25inter2, gate25inter3, gate25inter4, gate25inter5, gate25inter6, gate25inter7, gate25inter8, gate25inter9, gate25inter10, gate25inter11, gate25inter12, gate62inter0, gate62inter1, gate62inter2, gate62inter3, gate62inter4, gate62inter5, gate62inter6, gate62inter7, gate62inter8, gate62inter9, gate62inter10, gate62inter11, gate62inter12, gate64inter0, gate64inter1, gate64inter2, gate64inter3, gate64inter4, gate64inter5, gate64inter6, gate64inter7, gate64inter8, gate64inter9, gate64inter10, gate64inter11, gate64inter12, gate23inter0, gate23inter1, gate23inter2, gate23inter3, gate23inter4, gate23inter5, gate23inter6, gate23inter7, gate23inter8, gate23inter9, gate23inter10, gate23inter11, gate23inter12, gate106inter0, gate106inter1, gate106inter2, gate106inter3, gate106inter4, gate106inter5, gate106inter6, gate106inter7, gate106inter8, gate106inter9, gate106inter10, gate106inter11, gate106inter12;



inv1 gate1( .a(N1), .O(N118) );
inv1 gate2( .a(N4), .O(N119) );
inv1 gate3( .a(N11), .O(N122) );
inv1 gate4( .a(N17), .O(N123) );
inv1 gate5( .a(N24), .O(N126) );
inv1 gate6( .a(N30), .O(N127) );
inv1 gate7( .a(N37), .O(N130) );
inv1 gate8( .a(N43), .O(N131) );
inv1 gate9( .a(N50), .O(N134) );
inv1 gate10( .a(N56), .O(N135) );
inv1 gate11( .a(N63), .O(N138) );
inv1 gate12( .a(N69), .O(N139) );
inv1 gate13( .a(N76), .O(N142) );
inv1 gate14( .a(N82), .O(N143) );
inv1 gate15( .a(N89), .O(N146) );
inv1 gate16( .a(N95), .O(N147) );
inv1 gate17( .a(N102), .O(N150) );
inv1 gate18( .a(N108), .O(N151) );
nand2 gate19( .a(N118), .b(N4), .O(N154) );
nor2 gate20( .a(N8), .b(N119), .O(N157) );
nor2 gate21( .a(N14), .b(N119), .O(N158) );

  xor2  gate357(.a(N17), .b(N122), .O(gate22inter0));
  nand2 gate358(.a(gate22inter0), .b(s_28), .O(gate22inter1));
  and2  gate359(.a(N17), .b(N122), .O(gate22inter2));
  inv1  gate360(.a(s_28), .O(gate22inter3));
  inv1  gate361(.a(s_29), .O(gate22inter4));
  nand2 gate362(.a(gate22inter4), .b(gate22inter3), .O(gate22inter5));
  nor2  gate363(.a(gate22inter5), .b(gate22inter2), .O(gate22inter6));
  inv1  gate364(.a(N122), .O(gate22inter7));
  inv1  gate365(.a(N17), .O(gate22inter8));
  nand2 gate366(.a(gate22inter8), .b(gate22inter7), .O(gate22inter9));
  nand2 gate367(.a(s_29), .b(gate22inter3), .O(gate22inter10));
  nor2  gate368(.a(gate22inter10), .b(gate22inter9), .O(gate22inter11));
  nor2  gate369(.a(gate22inter11), .b(gate22inter6), .O(gate22inter12));
  nand2 gate370(.a(gate22inter12), .b(gate22inter1), .O(N159));

  xor2  gate637(.a(N30), .b(N126), .O(gate23inter0));
  nand2 gate638(.a(gate23inter0), .b(s_68), .O(gate23inter1));
  and2  gate639(.a(N30), .b(N126), .O(gate23inter2));
  inv1  gate640(.a(s_68), .O(gate23inter3));
  inv1  gate641(.a(s_69), .O(gate23inter4));
  nand2 gate642(.a(gate23inter4), .b(gate23inter3), .O(gate23inter5));
  nor2  gate643(.a(gate23inter5), .b(gate23inter2), .O(gate23inter6));
  inv1  gate644(.a(N126), .O(gate23inter7));
  inv1  gate645(.a(N30), .O(gate23inter8));
  nand2 gate646(.a(gate23inter8), .b(gate23inter7), .O(gate23inter9));
  nand2 gate647(.a(s_69), .b(gate23inter3), .O(gate23inter10));
  nor2  gate648(.a(gate23inter10), .b(gate23inter9), .O(gate23inter11));
  nor2  gate649(.a(gate23inter11), .b(gate23inter6), .O(gate23inter12));
  nand2 gate650(.a(gate23inter12), .b(gate23inter1), .O(N162));

  xor2  gate287(.a(N43), .b(N130), .O(gate24inter0));
  nand2 gate288(.a(gate24inter0), .b(s_18), .O(gate24inter1));
  and2  gate289(.a(N43), .b(N130), .O(gate24inter2));
  inv1  gate290(.a(s_18), .O(gate24inter3));
  inv1  gate291(.a(s_19), .O(gate24inter4));
  nand2 gate292(.a(gate24inter4), .b(gate24inter3), .O(gate24inter5));
  nor2  gate293(.a(gate24inter5), .b(gate24inter2), .O(gate24inter6));
  inv1  gate294(.a(N130), .O(gate24inter7));
  inv1  gate295(.a(N43), .O(gate24inter8));
  nand2 gate296(.a(gate24inter8), .b(gate24inter7), .O(gate24inter9));
  nand2 gate297(.a(s_19), .b(gate24inter3), .O(gate24inter10));
  nor2  gate298(.a(gate24inter10), .b(gate24inter9), .O(gate24inter11));
  nor2  gate299(.a(gate24inter11), .b(gate24inter6), .O(gate24inter12));
  nand2 gate300(.a(gate24inter12), .b(gate24inter1), .O(N165));

  xor2  gate595(.a(N56), .b(N134), .O(gate25inter0));
  nand2 gate596(.a(gate25inter0), .b(s_62), .O(gate25inter1));
  and2  gate597(.a(N56), .b(N134), .O(gate25inter2));
  inv1  gate598(.a(s_62), .O(gate25inter3));
  inv1  gate599(.a(s_63), .O(gate25inter4));
  nand2 gate600(.a(gate25inter4), .b(gate25inter3), .O(gate25inter5));
  nor2  gate601(.a(gate25inter5), .b(gate25inter2), .O(gate25inter6));
  inv1  gate602(.a(N134), .O(gate25inter7));
  inv1  gate603(.a(N56), .O(gate25inter8));
  nand2 gate604(.a(gate25inter8), .b(gate25inter7), .O(gate25inter9));
  nand2 gate605(.a(s_63), .b(gate25inter3), .O(gate25inter10));
  nor2  gate606(.a(gate25inter10), .b(gate25inter9), .O(gate25inter11));
  nor2  gate607(.a(gate25inter11), .b(gate25inter6), .O(gate25inter12));
  nand2 gate608(.a(gate25inter12), .b(gate25inter1), .O(N168));
nand2 gate26( .a(N138), .b(N69), .O(N171) );
nand2 gate27( .a(N142), .b(N82), .O(N174) );
nand2 gate28( .a(N146), .b(N95), .O(N177) );

  xor2  gate399(.a(N108), .b(N150), .O(gate29inter0));
  nand2 gate400(.a(gate29inter0), .b(s_34), .O(gate29inter1));
  and2  gate401(.a(N108), .b(N150), .O(gate29inter2));
  inv1  gate402(.a(s_34), .O(gate29inter3));
  inv1  gate403(.a(s_35), .O(gate29inter4));
  nand2 gate404(.a(gate29inter4), .b(gate29inter3), .O(gate29inter5));
  nor2  gate405(.a(gate29inter5), .b(gate29inter2), .O(gate29inter6));
  inv1  gate406(.a(N150), .O(gate29inter7));
  inv1  gate407(.a(N108), .O(gate29inter8));
  nand2 gate408(.a(gate29inter8), .b(gate29inter7), .O(gate29inter9));
  nand2 gate409(.a(s_35), .b(gate29inter3), .O(gate29inter10));
  nor2  gate410(.a(gate29inter10), .b(gate29inter9), .O(gate29inter11));
  nor2  gate411(.a(gate29inter11), .b(gate29inter6), .O(gate29inter12));
  nand2 gate412(.a(gate29inter12), .b(gate29inter1), .O(N180));

  xor2  gate413(.a(N123), .b(N21), .O(gate30inter0));
  nand2 gate414(.a(gate30inter0), .b(s_36), .O(gate30inter1));
  and2  gate415(.a(N123), .b(N21), .O(gate30inter2));
  inv1  gate416(.a(s_36), .O(gate30inter3));
  inv1  gate417(.a(s_37), .O(gate30inter4));
  nand2 gate418(.a(gate30inter4), .b(gate30inter3), .O(gate30inter5));
  nor2  gate419(.a(gate30inter5), .b(gate30inter2), .O(gate30inter6));
  inv1  gate420(.a(N21), .O(gate30inter7));
  inv1  gate421(.a(N123), .O(gate30inter8));
  nand2 gate422(.a(gate30inter8), .b(gate30inter7), .O(gate30inter9));
  nand2 gate423(.a(s_37), .b(gate30inter3), .O(gate30inter10));
  nor2  gate424(.a(gate30inter10), .b(gate30inter9), .O(gate30inter11));
  nor2  gate425(.a(gate30inter11), .b(gate30inter6), .O(gate30inter12));
  nand2 gate426(.a(gate30inter12), .b(gate30inter1), .O(N183));
nor2 gate31( .a(N27), .b(N123), .O(N184) );
nor2 gate32( .a(N34), .b(N127), .O(N185) );
nor2 gate33( .a(N40), .b(N127), .O(N186) );
nor2 gate34( .a(N47), .b(N131), .O(N187) );

  xor2  gate497(.a(N131), .b(N53), .O(gate35inter0));
  nand2 gate498(.a(gate35inter0), .b(s_48), .O(gate35inter1));
  and2  gate499(.a(N131), .b(N53), .O(gate35inter2));
  inv1  gate500(.a(s_48), .O(gate35inter3));
  inv1  gate501(.a(s_49), .O(gate35inter4));
  nand2 gate502(.a(gate35inter4), .b(gate35inter3), .O(gate35inter5));
  nor2  gate503(.a(gate35inter5), .b(gate35inter2), .O(gate35inter6));
  inv1  gate504(.a(N53), .O(gate35inter7));
  inv1  gate505(.a(N131), .O(gate35inter8));
  nand2 gate506(.a(gate35inter8), .b(gate35inter7), .O(gate35inter9));
  nand2 gate507(.a(s_49), .b(gate35inter3), .O(gate35inter10));
  nor2  gate508(.a(gate35inter10), .b(gate35inter9), .O(gate35inter11));
  nor2  gate509(.a(gate35inter11), .b(gate35inter6), .O(gate35inter12));
  nand2 gate510(.a(gate35inter12), .b(gate35inter1), .O(N188));
nor2 gate36( .a(N60), .b(N135), .O(N189) );
nor2 gate37( .a(N66), .b(N135), .O(N190) );
nor2 gate38( .a(N73), .b(N139), .O(N191) );
nor2 gate39( .a(N79), .b(N139), .O(N192) );
nor2 gate40( .a(N86), .b(N143), .O(N193) );

  xor2  gate455(.a(N143), .b(N92), .O(gate41inter0));
  nand2 gate456(.a(gate41inter0), .b(s_42), .O(gate41inter1));
  and2  gate457(.a(N143), .b(N92), .O(gate41inter2));
  inv1  gate458(.a(s_42), .O(gate41inter3));
  inv1  gate459(.a(s_43), .O(gate41inter4));
  nand2 gate460(.a(gate41inter4), .b(gate41inter3), .O(gate41inter5));
  nor2  gate461(.a(gate41inter5), .b(gate41inter2), .O(gate41inter6));
  inv1  gate462(.a(N92), .O(gate41inter7));
  inv1  gate463(.a(N143), .O(gate41inter8));
  nand2 gate464(.a(gate41inter8), .b(gate41inter7), .O(gate41inter9));
  nand2 gate465(.a(s_43), .b(gate41inter3), .O(gate41inter10));
  nor2  gate466(.a(gate41inter10), .b(gate41inter9), .O(gate41inter11));
  nor2  gate467(.a(gate41inter11), .b(gate41inter6), .O(gate41inter12));
  nand2 gate468(.a(gate41inter12), .b(gate41inter1), .O(N194));

  xor2  gate231(.a(N147), .b(N99), .O(gate42inter0));
  nand2 gate232(.a(gate42inter0), .b(s_10), .O(gate42inter1));
  and2  gate233(.a(N147), .b(N99), .O(gate42inter2));
  inv1  gate234(.a(s_10), .O(gate42inter3));
  inv1  gate235(.a(s_11), .O(gate42inter4));
  nand2 gate236(.a(gate42inter4), .b(gate42inter3), .O(gate42inter5));
  nor2  gate237(.a(gate42inter5), .b(gate42inter2), .O(gate42inter6));
  inv1  gate238(.a(N99), .O(gate42inter7));
  inv1  gate239(.a(N147), .O(gate42inter8));
  nand2 gate240(.a(gate42inter8), .b(gate42inter7), .O(gate42inter9));
  nand2 gate241(.a(s_11), .b(gate42inter3), .O(gate42inter10));
  nor2  gate242(.a(gate42inter10), .b(gate42inter9), .O(gate42inter11));
  nor2  gate243(.a(gate42inter11), .b(gate42inter6), .O(gate42inter12));
  nand2 gate244(.a(gate42inter12), .b(gate42inter1), .O(N195));
nor2 gate43( .a(N105), .b(N147), .O(N196) );
nor2 gate44( .a(N112), .b(N151), .O(N197) );
nor2 gate45( .a(N115), .b(N151), .O(N198) );
and9 gate46( .a(N154), .b(N159), .c(N162), .d(N165), .e(N168), .f(N171), .g(N174), .h(N177), .i(N180), .O(N199) );
inv1 gate47( .a(N199), .O(N203) );
inv1 gate48( .a(N199), .O(N213) );
inv1 gate49( .a(N199), .O(N223) );

  xor2  gate581(.a(N154), .b(N203), .O(gate50inter0));
  nand2 gate582(.a(gate50inter0), .b(s_60), .O(gate50inter1));
  and2  gate583(.a(N154), .b(N203), .O(gate50inter2));
  inv1  gate584(.a(s_60), .O(gate50inter3));
  inv1  gate585(.a(s_61), .O(gate50inter4));
  nand2 gate586(.a(gate50inter4), .b(gate50inter3), .O(gate50inter5));
  nor2  gate587(.a(gate50inter5), .b(gate50inter2), .O(gate50inter6));
  inv1  gate588(.a(N203), .O(gate50inter7));
  inv1  gate589(.a(N154), .O(gate50inter8));
  nand2 gate590(.a(gate50inter8), .b(gate50inter7), .O(gate50inter9));
  nand2 gate591(.a(s_61), .b(gate50inter3), .O(gate50inter10));
  nor2  gate592(.a(gate50inter10), .b(gate50inter9), .O(gate50inter11));
  nor2  gate593(.a(gate50inter11), .b(gate50inter6), .O(gate50inter12));
  nand2 gate594(.a(gate50inter12), .b(gate50inter1), .O(N224));
xor2 gate51( .a(N203), .b(N159), .O(N227) );

  xor2  gate301(.a(N162), .b(N203), .O(gate52inter0));
  nand2 gate302(.a(gate52inter0), .b(s_20), .O(gate52inter1));
  and2  gate303(.a(N162), .b(N203), .O(gate52inter2));
  inv1  gate304(.a(s_20), .O(gate52inter3));
  inv1  gate305(.a(s_21), .O(gate52inter4));
  nand2 gate306(.a(gate52inter4), .b(gate52inter3), .O(gate52inter5));
  nor2  gate307(.a(gate52inter5), .b(gate52inter2), .O(gate52inter6));
  inv1  gate308(.a(N203), .O(gate52inter7));
  inv1  gate309(.a(N162), .O(gate52inter8));
  nand2 gate310(.a(gate52inter8), .b(gate52inter7), .O(gate52inter9));
  nand2 gate311(.a(s_21), .b(gate52inter3), .O(gate52inter10));
  nor2  gate312(.a(gate52inter10), .b(gate52inter9), .O(gate52inter11));
  nor2  gate313(.a(gate52inter11), .b(gate52inter6), .O(gate52inter12));
  nand2 gate314(.a(gate52inter12), .b(gate52inter1), .O(N230));
xor2 gate53( .a(N203), .b(N165), .O(N233) );
xor2 gate54( .a(N203), .b(N168), .O(N236) );
xor2 gate55( .a(N203), .b(N171), .O(N239) );
nand2 gate56( .a(N1), .b(N213), .O(N242) );

  xor2  gate427(.a(N174), .b(N203), .O(gate57inter0));
  nand2 gate428(.a(gate57inter0), .b(s_38), .O(gate57inter1));
  and2  gate429(.a(N174), .b(N203), .O(gate57inter2));
  inv1  gate430(.a(s_38), .O(gate57inter3));
  inv1  gate431(.a(s_39), .O(gate57inter4));
  nand2 gate432(.a(gate57inter4), .b(gate57inter3), .O(gate57inter5));
  nor2  gate433(.a(gate57inter5), .b(gate57inter2), .O(gate57inter6));
  inv1  gate434(.a(N203), .O(gate57inter7));
  inv1  gate435(.a(N174), .O(gate57inter8));
  nand2 gate436(.a(gate57inter8), .b(gate57inter7), .O(gate57inter9));
  nand2 gate437(.a(s_39), .b(gate57inter3), .O(gate57inter10));
  nor2  gate438(.a(gate57inter10), .b(gate57inter9), .O(gate57inter11));
  nor2  gate439(.a(gate57inter11), .b(gate57inter6), .O(gate57inter12));
  nand2 gate440(.a(gate57inter12), .b(gate57inter1), .O(N243));
nand2 gate58( .a(N213), .b(N11), .O(N246) );
xor2 gate59( .a(N203), .b(N177), .O(N247) );

  xor2  gate273(.a(N24), .b(N213), .O(gate60inter0));
  nand2 gate274(.a(gate60inter0), .b(s_16), .O(gate60inter1));
  and2  gate275(.a(N24), .b(N213), .O(gate60inter2));
  inv1  gate276(.a(s_16), .O(gate60inter3));
  inv1  gate277(.a(s_17), .O(gate60inter4));
  nand2 gate278(.a(gate60inter4), .b(gate60inter3), .O(gate60inter5));
  nor2  gate279(.a(gate60inter5), .b(gate60inter2), .O(gate60inter6));
  inv1  gate280(.a(N213), .O(gate60inter7));
  inv1  gate281(.a(N24), .O(gate60inter8));
  nand2 gate282(.a(gate60inter8), .b(gate60inter7), .O(gate60inter9));
  nand2 gate283(.a(s_17), .b(gate60inter3), .O(gate60inter10));
  nor2  gate284(.a(gate60inter10), .b(gate60inter9), .O(gate60inter11));
  nor2  gate285(.a(gate60inter11), .b(gate60inter6), .O(gate60inter12));
  nand2 gate286(.a(gate60inter12), .b(gate60inter1), .O(N250));
xor2 gate61( .a(N203), .b(N180), .O(N251) );

  xor2  gate609(.a(N37), .b(N213), .O(gate62inter0));
  nand2 gate610(.a(gate62inter0), .b(s_64), .O(gate62inter1));
  and2  gate611(.a(N37), .b(N213), .O(gate62inter2));
  inv1  gate612(.a(s_64), .O(gate62inter3));
  inv1  gate613(.a(s_65), .O(gate62inter4));
  nand2 gate614(.a(gate62inter4), .b(gate62inter3), .O(gate62inter5));
  nor2  gate615(.a(gate62inter5), .b(gate62inter2), .O(gate62inter6));
  inv1  gate616(.a(N213), .O(gate62inter7));
  inv1  gate617(.a(N37), .O(gate62inter8));
  nand2 gate618(.a(gate62inter8), .b(gate62inter7), .O(gate62inter9));
  nand2 gate619(.a(s_65), .b(gate62inter3), .O(gate62inter10));
  nor2  gate620(.a(gate62inter10), .b(gate62inter9), .O(gate62inter11));
  nor2  gate621(.a(gate62inter11), .b(gate62inter6), .O(gate62inter12));
  nand2 gate622(.a(gate62inter12), .b(gate62inter1), .O(N254));

  xor2  gate525(.a(N50), .b(N213), .O(gate63inter0));
  nand2 gate526(.a(gate63inter0), .b(s_52), .O(gate63inter1));
  and2  gate527(.a(N50), .b(N213), .O(gate63inter2));
  inv1  gate528(.a(s_52), .O(gate63inter3));
  inv1  gate529(.a(s_53), .O(gate63inter4));
  nand2 gate530(.a(gate63inter4), .b(gate63inter3), .O(gate63inter5));
  nor2  gate531(.a(gate63inter5), .b(gate63inter2), .O(gate63inter6));
  inv1  gate532(.a(N213), .O(gate63inter7));
  inv1  gate533(.a(N50), .O(gate63inter8));
  nand2 gate534(.a(gate63inter8), .b(gate63inter7), .O(gate63inter9));
  nand2 gate535(.a(s_53), .b(gate63inter3), .O(gate63inter10));
  nor2  gate536(.a(gate63inter10), .b(gate63inter9), .O(gate63inter11));
  nor2  gate537(.a(gate63inter11), .b(gate63inter6), .O(gate63inter12));
  nand2 gate538(.a(gate63inter12), .b(gate63inter1), .O(N255));

  xor2  gate623(.a(N63), .b(N213), .O(gate64inter0));
  nand2 gate624(.a(gate64inter0), .b(s_66), .O(gate64inter1));
  and2  gate625(.a(N63), .b(N213), .O(gate64inter2));
  inv1  gate626(.a(s_66), .O(gate64inter3));
  inv1  gate627(.a(s_67), .O(gate64inter4));
  nand2 gate628(.a(gate64inter4), .b(gate64inter3), .O(gate64inter5));
  nor2  gate629(.a(gate64inter5), .b(gate64inter2), .O(gate64inter6));
  inv1  gate630(.a(N213), .O(gate64inter7));
  inv1  gate631(.a(N63), .O(gate64inter8));
  nand2 gate632(.a(gate64inter8), .b(gate64inter7), .O(gate64inter9));
  nand2 gate633(.a(s_67), .b(gate64inter3), .O(gate64inter10));
  nor2  gate634(.a(gate64inter10), .b(gate64inter9), .O(gate64inter11));
  nor2  gate635(.a(gate64inter11), .b(gate64inter6), .O(gate64inter12));
  nand2 gate636(.a(gate64inter12), .b(gate64inter1), .O(N256));

  xor2  gate469(.a(N76), .b(N213), .O(gate65inter0));
  nand2 gate470(.a(gate65inter0), .b(s_44), .O(gate65inter1));
  and2  gate471(.a(N76), .b(N213), .O(gate65inter2));
  inv1  gate472(.a(s_44), .O(gate65inter3));
  inv1  gate473(.a(s_45), .O(gate65inter4));
  nand2 gate474(.a(gate65inter4), .b(gate65inter3), .O(gate65inter5));
  nor2  gate475(.a(gate65inter5), .b(gate65inter2), .O(gate65inter6));
  inv1  gate476(.a(N213), .O(gate65inter7));
  inv1  gate477(.a(N76), .O(gate65inter8));
  nand2 gate478(.a(gate65inter8), .b(gate65inter7), .O(gate65inter9));
  nand2 gate479(.a(s_45), .b(gate65inter3), .O(gate65inter10));
  nor2  gate480(.a(gate65inter10), .b(gate65inter9), .O(gate65inter11));
  nor2  gate481(.a(gate65inter11), .b(gate65inter6), .O(gate65inter12));
  nand2 gate482(.a(gate65inter12), .b(gate65inter1), .O(N257));
nand2 gate66( .a(N213), .b(N89), .O(N258) );
nand2 gate67( .a(N213), .b(N102), .O(N259) );
nand2 gate68( .a(N224), .b(N157), .O(N260) );

  xor2  gate385(.a(N158), .b(N224), .O(gate69inter0));
  nand2 gate386(.a(gate69inter0), .b(s_32), .O(gate69inter1));
  and2  gate387(.a(N158), .b(N224), .O(gate69inter2));
  inv1  gate388(.a(s_32), .O(gate69inter3));
  inv1  gate389(.a(s_33), .O(gate69inter4));
  nand2 gate390(.a(gate69inter4), .b(gate69inter3), .O(gate69inter5));
  nor2  gate391(.a(gate69inter5), .b(gate69inter2), .O(gate69inter6));
  inv1  gate392(.a(N224), .O(gate69inter7));
  inv1  gate393(.a(N158), .O(gate69inter8));
  nand2 gate394(.a(gate69inter8), .b(gate69inter7), .O(gate69inter9));
  nand2 gate395(.a(s_33), .b(gate69inter3), .O(gate69inter10));
  nor2  gate396(.a(gate69inter10), .b(gate69inter9), .O(gate69inter11));
  nor2  gate397(.a(gate69inter11), .b(gate69inter6), .O(gate69inter12));
  nand2 gate398(.a(gate69inter12), .b(gate69inter1), .O(N263));

  xor2  gate259(.a(N183), .b(N227), .O(gate70inter0));
  nand2 gate260(.a(gate70inter0), .b(s_14), .O(gate70inter1));
  and2  gate261(.a(N183), .b(N227), .O(gate70inter2));
  inv1  gate262(.a(s_14), .O(gate70inter3));
  inv1  gate263(.a(s_15), .O(gate70inter4));
  nand2 gate264(.a(gate70inter4), .b(gate70inter3), .O(gate70inter5));
  nor2  gate265(.a(gate70inter5), .b(gate70inter2), .O(gate70inter6));
  inv1  gate266(.a(N227), .O(gate70inter7));
  inv1  gate267(.a(N183), .O(gate70inter8));
  nand2 gate268(.a(gate70inter8), .b(gate70inter7), .O(gate70inter9));
  nand2 gate269(.a(s_15), .b(gate70inter3), .O(gate70inter10));
  nor2  gate270(.a(gate70inter10), .b(gate70inter9), .O(gate70inter11));
  nor2  gate271(.a(gate70inter11), .b(gate70inter6), .O(gate70inter12));
  nand2 gate272(.a(gate70inter12), .b(gate70inter1), .O(N264));

  xor2  gate161(.a(N185), .b(N230), .O(gate71inter0));
  nand2 gate162(.a(gate71inter0), .b(s_0), .O(gate71inter1));
  and2  gate163(.a(N185), .b(N230), .O(gate71inter2));
  inv1  gate164(.a(s_0), .O(gate71inter3));
  inv1  gate165(.a(s_1), .O(gate71inter4));
  nand2 gate166(.a(gate71inter4), .b(gate71inter3), .O(gate71inter5));
  nor2  gate167(.a(gate71inter5), .b(gate71inter2), .O(gate71inter6));
  inv1  gate168(.a(N230), .O(gate71inter7));
  inv1  gate169(.a(N185), .O(gate71inter8));
  nand2 gate170(.a(gate71inter8), .b(gate71inter7), .O(gate71inter9));
  nand2 gate171(.a(s_1), .b(gate71inter3), .O(gate71inter10));
  nor2  gate172(.a(gate71inter10), .b(gate71inter9), .O(gate71inter11));
  nor2  gate173(.a(gate71inter11), .b(gate71inter6), .O(gate71inter12));
  nand2 gate174(.a(gate71inter12), .b(gate71inter1), .O(N267));

  xor2  gate203(.a(N187), .b(N233), .O(gate72inter0));
  nand2 gate204(.a(gate72inter0), .b(s_6), .O(gate72inter1));
  and2  gate205(.a(N187), .b(N233), .O(gate72inter2));
  inv1  gate206(.a(s_6), .O(gate72inter3));
  inv1  gate207(.a(s_7), .O(gate72inter4));
  nand2 gate208(.a(gate72inter4), .b(gate72inter3), .O(gate72inter5));
  nor2  gate209(.a(gate72inter5), .b(gate72inter2), .O(gate72inter6));
  inv1  gate210(.a(N233), .O(gate72inter7));
  inv1  gate211(.a(N187), .O(gate72inter8));
  nand2 gate212(.a(gate72inter8), .b(gate72inter7), .O(gate72inter9));
  nand2 gate213(.a(s_7), .b(gate72inter3), .O(gate72inter10));
  nor2  gate214(.a(gate72inter10), .b(gate72inter9), .O(gate72inter11));
  nor2  gate215(.a(gate72inter11), .b(gate72inter6), .O(gate72inter12));
  nand2 gate216(.a(gate72inter12), .b(gate72inter1), .O(N270));
nand2 gate73( .a(N236), .b(N189), .O(N273) );

  xor2  gate483(.a(N191), .b(N239), .O(gate74inter0));
  nand2 gate484(.a(gate74inter0), .b(s_46), .O(gate74inter1));
  and2  gate485(.a(N191), .b(N239), .O(gate74inter2));
  inv1  gate486(.a(s_46), .O(gate74inter3));
  inv1  gate487(.a(s_47), .O(gate74inter4));
  nand2 gate488(.a(gate74inter4), .b(gate74inter3), .O(gate74inter5));
  nor2  gate489(.a(gate74inter5), .b(gate74inter2), .O(gate74inter6));
  inv1  gate490(.a(N239), .O(gate74inter7));
  inv1  gate491(.a(N191), .O(gate74inter8));
  nand2 gate492(.a(gate74inter8), .b(gate74inter7), .O(gate74inter9));
  nand2 gate493(.a(s_47), .b(gate74inter3), .O(gate74inter10));
  nor2  gate494(.a(gate74inter10), .b(gate74inter9), .O(gate74inter11));
  nor2  gate495(.a(gate74inter11), .b(gate74inter6), .O(gate74inter12));
  nand2 gate496(.a(gate74inter12), .b(gate74inter1), .O(N276));
nand2 gate75( .a(N243), .b(N193), .O(N279) );
nand2 gate76( .a(N247), .b(N195), .O(N282) );

  xor2  gate343(.a(N197), .b(N251), .O(gate77inter0));
  nand2 gate344(.a(gate77inter0), .b(s_26), .O(gate77inter1));
  and2  gate345(.a(N197), .b(N251), .O(gate77inter2));
  inv1  gate346(.a(s_26), .O(gate77inter3));
  inv1  gate347(.a(s_27), .O(gate77inter4));
  nand2 gate348(.a(gate77inter4), .b(gate77inter3), .O(gate77inter5));
  nor2  gate349(.a(gate77inter5), .b(gate77inter2), .O(gate77inter6));
  inv1  gate350(.a(N251), .O(gate77inter7));
  inv1  gate351(.a(N197), .O(gate77inter8));
  nand2 gate352(.a(gate77inter8), .b(gate77inter7), .O(gate77inter9));
  nand2 gate353(.a(s_27), .b(gate77inter3), .O(gate77inter10));
  nor2  gate354(.a(gate77inter10), .b(gate77inter9), .O(gate77inter11));
  nor2  gate355(.a(gate77inter11), .b(gate77inter6), .O(gate77inter12));
  nand2 gate356(.a(gate77inter12), .b(gate77inter1), .O(N285));
nand2 gate78( .a(N227), .b(N184), .O(N288) );

  xor2  gate539(.a(N186), .b(N230), .O(gate79inter0));
  nand2 gate540(.a(gate79inter0), .b(s_54), .O(gate79inter1));
  and2  gate541(.a(N186), .b(N230), .O(gate79inter2));
  inv1  gate542(.a(s_54), .O(gate79inter3));
  inv1  gate543(.a(s_55), .O(gate79inter4));
  nand2 gate544(.a(gate79inter4), .b(gate79inter3), .O(gate79inter5));
  nor2  gate545(.a(gate79inter5), .b(gate79inter2), .O(gate79inter6));
  inv1  gate546(.a(N230), .O(gate79inter7));
  inv1  gate547(.a(N186), .O(gate79inter8));
  nand2 gate548(.a(gate79inter8), .b(gate79inter7), .O(gate79inter9));
  nand2 gate549(.a(s_55), .b(gate79inter3), .O(gate79inter10));
  nor2  gate550(.a(gate79inter10), .b(gate79inter9), .O(gate79inter11));
  nor2  gate551(.a(gate79inter11), .b(gate79inter6), .O(gate79inter12));
  nand2 gate552(.a(gate79inter12), .b(gate79inter1), .O(N289));
nand2 gate80( .a(N233), .b(N188), .O(N290) );
nand2 gate81( .a(N236), .b(N190), .O(N291) );
nand2 gate82( .a(N239), .b(N192), .O(N292) );

  xor2  gate175(.a(N194), .b(N243), .O(gate83inter0));
  nand2 gate176(.a(gate83inter0), .b(s_2), .O(gate83inter1));
  and2  gate177(.a(N194), .b(N243), .O(gate83inter2));
  inv1  gate178(.a(s_2), .O(gate83inter3));
  inv1  gate179(.a(s_3), .O(gate83inter4));
  nand2 gate180(.a(gate83inter4), .b(gate83inter3), .O(gate83inter5));
  nor2  gate181(.a(gate83inter5), .b(gate83inter2), .O(gate83inter6));
  inv1  gate182(.a(N243), .O(gate83inter7));
  inv1  gate183(.a(N194), .O(gate83inter8));
  nand2 gate184(.a(gate83inter8), .b(gate83inter7), .O(gate83inter9));
  nand2 gate185(.a(s_3), .b(gate83inter3), .O(gate83inter10));
  nor2  gate186(.a(gate83inter10), .b(gate83inter9), .O(gate83inter11));
  nor2  gate187(.a(gate83inter11), .b(gate83inter6), .O(gate83inter12));
  nand2 gate188(.a(gate83inter12), .b(gate83inter1), .O(N293));
nand2 gate84( .a(N247), .b(N196), .O(N294) );
nand2 gate85( .a(N251), .b(N198), .O(N295) );
and9 gate86( .a(N260), .b(N264), .c(N267), .d(N270), .e(N273), .f(N276), .g(N279), .h(N282), .i(N285), .O(N296) );
inv1 gate87( .a(N263), .O(N300) );
inv1 gate88( .a(N288), .O(N301) );
inv1 gate89( .a(N289), .O(N302) );
inv1 gate90( .a(N290), .O(N303) );
inv1 gate91( .a(N291), .O(N304) );
inv1 gate92( .a(N292), .O(N305) );
inv1 gate93( .a(N293), .O(N306) );
inv1 gate94( .a(N294), .O(N307) );
inv1 gate95( .a(N295), .O(N308) );
inv1 gate96( .a(N296), .O(N309) );
inv1 gate97( .a(N296), .O(N319) );
inv1 gate98( .a(N296), .O(N329) );
xor2 gate99( .a(N309), .b(N260), .O(N330) );

  xor2  gate511(.a(N264), .b(N309), .O(gate100inter0));
  nand2 gate512(.a(gate100inter0), .b(s_50), .O(gate100inter1));
  and2  gate513(.a(N264), .b(N309), .O(gate100inter2));
  inv1  gate514(.a(s_50), .O(gate100inter3));
  inv1  gate515(.a(s_51), .O(gate100inter4));
  nand2 gate516(.a(gate100inter4), .b(gate100inter3), .O(gate100inter5));
  nor2  gate517(.a(gate100inter5), .b(gate100inter2), .O(gate100inter6));
  inv1  gate518(.a(N309), .O(gate100inter7));
  inv1  gate519(.a(N264), .O(gate100inter8));
  nand2 gate520(.a(gate100inter8), .b(gate100inter7), .O(gate100inter9));
  nand2 gate521(.a(s_51), .b(gate100inter3), .O(gate100inter10));
  nor2  gate522(.a(gate100inter10), .b(gate100inter9), .O(gate100inter11));
  nor2  gate523(.a(gate100inter11), .b(gate100inter6), .O(gate100inter12));
  nand2 gate524(.a(gate100inter12), .b(gate100inter1), .O(N331));
xor2 gate101( .a(N309), .b(N267), .O(N332) );
xor2 gate102( .a(N309), .b(N270), .O(N333) );

  xor2  gate553(.a(N319), .b(N8), .O(gate103inter0));
  nand2 gate554(.a(gate103inter0), .b(s_56), .O(gate103inter1));
  and2  gate555(.a(N319), .b(N8), .O(gate103inter2));
  inv1  gate556(.a(s_56), .O(gate103inter3));
  inv1  gate557(.a(s_57), .O(gate103inter4));
  nand2 gate558(.a(gate103inter4), .b(gate103inter3), .O(gate103inter5));
  nor2  gate559(.a(gate103inter5), .b(gate103inter2), .O(gate103inter6));
  inv1  gate560(.a(N8), .O(gate103inter7));
  inv1  gate561(.a(N319), .O(gate103inter8));
  nand2 gate562(.a(gate103inter8), .b(gate103inter7), .O(gate103inter9));
  nand2 gate563(.a(s_57), .b(gate103inter3), .O(gate103inter10));
  nor2  gate564(.a(gate103inter10), .b(gate103inter9), .O(gate103inter11));
  nor2  gate565(.a(gate103inter11), .b(gate103inter6), .O(gate103inter12));
  nand2 gate566(.a(gate103inter12), .b(gate103inter1), .O(N334));
xor2 gate104( .a(N309), .b(N273), .O(N335) );
nand2 gate105( .a(N319), .b(N21), .O(N336) );

  xor2  gate651(.a(N276), .b(N309), .O(gate106inter0));
  nand2 gate652(.a(gate106inter0), .b(s_70), .O(gate106inter1));
  and2  gate653(.a(N276), .b(N309), .O(gate106inter2));
  inv1  gate654(.a(s_70), .O(gate106inter3));
  inv1  gate655(.a(s_71), .O(gate106inter4));
  nand2 gate656(.a(gate106inter4), .b(gate106inter3), .O(gate106inter5));
  nor2  gate657(.a(gate106inter5), .b(gate106inter2), .O(gate106inter6));
  inv1  gate658(.a(N309), .O(gate106inter7));
  inv1  gate659(.a(N276), .O(gate106inter8));
  nand2 gate660(.a(gate106inter8), .b(gate106inter7), .O(gate106inter9));
  nand2 gate661(.a(s_71), .b(gate106inter3), .O(gate106inter10));
  nor2  gate662(.a(gate106inter10), .b(gate106inter9), .O(gate106inter11));
  nor2  gate663(.a(gate106inter11), .b(gate106inter6), .O(gate106inter12));
  nand2 gate664(.a(gate106inter12), .b(gate106inter1), .O(N337));

  xor2  gate315(.a(N34), .b(N319), .O(gate107inter0));
  nand2 gate316(.a(gate107inter0), .b(s_22), .O(gate107inter1));
  and2  gate317(.a(N34), .b(N319), .O(gate107inter2));
  inv1  gate318(.a(s_22), .O(gate107inter3));
  inv1  gate319(.a(s_23), .O(gate107inter4));
  nand2 gate320(.a(gate107inter4), .b(gate107inter3), .O(gate107inter5));
  nor2  gate321(.a(gate107inter5), .b(gate107inter2), .O(gate107inter6));
  inv1  gate322(.a(N319), .O(gate107inter7));
  inv1  gate323(.a(N34), .O(gate107inter8));
  nand2 gate324(.a(gate107inter8), .b(gate107inter7), .O(gate107inter9));
  nand2 gate325(.a(s_23), .b(gate107inter3), .O(gate107inter10));
  nor2  gate326(.a(gate107inter10), .b(gate107inter9), .O(gate107inter11));
  nor2  gate327(.a(gate107inter11), .b(gate107inter6), .O(gate107inter12));
  nand2 gate328(.a(gate107inter12), .b(gate107inter1), .O(N338));
xor2 gate108( .a(N309), .b(N279), .O(N339) );
nand2 gate109( .a(N319), .b(N47), .O(N340) );
xor2 gate110( .a(N309), .b(N282), .O(N341) );
nand2 gate111( .a(N319), .b(N60), .O(N342) );

  xor2  gate441(.a(N285), .b(N309), .O(gate112inter0));
  nand2 gate442(.a(gate112inter0), .b(s_40), .O(gate112inter1));
  and2  gate443(.a(N285), .b(N309), .O(gate112inter2));
  inv1  gate444(.a(s_40), .O(gate112inter3));
  inv1  gate445(.a(s_41), .O(gate112inter4));
  nand2 gate446(.a(gate112inter4), .b(gate112inter3), .O(gate112inter5));
  nor2  gate447(.a(gate112inter5), .b(gate112inter2), .O(gate112inter6));
  inv1  gate448(.a(N309), .O(gate112inter7));
  inv1  gate449(.a(N285), .O(gate112inter8));
  nand2 gate450(.a(gate112inter8), .b(gate112inter7), .O(gate112inter9));
  nand2 gate451(.a(s_41), .b(gate112inter3), .O(gate112inter10));
  nor2  gate452(.a(gate112inter10), .b(gate112inter9), .O(gate112inter11));
  nor2  gate453(.a(gate112inter11), .b(gate112inter6), .O(gate112inter12));
  nand2 gate454(.a(gate112inter12), .b(gate112inter1), .O(N343));
nand2 gate113( .a(N319), .b(N73), .O(N344) );
nand2 gate114( .a(N319), .b(N86), .O(N345) );

  xor2  gate329(.a(N99), .b(N319), .O(gate115inter0));
  nand2 gate330(.a(gate115inter0), .b(s_24), .O(gate115inter1));
  and2  gate331(.a(N99), .b(N319), .O(gate115inter2));
  inv1  gate332(.a(s_24), .O(gate115inter3));
  inv1  gate333(.a(s_25), .O(gate115inter4));
  nand2 gate334(.a(gate115inter4), .b(gate115inter3), .O(gate115inter5));
  nor2  gate335(.a(gate115inter5), .b(gate115inter2), .O(gate115inter6));
  inv1  gate336(.a(N319), .O(gate115inter7));
  inv1  gate337(.a(N99), .O(gate115inter8));
  nand2 gate338(.a(gate115inter8), .b(gate115inter7), .O(gate115inter9));
  nand2 gate339(.a(s_25), .b(gate115inter3), .O(gate115inter10));
  nor2  gate340(.a(gate115inter10), .b(gate115inter9), .O(gate115inter11));
  nor2  gate341(.a(gate115inter11), .b(gate115inter6), .O(gate115inter12));
  nand2 gate342(.a(gate115inter12), .b(gate115inter1), .O(N346));
nand2 gate116( .a(N319), .b(N112), .O(N347) );

  xor2  gate217(.a(N300), .b(N330), .O(gate117inter0));
  nand2 gate218(.a(gate117inter0), .b(s_8), .O(gate117inter1));
  and2  gate219(.a(N300), .b(N330), .O(gate117inter2));
  inv1  gate220(.a(s_8), .O(gate117inter3));
  inv1  gate221(.a(s_9), .O(gate117inter4));
  nand2 gate222(.a(gate117inter4), .b(gate117inter3), .O(gate117inter5));
  nor2  gate223(.a(gate117inter5), .b(gate117inter2), .O(gate117inter6));
  inv1  gate224(.a(N330), .O(gate117inter7));
  inv1  gate225(.a(N300), .O(gate117inter8));
  nand2 gate226(.a(gate117inter8), .b(gate117inter7), .O(gate117inter9));
  nand2 gate227(.a(s_9), .b(gate117inter3), .O(gate117inter10));
  nor2  gate228(.a(gate117inter10), .b(gate117inter9), .O(gate117inter11));
  nor2  gate229(.a(gate117inter11), .b(gate117inter6), .O(gate117inter12));
  nand2 gate230(.a(gate117inter12), .b(gate117inter1), .O(N348));
nand2 gate118( .a(N331), .b(N301), .O(N349) );
nand2 gate119( .a(N332), .b(N302), .O(N350) );
nand2 gate120( .a(N333), .b(N303), .O(N351) );

  xor2  gate371(.a(N304), .b(N335), .O(gate121inter0));
  nand2 gate372(.a(gate121inter0), .b(s_30), .O(gate121inter1));
  and2  gate373(.a(N304), .b(N335), .O(gate121inter2));
  inv1  gate374(.a(s_30), .O(gate121inter3));
  inv1  gate375(.a(s_31), .O(gate121inter4));
  nand2 gate376(.a(gate121inter4), .b(gate121inter3), .O(gate121inter5));
  nor2  gate377(.a(gate121inter5), .b(gate121inter2), .O(gate121inter6));
  inv1  gate378(.a(N335), .O(gate121inter7));
  inv1  gate379(.a(N304), .O(gate121inter8));
  nand2 gate380(.a(gate121inter8), .b(gate121inter7), .O(gate121inter9));
  nand2 gate381(.a(s_31), .b(gate121inter3), .O(gate121inter10));
  nor2  gate382(.a(gate121inter10), .b(gate121inter9), .O(gate121inter11));
  nor2  gate383(.a(gate121inter11), .b(gate121inter6), .O(gate121inter12));
  nand2 gate384(.a(gate121inter12), .b(gate121inter1), .O(N352));

  xor2  gate567(.a(N305), .b(N337), .O(gate122inter0));
  nand2 gate568(.a(gate122inter0), .b(s_58), .O(gate122inter1));
  and2  gate569(.a(N305), .b(N337), .O(gate122inter2));
  inv1  gate570(.a(s_58), .O(gate122inter3));
  inv1  gate571(.a(s_59), .O(gate122inter4));
  nand2 gate572(.a(gate122inter4), .b(gate122inter3), .O(gate122inter5));
  nor2  gate573(.a(gate122inter5), .b(gate122inter2), .O(gate122inter6));
  inv1  gate574(.a(N337), .O(gate122inter7));
  inv1  gate575(.a(N305), .O(gate122inter8));
  nand2 gate576(.a(gate122inter8), .b(gate122inter7), .O(gate122inter9));
  nand2 gate577(.a(s_59), .b(gate122inter3), .O(gate122inter10));
  nor2  gate578(.a(gate122inter10), .b(gate122inter9), .O(gate122inter11));
  nor2  gate579(.a(gate122inter11), .b(gate122inter6), .O(gate122inter12));
  nand2 gate580(.a(gate122inter12), .b(gate122inter1), .O(N353));
nand2 gate123( .a(N339), .b(N306), .O(N354) );
nand2 gate124( .a(N341), .b(N307), .O(N355) );
nand2 gate125( .a(N343), .b(N308), .O(N356) );
and9 gate126( .a(N348), .b(N349), .c(N350), .d(N351), .e(N352), .f(N353), .g(N354), .h(N355), .i(N356), .O(N357) );
inv1 gate127( .a(N357), .O(N360) );
inv1 gate128( .a(N357), .O(N370) );
nand2 gate129( .a(N14), .b(N360), .O(N371) );

  xor2  gate245(.a(N27), .b(N360), .O(gate130inter0));
  nand2 gate246(.a(gate130inter0), .b(s_12), .O(gate130inter1));
  and2  gate247(.a(N27), .b(N360), .O(gate130inter2));
  inv1  gate248(.a(s_12), .O(gate130inter3));
  inv1  gate249(.a(s_13), .O(gate130inter4));
  nand2 gate250(.a(gate130inter4), .b(gate130inter3), .O(gate130inter5));
  nor2  gate251(.a(gate130inter5), .b(gate130inter2), .O(gate130inter6));
  inv1  gate252(.a(N360), .O(gate130inter7));
  inv1  gate253(.a(N27), .O(gate130inter8));
  nand2 gate254(.a(gate130inter8), .b(gate130inter7), .O(gate130inter9));
  nand2 gate255(.a(s_13), .b(gate130inter3), .O(gate130inter10));
  nor2  gate256(.a(gate130inter10), .b(gate130inter9), .O(gate130inter11));
  nor2  gate257(.a(gate130inter11), .b(gate130inter6), .O(gate130inter12));
  nand2 gate258(.a(gate130inter12), .b(gate130inter1), .O(N372));
nand2 gate131( .a(N360), .b(N40), .O(N373) );

  xor2  gate189(.a(N53), .b(N360), .O(gate132inter0));
  nand2 gate190(.a(gate132inter0), .b(s_4), .O(gate132inter1));
  and2  gate191(.a(N53), .b(N360), .O(gate132inter2));
  inv1  gate192(.a(s_4), .O(gate132inter3));
  inv1  gate193(.a(s_5), .O(gate132inter4));
  nand2 gate194(.a(gate132inter4), .b(gate132inter3), .O(gate132inter5));
  nor2  gate195(.a(gate132inter5), .b(gate132inter2), .O(gate132inter6));
  inv1  gate196(.a(N360), .O(gate132inter7));
  inv1  gate197(.a(N53), .O(gate132inter8));
  nand2 gate198(.a(gate132inter8), .b(gate132inter7), .O(gate132inter9));
  nand2 gate199(.a(s_5), .b(gate132inter3), .O(gate132inter10));
  nor2  gate200(.a(gate132inter10), .b(gate132inter9), .O(gate132inter11));
  nor2  gate201(.a(gate132inter11), .b(gate132inter6), .O(gate132inter12));
  nand2 gate202(.a(gate132inter12), .b(gate132inter1), .O(N374));
nand2 gate133( .a(N360), .b(N66), .O(N375) );
nand2 gate134( .a(N360), .b(N79), .O(N376) );
nand2 gate135( .a(N360), .b(N92), .O(N377) );
nand2 gate136( .a(N360), .b(N105), .O(N378) );
nand2 gate137( .a(N360), .b(N115), .O(N379) );
nand4 gate138( .a(N4), .b(N242), .c(N334), .d(N371), .O(N380) );
nand4 gate139( .a(N246), .b(N336), .c(N372), .d(N17), .O(N381) );
nand4 gate140( .a(N250), .b(N338), .c(N373), .d(N30), .O(N386) );
nand4 gate141( .a(N254), .b(N340), .c(N374), .d(N43), .O(N393) );
nand4 gate142( .a(N255), .b(N342), .c(N375), .d(N56), .O(N399) );
nand4 gate143( .a(N256), .b(N344), .c(N376), .d(N69), .O(N404) );
nand4 gate144( .a(N257), .b(N345), .c(N377), .d(N82), .O(N407) );
nand4 gate145( .a(N258), .b(N346), .c(N378), .d(N95), .O(N411) );
nand4 gate146( .a(N259), .b(N347), .c(N379), .d(N108), .O(N414) );
inv1 gate147( .a(N380), .O(N415) );
and8 gate148( .a(N381), .b(N386), .c(N393), .d(N399), .e(N404), .f(N407), .g(N411), .h(N414), .O(N416) );
inv1 gate149( .a(N393), .O(N417) );
inv1 gate150( .a(N404), .O(N418) );
inv1 gate151( .a(N407), .O(N419) );
inv1 gate152( .a(N411), .O(N420) );
nor2 gate153( .a(N415), .b(N416), .O(N421) );
nand2 gate154( .a(N386), .b(N417), .O(N422) );
nand4 gate155( .a(N386), .b(N393), .c(N418), .d(N399), .O(N425) );
nand3 gate156( .a(N399), .b(N393), .c(N419), .O(N428) );
nand4 gate157( .a(N386), .b(N393), .c(N407), .d(N420), .O(N429) );
nand4 gate158( .a(N381), .b(N386), .c(N422), .d(N399), .O(N430) );
nand4 gate159( .a(N381), .b(N386), .c(N425), .d(N428), .O(N431) );
nand4 gate160( .a(N381), .b(N422), .c(N425), .d(N429), .O(N432) );

endmodule