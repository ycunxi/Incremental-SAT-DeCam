module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);

input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;//RE__PI;

input s_0,s_1;//RE__ALLOW(00,01,10,11);
input s_2,s_3;//RE__ALLOW(00,01,10,11);
input s_4,s_5;//RE__ALLOW(00,01,10,11);
input s_6,s_7;//RE__ALLOW(00,01,10,11);
input s_8,s_9;//RE__ALLOW(00,01,10,11);
input s_10,s_11;//RE__ALLOW(00,01,10,11);
input s_12,s_13;//RE__ALLOW(00,01,10,11);
input s_14,s_15;//RE__ALLOW(00,01,10,11);
input s_16,s_17;//RE__ALLOW(00,01,10,11);
input s_18,s_19;//RE__ALLOW(00,01,10,11);
input s_20,s_21;//RE__ALLOW(00,01,10,11);
input s_22,s_23;//RE__ALLOW(00,01,10,11);
input s_24,s_25;//RE__ALLOW(00,01,10,11);
input s_26,s_27;//RE__ALLOW(00,01,10,11);
input s_28,s_29;//RE__ALLOW(00,01,10,11);
input s_30,s_31;//RE__ALLOW(00,01,10,11);
input s_32,s_33;//RE__ALLOW(00,01,10,11);
input s_34,s_35;//RE__ALLOW(00,01,10,11);
input s_36,s_37;//RE__ALLOW(00,01,10,11);
input s_38,s_39;//RE__ALLOW(00,01,10,11);
input s_40,s_41;//RE__ALLOW(00,01,10,11);
input s_42,s_43;//RE__ALLOW(00,01,10,11);
input s_44,s_45;//RE__ALLOW(00,01,10,11);
input s_46,s_47;//RE__ALLOW(00,01,10,11);
input s_48,s_49;//RE__ALLOW(00,01,10,11);
input s_50,s_51;//RE__ALLOW(00,01,10,11);
input s_52,s_53;//RE__ALLOW(00,01,10,11);
input s_54,s_55;//RE__ALLOW(00,01,10,11);
input s_56,s_57;//RE__ALLOW(00,01,10,11);
input s_58,s_59;//RE__ALLOW(00,01,10,11);
input s_60,s_61;//RE__ALLOW(00,01,10,11);
input s_62,s_63;//RE__ALLOW(00,01,10,11);
input s_64,s_65;//RE__ALLOW(00,01,10,11);
input s_66,s_67;//RE__ALLOW(00,01,10,11);
input s_68,s_69;//RE__ALLOW(00,01,10,11);
input s_70,s_71;//RE__ALLOW(00,01,10,11);
input s_72,s_73;//RE__ALLOW(00,01,10,11);
input s_74,s_75;//RE__ALLOW(00,01,10,11);
input s_76,s_77;//RE__ALLOW(00,01,10,11);
input s_78,s_79;//RE__ALLOW(00,01,10,11);
input s_80,s_81;//RE__ALLOW(00,01,10,11);
input s_82,s_83;//RE__ALLOW(00,01,10,11);
input s_84,s_85;//RE__ALLOW(00,01,10,11);
input s_86,s_87;//RE__ALLOW(00,01,10,11);
input s_88,s_89;//RE__ALLOW(00,01,10,11);
input s_90,s_91;//RE__ALLOW(00,01,10,11);
input s_92,s_93;//RE__ALLOW(00,01,10,11);
input s_94,s_95;//RE__ALLOW(00,01,10,11);
input s_96,s_97;//RE__ALLOW(00,01,10,11);
input s_98,s_99;//RE__ALLOW(00,01,10,11);
input s_100,s_101;//RE__ALLOW(00,01,10,11);
input s_102,s_103;//RE__ALLOW(00,01,10,11);
input s_104,s_105;//RE__ALLOW(00,01,10,11);
input s_106,s_107;//RE__ALLOW(00,01,10,11);
input s_108,s_109;//RE__ALLOW(00,01,10,11);
input s_110,s_111;//RE__ALLOW(00,01,10,11);
input s_112,s_113;//RE__ALLOW(00,01,10,11);
input s_114,s_115;//RE__ALLOW(00,01,10,11);
input s_116,s_117;//RE__ALLOW(00,01,10,11);
input s_118,s_119;//RE__ALLOW(00,01,10,11);
input s_120,s_121;//RE__ALLOW(00,01,10,11);
input s_122,s_123;//RE__ALLOW(00,01,10,11);
input s_124,s_125;//RE__ALLOW(00,01,10,11);
input s_126,s_127;//RE__ALLOW(00,01,10,11);
input s_128,s_129;//RE__ALLOW(00,01,10,11);
input s_130,s_131;//RE__ALLOW(00,01,10,11);
input s_132,s_133;//RE__ALLOW(00,01,10,11);
input s_134,s_135;//RE__ALLOW(00,01,10,11);
input s_136,s_137;//RE__ALLOW(00,01,10,11);
input s_138,s_139;//RE__ALLOW(00,01,10,11);
input s_140,s_141;//RE__ALLOW(00,01,10,11);
input s_142,s_143;//RE__ALLOW(00,01,10,11);
input s_144,s_145;//RE__ALLOW(00,01,10,11);
input s_146,s_147;//RE__ALLOW(00,01,10,11);
input s_148,s_149;//RE__ALLOW(00,01,10,11);
input s_150,s_151;//RE__ALLOW(00,01,10,11);
input s_152,s_153;//RE__ALLOW(00,01,10,11);
input s_154,s_155;//RE__ALLOW(00,01,10,11);
input s_156,s_157;//RE__ALLOW(00,01,10,11);
input s_158,s_159;//RE__ALLOW(00,01,10,11);
input s_160,s_161;//RE__ALLOW(00,01,10,11);
input s_162,s_163;//RE__ALLOW(00,01,10,11);
input s_164,s_165;//RE__ALLOW(00,01,10,11);
input s_166,s_167;//RE__ALLOW(00,01,10,11);
input s_168,s_169;//RE__ALLOW(00,01,10,11);
input s_170,s_171;//RE__ALLOW(00,01,10,11);
input s_172,s_173;//RE__ALLOW(00,01,10,11);
input s_174,s_175;//RE__ALLOW(00,01,10,11);
input s_176,s_177;//RE__ALLOW(00,01,10,11);
input s_178,s_179;//RE__ALLOW(00,01,10,11);
input s_180,s_181;//RE__ALLOW(00,01,10,11);
input s_182,s_183;//RE__ALLOW(00,01,10,11);
input s_184,s_185;//RE__ALLOW(00,01,10,11);
input s_186,s_187;//RE__ALLOW(00,01,10,11);
input s_188,s_189;//RE__ALLOW(00,01,10,11);
input s_190,s_191;//RE__ALLOW(00,01,10,11);
input s_192,s_193;//RE__ALLOW(00,01,10,11);
input s_194,s_195;//RE__ALLOW(00,01,10,11);
input s_196,s_197;//RE__ALLOW(00,01,10,11);
input s_198,s_199;//RE__ALLOW(00,01,10,11);
input s_200,s_201;//RE__ALLOW(00,01,10,11);
input s_202,s_203;//RE__ALLOW(00,01,10,11);
input s_204,s_205;//RE__ALLOW(00,01,10,11);
input s_206,s_207;//RE__ALLOW(00,01,10,11);
input s_208,s_209;//RE__ALLOW(00,01,10,11);
input s_210,s_211;//RE__ALLOW(00,01,10,11);
input s_212,s_213;//RE__ALLOW(00,01,10,11);
input s_214,s_215;//RE__ALLOW(00,01,10,11);
input s_216,s_217;//RE__ALLOW(00,01,10,11);
input s_218,s_219;//RE__ALLOW(00,01,10,11);
input s_220,s_221;//RE__ALLOW(00,01,10,11);
input s_222,s_223;//RE__ALLOW(00,01,10,11);
input s_224,s_225;//RE__ALLOW(00,01,10,11);
input s_226,s_227;//RE__ALLOW(00,01,10,11);
input s_228,s_229;//RE__ALLOW(00,01,10,11);
input s_230,s_231;//RE__ALLOW(00,01,10,11);
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;

  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate86inter0, gate86inter1, gate86inter2, gate86inter3, gate86inter4, gate86inter5, gate86inter6, gate86inter7, gate86inter8, gate86inter9, gate86inter10, gate86inter11, gate86inter12, gate292inter0, gate292inter1, gate292inter2, gate292inter3, gate292inter4, gate292inter5, gate292inter6, gate292inter7, gate292inter8, gate292inter9, gate292inter10, gate292inter11, gate292inter12, gate447inter0, gate447inter1, gate447inter2, gate447inter3, gate447inter4, gate447inter5, gate447inter6, gate447inter7, gate447inter8, gate447inter9, gate447inter10, gate447inter11, gate447inter12, gate193inter0, gate193inter1, gate193inter2, gate193inter3, gate193inter4, gate193inter5, gate193inter6, gate193inter7, gate193inter8, gate193inter9, gate193inter10, gate193inter11, gate193inter12, gate145inter0, gate145inter1, gate145inter2, gate145inter3, gate145inter4, gate145inter5, gate145inter6, gate145inter7, gate145inter8, gate145inter9, gate145inter10, gate145inter11, gate145inter12, gate464inter0, gate464inter1, gate464inter2, gate464inter3, gate464inter4, gate464inter5, gate464inter6, gate464inter7, gate464inter8, gate464inter9, gate464inter10, gate464inter11, gate464inter12, gate270inter0, gate270inter1, gate270inter2, gate270inter3, gate270inter4, gate270inter5, gate270inter6, gate270inter7, gate270inter8, gate270inter9, gate270inter10, gate270inter11, gate270inter12, gate494inter0, gate494inter1, gate494inter2, gate494inter3, gate494inter4, gate494inter5, gate494inter6, gate494inter7, gate494inter8, gate494inter9, gate494inter10, gate494inter11, gate494inter12, gate111inter0, gate111inter1, gate111inter2, gate111inter3, gate111inter4, gate111inter5, gate111inter6, gate111inter7, gate111inter8, gate111inter9, gate111inter10, gate111inter11, gate111inter12, gate445inter0, gate445inter1, gate445inter2, gate445inter3, gate445inter4, gate445inter5, gate445inter6, gate445inter7, gate445inter8, gate445inter9, gate445inter10, gate445inter11, gate445inter12, gate435inter0, gate435inter1, gate435inter2, gate435inter3, gate435inter4, gate435inter5, gate435inter6, gate435inter7, gate435inter8, gate435inter9, gate435inter10, gate435inter11, gate435inter12, gate418inter0, gate418inter1, gate418inter2, gate418inter3, gate418inter4, gate418inter5, gate418inter6, gate418inter7, gate418inter8, gate418inter9, gate418inter10, gate418inter11, gate418inter12, gate293inter0, gate293inter1, gate293inter2, gate293inter3, gate293inter4, gate293inter5, gate293inter6, gate293inter7, gate293inter8, gate293inter9, gate293inter10, gate293inter11, gate293inter12, gate212inter0, gate212inter1, gate212inter2, gate212inter3, gate212inter4, gate212inter5, gate212inter6, gate212inter7, gate212inter8, gate212inter9, gate212inter10, gate212inter11, gate212inter12, gate99inter0, gate99inter1, gate99inter2, gate99inter3, gate99inter4, gate99inter5, gate99inter6, gate99inter7, gate99inter8, gate99inter9, gate99inter10, gate99inter11, gate99inter12, gate261inter0, gate261inter1, gate261inter2, gate261inter3, gate261inter4, gate261inter5, gate261inter6, gate261inter7, gate261inter8, gate261inter9, gate261inter10, gate261inter11, gate261inter12, gate150inter0, gate150inter1, gate150inter2, gate150inter3, gate150inter4, gate150inter5, gate150inter6, gate150inter7, gate150inter8, gate150inter9, gate150inter10, gate150inter11, gate150inter12, gate226inter0, gate226inter1, gate226inter2, gate226inter3, gate226inter4, gate226inter5, gate226inter6, gate226inter7, gate226inter8, gate226inter9, gate226inter10, gate226inter11, gate226inter12, gate64inter0, gate64inter1, gate64inter2, gate64inter3, gate64inter4, gate64inter5, gate64inter6, gate64inter7, gate64inter8, gate64inter9, gate64inter10, gate64inter11, gate64inter12, gate207inter0, gate207inter1, gate207inter2, gate207inter3, gate207inter4, gate207inter5, gate207inter6, gate207inter7, gate207inter8, gate207inter9, gate207inter10, gate207inter11, gate207inter12, gate143inter0, gate143inter1, gate143inter2, gate143inter3, gate143inter4, gate143inter5, gate143inter6, gate143inter7, gate143inter8, gate143inter9, gate143inter10, gate143inter11, gate143inter12, gate41inter0, gate41inter1, gate41inter2, gate41inter3, gate41inter4, gate41inter5, gate41inter6, gate41inter7, gate41inter8, gate41inter9, gate41inter10, gate41inter11, gate41inter12, gate237inter0, gate237inter1, gate237inter2, gate237inter3, gate237inter4, gate237inter5, gate237inter6, gate237inter7, gate237inter8, gate237inter9, gate237inter10, gate237inter11, gate237inter12, gate403inter0, gate403inter1, gate403inter2, gate403inter3, gate403inter4, gate403inter5, gate403inter6, gate403inter7, gate403inter8, gate403inter9, gate403inter10, gate403inter11, gate403inter12, gate426inter0, gate426inter1, gate426inter2, gate426inter3, gate426inter4, gate426inter5, gate426inter6, gate426inter7, gate426inter8, gate426inter9, gate426inter10, gate426inter11, gate426inter12, gate408inter0, gate408inter1, gate408inter2, gate408inter3, gate408inter4, gate408inter5, gate408inter6, gate408inter7, gate408inter8, gate408inter9, gate408inter10, gate408inter11, gate408inter12, gate499inter0, gate499inter1, gate499inter2, gate499inter3, gate499inter4, gate499inter5, gate499inter6, gate499inter7, gate499inter8, gate499inter9, gate499inter10, gate499inter11, gate499inter12, gate423inter0, gate423inter1, gate423inter2, gate423inter3, gate423inter4, gate423inter5, gate423inter6, gate423inter7, gate423inter8, gate423inter9, gate423inter10, gate423inter11, gate423inter12, gate436inter0, gate436inter1, gate436inter2, gate436inter3, gate436inter4, gate436inter5, gate436inter6, gate436inter7, gate436inter8, gate436inter9, gate436inter10, gate436inter11, gate436inter12, gate250inter0, gate250inter1, gate250inter2, gate250inter3, gate250inter4, gate250inter5, gate250inter6, gate250inter7, gate250inter8, gate250inter9, gate250inter10, gate250inter11, gate250inter12, gate486inter0, gate486inter1, gate486inter2, gate486inter3, gate486inter4, gate486inter5, gate486inter6, gate486inter7, gate486inter8, gate486inter9, gate486inter10, gate486inter11, gate486inter12, gate504inter0, gate504inter1, gate504inter2, gate504inter3, gate504inter4, gate504inter5, gate504inter6, gate504inter7, gate504inter8, gate504inter9, gate504inter10, gate504inter11, gate504inter12, gate431inter0, gate431inter1, gate431inter2, gate431inter3, gate431inter4, gate431inter5, gate431inter6, gate431inter7, gate431inter8, gate431inter9, gate431inter10, gate431inter11, gate431inter12, gate153inter0, gate153inter1, gate153inter2, gate153inter3, gate153inter4, gate153inter5, gate153inter6, gate153inter7, gate153inter8, gate153inter9, gate153inter10, gate153inter11, gate153inter12, gate399inter0, gate399inter1, gate399inter2, gate399inter3, gate399inter4, gate399inter5, gate399inter6, gate399inter7, gate399inter8, gate399inter9, gate399inter10, gate399inter11, gate399inter12, gate454inter0, gate454inter1, gate454inter2, gate454inter3, gate454inter4, gate454inter5, gate454inter6, gate454inter7, gate454inter8, gate454inter9, gate454inter10, gate454inter11, gate454inter12, gate502inter0, gate502inter1, gate502inter2, gate502inter3, gate502inter4, gate502inter5, gate502inter6, gate502inter7, gate502inter8, gate502inter9, gate502inter10, gate502inter11, gate502inter12, gate444inter0, gate444inter1, gate444inter2, gate444inter3, gate444inter4, gate444inter5, gate444inter6, gate444inter7, gate444inter8, gate444inter9, gate444inter10, gate444inter11, gate444inter12, gate161inter0, gate161inter1, gate161inter2, gate161inter3, gate161inter4, gate161inter5, gate161inter6, gate161inter7, gate161inter8, gate161inter9, gate161inter10, gate161inter11, gate161inter12, gate201inter0, gate201inter1, gate201inter2, gate201inter3, gate201inter4, gate201inter5, gate201inter6, gate201inter7, gate201inter8, gate201inter9, gate201inter10, gate201inter11, gate201inter12, gate224inter0, gate224inter1, gate224inter2, gate224inter3, gate224inter4, gate224inter5, gate224inter6, gate224inter7, gate224inter8, gate224inter9, gate224inter10, gate224inter11, gate224inter12, gate108inter0, gate108inter1, gate108inter2, gate108inter3, gate108inter4, gate108inter5, gate108inter6, gate108inter7, gate108inter8, gate108inter9, gate108inter10, gate108inter11, gate108inter12, gate37inter0, gate37inter1, gate37inter2, gate37inter3, gate37inter4, gate37inter5, gate37inter6, gate37inter7, gate37inter8, gate37inter9, gate37inter10, gate37inter11, gate37inter12, gate157inter0, gate157inter1, gate157inter2, gate157inter3, gate157inter4, gate157inter5, gate157inter6, gate157inter7, gate157inter8, gate157inter9, gate157inter10, gate157inter11, gate157inter12, gate215inter0, gate215inter1, gate215inter2, gate215inter3, gate215inter4, gate215inter5, gate215inter6, gate215inter7, gate215inter8, gate215inter9, gate215inter10, gate215inter11, gate215inter12, gate420inter0, gate420inter1, gate420inter2, gate420inter3, gate420inter4, gate420inter5, gate420inter6, gate420inter7, gate420inter8, gate420inter9, gate420inter10, gate420inter11, gate420inter12, gate72inter0, gate72inter1, gate72inter2, gate72inter3, gate72inter4, gate72inter5, gate72inter6, gate72inter7, gate72inter8, gate72inter9, gate72inter10, gate72inter11, gate72inter12, gate10inter0, gate10inter1, gate10inter2, gate10inter3, gate10inter4, gate10inter5, gate10inter6, gate10inter7, gate10inter8, gate10inter9, gate10inter10, gate10inter11, gate10inter12, gate498inter0, gate498inter1, gate498inter2, gate498inter3, gate498inter4, gate498inter5, gate498inter6, gate498inter7, gate498inter8, gate498inter9, gate498inter10, gate498inter11, gate498inter12, gate59inter0, gate59inter1, gate59inter2, gate59inter3, gate59inter4, gate59inter5, gate59inter6, gate59inter7, gate59inter8, gate59inter9, gate59inter10, gate59inter11, gate59inter12, gate414inter0, gate414inter1, gate414inter2, gate414inter3, gate414inter4, gate414inter5, gate414inter6, gate414inter7, gate414inter8, gate414inter9, gate414inter10, gate414inter11, gate414inter12, gate24inter0, gate24inter1, gate24inter2, gate24inter3, gate24inter4, gate24inter5, gate24inter6, gate24inter7, gate24inter8, gate24inter9, gate24inter10, gate24inter11, gate24inter12, gate254inter0, gate254inter1, gate254inter2, gate254inter3, gate254inter4, gate254inter5, gate254inter6, gate254inter7, gate254inter8, gate254inter9, gate254inter10, gate254inter11, gate254inter12, gate222inter0, gate222inter1, gate222inter2, gate222inter3, gate222inter4, gate222inter5, gate222inter6, gate222inter7, gate222inter8, gate222inter9, gate222inter10, gate222inter11, gate222inter12, gate181inter0, gate181inter1, gate181inter2, gate181inter3, gate181inter4, gate181inter5, gate181inter6, gate181inter7, gate181inter8, gate181inter9, gate181inter10, gate181inter11, gate181inter12, gate467inter0, gate467inter1, gate467inter2, gate467inter3, gate467inter4, gate467inter5, gate467inter6, gate467inter7, gate467inter8, gate467inter9, gate467inter10, gate467inter11, gate467inter12, gate514inter0, gate514inter1, gate514inter2, gate514inter3, gate514inter4, gate514inter5, gate514inter6, gate514inter7, gate514inter8, gate514inter9, gate514inter10, gate514inter11, gate514inter12, gate53inter0, gate53inter1, gate53inter2, gate53inter3, gate53inter4, gate53inter5, gate53inter6, gate53inter7, gate53inter8, gate53inter9, gate53inter10, gate53inter11, gate53inter12, gate42inter0, gate42inter1, gate42inter2, gate42inter3, gate42inter4, gate42inter5, gate42inter6, gate42inter7, gate42inter8, gate42inter9, gate42inter10, gate42inter11, gate42inter12, gate47inter0, gate47inter1, gate47inter2, gate47inter3, gate47inter4, gate47inter5, gate47inter6, gate47inter7, gate47inter8, gate47inter9, gate47inter10, gate47inter11, gate47inter12, gate65inter0, gate65inter1, gate65inter2, gate65inter3, gate65inter4, gate65inter5, gate65inter6, gate65inter7, gate65inter8, gate65inter9, gate65inter10, gate65inter11, gate65inter12, gate276inter0, gate276inter1, gate276inter2, gate276inter3, gate276inter4, gate276inter5, gate276inter6, gate276inter7, gate276inter8, gate276inter9, gate276inter10, gate276inter11, gate276inter12, gate469inter0, gate469inter1, gate469inter2, gate469inter3, gate469inter4, gate469inter5, gate469inter6, gate469inter7, gate469inter8, gate469inter9, gate469inter10, gate469inter11, gate469inter12, gate186inter0, gate186inter1, gate186inter2, gate186inter3, gate186inter4, gate186inter5, gate186inter6, gate186inter7, gate186inter8, gate186inter9, gate186inter10, gate186inter11, gate186inter12, gate9inter0, gate9inter1, gate9inter2, gate9inter3, gate9inter4, gate9inter5, gate9inter6, gate9inter7, gate9inter8, gate9inter9, gate9inter10, gate9inter11, gate9inter12, gate274inter0, gate274inter1, gate274inter2, gate274inter3, gate274inter4, gate274inter5, gate274inter6, gate274inter7, gate274inter8, gate274inter9, gate274inter10, gate274inter11, gate274inter12, gate61inter0, gate61inter1, gate61inter2, gate61inter3, gate61inter4, gate61inter5, gate61inter6, gate61inter7, gate61inter8, gate61inter9, gate61inter10, gate61inter11, gate61inter12, gate170inter0, gate170inter1, gate170inter2, gate170inter3, gate170inter4, gate170inter5, gate170inter6, gate170inter7, gate170inter8, gate170inter9, gate170inter10, gate170inter11, gate170inter12, gate36inter0, gate36inter1, gate36inter2, gate36inter3, gate36inter4, gate36inter5, gate36inter6, gate36inter7, gate36inter8, gate36inter9, gate36inter10, gate36inter11, gate36inter12, gate452inter0, gate452inter1, gate452inter2, gate452inter3, gate452inter4, gate452inter5, gate452inter6, gate452inter7, gate452inter8, gate452inter9, gate452inter10, gate452inter11, gate452inter12, gate23inter0, gate23inter1, gate23inter2, gate23inter3, gate23inter4, gate23inter5, gate23inter6, gate23inter7, gate23inter8, gate23inter9, gate23inter10, gate23inter11, gate23inter12, gate440inter0, gate440inter1, gate440inter2, gate440inter3, gate440inter4, gate440inter5, gate440inter6, gate440inter7, gate440inter8, gate440inter9, gate440inter10, gate440inter11, gate440inter12, gate12inter0, gate12inter1, gate12inter2, gate12inter3, gate12inter4, gate12inter5, gate12inter6, gate12inter7, gate12inter8, gate12inter9, gate12inter10, gate12inter11, gate12inter12, gate74inter0, gate74inter1, gate74inter2, gate74inter3, gate74inter4, gate74inter5, gate74inter6, gate74inter7, gate74inter8, gate74inter9, gate74inter10, gate74inter11, gate74inter12, gate475inter0, gate475inter1, gate475inter2, gate475inter3, gate475inter4, gate475inter5, gate475inter6, gate475inter7, gate475inter8, gate475inter9, gate475inter10, gate475inter11, gate475inter12, gate220inter0, gate220inter1, gate220inter2, gate220inter3, gate220inter4, gate220inter5, gate220inter6, gate220inter7, gate220inter8, gate220inter9, gate220inter10, gate220inter11, gate220inter12, gate474inter0, gate474inter1, gate474inter2, gate474inter3, gate474inter4, gate474inter5, gate474inter6, gate474inter7, gate474inter8, gate474inter9, gate474inter10, gate474inter11, gate474inter12, gate25inter0, gate25inter1, gate25inter2, gate25inter3, gate25inter4, gate25inter5, gate25inter6, gate25inter7, gate25inter8, gate25inter9, gate25inter10, gate25inter11, gate25inter12, gate425inter0, gate425inter1, gate425inter2, gate425inter3, gate425inter4, gate425inter5, gate425inter6, gate425inter7, gate425inter8, gate425inter9, gate425inter10, gate425inter11, gate425inter12, gate122inter0, gate122inter1, gate122inter2, gate122inter3, gate122inter4, gate122inter5, gate122inter6, gate122inter7, gate122inter8, gate122inter9, gate122inter10, gate122inter11, gate122inter12, gate39inter0, gate39inter1, gate39inter2, gate39inter3, gate39inter4, gate39inter5, gate39inter6, gate39inter7, gate39inter8, gate39inter9, gate39inter10, gate39inter11, gate39inter12, gate268inter0, gate268inter1, gate268inter2, gate268inter3, gate268inter4, gate268inter5, gate268inter6, gate268inter7, gate268inter8, gate268inter9, gate268inter10, gate268inter11, gate268inter12, gate109inter0, gate109inter1, gate109inter2, gate109inter3, gate109inter4, gate109inter5, gate109inter6, gate109inter7, gate109inter8, gate109inter9, gate109inter10, gate109inter11, gate109inter12, gate233inter0, gate233inter1, gate233inter2, gate233inter3, gate233inter4, gate233inter5, gate233inter6, gate233inter7, gate233inter8, gate233inter9, gate233inter10, gate233inter11, gate233inter12, gate204inter0, gate204inter1, gate204inter2, gate204inter3, gate204inter4, gate204inter5, gate204inter6, gate204inter7, gate204inter8, gate204inter9, gate204inter10, gate204inter11, gate204inter12, gate409inter0, gate409inter1, gate409inter2, gate409inter3, gate409inter4, gate409inter5, gate409inter6, gate409inter7, gate409inter8, gate409inter9, gate409inter10, gate409inter11, gate409inter12, gate51inter0, gate51inter1, gate51inter2, gate51inter3, gate51inter4, gate51inter5, gate51inter6, gate51inter7, gate51inter8, gate51inter9, gate51inter10, gate51inter11, gate51inter12, gate154inter0, gate154inter1, gate154inter2, gate154inter3, gate154inter4, gate154inter5, gate154inter6, gate154inter7, gate154inter8, gate154inter9, gate154inter10, gate154inter11, gate154inter12, gate102inter0, gate102inter1, gate102inter2, gate102inter3, gate102inter4, gate102inter5, gate102inter6, gate102inter7, gate102inter8, gate102inter9, gate102inter10, gate102inter11, gate102inter12, gate396inter0, gate396inter1, gate396inter2, gate396inter3, gate396inter4, gate396inter5, gate396inter6, gate396inter7, gate396inter8, gate396inter9, gate396inter10, gate396inter11, gate396inter12, gate244inter0, gate244inter1, gate244inter2, gate244inter3, gate244inter4, gate244inter5, gate244inter6, gate244inter7, gate244inter8, gate244inter9, gate244inter10, gate244inter11, gate244inter12, gate217inter0, gate217inter1, gate217inter2, gate217inter3, gate217inter4, gate217inter5, gate217inter6, gate217inter7, gate217inter8, gate217inter9, gate217inter10, gate217inter11, gate217inter12, gate148inter0, gate148inter1, gate148inter2, gate148inter3, gate148inter4, gate148inter5, gate148inter6, gate148inter7, gate148inter8, gate148inter9, gate148inter10, gate148inter11, gate148inter12, gate180inter0, gate180inter1, gate180inter2, gate180inter3, gate180inter4, gate180inter5, gate180inter6, gate180inter7, gate180inter8, gate180inter9, gate180inter10, gate180inter11, gate180inter12, gate406inter0, gate406inter1, gate406inter2, gate406inter3, gate406inter4, gate406inter5, gate406inter6, gate406inter7, gate406inter8, gate406inter9, gate406inter10, gate406inter11, gate406inter12, gate26inter0, gate26inter1, gate26inter2, gate26inter3, gate26inter4, gate26inter5, gate26inter6, gate26inter7, gate26inter8, gate26inter9, gate26inter10, gate26inter11, gate26inter12, gate138inter0, gate138inter1, gate138inter2, gate138inter3, gate138inter4, gate138inter5, gate138inter6, gate138inter7, gate138inter8, gate138inter9, gate138inter10, gate138inter11, gate138inter12, gate107inter0, gate107inter1, gate107inter2, gate107inter3, gate107inter4, gate107inter5, gate107inter6, gate107inter7, gate107inter8, gate107inter9, gate107inter10, gate107inter11, gate107inter12, gate428inter0, gate428inter1, gate428inter2, gate428inter3, gate428inter4, gate428inter5, gate428inter6, gate428inter7, gate428inter8, gate428inter9, gate428inter10, gate428inter11, gate428inter12, gate255inter0, gate255inter1, gate255inter2, gate255inter3, gate255inter4, gate255inter5, gate255inter6, gate255inter7, gate255inter8, gate255inter9, gate255inter10, gate255inter11, gate255inter12, gate106inter0, gate106inter1, gate106inter2, gate106inter3, gate106inter4, gate106inter5, gate106inter6, gate106inter7, gate106inter8, gate106inter9, gate106inter10, gate106inter11, gate106inter12, gate97inter0, gate97inter1, gate97inter2, gate97inter3, gate97inter4, gate97inter5, gate97inter6, gate97inter7, gate97inter8, gate97inter9, gate97inter10, gate97inter11, gate97inter12, gate450inter0, gate450inter1, gate450inter2, gate450inter3, gate450inter4, gate450inter5, gate450inter6, gate450inter7, gate450inter8, gate450inter9, gate450inter10, gate450inter11, gate450inter12, gate14inter0, gate14inter1, gate14inter2, gate14inter3, gate14inter4, gate14inter5, gate14inter6, gate14inter7, gate14inter8, gate14inter9, gate14inter10, gate14inter11, gate14inter12, gate80inter0, gate80inter1, gate80inter2, gate80inter3, gate80inter4, gate80inter5, gate80inter6, gate80inter7, gate80inter8, gate80inter9, gate80inter10, gate80inter11, gate80inter12, gate151inter0, gate151inter1, gate151inter2, gate151inter3, gate151inter4, gate151inter5, gate151inter6, gate151inter7, gate151inter8, gate151inter9, gate151inter10, gate151inter11, gate151inter12, gate451inter0, gate451inter1, gate451inter2, gate451inter3, gate451inter4, gate451inter5, gate451inter6, gate451inter7, gate451inter8, gate451inter9, gate451inter10, gate451inter11, gate451inter12, gate124inter0, gate124inter1, gate124inter2, gate124inter3, gate124inter4, gate124inter5, gate124inter6, gate124inter7, gate124inter8, gate124inter9, gate124inter10, gate124inter11, gate124inter12, gate286inter0, gate286inter1, gate286inter2, gate286inter3, gate286inter4, gate286inter5, gate286inter6, gate286inter7, gate286inter8, gate286inter9, gate286inter10, gate286inter11, gate286inter12, gate219inter0, gate219inter1, gate219inter2, gate219inter3, gate219inter4, gate219inter5, gate219inter6, gate219inter7, gate219inter8, gate219inter9, gate219inter10, gate219inter11, gate219inter12, gate283inter0, gate283inter1, gate283inter2, gate283inter3, gate283inter4, gate283inter5, gate283inter6, gate283inter7, gate283inter8, gate283inter9, gate283inter10, gate283inter11, gate283inter12, gate156inter0, gate156inter1, gate156inter2, gate156inter3, gate156inter4, gate156inter5, gate156inter6, gate156inter7, gate156inter8, gate156inter9, gate156inter10, gate156inter11, gate156inter12, gate230inter0, gate230inter1, gate230inter2, gate230inter3, gate230inter4, gate230inter5, gate230inter6, gate230inter7, gate230inter8, gate230inter9, gate230inter10, gate230inter11, gate230inter12, gate459inter0, gate459inter1, gate459inter2, gate459inter3, gate459inter4, gate459inter5, gate459inter6, gate459inter7, gate459inter8, gate459inter9, gate459inter10, gate459inter11, gate459inter12, gate429inter0, gate429inter1, gate429inter2, gate429inter3, gate429inter4, gate429inter5, gate429inter6, gate429inter7, gate429inter8, gate429inter9, gate429inter10, gate429inter11, gate429inter12, gate85inter0, gate85inter1, gate85inter2, gate85inter3, gate85inter4, gate85inter5, gate85inter6, gate85inter7, gate85inter8, gate85inter9, gate85inter10, gate85inter11, gate85inter12;



and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );

  xor2  gate1443(.a(G2), .b(G1), .O(gate9inter0));
  nand2 gate1444(.a(gate9inter0), .b(s_128), .O(gate9inter1));
  and2  gate1445(.a(G2), .b(G1), .O(gate9inter2));
  inv1  gate1446(.a(s_128), .O(gate9inter3));
  inv1  gate1447(.a(s_129), .O(gate9inter4));
  nand2 gate1448(.a(gate9inter4), .b(gate9inter3), .O(gate9inter5));
  nor2  gate1449(.a(gate9inter5), .b(gate9inter2), .O(gate9inter6));
  inv1  gate1450(.a(G1), .O(gate9inter7));
  inv1  gate1451(.a(G2), .O(gate9inter8));
  nand2 gate1452(.a(gate9inter8), .b(gate9inter7), .O(gate9inter9));
  nand2 gate1453(.a(s_129), .b(gate9inter3), .O(gate9inter10));
  nor2  gate1454(.a(gate9inter10), .b(gate9inter9), .O(gate9inter11));
  nor2  gate1455(.a(gate9inter11), .b(gate9inter6), .O(gate9inter12));
  nand2 gate1456(.a(gate9inter12), .b(gate9inter1), .O(G266));

  xor2  gate1205(.a(G4), .b(G3), .O(gate10inter0));
  nand2 gate1206(.a(gate10inter0), .b(s_94), .O(gate10inter1));
  and2  gate1207(.a(G4), .b(G3), .O(gate10inter2));
  inv1  gate1208(.a(s_94), .O(gate10inter3));
  inv1  gate1209(.a(s_95), .O(gate10inter4));
  nand2 gate1210(.a(gate10inter4), .b(gate10inter3), .O(gate10inter5));
  nor2  gate1211(.a(gate10inter5), .b(gate10inter2), .O(gate10inter6));
  inv1  gate1212(.a(G3), .O(gate10inter7));
  inv1  gate1213(.a(G4), .O(gate10inter8));
  nand2 gate1214(.a(gate10inter8), .b(gate10inter7), .O(gate10inter9));
  nand2 gate1215(.a(s_95), .b(gate10inter3), .O(gate10inter10));
  nor2  gate1216(.a(gate10inter10), .b(gate10inter9), .O(gate10inter11));
  nor2  gate1217(.a(gate10inter11), .b(gate10inter6), .O(gate10inter12));
  nand2 gate1218(.a(gate10inter12), .b(gate10inter1), .O(G269));
nand2 gate11( .a(G5), .b(G6), .O(G272) );

  xor2  gate1555(.a(G8), .b(G7), .O(gate12inter0));
  nand2 gate1556(.a(gate12inter0), .b(s_144), .O(gate12inter1));
  and2  gate1557(.a(G8), .b(G7), .O(gate12inter2));
  inv1  gate1558(.a(s_144), .O(gate12inter3));
  inv1  gate1559(.a(s_145), .O(gate12inter4));
  nand2 gate1560(.a(gate12inter4), .b(gate12inter3), .O(gate12inter5));
  nor2  gate1561(.a(gate12inter5), .b(gate12inter2), .O(gate12inter6));
  inv1  gate1562(.a(G7), .O(gate12inter7));
  inv1  gate1563(.a(G8), .O(gate12inter8));
  nand2 gate1564(.a(gate12inter8), .b(gate12inter7), .O(gate12inter9));
  nand2 gate1565(.a(s_145), .b(gate12inter3), .O(gate12inter10));
  nor2  gate1566(.a(gate12inter10), .b(gate12inter9), .O(gate12inter11));
  nor2  gate1567(.a(gate12inter11), .b(gate12inter6), .O(gate12inter12));
  nand2 gate1568(.a(gate12inter12), .b(gate12inter1), .O(G275));
nand2 gate13( .a(G9), .b(G10), .O(G278) );

  xor2  gate1989(.a(G12), .b(G11), .O(gate14inter0));
  nand2 gate1990(.a(gate14inter0), .b(s_206), .O(gate14inter1));
  and2  gate1991(.a(G12), .b(G11), .O(gate14inter2));
  inv1  gate1992(.a(s_206), .O(gate14inter3));
  inv1  gate1993(.a(s_207), .O(gate14inter4));
  nand2 gate1994(.a(gate14inter4), .b(gate14inter3), .O(gate14inter5));
  nor2  gate1995(.a(gate14inter5), .b(gate14inter2), .O(gate14inter6));
  inv1  gate1996(.a(G11), .O(gate14inter7));
  inv1  gate1997(.a(G12), .O(gate14inter8));
  nand2 gate1998(.a(gate14inter8), .b(gate14inter7), .O(gate14inter9));
  nand2 gate1999(.a(s_207), .b(gate14inter3), .O(gate14inter10));
  nor2  gate2000(.a(gate14inter10), .b(gate14inter9), .O(gate14inter11));
  nor2  gate2001(.a(gate14inter11), .b(gate14inter6), .O(gate14inter12));
  nand2 gate2002(.a(gate14inter12), .b(gate14inter1), .O(G281));
nand2 gate15( .a(G13), .b(G14), .O(G284) );
nand2 gate16( .a(G15), .b(G16), .O(G287) );
nand2 gate17( .a(G17), .b(G18), .O(G290) );
nand2 gate18( .a(G19), .b(G20), .O(G293) );
nand2 gate19( .a(G21), .b(G22), .O(G296) );
nand2 gate20( .a(G23), .b(G24), .O(G299) );
nand2 gate21( .a(G25), .b(G26), .O(G302) );
nand2 gate22( .a(G27), .b(G28), .O(G305) );

  xor2  gate1527(.a(G30), .b(G29), .O(gate23inter0));
  nand2 gate1528(.a(gate23inter0), .b(s_140), .O(gate23inter1));
  and2  gate1529(.a(G30), .b(G29), .O(gate23inter2));
  inv1  gate1530(.a(s_140), .O(gate23inter3));
  inv1  gate1531(.a(s_141), .O(gate23inter4));
  nand2 gate1532(.a(gate23inter4), .b(gate23inter3), .O(gate23inter5));
  nor2  gate1533(.a(gate23inter5), .b(gate23inter2), .O(gate23inter6));
  inv1  gate1534(.a(G29), .O(gate23inter7));
  inv1  gate1535(.a(G30), .O(gate23inter8));
  nand2 gate1536(.a(gate23inter8), .b(gate23inter7), .O(gate23inter9));
  nand2 gate1537(.a(s_141), .b(gate23inter3), .O(gate23inter10));
  nor2  gate1538(.a(gate23inter10), .b(gate23inter9), .O(gate23inter11));
  nor2  gate1539(.a(gate23inter11), .b(gate23inter6), .O(gate23inter12));
  nand2 gate1540(.a(gate23inter12), .b(gate23inter1), .O(G308));

  xor2  gate1261(.a(G32), .b(G31), .O(gate24inter0));
  nand2 gate1262(.a(gate24inter0), .b(s_102), .O(gate24inter1));
  and2  gate1263(.a(G32), .b(G31), .O(gate24inter2));
  inv1  gate1264(.a(s_102), .O(gate24inter3));
  inv1  gate1265(.a(s_103), .O(gate24inter4));
  nand2 gate1266(.a(gate24inter4), .b(gate24inter3), .O(gate24inter5));
  nor2  gate1267(.a(gate24inter5), .b(gate24inter2), .O(gate24inter6));
  inv1  gate1268(.a(G31), .O(gate24inter7));
  inv1  gate1269(.a(G32), .O(gate24inter8));
  nand2 gate1270(.a(gate24inter8), .b(gate24inter7), .O(gate24inter9));
  nand2 gate1271(.a(s_103), .b(gate24inter3), .O(gate24inter10));
  nor2  gate1272(.a(gate24inter10), .b(gate24inter9), .O(gate24inter11));
  nor2  gate1273(.a(gate24inter11), .b(gate24inter6), .O(gate24inter12));
  nand2 gate1274(.a(gate24inter12), .b(gate24inter1), .O(G311));

  xor2  gate1625(.a(G5), .b(G1), .O(gate25inter0));
  nand2 gate1626(.a(gate25inter0), .b(s_154), .O(gate25inter1));
  and2  gate1627(.a(G5), .b(G1), .O(gate25inter2));
  inv1  gate1628(.a(s_154), .O(gate25inter3));
  inv1  gate1629(.a(s_155), .O(gate25inter4));
  nand2 gate1630(.a(gate25inter4), .b(gate25inter3), .O(gate25inter5));
  nor2  gate1631(.a(gate25inter5), .b(gate25inter2), .O(gate25inter6));
  inv1  gate1632(.a(G1), .O(gate25inter7));
  inv1  gate1633(.a(G5), .O(gate25inter8));
  nand2 gate1634(.a(gate25inter8), .b(gate25inter7), .O(gate25inter9));
  nand2 gate1635(.a(s_155), .b(gate25inter3), .O(gate25inter10));
  nor2  gate1636(.a(gate25inter10), .b(gate25inter9), .O(gate25inter11));
  nor2  gate1637(.a(gate25inter11), .b(gate25inter6), .O(gate25inter12));
  nand2 gate1638(.a(gate25inter12), .b(gate25inter1), .O(G314));

  xor2  gate1877(.a(G13), .b(G9), .O(gate26inter0));
  nand2 gate1878(.a(gate26inter0), .b(s_190), .O(gate26inter1));
  and2  gate1879(.a(G13), .b(G9), .O(gate26inter2));
  inv1  gate1880(.a(s_190), .O(gate26inter3));
  inv1  gate1881(.a(s_191), .O(gate26inter4));
  nand2 gate1882(.a(gate26inter4), .b(gate26inter3), .O(gate26inter5));
  nor2  gate1883(.a(gate26inter5), .b(gate26inter2), .O(gate26inter6));
  inv1  gate1884(.a(G9), .O(gate26inter7));
  inv1  gate1885(.a(G13), .O(gate26inter8));
  nand2 gate1886(.a(gate26inter8), .b(gate26inter7), .O(gate26inter9));
  nand2 gate1887(.a(s_191), .b(gate26inter3), .O(gate26inter10));
  nor2  gate1888(.a(gate26inter10), .b(gate26inter9), .O(gate26inter11));
  nor2  gate1889(.a(gate26inter11), .b(gate26inter6), .O(gate26inter12));
  nand2 gate1890(.a(gate26inter12), .b(gate26inter1), .O(G317));
nand2 gate27( .a(G2), .b(G6), .O(G320) );
nand2 gate28( .a(G10), .b(G14), .O(G323) );
nand2 gate29( .a(G3), .b(G7), .O(G326) );
nand2 gate30( .a(G11), .b(G15), .O(G329) );
nand2 gate31( .a(G4), .b(G8), .O(G332) );
nand2 gate32( .a(G12), .b(G16), .O(G335) );
nand2 gate33( .a(G17), .b(G21), .O(G338) );
nand2 gate34( .a(G25), .b(G29), .O(G341) );
nand2 gate35( .a(G18), .b(G22), .O(G344) );

  xor2  gate1499(.a(G30), .b(G26), .O(gate36inter0));
  nand2 gate1500(.a(gate36inter0), .b(s_136), .O(gate36inter1));
  and2  gate1501(.a(G30), .b(G26), .O(gate36inter2));
  inv1  gate1502(.a(s_136), .O(gate36inter3));
  inv1  gate1503(.a(s_137), .O(gate36inter4));
  nand2 gate1504(.a(gate36inter4), .b(gate36inter3), .O(gate36inter5));
  nor2  gate1505(.a(gate36inter5), .b(gate36inter2), .O(gate36inter6));
  inv1  gate1506(.a(G26), .O(gate36inter7));
  inv1  gate1507(.a(G30), .O(gate36inter8));
  nand2 gate1508(.a(gate36inter8), .b(gate36inter7), .O(gate36inter9));
  nand2 gate1509(.a(s_137), .b(gate36inter3), .O(gate36inter10));
  nor2  gate1510(.a(gate36inter10), .b(gate36inter9), .O(gate36inter11));
  nor2  gate1511(.a(gate36inter11), .b(gate36inter6), .O(gate36inter12));
  nand2 gate1512(.a(gate36inter12), .b(gate36inter1), .O(G347));

  xor2  gate1135(.a(G23), .b(G19), .O(gate37inter0));
  nand2 gate1136(.a(gate37inter0), .b(s_84), .O(gate37inter1));
  and2  gate1137(.a(G23), .b(G19), .O(gate37inter2));
  inv1  gate1138(.a(s_84), .O(gate37inter3));
  inv1  gate1139(.a(s_85), .O(gate37inter4));
  nand2 gate1140(.a(gate37inter4), .b(gate37inter3), .O(gate37inter5));
  nor2  gate1141(.a(gate37inter5), .b(gate37inter2), .O(gate37inter6));
  inv1  gate1142(.a(G19), .O(gate37inter7));
  inv1  gate1143(.a(G23), .O(gate37inter8));
  nand2 gate1144(.a(gate37inter8), .b(gate37inter7), .O(gate37inter9));
  nand2 gate1145(.a(s_85), .b(gate37inter3), .O(gate37inter10));
  nor2  gate1146(.a(gate37inter10), .b(gate37inter9), .O(gate37inter11));
  nor2  gate1147(.a(gate37inter11), .b(gate37inter6), .O(gate37inter12));
  nand2 gate1148(.a(gate37inter12), .b(gate37inter1), .O(G350));
nand2 gate38( .a(G27), .b(G31), .O(G353) );

  xor2  gate1667(.a(G24), .b(G20), .O(gate39inter0));
  nand2 gate1668(.a(gate39inter0), .b(s_160), .O(gate39inter1));
  and2  gate1669(.a(G24), .b(G20), .O(gate39inter2));
  inv1  gate1670(.a(s_160), .O(gate39inter3));
  inv1  gate1671(.a(s_161), .O(gate39inter4));
  nand2 gate1672(.a(gate39inter4), .b(gate39inter3), .O(gate39inter5));
  nor2  gate1673(.a(gate39inter5), .b(gate39inter2), .O(gate39inter6));
  inv1  gate1674(.a(G20), .O(gate39inter7));
  inv1  gate1675(.a(G24), .O(gate39inter8));
  nand2 gate1676(.a(gate39inter8), .b(gate39inter7), .O(gate39inter9));
  nand2 gate1677(.a(s_161), .b(gate39inter3), .O(gate39inter10));
  nor2  gate1678(.a(gate39inter10), .b(gate39inter9), .O(gate39inter11));
  nor2  gate1679(.a(gate39inter11), .b(gate39inter6), .O(gate39inter12));
  nand2 gate1680(.a(gate39inter12), .b(gate39inter1), .O(G356));
nand2 gate40( .a(G28), .b(G32), .O(G359) );

  xor2  gate841(.a(G266), .b(G1), .O(gate41inter0));
  nand2 gate842(.a(gate41inter0), .b(s_42), .O(gate41inter1));
  and2  gate843(.a(G266), .b(G1), .O(gate41inter2));
  inv1  gate844(.a(s_42), .O(gate41inter3));
  inv1  gate845(.a(s_43), .O(gate41inter4));
  nand2 gate846(.a(gate41inter4), .b(gate41inter3), .O(gate41inter5));
  nor2  gate847(.a(gate41inter5), .b(gate41inter2), .O(gate41inter6));
  inv1  gate848(.a(G1), .O(gate41inter7));
  inv1  gate849(.a(G266), .O(gate41inter8));
  nand2 gate850(.a(gate41inter8), .b(gate41inter7), .O(gate41inter9));
  nand2 gate851(.a(s_43), .b(gate41inter3), .O(gate41inter10));
  nor2  gate852(.a(gate41inter10), .b(gate41inter9), .O(gate41inter11));
  nor2  gate853(.a(gate41inter11), .b(gate41inter6), .O(gate41inter12));
  nand2 gate854(.a(gate41inter12), .b(gate41inter1), .O(G362));

  xor2  gate1359(.a(G266), .b(G2), .O(gate42inter0));
  nand2 gate1360(.a(gate42inter0), .b(s_116), .O(gate42inter1));
  and2  gate1361(.a(G266), .b(G2), .O(gate42inter2));
  inv1  gate1362(.a(s_116), .O(gate42inter3));
  inv1  gate1363(.a(s_117), .O(gate42inter4));
  nand2 gate1364(.a(gate42inter4), .b(gate42inter3), .O(gate42inter5));
  nor2  gate1365(.a(gate42inter5), .b(gate42inter2), .O(gate42inter6));
  inv1  gate1366(.a(G2), .O(gate42inter7));
  inv1  gate1367(.a(G266), .O(gate42inter8));
  nand2 gate1368(.a(gate42inter8), .b(gate42inter7), .O(gate42inter9));
  nand2 gate1369(.a(s_117), .b(gate42inter3), .O(gate42inter10));
  nor2  gate1370(.a(gate42inter10), .b(gate42inter9), .O(gate42inter11));
  nor2  gate1371(.a(gate42inter11), .b(gate42inter6), .O(gate42inter12));
  nand2 gate1372(.a(gate42inter12), .b(gate42inter1), .O(G363));
nand2 gate43( .a(G3), .b(G269), .O(G364) );
nand2 gate44( .a(G4), .b(G269), .O(G365) );
nand2 gate45( .a(G5), .b(G272), .O(G366) );
nand2 gate46( .a(G6), .b(G272), .O(G367) );

  xor2  gate1373(.a(G275), .b(G7), .O(gate47inter0));
  nand2 gate1374(.a(gate47inter0), .b(s_118), .O(gate47inter1));
  and2  gate1375(.a(G275), .b(G7), .O(gate47inter2));
  inv1  gate1376(.a(s_118), .O(gate47inter3));
  inv1  gate1377(.a(s_119), .O(gate47inter4));
  nand2 gate1378(.a(gate47inter4), .b(gate47inter3), .O(gate47inter5));
  nor2  gate1379(.a(gate47inter5), .b(gate47inter2), .O(gate47inter6));
  inv1  gate1380(.a(G7), .O(gate47inter7));
  inv1  gate1381(.a(G275), .O(gate47inter8));
  nand2 gate1382(.a(gate47inter8), .b(gate47inter7), .O(gate47inter9));
  nand2 gate1383(.a(s_119), .b(gate47inter3), .O(gate47inter10));
  nor2  gate1384(.a(gate47inter10), .b(gate47inter9), .O(gate47inter11));
  nor2  gate1385(.a(gate47inter11), .b(gate47inter6), .O(gate47inter12));
  nand2 gate1386(.a(gate47inter12), .b(gate47inter1), .O(G368));
nand2 gate48( .a(G8), .b(G275), .O(G369) );
nand2 gate49( .a(G9), .b(G278), .O(G370) );
nand2 gate50( .a(G10), .b(G278), .O(G371) );

  xor2  gate1751(.a(G281), .b(G11), .O(gate51inter0));
  nand2 gate1752(.a(gate51inter0), .b(s_172), .O(gate51inter1));
  and2  gate1753(.a(G281), .b(G11), .O(gate51inter2));
  inv1  gate1754(.a(s_172), .O(gate51inter3));
  inv1  gate1755(.a(s_173), .O(gate51inter4));
  nand2 gate1756(.a(gate51inter4), .b(gate51inter3), .O(gate51inter5));
  nor2  gate1757(.a(gate51inter5), .b(gate51inter2), .O(gate51inter6));
  inv1  gate1758(.a(G11), .O(gate51inter7));
  inv1  gate1759(.a(G281), .O(gate51inter8));
  nand2 gate1760(.a(gate51inter8), .b(gate51inter7), .O(gate51inter9));
  nand2 gate1761(.a(s_173), .b(gate51inter3), .O(gate51inter10));
  nor2  gate1762(.a(gate51inter10), .b(gate51inter9), .O(gate51inter11));
  nor2  gate1763(.a(gate51inter11), .b(gate51inter6), .O(gate51inter12));
  nand2 gate1764(.a(gate51inter12), .b(gate51inter1), .O(G372));
nand2 gate52( .a(G12), .b(G281), .O(G373) );

  xor2  gate1345(.a(G284), .b(G13), .O(gate53inter0));
  nand2 gate1346(.a(gate53inter0), .b(s_114), .O(gate53inter1));
  and2  gate1347(.a(G284), .b(G13), .O(gate53inter2));
  inv1  gate1348(.a(s_114), .O(gate53inter3));
  inv1  gate1349(.a(s_115), .O(gate53inter4));
  nand2 gate1350(.a(gate53inter4), .b(gate53inter3), .O(gate53inter5));
  nor2  gate1351(.a(gate53inter5), .b(gate53inter2), .O(gate53inter6));
  inv1  gate1352(.a(G13), .O(gate53inter7));
  inv1  gate1353(.a(G284), .O(gate53inter8));
  nand2 gate1354(.a(gate53inter8), .b(gate53inter7), .O(gate53inter9));
  nand2 gate1355(.a(s_115), .b(gate53inter3), .O(gate53inter10));
  nor2  gate1356(.a(gate53inter10), .b(gate53inter9), .O(gate53inter11));
  nor2  gate1357(.a(gate53inter11), .b(gate53inter6), .O(gate53inter12));
  nand2 gate1358(.a(gate53inter12), .b(gate53inter1), .O(G374));
nand2 gate54( .a(G14), .b(G284), .O(G375) );
nand2 gate55( .a(G15), .b(G287), .O(G376) );
nand2 gate56( .a(G16), .b(G287), .O(G377) );
nand2 gate57( .a(G17), .b(G290), .O(G378) );
nand2 gate58( .a(G18), .b(G290), .O(G379) );

  xor2  gate1233(.a(G293), .b(G19), .O(gate59inter0));
  nand2 gate1234(.a(gate59inter0), .b(s_98), .O(gate59inter1));
  and2  gate1235(.a(G293), .b(G19), .O(gate59inter2));
  inv1  gate1236(.a(s_98), .O(gate59inter3));
  inv1  gate1237(.a(s_99), .O(gate59inter4));
  nand2 gate1238(.a(gate59inter4), .b(gate59inter3), .O(gate59inter5));
  nor2  gate1239(.a(gate59inter5), .b(gate59inter2), .O(gate59inter6));
  inv1  gate1240(.a(G19), .O(gate59inter7));
  inv1  gate1241(.a(G293), .O(gate59inter8));
  nand2 gate1242(.a(gate59inter8), .b(gate59inter7), .O(gate59inter9));
  nand2 gate1243(.a(s_99), .b(gate59inter3), .O(gate59inter10));
  nor2  gate1244(.a(gate59inter10), .b(gate59inter9), .O(gate59inter11));
  nor2  gate1245(.a(gate59inter11), .b(gate59inter6), .O(gate59inter12));
  nand2 gate1246(.a(gate59inter12), .b(gate59inter1), .O(G380));
nand2 gate60( .a(G20), .b(G293), .O(G381) );

  xor2  gate1471(.a(G296), .b(G21), .O(gate61inter0));
  nand2 gate1472(.a(gate61inter0), .b(s_132), .O(gate61inter1));
  and2  gate1473(.a(G296), .b(G21), .O(gate61inter2));
  inv1  gate1474(.a(s_132), .O(gate61inter3));
  inv1  gate1475(.a(s_133), .O(gate61inter4));
  nand2 gate1476(.a(gate61inter4), .b(gate61inter3), .O(gate61inter5));
  nor2  gate1477(.a(gate61inter5), .b(gate61inter2), .O(gate61inter6));
  inv1  gate1478(.a(G21), .O(gate61inter7));
  inv1  gate1479(.a(G296), .O(gate61inter8));
  nand2 gate1480(.a(gate61inter8), .b(gate61inter7), .O(gate61inter9));
  nand2 gate1481(.a(s_133), .b(gate61inter3), .O(gate61inter10));
  nor2  gate1482(.a(gate61inter10), .b(gate61inter9), .O(gate61inter11));
  nor2  gate1483(.a(gate61inter11), .b(gate61inter6), .O(gate61inter12));
  nand2 gate1484(.a(gate61inter12), .b(gate61inter1), .O(G382));
nand2 gate62( .a(G22), .b(G296), .O(G383) );
nand2 gate63( .a(G23), .b(G299), .O(G384) );

  xor2  gate799(.a(G299), .b(G24), .O(gate64inter0));
  nand2 gate800(.a(gate64inter0), .b(s_36), .O(gate64inter1));
  and2  gate801(.a(G299), .b(G24), .O(gate64inter2));
  inv1  gate802(.a(s_36), .O(gate64inter3));
  inv1  gate803(.a(s_37), .O(gate64inter4));
  nand2 gate804(.a(gate64inter4), .b(gate64inter3), .O(gate64inter5));
  nor2  gate805(.a(gate64inter5), .b(gate64inter2), .O(gate64inter6));
  inv1  gate806(.a(G24), .O(gate64inter7));
  inv1  gate807(.a(G299), .O(gate64inter8));
  nand2 gate808(.a(gate64inter8), .b(gate64inter7), .O(gate64inter9));
  nand2 gate809(.a(s_37), .b(gate64inter3), .O(gate64inter10));
  nor2  gate810(.a(gate64inter10), .b(gate64inter9), .O(gate64inter11));
  nor2  gate811(.a(gate64inter11), .b(gate64inter6), .O(gate64inter12));
  nand2 gate812(.a(gate64inter12), .b(gate64inter1), .O(G385));

  xor2  gate1387(.a(G302), .b(G25), .O(gate65inter0));
  nand2 gate1388(.a(gate65inter0), .b(s_120), .O(gate65inter1));
  and2  gate1389(.a(G302), .b(G25), .O(gate65inter2));
  inv1  gate1390(.a(s_120), .O(gate65inter3));
  inv1  gate1391(.a(s_121), .O(gate65inter4));
  nand2 gate1392(.a(gate65inter4), .b(gate65inter3), .O(gate65inter5));
  nor2  gate1393(.a(gate65inter5), .b(gate65inter2), .O(gate65inter6));
  inv1  gate1394(.a(G25), .O(gate65inter7));
  inv1  gate1395(.a(G302), .O(gate65inter8));
  nand2 gate1396(.a(gate65inter8), .b(gate65inter7), .O(gate65inter9));
  nand2 gate1397(.a(s_121), .b(gate65inter3), .O(gate65inter10));
  nor2  gate1398(.a(gate65inter10), .b(gate65inter9), .O(gate65inter11));
  nor2  gate1399(.a(gate65inter11), .b(gate65inter6), .O(gate65inter12));
  nand2 gate1400(.a(gate65inter12), .b(gate65inter1), .O(G386));
nand2 gate66( .a(G26), .b(G302), .O(G387) );
nand2 gate67( .a(G27), .b(G305), .O(G388) );
nand2 gate68( .a(G28), .b(G305), .O(G389) );
nand2 gate69( .a(G29), .b(G308), .O(G390) );
nand2 gate70( .a(G30), .b(G308), .O(G391) );
nand2 gate71( .a(G31), .b(G311), .O(G392) );

  xor2  gate1191(.a(G311), .b(G32), .O(gate72inter0));
  nand2 gate1192(.a(gate72inter0), .b(s_92), .O(gate72inter1));
  and2  gate1193(.a(G311), .b(G32), .O(gate72inter2));
  inv1  gate1194(.a(s_92), .O(gate72inter3));
  inv1  gate1195(.a(s_93), .O(gate72inter4));
  nand2 gate1196(.a(gate72inter4), .b(gate72inter3), .O(gate72inter5));
  nor2  gate1197(.a(gate72inter5), .b(gate72inter2), .O(gate72inter6));
  inv1  gate1198(.a(G32), .O(gate72inter7));
  inv1  gate1199(.a(G311), .O(gate72inter8));
  nand2 gate1200(.a(gate72inter8), .b(gate72inter7), .O(gate72inter9));
  nand2 gate1201(.a(s_93), .b(gate72inter3), .O(gate72inter10));
  nor2  gate1202(.a(gate72inter10), .b(gate72inter9), .O(gate72inter11));
  nor2  gate1203(.a(gate72inter11), .b(gate72inter6), .O(gate72inter12));
  nand2 gate1204(.a(gate72inter12), .b(gate72inter1), .O(G393));
nand2 gate73( .a(G1), .b(G314), .O(G394) );

  xor2  gate1569(.a(G314), .b(G5), .O(gate74inter0));
  nand2 gate1570(.a(gate74inter0), .b(s_146), .O(gate74inter1));
  and2  gate1571(.a(G314), .b(G5), .O(gate74inter2));
  inv1  gate1572(.a(s_146), .O(gate74inter3));
  inv1  gate1573(.a(s_147), .O(gate74inter4));
  nand2 gate1574(.a(gate74inter4), .b(gate74inter3), .O(gate74inter5));
  nor2  gate1575(.a(gate74inter5), .b(gate74inter2), .O(gate74inter6));
  inv1  gate1576(.a(G5), .O(gate74inter7));
  inv1  gate1577(.a(G314), .O(gate74inter8));
  nand2 gate1578(.a(gate74inter8), .b(gate74inter7), .O(gate74inter9));
  nand2 gate1579(.a(s_147), .b(gate74inter3), .O(gate74inter10));
  nor2  gate1580(.a(gate74inter10), .b(gate74inter9), .O(gate74inter11));
  nor2  gate1581(.a(gate74inter11), .b(gate74inter6), .O(gate74inter12));
  nand2 gate1582(.a(gate74inter12), .b(gate74inter1), .O(G395));
nand2 gate75( .a(G9), .b(G317), .O(G396) );
nand2 gate76( .a(G13), .b(G317), .O(G397) );
nand2 gate77( .a(G2), .b(G320), .O(G398) );
nand2 gate78( .a(G6), .b(G320), .O(G399) );
nand2 gate79( .a(G10), .b(G323), .O(G400) );

  xor2  gate2003(.a(G323), .b(G14), .O(gate80inter0));
  nand2 gate2004(.a(gate80inter0), .b(s_208), .O(gate80inter1));
  and2  gate2005(.a(G323), .b(G14), .O(gate80inter2));
  inv1  gate2006(.a(s_208), .O(gate80inter3));
  inv1  gate2007(.a(s_209), .O(gate80inter4));
  nand2 gate2008(.a(gate80inter4), .b(gate80inter3), .O(gate80inter5));
  nor2  gate2009(.a(gate80inter5), .b(gate80inter2), .O(gate80inter6));
  inv1  gate2010(.a(G14), .O(gate80inter7));
  inv1  gate2011(.a(G323), .O(gate80inter8));
  nand2 gate2012(.a(gate80inter8), .b(gate80inter7), .O(gate80inter9));
  nand2 gate2013(.a(s_209), .b(gate80inter3), .O(gate80inter10));
  nor2  gate2014(.a(gate80inter10), .b(gate80inter9), .O(gate80inter11));
  nor2  gate2015(.a(gate80inter11), .b(gate80inter6), .O(gate80inter12));
  nand2 gate2016(.a(gate80inter12), .b(gate80inter1), .O(G401));
nand2 gate81( .a(G3), .b(G326), .O(G402) );
nand2 gate82( .a(G7), .b(G326), .O(G403) );
nand2 gate83( .a(G11), .b(G329), .O(G404) );
nand2 gate84( .a(G15), .b(G329), .O(G405) );

  xor2  gate2157(.a(G332), .b(G4), .O(gate85inter0));
  nand2 gate2158(.a(gate85inter0), .b(s_230), .O(gate85inter1));
  and2  gate2159(.a(G332), .b(G4), .O(gate85inter2));
  inv1  gate2160(.a(s_230), .O(gate85inter3));
  inv1  gate2161(.a(s_231), .O(gate85inter4));
  nand2 gate2162(.a(gate85inter4), .b(gate85inter3), .O(gate85inter5));
  nor2  gate2163(.a(gate85inter5), .b(gate85inter2), .O(gate85inter6));
  inv1  gate2164(.a(G4), .O(gate85inter7));
  inv1  gate2165(.a(G332), .O(gate85inter8));
  nand2 gate2166(.a(gate85inter8), .b(gate85inter7), .O(gate85inter9));
  nand2 gate2167(.a(s_231), .b(gate85inter3), .O(gate85inter10));
  nor2  gate2168(.a(gate85inter10), .b(gate85inter9), .O(gate85inter11));
  nor2  gate2169(.a(gate85inter11), .b(gate85inter6), .O(gate85inter12));
  nand2 gate2170(.a(gate85inter12), .b(gate85inter1), .O(G406));

  xor2  gate547(.a(G332), .b(G8), .O(gate86inter0));
  nand2 gate548(.a(gate86inter0), .b(s_0), .O(gate86inter1));
  and2  gate549(.a(G332), .b(G8), .O(gate86inter2));
  inv1  gate550(.a(s_0), .O(gate86inter3));
  inv1  gate551(.a(s_1), .O(gate86inter4));
  nand2 gate552(.a(gate86inter4), .b(gate86inter3), .O(gate86inter5));
  nor2  gate553(.a(gate86inter5), .b(gate86inter2), .O(gate86inter6));
  inv1  gate554(.a(G8), .O(gate86inter7));
  inv1  gate555(.a(G332), .O(gate86inter8));
  nand2 gate556(.a(gate86inter8), .b(gate86inter7), .O(gate86inter9));
  nand2 gate557(.a(s_1), .b(gate86inter3), .O(gate86inter10));
  nor2  gate558(.a(gate86inter10), .b(gate86inter9), .O(gate86inter11));
  nor2  gate559(.a(gate86inter11), .b(gate86inter6), .O(gate86inter12));
  nand2 gate560(.a(gate86inter12), .b(gate86inter1), .O(G407));
nand2 gate87( .a(G12), .b(G335), .O(G408) );
nand2 gate88( .a(G16), .b(G335), .O(G409) );
nand2 gate89( .a(G17), .b(G338), .O(G410) );
nand2 gate90( .a(G21), .b(G338), .O(G411) );
nand2 gate91( .a(G25), .b(G341), .O(G412) );
nand2 gate92( .a(G29), .b(G341), .O(G413) );
nand2 gate93( .a(G18), .b(G344), .O(G414) );
nand2 gate94( .a(G22), .b(G344), .O(G415) );
nand2 gate95( .a(G26), .b(G347), .O(G416) );
nand2 gate96( .a(G30), .b(G347), .O(G417) );

  xor2  gate1961(.a(G350), .b(G19), .O(gate97inter0));
  nand2 gate1962(.a(gate97inter0), .b(s_202), .O(gate97inter1));
  and2  gate1963(.a(G350), .b(G19), .O(gate97inter2));
  inv1  gate1964(.a(s_202), .O(gate97inter3));
  inv1  gate1965(.a(s_203), .O(gate97inter4));
  nand2 gate1966(.a(gate97inter4), .b(gate97inter3), .O(gate97inter5));
  nor2  gate1967(.a(gate97inter5), .b(gate97inter2), .O(gate97inter6));
  inv1  gate1968(.a(G19), .O(gate97inter7));
  inv1  gate1969(.a(G350), .O(gate97inter8));
  nand2 gate1970(.a(gate97inter8), .b(gate97inter7), .O(gate97inter9));
  nand2 gate1971(.a(s_203), .b(gate97inter3), .O(gate97inter10));
  nor2  gate1972(.a(gate97inter10), .b(gate97inter9), .O(gate97inter11));
  nor2  gate1973(.a(gate97inter11), .b(gate97inter6), .O(gate97inter12));
  nand2 gate1974(.a(gate97inter12), .b(gate97inter1), .O(G418));
nand2 gate98( .a(G23), .b(G350), .O(G419) );

  xor2  gate743(.a(G353), .b(G27), .O(gate99inter0));
  nand2 gate744(.a(gate99inter0), .b(s_28), .O(gate99inter1));
  and2  gate745(.a(G353), .b(G27), .O(gate99inter2));
  inv1  gate746(.a(s_28), .O(gate99inter3));
  inv1  gate747(.a(s_29), .O(gate99inter4));
  nand2 gate748(.a(gate99inter4), .b(gate99inter3), .O(gate99inter5));
  nor2  gate749(.a(gate99inter5), .b(gate99inter2), .O(gate99inter6));
  inv1  gate750(.a(G27), .O(gate99inter7));
  inv1  gate751(.a(G353), .O(gate99inter8));
  nand2 gate752(.a(gate99inter8), .b(gate99inter7), .O(gate99inter9));
  nand2 gate753(.a(s_29), .b(gate99inter3), .O(gate99inter10));
  nor2  gate754(.a(gate99inter10), .b(gate99inter9), .O(gate99inter11));
  nor2  gate755(.a(gate99inter11), .b(gate99inter6), .O(gate99inter12));
  nand2 gate756(.a(gate99inter12), .b(gate99inter1), .O(G420));
nand2 gate100( .a(G31), .b(G353), .O(G421) );
nand2 gate101( .a(G20), .b(G356), .O(G422) );

  xor2  gate1779(.a(G356), .b(G24), .O(gate102inter0));
  nand2 gate1780(.a(gate102inter0), .b(s_176), .O(gate102inter1));
  and2  gate1781(.a(G356), .b(G24), .O(gate102inter2));
  inv1  gate1782(.a(s_176), .O(gate102inter3));
  inv1  gate1783(.a(s_177), .O(gate102inter4));
  nand2 gate1784(.a(gate102inter4), .b(gate102inter3), .O(gate102inter5));
  nor2  gate1785(.a(gate102inter5), .b(gate102inter2), .O(gate102inter6));
  inv1  gate1786(.a(G24), .O(gate102inter7));
  inv1  gate1787(.a(G356), .O(gate102inter8));
  nand2 gate1788(.a(gate102inter8), .b(gate102inter7), .O(gate102inter9));
  nand2 gate1789(.a(s_177), .b(gate102inter3), .O(gate102inter10));
  nor2  gate1790(.a(gate102inter10), .b(gate102inter9), .O(gate102inter11));
  nor2  gate1791(.a(gate102inter11), .b(gate102inter6), .O(gate102inter12));
  nand2 gate1792(.a(gate102inter12), .b(gate102inter1), .O(G423));
nand2 gate103( .a(G28), .b(G359), .O(G424) );
nand2 gate104( .a(G32), .b(G359), .O(G425) );
nand2 gate105( .a(G362), .b(G363), .O(G426) );

  xor2  gate1947(.a(G365), .b(G364), .O(gate106inter0));
  nand2 gate1948(.a(gate106inter0), .b(s_200), .O(gate106inter1));
  and2  gate1949(.a(G365), .b(G364), .O(gate106inter2));
  inv1  gate1950(.a(s_200), .O(gate106inter3));
  inv1  gate1951(.a(s_201), .O(gate106inter4));
  nand2 gate1952(.a(gate106inter4), .b(gate106inter3), .O(gate106inter5));
  nor2  gate1953(.a(gate106inter5), .b(gate106inter2), .O(gate106inter6));
  inv1  gate1954(.a(G364), .O(gate106inter7));
  inv1  gate1955(.a(G365), .O(gate106inter8));
  nand2 gate1956(.a(gate106inter8), .b(gate106inter7), .O(gate106inter9));
  nand2 gate1957(.a(s_201), .b(gate106inter3), .O(gate106inter10));
  nor2  gate1958(.a(gate106inter10), .b(gate106inter9), .O(gate106inter11));
  nor2  gate1959(.a(gate106inter11), .b(gate106inter6), .O(gate106inter12));
  nand2 gate1960(.a(gate106inter12), .b(gate106inter1), .O(G429));

  xor2  gate1905(.a(G367), .b(G366), .O(gate107inter0));
  nand2 gate1906(.a(gate107inter0), .b(s_194), .O(gate107inter1));
  and2  gate1907(.a(G367), .b(G366), .O(gate107inter2));
  inv1  gate1908(.a(s_194), .O(gate107inter3));
  inv1  gate1909(.a(s_195), .O(gate107inter4));
  nand2 gate1910(.a(gate107inter4), .b(gate107inter3), .O(gate107inter5));
  nor2  gate1911(.a(gate107inter5), .b(gate107inter2), .O(gate107inter6));
  inv1  gate1912(.a(G366), .O(gate107inter7));
  inv1  gate1913(.a(G367), .O(gate107inter8));
  nand2 gate1914(.a(gate107inter8), .b(gate107inter7), .O(gate107inter9));
  nand2 gate1915(.a(s_195), .b(gate107inter3), .O(gate107inter10));
  nor2  gate1916(.a(gate107inter10), .b(gate107inter9), .O(gate107inter11));
  nor2  gate1917(.a(gate107inter11), .b(gate107inter6), .O(gate107inter12));
  nand2 gate1918(.a(gate107inter12), .b(gate107inter1), .O(G432));

  xor2  gate1121(.a(G369), .b(G368), .O(gate108inter0));
  nand2 gate1122(.a(gate108inter0), .b(s_82), .O(gate108inter1));
  and2  gate1123(.a(G369), .b(G368), .O(gate108inter2));
  inv1  gate1124(.a(s_82), .O(gate108inter3));
  inv1  gate1125(.a(s_83), .O(gate108inter4));
  nand2 gate1126(.a(gate108inter4), .b(gate108inter3), .O(gate108inter5));
  nor2  gate1127(.a(gate108inter5), .b(gate108inter2), .O(gate108inter6));
  inv1  gate1128(.a(G368), .O(gate108inter7));
  inv1  gate1129(.a(G369), .O(gate108inter8));
  nand2 gate1130(.a(gate108inter8), .b(gate108inter7), .O(gate108inter9));
  nand2 gate1131(.a(s_83), .b(gate108inter3), .O(gate108inter10));
  nor2  gate1132(.a(gate108inter10), .b(gate108inter9), .O(gate108inter11));
  nor2  gate1133(.a(gate108inter11), .b(gate108inter6), .O(gate108inter12));
  nand2 gate1134(.a(gate108inter12), .b(gate108inter1), .O(G435));

  xor2  gate1695(.a(G371), .b(G370), .O(gate109inter0));
  nand2 gate1696(.a(gate109inter0), .b(s_164), .O(gate109inter1));
  and2  gate1697(.a(G371), .b(G370), .O(gate109inter2));
  inv1  gate1698(.a(s_164), .O(gate109inter3));
  inv1  gate1699(.a(s_165), .O(gate109inter4));
  nand2 gate1700(.a(gate109inter4), .b(gate109inter3), .O(gate109inter5));
  nor2  gate1701(.a(gate109inter5), .b(gate109inter2), .O(gate109inter6));
  inv1  gate1702(.a(G370), .O(gate109inter7));
  inv1  gate1703(.a(G371), .O(gate109inter8));
  nand2 gate1704(.a(gate109inter8), .b(gate109inter7), .O(gate109inter9));
  nand2 gate1705(.a(s_165), .b(gate109inter3), .O(gate109inter10));
  nor2  gate1706(.a(gate109inter10), .b(gate109inter9), .O(gate109inter11));
  nor2  gate1707(.a(gate109inter11), .b(gate109inter6), .O(gate109inter12));
  nand2 gate1708(.a(gate109inter12), .b(gate109inter1), .O(G438));
nand2 gate110( .a(G372), .b(G373), .O(G441) );

  xor2  gate659(.a(G375), .b(G374), .O(gate111inter0));
  nand2 gate660(.a(gate111inter0), .b(s_16), .O(gate111inter1));
  and2  gate661(.a(G375), .b(G374), .O(gate111inter2));
  inv1  gate662(.a(s_16), .O(gate111inter3));
  inv1  gate663(.a(s_17), .O(gate111inter4));
  nand2 gate664(.a(gate111inter4), .b(gate111inter3), .O(gate111inter5));
  nor2  gate665(.a(gate111inter5), .b(gate111inter2), .O(gate111inter6));
  inv1  gate666(.a(G374), .O(gate111inter7));
  inv1  gate667(.a(G375), .O(gate111inter8));
  nand2 gate668(.a(gate111inter8), .b(gate111inter7), .O(gate111inter9));
  nand2 gate669(.a(s_17), .b(gate111inter3), .O(gate111inter10));
  nor2  gate670(.a(gate111inter10), .b(gate111inter9), .O(gate111inter11));
  nor2  gate671(.a(gate111inter11), .b(gate111inter6), .O(gate111inter12));
  nand2 gate672(.a(gate111inter12), .b(gate111inter1), .O(G444));
nand2 gate112( .a(G376), .b(G377), .O(G447) );
nand2 gate113( .a(G378), .b(G379), .O(G450) );
nand2 gate114( .a(G380), .b(G381), .O(G453) );
nand2 gate115( .a(G382), .b(G383), .O(G456) );
nand2 gate116( .a(G384), .b(G385), .O(G459) );
nand2 gate117( .a(G386), .b(G387), .O(G462) );
nand2 gate118( .a(G388), .b(G389), .O(G465) );
nand2 gate119( .a(G390), .b(G391), .O(G468) );
nand2 gate120( .a(G392), .b(G393), .O(G471) );
nand2 gate121( .a(G394), .b(G395), .O(G474) );

  xor2  gate1653(.a(G397), .b(G396), .O(gate122inter0));
  nand2 gate1654(.a(gate122inter0), .b(s_158), .O(gate122inter1));
  and2  gate1655(.a(G397), .b(G396), .O(gate122inter2));
  inv1  gate1656(.a(s_158), .O(gate122inter3));
  inv1  gate1657(.a(s_159), .O(gate122inter4));
  nand2 gate1658(.a(gate122inter4), .b(gate122inter3), .O(gate122inter5));
  nor2  gate1659(.a(gate122inter5), .b(gate122inter2), .O(gate122inter6));
  inv1  gate1660(.a(G396), .O(gate122inter7));
  inv1  gate1661(.a(G397), .O(gate122inter8));
  nand2 gate1662(.a(gate122inter8), .b(gate122inter7), .O(gate122inter9));
  nand2 gate1663(.a(s_159), .b(gate122inter3), .O(gate122inter10));
  nor2  gate1664(.a(gate122inter10), .b(gate122inter9), .O(gate122inter11));
  nor2  gate1665(.a(gate122inter11), .b(gate122inter6), .O(gate122inter12));
  nand2 gate1666(.a(gate122inter12), .b(gate122inter1), .O(G477));
nand2 gate123( .a(G398), .b(G399), .O(G480) );

  xor2  gate2045(.a(G401), .b(G400), .O(gate124inter0));
  nand2 gate2046(.a(gate124inter0), .b(s_214), .O(gate124inter1));
  and2  gate2047(.a(G401), .b(G400), .O(gate124inter2));
  inv1  gate2048(.a(s_214), .O(gate124inter3));
  inv1  gate2049(.a(s_215), .O(gate124inter4));
  nand2 gate2050(.a(gate124inter4), .b(gate124inter3), .O(gate124inter5));
  nor2  gate2051(.a(gate124inter5), .b(gate124inter2), .O(gate124inter6));
  inv1  gate2052(.a(G400), .O(gate124inter7));
  inv1  gate2053(.a(G401), .O(gate124inter8));
  nand2 gate2054(.a(gate124inter8), .b(gate124inter7), .O(gate124inter9));
  nand2 gate2055(.a(s_215), .b(gate124inter3), .O(gate124inter10));
  nor2  gate2056(.a(gate124inter10), .b(gate124inter9), .O(gate124inter11));
  nor2  gate2057(.a(gate124inter11), .b(gate124inter6), .O(gate124inter12));
  nand2 gate2058(.a(gate124inter12), .b(gate124inter1), .O(G483));
nand2 gate125( .a(G402), .b(G403), .O(G486) );
nand2 gate126( .a(G404), .b(G405), .O(G489) );
nand2 gate127( .a(G406), .b(G407), .O(G492) );
nand2 gate128( .a(G408), .b(G409), .O(G495) );
nand2 gate129( .a(G410), .b(G411), .O(G498) );
nand2 gate130( .a(G412), .b(G413), .O(G501) );
nand2 gate131( .a(G414), .b(G415), .O(G504) );
nand2 gate132( .a(G416), .b(G417), .O(G507) );
nand2 gate133( .a(G418), .b(G419), .O(G510) );
nand2 gate134( .a(G420), .b(G421), .O(G513) );
nand2 gate135( .a(G422), .b(G423), .O(G516) );
nand2 gate136( .a(G424), .b(G425), .O(G519) );
nand2 gate137( .a(G426), .b(G429), .O(G522) );

  xor2  gate1891(.a(G435), .b(G432), .O(gate138inter0));
  nand2 gate1892(.a(gate138inter0), .b(s_192), .O(gate138inter1));
  and2  gate1893(.a(G435), .b(G432), .O(gate138inter2));
  inv1  gate1894(.a(s_192), .O(gate138inter3));
  inv1  gate1895(.a(s_193), .O(gate138inter4));
  nand2 gate1896(.a(gate138inter4), .b(gate138inter3), .O(gate138inter5));
  nor2  gate1897(.a(gate138inter5), .b(gate138inter2), .O(gate138inter6));
  inv1  gate1898(.a(G432), .O(gate138inter7));
  inv1  gate1899(.a(G435), .O(gate138inter8));
  nand2 gate1900(.a(gate138inter8), .b(gate138inter7), .O(gate138inter9));
  nand2 gate1901(.a(s_193), .b(gate138inter3), .O(gate138inter10));
  nor2  gate1902(.a(gate138inter10), .b(gate138inter9), .O(gate138inter11));
  nor2  gate1903(.a(gate138inter11), .b(gate138inter6), .O(gate138inter12));
  nand2 gate1904(.a(gate138inter12), .b(gate138inter1), .O(G525));
nand2 gate139( .a(G438), .b(G441), .O(G528) );
nand2 gate140( .a(G444), .b(G447), .O(G531) );
nand2 gate141( .a(G450), .b(G453), .O(G534) );
nand2 gate142( .a(G456), .b(G459), .O(G537) );

  xor2  gate827(.a(G465), .b(G462), .O(gate143inter0));
  nand2 gate828(.a(gate143inter0), .b(s_40), .O(gate143inter1));
  and2  gate829(.a(G465), .b(G462), .O(gate143inter2));
  inv1  gate830(.a(s_40), .O(gate143inter3));
  inv1  gate831(.a(s_41), .O(gate143inter4));
  nand2 gate832(.a(gate143inter4), .b(gate143inter3), .O(gate143inter5));
  nor2  gate833(.a(gate143inter5), .b(gate143inter2), .O(gate143inter6));
  inv1  gate834(.a(G462), .O(gate143inter7));
  inv1  gate835(.a(G465), .O(gate143inter8));
  nand2 gate836(.a(gate143inter8), .b(gate143inter7), .O(gate143inter9));
  nand2 gate837(.a(s_41), .b(gate143inter3), .O(gate143inter10));
  nor2  gate838(.a(gate143inter10), .b(gate143inter9), .O(gate143inter11));
  nor2  gate839(.a(gate143inter11), .b(gate143inter6), .O(gate143inter12));
  nand2 gate840(.a(gate143inter12), .b(gate143inter1), .O(G540));
nand2 gate144( .a(G468), .b(G471), .O(G543) );

  xor2  gate603(.a(G477), .b(G474), .O(gate145inter0));
  nand2 gate604(.a(gate145inter0), .b(s_8), .O(gate145inter1));
  and2  gate605(.a(G477), .b(G474), .O(gate145inter2));
  inv1  gate606(.a(s_8), .O(gate145inter3));
  inv1  gate607(.a(s_9), .O(gate145inter4));
  nand2 gate608(.a(gate145inter4), .b(gate145inter3), .O(gate145inter5));
  nor2  gate609(.a(gate145inter5), .b(gate145inter2), .O(gate145inter6));
  inv1  gate610(.a(G474), .O(gate145inter7));
  inv1  gate611(.a(G477), .O(gate145inter8));
  nand2 gate612(.a(gate145inter8), .b(gate145inter7), .O(gate145inter9));
  nand2 gate613(.a(s_9), .b(gate145inter3), .O(gate145inter10));
  nor2  gate614(.a(gate145inter10), .b(gate145inter9), .O(gate145inter11));
  nor2  gate615(.a(gate145inter11), .b(gate145inter6), .O(gate145inter12));
  nand2 gate616(.a(gate145inter12), .b(gate145inter1), .O(G546));
nand2 gate146( .a(G480), .b(G483), .O(G549) );
nand2 gate147( .a(G486), .b(G489), .O(G552) );

  xor2  gate1835(.a(G495), .b(G492), .O(gate148inter0));
  nand2 gate1836(.a(gate148inter0), .b(s_184), .O(gate148inter1));
  and2  gate1837(.a(G495), .b(G492), .O(gate148inter2));
  inv1  gate1838(.a(s_184), .O(gate148inter3));
  inv1  gate1839(.a(s_185), .O(gate148inter4));
  nand2 gate1840(.a(gate148inter4), .b(gate148inter3), .O(gate148inter5));
  nor2  gate1841(.a(gate148inter5), .b(gate148inter2), .O(gate148inter6));
  inv1  gate1842(.a(G492), .O(gate148inter7));
  inv1  gate1843(.a(G495), .O(gate148inter8));
  nand2 gate1844(.a(gate148inter8), .b(gate148inter7), .O(gate148inter9));
  nand2 gate1845(.a(s_185), .b(gate148inter3), .O(gate148inter10));
  nor2  gate1846(.a(gate148inter10), .b(gate148inter9), .O(gate148inter11));
  nor2  gate1847(.a(gate148inter11), .b(gate148inter6), .O(gate148inter12));
  nand2 gate1848(.a(gate148inter12), .b(gate148inter1), .O(G555));
nand2 gate149( .a(G498), .b(G501), .O(G558) );

  xor2  gate771(.a(G507), .b(G504), .O(gate150inter0));
  nand2 gate772(.a(gate150inter0), .b(s_32), .O(gate150inter1));
  and2  gate773(.a(G507), .b(G504), .O(gate150inter2));
  inv1  gate774(.a(s_32), .O(gate150inter3));
  inv1  gate775(.a(s_33), .O(gate150inter4));
  nand2 gate776(.a(gate150inter4), .b(gate150inter3), .O(gate150inter5));
  nor2  gate777(.a(gate150inter5), .b(gate150inter2), .O(gate150inter6));
  inv1  gate778(.a(G504), .O(gate150inter7));
  inv1  gate779(.a(G507), .O(gate150inter8));
  nand2 gate780(.a(gate150inter8), .b(gate150inter7), .O(gate150inter9));
  nand2 gate781(.a(s_33), .b(gate150inter3), .O(gate150inter10));
  nor2  gate782(.a(gate150inter10), .b(gate150inter9), .O(gate150inter11));
  nor2  gate783(.a(gate150inter11), .b(gate150inter6), .O(gate150inter12));
  nand2 gate784(.a(gate150inter12), .b(gate150inter1), .O(G561));

  xor2  gate2017(.a(G513), .b(G510), .O(gate151inter0));
  nand2 gate2018(.a(gate151inter0), .b(s_210), .O(gate151inter1));
  and2  gate2019(.a(G513), .b(G510), .O(gate151inter2));
  inv1  gate2020(.a(s_210), .O(gate151inter3));
  inv1  gate2021(.a(s_211), .O(gate151inter4));
  nand2 gate2022(.a(gate151inter4), .b(gate151inter3), .O(gate151inter5));
  nor2  gate2023(.a(gate151inter5), .b(gate151inter2), .O(gate151inter6));
  inv1  gate2024(.a(G510), .O(gate151inter7));
  inv1  gate2025(.a(G513), .O(gate151inter8));
  nand2 gate2026(.a(gate151inter8), .b(gate151inter7), .O(gate151inter9));
  nand2 gate2027(.a(s_211), .b(gate151inter3), .O(gate151inter10));
  nor2  gate2028(.a(gate151inter10), .b(gate151inter9), .O(gate151inter11));
  nor2  gate2029(.a(gate151inter11), .b(gate151inter6), .O(gate151inter12));
  nand2 gate2030(.a(gate151inter12), .b(gate151inter1), .O(G564));
nand2 gate152( .a(G516), .b(G519), .O(G567) );

  xor2  gate1009(.a(G522), .b(G426), .O(gate153inter0));
  nand2 gate1010(.a(gate153inter0), .b(s_66), .O(gate153inter1));
  and2  gate1011(.a(G522), .b(G426), .O(gate153inter2));
  inv1  gate1012(.a(s_66), .O(gate153inter3));
  inv1  gate1013(.a(s_67), .O(gate153inter4));
  nand2 gate1014(.a(gate153inter4), .b(gate153inter3), .O(gate153inter5));
  nor2  gate1015(.a(gate153inter5), .b(gate153inter2), .O(gate153inter6));
  inv1  gate1016(.a(G426), .O(gate153inter7));
  inv1  gate1017(.a(G522), .O(gate153inter8));
  nand2 gate1018(.a(gate153inter8), .b(gate153inter7), .O(gate153inter9));
  nand2 gate1019(.a(s_67), .b(gate153inter3), .O(gate153inter10));
  nor2  gate1020(.a(gate153inter10), .b(gate153inter9), .O(gate153inter11));
  nor2  gate1021(.a(gate153inter11), .b(gate153inter6), .O(gate153inter12));
  nand2 gate1022(.a(gate153inter12), .b(gate153inter1), .O(G570));

  xor2  gate1765(.a(G522), .b(G429), .O(gate154inter0));
  nand2 gate1766(.a(gate154inter0), .b(s_174), .O(gate154inter1));
  and2  gate1767(.a(G522), .b(G429), .O(gate154inter2));
  inv1  gate1768(.a(s_174), .O(gate154inter3));
  inv1  gate1769(.a(s_175), .O(gate154inter4));
  nand2 gate1770(.a(gate154inter4), .b(gate154inter3), .O(gate154inter5));
  nor2  gate1771(.a(gate154inter5), .b(gate154inter2), .O(gate154inter6));
  inv1  gate1772(.a(G429), .O(gate154inter7));
  inv1  gate1773(.a(G522), .O(gate154inter8));
  nand2 gate1774(.a(gate154inter8), .b(gate154inter7), .O(gate154inter9));
  nand2 gate1775(.a(s_175), .b(gate154inter3), .O(gate154inter10));
  nor2  gate1776(.a(gate154inter10), .b(gate154inter9), .O(gate154inter11));
  nor2  gate1777(.a(gate154inter11), .b(gate154inter6), .O(gate154inter12));
  nand2 gate1778(.a(gate154inter12), .b(gate154inter1), .O(G571));
nand2 gate155( .a(G432), .b(G525), .O(G572) );

  xor2  gate2101(.a(G525), .b(G435), .O(gate156inter0));
  nand2 gate2102(.a(gate156inter0), .b(s_222), .O(gate156inter1));
  and2  gate2103(.a(G525), .b(G435), .O(gate156inter2));
  inv1  gate2104(.a(s_222), .O(gate156inter3));
  inv1  gate2105(.a(s_223), .O(gate156inter4));
  nand2 gate2106(.a(gate156inter4), .b(gate156inter3), .O(gate156inter5));
  nor2  gate2107(.a(gate156inter5), .b(gate156inter2), .O(gate156inter6));
  inv1  gate2108(.a(G435), .O(gate156inter7));
  inv1  gate2109(.a(G525), .O(gate156inter8));
  nand2 gate2110(.a(gate156inter8), .b(gate156inter7), .O(gate156inter9));
  nand2 gate2111(.a(s_223), .b(gate156inter3), .O(gate156inter10));
  nor2  gate2112(.a(gate156inter10), .b(gate156inter9), .O(gate156inter11));
  nor2  gate2113(.a(gate156inter11), .b(gate156inter6), .O(gate156inter12));
  nand2 gate2114(.a(gate156inter12), .b(gate156inter1), .O(G573));

  xor2  gate1149(.a(G528), .b(G438), .O(gate157inter0));
  nand2 gate1150(.a(gate157inter0), .b(s_86), .O(gate157inter1));
  and2  gate1151(.a(G528), .b(G438), .O(gate157inter2));
  inv1  gate1152(.a(s_86), .O(gate157inter3));
  inv1  gate1153(.a(s_87), .O(gate157inter4));
  nand2 gate1154(.a(gate157inter4), .b(gate157inter3), .O(gate157inter5));
  nor2  gate1155(.a(gate157inter5), .b(gate157inter2), .O(gate157inter6));
  inv1  gate1156(.a(G438), .O(gate157inter7));
  inv1  gate1157(.a(G528), .O(gate157inter8));
  nand2 gate1158(.a(gate157inter8), .b(gate157inter7), .O(gate157inter9));
  nand2 gate1159(.a(s_87), .b(gate157inter3), .O(gate157inter10));
  nor2  gate1160(.a(gate157inter10), .b(gate157inter9), .O(gate157inter11));
  nor2  gate1161(.a(gate157inter11), .b(gate157inter6), .O(gate157inter12));
  nand2 gate1162(.a(gate157inter12), .b(gate157inter1), .O(G574));
nand2 gate158( .a(G441), .b(G528), .O(G575) );
nand2 gate159( .a(G444), .b(G531), .O(G576) );
nand2 gate160( .a(G447), .b(G531), .O(G577) );

  xor2  gate1079(.a(G534), .b(G450), .O(gate161inter0));
  nand2 gate1080(.a(gate161inter0), .b(s_76), .O(gate161inter1));
  and2  gate1081(.a(G534), .b(G450), .O(gate161inter2));
  inv1  gate1082(.a(s_76), .O(gate161inter3));
  inv1  gate1083(.a(s_77), .O(gate161inter4));
  nand2 gate1084(.a(gate161inter4), .b(gate161inter3), .O(gate161inter5));
  nor2  gate1085(.a(gate161inter5), .b(gate161inter2), .O(gate161inter6));
  inv1  gate1086(.a(G450), .O(gate161inter7));
  inv1  gate1087(.a(G534), .O(gate161inter8));
  nand2 gate1088(.a(gate161inter8), .b(gate161inter7), .O(gate161inter9));
  nand2 gate1089(.a(s_77), .b(gate161inter3), .O(gate161inter10));
  nor2  gate1090(.a(gate161inter10), .b(gate161inter9), .O(gate161inter11));
  nor2  gate1091(.a(gate161inter11), .b(gate161inter6), .O(gate161inter12));
  nand2 gate1092(.a(gate161inter12), .b(gate161inter1), .O(G578));
nand2 gate162( .a(G453), .b(G534), .O(G579) );
nand2 gate163( .a(G456), .b(G537), .O(G580) );
nand2 gate164( .a(G459), .b(G537), .O(G581) );
nand2 gate165( .a(G462), .b(G540), .O(G582) );
nand2 gate166( .a(G465), .b(G540), .O(G583) );
nand2 gate167( .a(G468), .b(G543), .O(G584) );
nand2 gate168( .a(G471), .b(G543), .O(G585) );
nand2 gate169( .a(G474), .b(G546), .O(G586) );

  xor2  gate1485(.a(G546), .b(G477), .O(gate170inter0));
  nand2 gate1486(.a(gate170inter0), .b(s_134), .O(gate170inter1));
  and2  gate1487(.a(G546), .b(G477), .O(gate170inter2));
  inv1  gate1488(.a(s_134), .O(gate170inter3));
  inv1  gate1489(.a(s_135), .O(gate170inter4));
  nand2 gate1490(.a(gate170inter4), .b(gate170inter3), .O(gate170inter5));
  nor2  gate1491(.a(gate170inter5), .b(gate170inter2), .O(gate170inter6));
  inv1  gate1492(.a(G477), .O(gate170inter7));
  inv1  gate1493(.a(G546), .O(gate170inter8));
  nand2 gate1494(.a(gate170inter8), .b(gate170inter7), .O(gate170inter9));
  nand2 gate1495(.a(s_135), .b(gate170inter3), .O(gate170inter10));
  nor2  gate1496(.a(gate170inter10), .b(gate170inter9), .O(gate170inter11));
  nor2  gate1497(.a(gate170inter11), .b(gate170inter6), .O(gate170inter12));
  nand2 gate1498(.a(gate170inter12), .b(gate170inter1), .O(G587));
nand2 gate171( .a(G480), .b(G549), .O(G588) );
nand2 gate172( .a(G483), .b(G549), .O(G589) );
nand2 gate173( .a(G486), .b(G552), .O(G590) );
nand2 gate174( .a(G489), .b(G552), .O(G591) );
nand2 gate175( .a(G492), .b(G555), .O(G592) );
nand2 gate176( .a(G495), .b(G555), .O(G593) );
nand2 gate177( .a(G498), .b(G558), .O(G594) );
nand2 gate178( .a(G501), .b(G558), .O(G595) );
nand2 gate179( .a(G504), .b(G561), .O(G596) );

  xor2  gate1849(.a(G561), .b(G507), .O(gate180inter0));
  nand2 gate1850(.a(gate180inter0), .b(s_186), .O(gate180inter1));
  and2  gate1851(.a(G561), .b(G507), .O(gate180inter2));
  inv1  gate1852(.a(s_186), .O(gate180inter3));
  inv1  gate1853(.a(s_187), .O(gate180inter4));
  nand2 gate1854(.a(gate180inter4), .b(gate180inter3), .O(gate180inter5));
  nor2  gate1855(.a(gate180inter5), .b(gate180inter2), .O(gate180inter6));
  inv1  gate1856(.a(G507), .O(gate180inter7));
  inv1  gate1857(.a(G561), .O(gate180inter8));
  nand2 gate1858(.a(gate180inter8), .b(gate180inter7), .O(gate180inter9));
  nand2 gate1859(.a(s_187), .b(gate180inter3), .O(gate180inter10));
  nor2  gate1860(.a(gate180inter10), .b(gate180inter9), .O(gate180inter11));
  nor2  gate1861(.a(gate180inter11), .b(gate180inter6), .O(gate180inter12));
  nand2 gate1862(.a(gate180inter12), .b(gate180inter1), .O(G597));

  xor2  gate1303(.a(G564), .b(G510), .O(gate181inter0));
  nand2 gate1304(.a(gate181inter0), .b(s_108), .O(gate181inter1));
  and2  gate1305(.a(G564), .b(G510), .O(gate181inter2));
  inv1  gate1306(.a(s_108), .O(gate181inter3));
  inv1  gate1307(.a(s_109), .O(gate181inter4));
  nand2 gate1308(.a(gate181inter4), .b(gate181inter3), .O(gate181inter5));
  nor2  gate1309(.a(gate181inter5), .b(gate181inter2), .O(gate181inter6));
  inv1  gate1310(.a(G510), .O(gate181inter7));
  inv1  gate1311(.a(G564), .O(gate181inter8));
  nand2 gate1312(.a(gate181inter8), .b(gate181inter7), .O(gate181inter9));
  nand2 gate1313(.a(s_109), .b(gate181inter3), .O(gate181inter10));
  nor2  gate1314(.a(gate181inter10), .b(gate181inter9), .O(gate181inter11));
  nor2  gate1315(.a(gate181inter11), .b(gate181inter6), .O(gate181inter12));
  nand2 gate1316(.a(gate181inter12), .b(gate181inter1), .O(G598));
nand2 gate182( .a(G513), .b(G564), .O(G599) );
nand2 gate183( .a(G516), .b(G567), .O(G600) );
nand2 gate184( .a(G519), .b(G567), .O(G601) );
nand2 gate185( .a(G570), .b(G571), .O(G602) );

  xor2  gate1429(.a(G573), .b(G572), .O(gate186inter0));
  nand2 gate1430(.a(gate186inter0), .b(s_126), .O(gate186inter1));
  and2  gate1431(.a(G573), .b(G572), .O(gate186inter2));
  inv1  gate1432(.a(s_126), .O(gate186inter3));
  inv1  gate1433(.a(s_127), .O(gate186inter4));
  nand2 gate1434(.a(gate186inter4), .b(gate186inter3), .O(gate186inter5));
  nor2  gate1435(.a(gate186inter5), .b(gate186inter2), .O(gate186inter6));
  inv1  gate1436(.a(G572), .O(gate186inter7));
  inv1  gate1437(.a(G573), .O(gate186inter8));
  nand2 gate1438(.a(gate186inter8), .b(gate186inter7), .O(gate186inter9));
  nand2 gate1439(.a(s_127), .b(gate186inter3), .O(gate186inter10));
  nor2  gate1440(.a(gate186inter10), .b(gate186inter9), .O(gate186inter11));
  nor2  gate1441(.a(gate186inter11), .b(gate186inter6), .O(gate186inter12));
  nand2 gate1442(.a(gate186inter12), .b(gate186inter1), .O(G607));
nand2 gate187( .a(G574), .b(G575), .O(G612) );
nand2 gate188( .a(G576), .b(G577), .O(G617) );
nand2 gate189( .a(G578), .b(G579), .O(G622) );
nand2 gate190( .a(G580), .b(G581), .O(G627) );
nand2 gate191( .a(G582), .b(G583), .O(G632) );
nand2 gate192( .a(G584), .b(G585), .O(G637) );

  xor2  gate589(.a(G587), .b(G586), .O(gate193inter0));
  nand2 gate590(.a(gate193inter0), .b(s_6), .O(gate193inter1));
  and2  gate591(.a(G587), .b(G586), .O(gate193inter2));
  inv1  gate592(.a(s_6), .O(gate193inter3));
  inv1  gate593(.a(s_7), .O(gate193inter4));
  nand2 gate594(.a(gate193inter4), .b(gate193inter3), .O(gate193inter5));
  nor2  gate595(.a(gate193inter5), .b(gate193inter2), .O(gate193inter6));
  inv1  gate596(.a(G586), .O(gate193inter7));
  inv1  gate597(.a(G587), .O(gate193inter8));
  nand2 gate598(.a(gate193inter8), .b(gate193inter7), .O(gate193inter9));
  nand2 gate599(.a(s_7), .b(gate193inter3), .O(gate193inter10));
  nor2  gate600(.a(gate193inter10), .b(gate193inter9), .O(gate193inter11));
  nor2  gate601(.a(gate193inter11), .b(gate193inter6), .O(gate193inter12));
  nand2 gate602(.a(gate193inter12), .b(gate193inter1), .O(G642));
nand2 gate194( .a(G588), .b(G589), .O(G645) );
nand2 gate195( .a(G590), .b(G591), .O(G648) );
nand2 gate196( .a(G592), .b(G593), .O(G651) );
nand2 gate197( .a(G594), .b(G595), .O(G654) );
nand2 gate198( .a(G596), .b(G597), .O(G657) );
nand2 gate199( .a(G598), .b(G599), .O(G660) );
nand2 gate200( .a(G600), .b(G601), .O(G663) );

  xor2  gate1093(.a(G607), .b(G602), .O(gate201inter0));
  nand2 gate1094(.a(gate201inter0), .b(s_78), .O(gate201inter1));
  and2  gate1095(.a(G607), .b(G602), .O(gate201inter2));
  inv1  gate1096(.a(s_78), .O(gate201inter3));
  inv1  gate1097(.a(s_79), .O(gate201inter4));
  nand2 gate1098(.a(gate201inter4), .b(gate201inter3), .O(gate201inter5));
  nor2  gate1099(.a(gate201inter5), .b(gate201inter2), .O(gate201inter6));
  inv1  gate1100(.a(G602), .O(gate201inter7));
  inv1  gate1101(.a(G607), .O(gate201inter8));
  nand2 gate1102(.a(gate201inter8), .b(gate201inter7), .O(gate201inter9));
  nand2 gate1103(.a(s_79), .b(gate201inter3), .O(gate201inter10));
  nor2  gate1104(.a(gate201inter10), .b(gate201inter9), .O(gate201inter11));
  nor2  gate1105(.a(gate201inter11), .b(gate201inter6), .O(gate201inter12));
  nand2 gate1106(.a(gate201inter12), .b(gate201inter1), .O(G666));
nand2 gate202( .a(G612), .b(G617), .O(G669) );
nand2 gate203( .a(G602), .b(G612), .O(G672) );

  xor2  gate1723(.a(G617), .b(G607), .O(gate204inter0));
  nand2 gate1724(.a(gate204inter0), .b(s_168), .O(gate204inter1));
  and2  gate1725(.a(G617), .b(G607), .O(gate204inter2));
  inv1  gate1726(.a(s_168), .O(gate204inter3));
  inv1  gate1727(.a(s_169), .O(gate204inter4));
  nand2 gate1728(.a(gate204inter4), .b(gate204inter3), .O(gate204inter5));
  nor2  gate1729(.a(gate204inter5), .b(gate204inter2), .O(gate204inter6));
  inv1  gate1730(.a(G607), .O(gate204inter7));
  inv1  gate1731(.a(G617), .O(gate204inter8));
  nand2 gate1732(.a(gate204inter8), .b(gate204inter7), .O(gate204inter9));
  nand2 gate1733(.a(s_169), .b(gate204inter3), .O(gate204inter10));
  nor2  gate1734(.a(gate204inter10), .b(gate204inter9), .O(gate204inter11));
  nor2  gate1735(.a(gate204inter11), .b(gate204inter6), .O(gate204inter12));
  nand2 gate1736(.a(gate204inter12), .b(gate204inter1), .O(G675));
nand2 gate205( .a(G622), .b(G627), .O(G678) );
nand2 gate206( .a(G632), .b(G637), .O(G681) );

  xor2  gate813(.a(G632), .b(G622), .O(gate207inter0));
  nand2 gate814(.a(gate207inter0), .b(s_38), .O(gate207inter1));
  and2  gate815(.a(G632), .b(G622), .O(gate207inter2));
  inv1  gate816(.a(s_38), .O(gate207inter3));
  inv1  gate817(.a(s_39), .O(gate207inter4));
  nand2 gate818(.a(gate207inter4), .b(gate207inter3), .O(gate207inter5));
  nor2  gate819(.a(gate207inter5), .b(gate207inter2), .O(gate207inter6));
  inv1  gate820(.a(G622), .O(gate207inter7));
  inv1  gate821(.a(G632), .O(gate207inter8));
  nand2 gate822(.a(gate207inter8), .b(gate207inter7), .O(gate207inter9));
  nand2 gate823(.a(s_39), .b(gate207inter3), .O(gate207inter10));
  nor2  gate824(.a(gate207inter10), .b(gate207inter9), .O(gate207inter11));
  nor2  gate825(.a(gate207inter11), .b(gate207inter6), .O(gate207inter12));
  nand2 gate826(.a(gate207inter12), .b(gate207inter1), .O(G684));
nand2 gate208( .a(G627), .b(G637), .O(G687) );
nand2 gate209( .a(G602), .b(G666), .O(G690) );
nand2 gate210( .a(G607), .b(G666), .O(G691) );
nand2 gate211( .a(G612), .b(G669), .O(G692) );

  xor2  gate729(.a(G669), .b(G617), .O(gate212inter0));
  nand2 gate730(.a(gate212inter0), .b(s_26), .O(gate212inter1));
  and2  gate731(.a(G669), .b(G617), .O(gate212inter2));
  inv1  gate732(.a(s_26), .O(gate212inter3));
  inv1  gate733(.a(s_27), .O(gate212inter4));
  nand2 gate734(.a(gate212inter4), .b(gate212inter3), .O(gate212inter5));
  nor2  gate735(.a(gate212inter5), .b(gate212inter2), .O(gate212inter6));
  inv1  gate736(.a(G617), .O(gate212inter7));
  inv1  gate737(.a(G669), .O(gate212inter8));
  nand2 gate738(.a(gate212inter8), .b(gate212inter7), .O(gate212inter9));
  nand2 gate739(.a(s_27), .b(gate212inter3), .O(gate212inter10));
  nor2  gate740(.a(gate212inter10), .b(gate212inter9), .O(gate212inter11));
  nor2  gate741(.a(gate212inter11), .b(gate212inter6), .O(gate212inter12));
  nand2 gate742(.a(gate212inter12), .b(gate212inter1), .O(G693));
nand2 gate213( .a(G602), .b(G672), .O(G694) );
nand2 gate214( .a(G612), .b(G672), .O(G695) );

  xor2  gate1163(.a(G675), .b(G607), .O(gate215inter0));
  nand2 gate1164(.a(gate215inter0), .b(s_88), .O(gate215inter1));
  and2  gate1165(.a(G675), .b(G607), .O(gate215inter2));
  inv1  gate1166(.a(s_88), .O(gate215inter3));
  inv1  gate1167(.a(s_89), .O(gate215inter4));
  nand2 gate1168(.a(gate215inter4), .b(gate215inter3), .O(gate215inter5));
  nor2  gate1169(.a(gate215inter5), .b(gate215inter2), .O(gate215inter6));
  inv1  gate1170(.a(G607), .O(gate215inter7));
  inv1  gate1171(.a(G675), .O(gate215inter8));
  nand2 gate1172(.a(gate215inter8), .b(gate215inter7), .O(gate215inter9));
  nand2 gate1173(.a(s_89), .b(gate215inter3), .O(gate215inter10));
  nor2  gate1174(.a(gate215inter10), .b(gate215inter9), .O(gate215inter11));
  nor2  gate1175(.a(gate215inter11), .b(gate215inter6), .O(gate215inter12));
  nand2 gate1176(.a(gate215inter12), .b(gate215inter1), .O(G696));
nand2 gate216( .a(G617), .b(G675), .O(G697) );

  xor2  gate1821(.a(G678), .b(G622), .O(gate217inter0));
  nand2 gate1822(.a(gate217inter0), .b(s_182), .O(gate217inter1));
  and2  gate1823(.a(G678), .b(G622), .O(gate217inter2));
  inv1  gate1824(.a(s_182), .O(gate217inter3));
  inv1  gate1825(.a(s_183), .O(gate217inter4));
  nand2 gate1826(.a(gate217inter4), .b(gate217inter3), .O(gate217inter5));
  nor2  gate1827(.a(gate217inter5), .b(gate217inter2), .O(gate217inter6));
  inv1  gate1828(.a(G622), .O(gate217inter7));
  inv1  gate1829(.a(G678), .O(gate217inter8));
  nand2 gate1830(.a(gate217inter8), .b(gate217inter7), .O(gate217inter9));
  nand2 gate1831(.a(s_183), .b(gate217inter3), .O(gate217inter10));
  nor2  gate1832(.a(gate217inter10), .b(gate217inter9), .O(gate217inter11));
  nor2  gate1833(.a(gate217inter11), .b(gate217inter6), .O(gate217inter12));
  nand2 gate1834(.a(gate217inter12), .b(gate217inter1), .O(G698));
nand2 gate218( .a(G627), .b(G678), .O(G699) );

  xor2  gate2073(.a(G681), .b(G632), .O(gate219inter0));
  nand2 gate2074(.a(gate219inter0), .b(s_218), .O(gate219inter1));
  and2  gate2075(.a(G681), .b(G632), .O(gate219inter2));
  inv1  gate2076(.a(s_218), .O(gate219inter3));
  inv1  gate2077(.a(s_219), .O(gate219inter4));
  nand2 gate2078(.a(gate219inter4), .b(gate219inter3), .O(gate219inter5));
  nor2  gate2079(.a(gate219inter5), .b(gate219inter2), .O(gate219inter6));
  inv1  gate2080(.a(G632), .O(gate219inter7));
  inv1  gate2081(.a(G681), .O(gate219inter8));
  nand2 gate2082(.a(gate219inter8), .b(gate219inter7), .O(gate219inter9));
  nand2 gate2083(.a(s_219), .b(gate219inter3), .O(gate219inter10));
  nor2  gate2084(.a(gate219inter10), .b(gate219inter9), .O(gate219inter11));
  nor2  gate2085(.a(gate219inter11), .b(gate219inter6), .O(gate219inter12));
  nand2 gate2086(.a(gate219inter12), .b(gate219inter1), .O(G700));

  xor2  gate1597(.a(G681), .b(G637), .O(gate220inter0));
  nand2 gate1598(.a(gate220inter0), .b(s_150), .O(gate220inter1));
  and2  gate1599(.a(G681), .b(G637), .O(gate220inter2));
  inv1  gate1600(.a(s_150), .O(gate220inter3));
  inv1  gate1601(.a(s_151), .O(gate220inter4));
  nand2 gate1602(.a(gate220inter4), .b(gate220inter3), .O(gate220inter5));
  nor2  gate1603(.a(gate220inter5), .b(gate220inter2), .O(gate220inter6));
  inv1  gate1604(.a(G637), .O(gate220inter7));
  inv1  gate1605(.a(G681), .O(gate220inter8));
  nand2 gate1606(.a(gate220inter8), .b(gate220inter7), .O(gate220inter9));
  nand2 gate1607(.a(s_151), .b(gate220inter3), .O(gate220inter10));
  nor2  gate1608(.a(gate220inter10), .b(gate220inter9), .O(gate220inter11));
  nor2  gate1609(.a(gate220inter11), .b(gate220inter6), .O(gate220inter12));
  nand2 gate1610(.a(gate220inter12), .b(gate220inter1), .O(G701));
nand2 gate221( .a(G622), .b(G684), .O(G702) );

  xor2  gate1289(.a(G684), .b(G632), .O(gate222inter0));
  nand2 gate1290(.a(gate222inter0), .b(s_106), .O(gate222inter1));
  and2  gate1291(.a(G684), .b(G632), .O(gate222inter2));
  inv1  gate1292(.a(s_106), .O(gate222inter3));
  inv1  gate1293(.a(s_107), .O(gate222inter4));
  nand2 gate1294(.a(gate222inter4), .b(gate222inter3), .O(gate222inter5));
  nor2  gate1295(.a(gate222inter5), .b(gate222inter2), .O(gate222inter6));
  inv1  gate1296(.a(G632), .O(gate222inter7));
  inv1  gate1297(.a(G684), .O(gate222inter8));
  nand2 gate1298(.a(gate222inter8), .b(gate222inter7), .O(gate222inter9));
  nand2 gate1299(.a(s_107), .b(gate222inter3), .O(gate222inter10));
  nor2  gate1300(.a(gate222inter10), .b(gate222inter9), .O(gate222inter11));
  nor2  gate1301(.a(gate222inter11), .b(gate222inter6), .O(gate222inter12));
  nand2 gate1302(.a(gate222inter12), .b(gate222inter1), .O(G703));
nand2 gate223( .a(G627), .b(G687), .O(G704) );

  xor2  gate1107(.a(G687), .b(G637), .O(gate224inter0));
  nand2 gate1108(.a(gate224inter0), .b(s_80), .O(gate224inter1));
  and2  gate1109(.a(G687), .b(G637), .O(gate224inter2));
  inv1  gate1110(.a(s_80), .O(gate224inter3));
  inv1  gate1111(.a(s_81), .O(gate224inter4));
  nand2 gate1112(.a(gate224inter4), .b(gate224inter3), .O(gate224inter5));
  nor2  gate1113(.a(gate224inter5), .b(gate224inter2), .O(gate224inter6));
  inv1  gate1114(.a(G637), .O(gate224inter7));
  inv1  gate1115(.a(G687), .O(gate224inter8));
  nand2 gate1116(.a(gate224inter8), .b(gate224inter7), .O(gate224inter9));
  nand2 gate1117(.a(s_81), .b(gate224inter3), .O(gate224inter10));
  nor2  gate1118(.a(gate224inter10), .b(gate224inter9), .O(gate224inter11));
  nor2  gate1119(.a(gate224inter11), .b(gate224inter6), .O(gate224inter12));
  nand2 gate1120(.a(gate224inter12), .b(gate224inter1), .O(G705));
nand2 gate225( .a(G690), .b(G691), .O(G706) );

  xor2  gate785(.a(G693), .b(G692), .O(gate226inter0));
  nand2 gate786(.a(gate226inter0), .b(s_34), .O(gate226inter1));
  and2  gate787(.a(G693), .b(G692), .O(gate226inter2));
  inv1  gate788(.a(s_34), .O(gate226inter3));
  inv1  gate789(.a(s_35), .O(gate226inter4));
  nand2 gate790(.a(gate226inter4), .b(gate226inter3), .O(gate226inter5));
  nor2  gate791(.a(gate226inter5), .b(gate226inter2), .O(gate226inter6));
  inv1  gate792(.a(G692), .O(gate226inter7));
  inv1  gate793(.a(G693), .O(gate226inter8));
  nand2 gate794(.a(gate226inter8), .b(gate226inter7), .O(gate226inter9));
  nand2 gate795(.a(s_35), .b(gate226inter3), .O(gate226inter10));
  nor2  gate796(.a(gate226inter10), .b(gate226inter9), .O(gate226inter11));
  nor2  gate797(.a(gate226inter11), .b(gate226inter6), .O(gate226inter12));
  nand2 gate798(.a(gate226inter12), .b(gate226inter1), .O(G709));
nand2 gate227( .a(G694), .b(G695), .O(G712) );
nand2 gate228( .a(G696), .b(G697), .O(G715) );
nand2 gate229( .a(G698), .b(G699), .O(G718) );

  xor2  gate2115(.a(G701), .b(G700), .O(gate230inter0));
  nand2 gate2116(.a(gate230inter0), .b(s_224), .O(gate230inter1));
  and2  gate2117(.a(G701), .b(G700), .O(gate230inter2));
  inv1  gate2118(.a(s_224), .O(gate230inter3));
  inv1  gate2119(.a(s_225), .O(gate230inter4));
  nand2 gate2120(.a(gate230inter4), .b(gate230inter3), .O(gate230inter5));
  nor2  gate2121(.a(gate230inter5), .b(gate230inter2), .O(gate230inter6));
  inv1  gate2122(.a(G700), .O(gate230inter7));
  inv1  gate2123(.a(G701), .O(gate230inter8));
  nand2 gate2124(.a(gate230inter8), .b(gate230inter7), .O(gate230inter9));
  nand2 gate2125(.a(s_225), .b(gate230inter3), .O(gate230inter10));
  nor2  gate2126(.a(gate230inter10), .b(gate230inter9), .O(gate230inter11));
  nor2  gate2127(.a(gate230inter11), .b(gate230inter6), .O(gate230inter12));
  nand2 gate2128(.a(gate230inter12), .b(gate230inter1), .O(G721));
nand2 gate231( .a(G702), .b(G703), .O(G724) );
nand2 gate232( .a(G704), .b(G705), .O(G727) );

  xor2  gate1709(.a(G718), .b(G242), .O(gate233inter0));
  nand2 gate1710(.a(gate233inter0), .b(s_166), .O(gate233inter1));
  and2  gate1711(.a(G718), .b(G242), .O(gate233inter2));
  inv1  gate1712(.a(s_166), .O(gate233inter3));
  inv1  gate1713(.a(s_167), .O(gate233inter4));
  nand2 gate1714(.a(gate233inter4), .b(gate233inter3), .O(gate233inter5));
  nor2  gate1715(.a(gate233inter5), .b(gate233inter2), .O(gate233inter6));
  inv1  gate1716(.a(G242), .O(gate233inter7));
  inv1  gate1717(.a(G718), .O(gate233inter8));
  nand2 gate1718(.a(gate233inter8), .b(gate233inter7), .O(gate233inter9));
  nand2 gate1719(.a(s_167), .b(gate233inter3), .O(gate233inter10));
  nor2  gate1720(.a(gate233inter10), .b(gate233inter9), .O(gate233inter11));
  nor2  gate1721(.a(gate233inter11), .b(gate233inter6), .O(gate233inter12));
  nand2 gate1722(.a(gate233inter12), .b(gate233inter1), .O(G730));
nand2 gate234( .a(G245), .b(G721), .O(G733) );
nand2 gate235( .a(G248), .b(G724), .O(G736) );
nand2 gate236( .a(G251), .b(G727), .O(G739) );

  xor2  gate855(.a(G706), .b(G254), .O(gate237inter0));
  nand2 gate856(.a(gate237inter0), .b(s_44), .O(gate237inter1));
  and2  gate857(.a(G706), .b(G254), .O(gate237inter2));
  inv1  gate858(.a(s_44), .O(gate237inter3));
  inv1  gate859(.a(s_45), .O(gate237inter4));
  nand2 gate860(.a(gate237inter4), .b(gate237inter3), .O(gate237inter5));
  nor2  gate861(.a(gate237inter5), .b(gate237inter2), .O(gate237inter6));
  inv1  gate862(.a(G254), .O(gate237inter7));
  inv1  gate863(.a(G706), .O(gate237inter8));
  nand2 gate864(.a(gate237inter8), .b(gate237inter7), .O(gate237inter9));
  nand2 gate865(.a(s_45), .b(gate237inter3), .O(gate237inter10));
  nor2  gate866(.a(gate237inter10), .b(gate237inter9), .O(gate237inter11));
  nor2  gate867(.a(gate237inter11), .b(gate237inter6), .O(gate237inter12));
  nand2 gate868(.a(gate237inter12), .b(gate237inter1), .O(G742));
nand2 gate238( .a(G257), .b(G709), .O(G745) );
nand2 gate239( .a(G260), .b(G712), .O(G748) );
nand2 gate240( .a(G263), .b(G715), .O(G751) );
nand2 gate241( .a(G242), .b(G730), .O(G754) );
nand2 gate242( .a(G718), .b(G730), .O(G755) );
nand2 gate243( .a(G245), .b(G733), .O(G756) );

  xor2  gate1807(.a(G733), .b(G721), .O(gate244inter0));
  nand2 gate1808(.a(gate244inter0), .b(s_180), .O(gate244inter1));
  and2  gate1809(.a(G733), .b(G721), .O(gate244inter2));
  inv1  gate1810(.a(s_180), .O(gate244inter3));
  inv1  gate1811(.a(s_181), .O(gate244inter4));
  nand2 gate1812(.a(gate244inter4), .b(gate244inter3), .O(gate244inter5));
  nor2  gate1813(.a(gate244inter5), .b(gate244inter2), .O(gate244inter6));
  inv1  gate1814(.a(G721), .O(gate244inter7));
  inv1  gate1815(.a(G733), .O(gate244inter8));
  nand2 gate1816(.a(gate244inter8), .b(gate244inter7), .O(gate244inter9));
  nand2 gate1817(.a(s_181), .b(gate244inter3), .O(gate244inter10));
  nor2  gate1818(.a(gate244inter10), .b(gate244inter9), .O(gate244inter11));
  nor2  gate1819(.a(gate244inter11), .b(gate244inter6), .O(gate244inter12));
  nand2 gate1820(.a(gate244inter12), .b(gate244inter1), .O(G757));
nand2 gate245( .a(G248), .b(G736), .O(G758) );
nand2 gate246( .a(G724), .b(G736), .O(G759) );
nand2 gate247( .a(G251), .b(G739), .O(G760) );
nand2 gate248( .a(G727), .b(G739), .O(G761) );
nand2 gate249( .a(G254), .b(G742), .O(G762) );

  xor2  gate953(.a(G742), .b(G706), .O(gate250inter0));
  nand2 gate954(.a(gate250inter0), .b(s_58), .O(gate250inter1));
  and2  gate955(.a(G742), .b(G706), .O(gate250inter2));
  inv1  gate956(.a(s_58), .O(gate250inter3));
  inv1  gate957(.a(s_59), .O(gate250inter4));
  nand2 gate958(.a(gate250inter4), .b(gate250inter3), .O(gate250inter5));
  nor2  gate959(.a(gate250inter5), .b(gate250inter2), .O(gate250inter6));
  inv1  gate960(.a(G706), .O(gate250inter7));
  inv1  gate961(.a(G742), .O(gate250inter8));
  nand2 gate962(.a(gate250inter8), .b(gate250inter7), .O(gate250inter9));
  nand2 gate963(.a(s_59), .b(gate250inter3), .O(gate250inter10));
  nor2  gate964(.a(gate250inter10), .b(gate250inter9), .O(gate250inter11));
  nor2  gate965(.a(gate250inter11), .b(gate250inter6), .O(gate250inter12));
  nand2 gate966(.a(gate250inter12), .b(gate250inter1), .O(G763));
nand2 gate251( .a(G257), .b(G745), .O(G764) );
nand2 gate252( .a(G709), .b(G745), .O(G765) );
nand2 gate253( .a(G260), .b(G748), .O(G766) );

  xor2  gate1275(.a(G748), .b(G712), .O(gate254inter0));
  nand2 gate1276(.a(gate254inter0), .b(s_104), .O(gate254inter1));
  and2  gate1277(.a(G748), .b(G712), .O(gate254inter2));
  inv1  gate1278(.a(s_104), .O(gate254inter3));
  inv1  gate1279(.a(s_105), .O(gate254inter4));
  nand2 gate1280(.a(gate254inter4), .b(gate254inter3), .O(gate254inter5));
  nor2  gate1281(.a(gate254inter5), .b(gate254inter2), .O(gate254inter6));
  inv1  gate1282(.a(G712), .O(gate254inter7));
  inv1  gate1283(.a(G748), .O(gate254inter8));
  nand2 gate1284(.a(gate254inter8), .b(gate254inter7), .O(gate254inter9));
  nand2 gate1285(.a(s_105), .b(gate254inter3), .O(gate254inter10));
  nor2  gate1286(.a(gate254inter10), .b(gate254inter9), .O(gate254inter11));
  nor2  gate1287(.a(gate254inter11), .b(gate254inter6), .O(gate254inter12));
  nand2 gate1288(.a(gate254inter12), .b(gate254inter1), .O(G767));

  xor2  gate1933(.a(G751), .b(G263), .O(gate255inter0));
  nand2 gate1934(.a(gate255inter0), .b(s_198), .O(gate255inter1));
  and2  gate1935(.a(G751), .b(G263), .O(gate255inter2));
  inv1  gate1936(.a(s_198), .O(gate255inter3));
  inv1  gate1937(.a(s_199), .O(gate255inter4));
  nand2 gate1938(.a(gate255inter4), .b(gate255inter3), .O(gate255inter5));
  nor2  gate1939(.a(gate255inter5), .b(gate255inter2), .O(gate255inter6));
  inv1  gate1940(.a(G263), .O(gate255inter7));
  inv1  gate1941(.a(G751), .O(gate255inter8));
  nand2 gate1942(.a(gate255inter8), .b(gate255inter7), .O(gate255inter9));
  nand2 gate1943(.a(s_199), .b(gate255inter3), .O(gate255inter10));
  nor2  gate1944(.a(gate255inter10), .b(gate255inter9), .O(gate255inter11));
  nor2  gate1945(.a(gate255inter11), .b(gate255inter6), .O(gate255inter12));
  nand2 gate1946(.a(gate255inter12), .b(gate255inter1), .O(G768));
nand2 gate256( .a(G715), .b(G751), .O(G769) );
nand2 gate257( .a(G754), .b(G755), .O(G770) );
nand2 gate258( .a(G756), .b(G757), .O(G773) );
nand2 gate259( .a(G758), .b(G759), .O(G776) );
nand2 gate260( .a(G760), .b(G761), .O(G779) );

  xor2  gate757(.a(G763), .b(G762), .O(gate261inter0));
  nand2 gate758(.a(gate261inter0), .b(s_30), .O(gate261inter1));
  and2  gate759(.a(G763), .b(G762), .O(gate261inter2));
  inv1  gate760(.a(s_30), .O(gate261inter3));
  inv1  gate761(.a(s_31), .O(gate261inter4));
  nand2 gate762(.a(gate261inter4), .b(gate261inter3), .O(gate261inter5));
  nor2  gate763(.a(gate261inter5), .b(gate261inter2), .O(gate261inter6));
  inv1  gate764(.a(G762), .O(gate261inter7));
  inv1  gate765(.a(G763), .O(gate261inter8));
  nand2 gate766(.a(gate261inter8), .b(gate261inter7), .O(gate261inter9));
  nand2 gate767(.a(s_31), .b(gate261inter3), .O(gate261inter10));
  nor2  gate768(.a(gate261inter10), .b(gate261inter9), .O(gate261inter11));
  nor2  gate769(.a(gate261inter11), .b(gate261inter6), .O(gate261inter12));
  nand2 gate770(.a(gate261inter12), .b(gate261inter1), .O(G782));
nand2 gate262( .a(G764), .b(G765), .O(G785) );
nand2 gate263( .a(G766), .b(G767), .O(G788) );
nand2 gate264( .a(G768), .b(G769), .O(G791) );
nand2 gate265( .a(G642), .b(G770), .O(G794) );
nand2 gate266( .a(G645), .b(G773), .O(G797) );
nand2 gate267( .a(G648), .b(G776), .O(G800) );

  xor2  gate1681(.a(G779), .b(G651), .O(gate268inter0));
  nand2 gate1682(.a(gate268inter0), .b(s_162), .O(gate268inter1));
  and2  gate1683(.a(G779), .b(G651), .O(gate268inter2));
  inv1  gate1684(.a(s_162), .O(gate268inter3));
  inv1  gate1685(.a(s_163), .O(gate268inter4));
  nand2 gate1686(.a(gate268inter4), .b(gate268inter3), .O(gate268inter5));
  nor2  gate1687(.a(gate268inter5), .b(gate268inter2), .O(gate268inter6));
  inv1  gate1688(.a(G651), .O(gate268inter7));
  inv1  gate1689(.a(G779), .O(gate268inter8));
  nand2 gate1690(.a(gate268inter8), .b(gate268inter7), .O(gate268inter9));
  nand2 gate1691(.a(s_163), .b(gate268inter3), .O(gate268inter10));
  nor2  gate1692(.a(gate268inter10), .b(gate268inter9), .O(gate268inter11));
  nor2  gate1693(.a(gate268inter11), .b(gate268inter6), .O(gate268inter12));
  nand2 gate1694(.a(gate268inter12), .b(gate268inter1), .O(G803));
nand2 gate269( .a(G654), .b(G782), .O(G806) );

  xor2  gate631(.a(G785), .b(G657), .O(gate270inter0));
  nand2 gate632(.a(gate270inter0), .b(s_12), .O(gate270inter1));
  and2  gate633(.a(G785), .b(G657), .O(gate270inter2));
  inv1  gate634(.a(s_12), .O(gate270inter3));
  inv1  gate635(.a(s_13), .O(gate270inter4));
  nand2 gate636(.a(gate270inter4), .b(gate270inter3), .O(gate270inter5));
  nor2  gate637(.a(gate270inter5), .b(gate270inter2), .O(gate270inter6));
  inv1  gate638(.a(G657), .O(gate270inter7));
  inv1  gate639(.a(G785), .O(gate270inter8));
  nand2 gate640(.a(gate270inter8), .b(gate270inter7), .O(gate270inter9));
  nand2 gate641(.a(s_13), .b(gate270inter3), .O(gate270inter10));
  nor2  gate642(.a(gate270inter10), .b(gate270inter9), .O(gate270inter11));
  nor2  gate643(.a(gate270inter11), .b(gate270inter6), .O(gate270inter12));
  nand2 gate644(.a(gate270inter12), .b(gate270inter1), .O(G809));
nand2 gate271( .a(G660), .b(G788), .O(G812) );
nand2 gate272( .a(G663), .b(G791), .O(G815) );
nand2 gate273( .a(G642), .b(G794), .O(G818) );

  xor2  gate1457(.a(G794), .b(G770), .O(gate274inter0));
  nand2 gate1458(.a(gate274inter0), .b(s_130), .O(gate274inter1));
  and2  gate1459(.a(G794), .b(G770), .O(gate274inter2));
  inv1  gate1460(.a(s_130), .O(gate274inter3));
  inv1  gate1461(.a(s_131), .O(gate274inter4));
  nand2 gate1462(.a(gate274inter4), .b(gate274inter3), .O(gate274inter5));
  nor2  gate1463(.a(gate274inter5), .b(gate274inter2), .O(gate274inter6));
  inv1  gate1464(.a(G770), .O(gate274inter7));
  inv1  gate1465(.a(G794), .O(gate274inter8));
  nand2 gate1466(.a(gate274inter8), .b(gate274inter7), .O(gate274inter9));
  nand2 gate1467(.a(s_131), .b(gate274inter3), .O(gate274inter10));
  nor2  gate1468(.a(gate274inter10), .b(gate274inter9), .O(gate274inter11));
  nor2  gate1469(.a(gate274inter11), .b(gate274inter6), .O(gate274inter12));
  nand2 gate1470(.a(gate274inter12), .b(gate274inter1), .O(G819));
nand2 gate275( .a(G645), .b(G797), .O(G820) );

  xor2  gate1401(.a(G797), .b(G773), .O(gate276inter0));
  nand2 gate1402(.a(gate276inter0), .b(s_122), .O(gate276inter1));
  and2  gate1403(.a(G797), .b(G773), .O(gate276inter2));
  inv1  gate1404(.a(s_122), .O(gate276inter3));
  inv1  gate1405(.a(s_123), .O(gate276inter4));
  nand2 gate1406(.a(gate276inter4), .b(gate276inter3), .O(gate276inter5));
  nor2  gate1407(.a(gate276inter5), .b(gate276inter2), .O(gate276inter6));
  inv1  gate1408(.a(G773), .O(gate276inter7));
  inv1  gate1409(.a(G797), .O(gate276inter8));
  nand2 gate1410(.a(gate276inter8), .b(gate276inter7), .O(gate276inter9));
  nand2 gate1411(.a(s_123), .b(gate276inter3), .O(gate276inter10));
  nor2  gate1412(.a(gate276inter10), .b(gate276inter9), .O(gate276inter11));
  nor2  gate1413(.a(gate276inter11), .b(gate276inter6), .O(gate276inter12));
  nand2 gate1414(.a(gate276inter12), .b(gate276inter1), .O(G821));
nand2 gate277( .a(G648), .b(G800), .O(G822) );
nand2 gate278( .a(G776), .b(G800), .O(G823) );
nand2 gate279( .a(G651), .b(G803), .O(G824) );
nand2 gate280( .a(G779), .b(G803), .O(G825) );
nand2 gate281( .a(G654), .b(G806), .O(G826) );
nand2 gate282( .a(G782), .b(G806), .O(G827) );

  xor2  gate2087(.a(G809), .b(G657), .O(gate283inter0));
  nand2 gate2088(.a(gate283inter0), .b(s_220), .O(gate283inter1));
  and2  gate2089(.a(G809), .b(G657), .O(gate283inter2));
  inv1  gate2090(.a(s_220), .O(gate283inter3));
  inv1  gate2091(.a(s_221), .O(gate283inter4));
  nand2 gate2092(.a(gate283inter4), .b(gate283inter3), .O(gate283inter5));
  nor2  gate2093(.a(gate283inter5), .b(gate283inter2), .O(gate283inter6));
  inv1  gate2094(.a(G657), .O(gate283inter7));
  inv1  gate2095(.a(G809), .O(gate283inter8));
  nand2 gate2096(.a(gate283inter8), .b(gate283inter7), .O(gate283inter9));
  nand2 gate2097(.a(s_221), .b(gate283inter3), .O(gate283inter10));
  nor2  gate2098(.a(gate283inter10), .b(gate283inter9), .O(gate283inter11));
  nor2  gate2099(.a(gate283inter11), .b(gate283inter6), .O(gate283inter12));
  nand2 gate2100(.a(gate283inter12), .b(gate283inter1), .O(G828));
nand2 gate284( .a(G785), .b(G809), .O(G829) );
nand2 gate285( .a(G660), .b(G812), .O(G830) );

  xor2  gate2059(.a(G812), .b(G788), .O(gate286inter0));
  nand2 gate2060(.a(gate286inter0), .b(s_216), .O(gate286inter1));
  and2  gate2061(.a(G812), .b(G788), .O(gate286inter2));
  inv1  gate2062(.a(s_216), .O(gate286inter3));
  inv1  gate2063(.a(s_217), .O(gate286inter4));
  nand2 gate2064(.a(gate286inter4), .b(gate286inter3), .O(gate286inter5));
  nor2  gate2065(.a(gate286inter5), .b(gate286inter2), .O(gate286inter6));
  inv1  gate2066(.a(G788), .O(gate286inter7));
  inv1  gate2067(.a(G812), .O(gate286inter8));
  nand2 gate2068(.a(gate286inter8), .b(gate286inter7), .O(gate286inter9));
  nand2 gate2069(.a(s_217), .b(gate286inter3), .O(gate286inter10));
  nor2  gate2070(.a(gate286inter10), .b(gate286inter9), .O(gate286inter11));
  nor2  gate2071(.a(gate286inter11), .b(gate286inter6), .O(gate286inter12));
  nand2 gate2072(.a(gate286inter12), .b(gate286inter1), .O(G831));
nand2 gate287( .a(G663), .b(G815), .O(G832) );
nand2 gate288( .a(G791), .b(G815), .O(G833) );
nand2 gate289( .a(G818), .b(G819), .O(G834) );
nand2 gate290( .a(G820), .b(G821), .O(G847) );
nand2 gate291( .a(G822), .b(G823), .O(G860) );

  xor2  gate561(.a(G825), .b(G824), .O(gate292inter0));
  nand2 gate562(.a(gate292inter0), .b(s_2), .O(gate292inter1));
  and2  gate563(.a(G825), .b(G824), .O(gate292inter2));
  inv1  gate564(.a(s_2), .O(gate292inter3));
  inv1  gate565(.a(s_3), .O(gate292inter4));
  nand2 gate566(.a(gate292inter4), .b(gate292inter3), .O(gate292inter5));
  nor2  gate567(.a(gate292inter5), .b(gate292inter2), .O(gate292inter6));
  inv1  gate568(.a(G824), .O(gate292inter7));
  inv1  gate569(.a(G825), .O(gate292inter8));
  nand2 gate570(.a(gate292inter8), .b(gate292inter7), .O(gate292inter9));
  nand2 gate571(.a(s_3), .b(gate292inter3), .O(gate292inter10));
  nor2  gate572(.a(gate292inter10), .b(gate292inter9), .O(gate292inter11));
  nor2  gate573(.a(gate292inter11), .b(gate292inter6), .O(gate292inter12));
  nand2 gate574(.a(gate292inter12), .b(gate292inter1), .O(G873));

  xor2  gate715(.a(G829), .b(G828), .O(gate293inter0));
  nand2 gate716(.a(gate293inter0), .b(s_24), .O(gate293inter1));
  and2  gate717(.a(G829), .b(G828), .O(gate293inter2));
  inv1  gate718(.a(s_24), .O(gate293inter3));
  inv1  gate719(.a(s_25), .O(gate293inter4));
  nand2 gate720(.a(gate293inter4), .b(gate293inter3), .O(gate293inter5));
  nor2  gate721(.a(gate293inter5), .b(gate293inter2), .O(gate293inter6));
  inv1  gate722(.a(G828), .O(gate293inter7));
  inv1  gate723(.a(G829), .O(gate293inter8));
  nand2 gate724(.a(gate293inter8), .b(gate293inter7), .O(gate293inter9));
  nand2 gate725(.a(s_25), .b(gate293inter3), .O(gate293inter10));
  nor2  gate726(.a(gate293inter10), .b(gate293inter9), .O(gate293inter11));
  nor2  gate727(.a(gate293inter11), .b(gate293inter6), .O(gate293inter12));
  nand2 gate728(.a(gate293inter12), .b(gate293inter1), .O(G886));
nand2 gate294( .a(G832), .b(G833), .O(G899) );
nand2 gate295( .a(G830), .b(G831), .O(G912) );
nand2 gate296( .a(G826), .b(G827), .O(G925) );
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );
nand2 gate387( .a(G1), .b(G1036), .O(G1132) );
nand2 gate388( .a(G2), .b(G1039), .O(G1135) );
nand2 gate389( .a(G3), .b(G1042), .O(G1138) );
nand2 gate390( .a(G4), .b(G1045), .O(G1141) );
nand2 gate391( .a(G5), .b(G1048), .O(G1144) );
nand2 gate392( .a(G6), .b(G1051), .O(G1147) );
nand2 gate393( .a(G7), .b(G1054), .O(G1150) );
nand2 gate394( .a(G8), .b(G1057), .O(G1153) );
nand2 gate395( .a(G9), .b(G1060), .O(G1156) );

  xor2  gate1793(.a(G1063), .b(G10), .O(gate396inter0));
  nand2 gate1794(.a(gate396inter0), .b(s_178), .O(gate396inter1));
  and2  gate1795(.a(G1063), .b(G10), .O(gate396inter2));
  inv1  gate1796(.a(s_178), .O(gate396inter3));
  inv1  gate1797(.a(s_179), .O(gate396inter4));
  nand2 gate1798(.a(gate396inter4), .b(gate396inter3), .O(gate396inter5));
  nor2  gate1799(.a(gate396inter5), .b(gate396inter2), .O(gate396inter6));
  inv1  gate1800(.a(G10), .O(gate396inter7));
  inv1  gate1801(.a(G1063), .O(gate396inter8));
  nand2 gate1802(.a(gate396inter8), .b(gate396inter7), .O(gate396inter9));
  nand2 gate1803(.a(s_179), .b(gate396inter3), .O(gate396inter10));
  nor2  gate1804(.a(gate396inter10), .b(gate396inter9), .O(gate396inter11));
  nor2  gate1805(.a(gate396inter11), .b(gate396inter6), .O(gate396inter12));
  nand2 gate1806(.a(gate396inter12), .b(gate396inter1), .O(G1159));
nand2 gate397( .a(G11), .b(G1066), .O(G1162) );
nand2 gate398( .a(G12), .b(G1069), .O(G1165) );

  xor2  gate1023(.a(G1072), .b(G13), .O(gate399inter0));
  nand2 gate1024(.a(gate399inter0), .b(s_68), .O(gate399inter1));
  and2  gate1025(.a(G1072), .b(G13), .O(gate399inter2));
  inv1  gate1026(.a(s_68), .O(gate399inter3));
  inv1  gate1027(.a(s_69), .O(gate399inter4));
  nand2 gate1028(.a(gate399inter4), .b(gate399inter3), .O(gate399inter5));
  nor2  gate1029(.a(gate399inter5), .b(gate399inter2), .O(gate399inter6));
  inv1  gate1030(.a(G13), .O(gate399inter7));
  inv1  gate1031(.a(G1072), .O(gate399inter8));
  nand2 gate1032(.a(gate399inter8), .b(gate399inter7), .O(gate399inter9));
  nand2 gate1033(.a(s_69), .b(gate399inter3), .O(gate399inter10));
  nor2  gate1034(.a(gate399inter10), .b(gate399inter9), .O(gate399inter11));
  nor2  gate1035(.a(gate399inter11), .b(gate399inter6), .O(gate399inter12));
  nand2 gate1036(.a(gate399inter12), .b(gate399inter1), .O(G1168));
nand2 gate400( .a(G14), .b(G1075), .O(G1171) );
nand2 gate401( .a(G15), .b(G1078), .O(G1174) );
nand2 gate402( .a(G16), .b(G1081), .O(G1177) );

  xor2  gate869(.a(G1084), .b(G17), .O(gate403inter0));
  nand2 gate870(.a(gate403inter0), .b(s_46), .O(gate403inter1));
  and2  gate871(.a(G1084), .b(G17), .O(gate403inter2));
  inv1  gate872(.a(s_46), .O(gate403inter3));
  inv1  gate873(.a(s_47), .O(gate403inter4));
  nand2 gate874(.a(gate403inter4), .b(gate403inter3), .O(gate403inter5));
  nor2  gate875(.a(gate403inter5), .b(gate403inter2), .O(gate403inter6));
  inv1  gate876(.a(G17), .O(gate403inter7));
  inv1  gate877(.a(G1084), .O(gate403inter8));
  nand2 gate878(.a(gate403inter8), .b(gate403inter7), .O(gate403inter9));
  nand2 gate879(.a(s_47), .b(gate403inter3), .O(gate403inter10));
  nor2  gate880(.a(gate403inter10), .b(gate403inter9), .O(gate403inter11));
  nor2  gate881(.a(gate403inter11), .b(gate403inter6), .O(gate403inter12));
  nand2 gate882(.a(gate403inter12), .b(gate403inter1), .O(G1180));
nand2 gate404( .a(G18), .b(G1087), .O(G1183) );
nand2 gate405( .a(G19), .b(G1090), .O(G1186) );

  xor2  gate1863(.a(G1093), .b(G20), .O(gate406inter0));
  nand2 gate1864(.a(gate406inter0), .b(s_188), .O(gate406inter1));
  and2  gate1865(.a(G1093), .b(G20), .O(gate406inter2));
  inv1  gate1866(.a(s_188), .O(gate406inter3));
  inv1  gate1867(.a(s_189), .O(gate406inter4));
  nand2 gate1868(.a(gate406inter4), .b(gate406inter3), .O(gate406inter5));
  nor2  gate1869(.a(gate406inter5), .b(gate406inter2), .O(gate406inter6));
  inv1  gate1870(.a(G20), .O(gate406inter7));
  inv1  gate1871(.a(G1093), .O(gate406inter8));
  nand2 gate1872(.a(gate406inter8), .b(gate406inter7), .O(gate406inter9));
  nand2 gate1873(.a(s_189), .b(gate406inter3), .O(gate406inter10));
  nor2  gate1874(.a(gate406inter10), .b(gate406inter9), .O(gate406inter11));
  nor2  gate1875(.a(gate406inter11), .b(gate406inter6), .O(gate406inter12));
  nand2 gate1876(.a(gate406inter12), .b(gate406inter1), .O(G1189));
nand2 gate407( .a(G21), .b(G1096), .O(G1192) );

  xor2  gate897(.a(G1099), .b(G22), .O(gate408inter0));
  nand2 gate898(.a(gate408inter0), .b(s_50), .O(gate408inter1));
  and2  gate899(.a(G1099), .b(G22), .O(gate408inter2));
  inv1  gate900(.a(s_50), .O(gate408inter3));
  inv1  gate901(.a(s_51), .O(gate408inter4));
  nand2 gate902(.a(gate408inter4), .b(gate408inter3), .O(gate408inter5));
  nor2  gate903(.a(gate408inter5), .b(gate408inter2), .O(gate408inter6));
  inv1  gate904(.a(G22), .O(gate408inter7));
  inv1  gate905(.a(G1099), .O(gate408inter8));
  nand2 gate906(.a(gate408inter8), .b(gate408inter7), .O(gate408inter9));
  nand2 gate907(.a(s_51), .b(gate408inter3), .O(gate408inter10));
  nor2  gate908(.a(gate408inter10), .b(gate408inter9), .O(gate408inter11));
  nor2  gate909(.a(gate408inter11), .b(gate408inter6), .O(gate408inter12));
  nand2 gate910(.a(gate408inter12), .b(gate408inter1), .O(G1195));

  xor2  gate1737(.a(G1102), .b(G23), .O(gate409inter0));
  nand2 gate1738(.a(gate409inter0), .b(s_170), .O(gate409inter1));
  and2  gate1739(.a(G1102), .b(G23), .O(gate409inter2));
  inv1  gate1740(.a(s_170), .O(gate409inter3));
  inv1  gate1741(.a(s_171), .O(gate409inter4));
  nand2 gate1742(.a(gate409inter4), .b(gate409inter3), .O(gate409inter5));
  nor2  gate1743(.a(gate409inter5), .b(gate409inter2), .O(gate409inter6));
  inv1  gate1744(.a(G23), .O(gate409inter7));
  inv1  gate1745(.a(G1102), .O(gate409inter8));
  nand2 gate1746(.a(gate409inter8), .b(gate409inter7), .O(gate409inter9));
  nand2 gate1747(.a(s_171), .b(gate409inter3), .O(gate409inter10));
  nor2  gate1748(.a(gate409inter10), .b(gate409inter9), .O(gate409inter11));
  nor2  gate1749(.a(gate409inter11), .b(gate409inter6), .O(gate409inter12));
  nand2 gate1750(.a(gate409inter12), .b(gate409inter1), .O(G1198));
nand2 gate410( .a(G24), .b(G1105), .O(G1201) );
nand2 gate411( .a(G25), .b(G1108), .O(G1204) );
nand2 gate412( .a(G26), .b(G1111), .O(G1207) );
nand2 gate413( .a(G27), .b(G1114), .O(G1210) );

  xor2  gate1247(.a(G1117), .b(G28), .O(gate414inter0));
  nand2 gate1248(.a(gate414inter0), .b(s_100), .O(gate414inter1));
  and2  gate1249(.a(G1117), .b(G28), .O(gate414inter2));
  inv1  gate1250(.a(s_100), .O(gate414inter3));
  inv1  gate1251(.a(s_101), .O(gate414inter4));
  nand2 gate1252(.a(gate414inter4), .b(gate414inter3), .O(gate414inter5));
  nor2  gate1253(.a(gate414inter5), .b(gate414inter2), .O(gate414inter6));
  inv1  gate1254(.a(G28), .O(gate414inter7));
  inv1  gate1255(.a(G1117), .O(gate414inter8));
  nand2 gate1256(.a(gate414inter8), .b(gate414inter7), .O(gate414inter9));
  nand2 gate1257(.a(s_101), .b(gate414inter3), .O(gate414inter10));
  nor2  gate1258(.a(gate414inter10), .b(gate414inter9), .O(gate414inter11));
  nor2  gate1259(.a(gate414inter11), .b(gate414inter6), .O(gate414inter12));
  nand2 gate1260(.a(gate414inter12), .b(gate414inter1), .O(G1213));
nand2 gate415( .a(G29), .b(G1120), .O(G1216) );
nand2 gate416( .a(G30), .b(G1123), .O(G1219) );
nand2 gate417( .a(G31), .b(G1126), .O(G1222) );

  xor2  gate701(.a(G1129), .b(G32), .O(gate418inter0));
  nand2 gate702(.a(gate418inter0), .b(s_22), .O(gate418inter1));
  and2  gate703(.a(G1129), .b(G32), .O(gate418inter2));
  inv1  gate704(.a(s_22), .O(gate418inter3));
  inv1  gate705(.a(s_23), .O(gate418inter4));
  nand2 gate706(.a(gate418inter4), .b(gate418inter3), .O(gate418inter5));
  nor2  gate707(.a(gate418inter5), .b(gate418inter2), .O(gate418inter6));
  inv1  gate708(.a(G32), .O(gate418inter7));
  inv1  gate709(.a(G1129), .O(gate418inter8));
  nand2 gate710(.a(gate418inter8), .b(gate418inter7), .O(gate418inter9));
  nand2 gate711(.a(s_23), .b(gate418inter3), .O(gate418inter10));
  nor2  gate712(.a(gate418inter10), .b(gate418inter9), .O(gate418inter11));
  nor2  gate713(.a(gate418inter11), .b(gate418inter6), .O(gate418inter12));
  nand2 gate714(.a(gate418inter12), .b(gate418inter1), .O(G1225));
nand2 gate419( .a(G1), .b(G1132), .O(G1228) );

  xor2  gate1177(.a(G1132), .b(G1036), .O(gate420inter0));
  nand2 gate1178(.a(gate420inter0), .b(s_90), .O(gate420inter1));
  and2  gate1179(.a(G1132), .b(G1036), .O(gate420inter2));
  inv1  gate1180(.a(s_90), .O(gate420inter3));
  inv1  gate1181(.a(s_91), .O(gate420inter4));
  nand2 gate1182(.a(gate420inter4), .b(gate420inter3), .O(gate420inter5));
  nor2  gate1183(.a(gate420inter5), .b(gate420inter2), .O(gate420inter6));
  inv1  gate1184(.a(G1036), .O(gate420inter7));
  inv1  gate1185(.a(G1132), .O(gate420inter8));
  nand2 gate1186(.a(gate420inter8), .b(gate420inter7), .O(gate420inter9));
  nand2 gate1187(.a(s_91), .b(gate420inter3), .O(gate420inter10));
  nor2  gate1188(.a(gate420inter10), .b(gate420inter9), .O(gate420inter11));
  nor2  gate1189(.a(gate420inter11), .b(gate420inter6), .O(gate420inter12));
  nand2 gate1190(.a(gate420inter12), .b(gate420inter1), .O(G1229));
nand2 gate421( .a(G2), .b(G1135), .O(G1230) );
nand2 gate422( .a(G1039), .b(G1135), .O(G1231) );

  xor2  gate925(.a(G1138), .b(G3), .O(gate423inter0));
  nand2 gate926(.a(gate423inter0), .b(s_54), .O(gate423inter1));
  and2  gate927(.a(G1138), .b(G3), .O(gate423inter2));
  inv1  gate928(.a(s_54), .O(gate423inter3));
  inv1  gate929(.a(s_55), .O(gate423inter4));
  nand2 gate930(.a(gate423inter4), .b(gate423inter3), .O(gate423inter5));
  nor2  gate931(.a(gate423inter5), .b(gate423inter2), .O(gate423inter6));
  inv1  gate932(.a(G3), .O(gate423inter7));
  inv1  gate933(.a(G1138), .O(gate423inter8));
  nand2 gate934(.a(gate423inter8), .b(gate423inter7), .O(gate423inter9));
  nand2 gate935(.a(s_55), .b(gate423inter3), .O(gate423inter10));
  nor2  gate936(.a(gate423inter10), .b(gate423inter9), .O(gate423inter11));
  nor2  gate937(.a(gate423inter11), .b(gate423inter6), .O(gate423inter12));
  nand2 gate938(.a(gate423inter12), .b(gate423inter1), .O(G1232));
nand2 gate424( .a(G1042), .b(G1138), .O(G1233) );

  xor2  gate1639(.a(G1141), .b(G4), .O(gate425inter0));
  nand2 gate1640(.a(gate425inter0), .b(s_156), .O(gate425inter1));
  and2  gate1641(.a(G1141), .b(G4), .O(gate425inter2));
  inv1  gate1642(.a(s_156), .O(gate425inter3));
  inv1  gate1643(.a(s_157), .O(gate425inter4));
  nand2 gate1644(.a(gate425inter4), .b(gate425inter3), .O(gate425inter5));
  nor2  gate1645(.a(gate425inter5), .b(gate425inter2), .O(gate425inter6));
  inv1  gate1646(.a(G4), .O(gate425inter7));
  inv1  gate1647(.a(G1141), .O(gate425inter8));
  nand2 gate1648(.a(gate425inter8), .b(gate425inter7), .O(gate425inter9));
  nand2 gate1649(.a(s_157), .b(gate425inter3), .O(gate425inter10));
  nor2  gate1650(.a(gate425inter10), .b(gate425inter9), .O(gate425inter11));
  nor2  gate1651(.a(gate425inter11), .b(gate425inter6), .O(gate425inter12));
  nand2 gate1652(.a(gate425inter12), .b(gate425inter1), .O(G1234));

  xor2  gate883(.a(G1141), .b(G1045), .O(gate426inter0));
  nand2 gate884(.a(gate426inter0), .b(s_48), .O(gate426inter1));
  and2  gate885(.a(G1141), .b(G1045), .O(gate426inter2));
  inv1  gate886(.a(s_48), .O(gate426inter3));
  inv1  gate887(.a(s_49), .O(gate426inter4));
  nand2 gate888(.a(gate426inter4), .b(gate426inter3), .O(gate426inter5));
  nor2  gate889(.a(gate426inter5), .b(gate426inter2), .O(gate426inter6));
  inv1  gate890(.a(G1045), .O(gate426inter7));
  inv1  gate891(.a(G1141), .O(gate426inter8));
  nand2 gate892(.a(gate426inter8), .b(gate426inter7), .O(gate426inter9));
  nand2 gate893(.a(s_49), .b(gate426inter3), .O(gate426inter10));
  nor2  gate894(.a(gate426inter10), .b(gate426inter9), .O(gate426inter11));
  nor2  gate895(.a(gate426inter11), .b(gate426inter6), .O(gate426inter12));
  nand2 gate896(.a(gate426inter12), .b(gate426inter1), .O(G1235));
nand2 gate427( .a(G5), .b(G1144), .O(G1236) );

  xor2  gate1919(.a(G1144), .b(G1048), .O(gate428inter0));
  nand2 gate1920(.a(gate428inter0), .b(s_196), .O(gate428inter1));
  and2  gate1921(.a(G1144), .b(G1048), .O(gate428inter2));
  inv1  gate1922(.a(s_196), .O(gate428inter3));
  inv1  gate1923(.a(s_197), .O(gate428inter4));
  nand2 gate1924(.a(gate428inter4), .b(gate428inter3), .O(gate428inter5));
  nor2  gate1925(.a(gate428inter5), .b(gate428inter2), .O(gate428inter6));
  inv1  gate1926(.a(G1048), .O(gate428inter7));
  inv1  gate1927(.a(G1144), .O(gate428inter8));
  nand2 gate1928(.a(gate428inter8), .b(gate428inter7), .O(gate428inter9));
  nand2 gate1929(.a(s_197), .b(gate428inter3), .O(gate428inter10));
  nor2  gate1930(.a(gate428inter10), .b(gate428inter9), .O(gate428inter11));
  nor2  gate1931(.a(gate428inter11), .b(gate428inter6), .O(gate428inter12));
  nand2 gate1932(.a(gate428inter12), .b(gate428inter1), .O(G1237));

  xor2  gate2143(.a(G1147), .b(G6), .O(gate429inter0));
  nand2 gate2144(.a(gate429inter0), .b(s_228), .O(gate429inter1));
  and2  gate2145(.a(G1147), .b(G6), .O(gate429inter2));
  inv1  gate2146(.a(s_228), .O(gate429inter3));
  inv1  gate2147(.a(s_229), .O(gate429inter4));
  nand2 gate2148(.a(gate429inter4), .b(gate429inter3), .O(gate429inter5));
  nor2  gate2149(.a(gate429inter5), .b(gate429inter2), .O(gate429inter6));
  inv1  gate2150(.a(G6), .O(gate429inter7));
  inv1  gate2151(.a(G1147), .O(gate429inter8));
  nand2 gate2152(.a(gate429inter8), .b(gate429inter7), .O(gate429inter9));
  nand2 gate2153(.a(s_229), .b(gate429inter3), .O(gate429inter10));
  nor2  gate2154(.a(gate429inter10), .b(gate429inter9), .O(gate429inter11));
  nor2  gate2155(.a(gate429inter11), .b(gate429inter6), .O(gate429inter12));
  nand2 gate2156(.a(gate429inter12), .b(gate429inter1), .O(G1238));
nand2 gate430( .a(G1051), .b(G1147), .O(G1239) );

  xor2  gate995(.a(G1150), .b(G7), .O(gate431inter0));
  nand2 gate996(.a(gate431inter0), .b(s_64), .O(gate431inter1));
  and2  gate997(.a(G1150), .b(G7), .O(gate431inter2));
  inv1  gate998(.a(s_64), .O(gate431inter3));
  inv1  gate999(.a(s_65), .O(gate431inter4));
  nand2 gate1000(.a(gate431inter4), .b(gate431inter3), .O(gate431inter5));
  nor2  gate1001(.a(gate431inter5), .b(gate431inter2), .O(gate431inter6));
  inv1  gate1002(.a(G7), .O(gate431inter7));
  inv1  gate1003(.a(G1150), .O(gate431inter8));
  nand2 gate1004(.a(gate431inter8), .b(gate431inter7), .O(gate431inter9));
  nand2 gate1005(.a(s_65), .b(gate431inter3), .O(gate431inter10));
  nor2  gate1006(.a(gate431inter10), .b(gate431inter9), .O(gate431inter11));
  nor2  gate1007(.a(gate431inter11), .b(gate431inter6), .O(gate431inter12));
  nand2 gate1008(.a(gate431inter12), .b(gate431inter1), .O(G1240));
nand2 gate432( .a(G1054), .b(G1150), .O(G1241) );
nand2 gate433( .a(G8), .b(G1153), .O(G1242) );
nand2 gate434( .a(G1057), .b(G1153), .O(G1243) );

  xor2  gate687(.a(G1156), .b(G9), .O(gate435inter0));
  nand2 gate688(.a(gate435inter0), .b(s_20), .O(gate435inter1));
  and2  gate689(.a(G1156), .b(G9), .O(gate435inter2));
  inv1  gate690(.a(s_20), .O(gate435inter3));
  inv1  gate691(.a(s_21), .O(gate435inter4));
  nand2 gate692(.a(gate435inter4), .b(gate435inter3), .O(gate435inter5));
  nor2  gate693(.a(gate435inter5), .b(gate435inter2), .O(gate435inter6));
  inv1  gate694(.a(G9), .O(gate435inter7));
  inv1  gate695(.a(G1156), .O(gate435inter8));
  nand2 gate696(.a(gate435inter8), .b(gate435inter7), .O(gate435inter9));
  nand2 gate697(.a(s_21), .b(gate435inter3), .O(gate435inter10));
  nor2  gate698(.a(gate435inter10), .b(gate435inter9), .O(gate435inter11));
  nor2  gate699(.a(gate435inter11), .b(gate435inter6), .O(gate435inter12));
  nand2 gate700(.a(gate435inter12), .b(gate435inter1), .O(G1244));

  xor2  gate939(.a(G1156), .b(G1060), .O(gate436inter0));
  nand2 gate940(.a(gate436inter0), .b(s_56), .O(gate436inter1));
  and2  gate941(.a(G1156), .b(G1060), .O(gate436inter2));
  inv1  gate942(.a(s_56), .O(gate436inter3));
  inv1  gate943(.a(s_57), .O(gate436inter4));
  nand2 gate944(.a(gate436inter4), .b(gate436inter3), .O(gate436inter5));
  nor2  gate945(.a(gate436inter5), .b(gate436inter2), .O(gate436inter6));
  inv1  gate946(.a(G1060), .O(gate436inter7));
  inv1  gate947(.a(G1156), .O(gate436inter8));
  nand2 gate948(.a(gate436inter8), .b(gate436inter7), .O(gate436inter9));
  nand2 gate949(.a(s_57), .b(gate436inter3), .O(gate436inter10));
  nor2  gate950(.a(gate436inter10), .b(gate436inter9), .O(gate436inter11));
  nor2  gate951(.a(gate436inter11), .b(gate436inter6), .O(gate436inter12));
  nand2 gate952(.a(gate436inter12), .b(gate436inter1), .O(G1245));
nand2 gate437( .a(G10), .b(G1159), .O(G1246) );
nand2 gate438( .a(G1063), .b(G1159), .O(G1247) );
nand2 gate439( .a(G11), .b(G1162), .O(G1248) );

  xor2  gate1541(.a(G1162), .b(G1066), .O(gate440inter0));
  nand2 gate1542(.a(gate440inter0), .b(s_142), .O(gate440inter1));
  and2  gate1543(.a(G1162), .b(G1066), .O(gate440inter2));
  inv1  gate1544(.a(s_142), .O(gate440inter3));
  inv1  gate1545(.a(s_143), .O(gate440inter4));
  nand2 gate1546(.a(gate440inter4), .b(gate440inter3), .O(gate440inter5));
  nor2  gate1547(.a(gate440inter5), .b(gate440inter2), .O(gate440inter6));
  inv1  gate1548(.a(G1066), .O(gate440inter7));
  inv1  gate1549(.a(G1162), .O(gate440inter8));
  nand2 gate1550(.a(gate440inter8), .b(gate440inter7), .O(gate440inter9));
  nand2 gate1551(.a(s_143), .b(gate440inter3), .O(gate440inter10));
  nor2  gate1552(.a(gate440inter10), .b(gate440inter9), .O(gate440inter11));
  nor2  gate1553(.a(gate440inter11), .b(gate440inter6), .O(gate440inter12));
  nand2 gate1554(.a(gate440inter12), .b(gate440inter1), .O(G1249));
nand2 gate441( .a(G12), .b(G1165), .O(G1250) );
nand2 gate442( .a(G1069), .b(G1165), .O(G1251) );
nand2 gate443( .a(G13), .b(G1168), .O(G1252) );

  xor2  gate1065(.a(G1168), .b(G1072), .O(gate444inter0));
  nand2 gate1066(.a(gate444inter0), .b(s_74), .O(gate444inter1));
  and2  gate1067(.a(G1168), .b(G1072), .O(gate444inter2));
  inv1  gate1068(.a(s_74), .O(gate444inter3));
  inv1  gate1069(.a(s_75), .O(gate444inter4));
  nand2 gate1070(.a(gate444inter4), .b(gate444inter3), .O(gate444inter5));
  nor2  gate1071(.a(gate444inter5), .b(gate444inter2), .O(gate444inter6));
  inv1  gate1072(.a(G1072), .O(gate444inter7));
  inv1  gate1073(.a(G1168), .O(gate444inter8));
  nand2 gate1074(.a(gate444inter8), .b(gate444inter7), .O(gate444inter9));
  nand2 gate1075(.a(s_75), .b(gate444inter3), .O(gate444inter10));
  nor2  gate1076(.a(gate444inter10), .b(gate444inter9), .O(gate444inter11));
  nor2  gate1077(.a(gate444inter11), .b(gate444inter6), .O(gate444inter12));
  nand2 gate1078(.a(gate444inter12), .b(gate444inter1), .O(G1253));

  xor2  gate673(.a(G1171), .b(G14), .O(gate445inter0));
  nand2 gate674(.a(gate445inter0), .b(s_18), .O(gate445inter1));
  and2  gate675(.a(G1171), .b(G14), .O(gate445inter2));
  inv1  gate676(.a(s_18), .O(gate445inter3));
  inv1  gate677(.a(s_19), .O(gate445inter4));
  nand2 gate678(.a(gate445inter4), .b(gate445inter3), .O(gate445inter5));
  nor2  gate679(.a(gate445inter5), .b(gate445inter2), .O(gate445inter6));
  inv1  gate680(.a(G14), .O(gate445inter7));
  inv1  gate681(.a(G1171), .O(gate445inter8));
  nand2 gate682(.a(gate445inter8), .b(gate445inter7), .O(gate445inter9));
  nand2 gate683(.a(s_19), .b(gate445inter3), .O(gate445inter10));
  nor2  gate684(.a(gate445inter10), .b(gate445inter9), .O(gate445inter11));
  nor2  gate685(.a(gate445inter11), .b(gate445inter6), .O(gate445inter12));
  nand2 gate686(.a(gate445inter12), .b(gate445inter1), .O(G1254));
nand2 gate446( .a(G1075), .b(G1171), .O(G1255) );

  xor2  gate575(.a(G1174), .b(G15), .O(gate447inter0));
  nand2 gate576(.a(gate447inter0), .b(s_4), .O(gate447inter1));
  and2  gate577(.a(G1174), .b(G15), .O(gate447inter2));
  inv1  gate578(.a(s_4), .O(gate447inter3));
  inv1  gate579(.a(s_5), .O(gate447inter4));
  nand2 gate580(.a(gate447inter4), .b(gate447inter3), .O(gate447inter5));
  nor2  gate581(.a(gate447inter5), .b(gate447inter2), .O(gate447inter6));
  inv1  gate582(.a(G15), .O(gate447inter7));
  inv1  gate583(.a(G1174), .O(gate447inter8));
  nand2 gate584(.a(gate447inter8), .b(gate447inter7), .O(gate447inter9));
  nand2 gate585(.a(s_5), .b(gate447inter3), .O(gate447inter10));
  nor2  gate586(.a(gate447inter10), .b(gate447inter9), .O(gate447inter11));
  nor2  gate587(.a(gate447inter11), .b(gate447inter6), .O(gate447inter12));
  nand2 gate588(.a(gate447inter12), .b(gate447inter1), .O(G1256));
nand2 gate448( .a(G1078), .b(G1174), .O(G1257) );
nand2 gate449( .a(G16), .b(G1177), .O(G1258) );

  xor2  gate1975(.a(G1177), .b(G1081), .O(gate450inter0));
  nand2 gate1976(.a(gate450inter0), .b(s_204), .O(gate450inter1));
  and2  gate1977(.a(G1177), .b(G1081), .O(gate450inter2));
  inv1  gate1978(.a(s_204), .O(gate450inter3));
  inv1  gate1979(.a(s_205), .O(gate450inter4));
  nand2 gate1980(.a(gate450inter4), .b(gate450inter3), .O(gate450inter5));
  nor2  gate1981(.a(gate450inter5), .b(gate450inter2), .O(gate450inter6));
  inv1  gate1982(.a(G1081), .O(gate450inter7));
  inv1  gate1983(.a(G1177), .O(gate450inter8));
  nand2 gate1984(.a(gate450inter8), .b(gate450inter7), .O(gate450inter9));
  nand2 gate1985(.a(s_205), .b(gate450inter3), .O(gate450inter10));
  nor2  gate1986(.a(gate450inter10), .b(gate450inter9), .O(gate450inter11));
  nor2  gate1987(.a(gate450inter11), .b(gate450inter6), .O(gate450inter12));
  nand2 gate1988(.a(gate450inter12), .b(gate450inter1), .O(G1259));

  xor2  gate2031(.a(G1180), .b(G17), .O(gate451inter0));
  nand2 gate2032(.a(gate451inter0), .b(s_212), .O(gate451inter1));
  and2  gate2033(.a(G1180), .b(G17), .O(gate451inter2));
  inv1  gate2034(.a(s_212), .O(gate451inter3));
  inv1  gate2035(.a(s_213), .O(gate451inter4));
  nand2 gate2036(.a(gate451inter4), .b(gate451inter3), .O(gate451inter5));
  nor2  gate2037(.a(gate451inter5), .b(gate451inter2), .O(gate451inter6));
  inv1  gate2038(.a(G17), .O(gate451inter7));
  inv1  gate2039(.a(G1180), .O(gate451inter8));
  nand2 gate2040(.a(gate451inter8), .b(gate451inter7), .O(gate451inter9));
  nand2 gate2041(.a(s_213), .b(gate451inter3), .O(gate451inter10));
  nor2  gate2042(.a(gate451inter10), .b(gate451inter9), .O(gate451inter11));
  nor2  gate2043(.a(gate451inter11), .b(gate451inter6), .O(gate451inter12));
  nand2 gate2044(.a(gate451inter12), .b(gate451inter1), .O(G1260));

  xor2  gate1513(.a(G1180), .b(G1084), .O(gate452inter0));
  nand2 gate1514(.a(gate452inter0), .b(s_138), .O(gate452inter1));
  and2  gate1515(.a(G1180), .b(G1084), .O(gate452inter2));
  inv1  gate1516(.a(s_138), .O(gate452inter3));
  inv1  gate1517(.a(s_139), .O(gate452inter4));
  nand2 gate1518(.a(gate452inter4), .b(gate452inter3), .O(gate452inter5));
  nor2  gate1519(.a(gate452inter5), .b(gate452inter2), .O(gate452inter6));
  inv1  gate1520(.a(G1084), .O(gate452inter7));
  inv1  gate1521(.a(G1180), .O(gate452inter8));
  nand2 gate1522(.a(gate452inter8), .b(gate452inter7), .O(gate452inter9));
  nand2 gate1523(.a(s_139), .b(gate452inter3), .O(gate452inter10));
  nor2  gate1524(.a(gate452inter10), .b(gate452inter9), .O(gate452inter11));
  nor2  gate1525(.a(gate452inter11), .b(gate452inter6), .O(gate452inter12));
  nand2 gate1526(.a(gate452inter12), .b(gate452inter1), .O(G1261));
nand2 gate453( .a(G18), .b(G1183), .O(G1262) );

  xor2  gate1037(.a(G1183), .b(G1087), .O(gate454inter0));
  nand2 gate1038(.a(gate454inter0), .b(s_70), .O(gate454inter1));
  and2  gate1039(.a(G1183), .b(G1087), .O(gate454inter2));
  inv1  gate1040(.a(s_70), .O(gate454inter3));
  inv1  gate1041(.a(s_71), .O(gate454inter4));
  nand2 gate1042(.a(gate454inter4), .b(gate454inter3), .O(gate454inter5));
  nor2  gate1043(.a(gate454inter5), .b(gate454inter2), .O(gate454inter6));
  inv1  gate1044(.a(G1087), .O(gate454inter7));
  inv1  gate1045(.a(G1183), .O(gate454inter8));
  nand2 gate1046(.a(gate454inter8), .b(gate454inter7), .O(gate454inter9));
  nand2 gate1047(.a(s_71), .b(gate454inter3), .O(gate454inter10));
  nor2  gate1048(.a(gate454inter10), .b(gate454inter9), .O(gate454inter11));
  nor2  gate1049(.a(gate454inter11), .b(gate454inter6), .O(gate454inter12));
  nand2 gate1050(.a(gate454inter12), .b(gate454inter1), .O(G1263));
nand2 gate455( .a(G19), .b(G1186), .O(G1264) );
nand2 gate456( .a(G1090), .b(G1186), .O(G1265) );
nand2 gate457( .a(G20), .b(G1189), .O(G1266) );
nand2 gate458( .a(G1093), .b(G1189), .O(G1267) );

  xor2  gate2129(.a(G1192), .b(G21), .O(gate459inter0));
  nand2 gate2130(.a(gate459inter0), .b(s_226), .O(gate459inter1));
  and2  gate2131(.a(G1192), .b(G21), .O(gate459inter2));
  inv1  gate2132(.a(s_226), .O(gate459inter3));
  inv1  gate2133(.a(s_227), .O(gate459inter4));
  nand2 gate2134(.a(gate459inter4), .b(gate459inter3), .O(gate459inter5));
  nor2  gate2135(.a(gate459inter5), .b(gate459inter2), .O(gate459inter6));
  inv1  gate2136(.a(G21), .O(gate459inter7));
  inv1  gate2137(.a(G1192), .O(gate459inter8));
  nand2 gate2138(.a(gate459inter8), .b(gate459inter7), .O(gate459inter9));
  nand2 gate2139(.a(s_227), .b(gate459inter3), .O(gate459inter10));
  nor2  gate2140(.a(gate459inter10), .b(gate459inter9), .O(gate459inter11));
  nor2  gate2141(.a(gate459inter11), .b(gate459inter6), .O(gate459inter12));
  nand2 gate2142(.a(gate459inter12), .b(gate459inter1), .O(G1268));
nand2 gate460( .a(G1096), .b(G1192), .O(G1269) );
nand2 gate461( .a(G22), .b(G1195), .O(G1270) );
nand2 gate462( .a(G1099), .b(G1195), .O(G1271) );
nand2 gate463( .a(G23), .b(G1198), .O(G1272) );

  xor2  gate617(.a(G1198), .b(G1102), .O(gate464inter0));
  nand2 gate618(.a(gate464inter0), .b(s_10), .O(gate464inter1));
  and2  gate619(.a(G1198), .b(G1102), .O(gate464inter2));
  inv1  gate620(.a(s_10), .O(gate464inter3));
  inv1  gate621(.a(s_11), .O(gate464inter4));
  nand2 gate622(.a(gate464inter4), .b(gate464inter3), .O(gate464inter5));
  nor2  gate623(.a(gate464inter5), .b(gate464inter2), .O(gate464inter6));
  inv1  gate624(.a(G1102), .O(gate464inter7));
  inv1  gate625(.a(G1198), .O(gate464inter8));
  nand2 gate626(.a(gate464inter8), .b(gate464inter7), .O(gate464inter9));
  nand2 gate627(.a(s_11), .b(gate464inter3), .O(gate464inter10));
  nor2  gate628(.a(gate464inter10), .b(gate464inter9), .O(gate464inter11));
  nor2  gate629(.a(gate464inter11), .b(gate464inter6), .O(gate464inter12));
  nand2 gate630(.a(gate464inter12), .b(gate464inter1), .O(G1273));
nand2 gate465( .a(G24), .b(G1201), .O(G1274) );
nand2 gate466( .a(G1105), .b(G1201), .O(G1275) );

  xor2  gate1317(.a(G1204), .b(G25), .O(gate467inter0));
  nand2 gate1318(.a(gate467inter0), .b(s_110), .O(gate467inter1));
  and2  gate1319(.a(G1204), .b(G25), .O(gate467inter2));
  inv1  gate1320(.a(s_110), .O(gate467inter3));
  inv1  gate1321(.a(s_111), .O(gate467inter4));
  nand2 gate1322(.a(gate467inter4), .b(gate467inter3), .O(gate467inter5));
  nor2  gate1323(.a(gate467inter5), .b(gate467inter2), .O(gate467inter6));
  inv1  gate1324(.a(G25), .O(gate467inter7));
  inv1  gate1325(.a(G1204), .O(gate467inter8));
  nand2 gate1326(.a(gate467inter8), .b(gate467inter7), .O(gate467inter9));
  nand2 gate1327(.a(s_111), .b(gate467inter3), .O(gate467inter10));
  nor2  gate1328(.a(gate467inter10), .b(gate467inter9), .O(gate467inter11));
  nor2  gate1329(.a(gate467inter11), .b(gate467inter6), .O(gate467inter12));
  nand2 gate1330(.a(gate467inter12), .b(gate467inter1), .O(G1276));
nand2 gate468( .a(G1108), .b(G1204), .O(G1277) );

  xor2  gate1415(.a(G1207), .b(G26), .O(gate469inter0));
  nand2 gate1416(.a(gate469inter0), .b(s_124), .O(gate469inter1));
  and2  gate1417(.a(G1207), .b(G26), .O(gate469inter2));
  inv1  gate1418(.a(s_124), .O(gate469inter3));
  inv1  gate1419(.a(s_125), .O(gate469inter4));
  nand2 gate1420(.a(gate469inter4), .b(gate469inter3), .O(gate469inter5));
  nor2  gate1421(.a(gate469inter5), .b(gate469inter2), .O(gate469inter6));
  inv1  gate1422(.a(G26), .O(gate469inter7));
  inv1  gate1423(.a(G1207), .O(gate469inter8));
  nand2 gate1424(.a(gate469inter8), .b(gate469inter7), .O(gate469inter9));
  nand2 gate1425(.a(s_125), .b(gate469inter3), .O(gate469inter10));
  nor2  gate1426(.a(gate469inter10), .b(gate469inter9), .O(gate469inter11));
  nor2  gate1427(.a(gate469inter11), .b(gate469inter6), .O(gate469inter12));
  nand2 gate1428(.a(gate469inter12), .b(gate469inter1), .O(G1278));
nand2 gate470( .a(G1111), .b(G1207), .O(G1279) );
nand2 gate471( .a(G27), .b(G1210), .O(G1280) );
nand2 gate472( .a(G1114), .b(G1210), .O(G1281) );
nand2 gate473( .a(G28), .b(G1213), .O(G1282) );

  xor2  gate1611(.a(G1213), .b(G1117), .O(gate474inter0));
  nand2 gate1612(.a(gate474inter0), .b(s_152), .O(gate474inter1));
  and2  gate1613(.a(G1213), .b(G1117), .O(gate474inter2));
  inv1  gate1614(.a(s_152), .O(gate474inter3));
  inv1  gate1615(.a(s_153), .O(gate474inter4));
  nand2 gate1616(.a(gate474inter4), .b(gate474inter3), .O(gate474inter5));
  nor2  gate1617(.a(gate474inter5), .b(gate474inter2), .O(gate474inter6));
  inv1  gate1618(.a(G1117), .O(gate474inter7));
  inv1  gate1619(.a(G1213), .O(gate474inter8));
  nand2 gate1620(.a(gate474inter8), .b(gate474inter7), .O(gate474inter9));
  nand2 gate1621(.a(s_153), .b(gate474inter3), .O(gate474inter10));
  nor2  gate1622(.a(gate474inter10), .b(gate474inter9), .O(gate474inter11));
  nor2  gate1623(.a(gate474inter11), .b(gate474inter6), .O(gate474inter12));
  nand2 gate1624(.a(gate474inter12), .b(gate474inter1), .O(G1283));

  xor2  gate1583(.a(G1216), .b(G29), .O(gate475inter0));
  nand2 gate1584(.a(gate475inter0), .b(s_148), .O(gate475inter1));
  and2  gate1585(.a(G1216), .b(G29), .O(gate475inter2));
  inv1  gate1586(.a(s_148), .O(gate475inter3));
  inv1  gate1587(.a(s_149), .O(gate475inter4));
  nand2 gate1588(.a(gate475inter4), .b(gate475inter3), .O(gate475inter5));
  nor2  gate1589(.a(gate475inter5), .b(gate475inter2), .O(gate475inter6));
  inv1  gate1590(.a(G29), .O(gate475inter7));
  inv1  gate1591(.a(G1216), .O(gate475inter8));
  nand2 gate1592(.a(gate475inter8), .b(gate475inter7), .O(gate475inter9));
  nand2 gate1593(.a(s_149), .b(gate475inter3), .O(gate475inter10));
  nor2  gate1594(.a(gate475inter10), .b(gate475inter9), .O(gate475inter11));
  nor2  gate1595(.a(gate475inter11), .b(gate475inter6), .O(gate475inter12));
  nand2 gate1596(.a(gate475inter12), .b(gate475inter1), .O(G1284));
nand2 gate476( .a(G1120), .b(G1216), .O(G1285) );
nand2 gate477( .a(G30), .b(G1219), .O(G1286) );
nand2 gate478( .a(G1123), .b(G1219), .O(G1287) );
nand2 gate479( .a(G31), .b(G1222), .O(G1288) );
nand2 gate480( .a(G1126), .b(G1222), .O(G1289) );
nand2 gate481( .a(G32), .b(G1225), .O(G1290) );
nand2 gate482( .a(G1129), .b(G1225), .O(G1291) );
nand2 gate483( .a(G1228), .b(G1229), .O(G1292) );
nand2 gate484( .a(G1230), .b(G1231), .O(G1293) );
nand2 gate485( .a(G1232), .b(G1233), .O(G1294) );

  xor2  gate967(.a(G1235), .b(G1234), .O(gate486inter0));
  nand2 gate968(.a(gate486inter0), .b(s_60), .O(gate486inter1));
  and2  gate969(.a(G1235), .b(G1234), .O(gate486inter2));
  inv1  gate970(.a(s_60), .O(gate486inter3));
  inv1  gate971(.a(s_61), .O(gate486inter4));
  nand2 gate972(.a(gate486inter4), .b(gate486inter3), .O(gate486inter5));
  nor2  gate973(.a(gate486inter5), .b(gate486inter2), .O(gate486inter6));
  inv1  gate974(.a(G1234), .O(gate486inter7));
  inv1  gate975(.a(G1235), .O(gate486inter8));
  nand2 gate976(.a(gate486inter8), .b(gate486inter7), .O(gate486inter9));
  nand2 gate977(.a(s_61), .b(gate486inter3), .O(gate486inter10));
  nor2  gate978(.a(gate486inter10), .b(gate486inter9), .O(gate486inter11));
  nor2  gate979(.a(gate486inter11), .b(gate486inter6), .O(gate486inter12));
  nand2 gate980(.a(gate486inter12), .b(gate486inter1), .O(G1295));
nand2 gate487( .a(G1236), .b(G1237), .O(G1296) );
nand2 gate488( .a(G1238), .b(G1239), .O(G1297) );
nand2 gate489( .a(G1240), .b(G1241), .O(G1298) );
nand2 gate490( .a(G1242), .b(G1243), .O(G1299) );
nand2 gate491( .a(G1244), .b(G1245), .O(G1300) );
nand2 gate492( .a(G1246), .b(G1247), .O(G1301) );
nand2 gate493( .a(G1248), .b(G1249), .O(G1302) );

  xor2  gate645(.a(G1251), .b(G1250), .O(gate494inter0));
  nand2 gate646(.a(gate494inter0), .b(s_14), .O(gate494inter1));
  and2  gate647(.a(G1251), .b(G1250), .O(gate494inter2));
  inv1  gate648(.a(s_14), .O(gate494inter3));
  inv1  gate649(.a(s_15), .O(gate494inter4));
  nand2 gate650(.a(gate494inter4), .b(gate494inter3), .O(gate494inter5));
  nor2  gate651(.a(gate494inter5), .b(gate494inter2), .O(gate494inter6));
  inv1  gate652(.a(G1250), .O(gate494inter7));
  inv1  gate653(.a(G1251), .O(gate494inter8));
  nand2 gate654(.a(gate494inter8), .b(gate494inter7), .O(gate494inter9));
  nand2 gate655(.a(s_15), .b(gate494inter3), .O(gate494inter10));
  nor2  gate656(.a(gate494inter10), .b(gate494inter9), .O(gate494inter11));
  nor2  gate657(.a(gate494inter11), .b(gate494inter6), .O(gate494inter12));
  nand2 gate658(.a(gate494inter12), .b(gate494inter1), .O(G1303));
nand2 gate495( .a(G1252), .b(G1253), .O(G1304) );
nand2 gate496( .a(G1254), .b(G1255), .O(G1305) );
nand2 gate497( .a(G1256), .b(G1257), .O(G1306) );

  xor2  gate1219(.a(G1259), .b(G1258), .O(gate498inter0));
  nand2 gate1220(.a(gate498inter0), .b(s_96), .O(gate498inter1));
  and2  gate1221(.a(G1259), .b(G1258), .O(gate498inter2));
  inv1  gate1222(.a(s_96), .O(gate498inter3));
  inv1  gate1223(.a(s_97), .O(gate498inter4));
  nand2 gate1224(.a(gate498inter4), .b(gate498inter3), .O(gate498inter5));
  nor2  gate1225(.a(gate498inter5), .b(gate498inter2), .O(gate498inter6));
  inv1  gate1226(.a(G1258), .O(gate498inter7));
  inv1  gate1227(.a(G1259), .O(gate498inter8));
  nand2 gate1228(.a(gate498inter8), .b(gate498inter7), .O(gate498inter9));
  nand2 gate1229(.a(s_97), .b(gate498inter3), .O(gate498inter10));
  nor2  gate1230(.a(gate498inter10), .b(gate498inter9), .O(gate498inter11));
  nor2  gate1231(.a(gate498inter11), .b(gate498inter6), .O(gate498inter12));
  nand2 gate1232(.a(gate498inter12), .b(gate498inter1), .O(G1307));

  xor2  gate911(.a(G1261), .b(G1260), .O(gate499inter0));
  nand2 gate912(.a(gate499inter0), .b(s_52), .O(gate499inter1));
  and2  gate913(.a(G1261), .b(G1260), .O(gate499inter2));
  inv1  gate914(.a(s_52), .O(gate499inter3));
  inv1  gate915(.a(s_53), .O(gate499inter4));
  nand2 gate916(.a(gate499inter4), .b(gate499inter3), .O(gate499inter5));
  nor2  gate917(.a(gate499inter5), .b(gate499inter2), .O(gate499inter6));
  inv1  gate918(.a(G1260), .O(gate499inter7));
  inv1  gate919(.a(G1261), .O(gate499inter8));
  nand2 gate920(.a(gate499inter8), .b(gate499inter7), .O(gate499inter9));
  nand2 gate921(.a(s_53), .b(gate499inter3), .O(gate499inter10));
  nor2  gate922(.a(gate499inter10), .b(gate499inter9), .O(gate499inter11));
  nor2  gate923(.a(gate499inter11), .b(gate499inter6), .O(gate499inter12));
  nand2 gate924(.a(gate499inter12), .b(gate499inter1), .O(G1308));
nand2 gate500( .a(G1262), .b(G1263), .O(G1309) );
nand2 gate501( .a(G1264), .b(G1265), .O(G1310) );

  xor2  gate1051(.a(G1267), .b(G1266), .O(gate502inter0));
  nand2 gate1052(.a(gate502inter0), .b(s_72), .O(gate502inter1));
  and2  gate1053(.a(G1267), .b(G1266), .O(gate502inter2));
  inv1  gate1054(.a(s_72), .O(gate502inter3));
  inv1  gate1055(.a(s_73), .O(gate502inter4));
  nand2 gate1056(.a(gate502inter4), .b(gate502inter3), .O(gate502inter5));
  nor2  gate1057(.a(gate502inter5), .b(gate502inter2), .O(gate502inter6));
  inv1  gate1058(.a(G1266), .O(gate502inter7));
  inv1  gate1059(.a(G1267), .O(gate502inter8));
  nand2 gate1060(.a(gate502inter8), .b(gate502inter7), .O(gate502inter9));
  nand2 gate1061(.a(s_73), .b(gate502inter3), .O(gate502inter10));
  nor2  gate1062(.a(gate502inter10), .b(gate502inter9), .O(gate502inter11));
  nor2  gate1063(.a(gate502inter11), .b(gate502inter6), .O(gate502inter12));
  nand2 gate1064(.a(gate502inter12), .b(gate502inter1), .O(G1311));
nand2 gate503( .a(G1268), .b(G1269), .O(G1312) );

  xor2  gate981(.a(G1271), .b(G1270), .O(gate504inter0));
  nand2 gate982(.a(gate504inter0), .b(s_62), .O(gate504inter1));
  and2  gate983(.a(G1271), .b(G1270), .O(gate504inter2));
  inv1  gate984(.a(s_62), .O(gate504inter3));
  inv1  gate985(.a(s_63), .O(gate504inter4));
  nand2 gate986(.a(gate504inter4), .b(gate504inter3), .O(gate504inter5));
  nor2  gate987(.a(gate504inter5), .b(gate504inter2), .O(gate504inter6));
  inv1  gate988(.a(G1270), .O(gate504inter7));
  inv1  gate989(.a(G1271), .O(gate504inter8));
  nand2 gate990(.a(gate504inter8), .b(gate504inter7), .O(gate504inter9));
  nand2 gate991(.a(s_63), .b(gate504inter3), .O(gate504inter10));
  nor2  gate992(.a(gate504inter10), .b(gate504inter9), .O(gate504inter11));
  nor2  gate993(.a(gate504inter11), .b(gate504inter6), .O(gate504inter12));
  nand2 gate994(.a(gate504inter12), .b(gate504inter1), .O(G1313));
nand2 gate505( .a(G1272), .b(G1273), .O(G1314) );
nand2 gate506( .a(G1274), .b(G1275), .O(G1315) );
nand2 gate507( .a(G1276), .b(G1277), .O(G1316) );
nand2 gate508( .a(G1278), .b(G1279), .O(G1317) );
nand2 gate509( .a(G1280), .b(G1281), .O(G1318) );
nand2 gate510( .a(G1282), .b(G1283), .O(G1319) );
nand2 gate511( .a(G1284), .b(G1285), .O(G1320) );
nand2 gate512( .a(G1286), .b(G1287), .O(G1321) );
nand2 gate513( .a(G1288), .b(G1289), .O(G1322) );

  xor2  gate1331(.a(G1291), .b(G1290), .O(gate514inter0));
  nand2 gate1332(.a(gate514inter0), .b(s_112), .O(gate514inter1));
  and2  gate1333(.a(G1291), .b(G1290), .O(gate514inter2));
  inv1  gate1334(.a(s_112), .O(gate514inter3));
  inv1  gate1335(.a(s_113), .O(gate514inter4));
  nand2 gate1336(.a(gate514inter4), .b(gate514inter3), .O(gate514inter5));
  nor2  gate1337(.a(gate514inter5), .b(gate514inter2), .O(gate514inter6));
  inv1  gate1338(.a(G1290), .O(gate514inter7));
  inv1  gate1339(.a(G1291), .O(gate514inter8));
  nand2 gate1340(.a(gate514inter8), .b(gate514inter7), .O(gate514inter9));
  nand2 gate1341(.a(s_113), .b(gate514inter3), .O(gate514inter10));
  nor2  gate1342(.a(gate514inter10), .b(gate514inter9), .O(gate514inter11));
  nor2  gate1343(.a(gate514inter11), .b(gate514inter6), .O(gate514inter12));
  nand2 gate1344(.a(gate514inter12), .b(gate514inter1), .O(G1323));
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule