module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);

input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;//RE__PI;

input s_0,s_1;//RE__ALLOW(00,01,10,11);
input s_2,s_3;//RE__ALLOW(00,01,10,11);
input s_4,s_5;//RE__ALLOW(00,01,10,11);
input s_6,s_7;//RE__ALLOW(00,01,10,11);
input s_8,s_9;//RE__ALLOW(00,01,10,11);
input s_10,s_11;//RE__ALLOW(00,01,10,11);
input s_12,s_13;//RE__ALLOW(00,01,10,11);
input s_14,s_15;//RE__ALLOW(00,01,10,11);
input s_16,s_17;//RE__ALLOW(00,01,10,11);
input s_18,s_19;//RE__ALLOW(00,01,10,11);
input s_20,s_21;//RE__ALLOW(00,01,10,11);
input s_22,s_23;//RE__ALLOW(00,01,10,11);
input s_24,s_25;//RE__ALLOW(00,01,10,11);
input s_26,s_27;//RE__ALLOW(00,01,10,11);
input s_28,s_29;//RE__ALLOW(00,01,10,11);
input s_30,s_31;//RE__ALLOW(00,01,10,11);
input s_32,s_33;//RE__ALLOW(00,01,10,11);
input s_34,s_35;//RE__ALLOW(00,01,10,11);
input s_36,s_37;//RE__ALLOW(00,01,10,11);
input s_38,s_39;//RE__ALLOW(00,01,10,11);
input s_40,s_41;//RE__ALLOW(00,01,10,11);
input s_42,s_43;//RE__ALLOW(00,01,10,11);
input s_44,s_45;//RE__ALLOW(00,01,10,11);
input s_46,s_47;//RE__ALLOW(00,01,10,11);
input s_48,s_49;//RE__ALLOW(00,01,10,11);
input s_50,s_51;//RE__ALLOW(00,01,10,11);
input s_52,s_53;//RE__ALLOW(00,01,10,11);
input s_54,s_55;//RE__ALLOW(00,01,10,11);
input s_56,s_57;//RE__ALLOW(00,01,10,11);
input s_58,s_59;//RE__ALLOW(00,01,10,11);
input s_60,s_61;//RE__ALLOW(00,01,10,11);
input s_62,s_63;//RE__ALLOW(00,01,10,11);
input s_64,s_65;//RE__ALLOW(00,01,10,11);
input s_66,s_67;//RE__ALLOW(00,01,10,11);
input s_68,s_69;//RE__ALLOW(00,01,10,11);
input s_70,s_71;//RE__ALLOW(00,01,10,11);
input s_72,s_73;//RE__ALLOW(00,01,10,11);
input s_74,s_75;//RE__ALLOW(00,01,10,11);
input s_76,s_77;//RE__ALLOW(00,01,10,11);
input s_78,s_79;//RE__ALLOW(00,01,10,11);
input s_80,s_81;//RE__ALLOW(00,01,10,11);
input s_82,s_83;//RE__ALLOW(00,01,10,11);
input s_84,s_85;//RE__ALLOW(00,01,10,11);
input s_86,s_87;//RE__ALLOW(00,01,10,11);
input s_88,s_89;//RE__ALLOW(00,01,10,11);
input s_90,s_91;//RE__ALLOW(00,01,10,11);
input s_92,s_93;//RE__ALLOW(00,01,10,11);
input s_94,s_95;//RE__ALLOW(00,01,10,11);
input s_96,s_97;//RE__ALLOW(00,01,10,11);
input s_98,s_99;//RE__ALLOW(00,01,10,11);
input s_100,s_101;//RE__ALLOW(00,01,10,11);
input s_102,s_103;//RE__ALLOW(00,01,10,11);
input s_104,s_105;//RE__ALLOW(00,01,10,11);
input s_106,s_107;//RE__ALLOW(00,01,10,11);
input s_108,s_109;//RE__ALLOW(00,01,10,11);
input s_110,s_111;//RE__ALLOW(00,01,10,11);
input s_112,s_113;//RE__ALLOW(00,01,10,11);
input s_114,s_115;//RE__ALLOW(00,01,10,11);
input s_116,s_117;//RE__ALLOW(00,01,10,11);
input s_118,s_119;//RE__ALLOW(00,01,10,11);
input s_120,s_121;//RE__ALLOW(00,01,10,11);
input s_122,s_123;//RE__ALLOW(00,01,10,11);
input s_124,s_125;//RE__ALLOW(00,01,10,11);
input s_126,s_127;//RE__ALLOW(00,01,10,11);
input s_128,s_129;//RE__ALLOW(00,01,10,11);
input s_130,s_131;//RE__ALLOW(00,01,10,11);
input s_132,s_133;//RE__ALLOW(00,01,10,11);
input s_134,s_135;//RE__ALLOW(00,01,10,11);
input s_136,s_137;//RE__ALLOW(00,01,10,11);
input s_138,s_139;//RE__ALLOW(00,01,10,11);
input s_140,s_141;//RE__ALLOW(00,01,10,11);
input s_142,s_143;//RE__ALLOW(00,01,10,11);
input s_144,s_145;//RE__ALLOW(00,01,10,11);
input s_146,s_147;//RE__ALLOW(00,01,10,11);
input s_148,s_149;//RE__ALLOW(00,01,10,11);
input s_150,s_151;//RE__ALLOW(00,01,10,11);
input s_152,s_153;//RE__ALLOW(00,01,10,11);
input s_154,s_155;//RE__ALLOW(00,01,10,11);
input s_156,s_157;//RE__ALLOW(00,01,10,11);
input s_158,s_159;//RE__ALLOW(00,01,10,11);
input s_160,s_161;//RE__ALLOW(00,01,10,11);
input s_162,s_163;//RE__ALLOW(00,01,10,11);
input s_164,s_165;//RE__ALLOW(00,01,10,11);
input s_166,s_167;//RE__ALLOW(00,01,10,11);
input s_168,s_169;//RE__ALLOW(00,01,10,11);
input s_170,s_171;//RE__ALLOW(00,01,10,11);
input s_172,s_173;//RE__ALLOW(00,01,10,11);
input s_174,s_175;//RE__ALLOW(00,01,10,11);
input s_176,s_177;//RE__ALLOW(00,01,10,11);
input s_178,s_179;//RE__ALLOW(00,01,10,11);
input s_180,s_181;//RE__ALLOW(00,01,10,11);
input s_182,s_183;//RE__ALLOW(00,01,10,11);
input s_184,s_185;//RE__ALLOW(00,01,10,11);
input s_186,s_187;//RE__ALLOW(00,01,10,11);
input s_188,s_189;//RE__ALLOW(00,01,10,11);
input s_190,s_191;//RE__ALLOW(00,01,10,11);
input s_192,s_193;//RE__ALLOW(00,01,10,11);
input s_194,s_195;//RE__ALLOW(00,01,10,11);
input s_196,s_197;//RE__ALLOW(00,01,10,11);
input s_198,s_199;//RE__ALLOW(00,01,10,11);
input s_200,s_201;//RE__ALLOW(00,01,10,11);
input s_202,s_203;//RE__ALLOW(00,01,10,11);
input s_204,s_205;//RE__ALLOW(00,01,10,11);
input s_206,s_207;//RE__ALLOW(00,01,10,11);
input s_208,s_209;//RE__ALLOW(00,01,10,11);
input s_210,s_211;//RE__ALLOW(00,01,10,11);
input s_212,s_213;//RE__ALLOW(00,01,10,11);
input s_214,s_215;//RE__ALLOW(00,01,10,11);
input s_216,s_217;//RE__ALLOW(00,01,10,11);
input s_218,s_219;//RE__ALLOW(00,01,10,11);
input s_220,s_221;//RE__ALLOW(00,01,10,11);
input s_222,s_223;//RE__ALLOW(00,01,10,11);
input s_224,s_225;//RE__ALLOW(00,01,10,11);
input s_226,s_227;//RE__ALLOW(00,01,10,11);
input s_228,s_229;//RE__ALLOW(00,01,10,11);
input s_230,s_231;//RE__ALLOW(00,01,10,11);
input s_232,s_233;//RE__ALLOW(00,01,10,11);
input s_234,s_235;//RE__ALLOW(00,01,10,11);
input s_236,s_237;//RE__ALLOW(00,01,10,11);
input s_238,s_239;//RE__ALLOW(00,01,10,11);
input s_240,s_241;//RE__ALLOW(00,01,10,11);
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;

  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate471inter0, gate471inter1, gate471inter2, gate471inter3, gate471inter4, gate471inter5, gate471inter6, gate471inter7, gate471inter8, gate471inter9, gate471inter10, gate471inter11, gate471inter12, gate231inter0, gate231inter1, gate231inter2, gate231inter3, gate231inter4, gate231inter5, gate231inter6, gate231inter7, gate231inter8, gate231inter9, gate231inter10, gate231inter11, gate231inter12, gate270inter0, gate270inter1, gate270inter2, gate270inter3, gate270inter4, gate270inter5, gate270inter6, gate270inter7, gate270inter8, gate270inter9, gate270inter10, gate270inter11, gate270inter12, gate26inter0, gate26inter1, gate26inter2, gate26inter3, gate26inter4, gate26inter5, gate26inter6, gate26inter7, gate26inter8, gate26inter9, gate26inter10, gate26inter11, gate26inter12, gate160inter0, gate160inter1, gate160inter2, gate160inter3, gate160inter4, gate160inter5, gate160inter6, gate160inter7, gate160inter8, gate160inter9, gate160inter10, gate160inter11, gate160inter12, gate131inter0, gate131inter1, gate131inter2, gate131inter3, gate131inter4, gate131inter5, gate131inter6, gate131inter7, gate131inter8, gate131inter9, gate131inter10, gate131inter11, gate131inter12, gate18inter0, gate18inter1, gate18inter2, gate18inter3, gate18inter4, gate18inter5, gate18inter6, gate18inter7, gate18inter8, gate18inter9, gate18inter10, gate18inter11, gate18inter12, gate201inter0, gate201inter1, gate201inter2, gate201inter3, gate201inter4, gate201inter5, gate201inter6, gate201inter7, gate201inter8, gate201inter9, gate201inter10, gate201inter11, gate201inter12, gate61inter0, gate61inter1, gate61inter2, gate61inter3, gate61inter4, gate61inter5, gate61inter6, gate61inter7, gate61inter8, gate61inter9, gate61inter10, gate61inter11, gate61inter12, gate117inter0, gate117inter1, gate117inter2, gate117inter3, gate117inter4, gate117inter5, gate117inter6, gate117inter7, gate117inter8, gate117inter9, gate117inter10, gate117inter11, gate117inter12, gate418inter0, gate418inter1, gate418inter2, gate418inter3, gate418inter4, gate418inter5, gate418inter6, gate418inter7, gate418inter8, gate418inter9, gate418inter10, gate418inter11, gate418inter12, gate474inter0, gate474inter1, gate474inter2, gate474inter3, gate474inter4, gate474inter5, gate474inter6, gate474inter7, gate474inter8, gate474inter9, gate474inter10, gate474inter11, gate474inter12, gate449inter0, gate449inter1, gate449inter2, gate449inter3, gate449inter4, gate449inter5, gate449inter6, gate449inter7, gate449inter8, gate449inter9, gate449inter10, gate449inter11, gate449inter12, gate16inter0, gate16inter1, gate16inter2, gate16inter3, gate16inter4, gate16inter5, gate16inter6, gate16inter7, gate16inter8, gate16inter9, gate16inter10, gate16inter11, gate16inter12, gate143inter0, gate143inter1, gate143inter2, gate143inter3, gate143inter4, gate143inter5, gate143inter6, gate143inter7, gate143inter8, gate143inter9, gate143inter10, gate143inter11, gate143inter12, gate230inter0, gate230inter1, gate230inter2, gate230inter3, gate230inter4, gate230inter5, gate230inter6, gate230inter7, gate230inter8, gate230inter9, gate230inter10, gate230inter11, gate230inter12, gate393inter0, gate393inter1, gate393inter2, gate393inter3, gate393inter4, gate393inter5, gate393inter6, gate393inter7, gate393inter8, gate393inter9, gate393inter10, gate393inter11, gate393inter12, gate417inter0, gate417inter1, gate417inter2, gate417inter3, gate417inter4, gate417inter5, gate417inter6, gate417inter7, gate417inter8, gate417inter9, gate417inter10, gate417inter11, gate417inter12, gate190inter0, gate190inter1, gate190inter2, gate190inter3, gate190inter4, gate190inter5, gate190inter6, gate190inter7, gate190inter8, gate190inter9, gate190inter10, gate190inter11, gate190inter12, gate203inter0, gate203inter1, gate203inter2, gate203inter3, gate203inter4, gate203inter5, gate203inter6, gate203inter7, gate203inter8, gate203inter9, gate203inter10, gate203inter11, gate203inter12, gate511inter0, gate511inter1, gate511inter2, gate511inter3, gate511inter4, gate511inter5, gate511inter6, gate511inter7, gate511inter8, gate511inter9, gate511inter10, gate511inter11, gate511inter12, gate39inter0, gate39inter1, gate39inter2, gate39inter3, gate39inter4, gate39inter5, gate39inter6, gate39inter7, gate39inter8, gate39inter9, gate39inter10, gate39inter11, gate39inter12, gate35inter0, gate35inter1, gate35inter2, gate35inter3, gate35inter4, gate35inter5, gate35inter6, gate35inter7, gate35inter8, gate35inter9, gate35inter10, gate35inter11, gate35inter12, gate497inter0, gate497inter1, gate497inter2, gate497inter3, gate497inter4, gate497inter5, gate497inter6, gate497inter7, gate497inter8, gate497inter9, gate497inter10, gate497inter11, gate497inter12, gate251inter0, gate251inter1, gate251inter2, gate251inter3, gate251inter4, gate251inter5, gate251inter6, gate251inter7, gate251inter8, gate251inter9, gate251inter10, gate251inter11, gate251inter12, gate151inter0, gate151inter1, gate151inter2, gate151inter3, gate151inter4, gate151inter5, gate151inter6, gate151inter7, gate151inter8, gate151inter9, gate151inter10, gate151inter11, gate151inter12, gate104inter0, gate104inter1, gate104inter2, gate104inter3, gate104inter4, gate104inter5, gate104inter6, gate104inter7, gate104inter8, gate104inter9, gate104inter10, gate104inter11, gate104inter12, gate41inter0, gate41inter1, gate41inter2, gate41inter3, gate41inter4, gate41inter5, gate41inter6, gate41inter7, gate41inter8, gate41inter9, gate41inter10, gate41inter11, gate41inter12, gate81inter0, gate81inter1, gate81inter2, gate81inter3, gate81inter4, gate81inter5, gate81inter6, gate81inter7, gate81inter8, gate81inter9, gate81inter10, gate81inter11, gate81inter12, gate82inter0, gate82inter1, gate82inter2, gate82inter3, gate82inter4, gate82inter5, gate82inter6, gate82inter7, gate82inter8, gate82inter9, gate82inter10, gate82inter11, gate82inter12, gate65inter0, gate65inter1, gate65inter2, gate65inter3, gate65inter4, gate65inter5, gate65inter6, gate65inter7, gate65inter8, gate65inter9, gate65inter10, gate65inter11, gate65inter12, gate15inter0, gate15inter1, gate15inter2, gate15inter3, gate15inter4, gate15inter5, gate15inter6, gate15inter7, gate15inter8, gate15inter9, gate15inter10, gate15inter11, gate15inter12, gate169inter0, gate169inter1, gate169inter2, gate169inter3, gate169inter4, gate169inter5, gate169inter6, gate169inter7, gate169inter8, gate169inter9, gate169inter10, gate169inter11, gate169inter12, gate53inter0, gate53inter1, gate53inter2, gate53inter3, gate53inter4, gate53inter5, gate53inter6, gate53inter7, gate53inter8, gate53inter9, gate53inter10, gate53inter11, gate53inter12, gate429inter0, gate429inter1, gate429inter2, gate429inter3, gate429inter4, gate429inter5, gate429inter6, gate429inter7, gate429inter8, gate429inter9, gate429inter10, gate429inter11, gate429inter12, gate126inter0, gate126inter1, gate126inter2, gate126inter3, gate126inter4, gate126inter5, gate126inter6, gate126inter7, gate126inter8, gate126inter9, gate126inter10, gate126inter11, gate126inter12, gate408inter0, gate408inter1, gate408inter2, gate408inter3, gate408inter4, gate408inter5, gate408inter6, gate408inter7, gate408inter8, gate408inter9, gate408inter10, gate408inter11, gate408inter12, gate494inter0, gate494inter1, gate494inter2, gate494inter3, gate494inter4, gate494inter5, gate494inter6, gate494inter7, gate494inter8, gate494inter9, gate494inter10, gate494inter11, gate494inter12, gate109inter0, gate109inter1, gate109inter2, gate109inter3, gate109inter4, gate109inter5, gate109inter6, gate109inter7, gate109inter8, gate109inter9, gate109inter10, gate109inter11, gate109inter12, gate64inter0, gate64inter1, gate64inter2, gate64inter3, gate64inter4, gate64inter5, gate64inter6, gate64inter7, gate64inter8, gate64inter9, gate64inter10, gate64inter11, gate64inter12, gate477inter0, gate477inter1, gate477inter2, gate477inter3, gate477inter4, gate477inter5, gate477inter6, gate477inter7, gate477inter8, gate477inter9, gate477inter10, gate477inter11, gate477inter12, gate187inter0, gate187inter1, gate187inter2, gate187inter3, gate187inter4, gate187inter5, gate187inter6, gate187inter7, gate187inter8, gate187inter9, gate187inter10, gate187inter11, gate187inter12, gate406inter0, gate406inter1, gate406inter2, gate406inter3, gate406inter4, gate406inter5, gate406inter6, gate406inter7, gate406inter8, gate406inter9, gate406inter10, gate406inter11, gate406inter12, gate129inter0, gate129inter1, gate129inter2, gate129inter3, gate129inter4, gate129inter5, gate129inter6, gate129inter7, gate129inter8, gate129inter9, gate129inter10, gate129inter11, gate129inter12, gate186inter0, gate186inter1, gate186inter2, gate186inter3, gate186inter4, gate186inter5, gate186inter6, gate186inter7, gate186inter8, gate186inter9, gate186inter10, gate186inter11, gate186inter12, gate91inter0, gate91inter1, gate91inter2, gate91inter3, gate91inter4, gate91inter5, gate91inter6, gate91inter7, gate91inter8, gate91inter9, gate91inter10, gate91inter11, gate91inter12, gate253inter0, gate253inter1, gate253inter2, gate253inter3, gate253inter4, gate253inter5, gate253inter6, gate253inter7, gate253inter8, gate253inter9, gate253inter10, gate253inter11, gate253inter12, gate120inter0, gate120inter1, gate120inter2, gate120inter3, gate120inter4, gate120inter5, gate120inter6, gate120inter7, gate120inter8, gate120inter9, gate120inter10, gate120inter11, gate120inter12, gate77inter0, gate77inter1, gate77inter2, gate77inter3, gate77inter4, gate77inter5, gate77inter6, gate77inter7, gate77inter8, gate77inter9, gate77inter10, gate77inter11, gate77inter12, gate188inter0, gate188inter1, gate188inter2, gate188inter3, gate188inter4, gate188inter5, gate188inter6, gate188inter7, gate188inter8, gate188inter9, gate188inter10, gate188inter11, gate188inter12, gate96inter0, gate96inter1, gate96inter2, gate96inter3, gate96inter4, gate96inter5, gate96inter6, gate96inter7, gate96inter8, gate96inter9, gate96inter10, gate96inter11, gate96inter12, gate233inter0, gate233inter1, gate233inter2, gate233inter3, gate233inter4, gate233inter5, gate233inter6, gate233inter7, gate233inter8, gate233inter9, gate233inter10, gate233inter11, gate233inter12, gate496inter0, gate496inter1, gate496inter2, gate496inter3, gate496inter4, gate496inter5, gate496inter6, gate496inter7, gate496inter8, gate496inter9, gate496inter10, gate496inter11, gate496inter12, gate121inter0, gate121inter1, gate121inter2, gate121inter3, gate121inter4, gate121inter5, gate121inter6, gate121inter7, gate121inter8, gate121inter9, gate121inter10, gate121inter11, gate121inter12, gate426inter0, gate426inter1, gate426inter2, gate426inter3, gate426inter4, gate426inter5, gate426inter6, gate426inter7, gate426inter8, gate426inter9, gate426inter10, gate426inter11, gate426inter12, gate501inter0, gate501inter1, gate501inter2, gate501inter3, gate501inter4, gate501inter5, gate501inter6, gate501inter7, gate501inter8, gate501inter9, gate501inter10, gate501inter11, gate501inter12, gate63inter0, gate63inter1, gate63inter2, gate63inter3, gate63inter4, gate63inter5, gate63inter6, gate63inter7, gate63inter8, gate63inter9, gate63inter10, gate63inter11, gate63inter12, gate170inter0, gate170inter1, gate170inter2, gate170inter3, gate170inter4, gate170inter5, gate170inter6, gate170inter7, gate170inter8, gate170inter9, gate170inter10, gate170inter11, gate170inter12, gate38inter0, gate38inter1, gate38inter2, gate38inter3, gate38inter4, gate38inter5, gate38inter6, gate38inter7, gate38inter8, gate38inter9, gate38inter10, gate38inter11, gate38inter12, gate181inter0, gate181inter1, gate181inter2, gate181inter3, gate181inter4, gate181inter5, gate181inter6, gate181inter7, gate181inter8, gate181inter9, gate181inter10, gate181inter11, gate181inter12, gate249inter0, gate249inter1, gate249inter2, gate249inter3, gate249inter4, gate249inter5, gate249inter6, gate249inter7, gate249inter8, gate249inter9, gate249inter10, gate249inter11, gate249inter12, gate202inter0, gate202inter1, gate202inter2, gate202inter3, gate202inter4, gate202inter5, gate202inter6, gate202inter7, gate202inter8, gate202inter9, gate202inter10, gate202inter11, gate202inter12, gate261inter0, gate261inter1, gate261inter2, gate261inter3, gate261inter4, gate261inter5, gate261inter6, gate261inter7, gate261inter8, gate261inter9, gate261inter10, gate261inter11, gate261inter12, gate99inter0, gate99inter1, gate99inter2, gate99inter3, gate99inter4, gate99inter5, gate99inter6, gate99inter7, gate99inter8, gate99inter9, gate99inter10, gate99inter11, gate99inter12, gate439inter0, gate439inter1, gate439inter2, gate439inter3, gate439inter4, gate439inter5, gate439inter6, gate439inter7, gate439inter8, gate439inter9, gate439inter10, gate439inter11, gate439inter12, gate512inter0, gate512inter1, gate512inter2, gate512inter3, gate512inter4, gate512inter5, gate512inter6, gate512inter7, gate512inter8, gate512inter9, gate512inter10, gate512inter11, gate512inter12, gate94inter0, gate94inter1, gate94inter2, gate94inter3, gate94inter4, gate94inter5, gate94inter6, gate94inter7, gate94inter8, gate94inter9, gate94inter10, gate94inter11, gate94inter12, gate122inter0, gate122inter1, gate122inter2, gate122inter3, gate122inter4, gate122inter5, gate122inter6, gate122inter7, gate122inter8, gate122inter9, gate122inter10, gate122inter11, gate122inter12, gate51inter0, gate51inter1, gate51inter2, gate51inter3, gate51inter4, gate51inter5, gate51inter6, gate51inter7, gate51inter8, gate51inter9, gate51inter10, gate51inter11, gate51inter12, gate395inter0, gate395inter1, gate395inter2, gate395inter3, gate395inter4, gate395inter5, gate395inter6, gate395inter7, gate395inter8, gate395inter9, gate395inter10, gate395inter11, gate395inter12, gate75inter0, gate75inter1, gate75inter2, gate75inter3, gate75inter4, gate75inter5, gate75inter6, gate75inter7, gate75inter8, gate75inter9, gate75inter10, gate75inter11, gate75inter12, gate434inter0, gate434inter1, gate434inter2, gate434inter3, gate434inter4, gate434inter5, gate434inter6, gate434inter7, gate434inter8, gate434inter9, gate434inter10, gate434inter11, gate434inter12, gate206inter0, gate206inter1, gate206inter2, gate206inter3, gate206inter4, gate206inter5, gate206inter6, gate206inter7, gate206inter8, gate206inter9, gate206inter10, gate206inter11, gate206inter12, gate480inter0, gate480inter1, gate480inter2, gate480inter3, gate480inter4, gate480inter5, gate480inter6, gate480inter7, gate480inter8, gate480inter9, gate480inter10, gate480inter11, gate480inter12, gate413inter0, gate413inter1, gate413inter2, gate413inter3, gate413inter4, gate413inter5, gate413inter6, gate413inter7, gate413inter8, gate413inter9, gate413inter10, gate413inter11, gate413inter12, gate220inter0, gate220inter1, gate220inter2, gate220inter3, gate220inter4, gate220inter5, gate220inter6, gate220inter7, gate220inter8, gate220inter9, gate220inter10, gate220inter11, gate220inter12, gate419inter0, gate419inter1, gate419inter2, gate419inter3, gate419inter4, gate419inter5, gate419inter6, gate419inter7, gate419inter8, gate419inter9, gate419inter10, gate419inter11, gate419inter12, gate159inter0, gate159inter1, gate159inter2, gate159inter3, gate159inter4, gate159inter5, gate159inter6, gate159inter7, gate159inter8, gate159inter9, gate159inter10, gate159inter11, gate159inter12, gate272inter0, gate272inter1, gate272inter2, gate272inter3, gate272inter4, gate272inter5, gate272inter6, gate272inter7, gate272inter8, gate272inter9, gate272inter10, gate272inter11, gate272inter12, gate440inter0, gate440inter1, gate440inter2, gate440inter3, gate440inter4, gate440inter5, gate440inter6, gate440inter7, gate440inter8, gate440inter9, gate440inter10, gate440inter11, gate440inter12, gate172inter0, gate172inter1, gate172inter2, gate172inter3, gate172inter4, gate172inter5, gate172inter6, gate172inter7, gate172inter8, gate172inter9, gate172inter10, gate172inter11, gate172inter12, gate215inter0, gate215inter1, gate215inter2, gate215inter3, gate215inter4, gate215inter5, gate215inter6, gate215inter7, gate215inter8, gate215inter9, gate215inter10, gate215inter11, gate215inter12, gate43inter0, gate43inter1, gate43inter2, gate43inter3, gate43inter4, gate43inter5, gate43inter6, gate43inter7, gate43inter8, gate43inter9, gate43inter10, gate43inter11, gate43inter12, gate265inter0, gate265inter1, gate265inter2, gate265inter3, gate265inter4, gate265inter5, gate265inter6, gate265inter7, gate265inter8, gate265inter9, gate265inter10, gate265inter11, gate265inter12, gate240inter0, gate240inter1, gate240inter2, gate240inter3, gate240inter4, gate240inter5, gate240inter6, gate240inter7, gate240inter8, gate240inter9, gate240inter10, gate240inter11, gate240inter12, gate161inter0, gate161inter1, gate161inter2, gate161inter3, gate161inter4, gate161inter5, gate161inter6, gate161inter7, gate161inter8, gate161inter9, gate161inter10, gate161inter11, gate161inter12, gate280inter0, gate280inter1, gate280inter2, gate280inter3, gate280inter4, gate280inter5, gate280inter6, gate280inter7, gate280inter8, gate280inter9, gate280inter10, gate280inter11, gate280inter12, gate166inter0, gate166inter1, gate166inter2, gate166inter3, gate166inter4, gate166inter5, gate166inter6, gate166inter7, gate166inter8, gate166inter9, gate166inter10, gate166inter11, gate166inter12, gate74inter0, gate74inter1, gate74inter2, gate74inter3, gate74inter4, gate74inter5, gate74inter6, gate74inter7, gate74inter8, gate74inter9, gate74inter10, gate74inter11, gate74inter12, gate257inter0, gate257inter1, gate257inter2, gate257inter3, gate257inter4, gate257inter5, gate257inter6, gate257inter7, gate257inter8, gate257inter9, gate257inter10, gate257inter11, gate257inter12, gate432inter0, gate432inter1, gate432inter2, gate432inter3, gate432inter4, gate432inter5, gate432inter6, gate432inter7, gate432inter8, gate432inter9, gate432inter10, gate432inter11, gate432inter12, gate175inter0, gate175inter1, gate175inter2, gate175inter3, gate175inter4, gate175inter5, gate175inter6, gate175inter7, gate175inter8, gate175inter9, gate175inter10, gate175inter11, gate175inter12, gate468inter0, gate468inter1, gate468inter2, gate468inter3, gate468inter4, gate468inter5, gate468inter6, gate468inter7, gate468inter8, gate468inter9, gate468inter10, gate468inter11, gate468inter12, gate46inter0, gate46inter1, gate46inter2, gate46inter3, gate46inter4, gate46inter5, gate46inter6, gate46inter7, gate46inter8, gate46inter9, gate46inter10, gate46inter11, gate46inter12, gate113inter0, gate113inter1, gate113inter2, gate113inter3, gate113inter4, gate113inter5, gate113inter6, gate113inter7, gate113inter8, gate113inter9, gate113inter10, gate113inter11, gate113inter12, gate390inter0, gate390inter1, gate390inter2, gate390inter3, gate390inter4, gate390inter5, gate390inter6, gate390inter7, gate390inter8, gate390inter9, gate390inter10, gate390inter11, gate390inter12, gate278inter0, gate278inter1, gate278inter2, gate278inter3, gate278inter4, gate278inter5, gate278inter6, gate278inter7, gate278inter8, gate278inter9, gate278inter10, gate278inter11, gate278inter12, gate263inter0, gate263inter1, gate263inter2, gate263inter3, gate263inter4, gate263inter5, gate263inter6, gate263inter7, gate263inter8, gate263inter9, gate263inter10, gate263inter11, gate263inter12, gate425inter0, gate425inter1, gate425inter2, gate425inter3, gate425inter4, gate425inter5, gate425inter6, gate425inter7, gate425inter8, gate425inter9, gate425inter10, gate425inter11, gate425inter12, gate24inter0, gate24inter1, gate24inter2, gate24inter3, gate24inter4, gate24inter5, gate24inter6, gate24inter7, gate24inter8, gate24inter9, gate24inter10, gate24inter11, gate24inter12, gate97inter0, gate97inter1, gate97inter2, gate97inter3, gate97inter4, gate97inter5, gate97inter6, gate97inter7, gate97inter8, gate97inter9, gate97inter10, gate97inter11, gate97inter12, gate392inter0, gate392inter1, gate392inter2, gate392inter3, gate392inter4, gate392inter5, gate392inter6, gate392inter7, gate392inter8, gate392inter9, gate392inter10, gate392inter11, gate392inter12, gate437inter0, gate437inter1, gate437inter2, gate437inter3, gate437inter4, gate437inter5, gate437inter6, gate437inter7, gate437inter8, gate437inter9, gate437inter10, gate437inter11, gate437inter12, gate162inter0, gate162inter1, gate162inter2, gate162inter3, gate162inter4, gate162inter5, gate162inter6, gate162inter7, gate162inter8, gate162inter9, gate162inter10, gate162inter11, gate162inter12, gate134inter0, gate134inter1, gate134inter2, gate134inter3, gate134inter4, gate134inter5, gate134inter6, gate134inter7, gate134inter8, gate134inter9, gate134inter10, gate134inter11, gate134inter12, gate483inter0, gate483inter1, gate483inter2, gate483inter3, gate483inter4, gate483inter5, gate483inter6, gate483inter7, gate483inter8, gate483inter9, gate483inter10, gate483inter11, gate483inter12, gate37inter0, gate37inter1, gate37inter2, gate37inter3, gate37inter4, gate37inter5, gate37inter6, gate37inter7, gate37inter8, gate37inter9, gate37inter10, gate37inter11, gate37inter12, gate506inter0, gate506inter1, gate506inter2, gate506inter3, gate506inter4, gate506inter5, gate506inter6, gate506inter7, gate506inter8, gate506inter9, gate506inter10, gate506inter11, gate506inter12, gate179inter0, gate179inter1, gate179inter2, gate179inter3, gate179inter4, gate179inter5, gate179inter6, gate179inter7, gate179inter8, gate179inter9, gate179inter10, gate179inter11, gate179inter12, gate68inter0, gate68inter1, gate68inter2, gate68inter3, gate68inter4, gate68inter5, gate68inter6, gate68inter7, gate68inter8, gate68inter9, gate68inter10, gate68inter11, gate68inter12, gate87inter0, gate87inter1, gate87inter2, gate87inter3, gate87inter4, gate87inter5, gate87inter6, gate87inter7, gate87inter8, gate87inter9, gate87inter10, gate87inter11, gate87inter12, gate124inter0, gate124inter1, gate124inter2, gate124inter3, gate124inter4, gate124inter5, gate124inter6, gate124inter7, gate124inter8, gate124inter9, gate124inter10, gate124inter11, gate124inter12, gate510inter0, gate510inter1, gate510inter2, gate510inter3, gate510inter4, gate510inter5, gate510inter6, gate510inter7, gate510inter8, gate510inter9, gate510inter10, gate510inter11, gate510inter12, gate391inter0, gate391inter1, gate391inter2, gate391inter3, gate391inter4, gate391inter5, gate391inter6, gate391inter7, gate391inter8, gate391inter9, gate391inter10, gate391inter11, gate391inter12, gate416inter0, gate416inter1, gate416inter2, gate416inter3, gate416inter4, gate416inter5, gate416inter6, gate416inter7, gate416inter8, gate416inter9, gate416inter10, gate416inter11, gate416inter12, gate407inter0, gate407inter1, gate407inter2, gate407inter3, gate407inter4, gate407inter5, gate407inter6, gate407inter7, gate407inter8, gate407inter9, gate407inter10, gate407inter11, gate407inter12, gate30inter0, gate30inter1, gate30inter2, gate30inter3, gate30inter4, gate30inter5, gate30inter6, gate30inter7, gate30inter8, gate30inter9, gate30inter10, gate30inter11, gate30inter12, gate466inter0, gate466inter1, gate466inter2, gate466inter3, gate466inter4, gate466inter5, gate466inter6, gate466inter7, gate466inter8, gate466inter9, gate466inter10, gate466inter11, gate466inter12, gate290inter0, gate290inter1, gate290inter2, gate290inter3, gate290inter4, gate290inter5, gate290inter6, gate290inter7, gate290inter8, gate290inter9, gate290inter10, gate290inter11, gate290inter12, gate508inter0, gate508inter1, gate508inter2, gate508inter3, gate508inter4, gate508inter5, gate508inter6, gate508inter7, gate508inter8, gate508inter9, gate508inter10, gate508inter11, gate508inter12, gate125inter0, gate125inter1, gate125inter2, gate125inter3, gate125inter4, gate125inter5, gate125inter6, gate125inter7, gate125inter8, gate125inter9, gate125inter10, gate125inter11, gate125inter12;



and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );
nand2 gate9( .a(G1), .b(G2), .O(G266) );
nand2 gate10( .a(G3), .b(G4), .O(G269) );
nand2 gate11( .a(G5), .b(G6), .O(G272) );
nand2 gate12( .a(G7), .b(G8), .O(G275) );
nand2 gate13( .a(G9), .b(G10), .O(G278) );
nand2 gate14( .a(G11), .b(G12), .O(G281) );

  xor2  gate981(.a(G14), .b(G13), .O(gate15inter0));
  nand2 gate982(.a(gate15inter0), .b(s_62), .O(gate15inter1));
  and2  gate983(.a(G14), .b(G13), .O(gate15inter2));
  inv1  gate984(.a(s_62), .O(gate15inter3));
  inv1  gate985(.a(s_63), .O(gate15inter4));
  nand2 gate986(.a(gate15inter4), .b(gate15inter3), .O(gate15inter5));
  nor2  gate987(.a(gate15inter5), .b(gate15inter2), .O(gate15inter6));
  inv1  gate988(.a(G13), .O(gate15inter7));
  inv1  gate989(.a(G14), .O(gate15inter8));
  nand2 gate990(.a(gate15inter8), .b(gate15inter7), .O(gate15inter9));
  nand2 gate991(.a(s_63), .b(gate15inter3), .O(gate15inter10));
  nor2  gate992(.a(gate15inter10), .b(gate15inter9), .O(gate15inter11));
  nor2  gate993(.a(gate15inter11), .b(gate15inter6), .O(gate15inter12));
  nand2 gate994(.a(gate15inter12), .b(gate15inter1), .O(G284));

  xor2  gate729(.a(G16), .b(G15), .O(gate16inter0));
  nand2 gate730(.a(gate16inter0), .b(s_26), .O(gate16inter1));
  and2  gate731(.a(G16), .b(G15), .O(gate16inter2));
  inv1  gate732(.a(s_26), .O(gate16inter3));
  inv1  gate733(.a(s_27), .O(gate16inter4));
  nand2 gate734(.a(gate16inter4), .b(gate16inter3), .O(gate16inter5));
  nor2  gate735(.a(gate16inter5), .b(gate16inter2), .O(gate16inter6));
  inv1  gate736(.a(G15), .O(gate16inter7));
  inv1  gate737(.a(G16), .O(gate16inter8));
  nand2 gate738(.a(gate16inter8), .b(gate16inter7), .O(gate16inter9));
  nand2 gate739(.a(s_27), .b(gate16inter3), .O(gate16inter10));
  nor2  gate740(.a(gate16inter10), .b(gate16inter9), .O(gate16inter11));
  nor2  gate741(.a(gate16inter11), .b(gate16inter6), .O(gate16inter12));
  nand2 gate742(.a(gate16inter12), .b(gate16inter1), .O(G287));
nand2 gate17( .a(G17), .b(G18), .O(G290) );

  xor2  gate631(.a(G20), .b(G19), .O(gate18inter0));
  nand2 gate632(.a(gate18inter0), .b(s_12), .O(gate18inter1));
  and2  gate633(.a(G20), .b(G19), .O(gate18inter2));
  inv1  gate634(.a(s_12), .O(gate18inter3));
  inv1  gate635(.a(s_13), .O(gate18inter4));
  nand2 gate636(.a(gate18inter4), .b(gate18inter3), .O(gate18inter5));
  nor2  gate637(.a(gate18inter5), .b(gate18inter2), .O(gate18inter6));
  inv1  gate638(.a(G19), .O(gate18inter7));
  inv1  gate639(.a(G20), .O(gate18inter8));
  nand2 gate640(.a(gate18inter8), .b(gate18inter7), .O(gate18inter9));
  nand2 gate641(.a(s_13), .b(gate18inter3), .O(gate18inter10));
  nor2  gate642(.a(gate18inter10), .b(gate18inter9), .O(gate18inter11));
  nor2  gate643(.a(gate18inter11), .b(gate18inter6), .O(gate18inter12));
  nand2 gate644(.a(gate18inter12), .b(gate18inter1), .O(G293));
nand2 gate19( .a(G21), .b(G22), .O(G296) );
nand2 gate20( .a(G23), .b(G24), .O(G299) );
nand2 gate21( .a(G25), .b(G26), .O(G302) );
nand2 gate22( .a(G27), .b(G28), .O(G305) );
nand2 gate23( .a(G29), .b(G30), .O(G308) );

  xor2  gate1933(.a(G32), .b(G31), .O(gate24inter0));
  nand2 gate1934(.a(gate24inter0), .b(s_198), .O(gate24inter1));
  and2  gate1935(.a(G32), .b(G31), .O(gate24inter2));
  inv1  gate1936(.a(s_198), .O(gate24inter3));
  inv1  gate1937(.a(s_199), .O(gate24inter4));
  nand2 gate1938(.a(gate24inter4), .b(gate24inter3), .O(gate24inter5));
  nor2  gate1939(.a(gate24inter5), .b(gate24inter2), .O(gate24inter6));
  inv1  gate1940(.a(G31), .O(gate24inter7));
  inv1  gate1941(.a(G32), .O(gate24inter8));
  nand2 gate1942(.a(gate24inter8), .b(gate24inter7), .O(gate24inter9));
  nand2 gate1943(.a(s_199), .b(gate24inter3), .O(gate24inter10));
  nor2  gate1944(.a(gate24inter10), .b(gate24inter9), .O(gate24inter11));
  nor2  gate1945(.a(gate24inter11), .b(gate24inter6), .O(gate24inter12));
  nand2 gate1946(.a(gate24inter12), .b(gate24inter1), .O(G311));
nand2 gate25( .a(G1), .b(G5), .O(G314) );

  xor2  gate589(.a(G13), .b(G9), .O(gate26inter0));
  nand2 gate590(.a(gate26inter0), .b(s_6), .O(gate26inter1));
  and2  gate591(.a(G13), .b(G9), .O(gate26inter2));
  inv1  gate592(.a(s_6), .O(gate26inter3));
  inv1  gate593(.a(s_7), .O(gate26inter4));
  nand2 gate594(.a(gate26inter4), .b(gate26inter3), .O(gate26inter5));
  nor2  gate595(.a(gate26inter5), .b(gate26inter2), .O(gate26inter6));
  inv1  gate596(.a(G9), .O(gate26inter7));
  inv1  gate597(.a(G13), .O(gate26inter8));
  nand2 gate598(.a(gate26inter8), .b(gate26inter7), .O(gate26inter9));
  nand2 gate599(.a(s_7), .b(gate26inter3), .O(gate26inter10));
  nor2  gate600(.a(gate26inter10), .b(gate26inter9), .O(gate26inter11));
  nor2  gate601(.a(gate26inter11), .b(gate26inter6), .O(gate26inter12));
  nand2 gate602(.a(gate26inter12), .b(gate26inter1), .O(G317));
nand2 gate27( .a(G2), .b(G6), .O(G320) );
nand2 gate28( .a(G10), .b(G14), .O(G323) );
nand2 gate29( .a(G3), .b(G7), .O(G326) );

  xor2  gate2171(.a(G15), .b(G11), .O(gate30inter0));
  nand2 gate2172(.a(gate30inter0), .b(s_232), .O(gate30inter1));
  and2  gate2173(.a(G15), .b(G11), .O(gate30inter2));
  inv1  gate2174(.a(s_232), .O(gate30inter3));
  inv1  gate2175(.a(s_233), .O(gate30inter4));
  nand2 gate2176(.a(gate30inter4), .b(gate30inter3), .O(gate30inter5));
  nor2  gate2177(.a(gate30inter5), .b(gate30inter2), .O(gate30inter6));
  inv1  gate2178(.a(G11), .O(gate30inter7));
  inv1  gate2179(.a(G15), .O(gate30inter8));
  nand2 gate2180(.a(gate30inter8), .b(gate30inter7), .O(gate30inter9));
  nand2 gate2181(.a(s_233), .b(gate30inter3), .O(gate30inter10));
  nor2  gate2182(.a(gate30inter10), .b(gate30inter9), .O(gate30inter11));
  nor2  gate2183(.a(gate30inter11), .b(gate30inter6), .O(gate30inter12));
  nand2 gate2184(.a(gate30inter12), .b(gate30inter1), .O(G329));
nand2 gate31( .a(G4), .b(G8), .O(G332) );
nand2 gate32( .a(G12), .b(G16), .O(G335) );
nand2 gate33( .a(G17), .b(G21), .O(G338) );
nand2 gate34( .a(G25), .b(G29), .O(G341) );

  xor2  gate855(.a(G22), .b(G18), .O(gate35inter0));
  nand2 gate856(.a(gate35inter0), .b(s_44), .O(gate35inter1));
  and2  gate857(.a(G22), .b(G18), .O(gate35inter2));
  inv1  gate858(.a(s_44), .O(gate35inter3));
  inv1  gate859(.a(s_45), .O(gate35inter4));
  nand2 gate860(.a(gate35inter4), .b(gate35inter3), .O(gate35inter5));
  nor2  gate861(.a(gate35inter5), .b(gate35inter2), .O(gate35inter6));
  inv1  gate862(.a(G18), .O(gate35inter7));
  inv1  gate863(.a(G22), .O(gate35inter8));
  nand2 gate864(.a(gate35inter8), .b(gate35inter7), .O(gate35inter9));
  nand2 gate865(.a(s_45), .b(gate35inter3), .O(gate35inter10));
  nor2  gate866(.a(gate35inter10), .b(gate35inter9), .O(gate35inter11));
  nor2  gate867(.a(gate35inter11), .b(gate35inter6), .O(gate35inter12));
  nand2 gate868(.a(gate35inter12), .b(gate35inter1), .O(G344));
nand2 gate36( .a(G26), .b(G30), .O(G347) );

  xor2  gate2031(.a(G23), .b(G19), .O(gate37inter0));
  nand2 gate2032(.a(gate37inter0), .b(s_212), .O(gate37inter1));
  and2  gate2033(.a(G23), .b(G19), .O(gate37inter2));
  inv1  gate2034(.a(s_212), .O(gate37inter3));
  inv1  gate2035(.a(s_213), .O(gate37inter4));
  nand2 gate2036(.a(gate37inter4), .b(gate37inter3), .O(gate37inter5));
  nor2  gate2037(.a(gate37inter5), .b(gate37inter2), .O(gate37inter6));
  inv1  gate2038(.a(G19), .O(gate37inter7));
  inv1  gate2039(.a(G23), .O(gate37inter8));
  nand2 gate2040(.a(gate37inter8), .b(gate37inter7), .O(gate37inter9));
  nand2 gate2041(.a(s_213), .b(gate37inter3), .O(gate37inter10));
  nor2  gate2042(.a(gate37inter10), .b(gate37inter9), .O(gate37inter11));
  nor2  gate2043(.a(gate37inter11), .b(gate37inter6), .O(gate37inter12));
  nand2 gate2044(.a(gate37inter12), .b(gate37inter1), .O(G350));

  xor2  gate1359(.a(G31), .b(G27), .O(gate38inter0));
  nand2 gate1360(.a(gate38inter0), .b(s_116), .O(gate38inter1));
  and2  gate1361(.a(G31), .b(G27), .O(gate38inter2));
  inv1  gate1362(.a(s_116), .O(gate38inter3));
  inv1  gate1363(.a(s_117), .O(gate38inter4));
  nand2 gate1364(.a(gate38inter4), .b(gate38inter3), .O(gate38inter5));
  nor2  gate1365(.a(gate38inter5), .b(gate38inter2), .O(gate38inter6));
  inv1  gate1366(.a(G27), .O(gate38inter7));
  inv1  gate1367(.a(G31), .O(gate38inter8));
  nand2 gate1368(.a(gate38inter8), .b(gate38inter7), .O(gate38inter9));
  nand2 gate1369(.a(s_117), .b(gate38inter3), .O(gate38inter10));
  nor2  gate1370(.a(gate38inter10), .b(gate38inter9), .O(gate38inter11));
  nor2  gate1371(.a(gate38inter11), .b(gate38inter6), .O(gate38inter12));
  nand2 gate1372(.a(gate38inter12), .b(gate38inter1), .O(G353));

  xor2  gate841(.a(G24), .b(G20), .O(gate39inter0));
  nand2 gate842(.a(gate39inter0), .b(s_42), .O(gate39inter1));
  and2  gate843(.a(G24), .b(G20), .O(gate39inter2));
  inv1  gate844(.a(s_42), .O(gate39inter3));
  inv1  gate845(.a(s_43), .O(gate39inter4));
  nand2 gate846(.a(gate39inter4), .b(gate39inter3), .O(gate39inter5));
  nor2  gate847(.a(gate39inter5), .b(gate39inter2), .O(gate39inter6));
  inv1  gate848(.a(G20), .O(gate39inter7));
  inv1  gate849(.a(G24), .O(gate39inter8));
  nand2 gate850(.a(gate39inter8), .b(gate39inter7), .O(gate39inter9));
  nand2 gate851(.a(s_43), .b(gate39inter3), .O(gate39inter10));
  nor2  gate852(.a(gate39inter10), .b(gate39inter9), .O(gate39inter11));
  nor2  gate853(.a(gate39inter11), .b(gate39inter6), .O(gate39inter12));
  nand2 gate854(.a(gate39inter12), .b(gate39inter1), .O(G356));
nand2 gate40( .a(G28), .b(G32), .O(G359) );

  xor2  gate925(.a(G266), .b(G1), .O(gate41inter0));
  nand2 gate926(.a(gate41inter0), .b(s_54), .O(gate41inter1));
  and2  gate927(.a(G266), .b(G1), .O(gate41inter2));
  inv1  gate928(.a(s_54), .O(gate41inter3));
  inv1  gate929(.a(s_55), .O(gate41inter4));
  nand2 gate930(.a(gate41inter4), .b(gate41inter3), .O(gate41inter5));
  nor2  gate931(.a(gate41inter5), .b(gate41inter2), .O(gate41inter6));
  inv1  gate932(.a(G1), .O(gate41inter7));
  inv1  gate933(.a(G266), .O(gate41inter8));
  nand2 gate934(.a(gate41inter8), .b(gate41inter7), .O(gate41inter9));
  nand2 gate935(.a(s_55), .b(gate41inter3), .O(gate41inter10));
  nor2  gate936(.a(gate41inter10), .b(gate41inter9), .O(gate41inter11));
  nor2  gate937(.a(gate41inter11), .b(gate41inter6), .O(gate41inter12));
  nand2 gate938(.a(gate41inter12), .b(gate41inter1), .O(G362));
nand2 gate42( .a(G2), .b(G266), .O(G363) );

  xor2  gate1695(.a(G269), .b(G3), .O(gate43inter0));
  nand2 gate1696(.a(gate43inter0), .b(s_164), .O(gate43inter1));
  and2  gate1697(.a(G269), .b(G3), .O(gate43inter2));
  inv1  gate1698(.a(s_164), .O(gate43inter3));
  inv1  gate1699(.a(s_165), .O(gate43inter4));
  nand2 gate1700(.a(gate43inter4), .b(gate43inter3), .O(gate43inter5));
  nor2  gate1701(.a(gate43inter5), .b(gate43inter2), .O(gate43inter6));
  inv1  gate1702(.a(G3), .O(gate43inter7));
  inv1  gate1703(.a(G269), .O(gate43inter8));
  nand2 gate1704(.a(gate43inter8), .b(gate43inter7), .O(gate43inter9));
  nand2 gate1705(.a(s_165), .b(gate43inter3), .O(gate43inter10));
  nor2  gate1706(.a(gate43inter10), .b(gate43inter9), .O(gate43inter11));
  nor2  gate1707(.a(gate43inter11), .b(gate43inter6), .O(gate43inter12));
  nand2 gate1708(.a(gate43inter12), .b(gate43inter1), .O(G364));
nand2 gate44( .a(G4), .b(G269), .O(G365) );
nand2 gate45( .a(G5), .b(G272), .O(G366) );

  xor2  gate1849(.a(G272), .b(G6), .O(gate46inter0));
  nand2 gate1850(.a(gate46inter0), .b(s_186), .O(gate46inter1));
  and2  gate1851(.a(G272), .b(G6), .O(gate46inter2));
  inv1  gate1852(.a(s_186), .O(gate46inter3));
  inv1  gate1853(.a(s_187), .O(gate46inter4));
  nand2 gate1854(.a(gate46inter4), .b(gate46inter3), .O(gate46inter5));
  nor2  gate1855(.a(gate46inter5), .b(gate46inter2), .O(gate46inter6));
  inv1  gate1856(.a(G6), .O(gate46inter7));
  inv1  gate1857(.a(G272), .O(gate46inter8));
  nand2 gate1858(.a(gate46inter8), .b(gate46inter7), .O(gate46inter9));
  nand2 gate1859(.a(s_187), .b(gate46inter3), .O(gate46inter10));
  nor2  gate1860(.a(gate46inter10), .b(gate46inter9), .O(gate46inter11));
  nor2  gate1861(.a(gate46inter11), .b(gate46inter6), .O(gate46inter12));
  nand2 gate1862(.a(gate46inter12), .b(gate46inter1), .O(G367));
nand2 gate47( .a(G7), .b(G275), .O(G368) );
nand2 gate48( .a(G8), .b(G275), .O(G369) );
nand2 gate49( .a(G9), .b(G278), .O(G370) );
nand2 gate50( .a(G10), .b(G278), .O(G371) );

  xor2  gate1499(.a(G281), .b(G11), .O(gate51inter0));
  nand2 gate1500(.a(gate51inter0), .b(s_136), .O(gate51inter1));
  and2  gate1501(.a(G281), .b(G11), .O(gate51inter2));
  inv1  gate1502(.a(s_136), .O(gate51inter3));
  inv1  gate1503(.a(s_137), .O(gate51inter4));
  nand2 gate1504(.a(gate51inter4), .b(gate51inter3), .O(gate51inter5));
  nor2  gate1505(.a(gate51inter5), .b(gate51inter2), .O(gate51inter6));
  inv1  gate1506(.a(G11), .O(gate51inter7));
  inv1  gate1507(.a(G281), .O(gate51inter8));
  nand2 gate1508(.a(gate51inter8), .b(gate51inter7), .O(gate51inter9));
  nand2 gate1509(.a(s_137), .b(gate51inter3), .O(gate51inter10));
  nor2  gate1510(.a(gate51inter10), .b(gate51inter9), .O(gate51inter11));
  nor2  gate1511(.a(gate51inter11), .b(gate51inter6), .O(gate51inter12));
  nand2 gate1512(.a(gate51inter12), .b(gate51inter1), .O(G372));
nand2 gate52( .a(G12), .b(G281), .O(G373) );

  xor2  gate1009(.a(G284), .b(G13), .O(gate53inter0));
  nand2 gate1010(.a(gate53inter0), .b(s_66), .O(gate53inter1));
  and2  gate1011(.a(G284), .b(G13), .O(gate53inter2));
  inv1  gate1012(.a(s_66), .O(gate53inter3));
  inv1  gate1013(.a(s_67), .O(gate53inter4));
  nand2 gate1014(.a(gate53inter4), .b(gate53inter3), .O(gate53inter5));
  nor2  gate1015(.a(gate53inter5), .b(gate53inter2), .O(gate53inter6));
  inv1  gate1016(.a(G13), .O(gate53inter7));
  inv1  gate1017(.a(G284), .O(gate53inter8));
  nand2 gate1018(.a(gate53inter8), .b(gate53inter7), .O(gate53inter9));
  nand2 gate1019(.a(s_67), .b(gate53inter3), .O(gate53inter10));
  nor2  gate1020(.a(gate53inter10), .b(gate53inter9), .O(gate53inter11));
  nor2  gate1021(.a(gate53inter11), .b(gate53inter6), .O(gate53inter12));
  nand2 gate1022(.a(gate53inter12), .b(gate53inter1), .O(G374));
nand2 gate54( .a(G14), .b(G284), .O(G375) );
nand2 gate55( .a(G15), .b(G287), .O(G376) );
nand2 gate56( .a(G16), .b(G287), .O(G377) );
nand2 gate57( .a(G17), .b(G290), .O(G378) );
nand2 gate58( .a(G18), .b(G290), .O(G379) );
nand2 gate59( .a(G19), .b(G293), .O(G380) );
nand2 gate60( .a(G20), .b(G293), .O(G381) );

  xor2  gate659(.a(G296), .b(G21), .O(gate61inter0));
  nand2 gate660(.a(gate61inter0), .b(s_16), .O(gate61inter1));
  and2  gate661(.a(G296), .b(G21), .O(gate61inter2));
  inv1  gate662(.a(s_16), .O(gate61inter3));
  inv1  gate663(.a(s_17), .O(gate61inter4));
  nand2 gate664(.a(gate61inter4), .b(gate61inter3), .O(gate61inter5));
  nor2  gate665(.a(gate61inter5), .b(gate61inter2), .O(gate61inter6));
  inv1  gate666(.a(G21), .O(gate61inter7));
  inv1  gate667(.a(G296), .O(gate61inter8));
  nand2 gate668(.a(gate61inter8), .b(gate61inter7), .O(gate61inter9));
  nand2 gate669(.a(s_17), .b(gate61inter3), .O(gate61inter10));
  nor2  gate670(.a(gate61inter10), .b(gate61inter9), .O(gate61inter11));
  nor2  gate671(.a(gate61inter11), .b(gate61inter6), .O(gate61inter12));
  nand2 gate672(.a(gate61inter12), .b(gate61inter1), .O(G382));
nand2 gate62( .a(G22), .b(G296), .O(G383) );

  xor2  gate1331(.a(G299), .b(G23), .O(gate63inter0));
  nand2 gate1332(.a(gate63inter0), .b(s_112), .O(gate63inter1));
  and2  gate1333(.a(G299), .b(G23), .O(gate63inter2));
  inv1  gate1334(.a(s_112), .O(gate63inter3));
  inv1  gate1335(.a(s_113), .O(gate63inter4));
  nand2 gate1336(.a(gate63inter4), .b(gate63inter3), .O(gate63inter5));
  nor2  gate1337(.a(gate63inter5), .b(gate63inter2), .O(gate63inter6));
  inv1  gate1338(.a(G23), .O(gate63inter7));
  inv1  gate1339(.a(G299), .O(gate63inter8));
  nand2 gate1340(.a(gate63inter8), .b(gate63inter7), .O(gate63inter9));
  nand2 gate1341(.a(s_113), .b(gate63inter3), .O(gate63inter10));
  nor2  gate1342(.a(gate63inter10), .b(gate63inter9), .O(gate63inter11));
  nor2  gate1343(.a(gate63inter11), .b(gate63inter6), .O(gate63inter12));
  nand2 gate1344(.a(gate63inter12), .b(gate63inter1), .O(G384));

  xor2  gate1093(.a(G299), .b(G24), .O(gate64inter0));
  nand2 gate1094(.a(gate64inter0), .b(s_78), .O(gate64inter1));
  and2  gate1095(.a(G299), .b(G24), .O(gate64inter2));
  inv1  gate1096(.a(s_78), .O(gate64inter3));
  inv1  gate1097(.a(s_79), .O(gate64inter4));
  nand2 gate1098(.a(gate64inter4), .b(gate64inter3), .O(gate64inter5));
  nor2  gate1099(.a(gate64inter5), .b(gate64inter2), .O(gate64inter6));
  inv1  gate1100(.a(G24), .O(gate64inter7));
  inv1  gate1101(.a(G299), .O(gate64inter8));
  nand2 gate1102(.a(gate64inter8), .b(gate64inter7), .O(gate64inter9));
  nand2 gate1103(.a(s_79), .b(gate64inter3), .O(gate64inter10));
  nor2  gate1104(.a(gate64inter10), .b(gate64inter9), .O(gate64inter11));
  nor2  gate1105(.a(gate64inter11), .b(gate64inter6), .O(gate64inter12));
  nand2 gate1106(.a(gate64inter12), .b(gate64inter1), .O(G385));

  xor2  gate967(.a(G302), .b(G25), .O(gate65inter0));
  nand2 gate968(.a(gate65inter0), .b(s_60), .O(gate65inter1));
  and2  gate969(.a(G302), .b(G25), .O(gate65inter2));
  inv1  gate970(.a(s_60), .O(gate65inter3));
  inv1  gate971(.a(s_61), .O(gate65inter4));
  nand2 gate972(.a(gate65inter4), .b(gate65inter3), .O(gate65inter5));
  nor2  gate973(.a(gate65inter5), .b(gate65inter2), .O(gate65inter6));
  inv1  gate974(.a(G25), .O(gate65inter7));
  inv1  gate975(.a(G302), .O(gate65inter8));
  nand2 gate976(.a(gate65inter8), .b(gate65inter7), .O(gate65inter9));
  nand2 gate977(.a(s_61), .b(gate65inter3), .O(gate65inter10));
  nor2  gate978(.a(gate65inter10), .b(gate65inter9), .O(gate65inter11));
  nor2  gate979(.a(gate65inter11), .b(gate65inter6), .O(gate65inter12));
  nand2 gate980(.a(gate65inter12), .b(gate65inter1), .O(G386));
nand2 gate66( .a(G26), .b(G302), .O(G387) );
nand2 gate67( .a(G27), .b(G305), .O(G388) );

  xor2  gate2073(.a(G305), .b(G28), .O(gate68inter0));
  nand2 gate2074(.a(gate68inter0), .b(s_218), .O(gate68inter1));
  and2  gate2075(.a(G305), .b(G28), .O(gate68inter2));
  inv1  gate2076(.a(s_218), .O(gate68inter3));
  inv1  gate2077(.a(s_219), .O(gate68inter4));
  nand2 gate2078(.a(gate68inter4), .b(gate68inter3), .O(gate68inter5));
  nor2  gate2079(.a(gate68inter5), .b(gate68inter2), .O(gate68inter6));
  inv1  gate2080(.a(G28), .O(gate68inter7));
  inv1  gate2081(.a(G305), .O(gate68inter8));
  nand2 gate2082(.a(gate68inter8), .b(gate68inter7), .O(gate68inter9));
  nand2 gate2083(.a(s_219), .b(gate68inter3), .O(gate68inter10));
  nor2  gate2084(.a(gate68inter10), .b(gate68inter9), .O(gate68inter11));
  nor2  gate2085(.a(gate68inter11), .b(gate68inter6), .O(gate68inter12));
  nand2 gate2086(.a(gate68inter12), .b(gate68inter1), .O(G389));
nand2 gate69( .a(G29), .b(G308), .O(G390) );
nand2 gate70( .a(G30), .b(G308), .O(G391) );
nand2 gate71( .a(G31), .b(G311), .O(G392) );
nand2 gate72( .a(G32), .b(G311), .O(G393) );
nand2 gate73( .a(G1), .b(G314), .O(G394) );

  xor2  gate1779(.a(G314), .b(G5), .O(gate74inter0));
  nand2 gate1780(.a(gate74inter0), .b(s_176), .O(gate74inter1));
  and2  gate1781(.a(G314), .b(G5), .O(gate74inter2));
  inv1  gate1782(.a(s_176), .O(gate74inter3));
  inv1  gate1783(.a(s_177), .O(gate74inter4));
  nand2 gate1784(.a(gate74inter4), .b(gate74inter3), .O(gate74inter5));
  nor2  gate1785(.a(gate74inter5), .b(gate74inter2), .O(gate74inter6));
  inv1  gate1786(.a(G5), .O(gate74inter7));
  inv1  gate1787(.a(G314), .O(gate74inter8));
  nand2 gate1788(.a(gate74inter8), .b(gate74inter7), .O(gate74inter9));
  nand2 gate1789(.a(s_177), .b(gate74inter3), .O(gate74inter10));
  nor2  gate1790(.a(gate74inter10), .b(gate74inter9), .O(gate74inter11));
  nor2  gate1791(.a(gate74inter11), .b(gate74inter6), .O(gate74inter12));
  nand2 gate1792(.a(gate74inter12), .b(gate74inter1), .O(G395));

  xor2  gate1527(.a(G317), .b(G9), .O(gate75inter0));
  nand2 gate1528(.a(gate75inter0), .b(s_140), .O(gate75inter1));
  and2  gate1529(.a(G317), .b(G9), .O(gate75inter2));
  inv1  gate1530(.a(s_140), .O(gate75inter3));
  inv1  gate1531(.a(s_141), .O(gate75inter4));
  nand2 gate1532(.a(gate75inter4), .b(gate75inter3), .O(gate75inter5));
  nor2  gate1533(.a(gate75inter5), .b(gate75inter2), .O(gate75inter6));
  inv1  gate1534(.a(G9), .O(gate75inter7));
  inv1  gate1535(.a(G317), .O(gate75inter8));
  nand2 gate1536(.a(gate75inter8), .b(gate75inter7), .O(gate75inter9));
  nand2 gate1537(.a(s_141), .b(gate75inter3), .O(gate75inter10));
  nor2  gate1538(.a(gate75inter10), .b(gate75inter9), .O(gate75inter11));
  nor2  gate1539(.a(gate75inter11), .b(gate75inter6), .O(gate75inter12));
  nand2 gate1540(.a(gate75inter12), .b(gate75inter1), .O(G396));
nand2 gate76( .a(G13), .b(G317), .O(G397) );

  xor2  gate1219(.a(G320), .b(G2), .O(gate77inter0));
  nand2 gate1220(.a(gate77inter0), .b(s_96), .O(gate77inter1));
  and2  gate1221(.a(G320), .b(G2), .O(gate77inter2));
  inv1  gate1222(.a(s_96), .O(gate77inter3));
  inv1  gate1223(.a(s_97), .O(gate77inter4));
  nand2 gate1224(.a(gate77inter4), .b(gate77inter3), .O(gate77inter5));
  nor2  gate1225(.a(gate77inter5), .b(gate77inter2), .O(gate77inter6));
  inv1  gate1226(.a(G2), .O(gate77inter7));
  inv1  gate1227(.a(G320), .O(gate77inter8));
  nand2 gate1228(.a(gate77inter8), .b(gate77inter7), .O(gate77inter9));
  nand2 gate1229(.a(s_97), .b(gate77inter3), .O(gate77inter10));
  nor2  gate1230(.a(gate77inter10), .b(gate77inter9), .O(gate77inter11));
  nor2  gate1231(.a(gate77inter11), .b(gate77inter6), .O(gate77inter12));
  nand2 gate1232(.a(gate77inter12), .b(gate77inter1), .O(G398));
nand2 gate78( .a(G6), .b(G320), .O(G399) );
nand2 gate79( .a(G10), .b(G323), .O(G400) );
nand2 gate80( .a(G14), .b(G323), .O(G401) );

  xor2  gate939(.a(G326), .b(G3), .O(gate81inter0));
  nand2 gate940(.a(gate81inter0), .b(s_56), .O(gate81inter1));
  and2  gate941(.a(G326), .b(G3), .O(gate81inter2));
  inv1  gate942(.a(s_56), .O(gate81inter3));
  inv1  gate943(.a(s_57), .O(gate81inter4));
  nand2 gate944(.a(gate81inter4), .b(gate81inter3), .O(gate81inter5));
  nor2  gate945(.a(gate81inter5), .b(gate81inter2), .O(gate81inter6));
  inv1  gate946(.a(G3), .O(gate81inter7));
  inv1  gate947(.a(G326), .O(gate81inter8));
  nand2 gate948(.a(gate81inter8), .b(gate81inter7), .O(gate81inter9));
  nand2 gate949(.a(s_57), .b(gate81inter3), .O(gate81inter10));
  nor2  gate950(.a(gate81inter10), .b(gate81inter9), .O(gate81inter11));
  nor2  gate951(.a(gate81inter11), .b(gate81inter6), .O(gate81inter12));
  nand2 gate952(.a(gate81inter12), .b(gate81inter1), .O(G402));

  xor2  gate953(.a(G326), .b(G7), .O(gate82inter0));
  nand2 gate954(.a(gate82inter0), .b(s_58), .O(gate82inter1));
  and2  gate955(.a(G326), .b(G7), .O(gate82inter2));
  inv1  gate956(.a(s_58), .O(gate82inter3));
  inv1  gate957(.a(s_59), .O(gate82inter4));
  nand2 gate958(.a(gate82inter4), .b(gate82inter3), .O(gate82inter5));
  nor2  gate959(.a(gate82inter5), .b(gate82inter2), .O(gate82inter6));
  inv1  gate960(.a(G7), .O(gate82inter7));
  inv1  gate961(.a(G326), .O(gate82inter8));
  nand2 gate962(.a(gate82inter8), .b(gate82inter7), .O(gate82inter9));
  nand2 gate963(.a(s_59), .b(gate82inter3), .O(gate82inter10));
  nor2  gate964(.a(gate82inter10), .b(gate82inter9), .O(gate82inter11));
  nor2  gate965(.a(gate82inter11), .b(gate82inter6), .O(gate82inter12));
  nand2 gate966(.a(gate82inter12), .b(gate82inter1), .O(G403));
nand2 gate83( .a(G11), .b(G329), .O(G404) );
nand2 gate84( .a(G15), .b(G329), .O(G405) );
nand2 gate85( .a(G4), .b(G332), .O(G406) );
nand2 gate86( .a(G8), .b(G332), .O(G407) );

  xor2  gate2087(.a(G335), .b(G12), .O(gate87inter0));
  nand2 gate2088(.a(gate87inter0), .b(s_220), .O(gate87inter1));
  and2  gate2089(.a(G335), .b(G12), .O(gate87inter2));
  inv1  gate2090(.a(s_220), .O(gate87inter3));
  inv1  gate2091(.a(s_221), .O(gate87inter4));
  nand2 gate2092(.a(gate87inter4), .b(gate87inter3), .O(gate87inter5));
  nor2  gate2093(.a(gate87inter5), .b(gate87inter2), .O(gate87inter6));
  inv1  gate2094(.a(G12), .O(gate87inter7));
  inv1  gate2095(.a(G335), .O(gate87inter8));
  nand2 gate2096(.a(gate87inter8), .b(gate87inter7), .O(gate87inter9));
  nand2 gate2097(.a(s_221), .b(gate87inter3), .O(gate87inter10));
  nor2  gate2098(.a(gate87inter10), .b(gate87inter9), .O(gate87inter11));
  nor2  gate2099(.a(gate87inter11), .b(gate87inter6), .O(gate87inter12));
  nand2 gate2100(.a(gate87inter12), .b(gate87inter1), .O(G408));
nand2 gate88( .a(G16), .b(G335), .O(G409) );
nand2 gate89( .a(G17), .b(G338), .O(G410) );
nand2 gate90( .a(G21), .b(G338), .O(G411) );

  xor2  gate1177(.a(G341), .b(G25), .O(gate91inter0));
  nand2 gate1178(.a(gate91inter0), .b(s_90), .O(gate91inter1));
  and2  gate1179(.a(G341), .b(G25), .O(gate91inter2));
  inv1  gate1180(.a(s_90), .O(gate91inter3));
  inv1  gate1181(.a(s_91), .O(gate91inter4));
  nand2 gate1182(.a(gate91inter4), .b(gate91inter3), .O(gate91inter5));
  nor2  gate1183(.a(gate91inter5), .b(gate91inter2), .O(gate91inter6));
  inv1  gate1184(.a(G25), .O(gate91inter7));
  inv1  gate1185(.a(G341), .O(gate91inter8));
  nand2 gate1186(.a(gate91inter8), .b(gate91inter7), .O(gate91inter9));
  nand2 gate1187(.a(s_91), .b(gate91inter3), .O(gate91inter10));
  nor2  gate1188(.a(gate91inter10), .b(gate91inter9), .O(gate91inter11));
  nor2  gate1189(.a(gate91inter11), .b(gate91inter6), .O(gate91inter12));
  nand2 gate1190(.a(gate91inter12), .b(gate91inter1), .O(G412));
nand2 gate92( .a(G29), .b(G341), .O(G413) );
nand2 gate93( .a(G18), .b(G344), .O(G414) );

  xor2  gate1471(.a(G344), .b(G22), .O(gate94inter0));
  nand2 gate1472(.a(gate94inter0), .b(s_132), .O(gate94inter1));
  and2  gate1473(.a(G344), .b(G22), .O(gate94inter2));
  inv1  gate1474(.a(s_132), .O(gate94inter3));
  inv1  gate1475(.a(s_133), .O(gate94inter4));
  nand2 gate1476(.a(gate94inter4), .b(gate94inter3), .O(gate94inter5));
  nor2  gate1477(.a(gate94inter5), .b(gate94inter2), .O(gate94inter6));
  inv1  gate1478(.a(G22), .O(gate94inter7));
  inv1  gate1479(.a(G344), .O(gate94inter8));
  nand2 gate1480(.a(gate94inter8), .b(gate94inter7), .O(gate94inter9));
  nand2 gate1481(.a(s_133), .b(gate94inter3), .O(gate94inter10));
  nor2  gate1482(.a(gate94inter10), .b(gate94inter9), .O(gate94inter11));
  nor2  gate1483(.a(gate94inter11), .b(gate94inter6), .O(gate94inter12));
  nand2 gate1484(.a(gate94inter12), .b(gate94inter1), .O(G415));
nand2 gate95( .a(G26), .b(G347), .O(G416) );

  xor2  gate1247(.a(G347), .b(G30), .O(gate96inter0));
  nand2 gate1248(.a(gate96inter0), .b(s_100), .O(gate96inter1));
  and2  gate1249(.a(G347), .b(G30), .O(gate96inter2));
  inv1  gate1250(.a(s_100), .O(gate96inter3));
  inv1  gate1251(.a(s_101), .O(gate96inter4));
  nand2 gate1252(.a(gate96inter4), .b(gate96inter3), .O(gate96inter5));
  nor2  gate1253(.a(gate96inter5), .b(gate96inter2), .O(gate96inter6));
  inv1  gate1254(.a(G30), .O(gate96inter7));
  inv1  gate1255(.a(G347), .O(gate96inter8));
  nand2 gate1256(.a(gate96inter8), .b(gate96inter7), .O(gate96inter9));
  nand2 gate1257(.a(s_101), .b(gate96inter3), .O(gate96inter10));
  nor2  gate1258(.a(gate96inter10), .b(gate96inter9), .O(gate96inter11));
  nor2  gate1259(.a(gate96inter11), .b(gate96inter6), .O(gate96inter12));
  nand2 gate1260(.a(gate96inter12), .b(gate96inter1), .O(G417));

  xor2  gate1947(.a(G350), .b(G19), .O(gate97inter0));
  nand2 gate1948(.a(gate97inter0), .b(s_200), .O(gate97inter1));
  and2  gate1949(.a(G350), .b(G19), .O(gate97inter2));
  inv1  gate1950(.a(s_200), .O(gate97inter3));
  inv1  gate1951(.a(s_201), .O(gate97inter4));
  nand2 gate1952(.a(gate97inter4), .b(gate97inter3), .O(gate97inter5));
  nor2  gate1953(.a(gate97inter5), .b(gate97inter2), .O(gate97inter6));
  inv1  gate1954(.a(G19), .O(gate97inter7));
  inv1  gate1955(.a(G350), .O(gate97inter8));
  nand2 gate1956(.a(gate97inter8), .b(gate97inter7), .O(gate97inter9));
  nand2 gate1957(.a(s_201), .b(gate97inter3), .O(gate97inter10));
  nor2  gate1958(.a(gate97inter10), .b(gate97inter9), .O(gate97inter11));
  nor2  gate1959(.a(gate97inter11), .b(gate97inter6), .O(gate97inter12));
  nand2 gate1960(.a(gate97inter12), .b(gate97inter1), .O(G418));
nand2 gate98( .a(G23), .b(G350), .O(G419) );

  xor2  gate1429(.a(G353), .b(G27), .O(gate99inter0));
  nand2 gate1430(.a(gate99inter0), .b(s_126), .O(gate99inter1));
  and2  gate1431(.a(G353), .b(G27), .O(gate99inter2));
  inv1  gate1432(.a(s_126), .O(gate99inter3));
  inv1  gate1433(.a(s_127), .O(gate99inter4));
  nand2 gate1434(.a(gate99inter4), .b(gate99inter3), .O(gate99inter5));
  nor2  gate1435(.a(gate99inter5), .b(gate99inter2), .O(gate99inter6));
  inv1  gate1436(.a(G27), .O(gate99inter7));
  inv1  gate1437(.a(G353), .O(gate99inter8));
  nand2 gate1438(.a(gate99inter8), .b(gate99inter7), .O(gate99inter9));
  nand2 gate1439(.a(s_127), .b(gate99inter3), .O(gate99inter10));
  nor2  gate1440(.a(gate99inter10), .b(gate99inter9), .O(gate99inter11));
  nor2  gate1441(.a(gate99inter11), .b(gate99inter6), .O(gate99inter12));
  nand2 gate1442(.a(gate99inter12), .b(gate99inter1), .O(G420));
nand2 gate100( .a(G31), .b(G353), .O(G421) );
nand2 gate101( .a(G20), .b(G356), .O(G422) );
nand2 gate102( .a(G24), .b(G356), .O(G423) );
nand2 gate103( .a(G28), .b(G359), .O(G424) );

  xor2  gate911(.a(G359), .b(G32), .O(gate104inter0));
  nand2 gate912(.a(gate104inter0), .b(s_52), .O(gate104inter1));
  and2  gate913(.a(G359), .b(G32), .O(gate104inter2));
  inv1  gate914(.a(s_52), .O(gate104inter3));
  inv1  gate915(.a(s_53), .O(gate104inter4));
  nand2 gate916(.a(gate104inter4), .b(gate104inter3), .O(gate104inter5));
  nor2  gate917(.a(gate104inter5), .b(gate104inter2), .O(gate104inter6));
  inv1  gate918(.a(G32), .O(gate104inter7));
  inv1  gate919(.a(G359), .O(gate104inter8));
  nand2 gate920(.a(gate104inter8), .b(gate104inter7), .O(gate104inter9));
  nand2 gate921(.a(s_53), .b(gate104inter3), .O(gate104inter10));
  nor2  gate922(.a(gate104inter10), .b(gate104inter9), .O(gate104inter11));
  nor2  gate923(.a(gate104inter11), .b(gate104inter6), .O(gate104inter12));
  nand2 gate924(.a(gate104inter12), .b(gate104inter1), .O(G425));
nand2 gate105( .a(G362), .b(G363), .O(G426) );
nand2 gate106( .a(G364), .b(G365), .O(G429) );
nand2 gate107( .a(G366), .b(G367), .O(G432) );
nand2 gate108( .a(G368), .b(G369), .O(G435) );

  xor2  gate1079(.a(G371), .b(G370), .O(gate109inter0));
  nand2 gate1080(.a(gate109inter0), .b(s_76), .O(gate109inter1));
  and2  gate1081(.a(G371), .b(G370), .O(gate109inter2));
  inv1  gate1082(.a(s_76), .O(gate109inter3));
  inv1  gate1083(.a(s_77), .O(gate109inter4));
  nand2 gate1084(.a(gate109inter4), .b(gate109inter3), .O(gate109inter5));
  nor2  gate1085(.a(gate109inter5), .b(gate109inter2), .O(gate109inter6));
  inv1  gate1086(.a(G370), .O(gate109inter7));
  inv1  gate1087(.a(G371), .O(gate109inter8));
  nand2 gate1088(.a(gate109inter8), .b(gate109inter7), .O(gate109inter9));
  nand2 gate1089(.a(s_77), .b(gate109inter3), .O(gate109inter10));
  nor2  gate1090(.a(gate109inter10), .b(gate109inter9), .O(gate109inter11));
  nor2  gate1091(.a(gate109inter11), .b(gate109inter6), .O(gate109inter12));
  nand2 gate1092(.a(gate109inter12), .b(gate109inter1), .O(G438));
nand2 gate110( .a(G372), .b(G373), .O(G441) );
nand2 gate111( .a(G374), .b(G375), .O(G444) );
nand2 gate112( .a(G376), .b(G377), .O(G447) );

  xor2  gate1863(.a(G379), .b(G378), .O(gate113inter0));
  nand2 gate1864(.a(gate113inter0), .b(s_188), .O(gate113inter1));
  and2  gate1865(.a(G379), .b(G378), .O(gate113inter2));
  inv1  gate1866(.a(s_188), .O(gate113inter3));
  inv1  gate1867(.a(s_189), .O(gate113inter4));
  nand2 gate1868(.a(gate113inter4), .b(gate113inter3), .O(gate113inter5));
  nor2  gate1869(.a(gate113inter5), .b(gate113inter2), .O(gate113inter6));
  inv1  gate1870(.a(G378), .O(gate113inter7));
  inv1  gate1871(.a(G379), .O(gate113inter8));
  nand2 gate1872(.a(gate113inter8), .b(gate113inter7), .O(gate113inter9));
  nand2 gate1873(.a(s_189), .b(gate113inter3), .O(gate113inter10));
  nor2  gate1874(.a(gate113inter10), .b(gate113inter9), .O(gate113inter11));
  nor2  gate1875(.a(gate113inter11), .b(gate113inter6), .O(gate113inter12));
  nand2 gate1876(.a(gate113inter12), .b(gate113inter1), .O(G450));
nand2 gate114( .a(G380), .b(G381), .O(G453) );
nand2 gate115( .a(G382), .b(G383), .O(G456) );
nand2 gate116( .a(G384), .b(G385), .O(G459) );

  xor2  gate673(.a(G387), .b(G386), .O(gate117inter0));
  nand2 gate674(.a(gate117inter0), .b(s_18), .O(gate117inter1));
  and2  gate675(.a(G387), .b(G386), .O(gate117inter2));
  inv1  gate676(.a(s_18), .O(gate117inter3));
  inv1  gate677(.a(s_19), .O(gate117inter4));
  nand2 gate678(.a(gate117inter4), .b(gate117inter3), .O(gate117inter5));
  nor2  gate679(.a(gate117inter5), .b(gate117inter2), .O(gate117inter6));
  inv1  gate680(.a(G386), .O(gate117inter7));
  inv1  gate681(.a(G387), .O(gate117inter8));
  nand2 gate682(.a(gate117inter8), .b(gate117inter7), .O(gate117inter9));
  nand2 gate683(.a(s_19), .b(gate117inter3), .O(gate117inter10));
  nor2  gate684(.a(gate117inter10), .b(gate117inter9), .O(gate117inter11));
  nor2  gate685(.a(gate117inter11), .b(gate117inter6), .O(gate117inter12));
  nand2 gate686(.a(gate117inter12), .b(gate117inter1), .O(G462));
nand2 gate118( .a(G388), .b(G389), .O(G465) );
nand2 gate119( .a(G390), .b(G391), .O(G468) );

  xor2  gate1205(.a(G393), .b(G392), .O(gate120inter0));
  nand2 gate1206(.a(gate120inter0), .b(s_94), .O(gate120inter1));
  and2  gate1207(.a(G393), .b(G392), .O(gate120inter2));
  inv1  gate1208(.a(s_94), .O(gate120inter3));
  inv1  gate1209(.a(s_95), .O(gate120inter4));
  nand2 gate1210(.a(gate120inter4), .b(gate120inter3), .O(gate120inter5));
  nor2  gate1211(.a(gate120inter5), .b(gate120inter2), .O(gate120inter6));
  inv1  gate1212(.a(G392), .O(gate120inter7));
  inv1  gate1213(.a(G393), .O(gate120inter8));
  nand2 gate1214(.a(gate120inter8), .b(gate120inter7), .O(gate120inter9));
  nand2 gate1215(.a(s_95), .b(gate120inter3), .O(gate120inter10));
  nor2  gate1216(.a(gate120inter10), .b(gate120inter9), .O(gate120inter11));
  nor2  gate1217(.a(gate120inter11), .b(gate120inter6), .O(gate120inter12));
  nand2 gate1218(.a(gate120inter12), .b(gate120inter1), .O(G471));

  xor2  gate1289(.a(G395), .b(G394), .O(gate121inter0));
  nand2 gate1290(.a(gate121inter0), .b(s_106), .O(gate121inter1));
  and2  gate1291(.a(G395), .b(G394), .O(gate121inter2));
  inv1  gate1292(.a(s_106), .O(gate121inter3));
  inv1  gate1293(.a(s_107), .O(gate121inter4));
  nand2 gate1294(.a(gate121inter4), .b(gate121inter3), .O(gate121inter5));
  nor2  gate1295(.a(gate121inter5), .b(gate121inter2), .O(gate121inter6));
  inv1  gate1296(.a(G394), .O(gate121inter7));
  inv1  gate1297(.a(G395), .O(gate121inter8));
  nand2 gate1298(.a(gate121inter8), .b(gate121inter7), .O(gate121inter9));
  nand2 gate1299(.a(s_107), .b(gate121inter3), .O(gate121inter10));
  nor2  gate1300(.a(gate121inter10), .b(gate121inter9), .O(gate121inter11));
  nor2  gate1301(.a(gate121inter11), .b(gate121inter6), .O(gate121inter12));
  nand2 gate1302(.a(gate121inter12), .b(gate121inter1), .O(G474));

  xor2  gate1485(.a(G397), .b(G396), .O(gate122inter0));
  nand2 gate1486(.a(gate122inter0), .b(s_134), .O(gate122inter1));
  and2  gate1487(.a(G397), .b(G396), .O(gate122inter2));
  inv1  gate1488(.a(s_134), .O(gate122inter3));
  inv1  gate1489(.a(s_135), .O(gate122inter4));
  nand2 gate1490(.a(gate122inter4), .b(gate122inter3), .O(gate122inter5));
  nor2  gate1491(.a(gate122inter5), .b(gate122inter2), .O(gate122inter6));
  inv1  gate1492(.a(G396), .O(gate122inter7));
  inv1  gate1493(.a(G397), .O(gate122inter8));
  nand2 gate1494(.a(gate122inter8), .b(gate122inter7), .O(gate122inter9));
  nand2 gate1495(.a(s_135), .b(gate122inter3), .O(gate122inter10));
  nor2  gate1496(.a(gate122inter10), .b(gate122inter9), .O(gate122inter11));
  nor2  gate1497(.a(gate122inter11), .b(gate122inter6), .O(gate122inter12));
  nand2 gate1498(.a(gate122inter12), .b(gate122inter1), .O(G477));
nand2 gate123( .a(G398), .b(G399), .O(G480) );

  xor2  gate2101(.a(G401), .b(G400), .O(gate124inter0));
  nand2 gate2102(.a(gate124inter0), .b(s_222), .O(gate124inter1));
  and2  gate2103(.a(G401), .b(G400), .O(gate124inter2));
  inv1  gate2104(.a(s_222), .O(gate124inter3));
  inv1  gate2105(.a(s_223), .O(gate124inter4));
  nand2 gate2106(.a(gate124inter4), .b(gate124inter3), .O(gate124inter5));
  nor2  gate2107(.a(gate124inter5), .b(gate124inter2), .O(gate124inter6));
  inv1  gate2108(.a(G400), .O(gate124inter7));
  inv1  gate2109(.a(G401), .O(gate124inter8));
  nand2 gate2110(.a(gate124inter8), .b(gate124inter7), .O(gate124inter9));
  nand2 gate2111(.a(s_223), .b(gate124inter3), .O(gate124inter10));
  nor2  gate2112(.a(gate124inter10), .b(gate124inter9), .O(gate124inter11));
  nor2  gate2113(.a(gate124inter11), .b(gate124inter6), .O(gate124inter12));
  nand2 gate2114(.a(gate124inter12), .b(gate124inter1), .O(G483));

  xor2  gate2227(.a(G403), .b(G402), .O(gate125inter0));
  nand2 gate2228(.a(gate125inter0), .b(s_240), .O(gate125inter1));
  and2  gate2229(.a(G403), .b(G402), .O(gate125inter2));
  inv1  gate2230(.a(s_240), .O(gate125inter3));
  inv1  gate2231(.a(s_241), .O(gate125inter4));
  nand2 gate2232(.a(gate125inter4), .b(gate125inter3), .O(gate125inter5));
  nor2  gate2233(.a(gate125inter5), .b(gate125inter2), .O(gate125inter6));
  inv1  gate2234(.a(G402), .O(gate125inter7));
  inv1  gate2235(.a(G403), .O(gate125inter8));
  nand2 gate2236(.a(gate125inter8), .b(gate125inter7), .O(gate125inter9));
  nand2 gate2237(.a(s_241), .b(gate125inter3), .O(gate125inter10));
  nor2  gate2238(.a(gate125inter10), .b(gate125inter9), .O(gate125inter11));
  nor2  gate2239(.a(gate125inter11), .b(gate125inter6), .O(gate125inter12));
  nand2 gate2240(.a(gate125inter12), .b(gate125inter1), .O(G486));

  xor2  gate1037(.a(G405), .b(G404), .O(gate126inter0));
  nand2 gate1038(.a(gate126inter0), .b(s_70), .O(gate126inter1));
  and2  gate1039(.a(G405), .b(G404), .O(gate126inter2));
  inv1  gate1040(.a(s_70), .O(gate126inter3));
  inv1  gate1041(.a(s_71), .O(gate126inter4));
  nand2 gate1042(.a(gate126inter4), .b(gate126inter3), .O(gate126inter5));
  nor2  gate1043(.a(gate126inter5), .b(gate126inter2), .O(gate126inter6));
  inv1  gate1044(.a(G404), .O(gate126inter7));
  inv1  gate1045(.a(G405), .O(gate126inter8));
  nand2 gate1046(.a(gate126inter8), .b(gate126inter7), .O(gate126inter9));
  nand2 gate1047(.a(s_71), .b(gate126inter3), .O(gate126inter10));
  nor2  gate1048(.a(gate126inter10), .b(gate126inter9), .O(gate126inter11));
  nor2  gate1049(.a(gate126inter11), .b(gate126inter6), .O(gate126inter12));
  nand2 gate1050(.a(gate126inter12), .b(gate126inter1), .O(G489));
nand2 gate127( .a(G406), .b(G407), .O(G492) );
nand2 gate128( .a(G408), .b(G409), .O(G495) );

  xor2  gate1149(.a(G411), .b(G410), .O(gate129inter0));
  nand2 gate1150(.a(gate129inter0), .b(s_86), .O(gate129inter1));
  and2  gate1151(.a(G411), .b(G410), .O(gate129inter2));
  inv1  gate1152(.a(s_86), .O(gate129inter3));
  inv1  gate1153(.a(s_87), .O(gate129inter4));
  nand2 gate1154(.a(gate129inter4), .b(gate129inter3), .O(gate129inter5));
  nor2  gate1155(.a(gate129inter5), .b(gate129inter2), .O(gate129inter6));
  inv1  gate1156(.a(G410), .O(gate129inter7));
  inv1  gate1157(.a(G411), .O(gate129inter8));
  nand2 gate1158(.a(gate129inter8), .b(gate129inter7), .O(gate129inter9));
  nand2 gate1159(.a(s_87), .b(gate129inter3), .O(gate129inter10));
  nor2  gate1160(.a(gate129inter10), .b(gate129inter9), .O(gate129inter11));
  nor2  gate1161(.a(gate129inter11), .b(gate129inter6), .O(gate129inter12));
  nand2 gate1162(.a(gate129inter12), .b(gate129inter1), .O(G498));
nand2 gate130( .a(G412), .b(G413), .O(G501) );

  xor2  gate617(.a(G415), .b(G414), .O(gate131inter0));
  nand2 gate618(.a(gate131inter0), .b(s_10), .O(gate131inter1));
  and2  gate619(.a(G415), .b(G414), .O(gate131inter2));
  inv1  gate620(.a(s_10), .O(gate131inter3));
  inv1  gate621(.a(s_11), .O(gate131inter4));
  nand2 gate622(.a(gate131inter4), .b(gate131inter3), .O(gate131inter5));
  nor2  gate623(.a(gate131inter5), .b(gate131inter2), .O(gate131inter6));
  inv1  gate624(.a(G414), .O(gate131inter7));
  inv1  gate625(.a(G415), .O(gate131inter8));
  nand2 gate626(.a(gate131inter8), .b(gate131inter7), .O(gate131inter9));
  nand2 gate627(.a(s_11), .b(gate131inter3), .O(gate131inter10));
  nor2  gate628(.a(gate131inter10), .b(gate131inter9), .O(gate131inter11));
  nor2  gate629(.a(gate131inter11), .b(gate131inter6), .O(gate131inter12));
  nand2 gate630(.a(gate131inter12), .b(gate131inter1), .O(G504));
nand2 gate132( .a(G416), .b(G417), .O(G507) );
nand2 gate133( .a(G418), .b(G419), .O(G510) );

  xor2  gate2003(.a(G421), .b(G420), .O(gate134inter0));
  nand2 gate2004(.a(gate134inter0), .b(s_208), .O(gate134inter1));
  and2  gate2005(.a(G421), .b(G420), .O(gate134inter2));
  inv1  gate2006(.a(s_208), .O(gate134inter3));
  inv1  gate2007(.a(s_209), .O(gate134inter4));
  nand2 gate2008(.a(gate134inter4), .b(gate134inter3), .O(gate134inter5));
  nor2  gate2009(.a(gate134inter5), .b(gate134inter2), .O(gate134inter6));
  inv1  gate2010(.a(G420), .O(gate134inter7));
  inv1  gate2011(.a(G421), .O(gate134inter8));
  nand2 gate2012(.a(gate134inter8), .b(gate134inter7), .O(gate134inter9));
  nand2 gate2013(.a(s_209), .b(gate134inter3), .O(gate134inter10));
  nor2  gate2014(.a(gate134inter10), .b(gate134inter9), .O(gate134inter11));
  nor2  gate2015(.a(gate134inter11), .b(gate134inter6), .O(gate134inter12));
  nand2 gate2016(.a(gate134inter12), .b(gate134inter1), .O(G513));
nand2 gate135( .a(G422), .b(G423), .O(G516) );
nand2 gate136( .a(G424), .b(G425), .O(G519) );
nand2 gate137( .a(G426), .b(G429), .O(G522) );
nand2 gate138( .a(G432), .b(G435), .O(G525) );
nand2 gate139( .a(G438), .b(G441), .O(G528) );
nand2 gate140( .a(G444), .b(G447), .O(G531) );
nand2 gate141( .a(G450), .b(G453), .O(G534) );
nand2 gate142( .a(G456), .b(G459), .O(G537) );

  xor2  gate743(.a(G465), .b(G462), .O(gate143inter0));
  nand2 gate744(.a(gate143inter0), .b(s_28), .O(gate143inter1));
  and2  gate745(.a(G465), .b(G462), .O(gate143inter2));
  inv1  gate746(.a(s_28), .O(gate143inter3));
  inv1  gate747(.a(s_29), .O(gate143inter4));
  nand2 gate748(.a(gate143inter4), .b(gate143inter3), .O(gate143inter5));
  nor2  gate749(.a(gate143inter5), .b(gate143inter2), .O(gate143inter6));
  inv1  gate750(.a(G462), .O(gate143inter7));
  inv1  gate751(.a(G465), .O(gate143inter8));
  nand2 gate752(.a(gate143inter8), .b(gate143inter7), .O(gate143inter9));
  nand2 gate753(.a(s_29), .b(gate143inter3), .O(gate143inter10));
  nor2  gate754(.a(gate143inter10), .b(gate143inter9), .O(gate143inter11));
  nor2  gate755(.a(gate143inter11), .b(gate143inter6), .O(gate143inter12));
  nand2 gate756(.a(gate143inter12), .b(gate143inter1), .O(G540));
nand2 gate144( .a(G468), .b(G471), .O(G543) );
nand2 gate145( .a(G474), .b(G477), .O(G546) );
nand2 gate146( .a(G480), .b(G483), .O(G549) );
nand2 gate147( .a(G486), .b(G489), .O(G552) );
nand2 gate148( .a(G492), .b(G495), .O(G555) );
nand2 gate149( .a(G498), .b(G501), .O(G558) );
nand2 gate150( .a(G504), .b(G507), .O(G561) );

  xor2  gate897(.a(G513), .b(G510), .O(gate151inter0));
  nand2 gate898(.a(gate151inter0), .b(s_50), .O(gate151inter1));
  and2  gate899(.a(G513), .b(G510), .O(gate151inter2));
  inv1  gate900(.a(s_50), .O(gate151inter3));
  inv1  gate901(.a(s_51), .O(gate151inter4));
  nand2 gate902(.a(gate151inter4), .b(gate151inter3), .O(gate151inter5));
  nor2  gate903(.a(gate151inter5), .b(gate151inter2), .O(gate151inter6));
  inv1  gate904(.a(G510), .O(gate151inter7));
  inv1  gate905(.a(G513), .O(gate151inter8));
  nand2 gate906(.a(gate151inter8), .b(gate151inter7), .O(gate151inter9));
  nand2 gate907(.a(s_51), .b(gate151inter3), .O(gate151inter10));
  nor2  gate908(.a(gate151inter10), .b(gate151inter9), .O(gate151inter11));
  nor2  gate909(.a(gate151inter11), .b(gate151inter6), .O(gate151inter12));
  nand2 gate910(.a(gate151inter12), .b(gate151inter1), .O(G564));
nand2 gate152( .a(G516), .b(G519), .O(G567) );
nand2 gate153( .a(G426), .b(G522), .O(G570) );
nand2 gate154( .a(G429), .b(G522), .O(G571) );
nand2 gate155( .a(G432), .b(G525), .O(G572) );
nand2 gate156( .a(G435), .b(G525), .O(G573) );
nand2 gate157( .a(G438), .b(G528), .O(G574) );
nand2 gate158( .a(G441), .b(G528), .O(G575) );

  xor2  gate1625(.a(G531), .b(G444), .O(gate159inter0));
  nand2 gate1626(.a(gate159inter0), .b(s_154), .O(gate159inter1));
  and2  gate1627(.a(G531), .b(G444), .O(gate159inter2));
  inv1  gate1628(.a(s_154), .O(gate159inter3));
  inv1  gate1629(.a(s_155), .O(gate159inter4));
  nand2 gate1630(.a(gate159inter4), .b(gate159inter3), .O(gate159inter5));
  nor2  gate1631(.a(gate159inter5), .b(gate159inter2), .O(gate159inter6));
  inv1  gate1632(.a(G444), .O(gate159inter7));
  inv1  gate1633(.a(G531), .O(gate159inter8));
  nand2 gate1634(.a(gate159inter8), .b(gate159inter7), .O(gate159inter9));
  nand2 gate1635(.a(s_155), .b(gate159inter3), .O(gate159inter10));
  nor2  gate1636(.a(gate159inter10), .b(gate159inter9), .O(gate159inter11));
  nor2  gate1637(.a(gate159inter11), .b(gate159inter6), .O(gate159inter12));
  nand2 gate1638(.a(gate159inter12), .b(gate159inter1), .O(G576));

  xor2  gate603(.a(G531), .b(G447), .O(gate160inter0));
  nand2 gate604(.a(gate160inter0), .b(s_8), .O(gate160inter1));
  and2  gate605(.a(G531), .b(G447), .O(gate160inter2));
  inv1  gate606(.a(s_8), .O(gate160inter3));
  inv1  gate607(.a(s_9), .O(gate160inter4));
  nand2 gate608(.a(gate160inter4), .b(gate160inter3), .O(gate160inter5));
  nor2  gate609(.a(gate160inter5), .b(gate160inter2), .O(gate160inter6));
  inv1  gate610(.a(G447), .O(gate160inter7));
  inv1  gate611(.a(G531), .O(gate160inter8));
  nand2 gate612(.a(gate160inter8), .b(gate160inter7), .O(gate160inter9));
  nand2 gate613(.a(s_9), .b(gate160inter3), .O(gate160inter10));
  nor2  gate614(.a(gate160inter10), .b(gate160inter9), .O(gate160inter11));
  nor2  gate615(.a(gate160inter11), .b(gate160inter6), .O(gate160inter12));
  nand2 gate616(.a(gate160inter12), .b(gate160inter1), .O(G577));

  xor2  gate1737(.a(G534), .b(G450), .O(gate161inter0));
  nand2 gate1738(.a(gate161inter0), .b(s_170), .O(gate161inter1));
  and2  gate1739(.a(G534), .b(G450), .O(gate161inter2));
  inv1  gate1740(.a(s_170), .O(gate161inter3));
  inv1  gate1741(.a(s_171), .O(gate161inter4));
  nand2 gate1742(.a(gate161inter4), .b(gate161inter3), .O(gate161inter5));
  nor2  gate1743(.a(gate161inter5), .b(gate161inter2), .O(gate161inter6));
  inv1  gate1744(.a(G450), .O(gate161inter7));
  inv1  gate1745(.a(G534), .O(gate161inter8));
  nand2 gate1746(.a(gate161inter8), .b(gate161inter7), .O(gate161inter9));
  nand2 gate1747(.a(s_171), .b(gate161inter3), .O(gate161inter10));
  nor2  gate1748(.a(gate161inter10), .b(gate161inter9), .O(gate161inter11));
  nor2  gate1749(.a(gate161inter11), .b(gate161inter6), .O(gate161inter12));
  nand2 gate1750(.a(gate161inter12), .b(gate161inter1), .O(G578));

  xor2  gate1989(.a(G534), .b(G453), .O(gate162inter0));
  nand2 gate1990(.a(gate162inter0), .b(s_206), .O(gate162inter1));
  and2  gate1991(.a(G534), .b(G453), .O(gate162inter2));
  inv1  gate1992(.a(s_206), .O(gate162inter3));
  inv1  gate1993(.a(s_207), .O(gate162inter4));
  nand2 gate1994(.a(gate162inter4), .b(gate162inter3), .O(gate162inter5));
  nor2  gate1995(.a(gate162inter5), .b(gate162inter2), .O(gate162inter6));
  inv1  gate1996(.a(G453), .O(gate162inter7));
  inv1  gate1997(.a(G534), .O(gate162inter8));
  nand2 gate1998(.a(gate162inter8), .b(gate162inter7), .O(gate162inter9));
  nand2 gate1999(.a(s_207), .b(gate162inter3), .O(gate162inter10));
  nor2  gate2000(.a(gate162inter10), .b(gate162inter9), .O(gate162inter11));
  nor2  gate2001(.a(gate162inter11), .b(gate162inter6), .O(gate162inter12));
  nand2 gate2002(.a(gate162inter12), .b(gate162inter1), .O(G579));
nand2 gate163( .a(G456), .b(G537), .O(G580) );
nand2 gate164( .a(G459), .b(G537), .O(G581) );
nand2 gate165( .a(G462), .b(G540), .O(G582) );

  xor2  gate1765(.a(G540), .b(G465), .O(gate166inter0));
  nand2 gate1766(.a(gate166inter0), .b(s_174), .O(gate166inter1));
  and2  gate1767(.a(G540), .b(G465), .O(gate166inter2));
  inv1  gate1768(.a(s_174), .O(gate166inter3));
  inv1  gate1769(.a(s_175), .O(gate166inter4));
  nand2 gate1770(.a(gate166inter4), .b(gate166inter3), .O(gate166inter5));
  nor2  gate1771(.a(gate166inter5), .b(gate166inter2), .O(gate166inter6));
  inv1  gate1772(.a(G465), .O(gate166inter7));
  inv1  gate1773(.a(G540), .O(gate166inter8));
  nand2 gate1774(.a(gate166inter8), .b(gate166inter7), .O(gate166inter9));
  nand2 gate1775(.a(s_175), .b(gate166inter3), .O(gate166inter10));
  nor2  gate1776(.a(gate166inter10), .b(gate166inter9), .O(gate166inter11));
  nor2  gate1777(.a(gate166inter11), .b(gate166inter6), .O(gate166inter12));
  nand2 gate1778(.a(gate166inter12), .b(gate166inter1), .O(G583));
nand2 gate167( .a(G468), .b(G543), .O(G584) );
nand2 gate168( .a(G471), .b(G543), .O(G585) );

  xor2  gate995(.a(G546), .b(G474), .O(gate169inter0));
  nand2 gate996(.a(gate169inter0), .b(s_64), .O(gate169inter1));
  and2  gate997(.a(G546), .b(G474), .O(gate169inter2));
  inv1  gate998(.a(s_64), .O(gate169inter3));
  inv1  gate999(.a(s_65), .O(gate169inter4));
  nand2 gate1000(.a(gate169inter4), .b(gate169inter3), .O(gate169inter5));
  nor2  gate1001(.a(gate169inter5), .b(gate169inter2), .O(gate169inter6));
  inv1  gate1002(.a(G474), .O(gate169inter7));
  inv1  gate1003(.a(G546), .O(gate169inter8));
  nand2 gate1004(.a(gate169inter8), .b(gate169inter7), .O(gate169inter9));
  nand2 gate1005(.a(s_65), .b(gate169inter3), .O(gate169inter10));
  nor2  gate1006(.a(gate169inter10), .b(gate169inter9), .O(gate169inter11));
  nor2  gate1007(.a(gate169inter11), .b(gate169inter6), .O(gate169inter12));
  nand2 gate1008(.a(gate169inter12), .b(gate169inter1), .O(G586));

  xor2  gate1345(.a(G546), .b(G477), .O(gate170inter0));
  nand2 gate1346(.a(gate170inter0), .b(s_114), .O(gate170inter1));
  and2  gate1347(.a(G546), .b(G477), .O(gate170inter2));
  inv1  gate1348(.a(s_114), .O(gate170inter3));
  inv1  gate1349(.a(s_115), .O(gate170inter4));
  nand2 gate1350(.a(gate170inter4), .b(gate170inter3), .O(gate170inter5));
  nor2  gate1351(.a(gate170inter5), .b(gate170inter2), .O(gate170inter6));
  inv1  gate1352(.a(G477), .O(gate170inter7));
  inv1  gate1353(.a(G546), .O(gate170inter8));
  nand2 gate1354(.a(gate170inter8), .b(gate170inter7), .O(gate170inter9));
  nand2 gate1355(.a(s_115), .b(gate170inter3), .O(gate170inter10));
  nor2  gate1356(.a(gate170inter10), .b(gate170inter9), .O(gate170inter11));
  nor2  gate1357(.a(gate170inter11), .b(gate170inter6), .O(gate170inter12));
  nand2 gate1358(.a(gate170inter12), .b(gate170inter1), .O(G587));
nand2 gate171( .a(G480), .b(G549), .O(G588) );

  xor2  gate1667(.a(G549), .b(G483), .O(gate172inter0));
  nand2 gate1668(.a(gate172inter0), .b(s_160), .O(gate172inter1));
  and2  gate1669(.a(G549), .b(G483), .O(gate172inter2));
  inv1  gate1670(.a(s_160), .O(gate172inter3));
  inv1  gate1671(.a(s_161), .O(gate172inter4));
  nand2 gate1672(.a(gate172inter4), .b(gate172inter3), .O(gate172inter5));
  nor2  gate1673(.a(gate172inter5), .b(gate172inter2), .O(gate172inter6));
  inv1  gate1674(.a(G483), .O(gate172inter7));
  inv1  gate1675(.a(G549), .O(gate172inter8));
  nand2 gate1676(.a(gate172inter8), .b(gate172inter7), .O(gate172inter9));
  nand2 gate1677(.a(s_161), .b(gate172inter3), .O(gate172inter10));
  nor2  gate1678(.a(gate172inter10), .b(gate172inter9), .O(gate172inter11));
  nor2  gate1679(.a(gate172inter11), .b(gate172inter6), .O(gate172inter12));
  nand2 gate1680(.a(gate172inter12), .b(gate172inter1), .O(G589));
nand2 gate173( .a(G486), .b(G552), .O(G590) );
nand2 gate174( .a(G489), .b(G552), .O(G591) );

  xor2  gate1821(.a(G555), .b(G492), .O(gate175inter0));
  nand2 gate1822(.a(gate175inter0), .b(s_182), .O(gate175inter1));
  and2  gate1823(.a(G555), .b(G492), .O(gate175inter2));
  inv1  gate1824(.a(s_182), .O(gate175inter3));
  inv1  gate1825(.a(s_183), .O(gate175inter4));
  nand2 gate1826(.a(gate175inter4), .b(gate175inter3), .O(gate175inter5));
  nor2  gate1827(.a(gate175inter5), .b(gate175inter2), .O(gate175inter6));
  inv1  gate1828(.a(G492), .O(gate175inter7));
  inv1  gate1829(.a(G555), .O(gate175inter8));
  nand2 gate1830(.a(gate175inter8), .b(gate175inter7), .O(gate175inter9));
  nand2 gate1831(.a(s_183), .b(gate175inter3), .O(gate175inter10));
  nor2  gate1832(.a(gate175inter10), .b(gate175inter9), .O(gate175inter11));
  nor2  gate1833(.a(gate175inter11), .b(gate175inter6), .O(gate175inter12));
  nand2 gate1834(.a(gate175inter12), .b(gate175inter1), .O(G592));
nand2 gate176( .a(G495), .b(G555), .O(G593) );
nand2 gate177( .a(G498), .b(G558), .O(G594) );
nand2 gate178( .a(G501), .b(G558), .O(G595) );

  xor2  gate2059(.a(G561), .b(G504), .O(gate179inter0));
  nand2 gate2060(.a(gate179inter0), .b(s_216), .O(gate179inter1));
  and2  gate2061(.a(G561), .b(G504), .O(gate179inter2));
  inv1  gate2062(.a(s_216), .O(gate179inter3));
  inv1  gate2063(.a(s_217), .O(gate179inter4));
  nand2 gate2064(.a(gate179inter4), .b(gate179inter3), .O(gate179inter5));
  nor2  gate2065(.a(gate179inter5), .b(gate179inter2), .O(gate179inter6));
  inv1  gate2066(.a(G504), .O(gate179inter7));
  inv1  gate2067(.a(G561), .O(gate179inter8));
  nand2 gate2068(.a(gate179inter8), .b(gate179inter7), .O(gate179inter9));
  nand2 gate2069(.a(s_217), .b(gate179inter3), .O(gate179inter10));
  nor2  gate2070(.a(gate179inter10), .b(gate179inter9), .O(gate179inter11));
  nor2  gate2071(.a(gate179inter11), .b(gate179inter6), .O(gate179inter12));
  nand2 gate2072(.a(gate179inter12), .b(gate179inter1), .O(G596));
nand2 gate180( .a(G507), .b(G561), .O(G597) );

  xor2  gate1373(.a(G564), .b(G510), .O(gate181inter0));
  nand2 gate1374(.a(gate181inter0), .b(s_118), .O(gate181inter1));
  and2  gate1375(.a(G564), .b(G510), .O(gate181inter2));
  inv1  gate1376(.a(s_118), .O(gate181inter3));
  inv1  gate1377(.a(s_119), .O(gate181inter4));
  nand2 gate1378(.a(gate181inter4), .b(gate181inter3), .O(gate181inter5));
  nor2  gate1379(.a(gate181inter5), .b(gate181inter2), .O(gate181inter6));
  inv1  gate1380(.a(G510), .O(gate181inter7));
  inv1  gate1381(.a(G564), .O(gate181inter8));
  nand2 gate1382(.a(gate181inter8), .b(gate181inter7), .O(gate181inter9));
  nand2 gate1383(.a(s_119), .b(gate181inter3), .O(gate181inter10));
  nor2  gate1384(.a(gate181inter10), .b(gate181inter9), .O(gate181inter11));
  nor2  gate1385(.a(gate181inter11), .b(gate181inter6), .O(gate181inter12));
  nand2 gate1386(.a(gate181inter12), .b(gate181inter1), .O(G598));
nand2 gate182( .a(G513), .b(G564), .O(G599) );
nand2 gate183( .a(G516), .b(G567), .O(G600) );
nand2 gate184( .a(G519), .b(G567), .O(G601) );
nand2 gate185( .a(G570), .b(G571), .O(G602) );

  xor2  gate1163(.a(G573), .b(G572), .O(gate186inter0));
  nand2 gate1164(.a(gate186inter0), .b(s_88), .O(gate186inter1));
  and2  gate1165(.a(G573), .b(G572), .O(gate186inter2));
  inv1  gate1166(.a(s_88), .O(gate186inter3));
  inv1  gate1167(.a(s_89), .O(gate186inter4));
  nand2 gate1168(.a(gate186inter4), .b(gate186inter3), .O(gate186inter5));
  nor2  gate1169(.a(gate186inter5), .b(gate186inter2), .O(gate186inter6));
  inv1  gate1170(.a(G572), .O(gate186inter7));
  inv1  gate1171(.a(G573), .O(gate186inter8));
  nand2 gate1172(.a(gate186inter8), .b(gate186inter7), .O(gate186inter9));
  nand2 gate1173(.a(s_89), .b(gate186inter3), .O(gate186inter10));
  nor2  gate1174(.a(gate186inter10), .b(gate186inter9), .O(gate186inter11));
  nor2  gate1175(.a(gate186inter11), .b(gate186inter6), .O(gate186inter12));
  nand2 gate1176(.a(gate186inter12), .b(gate186inter1), .O(G607));

  xor2  gate1121(.a(G575), .b(G574), .O(gate187inter0));
  nand2 gate1122(.a(gate187inter0), .b(s_82), .O(gate187inter1));
  and2  gate1123(.a(G575), .b(G574), .O(gate187inter2));
  inv1  gate1124(.a(s_82), .O(gate187inter3));
  inv1  gate1125(.a(s_83), .O(gate187inter4));
  nand2 gate1126(.a(gate187inter4), .b(gate187inter3), .O(gate187inter5));
  nor2  gate1127(.a(gate187inter5), .b(gate187inter2), .O(gate187inter6));
  inv1  gate1128(.a(G574), .O(gate187inter7));
  inv1  gate1129(.a(G575), .O(gate187inter8));
  nand2 gate1130(.a(gate187inter8), .b(gate187inter7), .O(gate187inter9));
  nand2 gate1131(.a(s_83), .b(gate187inter3), .O(gate187inter10));
  nor2  gate1132(.a(gate187inter10), .b(gate187inter9), .O(gate187inter11));
  nor2  gate1133(.a(gate187inter11), .b(gate187inter6), .O(gate187inter12));
  nand2 gate1134(.a(gate187inter12), .b(gate187inter1), .O(G612));

  xor2  gate1233(.a(G577), .b(G576), .O(gate188inter0));
  nand2 gate1234(.a(gate188inter0), .b(s_98), .O(gate188inter1));
  and2  gate1235(.a(G577), .b(G576), .O(gate188inter2));
  inv1  gate1236(.a(s_98), .O(gate188inter3));
  inv1  gate1237(.a(s_99), .O(gate188inter4));
  nand2 gate1238(.a(gate188inter4), .b(gate188inter3), .O(gate188inter5));
  nor2  gate1239(.a(gate188inter5), .b(gate188inter2), .O(gate188inter6));
  inv1  gate1240(.a(G576), .O(gate188inter7));
  inv1  gate1241(.a(G577), .O(gate188inter8));
  nand2 gate1242(.a(gate188inter8), .b(gate188inter7), .O(gate188inter9));
  nand2 gate1243(.a(s_99), .b(gate188inter3), .O(gate188inter10));
  nor2  gate1244(.a(gate188inter10), .b(gate188inter9), .O(gate188inter11));
  nor2  gate1245(.a(gate188inter11), .b(gate188inter6), .O(gate188inter12));
  nand2 gate1246(.a(gate188inter12), .b(gate188inter1), .O(G617));
nand2 gate189( .a(G578), .b(G579), .O(G622) );

  xor2  gate799(.a(G581), .b(G580), .O(gate190inter0));
  nand2 gate800(.a(gate190inter0), .b(s_36), .O(gate190inter1));
  and2  gate801(.a(G581), .b(G580), .O(gate190inter2));
  inv1  gate802(.a(s_36), .O(gate190inter3));
  inv1  gate803(.a(s_37), .O(gate190inter4));
  nand2 gate804(.a(gate190inter4), .b(gate190inter3), .O(gate190inter5));
  nor2  gate805(.a(gate190inter5), .b(gate190inter2), .O(gate190inter6));
  inv1  gate806(.a(G580), .O(gate190inter7));
  inv1  gate807(.a(G581), .O(gate190inter8));
  nand2 gate808(.a(gate190inter8), .b(gate190inter7), .O(gate190inter9));
  nand2 gate809(.a(s_37), .b(gate190inter3), .O(gate190inter10));
  nor2  gate810(.a(gate190inter10), .b(gate190inter9), .O(gate190inter11));
  nor2  gate811(.a(gate190inter11), .b(gate190inter6), .O(gate190inter12));
  nand2 gate812(.a(gate190inter12), .b(gate190inter1), .O(G627));
nand2 gate191( .a(G582), .b(G583), .O(G632) );
nand2 gate192( .a(G584), .b(G585), .O(G637) );
nand2 gate193( .a(G586), .b(G587), .O(G642) );
nand2 gate194( .a(G588), .b(G589), .O(G645) );
nand2 gate195( .a(G590), .b(G591), .O(G648) );
nand2 gate196( .a(G592), .b(G593), .O(G651) );
nand2 gate197( .a(G594), .b(G595), .O(G654) );
nand2 gate198( .a(G596), .b(G597), .O(G657) );
nand2 gate199( .a(G598), .b(G599), .O(G660) );
nand2 gate200( .a(G600), .b(G601), .O(G663) );

  xor2  gate645(.a(G607), .b(G602), .O(gate201inter0));
  nand2 gate646(.a(gate201inter0), .b(s_14), .O(gate201inter1));
  and2  gate647(.a(G607), .b(G602), .O(gate201inter2));
  inv1  gate648(.a(s_14), .O(gate201inter3));
  inv1  gate649(.a(s_15), .O(gate201inter4));
  nand2 gate650(.a(gate201inter4), .b(gate201inter3), .O(gate201inter5));
  nor2  gate651(.a(gate201inter5), .b(gate201inter2), .O(gate201inter6));
  inv1  gate652(.a(G602), .O(gate201inter7));
  inv1  gate653(.a(G607), .O(gate201inter8));
  nand2 gate654(.a(gate201inter8), .b(gate201inter7), .O(gate201inter9));
  nand2 gate655(.a(s_15), .b(gate201inter3), .O(gate201inter10));
  nor2  gate656(.a(gate201inter10), .b(gate201inter9), .O(gate201inter11));
  nor2  gate657(.a(gate201inter11), .b(gate201inter6), .O(gate201inter12));
  nand2 gate658(.a(gate201inter12), .b(gate201inter1), .O(G666));

  xor2  gate1401(.a(G617), .b(G612), .O(gate202inter0));
  nand2 gate1402(.a(gate202inter0), .b(s_122), .O(gate202inter1));
  and2  gate1403(.a(G617), .b(G612), .O(gate202inter2));
  inv1  gate1404(.a(s_122), .O(gate202inter3));
  inv1  gate1405(.a(s_123), .O(gate202inter4));
  nand2 gate1406(.a(gate202inter4), .b(gate202inter3), .O(gate202inter5));
  nor2  gate1407(.a(gate202inter5), .b(gate202inter2), .O(gate202inter6));
  inv1  gate1408(.a(G612), .O(gate202inter7));
  inv1  gate1409(.a(G617), .O(gate202inter8));
  nand2 gate1410(.a(gate202inter8), .b(gate202inter7), .O(gate202inter9));
  nand2 gate1411(.a(s_123), .b(gate202inter3), .O(gate202inter10));
  nor2  gate1412(.a(gate202inter10), .b(gate202inter9), .O(gate202inter11));
  nor2  gate1413(.a(gate202inter11), .b(gate202inter6), .O(gate202inter12));
  nand2 gate1414(.a(gate202inter12), .b(gate202inter1), .O(G669));

  xor2  gate813(.a(G612), .b(G602), .O(gate203inter0));
  nand2 gate814(.a(gate203inter0), .b(s_38), .O(gate203inter1));
  and2  gate815(.a(G612), .b(G602), .O(gate203inter2));
  inv1  gate816(.a(s_38), .O(gate203inter3));
  inv1  gate817(.a(s_39), .O(gate203inter4));
  nand2 gate818(.a(gate203inter4), .b(gate203inter3), .O(gate203inter5));
  nor2  gate819(.a(gate203inter5), .b(gate203inter2), .O(gate203inter6));
  inv1  gate820(.a(G602), .O(gate203inter7));
  inv1  gate821(.a(G612), .O(gate203inter8));
  nand2 gate822(.a(gate203inter8), .b(gate203inter7), .O(gate203inter9));
  nand2 gate823(.a(s_39), .b(gate203inter3), .O(gate203inter10));
  nor2  gate824(.a(gate203inter10), .b(gate203inter9), .O(gate203inter11));
  nor2  gate825(.a(gate203inter11), .b(gate203inter6), .O(gate203inter12));
  nand2 gate826(.a(gate203inter12), .b(gate203inter1), .O(G672));
nand2 gate204( .a(G607), .b(G617), .O(G675) );
nand2 gate205( .a(G622), .b(G627), .O(G678) );

  xor2  gate1555(.a(G637), .b(G632), .O(gate206inter0));
  nand2 gate1556(.a(gate206inter0), .b(s_144), .O(gate206inter1));
  and2  gate1557(.a(G637), .b(G632), .O(gate206inter2));
  inv1  gate1558(.a(s_144), .O(gate206inter3));
  inv1  gate1559(.a(s_145), .O(gate206inter4));
  nand2 gate1560(.a(gate206inter4), .b(gate206inter3), .O(gate206inter5));
  nor2  gate1561(.a(gate206inter5), .b(gate206inter2), .O(gate206inter6));
  inv1  gate1562(.a(G632), .O(gate206inter7));
  inv1  gate1563(.a(G637), .O(gate206inter8));
  nand2 gate1564(.a(gate206inter8), .b(gate206inter7), .O(gate206inter9));
  nand2 gate1565(.a(s_145), .b(gate206inter3), .O(gate206inter10));
  nor2  gate1566(.a(gate206inter10), .b(gate206inter9), .O(gate206inter11));
  nor2  gate1567(.a(gate206inter11), .b(gate206inter6), .O(gate206inter12));
  nand2 gate1568(.a(gate206inter12), .b(gate206inter1), .O(G681));
nand2 gate207( .a(G622), .b(G632), .O(G684) );
nand2 gate208( .a(G627), .b(G637), .O(G687) );
nand2 gate209( .a(G602), .b(G666), .O(G690) );
nand2 gate210( .a(G607), .b(G666), .O(G691) );
nand2 gate211( .a(G612), .b(G669), .O(G692) );
nand2 gate212( .a(G617), .b(G669), .O(G693) );
nand2 gate213( .a(G602), .b(G672), .O(G694) );
nand2 gate214( .a(G612), .b(G672), .O(G695) );

  xor2  gate1681(.a(G675), .b(G607), .O(gate215inter0));
  nand2 gate1682(.a(gate215inter0), .b(s_162), .O(gate215inter1));
  and2  gate1683(.a(G675), .b(G607), .O(gate215inter2));
  inv1  gate1684(.a(s_162), .O(gate215inter3));
  inv1  gate1685(.a(s_163), .O(gate215inter4));
  nand2 gate1686(.a(gate215inter4), .b(gate215inter3), .O(gate215inter5));
  nor2  gate1687(.a(gate215inter5), .b(gate215inter2), .O(gate215inter6));
  inv1  gate1688(.a(G607), .O(gate215inter7));
  inv1  gate1689(.a(G675), .O(gate215inter8));
  nand2 gate1690(.a(gate215inter8), .b(gate215inter7), .O(gate215inter9));
  nand2 gate1691(.a(s_163), .b(gate215inter3), .O(gate215inter10));
  nor2  gate1692(.a(gate215inter10), .b(gate215inter9), .O(gate215inter11));
  nor2  gate1693(.a(gate215inter11), .b(gate215inter6), .O(gate215inter12));
  nand2 gate1694(.a(gate215inter12), .b(gate215inter1), .O(G696));
nand2 gate216( .a(G617), .b(G675), .O(G697) );
nand2 gate217( .a(G622), .b(G678), .O(G698) );
nand2 gate218( .a(G627), .b(G678), .O(G699) );
nand2 gate219( .a(G632), .b(G681), .O(G700) );

  xor2  gate1597(.a(G681), .b(G637), .O(gate220inter0));
  nand2 gate1598(.a(gate220inter0), .b(s_150), .O(gate220inter1));
  and2  gate1599(.a(G681), .b(G637), .O(gate220inter2));
  inv1  gate1600(.a(s_150), .O(gate220inter3));
  inv1  gate1601(.a(s_151), .O(gate220inter4));
  nand2 gate1602(.a(gate220inter4), .b(gate220inter3), .O(gate220inter5));
  nor2  gate1603(.a(gate220inter5), .b(gate220inter2), .O(gate220inter6));
  inv1  gate1604(.a(G637), .O(gate220inter7));
  inv1  gate1605(.a(G681), .O(gate220inter8));
  nand2 gate1606(.a(gate220inter8), .b(gate220inter7), .O(gate220inter9));
  nand2 gate1607(.a(s_151), .b(gate220inter3), .O(gate220inter10));
  nor2  gate1608(.a(gate220inter10), .b(gate220inter9), .O(gate220inter11));
  nor2  gate1609(.a(gate220inter11), .b(gate220inter6), .O(gate220inter12));
  nand2 gate1610(.a(gate220inter12), .b(gate220inter1), .O(G701));
nand2 gate221( .a(G622), .b(G684), .O(G702) );
nand2 gate222( .a(G632), .b(G684), .O(G703) );
nand2 gate223( .a(G627), .b(G687), .O(G704) );
nand2 gate224( .a(G637), .b(G687), .O(G705) );
nand2 gate225( .a(G690), .b(G691), .O(G706) );
nand2 gate226( .a(G692), .b(G693), .O(G709) );
nand2 gate227( .a(G694), .b(G695), .O(G712) );
nand2 gate228( .a(G696), .b(G697), .O(G715) );
nand2 gate229( .a(G698), .b(G699), .O(G718) );

  xor2  gate757(.a(G701), .b(G700), .O(gate230inter0));
  nand2 gate758(.a(gate230inter0), .b(s_30), .O(gate230inter1));
  and2  gate759(.a(G701), .b(G700), .O(gate230inter2));
  inv1  gate760(.a(s_30), .O(gate230inter3));
  inv1  gate761(.a(s_31), .O(gate230inter4));
  nand2 gate762(.a(gate230inter4), .b(gate230inter3), .O(gate230inter5));
  nor2  gate763(.a(gate230inter5), .b(gate230inter2), .O(gate230inter6));
  inv1  gate764(.a(G700), .O(gate230inter7));
  inv1  gate765(.a(G701), .O(gate230inter8));
  nand2 gate766(.a(gate230inter8), .b(gate230inter7), .O(gate230inter9));
  nand2 gate767(.a(s_31), .b(gate230inter3), .O(gate230inter10));
  nor2  gate768(.a(gate230inter10), .b(gate230inter9), .O(gate230inter11));
  nor2  gate769(.a(gate230inter11), .b(gate230inter6), .O(gate230inter12));
  nand2 gate770(.a(gate230inter12), .b(gate230inter1), .O(G721));

  xor2  gate561(.a(G703), .b(G702), .O(gate231inter0));
  nand2 gate562(.a(gate231inter0), .b(s_2), .O(gate231inter1));
  and2  gate563(.a(G703), .b(G702), .O(gate231inter2));
  inv1  gate564(.a(s_2), .O(gate231inter3));
  inv1  gate565(.a(s_3), .O(gate231inter4));
  nand2 gate566(.a(gate231inter4), .b(gate231inter3), .O(gate231inter5));
  nor2  gate567(.a(gate231inter5), .b(gate231inter2), .O(gate231inter6));
  inv1  gate568(.a(G702), .O(gate231inter7));
  inv1  gate569(.a(G703), .O(gate231inter8));
  nand2 gate570(.a(gate231inter8), .b(gate231inter7), .O(gate231inter9));
  nand2 gate571(.a(s_3), .b(gate231inter3), .O(gate231inter10));
  nor2  gate572(.a(gate231inter10), .b(gate231inter9), .O(gate231inter11));
  nor2  gate573(.a(gate231inter11), .b(gate231inter6), .O(gate231inter12));
  nand2 gate574(.a(gate231inter12), .b(gate231inter1), .O(G724));
nand2 gate232( .a(G704), .b(G705), .O(G727) );

  xor2  gate1261(.a(G718), .b(G242), .O(gate233inter0));
  nand2 gate1262(.a(gate233inter0), .b(s_102), .O(gate233inter1));
  and2  gate1263(.a(G718), .b(G242), .O(gate233inter2));
  inv1  gate1264(.a(s_102), .O(gate233inter3));
  inv1  gate1265(.a(s_103), .O(gate233inter4));
  nand2 gate1266(.a(gate233inter4), .b(gate233inter3), .O(gate233inter5));
  nor2  gate1267(.a(gate233inter5), .b(gate233inter2), .O(gate233inter6));
  inv1  gate1268(.a(G242), .O(gate233inter7));
  inv1  gate1269(.a(G718), .O(gate233inter8));
  nand2 gate1270(.a(gate233inter8), .b(gate233inter7), .O(gate233inter9));
  nand2 gate1271(.a(s_103), .b(gate233inter3), .O(gate233inter10));
  nor2  gate1272(.a(gate233inter10), .b(gate233inter9), .O(gate233inter11));
  nor2  gate1273(.a(gate233inter11), .b(gate233inter6), .O(gate233inter12));
  nand2 gate1274(.a(gate233inter12), .b(gate233inter1), .O(G730));
nand2 gate234( .a(G245), .b(G721), .O(G733) );
nand2 gate235( .a(G248), .b(G724), .O(G736) );
nand2 gate236( .a(G251), .b(G727), .O(G739) );
nand2 gate237( .a(G254), .b(G706), .O(G742) );
nand2 gate238( .a(G257), .b(G709), .O(G745) );
nand2 gate239( .a(G260), .b(G712), .O(G748) );

  xor2  gate1723(.a(G715), .b(G263), .O(gate240inter0));
  nand2 gate1724(.a(gate240inter0), .b(s_168), .O(gate240inter1));
  and2  gate1725(.a(G715), .b(G263), .O(gate240inter2));
  inv1  gate1726(.a(s_168), .O(gate240inter3));
  inv1  gate1727(.a(s_169), .O(gate240inter4));
  nand2 gate1728(.a(gate240inter4), .b(gate240inter3), .O(gate240inter5));
  nor2  gate1729(.a(gate240inter5), .b(gate240inter2), .O(gate240inter6));
  inv1  gate1730(.a(G263), .O(gate240inter7));
  inv1  gate1731(.a(G715), .O(gate240inter8));
  nand2 gate1732(.a(gate240inter8), .b(gate240inter7), .O(gate240inter9));
  nand2 gate1733(.a(s_169), .b(gate240inter3), .O(gate240inter10));
  nor2  gate1734(.a(gate240inter10), .b(gate240inter9), .O(gate240inter11));
  nor2  gate1735(.a(gate240inter11), .b(gate240inter6), .O(gate240inter12));
  nand2 gate1736(.a(gate240inter12), .b(gate240inter1), .O(G751));
nand2 gate241( .a(G242), .b(G730), .O(G754) );
nand2 gate242( .a(G718), .b(G730), .O(G755) );
nand2 gate243( .a(G245), .b(G733), .O(G756) );
nand2 gate244( .a(G721), .b(G733), .O(G757) );
nand2 gate245( .a(G248), .b(G736), .O(G758) );
nand2 gate246( .a(G724), .b(G736), .O(G759) );
nand2 gate247( .a(G251), .b(G739), .O(G760) );
nand2 gate248( .a(G727), .b(G739), .O(G761) );

  xor2  gate1387(.a(G742), .b(G254), .O(gate249inter0));
  nand2 gate1388(.a(gate249inter0), .b(s_120), .O(gate249inter1));
  and2  gate1389(.a(G742), .b(G254), .O(gate249inter2));
  inv1  gate1390(.a(s_120), .O(gate249inter3));
  inv1  gate1391(.a(s_121), .O(gate249inter4));
  nand2 gate1392(.a(gate249inter4), .b(gate249inter3), .O(gate249inter5));
  nor2  gate1393(.a(gate249inter5), .b(gate249inter2), .O(gate249inter6));
  inv1  gate1394(.a(G254), .O(gate249inter7));
  inv1  gate1395(.a(G742), .O(gate249inter8));
  nand2 gate1396(.a(gate249inter8), .b(gate249inter7), .O(gate249inter9));
  nand2 gate1397(.a(s_121), .b(gate249inter3), .O(gate249inter10));
  nor2  gate1398(.a(gate249inter10), .b(gate249inter9), .O(gate249inter11));
  nor2  gate1399(.a(gate249inter11), .b(gate249inter6), .O(gate249inter12));
  nand2 gate1400(.a(gate249inter12), .b(gate249inter1), .O(G762));
nand2 gate250( .a(G706), .b(G742), .O(G763) );

  xor2  gate883(.a(G745), .b(G257), .O(gate251inter0));
  nand2 gate884(.a(gate251inter0), .b(s_48), .O(gate251inter1));
  and2  gate885(.a(G745), .b(G257), .O(gate251inter2));
  inv1  gate886(.a(s_48), .O(gate251inter3));
  inv1  gate887(.a(s_49), .O(gate251inter4));
  nand2 gate888(.a(gate251inter4), .b(gate251inter3), .O(gate251inter5));
  nor2  gate889(.a(gate251inter5), .b(gate251inter2), .O(gate251inter6));
  inv1  gate890(.a(G257), .O(gate251inter7));
  inv1  gate891(.a(G745), .O(gate251inter8));
  nand2 gate892(.a(gate251inter8), .b(gate251inter7), .O(gate251inter9));
  nand2 gate893(.a(s_49), .b(gate251inter3), .O(gate251inter10));
  nor2  gate894(.a(gate251inter10), .b(gate251inter9), .O(gate251inter11));
  nor2  gate895(.a(gate251inter11), .b(gate251inter6), .O(gate251inter12));
  nand2 gate896(.a(gate251inter12), .b(gate251inter1), .O(G764));
nand2 gate252( .a(G709), .b(G745), .O(G765) );

  xor2  gate1191(.a(G748), .b(G260), .O(gate253inter0));
  nand2 gate1192(.a(gate253inter0), .b(s_92), .O(gate253inter1));
  and2  gate1193(.a(G748), .b(G260), .O(gate253inter2));
  inv1  gate1194(.a(s_92), .O(gate253inter3));
  inv1  gate1195(.a(s_93), .O(gate253inter4));
  nand2 gate1196(.a(gate253inter4), .b(gate253inter3), .O(gate253inter5));
  nor2  gate1197(.a(gate253inter5), .b(gate253inter2), .O(gate253inter6));
  inv1  gate1198(.a(G260), .O(gate253inter7));
  inv1  gate1199(.a(G748), .O(gate253inter8));
  nand2 gate1200(.a(gate253inter8), .b(gate253inter7), .O(gate253inter9));
  nand2 gate1201(.a(s_93), .b(gate253inter3), .O(gate253inter10));
  nor2  gate1202(.a(gate253inter10), .b(gate253inter9), .O(gate253inter11));
  nor2  gate1203(.a(gate253inter11), .b(gate253inter6), .O(gate253inter12));
  nand2 gate1204(.a(gate253inter12), .b(gate253inter1), .O(G766));
nand2 gate254( .a(G712), .b(G748), .O(G767) );
nand2 gate255( .a(G263), .b(G751), .O(G768) );
nand2 gate256( .a(G715), .b(G751), .O(G769) );

  xor2  gate1793(.a(G755), .b(G754), .O(gate257inter0));
  nand2 gate1794(.a(gate257inter0), .b(s_178), .O(gate257inter1));
  and2  gate1795(.a(G755), .b(G754), .O(gate257inter2));
  inv1  gate1796(.a(s_178), .O(gate257inter3));
  inv1  gate1797(.a(s_179), .O(gate257inter4));
  nand2 gate1798(.a(gate257inter4), .b(gate257inter3), .O(gate257inter5));
  nor2  gate1799(.a(gate257inter5), .b(gate257inter2), .O(gate257inter6));
  inv1  gate1800(.a(G754), .O(gate257inter7));
  inv1  gate1801(.a(G755), .O(gate257inter8));
  nand2 gate1802(.a(gate257inter8), .b(gate257inter7), .O(gate257inter9));
  nand2 gate1803(.a(s_179), .b(gate257inter3), .O(gate257inter10));
  nor2  gate1804(.a(gate257inter10), .b(gate257inter9), .O(gate257inter11));
  nor2  gate1805(.a(gate257inter11), .b(gate257inter6), .O(gate257inter12));
  nand2 gate1806(.a(gate257inter12), .b(gate257inter1), .O(G770));
nand2 gate258( .a(G756), .b(G757), .O(G773) );
nand2 gate259( .a(G758), .b(G759), .O(G776) );
nand2 gate260( .a(G760), .b(G761), .O(G779) );

  xor2  gate1415(.a(G763), .b(G762), .O(gate261inter0));
  nand2 gate1416(.a(gate261inter0), .b(s_124), .O(gate261inter1));
  and2  gate1417(.a(G763), .b(G762), .O(gate261inter2));
  inv1  gate1418(.a(s_124), .O(gate261inter3));
  inv1  gate1419(.a(s_125), .O(gate261inter4));
  nand2 gate1420(.a(gate261inter4), .b(gate261inter3), .O(gate261inter5));
  nor2  gate1421(.a(gate261inter5), .b(gate261inter2), .O(gate261inter6));
  inv1  gate1422(.a(G762), .O(gate261inter7));
  inv1  gate1423(.a(G763), .O(gate261inter8));
  nand2 gate1424(.a(gate261inter8), .b(gate261inter7), .O(gate261inter9));
  nand2 gate1425(.a(s_125), .b(gate261inter3), .O(gate261inter10));
  nor2  gate1426(.a(gate261inter10), .b(gate261inter9), .O(gate261inter11));
  nor2  gate1427(.a(gate261inter11), .b(gate261inter6), .O(gate261inter12));
  nand2 gate1428(.a(gate261inter12), .b(gate261inter1), .O(G782));
nand2 gate262( .a(G764), .b(G765), .O(G785) );

  xor2  gate1905(.a(G767), .b(G766), .O(gate263inter0));
  nand2 gate1906(.a(gate263inter0), .b(s_194), .O(gate263inter1));
  and2  gate1907(.a(G767), .b(G766), .O(gate263inter2));
  inv1  gate1908(.a(s_194), .O(gate263inter3));
  inv1  gate1909(.a(s_195), .O(gate263inter4));
  nand2 gate1910(.a(gate263inter4), .b(gate263inter3), .O(gate263inter5));
  nor2  gate1911(.a(gate263inter5), .b(gate263inter2), .O(gate263inter6));
  inv1  gate1912(.a(G766), .O(gate263inter7));
  inv1  gate1913(.a(G767), .O(gate263inter8));
  nand2 gate1914(.a(gate263inter8), .b(gate263inter7), .O(gate263inter9));
  nand2 gate1915(.a(s_195), .b(gate263inter3), .O(gate263inter10));
  nor2  gate1916(.a(gate263inter10), .b(gate263inter9), .O(gate263inter11));
  nor2  gate1917(.a(gate263inter11), .b(gate263inter6), .O(gate263inter12));
  nand2 gate1918(.a(gate263inter12), .b(gate263inter1), .O(G788));
nand2 gate264( .a(G768), .b(G769), .O(G791) );

  xor2  gate1709(.a(G770), .b(G642), .O(gate265inter0));
  nand2 gate1710(.a(gate265inter0), .b(s_166), .O(gate265inter1));
  and2  gate1711(.a(G770), .b(G642), .O(gate265inter2));
  inv1  gate1712(.a(s_166), .O(gate265inter3));
  inv1  gate1713(.a(s_167), .O(gate265inter4));
  nand2 gate1714(.a(gate265inter4), .b(gate265inter3), .O(gate265inter5));
  nor2  gate1715(.a(gate265inter5), .b(gate265inter2), .O(gate265inter6));
  inv1  gate1716(.a(G642), .O(gate265inter7));
  inv1  gate1717(.a(G770), .O(gate265inter8));
  nand2 gate1718(.a(gate265inter8), .b(gate265inter7), .O(gate265inter9));
  nand2 gate1719(.a(s_167), .b(gate265inter3), .O(gate265inter10));
  nor2  gate1720(.a(gate265inter10), .b(gate265inter9), .O(gate265inter11));
  nor2  gate1721(.a(gate265inter11), .b(gate265inter6), .O(gate265inter12));
  nand2 gate1722(.a(gate265inter12), .b(gate265inter1), .O(G794));
nand2 gate266( .a(G645), .b(G773), .O(G797) );
nand2 gate267( .a(G648), .b(G776), .O(G800) );
nand2 gate268( .a(G651), .b(G779), .O(G803) );
nand2 gate269( .a(G654), .b(G782), .O(G806) );

  xor2  gate575(.a(G785), .b(G657), .O(gate270inter0));
  nand2 gate576(.a(gate270inter0), .b(s_4), .O(gate270inter1));
  and2  gate577(.a(G785), .b(G657), .O(gate270inter2));
  inv1  gate578(.a(s_4), .O(gate270inter3));
  inv1  gate579(.a(s_5), .O(gate270inter4));
  nand2 gate580(.a(gate270inter4), .b(gate270inter3), .O(gate270inter5));
  nor2  gate581(.a(gate270inter5), .b(gate270inter2), .O(gate270inter6));
  inv1  gate582(.a(G657), .O(gate270inter7));
  inv1  gate583(.a(G785), .O(gate270inter8));
  nand2 gate584(.a(gate270inter8), .b(gate270inter7), .O(gate270inter9));
  nand2 gate585(.a(s_5), .b(gate270inter3), .O(gate270inter10));
  nor2  gate586(.a(gate270inter10), .b(gate270inter9), .O(gate270inter11));
  nor2  gate587(.a(gate270inter11), .b(gate270inter6), .O(gate270inter12));
  nand2 gate588(.a(gate270inter12), .b(gate270inter1), .O(G809));
nand2 gate271( .a(G660), .b(G788), .O(G812) );

  xor2  gate1639(.a(G791), .b(G663), .O(gate272inter0));
  nand2 gate1640(.a(gate272inter0), .b(s_156), .O(gate272inter1));
  and2  gate1641(.a(G791), .b(G663), .O(gate272inter2));
  inv1  gate1642(.a(s_156), .O(gate272inter3));
  inv1  gate1643(.a(s_157), .O(gate272inter4));
  nand2 gate1644(.a(gate272inter4), .b(gate272inter3), .O(gate272inter5));
  nor2  gate1645(.a(gate272inter5), .b(gate272inter2), .O(gate272inter6));
  inv1  gate1646(.a(G663), .O(gate272inter7));
  inv1  gate1647(.a(G791), .O(gate272inter8));
  nand2 gate1648(.a(gate272inter8), .b(gate272inter7), .O(gate272inter9));
  nand2 gate1649(.a(s_157), .b(gate272inter3), .O(gate272inter10));
  nor2  gate1650(.a(gate272inter10), .b(gate272inter9), .O(gate272inter11));
  nor2  gate1651(.a(gate272inter11), .b(gate272inter6), .O(gate272inter12));
  nand2 gate1652(.a(gate272inter12), .b(gate272inter1), .O(G815));
nand2 gate273( .a(G642), .b(G794), .O(G818) );
nand2 gate274( .a(G770), .b(G794), .O(G819) );
nand2 gate275( .a(G645), .b(G797), .O(G820) );
nand2 gate276( .a(G773), .b(G797), .O(G821) );
nand2 gate277( .a(G648), .b(G800), .O(G822) );

  xor2  gate1891(.a(G800), .b(G776), .O(gate278inter0));
  nand2 gate1892(.a(gate278inter0), .b(s_192), .O(gate278inter1));
  and2  gate1893(.a(G800), .b(G776), .O(gate278inter2));
  inv1  gate1894(.a(s_192), .O(gate278inter3));
  inv1  gate1895(.a(s_193), .O(gate278inter4));
  nand2 gate1896(.a(gate278inter4), .b(gate278inter3), .O(gate278inter5));
  nor2  gate1897(.a(gate278inter5), .b(gate278inter2), .O(gate278inter6));
  inv1  gate1898(.a(G776), .O(gate278inter7));
  inv1  gate1899(.a(G800), .O(gate278inter8));
  nand2 gate1900(.a(gate278inter8), .b(gate278inter7), .O(gate278inter9));
  nand2 gate1901(.a(s_193), .b(gate278inter3), .O(gate278inter10));
  nor2  gate1902(.a(gate278inter10), .b(gate278inter9), .O(gate278inter11));
  nor2  gate1903(.a(gate278inter11), .b(gate278inter6), .O(gate278inter12));
  nand2 gate1904(.a(gate278inter12), .b(gate278inter1), .O(G823));
nand2 gate279( .a(G651), .b(G803), .O(G824) );

  xor2  gate1751(.a(G803), .b(G779), .O(gate280inter0));
  nand2 gate1752(.a(gate280inter0), .b(s_172), .O(gate280inter1));
  and2  gate1753(.a(G803), .b(G779), .O(gate280inter2));
  inv1  gate1754(.a(s_172), .O(gate280inter3));
  inv1  gate1755(.a(s_173), .O(gate280inter4));
  nand2 gate1756(.a(gate280inter4), .b(gate280inter3), .O(gate280inter5));
  nor2  gate1757(.a(gate280inter5), .b(gate280inter2), .O(gate280inter6));
  inv1  gate1758(.a(G779), .O(gate280inter7));
  inv1  gate1759(.a(G803), .O(gate280inter8));
  nand2 gate1760(.a(gate280inter8), .b(gate280inter7), .O(gate280inter9));
  nand2 gate1761(.a(s_173), .b(gate280inter3), .O(gate280inter10));
  nor2  gate1762(.a(gate280inter10), .b(gate280inter9), .O(gate280inter11));
  nor2  gate1763(.a(gate280inter11), .b(gate280inter6), .O(gate280inter12));
  nand2 gate1764(.a(gate280inter12), .b(gate280inter1), .O(G825));
nand2 gate281( .a(G654), .b(G806), .O(G826) );
nand2 gate282( .a(G782), .b(G806), .O(G827) );
nand2 gate283( .a(G657), .b(G809), .O(G828) );
nand2 gate284( .a(G785), .b(G809), .O(G829) );
nand2 gate285( .a(G660), .b(G812), .O(G830) );
nand2 gate286( .a(G788), .b(G812), .O(G831) );
nand2 gate287( .a(G663), .b(G815), .O(G832) );
nand2 gate288( .a(G791), .b(G815), .O(G833) );
nand2 gate289( .a(G818), .b(G819), .O(G834) );

  xor2  gate2199(.a(G821), .b(G820), .O(gate290inter0));
  nand2 gate2200(.a(gate290inter0), .b(s_236), .O(gate290inter1));
  and2  gate2201(.a(G821), .b(G820), .O(gate290inter2));
  inv1  gate2202(.a(s_236), .O(gate290inter3));
  inv1  gate2203(.a(s_237), .O(gate290inter4));
  nand2 gate2204(.a(gate290inter4), .b(gate290inter3), .O(gate290inter5));
  nor2  gate2205(.a(gate290inter5), .b(gate290inter2), .O(gate290inter6));
  inv1  gate2206(.a(G820), .O(gate290inter7));
  inv1  gate2207(.a(G821), .O(gate290inter8));
  nand2 gate2208(.a(gate290inter8), .b(gate290inter7), .O(gate290inter9));
  nand2 gate2209(.a(s_237), .b(gate290inter3), .O(gate290inter10));
  nor2  gate2210(.a(gate290inter10), .b(gate290inter9), .O(gate290inter11));
  nor2  gate2211(.a(gate290inter11), .b(gate290inter6), .O(gate290inter12));
  nand2 gate2212(.a(gate290inter12), .b(gate290inter1), .O(G847));
nand2 gate291( .a(G822), .b(G823), .O(G860) );
nand2 gate292( .a(G824), .b(G825), .O(G873) );
nand2 gate293( .a(G828), .b(G829), .O(G886) );
nand2 gate294( .a(G832), .b(G833), .O(G899) );
nand2 gate295( .a(G830), .b(G831), .O(G912) );
nand2 gate296( .a(G826), .b(G827), .O(G925) );
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );
nand2 gate387( .a(G1), .b(G1036), .O(G1132) );
nand2 gate388( .a(G2), .b(G1039), .O(G1135) );
nand2 gate389( .a(G3), .b(G1042), .O(G1138) );

  xor2  gate1877(.a(G1045), .b(G4), .O(gate390inter0));
  nand2 gate1878(.a(gate390inter0), .b(s_190), .O(gate390inter1));
  and2  gate1879(.a(G1045), .b(G4), .O(gate390inter2));
  inv1  gate1880(.a(s_190), .O(gate390inter3));
  inv1  gate1881(.a(s_191), .O(gate390inter4));
  nand2 gate1882(.a(gate390inter4), .b(gate390inter3), .O(gate390inter5));
  nor2  gate1883(.a(gate390inter5), .b(gate390inter2), .O(gate390inter6));
  inv1  gate1884(.a(G4), .O(gate390inter7));
  inv1  gate1885(.a(G1045), .O(gate390inter8));
  nand2 gate1886(.a(gate390inter8), .b(gate390inter7), .O(gate390inter9));
  nand2 gate1887(.a(s_191), .b(gate390inter3), .O(gate390inter10));
  nor2  gate1888(.a(gate390inter10), .b(gate390inter9), .O(gate390inter11));
  nor2  gate1889(.a(gate390inter11), .b(gate390inter6), .O(gate390inter12));
  nand2 gate1890(.a(gate390inter12), .b(gate390inter1), .O(G1141));

  xor2  gate2129(.a(G1048), .b(G5), .O(gate391inter0));
  nand2 gate2130(.a(gate391inter0), .b(s_226), .O(gate391inter1));
  and2  gate2131(.a(G1048), .b(G5), .O(gate391inter2));
  inv1  gate2132(.a(s_226), .O(gate391inter3));
  inv1  gate2133(.a(s_227), .O(gate391inter4));
  nand2 gate2134(.a(gate391inter4), .b(gate391inter3), .O(gate391inter5));
  nor2  gate2135(.a(gate391inter5), .b(gate391inter2), .O(gate391inter6));
  inv1  gate2136(.a(G5), .O(gate391inter7));
  inv1  gate2137(.a(G1048), .O(gate391inter8));
  nand2 gate2138(.a(gate391inter8), .b(gate391inter7), .O(gate391inter9));
  nand2 gate2139(.a(s_227), .b(gate391inter3), .O(gate391inter10));
  nor2  gate2140(.a(gate391inter10), .b(gate391inter9), .O(gate391inter11));
  nor2  gate2141(.a(gate391inter11), .b(gate391inter6), .O(gate391inter12));
  nand2 gate2142(.a(gate391inter12), .b(gate391inter1), .O(G1144));

  xor2  gate1961(.a(G1051), .b(G6), .O(gate392inter0));
  nand2 gate1962(.a(gate392inter0), .b(s_202), .O(gate392inter1));
  and2  gate1963(.a(G1051), .b(G6), .O(gate392inter2));
  inv1  gate1964(.a(s_202), .O(gate392inter3));
  inv1  gate1965(.a(s_203), .O(gate392inter4));
  nand2 gate1966(.a(gate392inter4), .b(gate392inter3), .O(gate392inter5));
  nor2  gate1967(.a(gate392inter5), .b(gate392inter2), .O(gate392inter6));
  inv1  gate1968(.a(G6), .O(gate392inter7));
  inv1  gate1969(.a(G1051), .O(gate392inter8));
  nand2 gate1970(.a(gate392inter8), .b(gate392inter7), .O(gate392inter9));
  nand2 gate1971(.a(s_203), .b(gate392inter3), .O(gate392inter10));
  nor2  gate1972(.a(gate392inter10), .b(gate392inter9), .O(gate392inter11));
  nor2  gate1973(.a(gate392inter11), .b(gate392inter6), .O(gate392inter12));
  nand2 gate1974(.a(gate392inter12), .b(gate392inter1), .O(G1147));

  xor2  gate771(.a(G1054), .b(G7), .O(gate393inter0));
  nand2 gate772(.a(gate393inter0), .b(s_32), .O(gate393inter1));
  and2  gate773(.a(G1054), .b(G7), .O(gate393inter2));
  inv1  gate774(.a(s_32), .O(gate393inter3));
  inv1  gate775(.a(s_33), .O(gate393inter4));
  nand2 gate776(.a(gate393inter4), .b(gate393inter3), .O(gate393inter5));
  nor2  gate777(.a(gate393inter5), .b(gate393inter2), .O(gate393inter6));
  inv1  gate778(.a(G7), .O(gate393inter7));
  inv1  gate779(.a(G1054), .O(gate393inter8));
  nand2 gate780(.a(gate393inter8), .b(gate393inter7), .O(gate393inter9));
  nand2 gate781(.a(s_33), .b(gate393inter3), .O(gate393inter10));
  nor2  gate782(.a(gate393inter10), .b(gate393inter9), .O(gate393inter11));
  nor2  gate783(.a(gate393inter11), .b(gate393inter6), .O(gate393inter12));
  nand2 gate784(.a(gate393inter12), .b(gate393inter1), .O(G1150));
nand2 gate394( .a(G8), .b(G1057), .O(G1153) );

  xor2  gate1513(.a(G1060), .b(G9), .O(gate395inter0));
  nand2 gate1514(.a(gate395inter0), .b(s_138), .O(gate395inter1));
  and2  gate1515(.a(G1060), .b(G9), .O(gate395inter2));
  inv1  gate1516(.a(s_138), .O(gate395inter3));
  inv1  gate1517(.a(s_139), .O(gate395inter4));
  nand2 gate1518(.a(gate395inter4), .b(gate395inter3), .O(gate395inter5));
  nor2  gate1519(.a(gate395inter5), .b(gate395inter2), .O(gate395inter6));
  inv1  gate1520(.a(G9), .O(gate395inter7));
  inv1  gate1521(.a(G1060), .O(gate395inter8));
  nand2 gate1522(.a(gate395inter8), .b(gate395inter7), .O(gate395inter9));
  nand2 gate1523(.a(s_139), .b(gate395inter3), .O(gate395inter10));
  nor2  gate1524(.a(gate395inter10), .b(gate395inter9), .O(gate395inter11));
  nor2  gate1525(.a(gate395inter11), .b(gate395inter6), .O(gate395inter12));
  nand2 gate1526(.a(gate395inter12), .b(gate395inter1), .O(G1156));
nand2 gate396( .a(G10), .b(G1063), .O(G1159) );
nand2 gate397( .a(G11), .b(G1066), .O(G1162) );
nand2 gate398( .a(G12), .b(G1069), .O(G1165) );
nand2 gate399( .a(G13), .b(G1072), .O(G1168) );
nand2 gate400( .a(G14), .b(G1075), .O(G1171) );
nand2 gate401( .a(G15), .b(G1078), .O(G1174) );
nand2 gate402( .a(G16), .b(G1081), .O(G1177) );
nand2 gate403( .a(G17), .b(G1084), .O(G1180) );
nand2 gate404( .a(G18), .b(G1087), .O(G1183) );
nand2 gate405( .a(G19), .b(G1090), .O(G1186) );

  xor2  gate1135(.a(G1093), .b(G20), .O(gate406inter0));
  nand2 gate1136(.a(gate406inter0), .b(s_84), .O(gate406inter1));
  and2  gate1137(.a(G1093), .b(G20), .O(gate406inter2));
  inv1  gate1138(.a(s_84), .O(gate406inter3));
  inv1  gate1139(.a(s_85), .O(gate406inter4));
  nand2 gate1140(.a(gate406inter4), .b(gate406inter3), .O(gate406inter5));
  nor2  gate1141(.a(gate406inter5), .b(gate406inter2), .O(gate406inter6));
  inv1  gate1142(.a(G20), .O(gate406inter7));
  inv1  gate1143(.a(G1093), .O(gate406inter8));
  nand2 gate1144(.a(gate406inter8), .b(gate406inter7), .O(gate406inter9));
  nand2 gate1145(.a(s_85), .b(gate406inter3), .O(gate406inter10));
  nor2  gate1146(.a(gate406inter10), .b(gate406inter9), .O(gate406inter11));
  nor2  gate1147(.a(gate406inter11), .b(gate406inter6), .O(gate406inter12));
  nand2 gate1148(.a(gate406inter12), .b(gate406inter1), .O(G1189));

  xor2  gate2157(.a(G1096), .b(G21), .O(gate407inter0));
  nand2 gate2158(.a(gate407inter0), .b(s_230), .O(gate407inter1));
  and2  gate2159(.a(G1096), .b(G21), .O(gate407inter2));
  inv1  gate2160(.a(s_230), .O(gate407inter3));
  inv1  gate2161(.a(s_231), .O(gate407inter4));
  nand2 gate2162(.a(gate407inter4), .b(gate407inter3), .O(gate407inter5));
  nor2  gate2163(.a(gate407inter5), .b(gate407inter2), .O(gate407inter6));
  inv1  gate2164(.a(G21), .O(gate407inter7));
  inv1  gate2165(.a(G1096), .O(gate407inter8));
  nand2 gate2166(.a(gate407inter8), .b(gate407inter7), .O(gate407inter9));
  nand2 gate2167(.a(s_231), .b(gate407inter3), .O(gate407inter10));
  nor2  gate2168(.a(gate407inter10), .b(gate407inter9), .O(gate407inter11));
  nor2  gate2169(.a(gate407inter11), .b(gate407inter6), .O(gate407inter12));
  nand2 gate2170(.a(gate407inter12), .b(gate407inter1), .O(G1192));

  xor2  gate1051(.a(G1099), .b(G22), .O(gate408inter0));
  nand2 gate1052(.a(gate408inter0), .b(s_72), .O(gate408inter1));
  and2  gate1053(.a(G1099), .b(G22), .O(gate408inter2));
  inv1  gate1054(.a(s_72), .O(gate408inter3));
  inv1  gate1055(.a(s_73), .O(gate408inter4));
  nand2 gate1056(.a(gate408inter4), .b(gate408inter3), .O(gate408inter5));
  nor2  gate1057(.a(gate408inter5), .b(gate408inter2), .O(gate408inter6));
  inv1  gate1058(.a(G22), .O(gate408inter7));
  inv1  gate1059(.a(G1099), .O(gate408inter8));
  nand2 gate1060(.a(gate408inter8), .b(gate408inter7), .O(gate408inter9));
  nand2 gate1061(.a(s_73), .b(gate408inter3), .O(gate408inter10));
  nor2  gate1062(.a(gate408inter10), .b(gate408inter9), .O(gate408inter11));
  nor2  gate1063(.a(gate408inter11), .b(gate408inter6), .O(gate408inter12));
  nand2 gate1064(.a(gate408inter12), .b(gate408inter1), .O(G1195));
nand2 gate409( .a(G23), .b(G1102), .O(G1198) );
nand2 gate410( .a(G24), .b(G1105), .O(G1201) );
nand2 gate411( .a(G25), .b(G1108), .O(G1204) );
nand2 gate412( .a(G26), .b(G1111), .O(G1207) );

  xor2  gate1583(.a(G1114), .b(G27), .O(gate413inter0));
  nand2 gate1584(.a(gate413inter0), .b(s_148), .O(gate413inter1));
  and2  gate1585(.a(G1114), .b(G27), .O(gate413inter2));
  inv1  gate1586(.a(s_148), .O(gate413inter3));
  inv1  gate1587(.a(s_149), .O(gate413inter4));
  nand2 gate1588(.a(gate413inter4), .b(gate413inter3), .O(gate413inter5));
  nor2  gate1589(.a(gate413inter5), .b(gate413inter2), .O(gate413inter6));
  inv1  gate1590(.a(G27), .O(gate413inter7));
  inv1  gate1591(.a(G1114), .O(gate413inter8));
  nand2 gate1592(.a(gate413inter8), .b(gate413inter7), .O(gate413inter9));
  nand2 gate1593(.a(s_149), .b(gate413inter3), .O(gate413inter10));
  nor2  gate1594(.a(gate413inter10), .b(gate413inter9), .O(gate413inter11));
  nor2  gate1595(.a(gate413inter11), .b(gate413inter6), .O(gate413inter12));
  nand2 gate1596(.a(gate413inter12), .b(gate413inter1), .O(G1210));
nand2 gate414( .a(G28), .b(G1117), .O(G1213) );
nand2 gate415( .a(G29), .b(G1120), .O(G1216) );

  xor2  gate2143(.a(G1123), .b(G30), .O(gate416inter0));
  nand2 gate2144(.a(gate416inter0), .b(s_228), .O(gate416inter1));
  and2  gate2145(.a(G1123), .b(G30), .O(gate416inter2));
  inv1  gate2146(.a(s_228), .O(gate416inter3));
  inv1  gate2147(.a(s_229), .O(gate416inter4));
  nand2 gate2148(.a(gate416inter4), .b(gate416inter3), .O(gate416inter5));
  nor2  gate2149(.a(gate416inter5), .b(gate416inter2), .O(gate416inter6));
  inv1  gate2150(.a(G30), .O(gate416inter7));
  inv1  gate2151(.a(G1123), .O(gate416inter8));
  nand2 gate2152(.a(gate416inter8), .b(gate416inter7), .O(gate416inter9));
  nand2 gate2153(.a(s_229), .b(gate416inter3), .O(gate416inter10));
  nor2  gate2154(.a(gate416inter10), .b(gate416inter9), .O(gate416inter11));
  nor2  gate2155(.a(gate416inter11), .b(gate416inter6), .O(gate416inter12));
  nand2 gate2156(.a(gate416inter12), .b(gate416inter1), .O(G1219));

  xor2  gate785(.a(G1126), .b(G31), .O(gate417inter0));
  nand2 gate786(.a(gate417inter0), .b(s_34), .O(gate417inter1));
  and2  gate787(.a(G1126), .b(G31), .O(gate417inter2));
  inv1  gate788(.a(s_34), .O(gate417inter3));
  inv1  gate789(.a(s_35), .O(gate417inter4));
  nand2 gate790(.a(gate417inter4), .b(gate417inter3), .O(gate417inter5));
  nor2  gate791(.a(gate417inter5), .b(gate417inter2), .O(gate417inter6));
  inv1  gate792(.a(G31), .O(gate417inter7));
  inv1  gate793(.a(G1126), .O(gate417inter8));
  nand2 gate794(.a(gate417inter8), .b(gate417inter7), .O(gate417inter9));
  nand2 gate795(.a(s_35), .b(gate417inter3), .O(gate417inter10));
  nor2  gate796(.a(gate417inter10), .b(gate417inter9), .O(gate417inter11));
  nor2  gate797(.a(gate417inter11), .b(gate417inter6), .O(gate417inter12));
  nand2 gate798(.a(gate417inter12), .b(gate417inter1), .O(G1222));

  xor2  gate687(.a(G1129), .b(G32), .O(gate418inter0));
  nand2 gate688(.a(gate418inter0), .b(s_20), .O(gate418inter1));
  and2  gate689(.a(G1129), .b(G32), .O(gate418inter2));
  inv1  gate690(.a(s_20), .O(gate418inter3));
  inv1  gate691(.a(s_21), .O(gate418inter4));
  nand2 gate692(.a(gate418inter4), .b(gate418inter3), .O(gate418inter5));
  nor2  gate693(.a(gate418inter5), .b(gate418inter2), .O(gate418inter6));
  inv1  gate694(.a(G32), .O(gate418inter7));
  inv1  gate695(.a(G1129), .O(gate418inter8));
  nand2 gate696(.a(gate418inter8), .b(gate418inter7), .O(gate418inter9));
  nand2 gate697(.a(s_21), .b(gate418inter3), .O(gate418inter10));
  nor2  gate698(.a(gate418inter10), .b(gate418inter9), .O(gate418inter11));
  nor2  gate699(.a(gate418inter11), .b(gate418inter6), .O(gate418inter12));
  nand2 gate700(.a(gate418inter12), .b(gate418inter1), .O(G1225));

  xor2  gate1611(.a(G1132), .b(G1), .O(gate419inter0));
  nand2 gate1612(.a(gate419inter0), .b(s_152), .O(gate419inter1));
  and2  gate1613(.a(G1132), .b(G1), .O(gate419inter2));
  inv1  gate1614(.a(s_152), .O(gate419inter3));
  inv1  gate1615(.a(s_153), .O(gate419inter4));
  nand2 gate1616(.a(gate419inter4), .b(gate419inter3), .O(gate419inter5));
  nor2  gate1617(.a(gate419inter5), .b(gate419inter2), .O(gate419inter6));
  inv1  gate1618(.a(G1), .O(gate419inter7));
  inv1  gate1619(.a(G1132), .O(gate419inter8));
  nand2 gate1620(.a(gate419inter8), .b(gate419inter7), .O(gate419inter9));
  nand2 gate1621(.a(s_153), .b(gate419inter3), .O(gate419inter10));
  nor2  gate1622(.a(gate419inter10), .b(gate419inter9), .O(gate419inter11));
  nor2  gate1623(.a(gate419inter11), .b(gate419inter6), .O(gate419inter12));
  nand2 gate1624(.a(gate419inter12), .b(gate419inter1), .O(G1228));
nand2 gate420( .a(G1036), .b(G1132), .O(G1229) );
nand2 gate421( .a(G2), .b(G1135), .O(G1230) );
nand2 gate422( .a(G1039), .b(G1135), .O(G1231) );
nand2 gate423( .a(G3), .b(G1138), .O(G1232) );
nand2 gate424( .a(G1042), .b(G1138), .O(G1233) );

  xor2  gate1919(.a(G1141), .b(G4), .O(gate425inter0));
  nand2 gate1920(.a(gate425inter0), .b(s_196), .O(gate425inter1));
  and2  gate1921(.a(G1141), .b(G4), .O(gate425inter2));
  inv1  gate1922(.a(s_196), .O(gate425inter3));
  inv1  gate1923(.a(s_197), .O(gate425inter4));
  nand2 gate1924(.a(gate425inter4), .b(gate425inter3), .O(gate425inter5));
  nor2  gate1925(.a(gate425inter5), .b(gate425inter2), .O(gate425inter6));
  inv1  gate1926(.a(G4), .O(gate425inter7));
  inv1  gate1927(.a(G1141), .O(gate425inter8));
  nand2 gate1928(.a(gate425inter8), .b(gate425inter7), .O(gate425inter9));
  nand2 gate1929(.a(s_197), .b(gate425inter3), .O(gate425inter10));
  nor2  gate1930(.a(gate425inter10), .b(gate425inter9), .O(gate425inter11));
  nor2  gate1931(.a(gate425inter11), .b(gate425inter6), .O(gate425inter12));
  nand2 gate1932(.a(gate425inter12), .b(gate425inter1), .O(G1234));

  xor2  gate1303(.a(G1141), .b(G1045), .O(gate426inter0));
  nand2 gate1304(.a(gate426inter0), .b(s_108), .O(gate426inter1));
  and2  gate1305(.a(G1141), .b(G1045), .O(gate426inter2));
  inv1  gate1306(.a(s_108), .O(gate426inter3));
  inv1  gate1307(.a(s_109), .O(gate426inter4));
  nand2 gate1308(.a(gate426inter4), .b(gate426inter3), .O(gate426inter5));
  nor2  gate1309(.a(gate426inter5), .b(gate426inter2), .O(gate426inter6));
  inv1  gate1310(.a(G1045), .O(gate426inter7));
  inv1  gate1311(.a(G1141), .O(gate426inter8));
  nand2 gate1312(.a(gate426inter8), .b(gate426inter7), .O(gate426inter9));
  nand2 gate1313(.a(s_109), .b(gate426inter3), .O(gate426inter10));
  nor2  gate1314(.a(gate426inter10), .b(gate426inter9), .O(gate426inter11));
  nor2  gate1315(.a(gate426inter11), .b(gate426inter6), .O(gate426inter12));
  nand2 gate1316(.a(gate426inter12), .b(gate426inter1), .O(G1235));
nand2 gate427( .a(G5), .b(G1144), .O(G1236) );
nand2 gate428( .a(G1048), .b(G1144), .O(G1237) );

  xor2  gate1023(.a(G1147), .b(G6), .O(gate429inter0));
  nand2 gate1024(.a(gate429inter0), .b(s_68), .O(gate429inter1));
  and2  gate1025(.a(G1147), .b(G6), .O(gate429inter2));
  inv1  gate1026(.a(s_68), .O(gate429inter3));
  inv1  gate1027(.a(s_69), .O(gate429inter4));
  nand2 gate1028(.a(gate429inter4), .b(gate429inter3), .O(gate429inter5));
  nor2  gate1029(.a(gate429inter5), .b(gate429inter2), .O(gate429inter6));
  inv1  gate1030(.a(G6), .O(gate429inter7));
  inv1  gate1031(.a(G1147), .O(gate429inter8));
  nand2 gate1032(.a(gate429inter8), .b(gate429inter7), .O(gate429inter9));
  nand2 gate1033(.a(s_69), .b(gate429inter3), .O(gate429inter10));
  nor2  gate1034(.a(gate429inter10), .b(gate429inter9), .O(gate429inter11));
  nor2  gate1035(.a(gate429inter11), .b(gate429inter6), .O(gate429inter12));
  nand2 gate1036(.a(gate429inter12), .b(gate429inter1), .O(G1238));
nand2 gate430( .a(G1051), .b(G1147), .O(G1239) );
nand2 gate431( .a(G7), .b(G1150), .O(G1240) );

  xor2  gate1807(.a(G1150), .b(G1054), .O(gate432inter0));
  nand2 gate1808(.a(gate432inter0), .b(s_180), .O(gate432inter1));
  and2  gate1809(.a(G1150), .b(G1054), .O(gate432inter2));
  inv1  gate1810(.a(s_180), .O(gate432inter3));
  inv1  gate1811(.a(s_181), .O(gate432inter4));
  nand2 gate1812(.a(gate432inter4), .b(gate432inter3), .O(gate432inter5));
  nor2  gate1813(.a(gate432inter5), .b(gate432inter2), .O(gate432inter6));
  inv1  gate1814(.a(G1054), .O(gate432inter7));
  inv1  gate1815(.a(G1150), .O(gate432inter8));
  nand2 gate1816(.a(gate432inter8), .b(gate432inter7), .O(gate432inter9));
  nand2 gate1817(.a(s_181), .b(gate432inter3), .O(gate432inter10));
  nor2  gate1818(.a(gate432inter10), .b(gate432inter9), .O(gate432inter11));
  nor2  gate1819(.a(gate432inter11), .b(gate432inter6), .O(gate432inter12));
  nand2 gate1820(.a(gate432inter12), .b(gate432inter1), .O(G1241));
nand2 gate433( .a(G8), .b(G1153), .O(G1242) );

  xor2  gate1541(.a(G1153), .b(G1057), .O(gate434inter0));
  nand2 gate1542(.a(gate434inter0), .b(s_142), .O(gate434inter1));
  and2  gate1543(.a(G1153), .b(G1057), .O(gate434inter2));
  inv1  gate1544(.a(s_142), .O(gate434inter3));
  inv1  gate1545(.a(s_143), .O(gate434inter4));
  nand2 gate1546(.a(gate434inter4), .b(gate434inter3), .O(gate434inter5));
  nor2  gate1547(.a(gate434inter5), .b(gate434inter2), .O(gate434inter6));
  inv1  gate1548(.a(G1057), .O(gate434inter7));
  inv1  gate1549(.a(G1153), .O(gate434inter8));
  nand2 gate1550(.a(gate434inter8), .b(gate434inter7), .O(gate434inter9));
  nand2 gate1551(.a(s_143), .b(gate434inter3), .O(gate434inter10));
  nor2  gate1552(.a(gate434inter10), .b(gate434inter9), .O(gate434inter11));
  nor2  gate1553(.a(gate434inter11), .b(gate434inter6), .O(gate434inter12));
  nand2 gate1554(.a(gate434inter12), .b(gate434inter1), .O(G1243));
nand2 gate435( .a(G9), .b(G1156), .O(G1244) );
nand2 gate436( .a(G1060), .b(G1156), .O(G1245) );

  xor2  gate1975(.a(G1159), .b(G10), .O(gate437inter0));
  nand2 gate1976(.a(gate437inter0), .b(s_204), .O(gate437inter1));
  and2  gate1977(.a(G1159), .b(G10), .O(gate437inter2));
  inv1  gate1978(.a(s_204), .O(gate437inter3));
  inv1  gate1979(.a(s_205), .O(gate437inter4));
  nand2 gate1980(.a(gate437inter4), .b(gate437inter3), .O(gate437inter5));
  nor2  gate1981(.a(gate437inter5), .b(gate437inter2), .O(gate437inter6));
  inv1  gate1982(.a(G10), .O(gate437inter7));
  inv1  gate1983(.a(G1159), .O(gate437inter8));
  nand2 gate1984(.a(gate437inter8), .b(gate437inter7), .O(gate437inter9));
  nand2 gate1985(.a(s_205), .b(gate437inter3), .O(gate437inter10));
  nor2  gate1986(.a(gate437inter10), .b(gate437inter9), .O(gate437inter11));
  nor2  gate1987(.a(gate437inter11), .b(gate437inter6), .O(gate437inter12));
  nand2 gate1988(.a(gate437inter12), .b(gate437inter1), .O(G1246));
nand2 gate438( .a(G1063), .b(G1159), .O(G1247) );

  xor2  gate1443(.a(G1162), .b(G11), .O(gate439inter0));
  nand2 gate1444(.a(gate439inter0), .b(s_128), .O(gate439inter1));
  and2  gate1445(.a(G1162), .b(G11), .O(gate439inter2));
  inv1  gate1446(.a(s_128), .O(gate439inter3));
  inv1  gate1447(.a(s_129), .O(gate439inter4));
  nand2 gate1448(.a(gate439inter4), .b(gate439inter3), .O(gate439inter5));
  nor2  gate1449(.a(gate439inter5), .b(gate439inter2), .O(gate439inter6));
  inv1  gate1450(.a(G11), .O(gate439inter7));
  inv1  gate1451(.a(G1162), .O(gate439inter8));
  nand2 gate1452(.a(gate439inter8), .b(gate439inter7), .O(gate439inter9));
  nand2 gate1453(.a(s_129), .b(gate439inter3), .O(gate439inter10));
  nor2  gate1454(.a(gate439inter10), .b(gate439inter9), .O(gate439inter11));
  nor2  gate1455(.a(gate439inter11), .b(gate439inter6), .O(gate439inter12));
  nand2 gate1456(.a(gate439inter12), .b(gate439inter1), .O(G1248));

  xor2  gate1653(.a(G1162), .b(G1066), .O(gate440inter0));
  nand2 gate1654(.a(gate440inter0), .b(s_158), .O(gate440inter1));
  and2  gate1655(.a(G1162), .b(G1066), .O(gate440inter2));
  inv1  gate1656(.a(s_158), .O(gate440inter3));
  inv1  gate1657(.a(s_159), .O(gate440inter4));
  nand2 gate1658(.a(gate440inter4), .b(gate440inter3), .O(gate440inter5));
  nor2  gate1659(.a(gate440inter5), .b(gate440inter2), .O(gate440inter6));
  inv1  gate1660(.a(G1066), .O(gate440inter7));
  inv1  gate1661(.a(G1162), .O(gate440inter8));
  nand2 gate1662(.a(gate440inter8), .b(gate440inter7), .O(gate440inter9));
  nand2 gate1663(.a(s_159), .b(gate440inter3), .O(gate440inter10));
  nor2  gate1664(.a(gate440inter10), .b(gate440inter9), .O(gate440inter11));
  nor2  gate1665(.a(gate440inter11), .b(gate440inter6), .O(gate440inter12));
  nand2 gate1666(.a(gate440inter12), .b(gate440inter1), .O(G1249));
nand2 gate441( .a(G12), .b(G1165), .O(G1250) );
nand2 gate442( .a(G1069), .b(G1165), .O(G1251) );
nand2 gate443( .a(G13), .b(G1168), .O(G1252) );
nand2 gate444( .a(G1072), .b(G1168), .O(G1253) );
nand2 gate445( .a(G14), .b(G1171), .O(G1254) );
nand2 gate446( .a(G1075), .b(G1171), .O(G1255) );
nand2 gate447( .a(G15), .b(G1174), .O(G1256) );
nand2 gate448( .a(G1078), .b(G1174), .O(G1257) );

  xor2  gate715(.a(G1177), .b(G16), .O(gate449inter0));
  nand2 gate716(.a(gate449inter0), .b(s_24), .O(gate449inter1));
  and2  gate717(.a(G1177), .b(G16), .O(gate449inter2));
  inv1  gate718(.a(s_24), .O(gate449inter3));
  inv1  gate719(.a(s_25), .O(gate449inter4));
  nand2 gate720(.a(gate449inter4), .b(gate449inter3), .O(gate449inter5));
  nor2  gate721(.a(gate449inter5), .b(gate449inter2), .O(gate449inter6));
  inv1  gate722(.a(G16), .O(gate449inter7));
  inv1  gate723(.a(G1177), .O(gate449inter8));
  nand2 gate724(.a(gate449inter8), .b(gate449inter7), .O(gate449inter9));
  nand2 gate725(.a(s_25), .b(gate449inter3), .O(gate449inter10));
  nor2  gate726(.a(gate449inter10), .b(gate449inter9), .O(gate449inter11));
  nor2  gate727(.a(gate449inter11), .b(gate449inter6), .O(gate449inter12));
  nand2 gate728(.a(gate449inter12), .b(gate449inter1), .O(G1258));
nand2 gate450( .a(G1081), .b(G1177), .O(G1259) );
nand2 gate451( .a(G17), .b(G1180), .O(G1260) );
nand2 gate452( .a(G1084), .b(G1180), .O(G1261) );
nand2 gate453( .a(G18), .b(G1183), .O(G1262) );
nand2 gate454( .a(G1087), .b(G1183), .O(G1263) );
nand2 gate455( .a(G19), .b(G1186), .O(G1264) );
nand2 gate456( .a(G1090), .b(G1186), .O(G1265) );
nand2 gate457( .a(G20), .b(G1189), .O(G1266) );
nand2 gate458( .a(G1093), .b(G1189), .O(G1267) );
nand2 gate459( .a(G21), .b(G1192), .O(G1268) );
nand2 gate460( .a(G1096), .b(G1192), .O(G1269) );
nand2 gate461( .a(G22), .b(G1195), .O(G1270) );
nand2 gate462( .a(G1099), .b(G1195), .O(G1271) );
nand2 gate463( .a(G23), .b(G1198), .O(G1272) );
nand2 gate464( .a(G1102), .b(G1198), .O(G1273) );
nand2 gate465( .a(G24), .b(G1201), .O(G1274) );

  xor2  gate2185(.a(G1201), .b(G1105), .O(gate466inter0));
  nand2 gate2186(.a(gate466inter0), .b(s_234), .O(gate466inter1));
  and2  gate2187(.a(G1201), .b(G1105), .O(gate466inter2));
  inv1  gate2188(.a(s_234), .O(gate466inter3));
  inv1  gate2189(.a(s_235), .O(gate466inter4));
  nand2 gate2190(.a(gate466inter4), .b(gate466inter3), .O(gate466inter5));
  nor2  gate2191(.a(gate466inter5), .b(gate466inter2), .O(gate466inter6));
  inv1  gate2192(.a(G1105), .O(gate466inter7));
  inv1  gate2193(.a(G1201), .O(gate466inter8));
  nand2 gate2194(.a(gate466inter8), .b(gate466inter7), .O(gate466inter9));
  nand2 gate2195(.a(s_235), .b(gate466inter3), .O(gate466inter10));
  nor2  gate2196(.a(gate466inter10), .b(gate466inter9), .O(gate466inter11));
  nor2  gate2197(.a(gate466inter11), .b(gate466inter6), .O(gate466inter12));
  nand2 gate2198(.a(gate466inter12), .b(gate466inter1), .O(G1275));
nand2 gate467( .a(G25), .b(G1204), .O(G1276) );

  xor2  gate1835(.a(G1204), .b(G1108), .O(gate468inter0));
  nand2 gate1836(.a(gate468inter0), .b(s_184), .O(gate468inter1));
  and2  gate1837(.a(G1204), .b(G1108), .O(gate468inter2));
  inv1  gate1838(.a(s_184), .O(gate468inter3));
  inv1  gate1839(.a(s_185), .O(gate468inter4));
  nand2 gate1840(.a(gate468inter4), .b(gate468inter3), .O(gate468inter5));
  nor2  gate1841(.a(gate468inter5), .b(gate468inter2), .O(gate468inter6));
  inv1  gate1842(.a(G1108), .O(gate468inter7));
  inv1  gate1843(.a(G1204), .O(gate468inter8));
  nand2 gate1844(.a(gate468inter8), .b(gate468inter7), .O(gate468inter9));
  nand2 gate1845(.a(s_185), .b(gate468inter3), .O(gate468inter10));
  nor2  gate1846(.a(gate468inter10), .b(gate468inter9), .O(gate468inter11));
  nor2  gate1847(.a(gate468inter11), .b(gate468inter6), .O(gate468inter12));
  nand2 gate1848(.a(gate468inter12), .b(gate468inter1), .O(G1277));
nand2 gate469( .a(G26), .b(G1207), .O(G1278) );
nand2 gate470( .a(G1111), .b(G1207), .O(G1279) );

  xor2  gate547(.a(G1210), .b(G27), .O(gate471inter0));
  nand2 gate548(.a(gate471inter0), .b(s_0), .O(gate471inter1));
  and2  gate549(.a(G1210), .b(G27), .O(gate471inter2));
  inv1  gate550(.a(s_0), .O(gate471inter3));
  inv1  gate551(.a(s_1), .O(gate471inter4));
  nand2 gate552(.a(gate471inter4), .b(gate471inter3), .O(gate471inter5));
  nor2  gate553(.a(gate471inter5), .b(gate471inter2), .O(gate471inter6));
  inv1  gate554(.a(G27), .O(gate471inter7));
  inv1  gate555(.a(G1210), .O(gate471inter8));
  nand2 gate556(.a(gate471inter8), .b(gate471inter7), .O(gate471inter9));
  nand2 gate557(.a(s_1), .b(gate471inter3), .O(gate471inter10));
  nor2  gate558(.a(gate471inter10), .b(gate471inter9), .O(gate471inter11));
  nor2  gate559(.a(gate471inter11), .b(gate471inter6), .O(gate471inter12));
  nand2 gate560(.a(gate471inter12), .b(gate471inter1), .O(G1280));
nand2 gate472( .a(G1114), .b(G1210), .O(G1281) );
nand2 gate473( .a(G28), .b(G1213), .O(G1282) );

  xor2  gate701(.a(G1213), .b(G1117), .O(gate474inter0));
  nand2 gate702(.a(gate474inter0), .b(s_22), .O(gate474inter1));
  and2  gate703(.a(G1213), .b(G1117), .O(gate474inter2));
  inv1  gate704(.a(s_22), .O(gate474inter3));
  inv1  gate705(.a(s_23), .O(gate474inter4));
  nand2 gate706(.a(gate474inter4), .b(gate474inter3), .O(gate474inter5));
  nor2  gate707(.a(gate474inter5), .b(gate474inter2), .O(gate474inter6));
  inv1  gate708(.a(G1117), .O(gate474inter7));
  inv1  gate709(.a(G1213), .O(gate474inter8));
  nand2 gate710(.a(gate474inter8), .b(gate474inter7), .O(gate474inter9));
  nand2 gate711(.a(s_23), .b(gate474inter3), .O(gate474inter10));
  nor2  gate712(.a(gate474inter10), .b(gate474inter9), .O(gate474inter11));
  nor2  gate713(.a(gate474inter11), .b(gate474inter6), .O(gate474inter12));
  nand2 gate714(.a(gate474inter12), .b(gate474inter1), .O(G1283));
nand2 gate475( .a(G29), .b(G1216), .O(G1284) );
nand2 gate476( .a(G1120), .b(G1216), .O(G1285) );

  xor2  gate1107(.a(G1219), .b(G30), .O(gate477inter0));
  nand2 gate1108(.a(gate477inter0), .b(s_80), .O(gate477inter1));
  and2  gate1109(.a(G1219), .b(G30), .O(gate477inter2));
  inv1  gate1110(.a(s_80), .O(gate477inter3));
  inv1  gate1111(.a(s_81), .O(gate477inter4));
  nand2 gate1112(.a(gate477inter4), .b(gate477inter3), .O(gate477inter5));
  nor2  gate1113(.a(gate477inter5), .b(gate477inter2), .O(gate477inter6));
  inv1  gate1114(.a(G30), .O(gate477inter7));
  inv1  gate1115(.a(G1219), .O(gate477inter8));
  nand2 gate1116(.a(gate477inter8), .b(gate477inter7), .O(gate477inter9));
  nand2 gate1117(.a(s_81), .b(gate477inter3), .O(gate477inter10));
  nor2  gate1118(.a(gate477inter10), .b(gate477inter9), .O(gate477inter11));
  nor2  gate1119(.a(gate477inter11), .b(gate477inter6), .O(gate477inter12));
  nand2 gate1120(.a(gate477inter12), .b(gate477inter1), .O(G1286));
nand2 gate478( .a(G1123), .b(G1219), .O(G1287) );
nand2 gate479( .a(G31), .b(G1222), .O(G1288) );

  xor2  gate1569(.a(G1222), .b(G1126), .O(gate480inter0));
  nand2 gate1570(.a(gate480inter0), .b(s_146), .O(gate480inter1));
  and2  gate1571(.a(G1222), .b(G1126), .O(gate480inter2));
  inv1  gate1572(.a(s_146), .O(gate480inter3));
  inv1  gate1573(.a(s_147), .O(gate480inter4));
  nand2 gate1574(.a(gate480inter4), .b(gate480inter3), .O(gate480inter5));
  nor2  gate1575(.a(gate480inter5), .b(gate480inter2), .O(gate480inter6));
  inv1  gate1576(.a(G1126), .O(gate480inter7));
  inv1  gate1577(.a(G1222), .O(gate480inter8));
  nand2 gate1578(.a(gate480inter8), .b(gate480inter7), .O(gate480inter9));
  nand2 gate1579(.a(s_147), .b(gate480inter3), .O(gate480inter10));
  nor2  gate1580(.a(gate480inter10), .b(gate480inter9), .O(gate480inter11));
  nor2  gate1581(.a(gate480inter11), .b(gate480inter6), .O(gate480inter12));
  nand2 gate1582(.a(gate480inter12), .b(gate480inter1), .O(G1289));
nand2 gate481( .a(G32), .b(G1225), .O(G1290) );
nand2 gate482( .a(G1129), .b(G1225), .O(G1291) );

  xor2  gate2017(.a(G1229), .b(G1228), .O(gate483inter0));
  nand2 gate2018(.a(gate483inter0), .b(s_210), .O(gate483inter1));
  and2  gate2019(.a(G1229), .b(G1228), .O(gate483inter2));
  inv1  gate2020(.a(s_210), .O(gate483inter3));
  inv1  gate2021(.a(s_211), .O(gate483inter4));
  nand2 gate2022(.a(gate483inter4), .b(gate483inter3), .O(gate483inter5));
  nor2  gate2023(.a(gate483inter5), .b(gate483inter2), .O(gate483inter6));
  inv1  gate2024(.a(G1228), .O(gate483inter7));
  inv1  gate2025(.a(G1229), .O(gate483inter8));
  nand2 gate2026(.a(gate483inter8), .b(gate483inter7), .O(gate483inter9));
  nand2 gate2027(.a(s_211), .b(gate483inter3), .O(gate483inter10));
  nor2  gate2028(.a(gate483inter10), .b(gate483inter9), .O(gate483inter11));
  nor2  gate2029(.a(gate483inter11), .b(gate483inter6), .O(gate483inter12));
  nand2 gate2030(.a(gate483inter12), .b(gate483inter1), .O(G1292));
nand2 gate484( .a(G1230), .b(G1231), .O(G1293) );
nand2 gate485( .a(G1232), .b(G1233), .O(G1294) );
nand2 gate486( .a(G1234), .b(G1235), .O(G1295) );
nand2 gate487( .a(G1236), .b(G1237), .O(G1296) );
nand2 gate488( .a(G1238), .b(G1239), .O(G1297) );
nand2 gate489( .a(G1240), .b(G1241), .O(G1298) );
nand2 gate490( .a(G1242), .b(G1243), .O(G1299) );
nand2 gate491( .a(G1244), .b(G1245), .O(G1300) );
nand2 gate492( .a(G1246), .b(G1247), .O(G1301) );
nand2 gate493( .a(G1248), .b(G1249), .O(G1302) );

  xor2  gate1065(.a(G1251), .b(G1250), .O(gate494inter0));
  nand2 gate1066(.a(gate494inter0), .b(s_74), .O(gate494inter1));
  and2  gate1067(.a(G1251), .b(G1250), .O(gate494inter2));
  inv1  gate1068(.a(s_74), .O(gate494inter3));
  inv1  gate1069(.a(s_75), .O(gate494inter4));
  nand2 gate1070(.a(gate494inter4), .b(gate494inter3), .O(gate494inter5));
  nor2  gate1071(.a(gate494inter5), .b(gate494inter2), .O(gate494inter6));
  inv1  gate1072(.a(G1250), .O(gate494inter7));
  inv1  gate1073(.a(G1251), .O(gate494inter8));
  nand2 gate1074(.a(gate494inter8), .b(gate494inter7), .O(gate494inter9));
  nand2 gate1075(.a(s_75), .b(gate494inter3), .O(gate494inter10));
  nor2  gate1076(.a(gate494inter10), .b(gate494inter9), .O(gate494inter11));
  nor2  gate1077(.a(gate494inter11), .b(gate494inter6), .O(gate494inter12));
  nand2 gate1078(.a(gate494inter12), .b(gate494inter1), .O(G1303));
nand2 gate495( .a(G1252), .b(G1253), .O(G1304) );

  xor2  gate1275(.a(G1255), .b(G1254), .O(gate496inter0));
  nand2 gate1276(.a(gate496inter0), .b(s_104), .O(gate496inter1));
  and2  gate1277(.a(G1255), .b(G1254), .O(gate496inter2));
  inv1  gate1278(.a(s_104), .O(gate496inter3));
  inv1  gate1279(.a(s_105), .O(gate496inter4));
  nand2 gate1280(.a(gate496inter4), .b(gate496inter3), .O(gate496inter5));
  nor2  gate1281(.a(gate496inter5), .b(gate496inter2), .O(gate496inter6));
  inv1  gate1282(.a(G1254), .O(gate496inter7));
  inv1  gate1283(.a(G1255), .O(gate496inter8));
  nand2 gate1284(.a(gate496inter8), .b(gate496inter7), .O(gate496inter9));
  nand2 gate1285(.a(s_105), .b(gate496inter3), .O(gate496inter10));
  nor2  gate1286(.a(gate496inter10), .b(gate496inter9), .O(gate496inter11));
  nor2  gate1287(.a(gate496inter11), .b(gate496inter6), .O(gate496inter12));
  nand2 gate1288(.a(gate496inter12), .b(gate496inter1), .O(G1305));

  xor2  gate869(.a(G1257), .b(G1256), .O(gate497inter0));
  nand2 gate870(.a(gate497inter0), .b(s_46), .O(gate497inter1));
  and2  gate871(.a(G1257), .b(G1256), .O(gate497inter2));
  inv1  gate872(.a(s_46), .O(gate497inter3));
  inv1  gate873(.a(s_47), .O(gate497inter4));
  nand2 gate874(.a(gate497inter4), .b(gate497inter3), .O(gate497inter5));
  nor2  gate875(.a(gate497inter5), .b(gate497inter2), .O(gate497inter6));
  inv1  gate876(.a(G1256), .O(gate497inter7));
  inv1  gate877(.a(G1257), .O(gate497inter8));
  nand2 gate878(.a(gate497inter8), .b(gate497inter7), .O(gate497inter9));
  nand2 gate879(.a(s_47), .b(gate497inter3), .O(gate497inter10));
  nor2  gate880(.a(gate497inter10), .b(gate497inter9), .O(gate497inter11));
  nor2  gate881(.a(gate497inter11), .b(gate497inter6), .O(gate497inter12));
  nand2 gate882(.a(gate497inter12), .b(gate497inter1), .O(G1306));
nand2 gate498( .a(G1258), .b(G1259), .O(G1307) );
nand2 gate499( .a(G1260), .b(G1261), .O(G1308) );
nand2 gate500( .a(G1262), .b(G1263), .O(G1309) );

  xor2  gate1317(.a(G1265), .b(G1264), .O(gate501inter0));
  nand2 gate1318(.a(gate501inter0), .b(s_110), .O(gate501inter1));
  and2  gate1319(.a(G1265), .b(G1264), .O(gate501inter2));
  inv1  gate1320(.a(s_110), .O(gate501inter3));
  inv1  gate1321(.a(s_111), .O(gate501inter4));
  nand2 gate1322(.a(gate501inter4), .b(gate501inter3), .O(gate501inter5));
  nor2  gate1323(.a(gate501inter5), .b(gate501inter2), .O(gate501inter6));
  inv1  gate1324(.a(G1264), .O(gate501inter7));
  inv1  gate1325(.a(G1265), .O(gate501inter8));
  nand2 gate1326(.a(gate501inter8), .b(gate501inter7), .O(gate501inter9));
  nand2 gate1327(.a(s_111), .b(gate501inter3), .O(gate501inter10));
  nor2  gate1328(.a(gate501inter10), .b(gate501inter9), .O(gate501inter11));
  nor2  gate1329(.a(gate501inter11), .b(gate501inter6), .O(gate501inter12));
  nand2 gate1330(.a(gate501inter12), .b(gate501inter1), .O(G1310));
nand2 gate502( .a(G1266), .b(G1267), .O(G1311) );
nand2 gate503( .a(G1268), .b(G1269), .O(G1312) );
nand2 gate504( .a(G1270), .b(G1271), .O(G1313) );
nand2 gate505( .a(G1272), .b(G1273), .O(G1314) );

  xor2  gate2045(.a(G1275), .b(G1274), .O(gate506inter0));
  nand2 gate2046(.a(gate506inter0), .b(s_214), .O(gate506inter1));
  and2  gate2047(.a(G1275), .b(G1274), .O(gate506inter2));
  inv1  gate2048(.a(s_214), .O(gate506inter3));
  inv1  gate2049(.a(s_215), .O(gate506inter4));
  nand2 gate2050(.a(gate506inter4), .b(gate506inter3), .O(gate506inter5));
  nor2  gate2051(.a(gate506inter5), .b(gate506inter2), .O(gate506inter6));
  inv1  gate2052(.a(G1274), .O(gate506inter7));
  inv1  gate2053(.a(G1275), .O(gate506inter8));
  nand2 gate2054(.a(gate506inter8), .b(gate506inter7), .O(gate506inter9));
  nand2 gate2055(.a(s_215), .b(gate506inter3), .O(gate506inter10));
  nor2  gate2056(.a(gate506inter10), .b(gate506inter9), .O(gate506inter11));
  nor2  gate2057(.a(gate506inter11), .b(gate506inter6), .O(gate506inter12));
  nand2 gate2058(.a(gate506inter12), .b(gate506inter1), .O(G1315));
nand2 gate507( .a(G1276), .b(G1277), .O(G1316) );

  xor2  gate2213(.a(G1279), .b(G1278), .O(gate508inter0));
  nand2 gate2214(.a(gate508inter0), .b(s_238), .O(gate508inter1));
  and2  gate2215(.a(G1279), .b(G1278), .O(gate508inter2));
  inv1  gate2216(.a(s_238), .O(gate508inter3));
  inv1  gate2217(.a(s_239), .O(gate508inter4));
  nand2 gate2218(.a(gate508inter4), .b(gate508inter3), .O(gate508inter5));
  nor2  gate2219(.a(gate508inter5), .b(gate508inter2), .O(gate508inter6));
  inv1  gate2220(.a(G1278), .O(gate508inter7));
  inv1  gate2221(.a(G1279), .O(gate508inter8));
  nand2 gate2222(.a(gate508inter8), .b(gate508inter7), .O(gate508inter9));
  nand2 gate2223(.a(s_239), .b(gate508inter3), .O(gate508inter10));
  nor2  gate2224(.a(gate508inter10), .b(gate508inter9), .O(gate508inter11));
  nor2  gate2225(.a(gate508inter11), .b(gate508inter6), .O(gate508inter12));
  nand2 gate2226(.a(gate508inter12), .b(gate508inter1), .O(G1317));
nand2 gate509( .a(G1280), .b(G1281), .O(G1318) );

  xor2  gate2115(.a(G1283), .b(G1282), .O(gate510inter0));
  nand2 gate2116(.a(gate510inter0), .b(s_224), .O(gate510inter1));
  and2  gate2117(.a(G1283), .b(G1282), .O(gate510inter2));
  inv1  gate2118(.a(s_224), .O(gate510inter3));
  inv1  gate2119(.a(s_225), .O(gate510inter4));
  nand2 gate2120(.a(gate510inter4), .b(gate510inter3), .O(gate510inter5));
  nor2  gate2121(.a(gate510inter5), .b(gate510inter2), .O(gate510inter6));
  inv1  gate2122(.a(G1282), .O(gate510inter7));
  inv1  gate2123(.a(G1283), .O(gate510inter8));
  nand2 gate2124(.a(gate510inter8), .b(gate510inter7), .O(gate510inter9));
  nand2 gate2125(.a(s_225), .b(gate510inter3), .O(gate510inter10));
  nor2  gate2126(.a(gate510inter10), .b(gate510inter9), .O(gate510inter11));
  nor2  gate2127(.a(gate510inter11), .b(gate510inter6), .O(gate510inter12));
  nand2 gate2128(.a(gate510inter12), .b(gate510inter1), .O(G1319));

  xor2  gate827(.a(G1285), .b(G1284), .O(gate511inter0));
  nand2 gate828(.a(gate511inter0), .b(s_40), .O(gate511inter1));
  and2  gate829(.a(G1285), .b(G1284), .O(gate511inter2));
  inv1  gate830(.a(s_40), .O(gate511inter3));
  inv1  gate831(.a(s_41), .O(gate511inter4));
  nand2 gate832(.a(gate511inter4), .b(gate511inter3), .O(gate511inter5));
  nor2  gate833(.a(gate511inter5), .b(gate511inter2), .O(gate511inter6));
  inv1  gate834(.a(G1284), .O(gate511inter7));
  inv1  gate835(.a(G1285), .O(gate511inter8));
  nand2 gate836(.a(gate511inter8), .b(gate511inter7), .O(gate511inter9));
  nand2 gate837(.a(s_41), .b(gate511inter3), .O(gate511inter10));
  nor2  gate838(.a(gate511inter10), .b(gate511inter9), .O(gate511inter11));
  nor2  gate839(.a(gate511inter11), .b(gate511inter6), .O(gate511inter12));
  nand2 gate840(.a(gate511inter12), .b(gate511inter1), .O(G1320));

  xor2  gate1457(.a(G1287), .b(G1286), .O(gate512inter0));
  nand2 gate1458(.a(gate512inter0), .b(s_130), .O(gate512inter1));
  and2  gate1459(.a(G1287), .b(G1286), .O(gate512inter2));
  inv1  gate1460(.a(s_130), .O(gate512inter3));
  inv1  gate1461(.a(s_131), .O(gate512inter4));
  nand2 gate1462(.a(gate512inter4), .b(gate512inter3), .O(gate512inter5));
  nor2  gate1463(.a(gate512inter5), .b(gate512inter2), .O(gate512inter6));
  inv1  gate1464(.a(G1286), .O(gate512inter7));
  inv1  gate1465(.a(G1287), .O(gate512inter8));
  nand2 gate1466(.a(gate512inter8), .b(gate512inter7), .O(gate512inter9));
  nand2 gate1467(.a(s_131), .b(gate512inter3), .O(gate512inter10));
  nor2  gate1468(.a(gate512inter10), .b(gate512inter9), .O(gate512inter11));
  nor2  gate1469(.a(gate512inter11), .b(gate512inter6), .O(gate512inter12));
  nand2 gate1470(.a(gate512inter12), .b(gate512inter1), .O(G1321));
nand2 gate513( .a(G1288), .b(G1289), .O(G1322) );
nand2 gate514( .a(G1290), .b(G1291), .O(G1323) );
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule