module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);

input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;//RE__PI;

input s_0,s_1;//RE__ALLOW(00,01,10,11);
input s_2,s_3;//RE__ALLOW(00,01,10,11);
input s_4,s_5;//RE__ALLOW(00,01,10,11);
input s_6,s_7;//RE__ALLOW(00,01,10,11);
input s_8,s_9;//RE__ALLOW(00,01,10,11);
input s_10,s_11;//RE__ALLOW(00,01,10,11);
input s_12,s_13;//RE__ALLOW(00,01,10,11);
input s_14,s_15;//RE__ALLOW(00,01,10,11);
input s_16,s_17;//RE__ALLOW(00,01,10,11);
input s_18,s_19;//RE__ALLOW(00,01,10,11);
input s_20,s_21;//RE__ALLOW(00,01,10,11);
input s_22,s_23;//RE__ALLOW(00,01,10,11);
input s_24,s_25;//RE__ALLOW(00,01,10,11);
input s_26,s_27;//RE__ALLOW(00,01,10,11);
input s_28,s_29;//RE__ALLOW(00,01,10,11);
input s_30,s_31;//RE__ALLOW(00,01,10,11);
input s_32,s_33;//RE__ALLOW(00,01,10,11);
input s_34,s_35;//RE__ALLOW(00,01,10,11);
input s_36,s_37;//RE__ALLOW(00,01,10,11);
input s_38,s_39;//RE__ALLOW(00,01,10,11);
input s_40,s_41;//RE__ALLOW(00,01,10,11);
input s_42,s_43;//RE__ALLOW(00,01,10,11);
input s_44,s_45;//RE__ALLOW(00,01,10,11);
input s_46,s_47;//RE__ALLOW(00,01,10,11);
input s_48,s_49;//RE__ALLOW(00,01,10,11);
input s_50,s_51;//RE__ALLOW(00,01,10,11);
input s_52,s_53;//RE__ALLOW(00,01,10,11);
input s_54,s_55;//RE__ALLOW(00,01,10,11);
input s_56,s_57;//RE__ALLOW(00,01,10,11);
input s_58,s_59;//RE__ALLOW(00,01,10,11);
input s_60,s_61;//RE__ALLOW(00,01,10,11);
input s_62,s_63;//RE__ALLOW(00,01,10,11);
input s_64,s_65;//RE__ALLOW(00,01,10,11);
input s_66,s_67;//RE__ALLOW(00,01,10,11);
input s_68,s_69;//RE__ALLOW(00,01,10,11);
input s_70,s_71;//RE__ALLOW(00,01,10,11);
input s_72,s_73;//RE__ALLOW(00,01,10,11);
input s_74,s_75;//RE__ALLOW(00,01,10,11);
input s_76,s_77;//RE__ALLOW(00,01,10,11);
input s_78,s_79;//RE__ALLOW(00,01,10,11);
input s_80,s_81;//RE__ALLOW(00,01,10,11);
input s_82,s_83;//RE__ALLOW(00,01,10,11);
input s_84,s_85;//RE__ALLOW(00,01,10,11);
input s_86,s_87;//RE__ALLOW(00,01,10,11);
input s_88,s_89;//RE__ALLOW(00,01,10,11);
input s_90,s_91;//RE__ALLOW(00,01,10,11);
input s_92,s_93;//RE__ALLOW(00,01,10,11);
input s_94,s_95;//RE__ALLOW(00,01,10,11);
input s_96,s_97;//RE__ALLOW(00,01,10,11);
input s_98,s_99;//RE__ALLOW(00,01,10,11);
input s_100,s_101;//RE__ALLOW(00,01,10,11);
input s_102,s_103;//RE__ALLOW(00,01,10,11);
input s_104,s_105;//RE__ALLOW(00,01,10,11);
input s_106,s_107;//RE__ALLOW(00,01,10,11);
input s_108,s_109;//RE__ALLOW(00,01,10,11);
input s_110,s_111;//RE__ALLOW(00,01,10,11);
input s_112,s_113;//RE__ALLOW(00,01,10,11);
input s_114,s_115;//RE__ALLOW(00,01,10,11);
input s_116,s_117;//RE__ALLOW(00,01,10,11);
input s_118,s_119;//RE__ALLOW(00,01,10,11);
input s_120,s_121;//RE__ALLOW(00,01,10,11);
input s_122,s_123;//RE__ALLOW(00,01,10,11);
input s_124,s_125;//RE__ALLOW(00,01,10,11);
input s_126,s_127;//RE__ALLOW(00,01,10,11);
input s_128,s_129;//RE__ALLOW(00,01,10,11);
input s_130,s_131;//RE__ALLOW(00,01,10,11);
input s_132,s_133;//RE__ALLOW(00,01,10,11);
input s_134,s_135;//RE__ALLOW(00,01,10,11);
input s_136,s_137;//RE__ALLOW(00,01,10,11);
input s_138,s_139;//RE__ALLOW(00,01,10,11);
input s_140,s_141;//RE__ALLOW(00,01,10,11);
input s_142,s_143;//RE__ALLOW(00,01,10,11);
input s_144,s_145;//RE__ALLOW(00,01,10,11);
input s_146,s_147;//RE__ALLOW(00,01,10,11);
input s_148,s_149;//RE__ALLOW(00,01,10,11);
input s_150,s_151;//RE__ALLOW(00,01,10,11);
input s_152,s_153;//RE__ALLOW(00,01,10,11);
input s_154,s_155;//RE__ALLOW(00,01,10,11);
input s_156,s_157;//RE__ALLOW(00,01,10,11);
input s_158,s_159;//RE__ALLOW(00,01,10,11);
input s_160,s_161;//RE__ALLOW(00,01,10,11);
input s_162,s_163;//RE__ALLOW(00,01,10,11);
input s_164,s_165;//RE__ALLOW(00,01,10,11);
input s_166,s_167;//RE__ALLOW(00,01,10,11);
input s_168,s_169;//RE__ALLOW(00,01,10,11);
input s_170,s_171;//RE__ALLOW(00,01,10,11);
input s_172,s_173;//RE__ALLOW(00,01,10,11);
input s_174,s_175;//RE__ALLOW(00,01,10,11);
input s_176,s_177;//RE__ALLOW(00,01,10,11);
input s_178,s_179;//RE__ALLOW(00,01,10,11);
input s_180,s_181;//RE__ALLOW(00,01,10,11);
input s_182,s_183;//RE__ALLOW(00,01,10,11);
input s_184,s_185;//RE__ALLOW(00,01,10,11);
input s_186,s_187;//RE__ALLOW(00,01,10,11);
input s_188,s_189;//RE__ALLOW(00,01,10,11);
input s_190,s_191;//RE__ALLOW(00,01,10,11);
input s_192,s_193;//RE__ALLOW(00,01,10,11);
input s_194,s_195;//RE__ALLOW(00,01,10,11);
input s_196,s_197;//RE__ALLOW(00,01,10,11);
input s_198,s_199;//RE__ALLOW(00,01,10,11);
input s_200,s_201;//RE__ALLOW(00,01,10,11);
input s_202,s_203;//RE__ALLOW(00,01,10,11);
input s_204,s_205;//RE__ALLOW(00,01,10,11);
input s_206,s_207;//RE__ALLOW(00,01,10,11);
input s_208,s_209;//RE__ALLOW(00,01,10,11);
input s_210,s_211;//RE__ALLOW(00,01,10,11);
input s_212,s_213;//RE__ALLOW(00,01,10,11);
input s_214,s_215;//RE__ALLOW(00,01,10,11);
input s_216,s_217;//RE__ALLOW(00,01,10,11);
input s_218,s_219;//RE__ALLOW(00,01,10,11);
input s_220,s_221;//RE__ALLOW(00,01,10,11);
input s_222,s_223;//RE__ALLOW(00,01,10,11);
input s_224,s_225;//RE__ALLOW(00,01,10,11);
input s_226,s_227;//RE__ALLOW(00,01,10,11);
input s_228,s_229;//RE__ALLOW(00,01,10,11);
input s_230,s_231;//RE__ALLOW(00,01,10,11);
input s_232,s_233;//RE__ALLOW(00,01,10,11);
input s_234,s_235;//RE__ALLOW(00,01,10,11);
input s_236,s_237;//RE__ALLOW(00,01,10,11);
input s_238,s_239;//RE__ALLOW(00,01,10,11);
input s_240,s_241;//RE__ALLOW(00,01,10,11);
input s_242,s_243;//RE__ALLOW(00,01,10,11);
input s_244,s_245;//RE__ALLOW(00,01,10,11);
input s_246,s_247;//RE__ALLOW(00,01,10,11);
input s_248,s_249;//RE__ALLOW(00,01,10,11);
input s_250,s_251;//RE__ALLOW(00,01,10,11);
input s_252,s_253;//RE__ALLOW(00,01,10,11);
input s_254,s_255;//RE__ALLOW(00,01,10,11);
input s_256,s_257;//RE__ALLOW(00,01,10,11);
input s_258,s_259;//RE__ALLOW(00,01,10,11);
input s_260,s_261;//RE__ALLOW(00,01,10,11);
input s_262,s_263;//RE__ALLOW(00,01,10,11);
input s_264,s_265;//RE__ALLOW(00,01,10,11);
input s_266,s_267;//RE__ALLOW(00,01,10,11);
input s_268,s_269;//RE__ALLOW(00,01,10,11);
input s_270,s_271;//RE__ALLOW(00,01,10,11);
input s_272,s_273;//RE__ALLOW(00,01,10,11);
input s_274,s_275;//RE__ALLOW(00,01,10,11);
input s_276,s_277;//RE__ALLOW(00,01,10,11);
input s_278,s_279;//RE__ALLOW(00,01,10,11);
input s_280,s_281;//RE__ALLOW(00,01,10,11);
input s_282,s_283;//RE__ALLOW(00,01,10,11);
input s_284,s_285;//RE__ALLOW(00,01,10,11);
input s_286,s_287;//RE__ALLOW(00,01,10,11);
input s_288,s_289;//RE__ALLOW(00,01,10,11);
input s_290,s_291;//RE__ALLOW(00,01,10,11);
input s_292,s_293;//RE__ALLOW(00,01,10,11);
input s_294,s_295;//RE__ALLOW(00,01,10,11);
input s_296,s_297;//RE__ALLOW(00,01,10,11);
input s_298,s_299;//RE__ALLOW(00,01,10,11);
input s_300,s_301;//RE__ALLOW(00,01,10,11);
input s_302,s_303;//RE__ALLOW(00,01,10,11);
input s_304,s_305;//RE__ALLOW(00,01,10,11);
input s_306,s_307;//RE__ALLOW(00,01,10,11);
input s_308,s_309;//RE__ALLOW(00,01,10,11);
input s_310,s_311;//RE__ALLOW(00,01,10,11);
input s_312,s_313;//RE__ALLOW(00,01,10,11);
input s_314,s_315;//RE__ALLOW(00,01,10,11);
input s_316,s_317;//RE__ALLOW(00,01,10,11);
input s_318,s_319;//RE__ALLOW(00,01,10,11);
input s_320,s_321;//RE__ALLOW(00,01,10,11);
input s_322,s_323;//RE__ALLOW(00,01,10,11);
input s_324,s_325;//RE__ALLOW(00,01,10,11);
input s_326,s_327;//RE__ALLOW(00,01,10,11);
input s_328,s_329;//RE__ALLOW(00,01,10,11);
input s_330,s_331;//RE__ALLOW(00,01,10,11);
input s_332,s_333;//RE__ALLOW(00,01,10,11);
input s_334,s_335;//RE__ALLOW(00,01,10,11);
input s_336,s_337;//RE__ALLOW(00,01,10,11);
input s_338,s_339;//RE__ALLOW(00,01,10,11);
input s_340,s_341;//RE__ALLOW(00,01,10,11);
input s_342,s_343;//RE__ALLOW(00,01,10,11);
input s_344,s_345;//RE__ALLOW(00,01,10,11);
input s_346,s_347;//RE__ALLOW(00,01,10,11);
input s_348,s_349;//RE__ALLOW(00,01,10,11);
input s_350,s_351;//RE__ALLOW(00,01,10,11);
input s_352,s_353;//RE__ALLOW(00,01,10,11);
input s_354,s_355;//RE__ALLOW(00,01,10,11);
input s_356,s_357;//RE__ALLOW(00,01,10,11);
input s_358,s_359;//RE__ALLOW(00,01,10,11);
input s_360,s_361;//RE__ALLOW(00,01,10,11);
input s_362,s_363;//RE__ALLOW(00,01,10,11);
input s_364,s_365;//RE__ALLOW(00,01,10,11);
input s_366,s_367;//RE__ALLOW(00,01,10,11);
input s_368,s_369;//RE__ALLOW(00,01,10,11);
input s_370,s_371;//RE__ALLOW(00,01,10,11);
input s_372,s_373;//RE__ALLOW(00,01,10,11);
input s_374,s_375;//RE__ALLOW(00,01,10,11);
input s_376,s_377;//RE__ALLOW(00,01,10,11);
input s_378,s_379;//RE__ALLOW(00,01,10,11);
input s_380,s_381;//RE__ALLOW(00,01,10,11);
input s_382,s_383;//RE__ALLOW(00,01,10,11);
input s_384,s_385;//RE__ALLOW(00,01,10,11);
input s_386,s_387;//RE__ALLOW(00,01,10,11);
input s_388,s_389;//RE__ALLOW(00,01,10,11);
input s_390,s_391;//RE__ALLOW(00,01,10,11);
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;

  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate494inter0, gate494inter1, gate494inter2, gate494inter3, gate494inter4, gate494inter5, gate494inter6, gate494inter7, gate494inter8, gate494inter9, gate494inter10, gate494inter11, gate494inter12, gate443inter0, gate443inter1, gate443inter2, gate443inter3, gate443inter4, gate443inter5, gate443inter6, gate443inter7, gate443inter8, gate443inter9, gate443inter10, gate443inter11, gate443inter12, gate421inter0, gate421inter1, gate421inter2, gate421inter3, gate421inter4, gate421inter5, gate421inter6, gate421inter7, gate421inter8, gate421inter9, gate421inter10, gate421inter11, gate421inter12, gate428inter0, gate428inter1, gate428inter2, gate428inter3, gate428inter4, gate428inter5, gate428inter6, gate428inter7, gate428inter8, gate428inter9, gate428inter10, gate428inter11, gate428inter12, gate138inter0, gate138inter1, gate138inter2, gate138inter3, gate138inter4, gate138inter5, gate138inter6, gate138inter7, gate138inter8, gate138inter9, gate138inter10, gate138inter11, gate138inter12, gate419inter0, gate419inter1, gate419inter2, gate419inter3, gate419inter4, gate419inter5, gate419inter6, gate419inter7, gate419inter8, gate419inter9, gate419inter10, gate419inter11, gate419inter12, gate66inter0, gate66inter1, gate66inter2, gate66inter3, gate66inter4, gate66inter5, gate66inter6, gate66inter7, gate66inter8, gate66inter9, gate66inter10, gate66inter11, gate66inter12, gate222inter0, gate222inter1, gate222inter2, gate222inter3, gate222inter4, gate222inter5, gate222inter6, gate222inter7, gate222inter8, gate222inter9, gate222inter10, gate222inter11, gate222inter12, gate441inter0, gate441inter1, gate441inter2, gate441inter3, gate441inter4, gate441inter5, gate441inter6, gate441inter7, gate441inter8, gate441inter9, gate441inter10, gate441inter11, gate441inter12, gate94inter0, gate94inter1, gate94inter2, gate94inter3, gate94inter4, gate94inter5, gate94inter6, gate94inter7, gate94inter8, gate94inter9, gate94inter10, gate94inter11, gate94inter12, gate296inter0, gate296inter1, gate296inter2, gate296inter3, gate296inter4, gate296inter5, gate296inter6, gate296inter7, gate296inter8, gate296inter9, gate296inter10, gate296inter11, gate296inter12, gate513inter0, gate513inter1, gate513inter2, gate513inter3, gate513inter4, gate513inter5, gate513inter6, gate513inter7, gate513inter8, gate513inter9, gate513inter10, gate513inter11, gate513inter12, gate82inter0, gate82inter1, gate82inter2, gate82inter3, gate82inter4, gate82inter5, gate82inter6, gate82inter7, gate82inter8, gate82inter9, gate82inter10, gate82inter11, gate82inter12, gate246inter0, gate246inter1, gate246inter2, gate246inter3, gate246inter4, gate246inter5, gate246inter6, gate246inter7, gate246inter8, gate246inter9, gate246inter10, gate246inter11, gate246inter12, gate470inter0, gate470inter1, gate470inter2, gate470inter3, gate470inter4, gate470inter5, gate470inter6, gate470inter7, gate470inter8, gate470inter9, gate470inter10, gate470inter11, gate470inter12, gate407inter0, gate407inter1, gate407inter2, gate407inter3, gate407inter4, gate407inter5, gate407inter6, gate407inter7, gate407inter8, gate407inter9, gate407inter10, gate407inter11, gate407inter12, gate512inter0, gate512inter1, gate512inter2, gate512inter3, gate512inter4, gate512inter5, gate512inter6, gate512inter7, gate512inter8, gate512inter9, gate512inter10, gate512inter11, gate512inter12, gate64inter0, gate64inter1, gate64inter2, gate64inter3, gate64inter4, gate64inter5, gate64inter6, gate64inter7, gate64inter8, gate64inter9, gate64inter10, gate64inter11, gate64inter12, gate11inter0, gate11inter1, gate11inter2, gate11inter3, gate11inter4, gate11inter5, gate11inter6, gate11inter7, gate11inter8, gate11inter9, gate11inter10, gate11inter11, gate11inter12, gate417inter0, gate417inter1, gate417inter2, gate417inter3, gate417inter4, gate417inter5, gate417inter6, gate417inter7, gate417inter8, gate417inter9, gate417inter10, gate417inter11, gate417inter12, gate459inter0, gate459inter1, gate459inter2, gate459inter3, gate459inter4, gate459inter5, gate459inter6, gate459inter7, gate459inter8, gate459inter9, gate459inter10, gate459inter11, gate459inter12, gate41inter0, gate41inter1, gate41inter2, gate41inter3, gate41inter4, gate41inter5, gate41inter6, gate41inter7, gate41inter8, gate41inter9, gate41inter10, gate41inter11, gate41inter12, gate281inter0, gate281inter1, gate281inter2, gate281inter3, gate281inter4, gate281inter5, gate281inter6, gate281inter7, gate281inter8, gate281inter9, gate281inter10, gate281inter11, gate281inter12, gate34inter0, gate34inter1, gate34inter2, gate34inter3, gate34inter4, gate34inter5, gate34inter6, gate34inter7, gate34inter8, gate34inter9, gate34inter10, gate34inter11, gate34inter12, gate198inter0, gate198inter1, gate198inter2, gate198inter3, gate198inter4, gate198inter5, gate198inter6, gate198inter7, gate198inter8, gate198inter9, gate198inter10, gate198inter11, gate198inter12, gate402inter0, gate402inter1, gate402inter2, gate402inter3, gate402inter4, gate402inter5, gate402inter6, gate402inter7, gate402inter8, gate402inter9, gate402inter10, gate402inter11, gate402inter12, gate289inter0, gate289inter1, gate289inter2, gate289inter3, gate289inter4, gate289inter5, gate289inter6, gate289inter7, gate289inter8, gate289inter9, gate289inter10, gate289inter11, gate289inter12, gate473inter0, gate473inter1, gate473inter2, gate473inter3, gate473inter4, gate473inter5, gate473inter6, gate473inter7, gate473inter8, gate473inter9, gate473inter10, gate473inter11, gate473inter12, gate221inter0, gate221inter1, gate221inter2, gate221inter3, gate221inter4, gate221inter5, gate221inter6, gate221inter7, gate221inter8, gate221inter9, gate221inter10, gate221inter11, gate221inter12, gate204inter0, gate204inter1, gate204inter2, gate204inter3, gate204inter4, gate204inter5, gate204inter6, gate204inter7, gate204inter8, gate204inter9, gate204inter10, gate204inter11, gate204inter12, gate190inter0, gate190inter1, gate190inter2, gate190inter3, gate190inter4, gate190inter5, gate190inter6, gate190inter7, gate190inter8, gate190inter9, gate190inter10, gate190inter11, gate190inter12, gate458inter0, gate458inter1, gate458inter2, gate458inter3, gate458inter4, gate458inter5, gate458inter6, gate458inter7, gate458inter8, gate458inter9, gate458inter10, gate458inter11, gate458inter12, gate411inter0, gate411inter1, gate411inter2, gate411inter3, gate411inter4, gate411inter5, gate411inter6, gate411inter7, gate411inter8, gate411inter9, gate411inter10, gate411inter11, gate411inter12, gate159inter0, gate159inter1, gate159inter2, gate159inter3, gate159inter4, gate159inter5, gate159inter6, gate159inter7, gate159inter8, gate159inter9, gate159inter10, gate159inter11, gate159inter12, gate192inter0, gate192inter1, gate192inter2, gate192inter3, gate192inter4, gate192inter5, gate192inter6, gate192inter7, gate192inter8, gate192inter9, gate192inter10, gate192inter11, gate192inter12, gate239inter0, gate239inter1, gate239inter2, gate239inter3, gate239inter4, gate239inter5, gate239inter6, gate239inter7, gate239inter8, gate239inter9, gate239inter10, gate239inter11, gate239inter12, gate217inter0, gate217inter1, gate217inter2, gate217inter3, gate217inter4, gate217inter5, gate217inter6, gate217inter7, gate217inter8, gate217inter9, gate217inter10, gate217inter11, gate217inter12, gate39inter0, gate39inter1, gate39inter2, gate39inter3, gate39inter4, gate39inter5, gate39inter6, gate39inter7, gate39inter8, gate39inter9, gate39inter10, gate39inter11, gate39inter12, gate227inter0, gate227inter1, gate227inter2, gate227inter3, gate227inter4, gate227inter5, gate227inter6, gate227inter7, gate227inter8, gate227inter9, gate227inter10, gate227inter11, gate227inter12, gate475inter0, gate475inter1, gate475inter2, gate475inter3, gate475inter4, gate475inter5, gate475inter6, gate475inter7, gate475inter8, gate475inter9, gate475inter10, gate475inter11, gate475inter12, gate413inter0, gate413inter1, gate413inter2, gate413inter3, gate413inter4, gate413inter5, gate413inter6, gate413inter7, gate413inter8, gate413inter9, gate413inter10, gate413inter11, gate413inter12, gate249inter0, gate249inter1, gate249inter2, gate249inter3, gate249inter4, gate249inter5, gate249inter6, gate249inter7, gate249inter8, gate249inter9, gate249inter10, gate249inter11, gate249inter12, gate98inter0, gate98inter1, gate98inter2, gate98inter3, gate98inter4, gate98inter5, gate98inter6, gate98inter7, gate98inter8, gate98inter9, gate98inter10, gate98inter11, gate98inter12, gate85inter0, gate85inter1, gate85inter2, gate85inter3, gate85inter4, gate85inter5, gate85inter6, gate85inter7, gate85inter8, gate85inter9, gate85inter10, gate85inter11, gate85inter12, gate460inter0, gate460inter1, gate460inter2, gate460inter3, gate460inter4, gate460inter5, gate460inter6, gate460inter7, gate460inter8, gate460inter9, gate460inter10, gate460inter11, gate460inter12, gate15inter0, gate15inter1, gate15inter2, gate15inter3, gate15inter4, gate15inter5, gate15inter6, gate15inter7, gate15inter8, gate15inter9, gate15inter10, gate15inter11, gate15inter12, gate127inter0, gate127inter1, gate127inter2, gate127inter3, gate127inter4, gate127inter5, gate127inter6, gate127inter7, gate127inter8, gate127inter9, gate127inter10, gate127inter11, gate127inter12, gate391inter0, gate391inter1, gate391inter2, gate391inter3, gate391inter4, gate391inter5, gate391inter6, gate391inter7, gate391inter8, gate391inter9, gate391inter10, gate391inter11, gate391inter12, gate425inter0, gate425inter1, gate425inter2, gate425inter3, gate425inter4, gate425inter5, gate425inter6, gate425inter7, gate425inter8, gate425inter9, gate425inter10, gate425inter11, gate425inter12, gate254inter0, gate254inter1, gate254inter2, gate254inter3, gate254inter4, gate254inter5, gate254inter6, gate254inter7, gate254inter8, gate254inter9, gate254inter10, gate254inter11, gate254inter12, gate175inter0, gate175inter1, gate175inter2, gate175inter3, gate175inter4, gate175inter5, gate175inter6, gate175inter7, gate175inter8, gate175inter9, gate175inter10, gate175inter11, gate175inter12, gate251inter0, gate251inter1, gate251inter2, gate251inter3, gate251inter4, gate251inter5, gate251inter6, gate251inter7, gate251inter8, gate251inter9, gate251inter10, gate251inter11, gate251inter12, gate492inter0, gate492inter1, gate492inter2, gate492inter3, gate492inter4, gate492inter5, gate492inter6, gate492inter7, gate492inter8, gate492inter9, gate492inter10, gate492inter11, gate492inter12, gate137inter0, gate137inter1, gate137inter2, gate137inter3, gate137inter4, gate137inter5, gate137inter6, gate137inter7, gate137inter8, gate137inter9, gate137inter10, gate137inter11, gate137inter12, gate178inter0, gate178inter1, gate178inter2, gate178inter3, gate178inter4, gate178inter5, gate178inter6, gate178inter7, gate178inter8, gate178inter9, gate178inter10, gate178inter11, gate178inter12, gate157inter0, gate157inter1, gate157inter2, gate157inter3, gate157inter4, gate157inter5, gate157inter6, gate157inter7, gate157inter8, gate157inter9, gate157inter10, gate157inter11, gate157inter12, gate139inter0, gate139inter1, gate139inter2, gate139inter3, gate139inter4, gate139inter5, gate139inter6, gate139inter7, gate139inter8, gate139inter9, gate139inter10, gate139inter11, gate139inter12, gate185inter0, gate185inter1, gate185inter2, gate185inter3, gate185inter4, gate185inter5, gate185inter6, gate185inter7, gate185inter8, gate185inter9, gate185inter10, gate185inter11, gate185inter12, gate240inter0, gate240inter1, gate240inter2, gate240inter3, gate240inter4, gate240inter5, gate240inter6, gate240inter7, gate240inter8, gate240inter9, gate240inter10, gate240inter11, gate240inter12, gate268inter0, gate268inter1, gate268inter2, gate268inter3, gate268inter4, gate268inter5, gate268inter6, gate268inter7, gate268inter8, gate268inter9, gate268inter10, gate268inter11, gate268inter12, gate117inter0, gate117inter1, gate117inter2, gate117inter3, gate117inter4, gate117inter5, gate117inter6, gate117inter7, gate117inter8, gate117inter9, gate117inter10, gate117inter11, gate117inter12, gate514inter0, gate514inter1, gate514inter2, gate514inter3, gate514inter4, gate514inter5, gate514inter6, gate514inter7, gate514inter8, gate514inter9, gate514inter10, gate514inter11, gate514inter12, gate434inter0, gate434inter1, gate434inter2, gate434inter3, gate434inter4, gate434inter5, gate434inter6, gate434inter7, gate434inter8, gate434inter9, gate434inter10, gate434inter11, gate434inter12, gate129inter0, gate129inter1, gate129inter2, gate129inter3, gate129inter4, gate129inter5, gate129inter6, gate129inter7, gate129inter8, gate129inter9, gate129inter10, gate129inter11, gate129inter12, gate266inter0, gate266inter1, gate266inter2, gate266inter3, gate266inter4, gate266inter5, gate266inter6, gate266inter7, gate266inter8, gate266inter9, gate266inter10, gate266inter11, gate266inter12, gate481inter0, gate481inter1, gate481inter2, gate481inter3, gate481inter4, gate481inter5, gate481inter6, gate481inter7, gate481inter8, gate481inter9, gate481inter10, gate481inter11, gate481inter12, gate244inter0, gate244inter1, gate244inter2, gate244inter3, gate244inter4, gate244inter5, gate244inter6, gate244inter7, gate244inter8, gate244inter9, gate244inter10, gate244inter11, gate244inter12, gate23inter0, gate23inter1, gate23inter2, gate23inter3, gate23inter4, gate23inter5, gate23inter6, gate23inter7, gate23inter8, gate23inter9, gate23inter10, gate23inter11, gate23inter12, gate457inter0, gate457inter1, gate457inter2, gate457inter3, gate457inter4, gate457inter5, gate457inter6, gate457inter7, gate457inter8, gate457inter9, gate457inter10, gate457inter11, gate457inter12, gate245inter0, gate245inter1, gate245inter2, gate245inter3, gate245inter4, gate245inter5, gate245inter6, gate245inter7, gate245inter8, gate245inter9, gate245inter10, gate245inter11, gate245inter12, gate295inter0, gate295inter1, gate295inter2, gate295inter3, gate295inter4, gate295inter5, gate295inter6, gate295inter7, gate295inter8, gate295inter9, gate295inter10, gate295inter11, gate295inter12, gate107inter0, gate107inter1, gate107inter2, gate107inter3, gate107inter4, gate107inter5, gate107inter6, gate107inter7, gate107inter8, gate107inter9, gate107inter10, gate107inter11, gate107inter12, gate135inter0, gate135inter1, gate135inter2, gate135inter3, gate135inter4, gate135inter5, gate135inter6, gate135inter7, gate135inter8, gate135inter9, gate135inter10, gate135inter11, gate135inter12, gate395inter0, gate395inter1, gate395inter2, gate395inter3, gate395inter4, gate395inter5, gate395inter6, gate395inter7, gate395inter8, gate395inter9, gate395inter10, gate395inter11, gate395inter12, gate387inter0, gate387inter1, gate387inter2, gate387inter3, gate387inter4, gate387inter5, gate387inter6, gate387inter7, gate387inter8, gate387inter9, gate387inter10, gate387inter11, gate387inter12, gate261inter0, gate261inter1, gate261inter2, gate261inter3, gate261inter4, gate261inter5, gate261inter6, gate261inter7, gate261inter8, gate261inter9, gate261inter10, gate261inter11, gate261inter12, gate68inter0, gate68inter1, gate68inter2, gate68inter3, gate68inter4, gate68inter5, gate68inter6, gate68inter7, gate68inter8, gate68inter9, gate68inter10, gate68inter11, gate68inter12, gate482inter0, gate482inter1, gate482inter2, gate482inter3, gate482inter4, gate482inter5, gate482inter6, gate482inter7, gate482inter8, gate482inter9, gate482inter10, gate482inter11, gate482inter12, gate272inter0, gate272inter1, gate272inter2, gate272inter3, gate272inter4, gate272inter5, gate272inter6, gate272inter7, gate272inter8, gate272inter9, gate272inter10, gate272inter11, gate272inter12, gate183inter0, gate183inter1, gate183inter2, gate183inter3, gate183inter4, gate183inter5, gate183inter6, gate183inter7, gate183inter8, gate183inter9, gate183inter10, gate183inter11, gate183inter12, gate433inter0, gate433inter1, gate433inter2, gate433inter3, gate433inter4, gate433inter5, gate433inter6, gate433inter7, gate433inter8, gate433inter9, gate433inter10, gate433inter11, gate433inter12, gate191inter0, gate191inter1, gate191inter2, gate191inter3, gate191inter4, gate191inter5, gate191inter6, gate191inter7, gate191inter8, gate191inter9, gate191inter10, gate191inter11, gate191inter12, gate10inter0, gate10inter1, gate10inter2, gate10inter3, gate10inter4, gate10inter5, gate10inter6, gate10inter7, gate10inter8, gate10inter9, gate10inter10, gate10inter11, gate10inter12, gate20inter0, gate20inter1, gate20inter2, gate20inter3, gate20inter4, gate20inter5, gate20inter6, gate20inter7, gate20inter8, gate20inter9, gate20inter10, gate20inter11, gate20inter12, gate396inter0, gate396inter1, gate396inter2, gate396inter3, gate396inter4, gate396inter5, gate396inter6, gate396inter7, gate396inter8, gate396inter9, gate396inter10, gate396inter11, gate396inter12, gate90inter0, gate90inter1, gate90inter2, gate90inter3, gate90inter4, gate90inter5, gate90inter6, gate90inter7, gate90inter8, gate90inter9, gate90inter10, gate90inter11, gate90inter12, gate49inter0, gate49inter1, gate49inter2, gate49inter3, gate49inter4, gate49inter5, gate49inter6, gate49inter7, gate49inter8, gate49inter9, gate49inter10, gate49inter11, gate49inter12, gate76inter0, gate76inter1, gate76inter2, gate76inter3, gate76inter4, gate76inter5, gate76inter6, gate76inter7, gate76inter8, gate76inter9, gate76inter10, gate76inter11, gate76inter12, gate173inter0, gate173inter1, gate173inter2, gate173inter3, gate173inter4, gate173inter5, gate173inter6, gate173inter7, gate173inter8, gate173inter9, gate173inter10, gate173inter11, gate173inter12, gate445inter0, gate445inter1, gate445inter2, gate445inter3, gate445inter4, gate445inter5, gate445inter6, gate445inter7, gate445inter8, gate445inter9, gate445inter10, gate445inter11, gate445inter12, gate225inter0, gate225inter1, gate225inter2, gate225inter3, gate225inter4, gate225inter5, gate225inter6, gate225inter7, gate225inter8, gate225inter9, gate225inter10, gate225inter11, gate225inter12, gate150inter0, gate150inter1, gate150inter2, gate150inter3, gate150inter4, gate150inter5, gate150inter6, gate150inter7, gate150inter8, gate150inter9, gate150inter10, gate150inter11, gate150inter12, gate168inter0, gate168inter1, gate168inter2, gate168inter3, gate168inter4, gate168inter5, gate168inter6, gate168inter7, gate168inter8, gate168inter9, gate168inter10, gate168inter11, gate168inter12, gate142inter0, gate142inter1, gate142inter2, gate142inter3, gate142inter4, gate142inter5, gate142inter6, gate142inter7, gate142inter8, gate142inter9, gate142inter10, gate142inter11, gate142inter12, gate279inter0, gate279inter1, gate279inter2, gate279inter3, gate279inter4, gate279inter5, gate279inter6, gate279inter7, gate279inter8, gate279inter9, gate279inter10, gate279inter11, gate279inter12, gate415inter0, gate415inter1, gate415inter2, gate415inter3, gate415inter4, gate415inter5, gate415inter6, gate415inter7, gate415inter8, gate415inter9, gate415inter10, gate415inter11, gate415inter12, gate483inter0, gate483inter1, gate483inter2, gate483inter3, gate483inter4, gate483inter5, gate483inter6, gate483inter7, gate483inter8, gate483inter9, gate483inter10, gate483inter11, gate483inter12, gate287inter0, gate287inter1, gate287inter2, gate287inter3, gate287inter4, gate287inter5, gate287inter6, gate287inter7, gate287inter8, gate287inter9, gate287inter10, gate287inter11, gate287inter12, gate70inter0, gate70inter1, gate70inter2, gate70inter3, gate70inter4, gate70inter5, gate70inter6, gate70inter7, gate70inter8, gate70inter9, gate70inter10, gate70inter11, gate70inter12, gate203inter0, gate203inter1, gate203inter2, gate203inter3, gate203inter4, gate203inter5, gate203inter6, gate203inter7, gate203inter8, gate203inter9, gate203inter10, gate203inter11, gate203inter12, gate110inter0, gate110inter1, gate110inter2, gate110inter3, gate110inter4, gate110inter5, gate110inter6, gate110inter7, gate110inter8, gate110inter9, gate110inter10, gate110inter11, gate110inter12, gate89inter0, gate89inter1, gate89inter2, gate89inter3, gate89inter4, gate89inter5, gate89inter6, gate89inter7, gate89inter8, gate89inter9, gate89inter10, gate89inter11, gate89inter12, gate278inter0, gate278inter1, gate278inter2, gate278inter3, gate278inter4, gate278inter5, gate278inter6, gate278inter7, gate278inter8, gate278inter9, gate278inter10, gate278inter11, gate278inter12, gate462inter0, gate462inter1, gate462inter2, gate462inter3, gate462inter4, gate462inter5, gate462inter6, gate462inter7, gate462inter8, gate462inter9, gate462inter10, gate462inter11, gate462inter12, gate211inter0, gate211inter1, gate211inter2, gate211inter3, gate211inter4, gate211inter5, gate211inter6, gate211inter7, gate211inter8, gate211inter9, gate211inter10, gate211inter11, gate211inter12, gate40inter0, gate40inter1, gate40inter2, gate40inter3, gate40inter4, gate40inter5, gate40inter6, gate40inter7, gate40inter8, gate40inter9, gate40inter10, gate40inter11, gate40inter12, gate9inter0, gate9inter1, gate9inter2, gate9inter3, gate9inter4, gate9inter5, gate9inter6, gate9inter7, gate9inter8, gate9inter9, gate9inter10, gate9inter11, gate9inter12, gate102inter0, gate102inter1, gate102inter2, gate102inter3, gate102inter4, gate102inter5, gate102inter6, gate102inter7, gate102inter8, gate102inter9, gate102inter10, gate102inter11, gate102inter12, gate501inter0, gate501inter1, gate501inter2, gate501inter3, gate501inter4, gate501inter5, gate501inter6, gate501inter7, gate501inter8, gate501inter9, gate501inter10, gate501inter11, gate501inter12, gate162inter0, gate162inter1, gate162inter2, gate162inter3, gate162inter4, gate162inter5, gate162inter6, gate162inter7, gate162inter8, gate162inter9, gate162inter10, gate162inter11, gate162inter12, gate493inter0, gate493inter1, gate493inter2, gate493inter3, gate493inter4, gate493inter5, gate493inter6, gate493inter7, gate493inter8, gate493inter9, gate493inter10, gate493inter11, gate493inter12, gate453inter0, gate453inter1, gate453inter2, gate453inter3, gate453inter4, gate453inter5, gate453inter6, gate453inter7, gate453inter8, gate453inter9, gate453inter10, gate453inter11, gate453inter12, gate31inter0, gate31inter1, gate31inter2, gate31inter3, gate31inter4, gate31inter5, gate31inter6, gate31inter7, gate31inter8, gate31inter9, gate31inter10, gate31inter11, gate31inter12, gate27inter0, gate27inter1, gate27inter2, gate27inter3, gate27inter4, gate27inter5, gate27inter6, gate27inter7, gate27inter8, gate27inter9, gate27inter10, gate27inter11, gate27inter12, gate12inter0, gate12inter1, gate12inter2, gate12inter3, gate12inter4, gate12inter5, gate12inter6, gate12inter7, gate12inter8, gate12inter9, gate12inter10, gate12inter11, gate12inter12, gate194inter0, gate194inter1, gate194inter2, gate194inter3, gate194inter4, gate194inter5, gate194inter6, gate194inter7, gate194inter8, gate194inter9, gate194inter10, gate194inter11, gate194inter12, gate509inter0, gate509inter1, gate509inter2, gate509inter3, gate509inter4, gate509inter5, gate509inter6, gate509inter7, gate509inter8, gate509inter9, gate509inter10, gate509inter11, gate509inter12, gate426inter0, gate426inter1, gate426inter2, gate426inter3, gate426inter4, gate426inter5, gate426inter6, gate426inter7, gate426inter8, gate426inter9, gate426inter10, gate426inter11, gate426inter12, gate103inter0, gate103inter1, gate103inter2, gate103inter3, gate103inter4, gate103inter5, gate103inter6, gate103inter7, gate103inter8, gate103inter9, gate103inter10, gate103inter11, gate103inter12, gate126inter0, gate126inter1, gate126inter2, gate126inter3, gate126inter4, gate126inter5, gate126inter6, gate126inter7, gate126inter8, gate126inter9, gate126inter10, gate126inter11, gate126inter12, gate394inter0, gate394inter1, gate394inter2, gate394inter3, gate394inter4, gate394inter5, gate394inter6, gate394inter7, gate394inter8, gate394inter9, gate394inter10, gate394inter11, gate394inter12, gate62inter0, gate62inter1, gate62inter2, gate62inter3, gate62inter4, gate62inter5, gate62inter6, gate62inter7, gate62inter8, gate62inter9, gate62inter10, gate62inter11, gate62inter12, gate248inter0, gate248inter1, gate248inter2, gate248inter3, gate248inter4, gate248inter5, gate248inter6, gate248inter7, gate248inter8, gate248inter9, gate248inter10, gate248inter11, gate248inter12, gate147inter0, gate147inter1, gate147inter2, gate147inter3, gate147inter4, gate147inter5, gate147inter6, gate147inter7, gate147inter8, gate147inter9, gate147inter10, gate147inter11, gate147inter12, gate154inter0, gate154inter1, gate154inter2, gate154inter3, gate154inter4, gate154inter5, gate154inter6, gate154inter7, gate154inter8, gate154inter9, gate154inter10, gate154inter11, gate154inter12, gate104inter0, gate104inter1, gate104inter2, gate104inter3, gate104inter4, gate104inter5, gate104inter6, gate104inter7, gate104inter8, gate104inter9, gate104inter10, gate104inter11, gate104inter12, gate13inter0, gate13inter1, gate13inter2, gate13inter3, gate13inter4, gate13inter5, gate13inter6, gate13inter7, gate13inter8, gate13inter9, gate13inter10, gate13inter11, gate13inter12, gate488inter0, gate488inter1, gate488inter2, gate488inter3, gate488inter4, gate488inter5, gate488inter6, gate488inter7, gate488inter8, gate488inter9, gate488inter10, gate488inter11, gate488inter12, gate467inter0, gate467inter1, gate467inter2, gate467inter3, gate467inter4, gate467inter5, gate467inter6, gate467inter7, gate467inter8, gate467inter9, gate467inter10, gate467inter11, gate467inter12, gate99inter0, gate99inter1, gate99inter2, gate99inter3, gate99inter4, gate99inter5, gate99inter6, gate99inter7, gate99inter8, gate99inter9, gate99inter10, gate99inter11, gate99inter12, gate215inter0, gate215inter1, gate215inter2, gate215inter3, gate215inter4, gate215inter5, gate215inter6, gate215inter7, gate215inter8, gate215inter9, gate215inter10, gate215inter11, gate215inter12, gate14inter0, gate14inter1, gate14inter2, gate14inter3, gate14inter4, gate14inter5, gate14inter6, gate14inter7, gate14inter8, gate14inter9, gate14inter10, gate14inter11, gate14inter12, gate38inter0, gate38inter1, gate38inter2, gate38inter3, gate38inter4, gate38inter5, gate38inter6, gate38inter7, gate38inter8, gate38inter9, gate38inter10, gate38inter11, gate38inter12, gate269inter0, gate269inter1, gate269inter2, gate269inter3, gate269inter4, gate269inter5, gate269inter6, gate269inter7, gate269inter8, gate269inter9, gate269inter10, gate269inter11, gate269inter12, gate179inter0, gate179inter1, gate179inter2, gate179inter3, gate179inter4, gate179inter5, gate179inter6, gate179inter7, gate179inter8, gate179inter9, gate179inter10, gate179inter11, gate179inter12, gate435inter0, gate435inter1, gate435inter2, gate435inter3, gate435inter4, gate435inter5, gate435inter6, gate435inter7, gate435inter8, gate435inter9, gate435inter10, gate435inter11, gate435inter12, gate409inter0, gate409inter1, gate409inter2, gate409inter3, gate409inter4, gate409inter5, gate409inter6, gate409inter7, gate409inter8, gate409inter9, gate409inter10, gate409inter11, gate409inter12, gate444inter0, gate444inter1, gate444inter2, gate444inter3, gate444inter4, gate444inter5, gate444inter6, gate444inter7, gate444inter8, gate444inter9, gate444inter10, gate444inter11, gate444inter12, gate271inter0, gate271inter1, gate271inter2, gate271inter3, gate271inter4, gate271inter5, gate271inter6, gate271inter7, gate271inter8, gate271inter9, gate271inter10, gate271inter11, gate271inter12, gate250inter0, gate250inter1, gate250inter2, gate250inter3, gate250inter4, gate250inter5, gate250inter6, gate250inter7, gate250inter8, gate250inter9, gate250inter10, gate250inter11, gate250inter12, gate47inter0, gate47inter1, gate47inter2, gate47inter3, gate47inter4, gate47inter5, gate47inter6, gate47inter7, gate47inter8, gate47inter9, gate47inter10, gate47inter11, gate47inter12, gate510inter0, gate510inter1, gate510inter2, gate510inter3, gate510inter4, gate510inter5, gate510inter6, gate510inter7, gate510inter8, gate510inter9, gate510inter10, gate510inter11, gate510inter12, gate241inter0, gate241inter1, gate241inter2, gate241inter3, gate241inter4, gate241inter5, gate241inter6, gate241inter7, gate241inter8, gate241inter9, gate241inter10, gate241inter11, gate241inter12, gate404inter0, gate404inter1, gate404inter2, gate404inter3, gate404inter4, gate404inter5, gate404inter6, gate404inter7, gate404inter8, gate404inter9, gate404inter10, gate404inter11, gate404inter12, gate430inter0, gate430inter1, gate430inter2, gate430inter3, gate430inter4, gate430inter5, gate430inter6, gate430inter7, gate430inter8, gate430inter9, gate430inter10, gate430inter11, gate430inter12, gate37inter0, gate37inter1, gate37inter2, gate37inter3, gate37inter4, gate37inter5, gate37inter6, gate37inter7, gate37inter8, gate37inter9, gate37inter10, gate37inter11, gate37inter12, gate195inter0, gate195inter1, gate195inter2, gate195inter3, gate195inter4, gate195inter5, gate195inter6, gate195inter7, gate195inter8, gate195inter9, gate195inter10, gate195inter11, gate195inter12, gate155inter0, gate155inter1, gate155inter2, gate155inter3, gate155inter4, gate155inter5, gate155inter6, gate155inter7, gate155inter8, gate155inter9, gate155inter10, gate155inter11, gate155inter12, gate88inter0, gate88inter1, gate88inter2, gate88inter3, gate88inter4, gate88inter5, gate88inter6, gate88inter7, gate88inter8, gate88inter9, gate88inter10, gate88inter11, gate88inter12, gate292inter0, gate292inter1, gate292inter2, gate292inter3, gate292inter4, gate292inter5, gate292inter6, gate292inter7, gate292inter8, gate292inter9, gate292inter10, gate292inter11, gate292inter12, gate188inter0, gate188inter1, gate188inter2, gate188inter3, gate188inter4, gate188inter5, gate188inter6, gate188inter7, gate188inter8, gate188inter9, gate188inter10, gate188inter11, gate188inter12, gate234inter0, gate234inter1, gate234inter2, gate234inter3, gate234inter4, gate234inter5, gate234inter6, gate234inter7, gate234inter8, gate234inter9, gate234inter10, gate234inter11, gate234inter12, gate449inter0, gate449inter1, gate449inter2, gate449inter3, gate449inter4, gate449inter5, gate449inter6, gate449inter7, gate449inter8, gate449inter9, gate449inter10, gate449inter11, gate449inter12, gate485inter0, gate485inter1, gate485inter2, gate485inter3, gate485inter4, gate485inter5, gate485inter6, gate485inter7, gate485inter8, gate485inter9, gate485inter10, gate485inter11, gate485inter12, gate143inter0, gate143inter1, gate143inter2, gate143inter3, gate143inter4, gate143inter5, gate143inter6, gate143inter7, gate143inter8, gate143inter9, gate143inter10, gate143inter11, gate143inter12, gate410inter0, gate410inter1, gate410inter2, gate410inter3, gate410inter4, gate410inter5, gate410inter6, gate410inter7, gate410inter8, gate410inter9, gate410inter10, gate410inter11, gate410inter12, gate270inter0, gate270inter1, gate270inter2, gate270inter3, gate270inter4, gate270inter5, gate270inter6, gate270inter7, gate270inter8, gate270inter9, gate270inter10, gate270inter11, gate270inter12, gate216inter0, gate216inter1, gate216inter2, gate216inter3, gate216inter4, gate216inter5, gate216inter6, gate216inter7, gate216inter8, gate216inter9, gate216inter10, gate216inter11, gate216inter12, gate506inter0, gate506inter1, gate506inter2, gate506inter3, gate506inter4, gate506inter5, gate506inter6, gate506inter7, gate506inter8, gate506inter9, gate506inter10, gate506inter11, gate506inter12, gate219inter0, gate219inter1, gate219inter2, gate219inter3, gate219inter4, gate219inter5, gate219inter6, gate219inter7, gate219inter8, gate219inter9, gate219inter10, gate219inter11, gate219inter12, gate111inter0, gate111inter1, gate111inter2, gate111inter3, gate111inter4, gate111inter5, gate111inter6, gate111inter7, gate111inter8, gate111inter9, gate111inter10, gate111inter11, gate111inter12, gate400inter0, gate400inter1, gate400inter2, gate400inter3, gate400inter4, gate400inter5, gate400inter6, gate400inter7, gate400inter8, gate400inter9, gate400inter10, gate400inter11, gate400inter12, gate128inter0, gate128inter1, gate128inter2, gate128inter3, gate128inter4, gate128inter5, gate128inter6, gate128inter7, gate128inter8, gate128inter9, gate128inter10, gate128inter11, gate128inter12, gate160inter0, gate160inter1, gate160inter2, gate160inter3, gate160inter4, gate160inter5, gate160inter6, gate160inter7, gate160inter8, gate160inter9, gate160inter10, gate160inter11, gate160inter12, gate463inter0, gate463inter1, gate463inter2, gate463inter3, gate463inter4, gate463inter5, gate463inter6, gate463inter7, gate463inter8, gate463inter9, gate463inter10, gate463inter11, gate463inter12, gate247inter0, gate247inter1, gate247inter2, gate247inter3, gate247inter4, gate247inter5, gate247inter6, gate247inter7, gate247inter8, gate247inter9, gate247inter10, gate247inter11, gate247inter12, gate461inter0, gate461inter1, gate461inter2, gate461inter3, gate461inter4, gate461inter5, gate461inter6, gate461inter7, gate461inter8, gate461inter9, gate461inter10, gate461inter11, gate461inter12, gate123inter0, gate123inter1, gate123inter2, gate123inter3, gate123inter4, gate123inter5, gate123inter6, gate123inter7, gate123inter8, gate123inter9, gate123inter10, gate123inter11, gate123inter12, gate446inter0, gate446inter1, gate446inter2, gate446inter3, gate446inter4, gate446inter5, gate446inter6, gate446inter7, gate446inter8, gate446inter9, gate446inter10, gate446inter11, gate446inter12, gate101inter0, gate101inter1, gate101inter2, gate101inter3, gate101inter4, gate101inter5, gate101inter6, gate101inter7, gate101inter8, gate101inter9, gate101inter10, gate101inter11, gate101inter12, gate96inter0, gate96inter1, gate96inter2, gate96inter3, gate96inter4, gate96inter5, gate96inter6, gate96inter7, gate96inter8, gate96inter9, gate96inter10, gate96inter11, gate96inter12, gate422inter0, gate422inter1, gate422inter2, gate422inter3, gate422inter4, gate422inter5, gate422inter6, gate422inter7, gate422inter8, gate422inter9, gate422inter10, gate422inter11, gate422inter12, gate130inter0, gate130inter1, gate130inter2, gate130inter3, gate130inter4, gate130inter5, gate130inter6, gate130inter7, gate130inter8, gate130inter9, gate130inter10, gate130inter11, gate130inter12, gate84inter0, gate84inter1, gate84inter2, gate84inter3, gate84inter4, gate84inter5, gate84inter6, gate84inter7, gate84inter8, gate84inter9, gate84inter10, gate84inter11, gate84inter12, gate69inter0, gate69inter1, gate69inter2, gate69inter3, gate69inter4, gate69inter5, gate69inter6, gate69inter7, gate69inter8, gate69inter9, gate69inter10, gate69inter11, gate69inter12, gate447inter0, gate447inter1, gate447inter2, gate447inter3, gate447inter4, gate447inter5, gate447inter6, gate447inter7, gate447inter8, gate447inter9, gate447inter10, gate447inter11, gate447inter12, gate171inter0, gate171inter1, gate171inter2, gate171inter3, gate171inter4, gate171inter5, gate171inter6, gate171inter7, gate171inter8, gate171inter9, gate171inter10, gate171inter11, gate171inter12, gate264inter0, gate264inter1, gate264inter2, gate264inter3, gate264inter4, gate264inter5, gate264inter6, gate264inter7, gate264inter8, gate264inter9, gate264inter10, gate264inter11, gate264inter12, gate86inter0, gate86inter1, gate86inter2, gate86inter3, gate86inter4, gate86inter5, gate86inter6, gate86inter7, gate86inter8, gate86inter9, gate86inter10, gate86inter11, gate86inter12, gate416inter0, gate416inter1, gate416inter2, gate416inter3, gate416inter4, gate416inter5, gate416inter6, gate416inter7, gate416inter8, gate416inter9, gate416inter10, gate416inter11, gate416inter12, gate24inter0, gate24inter1, gate24inter2, gate24inter3, gate24inter4, gate24inter5, gate24inter6, gate24inter7, gate24inter8, gate24inter9, gate24inter10, gate24inter11, gate24inter12, gate405inter0, gate405inter1, gate405inter2, gate405inter3, gate405inter4, gate405inter5, gate405inter6, gate405inter7, gate405inter8, gate405inter9, gate405inter10, gate405inter11, gate405inter12, gate79inter0, gate79inter1, gate79inter2, gate79inter3, gate79inter4, gate79inter5, gate79inter6, gate79inter7, gate79inter8, gate79inter9, gate79inter10, gate79inter11, gate79inter12, gate502inter0, gate502inter1, gate502inter2, gate502inter3, gate502inter4, gate502inter5, gate502inter6, gate502inter7, gate502inter8, gate502inter9, gate502inter10, gate502inter11, gate502inter12, gate399inter0, gate399inter1, gate399inter2, gate399inter3, gate399inter4, gate399inter5, gate399inter6, gate399inter7, gate399inter8, gate399inter9, gate399inter10, gate399inter11, gate399inter12, gate392inter0, gate392inter1, gate392inter2, gate392inter3, gate392inter4, gate392inter5, gate392inter6, gate392inter7, gate392inter8, gate392inter9, gate392inter10, gate392inter11, gate392inter12, gate124inter0, gate124inter1, gate124inter2, gate124inter3, gate124inter4, gate124inter5, gate124inter6, gate124inter7, gate124inter8, gate124inter9, gate124inter10, gate124inter11, gate124inter12, gate83inter0, gate83inter1, gate83inter2, gate83inter3, gate83inter4, gate83inter5, gate83inter6, gate83inter7, gate83inter8, gate83inter9, gate83inter10, gate83inter11, gate83inter12, gate507inter0, gate507inter1, gate507inter2, gate507inter3, gate507inter4, gate507inter5, gate507inter6, gate507inter7, gate507inter8, gate507inter9, gate507inter10, gate507inter11, gate507inter12, gate468inter0, gate468inter1, gate468inter2, gate468inter3, gate468inter4, gate468inter5, gate468inter6, gate468inter7, gate468inter8, gate468inter9, gate468inter10, gate468inter11, gate468inter12, gate496inter0, gate496inter1, gate496inter2, gate496inter3, gate496inter4, gate496inter5, gate496inter6, gate496inter7, gate496inter8, gate496inter9, gate496inter10, gate496inter11, gate496inter12, gate438inter0, gate438inter1, gate438inter2, gate438inter3, gate438inter4, gate438inter5, gate438inter6, gate438inter7, gate438inter8, gate438inter9, gate438inter10, gate438inter11, gate438inter12, gate202inter0, gate202inter1, gate202inter2, gate202inter3, gate202inter4, gate202inter5, gate202inter6, gate202inter7, gate202inter8, gate202inter9, gate202inter10, gate202inter11, gate202inter12, gate153inter0, gate153inter1, gate153inter2, gate153inter3, gate153inter4, gate153inter5, gate153inter6, gate153inter7, gate153inter8, gate153inter9, gate153inter10, gate153inter11, gate153inter12, gate167inter0, gate167inter1, gate167inter2, gate167inter3, gate167inter4, gate167inter5, gate167inter6, gate167inter7, gate167inter8, gate167inter9, gate167inter10, gate167inter11, gate167inter12, gate177inter0, gate177inter1, gate177inter2, gate177inter3, gate177inter4, gate177inter5, gate177inter6, gate177inter7, gate177inter8, gate177inter9, gate177inter10, gate177inter11, gate177inter12;



and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );

  xor2  gate2031(.a(G2), .b(G1), .O(gate9inter0));
  nand2 gate2032(.a(gate9inter0), .b(s_212), .O(gate9inter1));
  and2  gate2033(.a(G2), .b(G1), .O(gate9inter2));
  inv1  gate2034(.a(s_212), .O(gate9inter3));
  inv1  gate2035(.a(s_213), .O(gate9inter4));
  nand2 gate2036(.a(gate9inter4), .b(gate9inter3), .O(gate9inter5));
  nor2  gate2037(.a(gate9inter5), .b(gate9inter2), .O(gate9inter6));
  inv1  gate2038(.a(G1), .O(gate9inter7));
  inv1  gate2039(.a(G2), .O(gate9inter8));
  nand2 gate2040(.a(gate9inter8), .b(gate9inter7), .O(gate9inter9));
  nand2 gate2041(.a(s_213), .b(gate9inter3), .O(gate9inter10));
  nor2  gate2042(.a(gate9inter10), .b(gate9inter9), .O(gate9inter11));
  nor2  gate2043(.a(gate9inter11), .b(gate9inter6), .O(gate9inter12));
  nand2 gate2044(.a(gate9inter12), .b(gate9inter1), .O(G266));

  xor2  gate1695(.a(G4), .b(G3), .O(gate10inter0));
  nand2 gate1696(.a(gate10inter0), .b(s_164), .O(gate10inter1));
  and2  gate1697(.a(G4), .b(G3), .O(gate10inter2));
  inv1  gate1698(.a(s_164), .O(gate10inter3));
  inv1  gate1699(.a(s_165), .O(gate10inter4));
  nand2 gate1700(.a(gate10inter4), .b(gate10inter3), .O(gate10inter5));
  nor2  gate1701(.a(gate10inter5), .b(gate10inter2), .O(gate10inter6));
  inv1  gate1702(.a(G3), .O(gate10inter7));
  inv1  gate1703(.a(G4), .O(gate10inter8));
  nand2 gate1704(.a(gate10inter8), .b(gate10inter7), .O(gate10inter9));
  nand2 gate1705(.a(s_165), .b(gate10inter3), .O(gate10inter10));
  nor2  gate1706(.a(gate10inter10), .b(gate10inter9), .O(gate10inter11));
  nor2  gate1707(.a(gate10inter11), .b(gate10inter6), .O(gate10inter12));
  nand2 gate1708(.a(gate10inter12), .b(gate10inter1), .O(G269));

  xor2  gate799(.a(G6), .b(G5), .O(gate11inter0));
  nand2 gate800(.a(gate11inter0), .b(s_36), .O(gate11inter1));
  and2  gate801(.a(G6), .b(G5), .O(gate11inter2));
  inv1  gate802(.a(s_36), .O(gate11inter3));
  inv1  gate803(.a(s_37), .O(gate11inter4));
  nand2 gate804(.a(gate11inter4), .b(gate11inter3), .O(gate11inter5));
  nor2  gate805(.a(gate11inter5), .b(gate11inter2), .O(gate11inter6));
  inv1  gate806(.a(G5), .O(gate11inter7));
  inv1  gate807(.a(G6), .O(gate11inter8));
  nand2 gate808(.a(gate11inter8), .b(gate11inter7), .O(gate11inter9));
  nand2 gate809(.a(s_37), .b(gate11inter3), .O(gate11inter10));
  nor2  gate810(.a(gate11inter10), .b(gate11inter9), .O(gate11inter11));
  nor2  gate811(.a(gate11inter11), .b(gate11inter6), .O(gate11inter12));
  nand2 gate812(.a(gate11inter12), .b(gate11inter1), .O(G272));

  xor2  gate2143(.a(G8), .b(G7), .O(gate12inter0));
  nand2 gate2144(.a(gate12inter0), .b(s_228), .O(gate12inter1));
  and2  gate2145(.a(G8), .b(G7), .O(gate12inter2));
  inv1  gate2146(.a(s_228), .O(gate12inter3));
  inv1  gate2147(.a(s_229), .O(gate12inter4));
  nand2 gate2148(.a(gate12inter4), .b(gate12inter3), .O(gate12inter5));
  nor2  gate2149(.a(gate12inter5), .b(gate12inter2), .O(gate12inter6));
  inv1  gate2150(.a(G7), .O(gate12inter7));
  inv1  gate2151(.a(G8), .O(gate12inter8));
  nand2 gate2152(.a(gate12inter8), .b(gate12inter7), .O(gate12inter9));
  nand2 gate2153(.a(s_229), .b(gate12inter3), .O(gate12inter10));
  nor2  gate2154(.a(gate12inter10), .b(gate12inter9), .O(gate12inter11));
  nor2  gate2155(.a(gate12inter11), .b(gate12inter6), .O(gate12inter12));
  nand2 gate2156(.a(gate12inter12), .b(gate12inter1), .O(G275));

  xor2  gate2311(.a(G10), .b(G9), .O(gate13inter0));
  nand2 gate2312(.a(gate13inter0), .b(s_252), .O(gate13inter1));
  and2  gate2313(.a(G10), .b(G9), .O(gate13inter2));
  inv1  gate2314(.a(s_252), .O(gate13inter3));
  inv1  gate2315(.a(s_253), .O(gate13inter4));
  nand2 gate2316(.a(gate13inter4), .b(gate13inter3), .O(gate13inter5));
  nor2  gate2317(.a(gate13inter5), .b(gate13inter2), .O(gate13inter6));
  inv1  gate2318(.a(G9), .O(gate13inter7));
  inv1  gate2319(.a(G10), .O(gate13inter8));
  nand2 gate2320(.a(gate13inter8), .b(gate13inter7), .O(gate13inter9));
  nand2 gate2321(.a(s_253), .b(gate13inter3), .O(gate13inter10));
  nor2  gate2322(.a(gate13inter10), .b(gate13inter9), .O(gate13inter11));
  nor2  gate2323(.a(gate13inter11), .b(gate13inter6), .O(gate13inter12));
  nand2 gate2324(.a(gate13inter12), .b(gate13inter1), .O(G278));

  xor2  gate2381(.a(G12), .b(G11), .O(gate14inter0));
  nand2 gate2382(.a(gate14inter0), .b(s_262), .O(gate14inter1));
  and2  gate2383(.a(G12), .b(G11), .O(gate14inter2));
  inv1  gate2384(.a(s_262), .O(gate14inter3));
  inv1  gate2385(.a(s_263), .O(gate14inter4));
  nand2 gate2386(.a(gate14inter4), .b(gate14inter3), .O(gate14inter5));
  nor2  gate2387(.a(gate14inter5), .b(gate14inter2), .O(gate14inter6));
  inv1  gate2388(.a(G11), .O(gate14inter7));
  inv1  gate2389(.a(G12), .O(gate14inter8));
  nand2 gate2390(.a(gate14inter8), .b(gate14inter7), .O(gate14inter9));
  nand2 gate2391(.a(s_263), .b(gate14inter3), .O(gate14inter10));
  nor2  gate2392(.a(gate14inter10), .b(gate14inter9), .O(gate14inter11));
  nor2  gate2393(.a(gate14inter11), .b(gate14inter6), .O(gate14inter12));
  nand2 gate2394(.a(gate14inter12), .b(gate14inter1), .O(G281));

  xor2  gate1177(.a(G14), .b(G13), .O(gate15inter0));
  nand2 gate1178(.a(gate15inter0), .b(s_90), .O(gate15inter1));
  and2  gate1179(.a(G14), .b(G13), .O(gate15inter2));
  inv1  gate1180(.a(s_90), .O(gate15inter3));
  inv1  gate1181(.a(s_91), .O(gate15inter4));
  nand2 gate1182(.a(gate15inter4), .b(gate15inter3), .O(gate15inter5));
  nor2  gate1183(.a(gate15inter5), .b(gate15inter2), .O(gate15inter6));
  inv1  gate1184(.a(G13), .O(gate15inter7));
  inv1  gate1185(.a(G14), .O(gate15inter8));
  nand2 gate1186(.a(gate15inter8), .b(gate15inter7), .O(gate15inter9));
  nand2 gate1187(.a(s_91), .b(gate15inter3), .O(gate15inter10));
  nor2  gate1188(.a(gate15inter10), .b(gate15inter9), .O(gate15inter11));
  nor2  gate1189(.a(gate15inter11), .b(gate15inter6), .O(gate15inter12));
  nand2 gate1190(.a(gate15inter12), .b(gate15inter1), .O(G284));
nand2 gate16( .a(G15), .b(G16), .O(G287) );
nand2 gate17( .a(G17), .b(G18), .O(G290) );
nand2 gate18( .a(G19), .b(G20), .O(G293) );
nand2 gate19( .a(G21), .b(G22), .O(G296) );

  xor2  gate1709(.a(G24), .b(G23), .O(gate20inter0));
  nand2 gate1710(.a(gate20inter0), .b(s_166), .O(gate20inter1));
  and2  gate1711(.a(G24), .b(G23), .O(gate20inter2));
  inv1  gate1712(.a(s_166), .O(gate20inter3));
  inv1  gate1713(.a(s_167), .O(gate20inter4));
  nand2 gate1714(.a(gate20inter4), .b(gate20inter3), .O(gate20inter5));
  nor2  gate1715(.a(gate20inter5), .b(gate20inter2), .O(gate20inter6));
  inv1  gate1716(.a(G23), .O(gate20inter7));
  inv1  gate1717(.a(G24), .O(gate20inter8));
  nand2 gate1718(.a(gate20inter8), .b(gate20inter7), .O(gate20inter9));
  nand2 gate1719(.a(s_167), .b(gate20inter3), .O(gate20inter10));
  nor2  gate1720(.a(gate20inter10), .b(gate20inter9), .O(gate20inter11));
  nor2  gate1721(.a(gate20inter11), .b(gate20inter6), .O(gate20inter12));
  nand2 gate1722(.a(gate20inter12), .b(gate20inter1), .O(G299));
nand2 gate21( .a(G25), .b(G26), .O(G302) );
nand2 gate22( .a(G27), .b(G28), .O(G305) );

  xor2  gate1485(.a(G30), .b(G29), .O(gate23inter0));
  nand2 gate1486(.a(gate23inter0), .b(s_134), .O(gate23inter1));
  and2  gate1487(.a(G30), .b(G29), .O(gate23inter2));
  inv1  gate1488(.a(s_134), .O(gate23inter3));
  inv1  gate1489(.a(s_135), .O(gate23inter4));
  nand2 gate1490(.a(gate23inter4), .b(gate23inter3), .O(gate23inter5));
  nor2  gate1491(.a(gate23inter5), .b(gate23inter2), .O(gate23inter6));
  inv1  gate1492(.a(G29), .O(gate23inter7));
  inv1  gate1493(.a(G30), .O(gate23inter8));
  nand2 gate1494(.a(gate23inter8), .b(gate23inter7), .O(gate23inter9));
  nand2 gate1495(.a(s_135), .b(gate23inter3), .O(gate23inter10));
  nor2  gate1496(.a(gate23inter10), .b(gate23inter9), .O(gate23inter11));
  nor2  gate1497(.a(gate23inter11), .b(gate23inter6), .O(gate23inter12));
  nand2 gate1498(.a(gate23inter12), .b(gate23inter1), .O(G308));

  xor2  gate3067(.a(G32), .b(G31), .O(gate24inter0));
  nand2 gate3068(.a(gate24inter0), .b(s_360), .O(gate24inter1));
  and2  gate3069(.a(G32), .b(G31), .O(gate24inter2));
  inv1  gate3070(.a(s_360), .O(gate24inter3));
  inv1  gate3071(.a(s_361), .O(gate24inter4));
  nand2 gate3072(.a(gate24inter4), .b(gate24inter3), .O(gate24inter5));
  nor2  gate3073(.a(gate24inter5), .b(gate24inter2), .O(gate24inter6));
  inv1  gate3074(.a(G31), .O(gate24inter7));
  inv1  gate3075(.a(G32), .O(gate24inter8));
  nand2 gate3076(.a(gate24inter8), .b(gate24inter7), .O(gate24inter9));
  nand2 gate3077(.a(s_361), .b(gate24inter3), .O(gate24inter10));
  nor2  gate3078(.a(gate24inter10), .b(gate24inter9), .O(gate24inter11));
  nor2  gate3079(.a(gate24inter11), .b(gate24inter6), .O(gate24inter12));
  nand2 gate3080(.a(gate24inter12), .b(gate24inter1), .O(G311));
nand2 gate25( .a(G1), .b(G5), .O(G314) );
nand2 gate26( .a(G9), .b(G13), .O(G317) );

  xor2  gate2129(.a(G6), .b(G2), .O(gate27inter0));
  nand2 gate2130(.a(gate27inter0), .b(s_226), .O(gate27inter1));
  and2  gate2131(.a(G6), .b(G2), .O(gate27inter2));
  inv1  gate2132(.a(s_226), .O(gate27inter3));
  inv1  gate2133(.a(s_227), .O(gate27inter4));
  nand2 gate2134(.a(gate27inter4), .b(gate27inter3), .O(gate27inter5));
  nor2  gate2135(.a(gate27inter5), .b(gate27inter2), .O(gate27inter6));
  inv1  gate2136(.a(G2), .O(gate27inter7));
  inv1  gate2137(.a(G6), .O(gate27inter8));
  nand2 gate2138(.a(gate27inter8), .b(gate27inter7), .O(gate27inter9));
  nand2 gate2139(.a(s_227), .b(gate27inter3), .O(gate27inter10));
  nor2  gate2140(.a(gate27inter10), .b(gate27inter9), .O(gate27inter11));
  nor2  gate2141(.a(gate27inter11), .b(gate27inter6), .O(gate27inter12));
  nand2 gate2142(.a(gate27inter12), .b(gate27inter1), .O(G320));
nand2 gate28( .a(G10), .b(G14), .O(G323) );
nand2 gate29( .a(G3), .b(G7), .O(G326) );
nand2 gate30( .a(G11), .b(G15), .O(G329) );

  xor2  gate2115(.a(G8), .b(G4), .O(gate31inter0));
  nand2 gate2116(.a(gate31inter0), .b(s_224), .O(gate31inter1));
  and2  gate2117(.a(G8), .b(G4), .O(gate31inter2));
  inv1  gate2118(.a(s_224), .O(gate31inter3));
  inv1  gate2119(.a(s_225), .O(gate31inter4));
  nand2 gate2120(.a(gate31inter4), .b(gate31inter3), .O(gate31inter5));
  nor2  gate2121(.a(gate31inter5), .b(gate31inter2), .O(gate31inter6));
  inv1  gate2122(.a(G4), .O(gate31inter7));
  inv1  gate2123(.a(G8), .O(gate31inter8));
  nand2 gate2124(.a(gate31inter8), .b(gate31inter7), .O(gate31inter9));
  nand2 gate2125(.a(s_225), .b(gate31inter3), .O(gate31inter10));
  nor2  gate2126(.a(gate31inter10), .b(gate31inter9), .O(gate31inter11));
  nor2  gate2127(.a(gate31inter11), .b(gate31inter6), .O(gate31inter12));
  nand2 gate2128(.a(gate31inter12), .b(gate31inter1), .O(G332));
nand2 gate32( .a(G12), .b(G16), .O(G335) );
nand2 gate33( .a(G17), .b(G21), .O(G338) );

  xor2  gate869(.a(G29), .b(G25), .O(gate34inter0));
  nand2 gate870(.a(gate34inter0), .b(s_46), .O(gate34inter1));
  and2  gate871(.a(G29), .b(G25), .O(gate34inter2));
  inv1  gate872(.a(s_46), .O(gate34inter3));
  inv1  gate873(.a(s_47), .O(gate34inter4));
  nand2 gate874(.a(gate34inter4), .b(gate34inter3), .O(gate34inter5));
  nor2  gate875(.a(gate34inter5), .b(gate34inter2), .O(gate34inter6));
  inv1  gate876(.a(G25), .O(gate34inter7));
  inv1  gate877(.a(G29), .O(gate34inter8));
  nand2 gate878(.a(gate34inter8), .b(gate34inter7), .O(gate34inter9));
  nand2 gate879(.a(s_47), .b(gate34inter3), .O(gate34inter10));
  nor2  gate880(.a(gate34inter10), .b(gate34inter9), .O(gate34inter11));
  nor2  gate881(.a(gate34inter11), .b(gate34inter6), .O(gate34inter12));
  nand2 gate882(.a(gate34inter12), .b(gate34inter1), .O(G341));
nand2 gate35( .a(G18), .b(G22), .O(G344) );
nand2 gate36( .a(G26), .b(G30), .O(G347) );

  xor2  gate2577(.a(G23), .b(G19), .O(gate37inter0));
  nand2 gate2578(.a(gate37inter0), .b(s_290), .O(gate37inter1));
  and2  gate2579(.a(G23), .b(G19), .O(gate37inter2));
  inv1  gate2580(.a(s_290), .O(gate37inter3));
  inv1  gate2581(.a(s_291), .O(gate37inter4));
  nand2 gate2582(.a(gate37inter4), .b(gate37inter3), .O(gate37inter5));
  nor2  gate2583(.a(gate37inter5), .b(gate37inter2), .O(gate37inter6));
  inv1  gate2584(.a(G19), .O(gate37inter7));
  inv1  gate2585(.a(G23), .O(gate37inter8));
  nand2 gate2586(.a(gate37inter8), .b(gate37inter7), .O(gate37inter9));
  nand2 gate2587(.a(s_291), .b(gate37inter3), .O(gate37inter10));
  nor2  gate2588(.a(gate37inter10), .b(gate37inter9), .O(gate37inter11));
  nor2  gate2589(.a(gate37inter11), .b(gate37inter6), .O(gate37inter12));
  nand2 gate2590(.a(gate37inter12), .b(gate37inter1), .O(G350));

  xor2  gate2395(.a(G31), .b(G27), .O(gate38inter0));
  nand2 gate2396(.a(gate38inter0), .b(s_264), .O(gate38inter1));
  and2  gate2397(.a(G31), .b(G27), .O(gate38inter2));
  inv1  gate2398(.a(s_264), .O(gate38inter3));
  inv1  gate2399(.a(s_265), .O(gate38inter4));
  nand2 gate2400(.a(gate38inter4), .b(gate38inter3), .O(gate38inter5));
  nor2  gate2401(.a(gate38inter5), .b(gate38inter2), .O(gate38inter6));
  inv1  gate2402(.a(G27), .O(gate38inter7));
  inv1  gate2403(.a(G31), .O(gate38inter8));
  nand2 gate2404(.a(gate38inter8), .b(gate38inter7), .O(gate38inter9));
  nand2 gate2405(.a(s_265), .b(gate38inter3), .O(gate38inter10));
  nor2  gate2406(.a(gate38inter10), .b(gate38inter9), .O(gate38inter11));
  nor2  gate2407(.a(gate38inter11), .b(gate38inter6), .O(gate38inter12));
  nand2 gate2408(.a(gate38inter12), .b(gate38inter1), .O(G353));

  xor2  gate1065(.a(G24), .b(G20), .O(gate39inter0));
  nand2 gate1066(.a(gate39inter0), .b(s_74), .O(gate39inter1));
  and2  gate1067(.a(G24), .b(G20), .O(gate39inter2));
  inv1  gate1068(.a(s_74), .O(gate39inter3));
  inv1  gate1069(.a(s_75), .O(gate39inter4));
  nand2 gate1070(.a(gate39inter4), .b(gate39inter3), .O(gate39inter5));
  nor2  gate1071(.a(gate39inter5), .b(gate39inter2), .O(gate39inter6));
  inv1  gate1072(.a(G20), .O(gate39inter7));
  inv1  gate1073(.a(G24), .O(gate39inter8));
  nand2 gate1074(.a(gate39inter8), .b(gate39inter7), .O(gate39inter9));
  nand2 gate1075(.a(s_75), .b(gate39inter3), .O(gate39inter10));
  nor2  gate1076(.a(gate39inter10), .b(gate39inter9), .O(gate39inter11));
  nor2  gate1077(.a(gate39inter11), .b(gate39inter6), .O(gate39inter12));
  nand2 gate1078(.a(gate39inter12), .b(gate39inter1), .O(G356));

  xor2  gate2017(.a(G32), .b(G28), .O(gate40inter0));
  nand2 gate2018(.a(gate40inter0), .b(s_210), .O(gate40inter1));
  and2  gate2019(.a(G32), .b(G28), .O(gate40inter2));
  inv1  gate2020(.a(s_210), .O(gate40inter3));
  inv1  gate2021(.a(s_211), .O(gate40inter4));
  nand2 gate2022(.a(gate40inter4), .b(gate40inter3), .O(gate40inter5));
  nor2  gate2023(.a(gate40inter5), .b(gate40inter2), .O(gate40inter6));
  inv1  gate2024(.a(G28), .O(gate40inter7));
  inv1  gate2025(.a(G32), .O(gate40inter8));
  nand2 gate2026(.a(gate40inter8), .b(gate40inter7), .O(gate40inter9));
  nand2 gate2027(.a(s_211), .b(gate40inter3), .O(gate40inter10));
  nor2  gate2028(.a(gate40inter10), .b(gate40inter9), .O(gate40inter11));
  nor2  gate2029(.a(gate40inter11), .b(gate40inter6), .O(gate40inter12));
  nand2 gate2030(.a(gate40inter12), .b(gate40inter1), .O(G359));

  xor2  gate841(.a(G266), .b(G1), .O(gate41inter0));
  nand2 gate842(.a(gate41inter0), .b(s_42), .O(gate41inter1));
  and2  gate843(.a(G266), .b(G1), .O(gate41inter2));
  inv1  gate844(.a(s_42), .O(gate41inter3));
  inv1  gate845(.a(s_43), .O(gate41inter4));
  nand2 gate846(.a(gate41inter4), .b(gate41inter3), .O(gate41inter5));
  nor2  gate847(.a(gate41inter5), .b(gate41inter2), .O(gate41inter6));
  inv1  gate848(.a(G1), .O(gate41inter7));
  inv1  gate849(.a(G266), .O(gate41inter8));
  nand2 gate850(.a(gate41inter8), .b(gate41inter7), .O(gate41inter9));
  nand2 gate851(.a(s_43), .b(gate41inter3), .O(gate41inter10));
  nor2  gate852(.a(gate41inter10), .b(gate41inter9), .O(gate41inter11));
  nor2  gate853(.a(gate41inter11), .b(gate41inter6), .O(gate41inter12));
  nand2 gate854(.a(gate41inter12), .b(gate41inter1), .O(G362));
nand2 gate42( .a(G2), .b(G266), .O(G363) );
nand2 gate43( .a(G3), .b(G269), .O(G364) );
nand2 gate44( .a(G4), .b(G269), .O(G365) );
nand2 gate45( .a(G5), .b(G272), .O(G366) );
nand2 gate46( .a(G6), .b(G272), .O(G367) );

  xor2  gate2507(.a(G275), .b(G7), .O(gate47inter0));
  nand2 gate2508(.a(gate47inter0), .b(s_280), .O(gate47inter1));
  and2  gate2509(.a(G275), .b(G7), .O(gate47inter2));
  inv1  gate2510(.a(s_280), .O(gate47inter3));
  inv1  gate2511(.a(s_281), .O(gate47inter4));
  nand2 gate2512(.a(gate47inter4), .b(gate47inter3), .O(gate47inter5));
  nor2  gate2513(.a(gate47inter5), .b(gate47inter2), .O(gate47inter6));
  inv1  gate2514(.a(G7), .O(gate47inter7));
  inv1  gate2515(.a(G275), .O(gate47inter8));
  nand2 gate2516(.a(gate47inter8), .b(gate47inter7), .O(gate47inter9));
  nand2 gate2517(.a(s_281), .b(gate47inter3), .O(gate47inter10));
  nor2  gate2518(.a(gate47inter10), .b(gate47inter9), .O(gate47inter11));
  nor2  gate2519(.a(gate47inter11), .b(gate47inter6), .O(gate47inter12));
  nand2 gate2520(.a(gate47inter12), .b(gate47inter1), .O(G368));
nand2 gate48( .a(G8), .b(G275), .O(G369) );

  xor2  gate1751(.a(G278), .b(G9), .O(gate49inter0));
  nand2 gate1752(.a(gate49inter0), .b(s_172), .O(gate49inter1));
  and2  gate1753(.a(G278), .b(G9), .O(gate49inter2));
  inv1  gate1754(.a(s_172), .O(gate49inter3));
  inv1  gate1755(.a(s_173), .O(gate49inter4));
  nand2 gate1756(.a(gate49inter4), .b(gate49inter3), .O(gate49inter5));
  nor2  gate1757(.a(gate49inter5), .b(gate49inter2), .O(gate49inter6));
  inv1  gate1758(.a(G9), .O(gate49inter7));
  inv1  gate1759(.a(G278), .O(gate49inter8));
  nand2 gate1760(.a(gate49inter8), .b(gate49inter7), .O(gate49inter9));
  nand2 gate1761(.a(s_173), .b(gate49inter3), .O(gate49inter10));
  nor2  gate1762(.a(gate49inter10), .b(gate49inter9), .O(gate49inter11));
  nor2  gate1763(.a(gate49inter11), .b(gate49inter6), .O(gate49inter12));
  nand2 gate1764(.a(gate49inter12), .b(gate49inter1), .O(G370));
nand2 gate50( .a(G10), .b(G278), .O(G371) );
nand2 gate51( .a(G11), .b(G281), .O(G372) );
nand2 gate52( .a(G12), .b(G281), .O(G373) );
nand2 gate53( .a(G13), .b(G284), .O(G374) );
nand2 gate54( .a(G14), .b(G284), .O(G375) );
nand2 gate55( .a(G15), .b(G287), .O(G376) );
nand2 gate56( .a(G16), .b(G287), .O(G377) );
nand2 gate57( .a(G17), .b(G290), .O(G378) );
nand2 gate58( .a(G18), .b(G290), .O(G379) );
nand2 gate59( .a(G19), .b(G293), .O(G380) );
nand2 gate60( .a(G20), .b(G293), .O(G381) );
nand2 gate61( .a(G21), .b(G296), .O(G382) );

  xor2  gate2241(.a(G296), .b(G22), .O(gate62inter0));
  nand2 gate2242(.a(gate62inter0), .b(s_242), .O(gate62inter1));
  and2  gate2243(.a(G296), .b(G22), .O(gate62inter2));
  inv1  gate2244(.a(s_242), .O(gate62inter3));
  inv1  gate2245(.a(s_243), .O(gate62inter4));
  nand2 gate2246(.a(gate62inter4), .b(gate62inter3), .O(gate62inter5));
  nor2  gate2247(.a(gate62inter5), .b(gate62inter2), .O(gate62inter6));
  inv1  gate2248(.a(G22), .O(gate62inter7));
  inv1  gate2249(.a(G296), .O(gate62inter8));
  nand2 gate2250(.a(gate62inter8), .b(gate62inter7), .O(gate62inter9));
  nand2 gate2251(.a(s_243), .b(gate62inter3), .O(gate62inter10));
  nor2  gate2252(.a(gate62inter10), .b(gate62inter9), .O(gate62inter11));
  nor2  gate2253(.a(gate62inter11), .b(gate62inter6), .O(gate62inter12));
  nand2 gate2254(.a(gate62inter12), .b(gate62inter1), .O(G383));
nand2 gate63( .a(G23), .b(G299), .O(G384) );

  xor2  gate785(.a(G299), .b(G24), .O(gate64inter0));
  nand2 gate786(.a(gate64inter0), .b(s_34), .O(gate64inter1));
  and2  gate787(.a(G299), .b(G24), .O(gate64inter2));
  inv1  gate788(.a(s_34), .O(gate64inter3));
  inv1  gate789(.a(s_35), .O(gate64inter4));
  nand2 gate790(.a(gate64inter4), .b(gate64inter3), .O(gate64inter5));
  nor2  gate791(.a(gate64inter5), .b(gate64inter2), .O(gate64inter6));
  inv1  gate792(.a(G24), .O(gate64inter7));
  inv1  gate793(.a(G299), .O(gate64inter8));
  nand2 gate794(.a(gate64inter8), .b(gate64inter7), .O(gate64inter9));
  nand2 gate795(.a(s_35), .b(gate64inter3), .O(gate64inter10));
  nor2  gate796(.a(gate64inter10), .b(gate64inter9), .O(gate64inter11));
  nor2  gate797(.a(gate64inter11), .b(gate64inter6), .O(gate64inter12));
  nand2 gate798(.a(gate64inter12), .b(gate64inter1), .O(G385));
nand2 gate65( .a(G25), .b(G302), .O(G386) );

  xor2  gate631(.a(G302), .b(G26), .O(gate66inter0));
  nand2 gate632(.a(gate66inter0), .b(s_12), .O(gate66inter1));
  and2  gate633(.a(G302), .b(G26), .O(gate66inter2));
  inv1  gate634(.a(s_12), .O(gate66inter3));
  inv1  gate635(.a(s_13), .O(gate66inter4));
  nand2 gate636(.a(gate66inter4), .b(gate66inter3), .O(gate66inter5));
  nor2  gate637(.a(gate66inter5), .b(gate66inter2), .O(gate66inter6));
  inv1  gate638(.a(G26), .O(gate66inter7));
  inv1  gate639(.a(G302), .O(gate66inter8));
  nand2 gate640(.a(gate66inter8), .b(gate66inter7), .O(gate66inter9));
  nand2 gate641(.a(s_13), .b(gate66inter3), .O(gate66inter10));
  nor2  gate642(.a(gate66inter10), .b(gate66inter9), .O(gate66inter11));
  nor2  gate643(.a(gate66inter11), .b(gate66inter6), .O(gate66inter12));
  nand2 gate644(.a(gate66inter12), .b(gate66inter1), .O(G387));
nand2 gate67( .a(G27), .b(G305), .O(G388) );

  xor2  gate1611(.a(G305), .b(G28), .O(gate68inter0));
  nand2 gate1612(.a(gate68inter0), .b(s_152), .O(gate68inter1));
  and2  gate1613(.a(G305), .b(G28), .O(gate68inter2));
  inv1  gate1614(.a(s_152), .O(gate68inter3));
  inv1  gate1615(.a(s_153), .O(gate68inter4));
  nand2 gate1616(.a(gate68inter4), .b(gate68inter3), .O(gate68inter5));
  nor2  gate1617(.a(gate68inter5), .b(gate68inter2), .O(gate68inter6));
  inv1  gate1618(.a(G28), .O(gate68inter7));
  inv1  gate1619(.a(G305), .O(gate68inter8));
  nand2 gate1620(.a(gate68inter8), .b(gate68inter7), .O(gate68inter9));
  nand2 gate1621(.a(s_153), .b(gate68inter3), .O(gate68inter10));
  nor2  gate1622(.a(gate68inter10), .b(gate68inter9), .O(gate68inter11));
  nor2  gate1623(.a(gate68inter11), .b(gate68inter6), .O(gate68inter12));
  nand2 gate1624(.a(gate68inter12), .b(gate68inter1), .O(G389));

  xor2  gate2983(.a(G308), .b(G29), .O(gate69inter0));
  nand2 gate2984(.a(gate69inter0), .b(s_348), .O(gate69inter1));
  and2  gate2985(.a(G308), .b(G29), .O(gate69inter2));
  inv1  gate2986(.a(s_348), .O(gate69inter3));
  inv1  gate2987(.a(s_349), .O(gate69inter4));
  nand2 gate2988(.a(gate69inter4), .b(gate69inter3), .O(gate69inter5));
  nor2  gate2989(.a(gate69inter5), .b(gate69inter2), .O(gate69inter6));
  inv1  gate2990(.a(G29), .O(gate69inter7));
  inv1  gate2991(.a(G308), .O(gate69inter8));
  nand2 gate2992(.a(gate69inter8), .b(gate69inter7), .O(gate69inter9));
  nand2 gate2993(.a(s_349), .b(gate69inter3), .O(gate69inter10));
  nor2  gate2994(.a(gate69inter10), .b(gate69inter9), .O(gate69inter11));
  nor2  gate2995(.a(gate69inter11), .b(gate69inter6), .O(gate69inter12));
  nand2 gate2996(.a(gate69inter12), .b(gate69inter1), .O(G390));

  xor2  gate1919(.a(G308), .b(G30), .O(gate70inter0));
  nand2 gate1920(.a(gate70inter0), .b(s_196), .O(gate70inter1));
  and2  gate1921(.a(G308), .b(G30), .O(gate70inter2));
  inv1  gate1922(.a(s_196), .O(gate70inter3));
  inv1  gate1923(.a(s_197), .O(gate70inter4));
  nand2 gate1924(.a(gate70inter4), .b(gate70inter3), .O(gate70inter5));
  nor2  gate1925(.a(gate70inter5), .b(gate70inter2), .O(gate70inter6));
  inv1  gate1926(.a(G30), .O(gate70inter7));
  inv1  gate1927(.a(G308), .O(gate70inter8));
  nand2 gate1928(.a(gate70inter8), .b(gate70inter7), .O(gate70inter9));
  nand2 gate1929(.a(s_197), .b(gate70inter3), .O(gate70inter10));
  nor2  gate1930(.a(gate70inter10), .b(gate70inter9), .O(gate70inter11));
  nor2  gate1931(.a(gate70inter11), .b(gate70inter6), .O(gate70inter12));
  nand2 gate1932(.a(gate70inter12), .b(gate70inter1), .O(G391));
nand2 gate71( .a(G31), .b(G311), .O(G392) );
nand2 gate72( .a(G32), .b(G311), .O(G393) );
nand2 gate73( .a(G1), .b(G314), .O(G394) );
nand2 gate74( .a(G5), .b(G314), .O(G395) );
nand2 gate75( .a(G9), .b(G317), .O(G396) );

  xor2  gate1765(.a(G317), .b(G13), .O(gate76inter0));
  nand2 gate1766(.a(gate76inter0), .b(s_174), .O(gate76inter1));
  and2  gate1767(.a(G317), .b(G13), .O(gate76inter2));
  inv1  gate1768(.a(s_174), .O(gate76inter3));
  inv1  gate1769(.a(s_175), .O(gate76inter4));
  nand2 gate1770(.a(gate76inter4), .b(gate76inter3), .O(gate76inter5));
  nor2  gate1771(.a(gate76inter5), .b(gate76inter2), .O(gate76inter6));
  inv1  gate1772(.a(G13), .O(gate76inter7));
  inv1  gate1773(.a(G317), .O(gate76inter8));
  nand2 gate1774(.a(gate76inter8), .b(gate76inter7), .O(gate76inter9));
  nand2 gate1775(.a(s_175), .b(gate76inter3), .O(gate76inter10));
  nor2  gate1776(.a(gate76inter10), .b(gate76inter9), .O(gate76inter11));
  nor2  gate1777(.a(gate76inter11), .b(gate76inter6), .O(gate76inter12));
  nand2 gate1778(.a(gate76inter12), .b(gate76inter1), .O(G397));
nand2 gate77( .a(G2), .b(G320), .O(G398) );
nand2 gate78( .a(G6), .b(G320), .O(G399) );

  xor2  gate3095(.a(G323), .b(G10), .O(gate79inter0));
  nand2 gate3096(.a(gate79inter0), .b(s_364), .O(gate79inter1));
  and2  gate3097(.a(G323), .b(G10), .O(gate79inter2));
  inv1  gate3098(.a(s_364), .O(gate79inter3));
  inv1  gate3099(.a(s_365), .O(gate79inter4));
  nand2 gate3100(.a(gate79inter4), .b(gate79inter3), .O(gate79inter5));
  nor2  gate3101(.a(gate79inter5), .b(gate79inter2), .O(gate79inter6));
  inv1  gate3102(.a(G10), .O(gate79inter7));
  inv1  gate3103(.a(G323), .O(gate79inter8));
  nand2 gate3104(.a(gate79inter8), .b(gate79inter7), .O(gate79inter9));
  nand2 gate3105(.a(s_365), .b(gate79inter3), .O(gate79inter10));
  nor2  gate3106(.a(gate79inter10), .b(gate79inter9), .O(gate79inter11));
  nor2  gate3107(.a(gate79inter11), .b(gate79inter6), .O(gate79inter12));
  nand2 gate3108(.a(gate79inter12), .b(gate79inter1), .O(G400));
nand2 gate80( .a(G14), .b(G323), .O(G401) );
nand2 gate81( .a(G3), .b(G326), .O(G402) );

  xor2  gate715(.a(G326), .b(G7), .O(gate82inter0));
  nand2 gate716(.a(gate82inter0), .b(s_24), .O(gate82inter1));
  and2  gate717(.a(G326), .b(G7), .O(gate82inter2));
  inv1  gate718(.a(s_24), .O(gate82inter3));
  inv1  gate719(.a(s_25), .O(gate82inter4));
  nand2 gate720(.a(gate82inter4), .b(gate82inter3), .O(gate82inter5));
  nor2  gate721(.a(gate82inter5), .b(gate82inter2), .O(gate82inter6));
  inv1  gate722(.a(G7), .O(gate82inter7));
  inv1  gate723(.a(G326), .O(gate82inter8));
  nand2 gate724(.a(gate82inter8), .b(gate82inter7), .O(gate82inter9));
  nand2 gate725(.a(s_25), .b(gate82inter3), .O(gate82inter10));
  nor2  gate726(.a(gate82inter10), .b(gate82inter9), .O(gate82inter11));
  nor2  gate727(.a(gate82inter11), .b(gate82inter6), .O(gate82inter12));
  nand2 gate728(.a(gate82inter12), .b(gate82inter1), .O(G403));

  xor2  gate3165(.a(G329), .b(G11), .O(gate83inter0));
  nand2 gate3166(.a(gate83inter0), .b(s_374), .O(gate83inter1));
  and2  gate3167(.a(G329), .b(G11), .O(gate83inter2));
  inv1  gate3168(.a(s_374), .O(gate83inter3));
  inv1  gate3169(.a(s_375), .O(gate83inter4));
  nand2 gate3170(.a(gate83inter4), .b(gate83inter3), .O(gate83inter5));
  nor2  gate3171(.a(gate83inter5), .b(gate83inter2), .O(gate83inter6));
  inv1  gate3172(.a(G11), .O(gate83inter7));
  inv1  gate3173(.a(G329), .O(gate83inter8));
  nand2 gate3174(.a(gate83inter8), .b(gate83inter7), .O(gate83inter9));
  nand2 gate3175(.a(s_375), .b(gate83inter3), .O(gate83inter10));
  nor2  gate3176(.a(gate83inter10), .b(gate83inter9), .O(gate83inter11));
  nor2  gate3177(.a(gate83inter11), .b(gate83inter6), .O(gate83inter12));
  nand2 gate3178(.a(gate83inter12), .b(gate83inter1), .O(G404));

  xor2  gate2969(.a(G329), .b(G15), .O(gate84inter0));
  nand2 gate2970(.a(gate84inter0), .b(s_346), .O(gate84inter1));
  and2  gate2971(.a(G329), .b(G15), .O(gate84inter2));
  inv1  gate2972(.a(s_346), .O(gate84inter3));
  inv1  gate2973(.a(s_347), .O(gate84inter4));
  nand2 gate2974(.a(gate84inter4), .b(gate84inter3), .O(gate84inter5));
  nor2  gate2975(.a(gate84inter5), .b(gate84inter2), .O(gate84inter6));
  inv1  gate2976(.a(G15), .O(gate84inter7));
  inv1  gate2977(.a(G329), .O(gate84inter8));
  nand2 gate2978(.a(gate84inter8), .b(gate84inter7), .O(gate84inter9));
  nand2 gate2979(.a(s_347), .b(gate84inter3), .O(gate84inter10));
  nor2  gate2980(.a(gate84inter10), .b(gate84inter9), .O(gate84inter11));
  nor2  gate2981(.a(gate84inter11), .b(gate84inter6), .O(gate84inter12));
  nand2 gate2982(.a(gate84inter12), .b(gate84inter1), .O(G405));

  xor2  gate1149(.a(G332), .b(G4), .O(gate85inter0));
  nand2 gate1150(.a(gate85inter0), .b(s_86), .O(gate85inter1));
  and2  gate1151(.a(G332), .b(G4), .O(gate85inter2));
  inv1  gate1152(.a(s_86), .O(gate85inter3));
  inv1  gate1153(.a(s_87), .O(gate85inter4));
  nand2 gate1154(.a(gate85inter4), .b(gate85inter3), .O(gate85inter5));
  nor2  gate1155(.a(gate85inter5), .b(gate85inter2), .O(gate85inter6));
  inv1  gate1156(.a(G4), .O(gate85inter7));
  inv1  gate1157(.a(G332), .O(gate85inter8));
  nand2 gate1158(.a(gate85inter8), .b(gate85inter7), .O(gate85inter9));
  nand2 gate1159(.a(s_87), .b(gate85inter3), .O(gate85inter10));
  nor2  gate1160(.a(gate85inter10), .b(gate85inter9), .O(gate85inter11));
  nor2  gate1161(.a(gate85inter11), .b(gate85inter6), .O(gate85inter12));
  nand2 gate1162(.a(gate85inter12), .b(gate85inter1), .O(G406));

  xor2  gate3039(.a(G332), .b(G8), .O(gate86inter0));
  nand2 gate3040(.a(gate86inter0), .b(s_356), .O(gate86inter1));
  and2  gate3041(.a(G332), .b(G8), .O(gate86inter2));
  inv1  gate3042(.a(s_356), .O(gate86inter3));
  inv1  gate3043(.a(s_357), .O(gate86inter4));
  nand2 gate3044(.a(gate86inter4), .b(gate86inter3), .O(gate86inter5));
  nor2  gate3045(.a(gate86inter5), .b(gate86inter2), .O(gate86inter6));
  inv1  gate3046(.a(G8), .O(gate86inter7));
  inv1  gate3047(.a(G332), .O(gate86inter8));
  nand2 gate3048(.a(gate86inter8), .b(gate86inter7), .O(gate86inter9));
  nand2 gate3049(.a(s_357), .b(gate86inter3), .O(gate86inter10));
  nor2  gate3050(.a(gate86inter10), .b(gate86inter9), .O(gate86inter11));
  nor2  gate3051(.a(gate86inter11), .b(gate86inter6), .O(gate86inter12));
  nand2 gate3052(.a(gate86inter12), .b(gate86inter1), .O(G407));
nand2 gate87( .a(G12), .b(G335), .O(G408) );

  xor2  gate2619(.a(G335), .b(G16), .O(gate88inter0));
  nand2 gate2620(.a(gate88inter0), .b(s_296), .O(gate88inter1));
  and2  gate2621(.a(G335), .b(G16), .O(gate88inter2));
  inv1  gate2622(.a(s_296), .O(gate88inter3));
  inv1  gate2623(.a(s_297), .O(gate88inter4));
  nand2 gate2624(.a(gate88inter4), .b(gate88inter3), .O(gate88inter5));
  nor2  gate2625(.a(gate88inter5), .b(gate88inter2), .O(gate88inter6));
  inv1  gate2626(.a(G16), .O(gate88inter7));
  inv1  gate2627(.a(G335), .O(gate88inter8));
  nand2 gate2628(.a(gate88inter8), .b(gate88inter7), .O(gate88inter9));
  nand2 gate2629(.a(s_297), .b(gate88inter3), .O(gate88inter10));
  nor2  gate2630(.a(gate88inter10), .b(gate88inter9), .O(gate88inter11));
  nor2  gate2631(.a(gate88inter11), .b(gate88inter6), .O(gate88inter12));
  nand2 gate2632(.a(gate88inter12), .b(gate88inter1), .O(G409));

  xor2  gate1961(.a(G338), .b(G17), .O(gate89inter0));
  nand2 gate1962(.a(gate89inter0), .b(s_202), .O(gate89inter1));
  and2  gate1963(.a(G338), .b(G17), .O(gate89inter2));
  inv1  gate1964(.a(s_202), .O(gate89inter3));
  inv1  gate1965(.a(s_203), .O(gate89inter4));
  nand2 gate1966(.a(gate89inter4), .b(gate89inter3), .O(gate89inter5));
  nor2  gate1967(.a(gate89inter5), .b(gate89inter2), .O(gate89inter6));
  inv1  gate1968(.a(G17), .O(gate89inter7));
  inv1  gate1969(.a(G338), .O(gate89inter8));
  nand2 gate1970(.a(gate89inter8), .b(gate89inter7), .O(gate89inter9));
  nand2 gate1971(.a(s_203), .b(gate89inter3), .O(gate89inter10));
  nor2  gate1972(.a(gate89inter10), .b(gate89inter9), .O(gate89inter11));
  nor2  gate1973(.a(gate89inter11), .b(gate89inter6), .O(gate89inter12));
  nand2 gate1974(.a(gate89inter12), .b(gate89inter1), .O(G410));

  xor2  gate1737(.a(G338), .b(G21), .O(gate90inter0));
  nand2 gate1738(.a(gate90inter0), .b(s_170), .O(gate90inter1));
  and2  gate1739(.a(G338), .b(G21), .O(gate90inter2));
  inv1  gate1740(.a(s_170), .O(gate90inter3));
  inv1  gate1741(.a(s_171), .O(gate90inter4));
  nand2 gate1742(.a(gate90inter4), .b(gate90inter3), .O(gate90inter5));
  nor2  gate1743(.a(gate90inter5), .b(gate90inter2), .O(gate90inter6));
  inv1  gate1744(.a(G21), .O(gate90inter7));
  inv1  gate1745(.a(G338), .O(gate90inter8));
  nand2 gate1746(.a(gate90inter8), .b(gate90inter7), .O(gate90inter9));
  nand2 gate1747(.a(s_171), .b(gate90inter3), .O(gate90inter10));
  nor2  gate1748(.a(gate90inter10), .b(gate90inter9), .O(gate90inter11));
  nor2  gate1749(.a(gate90inter11), .b(gate90inter6), .O(gate90inter12));
  nand2 gate1750(.a(gate90inter12), .b(gate90inter1), .O(G411));
nand2 gate91( .a(G25), .b(G341), .O(G412) );
nand2 gate92( .a(G29), .b(G341), .O(G413) );
nand2 gate93( .a(G18), .b(G344), .O(G414) );

  xor2  gate673(.a(G344), .b(G22), .O(gate94inter0));
  nand2 gate674(.a(gate94inter0), .b(s_18), .O(gate94inter1));
  and2  gate675(.a(G344), .b(G22), .O(gate94inter2));
  inv1  gate676(.a(s_18), .O(gate94inter3));
  inv1  gate677(.a(s_19), .O(gate94inter4));
  nand2 gate678(.a(gate94inter4), .b(gate94inter3), .O(gate94inter5));
  nor2  gate679(.a(gate94inter5), .b(gate94inter2), .O(gate94inter6));
  inv1  gate680(.a(G22), .O(gate94inter7));
  inv1  gate681(.a(G344), .O(gate94inter8));
  nand2 gate682(.a(gate94inter8), .b(gate94inter7), .O(gate94inter9));
  nand2 gate683(.a(s_19), .b(gate94inter3), .O(gate94inter10));
  nor2  gate684(.a(gate94inter10), .b(gate94inter9), .O(gate94inter11));
  nor2  gate685(.a(gate94inter11), .b(gate94inter6), .O(gate94inter12));
  nand2 gate686(.a(gate94inter12), .b(gate94inter1), .O(G415));
nand2 gate95( .a(G26), .b(G347), .O(G416) );

  xor2  gate2927(.a(G347), .b(G30), .O(gate96inter0));
  nand2 gate2928(.a(gate96inter0), .b(s_340), .O(gate96inter1));
  and2  gate2929(.a(G347), .b(G30), .O(gate96inter2));
  inv1  gate2930(.a(s_340), .O(gate96inter3));
  inv1  gate2931(.a(s_341), .O(gate96inter4));
  nand2 gate2932(.a(gate96inter4), .b(gate96inter3), .O(gate96inter5));
  nor2  gate2933(.a(gate96inter5), .b(gate96inter2), .O(gate96inter6));
  inv1  gate2934(.a(G30), .O(gate96inter7));
  inv1  gate2935(.a(G347), .O(gate96inter8));
  nand2 gate2936(.a(gate96inter8), .b(gate96inter7), .O(gate96inter9));
  nand2 gate2937(.a(s_341), .b(gate96inter3), .O(gate96inter10));
  nor2  gate2938(.a(gate96inter10), .b(gate96inter9), .O(gate96inter11));
  nor2  gate2939(.a(gate96inter11), .b(gate96inter6), .O(gate96inter12));
  nand2 gate2940(.a(gate96inter12), .b(gate96inter1), .O(G417));
nand2 gate97( .a(G19), .b(G350), .O(G418) );

  xor2  gate1135(.a(G350), .b(G23), .O(gate98inter0));
  nand2 gate1136(.a(gate98inter0), .b(s_84), .O(gate98inter1));
  and2  gate1137(.a(G350), .b(G23), .O(gate98inter2));
  inv1  gate1138(.a(s_84), .O(gate98inter3));
  inv1  gate1139(.a(s_85), .O(gate98inter4));
  nand2 gate1140(.a(gate98inter4), .b(gate98inter3), .O(gate98inter5));
  nor2  gate1141(.a(gate98inter5), .b(gate98inter2), .O(gate98inter6));
  inv1  gate1142(.a(G23), .O(gate98inter7));
  inv1  gate1143(.a(G350), .O(gate98inter8));
  nand2 gate1144(.a(gate98inter8), .b(gate98inter7), .O(gate98inter9));
  nand2 gate1145(.a(s_85), .b(gate98inter3), .O(gate98inter10));
  nor2  gate1146(.a(gate98inter10), .b(gate98inter9), .O(gate98inter11));
  nor2  gate1147(.a(gate98inter11), .b(gate98inter6), .O(gate98inter12));
  nand2 gate1148(.a(gate98inter12), .b(gate98inter1), .O(G419));

  xor2  gate2353(.a(G353), .b(G27), .O(gate99inter0));
  nand2 gate2354(.a(gate99inter0), .b(s_258), .O(gate99inter1));
  and2  gate2355(.a(G353), .b(G27), .O(gate99inter2));
  inv1  gate2356(.a(s_258), .O(gate99inter3));
  inv1  gate2357(.a(s_259), .O(gate99inter4));
  nand2 gate2358(.a(gate99inter4), .b(gate99inter3), .O(gate99inter5));
  nor2  gate2359(.a(gate99inter5), .b(gate99inter2), .O(gate99inter6));
  inv1  gate2360(.a(G27), .O(gate99inter7));
  inv1  gate2361(.a(G353), .O(gate99inter8));
  nand2 gate2362(.a(gate99inter8), .b(gate99inter7), .O(gate99inter9));
  nand2 gate2363(.a(s_259), .b(gate99inter3), .O(gate99inter10));
  nor2  gate2364(.a(gate99inter10), .b(gate99inter9), .O(gate99inter11));
  nor2  gate2365(.a(gate99inter11), .b(gate99inter6), .O(gate99inter12));
  nand2 gate2366(.a(gate99inter12), .b(gate99inter1), .O(G420));
nand2 gate100( .a(G31), .b(G353), .O(G421) );

  xor2  gate2913(.a(G356), .b(G20), .O(gate101inter0));
  nand2 gate2914(.a(gate101inter0), .b(s_338), .O(gate101inter1));
  and2  gate2915(.a(G356), .b(G20), .O(gate101inter2));
  inv1  gate2916(.a(s_338), .O(gate101inter3));
  inv1  gate2917(.a(s_339), .O(gate101inter4));
  nand2 gate2918(.a(gate101inter4), .b(gate101inter3), .O(gate101inter5));
  nor2  gate2919(.a(gate101inter5), .b(gate101inter2), .O(gate101inter6));
  inv1  gate2920(.a(G20), .O(gate101inter7));
  inv1  gate2921(.a(G356), .O(gate101inter8));
  nand2 gate2922(.a(gate101inter8), .b(gate101inter7), .O(gate101inter9));
  nand2 gate2923(.a(s_339), .b(gate101inter3), .O(gate101inter10));
  nor2  gate2924(.a(gate101inter10), .b(gate101inter9), .O(gate101inter11));
  nor2  gate2925(.a(gate101inter11), .b(gate101inter6), .O(gate101inter12));
  nand2 gate2926(.a(gate101inter12), .b(gate101inter1), .O(G422));

  xor2  gate2045(.a(G356), .b(G24), .O(gate102inter0));
  nand2 gate2046(.a(gate102inter0), .b(s_214), .O(gate102inter1));
  and2  gate2047(.a(G356), .b(G24), .O(gate102inter2));
  inv1  gate2048(.a(s_214), .O(gate102inter3));
  inv1  gate2049(.a(s_215), .O(gate102inter4));
  nand2 gate2050(.a(gate102inter4), .b(gate102inter3), .O(gate102inter5));
  nor2  gate2051(.a(gate102inter5), .b(gate102inter2), .O(gate102inter6));
  inv1  gate2052(.a(G24), .O(gate102inter7));
  inv1  gate2053(.a(G356), .O(gate102inter8));
  nand2 gate2054(.a(gate102inter8), .b(gate102inter7), .O(gate102inter9));
  nand2 gate2055(.a(s_215), .b(gate102inter3), .O(gate102inter10));
  nor2  gate2056(.a(gate102inter10), .b(gate102inter9), .O(gate102inter11));
  nor2  gate2057(.a(gate102inter11), .b(gate102inter6), .O(gate102inter12));
  nand2 gate2058(.a(gate102inter12), .b(gate102inter1), .O(G423));

  xor2  gate2199(.a(G359), .b(G28), .O(gate103inter0));
  nand2 gate2200(.a(gate103inter0), .b(s_236), .O(gate103inter1));
  and2  gate2201(.a(G359), .b(G28), .O(gate103inter2));
  inv1  gate2202(.a(s_236), .O(gate103inter3));
  inv1  gate2203(.a(s_237), .O(gate103inter4));
  nand2 gate2204(.a(gate103inter4), .b(gate103inter3), .O(gate103inter5));
  nor2  gate2205(.a(gate103inter5), .b(gate103inter2), .O(gate103inter6));
  inv1  gate2206(.a(G28), .O(gate103inter7));
  inv1  gate2207(.a(G359), .O(gate103inter8));
  nand2 gate2208(.a(gate103inter8), .b(gate103inter7), .O(gate103inter9));
  nand2 gate2209(.a(s_237), .b(gate103inter3), .O(gate103inter10));
  nor2  gate2210(.a(gate103inter10), .b(gate103inter9), .O(gate103inter11));
  nor2  gate2211(.a(gate103inter11), .b(gate103inter6), .O(gate103inter12));
  nand2 gate2212(.a(gate103inter12), .b(gate103inter1), .O(G424));

  xor2  gate2297(.a(G359), .b(G32), .O(gate104inter0));
  nand2 gate2298(.a(gate104inter0), .b(s_250), .O(gate104inter1));
  and2  gate2299(.a(G359), .b(G32), .O(gate104inter2));
  inv1  gate2300(.a(s_250), .O(gate104inter3));
  inv1  gate2301(.a(s_251), .O(gate104inter4));
  nand2 gate2302(.a(gate104inter4), .b(gate104inter3), .O(gate104inter5));
  nor2  gate2303(.a(gate104inter5), .b(gate104inter2), .O(gate104inter6));
  inv1  gate2304(.a(G32), .O(gate104inter7));
  inv1  gate2305(.a(G359), .O(gate104inter8));
  nand2 gate2306(.a(gate104inter8), .b(gate104inter7), .O(gate104inter9));
  nand2 gate2307(.a(s_251), .b(gate104inter3), .O(gate104inter10));
  nor2  gate2308(.a(gate104inter10), .b(gate104inter9), .O(gate104inter11));
  nor2  gate2309(.a(gate104inter11), .b(gate104inter6), .O(gate104inter12));
  nand2 gate2310(.a(gate104inter12), .b(gate104inter1), .O(G425));
nand2 gate105( .a(G362), .b(G363), .O(G426) );
nand2 gate106( .a(G364), .b(G365), .O(G429) );

  xor2  gate1541(.a(G367), .b(G366), .O(gate107inter0));
  nand2 gate1542(.a(gate107inter0), .b(s_142), .O(gate107inter1));
  and2  gate1543(.a(G367), .b(G366), .O(gate107inter2));
  inv1  gate1544(.a(s_142), .O(gate107inter3));
  inv1  gate1545(.a(s_143), .O(gate107inter4));
  nand2 gate1546(.a(gate107inter4), .b(gate107inter3), .O(gate107inter5));
  nor2  gate1547(.a(gate107inter5), .b(gate107inter2), .O(gate107inter6));
  inv1  gate1548(.a(G366), .O(gate107inter7));
  inv1  gate1549(.a(G367), .O(gate107inter8));
  nand2 gate1550(.a(gate107inter8), .b(gate107inter7), .O(gate107inter9));
  nand2 gate1551(.a(s_143), .b(gate107inter3), .O(gate107inter10));
  nor2  gate1552(.a(gate107inter10), .b(gate107inter9), .O(gate107inter11));
  nor2  gate1553(.a(gate107inter11), .b(gate107inter6), .O(gate107inter12));
  nand2 gate1554(.a(gate107inter12), .b(gate107inter1), .O(G432));
nand2 gate108( .a(G368), .b(G369), .O(G435) );
nand2 gate109( .a(G370), .b(G371), .O(G438) );

  xor2  gate1947(.a(G373), .b(G372), .O(gate110inter0));
  nand2 gate1948(.a(gate110inter0), .b(s_200), .O(gate110inter1));
  and2  gate1949(.a(G373), .b(G372), .O(gate110inter2));
  inv1  gate1950(.a(s_200), .O(gate110inter3));
  inv1  gate1951(.a(s_201), .O(gate110inter4));
  nand2 gate1952(.a(gate110inter4), .b(gate110inter3), .O(gate110inter5));
  nor2  gate1953(.a(gate110inter5), .b(gate110inter2), .O(gate110inter6));
  inv1  gate1954(.a(G372), .O(gate110inter7));
  inv1  gate1955(.a(G373), .O(gate110inter8));
  nand2 gate1956(.a(gate110inter8), .b(gate110inter7), .O(gate110inter9));
  nand2 gate1957(.a(s_201), .b(gate110inter3), .O(gate110inter10));
  nor2  gate1958(.a(gate110inter10), .b(gate110inter9), .O(gate110inter11));
  nor2  gate1959(.a(gate110inter11), .b(gate110inter6), .O(gate110inter12));
  nand2 gate1960(.a(gate110inter12), .b(gate110inter1), .O(G441));

  xor2  gate2787(.a(G375), .b(G374), .O(gate111inter0));
  nand2 gate2788(.a(gate111inter0), .b(s_320), .O(gate111inter1));
  and2  gate2789(.a(G375), .b(G374), .O(gate111inter2));
  inv1  gate2790(.a(s_320), .O(gate111inter3));
  inv1  gate2791(.a(s_321), .O(gate111inter4));
  nand2 gate2792(.a(gate111inter4), .b(gate111inter3), .O(gate111inter5));
  nor2  gate2793(.a(gate111inter5), .b(gate111inter2), .O(gate111inter6));
  inv1  gate2794(.a(G374), .O(gate111inter7));
  inv1  gate2795(.a(G375), .O(gate111inter8));
  nand2 gate2796(.a(gate111inter8), .b(gate111inter7), .O(gate111inter9));
  nand2 gate2797(.a(s_321), .b(gate111inter3), .O(gate111inter10));
  nor2  gate2798(.a(gate111inter10), .b(gate111inter9), .O(gate111inter11));
  nor2  gate2799(.a(gate111inter11), .b(gate111inter6), .O(gate111inter12));
  nand2 gate2800(.a(gate111inter12), .b(gate111inter1), .O(G444));
nand2 gate112( .a(G376), .b(G377), .O(G447) );
nand2 gate113( .a(G378), .b(G379), .O(G450) );
nand2 gate114( .a(G380), .b(G381), .O(G453) );
nand2 gate115( .a(G382), .b(G383), .O(G456) );
nand2 gate116( .a(G384), .b(G385), .O(G459) );

  xor2  gate1387(.a(G387), .b(G386), .O(gate117inter0));
  nand2 gate1388(.a(gate117inter0), .b(s_120), .O(gate117inter1));
  and2  gate1389(.a(G387), .b(G386), .O(gate117inter2));
  inv1  gate1390(.a(s_120), .O(gate117inter3));
  inv1  gate1391(.a(s_121), .O(gate117inter4));
  nand2 gate1392(.a(gate117inter4), .b(gate117inter3), .O(gate117inter5));
  nor2  gate1393(.a(gate117inter5), .b(gate117inter2), .O(gate117inter6));
  inv1  gate1394(.a(G386), .O(gate117inter7));
  inv1  gate1395(.a(G387), .O(gate117inter8));
  nand2 gate1396(.a(gate117inter8), .b(gate117inter7), .O(gate117inter9));
  nand2 gate1397(.a(s_121), .b(gate117inter3), .O(gate117inter10));
  nor2  gate1398(.a(gate117inter10), .b(gate117inter9), .O(gate117inter11));
  nor2  gate1399(.a(gate117inter11), .b(gate117inter6), .O(gate117inter12));
  nand2 gate1400(.a(gate117inter12), .b(gate117inter1), .O(G462));
nand2 gate118( .a(G388), .b(G389), .O(G465) );
nand2 gate119( .a(G390), .b(G391), .O(G468) );
nand2 gate120( .a(G392), .b(G393), .O(G471) );
nand2 gate121( .a(G394), .b(G395), .O(G474) );
nand2 gate122( .a(G396), .b(G397), .O(G477) );

  xor2  gate2885(.a(G399), .b(G398), .O(gate123inter0));
  nand2 gate2886(.a(gate123inter0), .b(s_334), .O(gate123inter1));
  and2  gate2887(.a(G399), .b(G398), .O(gate123inter2));
  inv1  gate2888(.a(s_334), .O(gate123inter3));
  inv1  gate2889(.a(s_335), .O(gate123inter4));
  nand2 gate2890(.a(gate123inter4), .b(gate123inter3), .O(gate123inter5));
  nor2  gate2891(.a(gate123inter5), .b(gate123inter2), .O(gate123inter6));
  inv1  gate2892(.a(G398), .O(gate123inter7));
  inv1  gate2893(.a(G399), .O(gate123inter8));
  nand2 gate2894(.a(gate123inter8), .b(gate123inter7), .O(gate123inter9));
  nand2 gate2895(.a(s_335), .b(gate123inter3), .O(gate123inter10));
  nor2  gate2896(.a(gate123inter10), .b(gate123inter9), .O(gate123inter11));
  nor2  gate2897(.a(gate123inter11), .b(gate123inter6), .O(gate123inter12));
  nand2 gate2898(.a(gate123inter12), .b(gate123inter1), .O(G480));

  xor2  gate3151(.a(G401), .b(G400), .O(gate124inter0));
  nand2 gate3152(.a(gate124inter0), .b(s_372), .O(gate124inter1));
  and2  gate3153(.a(G401), .b(G400), .O(gate124inter2));
  inv1  gate3154(.a(s_372), .O(gate124inter3));
  inv1  gate3155(.a(s_373), .O(gate124inter4));
  nand2 gate3156(.a(gate124inter4), .b(gate124inter3), .O(gate124inter5));
  nor2  gate3157(.a(gate124inter5), .b(gate124inter2), .O(gate124inter6));
  inv1  gate3158(.a(G400), .O(gate124inter7));
  inv1  gate3159(.a(G401), .O(gate124inter8));
  nand2 gate3160(.a(gate124inter8), .b(gate124inter7), .O(gate124inter9));
  nand2 gate3161(.a(s_373), .b(gate124inter3), .O(gate124inter10));
  nor2  gate3162(.a(gate124inter10), .b(gate124inter9), .O(gate124inter11));
  nor2  gate3163(.a(gate124inter11), .b(gate124inter6), .O(gate124inter12));
  nand2 gate3164(.a(gate124inter12), .b(gate124inter1), .O(G483));
nand2 gate125( .a(G402), .b(G403), .O(G486) );

  xor2  gate2213(.a(G405), .b(G404), .O(gate126inter0));
  nand2 gate2214(.a(gate126inter0), .b(s_238), .O(gate126inter1));
  and2  gate2215(.a(G405), .b(G404), .O(gate126inter2));
  inv1  gate2216(.a(s_238), .O(gate126inter3));
  inv1  gate2217(.a(s_239), .O(gate126inter4));
  nand2 gate2218(.a(gate126inter4), .b(gate126inter3), .O(gate126inter5));
  nor2  gate2219(.a(gate126inter5), .b(gate126inter2), .O(gate126inter6));
  inv1  gate2220(.a(G404), .O(gate126inter7));
  inv1  gate2221(.a(G405), .O(gate126inter8));
  nand2 gate2222(.a(gate126inter8), .b(gate126inter7), .O(gate126inter9));
  nand2 gate2223(.a(s_239), .b(gate126inter3), .O(gate126inter10));
  nor2  gate2224(.a(gate126inter10), .b(gate126inter9), .O(gate126inter11));
  nor2  gate2225(.a(gate126inter11), .b(gate126inter6), .O(gate126inter12));
  nand2 gate2226(.a(gate126inter12), .b(gate126inter1), .O(G489));

  xor2  gate1191(.a(G407), .b(G406), .O(gate127inter0));
  nand2 gate1192(.a(gate127inter0), .b(s_92), .O(gate127inter1));
  and2  gate1193(.a(G407), .b(G406), .O(gate127inter2));
  inv1  gate1194(.a(s_92), .O(gate127inter3));
  inv1  gate1195(.a(s_93), .O(gate127inter4));
  nand2 gate1196(.a(gate127inter4), .b(gate127inter3), .O(gate127inter5));
  nor2  gate1197(.a(gate127inter5), .b(gate127inter2), .O(gate127inter6));
  inv1  gate1198(.a(G406), .O(gate127inter7));
  inv1  gate1199(.a(G407), .O(gate127inter8));
  nand2 gate1200(.a(gate127inter8), .b(gate127inter7), .O(gate127inter9));
  nand2 gate1201(.a(s_93), .b(gate127inter3), .O(gate127inter10));
  nor2  gate1202(.a(gate127inter10), .b(gate127inter9), .O(gate127inter11));
  nor2  gate1203(.a(gate127inter11), .b(gate127inter6), .O(gate127inter12));
  nand2 gate1204(.a(gate127inter12), .b(gate127inter1), .O(G492));

  xor2  gate2815(.a(G409), .b(G408), .O(gate128inter0));
  nand2 gate2816(.a(gate128inter0), .b(s_324), .O(gate128inter1));
  and2  gate2817(.a(G409), .b(G408), .O(gate128inter2));
  inv1  gate2818(.a(s_324), .O(gate128inter3));
  inv1  gate2819(.a(s_325), .O(gate128inter4));
  nand2 gate2820(.a(gate128inter4), .b(gate128inter3), .O(gate128inter5));
  nor2  gate2821(.a(gate128inter5), .b(gate128inter2), .O(gate128inter6));
  inv1  gate2822(.a(G408), .O(gate128inter7));
  inv1  gate2823(.a(G409), .O(gate128inter8));
  nand2 gate2824(.a(gate128inter8), .b(gate128inter7), .O(gate128inter9));
  nand2 gate2825(.a(s_325), .b(gate128inter3), .O(gate128inter10));
  nor2  gate2826(.a(gate128inter10), .b(gate128inter9), .O(gate128inter11));
  nor2  gate2827(.a(gate128inter11), .b(gate128inter6), .O(gate128inter12));
  nand2 gate2828(.a(gate128inter12), .b(gate128inter1), .O(G495));

  xor2  gate1429(.a(G411), .b(G410), .O(gate129inter0));
  nand2 gate1430(.a(gate129inter0), .b(s_126), .O(gate129inter1));
  and2  gate1431(.a(G411), .b(G410), .O(gate129inter2));
  inv1  gate1432(.a(s_126), .O(gate129inter3));
  inv1  gate1433(.a(s_127), .O(gate129inter4));
  nand2 gate1434(.a(gate129inter4), .b(gate129inter3), .O(gate129inter5));
  nor2  gate1435(.a(gate129inter5), .b(gate129inter2), .O(gate129inter6));
  inv1  gate1436(.a(G410), .O(gate129inter7));
  inv1  gate1437(.a(G411), .O(gate129inter8));
  nand2 gate1438(.a(gate129inter8), .b(gate129inter7), .O(gate129inter9));
  nand2 gate1439(.a(s_127), .b(gate129inter3), .O(gate129inter10));
  nor2  gate1440(.a(gate129inter10), .b(gate129inter9), .O(gate129inter11));
  nor2  gate1441(.a(gate129inter11), .b(gate129inter6), .O(gate129inter12));
  nand2 gate1442(.a(gate129inter12), .b(gate129inter1), .O(G498));

  xor2  gate2955(.a(G413), .b(G412), .O(gate130inter0));
  nand2 gate2956(.a(gate130inter0), .b(s_344), .O(gate130inter1));
  and2  gate2957(.a(G413), .b(G412), .O(gate130inter2));
  inv1  gate2958(.a(s_344), .O(gate130inter3));
  inv1  gate2959(.a(s_345), .O(gate130inter4));
  nand2 gate2960(.a(gate130inter4), .b(gate130inter3), .O(gate130inter5));
  nor2  gate2961(.a(gate130inter5), .b(gate130inter2), .O(gate130inter6));
  inv1  gate2962(.a(G412), .O(gate130inter7));
  inv1  gate2963(.a(G413), .O(gate130inter8));
  nand2 gate2964(.a(gate130inter8), .b(gate130inter7), .O(gate130inter9));
  nand2 gate2965(.a(s_345), .b(gate130inter3), .O(gate130inter10));
  nor2  gate2966(.a(gate130inter10), .b(gate130inter9), .O(gate130inter11));
  nor2  gate2967(.a(gate130inter11), .b(gate130inter6), .O(gate130inter12));
  nand2 gate2968(.a(gate130inter12), .b(gate130inter1), .O(G501));
nand2 gate131( .a(G414), .b(G415), .O(G504) );
nand2 gate132( .a(G416), .b(G417), .O(G507) );
nand2 gate133( .a(G418), .b(G419), .O(G510) );
nand2 gate134( .a(G420), .b(G421), .O(G513) );

  xor2  gate1555(.a(G423), .b(G422), .O(gate135inter0));
  nand2 gate1556(.a(gate135inter0), .b(s_144), .O(gate135inter1));
  and2  gate1557(.a(G423), .b(G422), .O(gate135inter2));
  inv1  gate1558(.a(s_144), .O(gate135inter3));
  inv1  gate1559(.a(s_145), .O(gate135inter4));
  nand2 gate1560(.a(gate135inter4), .b(gate135inter3), .O(gate135inter5));
  nor2  gate1561(.a(gate135inter5), .b(gate135inter2), .O(gate135inter6));
  inv1  gate1562(.a(G422), .O(gate135inter7));
  inv1  gate1563(.a(G423), .O(gate135inter8));
  nand2 gate1564(.a(gate135inter8), .b(gate135inter7), .O(gate135inter9));
  nand2 gate1565(.a(s_145), .b(gate135inter3), .O(gate135inter10));
  nor2  gate1566(.a(gate135inter10), .b(gate135inter9), .O(gate135inter11));
  nor2  gate1567(.a(gate135inter11), .b(gate135inter6), .O(gate135inter12));
  nand2 gate1568(.a(gate135inter12), .b(gate135inter1), .O(G516));
nand2 gate136( .a(G424), .b(G425), .O(G519) );

  xor2  gate1289(.a(G429), .b(G426), .O(gate137inter0));
  nand2 gate1290(.a(gate137inter0), .b(s_106), .O(gate137inter1));
  and2  gate1291(.a(G429), .b(G426), .O(gate137inter2));
  inv1  gate1292(.a(s_106), .O(gate137inter3));
  inv1  gate1293(.a(s_107), .O(gate137inter4));
  nand2 gate1294(.a(gate137inter4), .b(gate137inter3), .O(gate137inter5));
  nor2  gate1295(.a(gate137inter5), .b(gate137inter2), .O(gate137inter6));
  inv1  gate1296(.a(G426), .O(gate137inter7));
  inv1  gate1297(.a(G429), .O(gate137inter8));
  nand2 gate1298(.a(gate137inter8), .b(gate137inter7), .O(gate137inter9));
  nand2 gate1299(.a(s_107), .b(gate137inter3), .O(gate137inter10));
  nor2  gate1300(.a(gate137inter10), .b(gate137inter9), .O(gate137inter11));
  nor2  gate1301(.a(gate137inter11), .b(gate137inter6), .O(gate137inter12));
  nand2 gate1302(.a(gate137inter12), .b(gate137inter1), .O(G522));

  xor2  gate603(.a(G435), .b(G432), .O(gate138inter0));
  nand2 gate604(.a(gate138inter0), .b(s_8), .O(gate138inter1));
  and2  gate605(.a(G435), .b(G432), .O(gate138inter2));
  inv1  gate606(.a(s_8), .O(gate138inter3));
  inv1  gate607(.a(s_9), .O(gate138inter4));
  nand2 gate608(.a(gate138inter4), .b(gate138inter3), .O(gate138inter5));
  nor2  gate609(.a(gate138inter5), .b(gate138inter2), .O(gate138inter6));
  inv1  gate610(.a(G432), .O(gate138inter7));
  inv1  gate611(.a(G435), .O(gate138inter8));
  nand2 gate612(.a(gate138inter8), .b(gate138inter7), .O(gate138inter9));
  nand2 gate613(.a(s_9), .b(gate138inter3), .O(gate138inter10));
  nor2  gate614(.a(gate138inter10), .b(gate138inter9), .O(gate138inter11));
  nor2  gate615(.a(gate138inter11), .b(gate138inter6), .O(gate138inter12));
  nand2 gate616(.a(gate138inter12), .b(gate138inter1), .O(G525));

  xor2  gate1331(.a(G441), .b(G438), .O(gate139inter0));
  nand2 gate1332(.a(gate139inter0), .b(s_112), .O(gate139inter1));
  and2  gate1333(.a(G441), .b(G438), .O(gate139inter2));
  inv1  gate1334(.a(s_112), .O(gate139inter3));
  inv1  gate1335(.a(s_113), .O(gate139inter4));
  nand2 gate1336(.a(gate139inter4), .b(gate139inter3), .O(gate139inter5));
  nor2  gate1337(.a(gate139inter5), .b(gate139inter2), .O(gate139inter6));
  inv1  gate1338(.a(G438), .O(gate139inter7));
  inv1  gate1339(.a(G441), .O(gate139inter8));
  nand2 gate1340(.a(gate139inter8), .b(gate139inter7), .O(gate139inter9));
  nand2 gate1341(.a(s_113), .b(gate139inter3), .O(gate139inter10));
  nor2  gate1342(.a(gate139inter10), .b(gate139inter9), .O(gate139inter11));
  nor2  gate1343(.a(gate139inter11), .b(gate139inter6), .O(gate139inter12));
  nand2 gate1344(.a(gate139inter12), .b(gate139inter1), .O(G528));
nand2 gate140( .a(G444), .b(G447), .O(G531) );
nand2 gate141( .a(G450), .b(G453), .O(G534) );

  xor2  gate1849(.a(G459), .b(G456), .O(gate142inter0));
  nand2 gate1850(.a(gate142inter0), .b(s_186), .O(gate142inter1));
  and2  gate1851(.a(G459), .b(G456), .O(gate142inter2));
  inv1  gate1852(.a(s_186), .O(gate142inter3));
  inv1  gate1853(.a(s_187), .O(gate142inter4));
  nand2 gate1854(.a(gate142inter4), .b(gate142inter3), .O(gate142inter5));
  nor2  gate1855(.a(gate142inter5), .b(gate142inter2), .O(gate142inter6));
  inv1  gate1856(.a(G456), .O(gate142inter7));
  inv1  gate1857(.a(G459), .O(gate142inter8));
  nand2 gate1858(.a(gate142inter8), .b(gate142inter7), .O(gate142inter9));
  nand2 gate1859(.a(s_187), .b(gate142inter3), .O(gate142inter10));
  nor2  gate1860(.a(gate142inter10), .b(gate142inter9), .O(gate142inter11));
  nor2  gate1861(.a(gate142inter11), .b(gate142inter6), .O(gate142inter12));
  nand2 gate1862(.a(gate142inter12), .b(gate142inter1), .O(G537));

  xor2  gate2703(.a(G465), .b(G462), .O(gate143inter0));
  nand2 gate2704(.a(gate143inter0), .b(s_308), .O(gate143inter1));
  and2  gate2705(.a(G465), .b(G462), .O(gate143inter2));
  inv1  gate2706(.a(s_308), .O(gate143inter3));
  inv1  gate2707(.a(s_309), .O(gate143inter4));
  nand2 gate2708(.a(gate143inter4), .b(gate143inter3), .O(gate143inter5));
  nor2  gate2709(.a(gate143inter5), .b(gate143inter2), .O(gate143inter6));
  inv1  gate2710(.a(G462), .O(gate143inter7));
  inv1  gate2711(.a(G465), .O(gate143inter8));
  nand2 gate2712(.a(gate143inter8), .b(gate143inter7), .O(gate143inter9));
  nand2 gate2713(.a(s_309), .b(gate143inter3), .O(gate143inter10));
  nor2  gate2714(.a(gate143inter10), .b(gate143inter9), .O(gate143inter11));
  nor2  gate2715(.a(gate143inter11), .b(gate143inter6), .O(gate143inter12));
  nand2 gate2716(.a(gate143inter12), .b(gate143inter1), .O(G540));
nand2 gate144( .a(G468), .b(G471), .O(G543) );
nand2 gate145( .a(G474), .b(G477), .O(G546) );
nand2 gate146( .a(G480), .b(G483), .O(G549) );

  xor2  gate2269(.a(G489), .b(G486), .O(gate147inter0));
  nand2 gate2270(.a(gate147inter0), .b(s_246), .O(gate147inter1));
  and2  gate2271(.a(G489), .b(G486), .O(gate147inter2));
  inv1  gate2272(.a(s_246), .O(gate147inter3));
  inv1  gate2273(.a(s_247), .O(gate147inter4));
  nand2 gate2274(.a(gate147inter4), .b(gate147inter3), .O(gate147inter5));
  nor2  gate2275(.a(gate147inter5), .b(gate147inter2), .O(gate147inter6));
  inv1  gate2276(.a(G486), .O(gate147inter7));
  inv1  gate2277(.a(G489), .O(gate147inter8));
  nand2 gate2278(.a(gate147inter8), .b(gate147inter7), .O(gate147inter9));
  nand2 gate2279(.a(s_247), .b(gate147inter3), .O(gate147inter10));
  nor2  gate2280(.a(gate147inter10), .b(gate147inter9), .O(gate147inter11));
  nor2  gate2281(.a(gate147inter11), .b(gate147inter6), .O(gate147inter12));
  nand2 gate2282(.a(gate147inter12), .b(gate147inter1), .O(G552));
nand2 gate148( .a(G492), .b(G495), .O(G555) );
nand2 gate149( .a(G498), .b(G501), .O(G558) );

  xor2  gate1821(.a(G507), .b(G504), .O(gate150inter0));
  nand2 gate1822(.a(gate150inter0), .b(s_182), .O(gate150inter1));
  and2  gate1823(.a(G507), .b(G504), .O(gate150inter2));
  inv1  gate1824(.a(s_182), .O(gate150inter3));
  inv1  gate1825(.a(s_183), .O(gate150inter4));
  nand2 gate1826(.a(gate150inter4), .b(gate150inter3), .O(gate150inter5));
  nor2  gate1827(.a(gate150inter5), .b(gate150inter2), .O(gate150inter6));
  inv1  gate1828(.a(G504), .O(gate150inter7));
  inv1  gate1829(.a(G507), .O(gate150inter8));
  nand2 gate1830(.a(gate150inter8), .b(gate150inter7), .O(gate150inter9));
  nand2 gate1831(.a(s_183), .b(gate150inter3), .O(gate150inter10));
  nor2  gate1832(.a(gate150inter10), .b(gate150inter9), .O(gate150inter11));
  nor2  gate1833(.a(gate150inter11), .b(gate150inter6), .O(gate150inter12));
  nand2 gate1834(.a(gate150inter12), .b(gate150inter1), .O(G561));
nand2 gate151( .a(G510), .b(G513), .O(G564) );
nand2 gate152( .a(G516), .b(G519), .O(G567) );

  xor2  gate3249(.a(G522), .b(G426), .O(gate153inter0));
  nand2 gate3250(.a(gate153inter0), .b(s_386), .O(gate153inter1));
  and2  gate3251(.a(G522), .b(G426), .O(gate153inter2));
  inv1  gate3252(.a(s_386), .O(gate153inter3));
  inv1  gate3253(.a(s_387), .O(gate153inter4));
  nand2 gate3254(.a(gate153inter4), .b(gate153inter3), .O(gate153inter5));
  nor2  gate3255(.a(gate153inter5), .b(gate153inter2), .O(gate153inter6));
  inv1  gate3256(.a(G426), .O(gate153inter7));
  inv1  gate3257(.a(G522), .O(gate153inter8));
  nand2 gate3258(.a(gate153inter8), .b(gate153inter7), .O(gate153inter9));
  nand2 gate3259(.a(s_387), .b(gate153inter3), .O(gate153inter10));
  nor2  gate3260(.a(gate153inter10), .b(gate153inter9), .O(gate153inter11));
  nor2  gate3261(.a(gate153inter11), .b(gate153inter6), .O(gate153inter12));
  nand2 gate3262(.a(gate153inter12), .b(gate153inter1), .O(G570));

  xor2  gate2283(.a(G522), .b(G429), .O(gate154inter0));
  nand2 gate2284(.a(gate154inter0), .b(s_248), .O(gate154inter1));
  and2  gate2285(.a(G522), .b(G429), .O(gate154inter2));
  inv1  gate2286(.a(s_248), .O(gate154inter3));
  inv1  gate2287(.a(s_249), .O(gate154inter4));
  nand2 gate2288(.a(gate154inter4), .b(gate154inter3), .O(gate154inter5));
  nor2  gate2289(.a(gate154inter5), .b(gate154inter2), .O(gate154inter6));
  inv1  gate2290(.a(G429), .O(gate154inter7));
  inv1  gate2291(.a(G522), .O(gate154inter8));
  nand2 gate2292(.a(gate154inter8), .b(gate154inter7), .O(gate154inter9));
  nand2 gate2293(.a(s_249), .b(gate154inter3), .O(gate154inter10));
  nor2  gate2294(.a(gate154inter10), .b(gate154inter9), .O(gate154inter11));
  nor2  gate2295(.a(gate154inter11), .b(gate154inter6), .O(gate154inter12));
  nand2 gate2296(.a(gate154inter12), .b(gate154inter1), .O(G571));

  xor2  gate2605(.a(G525), .b(G432), .O(gate155inter0));
  nand2 gate2606(.a(gate155inter0), .b(s_294), .O(gate155inter1));
  and2  gate2607(.a(G525), .b(G432), .O(gate155inter2));
  inv1  gate2608(.a(s_294), .O(gate155inter3));
  inv1  gate2609(.a(s_295), .O(gate155inter4));
  nand2 gate2610(.a(gate155inter4), .b(gate155inter3), .O(gate155inter5));
  nor2  gate2611(.a(gate155inter5), .b(gate155inter2), .O(gate155inter6));
  inv1  gate2612(.a(G432), .O(gate155inter7));
  inv1  gate2613(.a(G525), .O(gate155inter8));
  nand2 gate2614(.a(gate155inter8), .b(gate155inter7), .O(gate155inter9));
  nand2 gate2615(.a(s_295), .b(gate155inter3), .O(gate155inter10));
  nor2  gate2616(.a(gate155inter10), .b(gate155inter9), .O(gate155inter11));
  nor2  gate2617(.a(gate155inter11), .b(gate155inter6), .O(gate155inter12));
  nand2 gate2618(.a(gate155inter12), .b(gate155inter1), .O(G572));
nand2 gate156( .a(G435), .b(G525), .O(G573) );

  xor2  gate1317(.a(G528), .b(G438), .O(gate157inter0));
  nand2 gate1318(.a(gate157inter0), .b(s_110), .O(gate157inter1));
  and2  gate1319(.a(G528), .b(G438), .O(gate157inter2));
  inv1  gate1320(.a(s_110), .O(gate157inter3));
  inv1  gate1321(.a(s_111), .O(gate157inter4));
  nand2 gate1322(.a(gate157inter4), .b(gate157inter3), .O(gate157inter5));
  nor2  gate1323(.a(gate157inter5), .b(gate157inter2), .O(gate157inter6));
  inv1  gate1324(.a(G438), .O(gate157inter7));
  inv1  gate1325(.a(G528), .O(gate157inter8));
  nand2 gate1326(.a(gate157inter8), .b(gate157inter7), .O(gate157inter9));
  nand2 gate1327(.a(s_111), .b(gate157inter3), .O(gate157inter10));
  nor2  gate1328(.a(gate157inter10), .b(gate157inter9), .O(gate157inter11));
  nor2  gate1329(.a(gate157inter11), .b(gate157inter6), .O(gate157inter12));
  nand2 gate1330(.a(gate157inter12), .b(gate157inter1), .O(G574));
nand2 gate158( .a(G441), .b(G528), .O(G575) );

  xor2  gate1009(.a(G531), .b(G444), .O(gate159inter0));
  nand2 gate1010(.a(gate159inter0), .b(s_66), .O(gate159inter1));
  and2  gate1011(.a(G531), .b(G444), .O(gate159inter2));
  inv1  gate1012(.a(s_66), .O(gate159inter3));
  inv1  gate1013(.a(s_67), .O(gate159inter4));
  nand2 gate1014(.a(gate159inter4), .b(gate159inter3), .O(gate159inter5));
  nor2  gate1015(.a(gate159inter5), .b(gate159inter2), .O(gate159inter6));
  inv1  gate1016(.a(G444), .O(gate159inter7));
  inv1  gate1017(.a(G531), .O(gate159inter8));
  nand2 gate1018(.a(gate159inter8), .b(gate159inter7), .O(gate159inter9));
  nand2 gate1019(.a(s_67), .b(gate159inter3), .O(gate159inter10));
  nor2  gate1020(.a(gate159inter10), .b(gate159inter9), .O(gate159inter11));
  nor2  gate1021(.a(gate159inter11), .b(gate159inter6), .O(gate159inter12));
  nand2 gate1022(.a(gate159inter12), .b(gate159inter1), .O(G576));

  xor2  gate2829(.a(G531), .b(G447), .O(gate160inter0));
  nand2 gate2830(.a(gate160inter0), .b(s_326), .O(gate160inter1));
  and2  gate2831(.a(G531), .b(G447), .O(gate160inter2));
  inv1  gate2832(.a(s_326), .O(gate160inter3));
  inv1  gate2833(.a(s_327), .O(gate160inter4));
  nand2 gate2834(.a(gate160inter4), .b(gate160inter3), .O(gate160inter5));
  nor2  gate2835(.a(gate160inter5), .b(gate160inter2), .O(gate160inter6));
  inv1  gate2836(.a(G447), .O(gate160inter7));
  inv1  gate2837(.a(G531), .O(gate160inter8));
  nand2 gate2838(.a(gate160inter8), .b(gate160inter7), .O(gate160inter9));
  nand2 gate2839(.a(s_327), .b(gate160inter3), .O(gate160inter10));
  nor2  gate2840(.a(gate160inter10), .b(gate160inter9), .O(gate160inter11));
  nor2  gate2841(.a(gate160inter11), .b(gate160inter6), .O(gate160inter12));
  nand2 gate2842(.a(gate160inter12), .b(gate160inter1), .O(G577));
nand2 gate161( .a(G450), .b(G534), .O(G578) );

  xor2  gate2073(.a(G534), .b(G453), .O(gate162inter0));
  nand2 gate2074(.a(gate162inter0), .b(s_218), .O(gate162inter1));
  and2  gate2075(.a(G534), .b(G453), .O(gate162inter2));
  inv1  gate2076(.a(s_218), .O(gate162inter3));
  inv1  gate2077(.a(s_219), .O(gate162inter4));
  nand2 gate2078(.a(gate162inter4), .b(gate162inter3), .O(gate162inter5));
  nor2  gate2079(.a(gate162inter5), .b(gate162inter2), .O(gate162inter6));
  inv1  gate2080(.a(G453), .O(gate162inter7));
  inv1  gate2081(.a(G534), .O(gate162inter8));
  nand2 gate2082(.a(gate162inter8), .b(gate162inter7), .O(gate162inter9));
  nand2 gate2083(.a(s_219), .b(gate162inter3), .O(gate162inter10));
  nor2  gate2084(.a(gate162inter10), .b(gate162inter9), .O(gate162inter11));
  nor2  gate2085(.a(gate162inter11), .b(gate162inter6), .O(gate162inter12));
  nand2 gate2086(.a(gate162inter12), .b(gate162inter1), .O(G579));
nand2 gate163( .a(G456), .b(G537), .O(G580) );
nand2 gate164( .a(G459), .b(G537), .O(G581) );
nand2 gate165( .a(G462), .b(G540), .O(G582) );
nand2 gate166( .a(G465), .b(G540), .O(G583) );

  xor2  gate3263(.a(G543), .b(G468), .O(gate167inter0));
  nand2 gate3264(.a(gate167inter0), .b(s_388), .O(gate167inter1));
  and2  gate3265(.a(G543), .b(G468), .O(gate167inter2));
  inv1  gate3266(.a(s_388), .O(gate167inter3));
  inv1  gate3267(.a(s_389), .O(gate167inter4));
  nand2 gate3268(.a(gate167inter4), .b(gate167inter3), .O(gate167inter5));
  nor2  gate3269(.a(gate167inter5), .b(gate167inter2), .O(gate167inter6));
  inv1  gate3270(.a(G468), .O(gate167inter7));
  inv1  gate3271(.a(G543), .O(gate167inter8));
  nand2 gate3272(.a(gate167inter8), .b(gate167inter7), .O(gate167inter9));
  nand2 gate3273(.a(s_389), .b(gate167inter3), .O(gate167inter10));
  nor2  gate3274(.a(gate167inter10), .b(gate167inter9), .O(gate167inter11));
  nor2  gate3275(.a(gate167inter11), .b(gate167inter6), .O(gate167inter12));
  nand2 gate3276(.a(gate167inter12), .b(gate167inter1), .O(G584));

  xor2  gate1835(.a(G543), .b(G471), .O(gate168inter0));
  nand2 gate1836(.a(gate168inter0), .b(s_184), .O(gate168inter1));
  and2  gate1837(.a(G543), .b(G471), .O(gate168inter2));
  inv1  gate1838(.a(s_184), .O(gate168inter3));
  inv1  gate1839(.a(s_185), .O(gate168inter4));
  nand2 gate1840(.a(gate168inter4), .b(gate168inter3), .O(gate168inter5));
  nor2  gate1841(.a(gate168inter5), .b(gate168inter2), .O(gate168inter6));
  inv1  gate1842(.a(G471), .O(gate168inter7));
  inv1  gate1843(.a(G543), .O(gate168inter8));
  nand2 gate1844(.a(gate168inter8), .b(gate168inter7), .O(gate168inter9));
  nand2 gate1845(.a(s_185), .b(gate168inter3), .O(gate168inter10));
  nor2  gate1846(.a(gate168inter10), .b(gate168inter9), .O(gate168inter11));
  nor2  gate1847(.a(gate168inter11), .b(gate168inter6), .O(gate168inter12));
  nand2 gate1848(.a(gate168inter12), .b(gate168inter1), .O(G585));
nand2 gate169( .a(G474), .b(G546), .O(G586) );
nand2 gate170( .a(G477), .b(G546), .O(G587) );

  xor2  gate3011(.a(G549), .b(G480), .O(gate171inter0));
  nand2 gate3012(.a(gate171inter0), .b(s_352), .O(gate171inter1));
  and2  gate3013(.a(G549), .b(G480), .O(gate171inter2));
  inv1  gate3014(.a(s_352), .O(gate171inter3));
  inv1  gate3015(.a(s_353), .O(gate171inter4));
  nand2 gate3016(.a(gate171inter4), .b(gate171inter3), .O(gate171inter5));
  nor2  gate3017(.a(gate171inter5), .b(gate171inter2), .O(gate171inter6));
  inv1  gate3018(.a(G480), .O(gate171inter7));
  inv1  gate3019(.a(G549), .O(gate171inter8));
  nand2 gate3020(.a(gate171inter8), .b(gate171inter7), .O(gate171inter9));
  nand2 gate3021(.a(s_353), .b(gate171inter3), .O(gate171inter10));
  nor2  gate3022(.a(gate171inter10), .b(gate171inter9), .O(gate171inter11));
  nor2  gate3023(.a(gate171inter11), .b(gate171inter6), .O(gate171inter12));
  nand2 gate3024(.a(gate171inter12), .b(gate171inter1), .O(G588));
nand2 gate172( .a(G483), .b(G549), .O(G589) );

  xor2  gate1779(.a(G552), .b(G486), .O(gate173inter0));
  nand2 gate1780(.a(gate173inter0), .b(s_176), .O(gate173inter1));
  and2  gate1781(.a(G552), .b(G486), .O(gate173inter2));
  inv1  gate1782(.a(s_176), .O(gate173inter3));
  inv1  gate1783(.a(s_177), .O(gate173inter4));
  nand2 gate1784(.a(gate173inter4), .b(gate173inter3), .O(gate173inter5));
  nor2  gate1785(.a(gate173inter5), .b(gate173inter2), .O(gate173inter6));
  inv1  gate1786(.a(G486), .O(gate173inter7));
  inv1  gate1787(.a(G552), .O(gate173inter8));
  nand2 gate1788(.a(gate173inter8), .b(gate173inter7), .O(gate173inter9));
  nand2 gate1789(.a(s_177), .b(gate173inter3), .O(gate173inter10));
  nor2  gate1790(.a(gate173inter10), .b(gate173inter9), .O(gate173inter11));
  nor2  gate1791(.a(gate173inter11), .b(gate173inter6), .O(gate173inter12));
  nand2 gate1792(.a(gate173inter12), .b(gate173inter1), .O(G590));
nand2 gate174( .a(G489), .b(G552), .O(G591) );

  xor2  gate1247(.a(G555), .b(G492), .O(gate175inter0));
  nand2 gate1248(.a(gate175inter0), .b(s_100), .O(gate175inter1));
  and2  gate1249(.a(G555), .b(G492), .O(gate175inter2));
  inv1  gate1250(.a(s_100), .O(gate175inter3));
  inv1  gate1251(.a(s_101), .O(gate175inter4));
  nand2 gate1252(.a(gate175inter4), .b(gate175inter3), .O(gate175inter5));
  nor2  gate1253(.a(gate175inter5), .b(gate175inter2), .O(gate175inter6));
  inv1  gate1254(.a(G492), .O(gate175inter7));
  inv1  gate1255(.a(G555), .O(gate175inter8));
  nand2 gate1256(.a(gate175inter8), .b(gate175inter7), .O(gate175inter9));
  nand2 gate1257(.a(s_101), .b(gate175inter3), .O(gate175inter10));
  nor2  gate1258(.a(gate175inter10), .b(gate175inter9), .O(gate175inter11));
  nor2  gate1259(.a(gate175inter11), .b(gate175inter6), .O(gate175inter12));
  nand2 gate1260(.a(gate175inter12), .b(gate175inter1), .O(G592));
nand2 gate176( .a(G495), .b(G555), .O(G593) );

  xor2  gate3277(.a(G558), .b(G498), .O(gate177inter0));
  nand2 gate3278(.a(gate177inter0), .b(s_390), .O(gate177inter1));
  and2  gate3279(.a(G558), .b(G498), .O(gate177inter2));
  inv1  gate3280(.a(s_390), .O(gate177inter3));
  inv1  gate3281(.a(s_391), .O(gate177inter4));
  nand2 gate3282(.a(gate177inter4), .b(gate177inter3), .O(gate177inter5));
  nor2  gate3283(.a(gate177inter5), .b(gate177inter2), .O(gate177inter6));
  inv1  gate3284(.a(G498), .O(gate177inter7));
  inv1  gate3285(.a(G558), .O(gate177inter8));
  nand2 gate3286(.a(gate177inter8), .b(gate177inter7), .O(gate177inter9));
  nand2 gate3287(.a(s_391), .b(gate177inter3), .O(gate177inter10));
  nor2  gate3288(.a(gate177inter10), .b(gate177inter9), .O(gate177inter11));
  nor2  gate3289(.a(gate177inter11), .b(gate177inter6), .O(gate177inter12));
  nand2 gate3290(.a(gate177inter12), .b(gate177inter1), .O(G594));

  xor2  gate1303(.a(G558), .b(G501), .O(gate178inter0));
  nand2 gate1304(.a(gate178inter0), .b(s_108), .O(gate178inter1));
  and2  gate1305(.a(G558), .b(G501), .O(gate178inter2));
  inv1  gate1306(.a(s_108), .O(gate178inter3));
  inv1  gate1307(.a(s_109), .O(gate178inter4));
  nand2 gate1308(.a(gate178inter4), .b(gate178inter3), .O(gate178inter5));
  nor2  gate1309(.a(gate178inter5), .b(gate178inter2), .O(gate178inter6));
  inv1  gate1310(.a(G501), .O(gate178inter7));
  inv1  gate1311(.a(G558), .O(gate178inter8));
  nand2 gate1312(.a(gate178inter8), .b(gate178inter7), .O(gate178inter9));
  nand2 gate1313(.a(s_109), .b(gate178inter3), .O(gate178inter10));
  nor2  gate1314(.a(gate178inter10), .b(gate178inter9), .O(gate178inter11));
  nor2  gate1315(.a(gate178inter11), .b(gate178inter6), .O(gate178inter12));
  nand2 gate1316(.a(gate178inter12), .b(gate178inter1), .O(G595));

  xor2  gate2423(.a(G561), .b(G504), .O(gate179inter0));
  nand2 gate2424(.a(gate179inter0), .b(s_268), .O(gate179inter1));
  and2  gate2425(.a(G561), .b(G504), .O(gate179inter2));
  inv1  gate2426(.a(s_268), .O(gate179inter3));
  inv1  gate2427(.a(s_269), .O(gate179inter4));
  nand2 gate2428(.a(gate179inter4), .b(gate179inter3), .O(gate179inter5));
  nor2  gate2429(.a(gate179inter5), .b(gate179inter2), .O(gate179inter6));
  inv1  gate2430(.a(G504), .O(gate179inter7));
  inv1  gate2431(.a(G561), .O(gate179inter8));
  nand2 gate2432(.a(gate179inter8), .b(gate179inter7), .O(gate179inter9));
  nand2 gate2433(.a(s_269), .b(gate179inter3), .O(gate179inter10));
  nor2  gate2434(.a(gate179inter10), .b(gate179inter9), .O(gate179inter11));
  nor2  gate2435(.a(gate179inter11), .b(gate179inter6), .O(gate179inter12));
  nand2 gate2436(.a(gate179inter12), .b(gate179inter1), .O(G596));
nand2 gate180( .a(G507), .b(G561), .O(G597) );
nand2 gate181( .a(G510), .b(G564), .O(G598) );
nand2 gate182( .a(G513), .b(G564), .O(G599) );

  xor2  gate1653(.a(G567), .b(G516), .O(gate183inter0));
  nand2 gate1654(.a(gate183inter0), .b(s_158), .O(gate183inter1));
  and2  gate1655(.a(G567), .b(G516), .O(gate183inter2));
  inv1  gate1656(.a(s_158), .O(gate183inter3));
  inv1  gate1657(.a(s_159), .O(gate183inter4));
  nand2 gate1658(.a(gate183inter4), .b(gate183inter3), .O(gate183inter5));
  nor2  gate1659(.a(gate183inter5), .b(gate183inter2), .O(gate183inter6));
  inv1  gate1660(.a(G516), .O(gate183inter7));
  inv1  gate1661(.a(G567), .O(gate183inter8));
  nand2 gate1662(.a(gate183inter8), .b(gate183inter7), .O(gate183inter9));
  nand2 gate1663(.a(s_159), .b(gate183inter3), .O(gate183inter10));
  nor2  gate1664(.a(gate183inter10), .b(gate183inter9), .O(gate183inter11));
  nor2  gate1665(.a(gate183inter11), .b(gate183inter6), .O(gate183inter12));
  nand2 gate1666(.a(gate183inter12), .b(gate183inter1), .O(G600));
nand2 gate184( .a(G519), .b(G567), .O(G601) );

  xor2  gate1345(.a(G571), .b(G570), .O(gate185inter0));
  nand2 gate1346(.a(gate185inter0), .b(s_114), .O(gate185inter1));
  and2  gate1347(.a(G571), .b(G570), .O(gate185inter2));
  inv1  gate1348(.a(s_114), .O(gate185inter3));
  inv1  gate1349(.a(s_115), .O(gate185inter4));
  nand2 gate1350(.a(gate185inter4), .b(gate185inter3), .O(gate185inter5));
  nor2  gate1351(.a(gate185inter5), .b(gate185inter2), .O(gate185inter6));
  inv1  gate1352(.a(G570), .O(gate185inter7));
  inv1  gate1353(.a(G571), .O(gate185inter8));
  nand2 gate1354(.a(gate185inter8), .b(gate185inter7), .O(gate185inter9));
  nand2 gate1355(.a(s_115), .b(gate185inter3), .O(gate185inter10));
  nor2  gate1356(.a(gate185inter10), .b(gate185inter9), .O(gate185inter11));
  nor2  gate1357(.a(gate185inter11), .b(gate185inter6), .O(gate185inter12));
  nand2 gate1358(.a(gate185inter12), .b(gate185inter1), .O(G602));
nand2 gate186( .a(G572), .b(G573), .O(G607) );
nand2 gate187( .a(G574), .b(G575), .O(G612) );

  xor2  gate2647(.a(G577), .b(G576), .O(gate188inter0));
  nand2 gate2648(.a(gate188inter0), .b(s_300), .O(gate188inter1));
  and2  gate2649(.a(G577), .b(G576), .O(gate188inter2));
  inv1  gate2650(.a(s_300), .O(gate188inter3));
  inv1  gate2651(.a(s_301), .O(gate188inter4));
  nand2 gate2652(.a(gate188inter4), .b(gate188inter3), .O(gate188inter5));
  nor2  gate2653(.a(gate188inter5), .b(gate188inter2), .O(gate188inter6));
  inv1  gate2654(.a(G576), .O(gate188inter7));
  inv1  gate2655(.a(G577), .O(gate188inter8));
  nand2 gate2656(.a(gate188inter8), .b(gate188inter7), .O(gate188inter9));
  nand2 gate2657(.a(s_301), .b(gate188inter3), .O(gate188inter10));
  nor2  gate2658(.a(gate188inter10), .b(gate188inter9), .O(gate188inter11));
  nor2  gate2659(.a(gate188inter11), .b(gate188inter6), .O(gate188inter12));
  nand2 gate2660(.a(gate188inter12), .b(gate188inter1), .O(G617));
nand2 gate189( .a(G578), .b(G579), .O(G622) );

  xor2  gate967(.a(G581), .b(G580), .O(gate190inter0));
  nand2 gate968(.a(gate190inter0), .b(s_60), .O(gate190inter1));
  and2  gate969(.a(G581), .b(G580), .O(gate190inter2));
  inv1  gate970(.a(s_60), .O(gate190inter3));
  inv1  gate971(.a(s_61), .O(gate190inter4));
  nand2 gate972(.a(gate190inter4), .b(gate190inter3), .O(gate190inter5));
  nor2  gate973(.a(gate190inter5), .b(gate190inter2), .O(gate190inter6));
  inv1  gate974(.a(G580), .O(gate190inter7));
  inv1  gate975(.a(G581), .O(gate190inter8));
  nand2 gate976(.a(gate190inter8), .b(gate190inter7), .O(gate190inter9));
  nand2 gate977(.a(s_61), .b(gate190inter3), .O(gate190inter10));
  nor2  gate978(.a(gate190inter10), .b(gate190inter9), .O(gate190inter11));
  nor2  gate979(.a(gate190inter11), .b(gate190inter6), .O(gate190inter12));
  nand2 gate980(.a(gate190inter12), .b(gate190inter1), .O(G627));

  xor2  gate1681(.a(G583), .b(G582), .O(gate191inter0));
  nand2 gate1682(.a(gate191inter0), .b(s_162), .O(gate191inter1));
  and2  gate1683(.a(G583), .b(G582), .O(gate191inter2));
  inv1  gate1684(.a(s_162), .O(gate191inter3));
  inv1  gate1685(.a(s_163), .O(gate191inter4));
  nand2 gate1686(.a(gate191inter4), .b(gate191inter3), .O(gate191inter5));
  nor2  gate1687(.a(gate191inter5), .b(gate191inter2), .O(gate191inter6));
  inv1  gate1688(.a(G582), .O(gate191inter7));
  inv1  gate1689(.a(G583), .O(gate191inter8));
  nand2 gate1690(.a(gate191inter8), .b(gate191inter7), .O(gate191inter9));
  nand2 gate1691(.a(s_163), .b(gate191inter3), .O(gate191inter10));
  nor2  gate1692(.a(gate191inter10), .b(gate191inter9), .O(gate191inter11));
  nor2  gate1693(.a(gate191inter11), .b(gate191inter6), .O(gate191inter12));
  nand2 gate1694(.a(gate191inter12), .b(gate191inter1), .O(G632));

  xor2  gate1023(.a(G585), .b(G584), .O(gate192inter0));
  nand2 gate1024(.a(gate192inter0), .b(s_68), .O(gate192inter1));
  and2  gate1025(.a(G585), .b(G584), .O(gate192inter2));
  inv1  gate1026(.a(s_68), .O(gate192inter3));
  inv1  gate1027(.a(s_69), .O(gate192inter4));
  nand2 gate1028(.a(gate192inter4), .b(gate192inter3), .O(gate192inter5));
  nor2  gate1029(.a(gate192inter5), .b(gate192inter2), .O(gate192inter6));
  inv1  gate1030(.a(G584), .O(gate192inter7));
  inv1  gate1031(.a(G585), .O(gate192inter8));
  nand2 gate1032(.a(gate192inter8), .b(gate192inter7), .O(gate192inter9));
  nand2 gate1033(.a(s_69), .b(gate192inter3), .O(gate192inter10));
  nor2  gate1034(.a(gate192inter10), .b(gate192inter9), .O(gate192inter11));
  nor2  gate1035(.a(gate192inter11), .b(gate192inter6), .O(gate192inter12));
  nand2 gate1036(.a(gate192inter12), .b(gate192inter1), .O(G637));
nand2 gate193( .a(G586), .b(G587), .O(G642) );

  xor2  gate2157(.a(G589), .b(G588), .O(gate194inter0));
  nand2 gate2158(.a(gate194inter0), .b(s_230), .O(gate194inter1));
  and2  gate2159(.a(G589), .b(G588), .O(gate194inter2));
  inv1  gate2160(.a(s_230), .O(gate194inter3));
  inv1  gate2161(.a(s_231), .O(gate194inter4));
  nand2 gate2162(.a(gate194inter4), .b(gate194inter3), .O(gate194inter5));
  nor2  gate2163(.a(gate194inter5), .b(gate194inter2), .O(gate194inter6));
  inv1  gate2164(.a(G588), .O(gate194inter7));
  inv1  gate2165(.a(G589), .O(gate194inter8));
  nand2 gate2166(.a(gate194inter8), .b(gate194inter7), .O(gate194inter9));
  nand2 gate2167(.a(s_231), .b(gate194inter3), .O(gate194inter10));
  nor2  gate2168(.a(gate194inter10), .b(gate194inter9), .O(gate194inter11));
  nor2  gate2169(.a(gate194inter11), .b(gate194inter6), .O(gate194inter12));
  nand2 gate2170(.a(gate194inter12), .b(gate194inter1), .O(G645));

  xor2  gate2591(.a(G591), .b(G590), .O(gate195inter0));
  nand2 gate2592(.a(gate195inter0), .b(s_292), .O(gate195inter1));
  and2  gate2593(.a(G591), .b(G590), .O(gate195inter2));
  inv1  gate2594(.a(s_292), .O(gate195inter3));
  inv1  gate2595(.a(s_293), .O(gate195inter4));
  nand2 gate2596(.a(gate195inter4), .b(gate195inter3), .O(gate195inter5));
  nor2  gate2597(.a(gate195inter5), .b(gate195inter2), .O(gate195inter6));
  inv1  gate2598(.a(G590), .O(gate195inter7));
  inv1  gate2599(.a(G591), .O(gate195inter8));
  nand2 gate2600(.a(gate195inter8), .b(gate195inter7), .O(gate195inter9));
  nand2 gate2601(.a(s_293), .b(gate195inter3), .O(gate195inter10));
  nor2  gate2602(.a(gate195inter10), .b(gate195inter9), .O(gate195inter11));
  nor2  gate2603(.a(gate195inter11), .b(gate195inter6), .O(gate195inter12));
  nand2 gate2604(.a(gate195inter12), .b(gate195inter1), .O(G648));
nand2 gate196( .a(G592), .b(G593), .O(G651) );
nand2 gate197( .a(G594), .b(G595), .O(G654) );

  xor2  gate883(.a(G597), .b(G596), .O(gate198inter0));
  nand2 gate884(.a(gate198inter0), .b(s_48), .O(gate198inter1));
  and2  gate885(.a(G597), .b(G596), .O(gate198inter2));
  inv1  gate886(.a(s_48), .O(gate198inter3));
  inv1  gate887(.a(s_49), .O(gate198inter4));
  nand2 gate888(.a(gate198inter4), .b(gate198inter3), .O(gate198inter5));
  nor2  gate889(.a(gate198inter5), .b(gate198inter2), .O(gate198inter6));
  inv1  gate890(.a(G596), .O(gate198inter7));
  inv1  gate891(.a(G597), .O(gate198inter8));
  nand2 gate892(.a(gate198inter8), .b(gate198inter7), .O(gate198inter9));
  nand2 gate893(.a(s_49), .b(gate198inter3), .O(gate198inter10));
  nor2  gate894(.a(gate198inter10), .b(gate198inter9), .O(gate198inter11));
  nor2  gate895(.a(gate198inter11), .b(gate198inter6), .O(gate198inter12));
  nand2 gate896(.a(gate198inter12), .b(gate198inter1), .O(G657));
nand2 gate199( .a(G598), .b(G599), .O(G660) );
nand2 gate200( .a(G600), .b(G601), .O(G663) );
nand2 gate201( .a(G602), .b(G607), .O(G666) );

  xor2  gate3235(.a(G617), .b(G612), .O(gate202inter0));
  nand2 gate3236(.a(gate202inter0), .b(s_384), .O(gate202inter1));
  and2  gate3237(.a(G617), .b(G612), .O(gate202inter2));
  inv1  gate3238(.a(s_384), .O(gate202inter3));
  inv1  gate3239(.a(s_385), .O(gate202inter4));
  nand2 gate3240(.a(gate202inter4), .b(gate202inter3), .O(gate202inter5));
  nor2  gate3241(.a(gate202inter5), .b(gate202inter2), .O(gate202inter6));
  inv1  gate3242(.a(G612), .O(gate202inter7));
  inv1  gate3243(.a(G617), .O(gate202inter8));
  nand2 gate3244(.a(gate202inter8), .b(gate202inter7), .O(gate202inter9));
  nand2 gate3245(.a(s_385), .b(gate202inter3), .O(gate202inter10));
  nor2  gate3246(.a(gate202inter10), .b(gate202inter9), .O(gate202inter11));
  nor2  gate3247(.a(gate202inter11), .b(gate202inter6), .O(gate202inter12));
  nand2 gate3248(.a(gate202inter12), .b(gate202inter1), .O(G669));

  xor2  gate1933(.a(G612), .b(G602), .O(gate203inter0));
  nand2 gate1934(.a(gate203inter0), .b(s_198), .O(gate203inter1));
  and2  gate1935(.a(G612), .b(G602), .O(gate203inter2));
  inv1  gate1936(.a(s_198), .O(gate203inter3));
  inv1  gate1937(.a(s_199), .O(gate203inter4));
  nand2 gate1938(.a(gate203inter4), .b(gate203inter3), .O(gate203inter5));
  nor2  gate1939(.a(gate203inter5), .b(gate203inter2), .O(gate203inter6));
  inv1  gate1940(.a(G602), .O(gate203inter7));
  inv1  gate1941(.a(G612), .O(gate203inter8));
  nand2 gate1942(.a(gate203inter8), .b(gate203inter7), .O(gate203inter9));
  nand2 gate1943(.a(s_199), .b(gate203inter3), .O(gate203inter10));
  nor2  gate1944(.a(gate203inter10), .b(gate203inter9), .O(gate203inter11));
  nor2  gate1945(.a(gate203inter11), .b(gate203inter6), .O(gate203inter12));
  nand2 gate1946(.a(gate203inter12), .b(gate203inter1), .O(G672));

  xor2  gate953(.a(G617), .b(G607), .O(gate204inter0));
  nand2 gate954(.a(gate204inter0), .b(s_58), .O(gate204inter1));
  and2  gate955(.a(G617), .b(G607), .O(gate204inter2));
  inv1  gate956(.a(s_58), .O(gate204inter3));
  inv1  gate957(.a(s_59), .O(gate204inter4));
  nand2 gate958(.a(gate204inter4), .b(gate204inter3), .O(gate204inter5));
  nor2  gate959(.a(gate204inter5), .b(gate204inter2), .O(gate204inter6));
  inv1  gate960(.a(G607), .O(gate204inter7));
  inv1  gate961(.a(G617), .O(gate204inter8));
  nand2 gate962(.a(gate204inter8), .b(gate204inter7), .O(gate204inter9));
  nand2 gate963(.a(s_59), .b(gate204inter3), .O(gate204inter10));
  nor2  gate964(.a(gate204inter10), .b(gate204inter9), .O(gate204inter11));
  nor2  gate965(.a(gate204inter11), .b(gate204inter6), .O(gate204inter12));
  nand2 gate966(.a(gate204inter12), .b(gate204inter1), .O(G675));
nand2 gate205( .a(G622), .b(G627), .O(G678) );
nand2 gate206( .a(G632), .b(G637), .O(G681) );
nand2 gate207( .a(G622), .b(G632), .O(G684) );
nand2 gate208( .a(G627), .b(G637), .O(G687) );
nand2 gate209( .a(G602), .b(G666), .O(G690) );
nand2 gate210( .a(G607), .b(G666), .O(G691) );

  xor2  gate2003(.a(G669), .b(G612), .O(gate211inter0));
  nand2 gate2004(.a(gate211inter0), .b(s_208), .O(gate211inter1));
  and2  gate2005(.a(G669), .b(G612), .O(gate211inter2));
  inv1  gate2006(.a(s_208), .O(gate211inter3));
  inv1  gate2007(.a(s_209), .O(gate211inter4));
  nand2 gate2008(.a(gate211inter4), .b(gate211inter3), .O(gate211inter5));
  nor2  gate2009(.a(gate211inter5), .b(gate211inter2), .O(gate211inter6));
  inv1  gate2010(.a(G612), .O(gate211inter7));
  inv1  gate2011(.a(G669), .O(gate211inter8));
  nand2 gate2012(.a(gate211inter8), .b(gate211inter7), .O(gate211inter9));
  nand2 gate2013(.a(s_209), .b(gate211inter3), .O(gate211inter10));
  nor2  gate2014(.a(gate211inter10), .b(gate211inter9), .O(gate211inter11));
  nor2  gate2015(.a(gate211inter11), .b(gate211inter6), .O(gate211inter12));
  nand2 gate2016(.a(gate211inter12), .b(gate211inter1), .O(G692));
nand2 gate212( .a(G617), .b(G669), .O(G693) );
nand2 gate213( .a(G602), .b(G672), .O(G694) );
nand2 gate214( .a(G612), .b(G672), .O(G695) );

  xor2  gate2367(.a(G675), .b(G607), .O(gate215inter0));
  nand2 gate2368(.a(gate215inter0), .b(s_260), .O(gate215inter1));
  and2  gate2369(.a(G675), .b(G607), .O(gate215inter2));
  inv1  gate2370(.a(s_260), .O(gate215inter3));
  inv1  gate2371(.a(s_261), .O(gate215inter4));
  nand2 gate2372(.a(gate215inter4), .b(gate215inter3), .O(gate215inter5));
  nor2  gate2373(.a(gate215inter5), .b(gate215inter2), .O(gate215inter6));
  inv1  gate2374(.a(G607), .O(gate215inter7));
  inv1  gate2375(.a(G675), .O(gate215inter8));
  nand2 gate2376(.a(gate215inter8), .b(gate215inter7), .O(gate215inter9));
  nand2 gate2377(.a(s_261), .b(gate215inter3), .O(gate215inter10));
  nor2  gate2378(.a(gate215inter10), .b(gate215inter9), .O(gate215inter11));
  nor2  gate2379(.a(gate215inter11), .b(gate215inter6), .O(gate215inter12));
  nand2 gate2380(.a(gate215inter12), .b(gate215inter1), .O(G696));

  xor2  gate2745(.a(G675), .b(G617), .O(gate216inter0));
  nand2 gate2746(.a(gate216inter0), .b(s_314), .O(gate216inter1));
  and2  gate2747(.a(G675), .b(G617), .O(gate216inter2));
  inv1  gate2748(.a(s_314), .O(gate216inter3));
  inv1  gate2749(.a(s_315), .O(gate216inter4));
  nand2 gate2750(.a(gate216inter4), .b(gate216inter3), .O(gate216inter5));
  nor2  gate2751(.a(gate216inter5), .b(gate216inter2), .O(gate216inter6));
  inv1  gate2752(.a(G617), .O(gate216inter7));
  inv1  gate2753(.a(G675), .O(gate216inter8));
  nand2 gate2754(.a(gate216inter8), .b(gate216inter7), .O(gate216inter9));
  nand2 gate2755(.a(s_315), .b(gate216inter3), .O(gate216inter10));
  nor2  gate2756(.a(gate216inter10), .b(gate216inter9), .O(gate216inter11));
  nor2  gate2757(.a(gate216inter11), .b(gate216inter6), .O(gate216inter12));
  nand2 gate2758(.a(gate216inter12), .b(gate216inter1), .O(G697));

  xor2  gate1051(.a(G678), .b(G622), .O(gate217inter0));
  nand2 gate1052(.a(gate217inter0), .b(s_72), .O(gate217inter1));
  and2  gate1053(.a(G678), .b(G622), .O(gate217inter2));
  inv1  gate1054(.a(s_72), .O(gate217inter3));
  inv1  gate1055(.a(s_73), .O(gate217inter4));
  nand2 gate1056(.a(gate217inter4), .b(gate217inter3), .O(gate217inter5));
  nor2  gate1057(.a(gate217inter5), .b(gate217inter2), .O(gate217inter6));
  inv1  gate1058(.a(G622), .O(gate217inter7));
  inv1  gate1059(.a(G678), .O(gate217inter8));
  nand2 gate1060(.a(gate217inter8), .b(gate217inter7), .O(gate217inter9));
  nand2 gate1061(.a(s_73), .b(gate217inter3), .O(gate217inter10));
  nor2  gate1062(.a(gate217inter10), .b(gate217inter9), .O(gate217inter11));
  nor2  gate1063(.a(gate217inter11), .b(gate217inter6), .O(gate217inter12));
  nand2 gate1064(.a(gate217inter12), .b(gate217inter1), .O(G698));
nand2 gate218( .a(G627), .b(G678), .O(G699) );

  xor2  gate2773(.a(G681), .b(G632), .O(gate219inter0));
  nand2 gate2774(.a(gate219inter0), .b(s_318), .O(gate219inter1));
  and2  gate2775(.a(G681), .b(G632), .O(gate219inter2));
  inv1  gate2776(.a(s_318), .O(gate219inter3));
  inv1  gate2777(.a(s_319), .O(gate219inter4));
  nand2 gate2778(.a(gate219inter4), .b(gate219inter3), .O(gate219inter5));
  nor2  gate2779(.a(gate219inter5), .b(gate219inter2), .O(gate219inter6));
  inv1  gate2780(.a(G632), .O(gate219inter7));
  inv1  gate2781(.a(G681), .O(gate219inter8));
  nand2 gate2782(.a(gate219inter8), .b(gate219inter7), .O(gate219inter9));
  nand2 gate2783(.a(s_319), .b(gate219inter3), .O(gate219inter10));
  nor2  gate2784(.a(gate219inter10), .b(gate219inter9), .O(gate219inter11));
  nor2  gate2785(.a(gate219inter11), .b(gate219inter6), .O(gate219inter12));
  nand2 gate2786(.a(gate219inter12), .b(gate219inter1), .O(G700));
nand2 gate220( .a(G637), .b(G681), .O(G701) );

  xor2  gate939(.a(G684), .b(G622), .O(gate221inter0));
  nand2 gate940(.a(gate221inter0), .b(s_56), .O(gate221inter1));
  and2  gate941(.a(G684), .b(G622), .O(gate221inter2));
  inv1  gate942(.a(s_56), .O(gate221inter3));
  inv1  gate943(.a(s_57), .O(gate221inter4));
  nand2 gate944(.a(gate221inter4), .b(gate221inter3), .O(gate221inter5));
  nor2  gate945(.a(gate221inter5), .b(gate221inter2), .O(gate221inter6));
  inv1  gate946(.a(G622), .O(gate221inter7));
  inv1  gate947(.a(G684), .O(gate221inter8));
  nand2 gate948(.a(gate221inter8), .b(gate221inter7), .O(gate221inter9));
  nand2 gate949(.a(s_57), .b(gate221inter3), .O(gate221inter10));
  nor2  gate950(.a(gate221inter10), .b(gate221inter9), .O(gate221inter11));
  nor2  gate951(.a(gate221inter11), .b(gate221inter6), .O(gate221inter12));
  nand2 gate952(.a(gate221inter12), .b(gate221inter1), .O(G702));

  xor2  gate645(.a(G684), .b(G632), .O(gate222inter0));
  nand2 gate646(.a(gate222inter0), .b(s_14), .O(gate222inter1));
  and2  gate647(.a(G684), .b(G632), .O(gate222inter2));
  inv1  gate648(.a(s_14), .O(gate222inter3));
  inv1  gate649(.a(s_15), .O(gate222inter4));
  nand2 gate650(.a(gate222inter4), .b(gate222inter3), .O(gate222inter5));
  nor2  gate651(.a(gate222inter5), .b(gate222inter2), .O(gate222inter6));
  inv1  gate652(.a(G632), .O(gate222inter7));
  inv1  gate653(.a(G684), .O(gate222inter8));
  nand2 gate654(.a(gate222inter8), .b(gate222inter7), .O(gate222inter9));
  nand2 gate655(.a(s_15), .b(gate222inter3), .O(gate222inter10));
  nor2  gate656(.a(gate222inter10), .b(gate222inter9), .O(gate222inter11));
  nor2  gate657(.a(gate222inter11), .b(gate222inter6), .O(gate222inter12));
  nand2 gate658(.a(gate222inter12), .b(gate222inter1), .O(G703));
nand2 gate223( .a(G627), .b(G687), .O(G704) );
nand2 gate224( .a(G637), .b(G687), .O(G705) );

  xor2  gate1807(.a(G691), .b(G690), .O(gate225inter0));
  nand2 gate1808(.a(gate225inter0), .b(s_180), .O(gate225inter1));
  and2  gate1809(.a(G691), .b(G690), .O(gate225inter2));
  inv1  gate1810(.a(s_180), .O(gate225inter3));
  inv1  gate1811(.a(s_181), .O(gate225inter4));
  nand2 gate1812(.a(gate225inter4), .b(gate225inter3), .O(gate225inter5));
  nor2  gate1813(.a(gate225inter5), .b(gate225inter2), .O(gate225inter6));
  inv1  gate1814(.a(G690), .O(gate225inter7));
  inv1  gate1815(.a(G691), .O(gate225inter8));
  nand2 gate1816(.a(gate225inter8), .b(gate225inter7), .O(gate225inter9));
  nand2 gate1817(.a(s_181), .b(gate225inter3), .O(gate225inter10));
  nor2  gate1818(.a(gate225inter10), .b(gate225inter9), .O(gate225inter11));
  nor2  gate1819(.a(gate225inter11), .b(gate225inter6), .O(gate225inter12));
  nand2 gate1820(.a(gate225inter12), .b(gate225inter1), .O(G706));
nand2 gate226( .a(G692), .b(G693), .O(G709) );

  xor2  gate1079(.a(G695), .b(G694), .O(gate227inter0));
  nand2 gate1080(.a(gate227inter0), .b(s_76), .O(gate227inter1));
  and2  gate1081(.a(G695), .b(G694), .O(gate227inter2));
  inv1  gate1082(.a(s_76), .O(gate227inter3));
  inv1  gate1083(.a(s_77), .O(gate227inter4));
  nand2 gate1084(.a(gate227inter4), .b(gate227inter3), .O(gate227inter5));
  nor2  gate1085(.a(gate227inter5), .b(gate227inter2), .O(gate227inter6));
  inv1  gate1086(.a(G694), .O(gate227inter7));
  inv1  gate1087(.a(G695), .O(gate227inter8));
  nand2 gate1088(.a(gate227inter8), .b(gate227inter7), .O(gate227inter9));
  nand2 gate1089(.a(s_77), .b(gate227inter3), .O(gate227inter10));
  nor2  gate1090(.a(gate227inter10), .b(gate227inter9), .O(gate227inter11));
  nor2  gate1091(.a(gate227inter11), .b(gate227inter6), .O(gate227inter12));
  nand2 gate1092(.a(gate227inter12), .b(gate227inter1), .O(G712));
nand2 gate228( .a(G696), .b(G697), .O(G715) );
nand2 gate229( .a(G698), .b(G699), .O(G718) );
nand2 gate230( .a(G700), .b(G701), .O(G721) );
nand2 gate231( .a(G702), .b(G703), .O(G724) );
nand2 gate232( .a(G704), .b(G705), .O(G727) );
nand2 gate233( .a(G242), .b(G718), .O(G730) );

  xor2  gate2661(.a(G721), .b(G245), .O(gate234inter0));
  nand2 gate2662(.a(gate234inter0), .b(s_302), .O(gate234inter1));
  and2  gate2663(.a(G721), .b(G245), .O(gate234inter2));
  inv1  gate2664(.a(s_302), .O(gate234inter3));
  inv1  gate2665(.a(s_303), .O(gate234inter4));
  nand2 gate2666(.a(gate234inter4), .b(gate234inter3), .O(gate234inter5));
  nor2  gate2667(.a(gate234inter5), .b(gate234inter2), .O(gate234inter6));
  inv1  gate2668(.a(G245), .O(gate234inter7));
  inv1  gate2669(.a(G721), .O(gate234inter8));
  nand2 gate2670(.a(gate234inter8), .b(gate234inter7), .O(gate234inter9));
  nand2 gate2671(.a(s_303), .b(gate234inter3), .O(gate234inter10));
  nor2  gate2672(.a(gate234inter10), .b(gate234inter9), .O(gate234inter11));
  nor2  gate2673(.a(gate234inter11), .b(gate234inter6), .O(gate234inter12));
  nand2 gate2674(.a(gate234inter12), .b(gate234inter1), .O(G733));
nand2 gate235( .a(G248), .b(G724), .O(G736) );
nand2 gate236( .a(G251), .b(G727), .O(G739) );
nand2 gate237( .a(G254), .b(G706), .O(G742) );
nand2 gate238( .a(G257), .b(G709), .O(G745) );

  xor2  gate1037(.a(G712), .b(G260), .O(gate239inter0));
  nand2 gate1038(.a(gate239inter0), .b(s_70), .O(gate239inter1));
  and2  gate1039(.a(G712), .b(G260), .O(gate239inter2));
  inv1  gate1040(.a(s_70), .O(gate239inter3));
  inv1  gate1041(.a(s_71), .O(gate239inter4));
  nand2 gate1042(.a(gate239inter4), .b(gate239inter3), .O(gate239inter5));
  nor2  gate1043(.a(gate239inter5), .b(gate239inter2), .O(gate239inter6));
  inv1  gate1044(.a(G260), .O(gate239inter7));
  inv1  gate1045(.a(G712), .O(gate239inter8));
  nand2 gate1046(.a(gate239inter8), .b(gate239inter7), .O(gate239inter9));
  nand2 gate1047(.a(s_71), .b(gate239inter3), .O(gate239inter10));
  nor2  gate1048(.a(gate239inter10), .b(gate239inter9), .O(gate239inter11));
  nor2  gate1049(.a(gate239inter11), .b(gate239inter6), .O(gate239inter12));
  nand2 gate1050(.a(gate239inter12), .b(gate239inter1), .O(G748));

  xor2  gate1359(.a(G715), .b(G263), .O(gate240inter0));
  nand2 gate1360(.a(gate240inter0), .b(s_116), .O(gate240inter1));
  and2  gate1361(.a(G715), .b(G263), .O(gate240inter2));
  inv1  gate1362(.a(s_116), .O(gate240inter3));
  inv1  gate1363(.a(s_117), .O(gate240inter4));
  nand2 gate1364(.a(gate240inter4), .b(gate240inter3), .O(gate240inter5));
  nor2  gate1365(.a(gate240inter5), .b(gate240inter2), .O(gate240inter6));
  inv1  gate1366(.a(G263), .O(gate240inter7));
  inv1  gate1367(.a(G715), .O(gate240inter8));
  nand2 gate1368(.a(gate240inter8), .b(gate240inter7), .O(gate240inter9));
  nand2 gate1369(.a(s_117), .b(gate240inter3), .O(gate240inter10));
  nor2  gate1370(.a(gate240inter10), .b(gate240inter9), .O(gate240inter11));
  nor2  gate1371(.a(gate240inter11), .b(gate240inter6), .O(gate240inter12));
  nand2 gate1372(.a(gate240inter12), .b(gate240inter1), .O(G751));

  xor2  gate2535(.a(G730), .b(G242), .O(gate241inter0));
  nand2 gate2536(.a(gate241inter0), .b(s_284), .O(gate241inter1));
  and2  gate2537(.a(G730), .b(G242), .O(gate241inter2));
  inv1  gate2538(.a(s_284), .O(gate241inter3));
  inv1  gate2539(.a(s_285), .O(gate241inter4));
  nand2 gate2540(.a(gate241inter4), .b(gate241inter3), .O(gate241inter5));
  nor2  gate2541(.a(gate241inter5), .b(gate241inter2), .O(gate241inter6));
  inv1  gate2542(.a(G242), .O(gate241inter7));
  inv1  gate2543(.a(G730), .O(gate241inter8));
  nand2 gate2544(.a(gate241inter8), .b(gate241inter7), .O(gate241inter9));
  nand2 gate2545(.a(s_285), .b(gate241inter3), .O(gate241inter10));
  nor2  gate2546(.a(gate241inter10), .b(gate241inter9), .O(gate241inter11));
  nor2  gate2547(.a(gate241inter11), .b(gate241inter6), .O(gate241inter12));
  nand2 gate2548(.a(gate241inter12), .b(gate241inter1), .O(G754));
nand2 gate242( .a(G718), .b(G730), .O(G755) );
nand2 gate243( .a(G245), .b(G733), .O(G756) );

  xor2  gate1471(.a(G733), .b(G721), .O(gate244inter0));
  nand2 gate1472(.a(gate244inter0), .b(s_132), .O(gate244inter1));
  and2  gate1473(.a(G733), .b(G721), .O(gate244inter2));
  inv1  gate1474(.a(s_132), .O(gate244inter3));
  inv1  gate1475(.a(s_133), .O(gate244inter4));
  nand2 gate1476(.a(gate244inter4), .b(gate244inter3), .O(gate244inter5));
  nor2  gate1477(.a(gate244inter5), .b(gate244inter2), .O(gate244inter6));
  inv1  gate1478(.a(G721), .O(gate244inter7));
  inv1  gate1479(.a(G733), .O(gate244inter8));
  nand2 gate1480(.a(gate244inter8), .b(gate244inter7), .O(gate244inter9));
  nand2 gate1481(.a(s_133), .b(gate244inter3), .O(gate244inter10));
  nor2  gate1482(.a(gate244inter10), .b(gate244inter9), .O(gate244inter11));
  nor2  gate1483(.a(gate244inter11), .b(gate244inter6), .O(gate244inter12));
  nand2 gate1484(.a(gate244inter12), .b(gate244inter1), .O(G757));

  xor2  gate1513(.a(G736), .b(G248), .O(gate245inter0));
  nand2 gate1514(.a(gate245inter0), .b(s_138), .O(gate245inter1));
  and2  gate1515(.a(G736), .b(G248), .O(gate245inter2));
  inv1  gate1516(.a(s_138), .O(gate245inter3));
  inv1  gate1517(.a(s_139), .O(gate245inter4));
  nand2 gate1518(.a(gate245inter4), .b(gate245inter3), .O(gate245inter5));
  nor2  gate1519(.a(gate245inter5), .b(gate245inter2), .O(gate245inter6));
  inv1  gate1520(.a(G248), .O(gate245inter7));
  inv1  gate1521(.a(G736), .O(gate245inter8));
  nand2 gate1522(.a(gate245inter8), .b(gate245inter7), .O(gate245inter9));
  nand2 gate1523(.a(s_139), .b(gate245inter3), .O(gate245inter10));
  nor2  gate1524(.a(gate245inter10), .b(gate245inter9), .O(gate245inter11));
  nor2  gate1525(.a(gate245inter11), .b(gate245inter6), .O(gate245inter12));
  nand2 gate1526(.a(gate245inter12), .b(gate245inter1), .O(G758));

  xor2  gate729(.a(G736), .b(G724), .O(gate246inter0));
  nand2 gate730(.a(gate246inter0), .b(s_26), .O(gate246inter1));
  and2  gate731(.a(G736), .b(G724), .O(gate246inter2));
  inv1  gate732(.a(s_26), .O(gate246inter3));
  inv1  gate733(.a(s_27), .O(gate246inter4));
  nand2 gate734(.a(gate246inter4), .b(gate246inter3), .O(gate246inter5));
  nor2  gate735(.a(gate246inter5), .b(gate246inter2), .O(gate246inter6));
  inv1  gate736(.a(G724), .O(gate246inter7));
  inv1  gate737(.a(G736), .O(gate246inter8));
  nand2 gate738(.a(gate246inter8), .b(gate246inter7), .O(gate246inter9));
  nand2 gate739(.a(s_27), .b(gate246inter3), .O(gate246inter10));
  nor2  gate740(.a(gate246inter10), .b(gate246inter9), .O(gate246inter11));
  nor2  gate741(.a(gate246inter11), .b(gate246inter6), .O(gate246inter12));
  nand2 gate742(.a(gate246inter12), .b(gate246inter1), .O(G759));

  xor2  gate2857(.a(G739), .b(G251), .O(gate247inter0));
  nand2 gate2858(.a(gate247inter0), .b(s_330), .O(gate247inter1));
  and2  gate2859(.a(G739), .b(G251), .O(gate247inter2));
  inv1  gate2860(.a(s_330), .O(gate247inter3));
  inv1  gate2861(.a(s_331), .O(gate247inter4));
  nand2 gate2862(.a(gate247inter4), .b(gate247inter3), .O(gate247inter5));
  nor2  gate2863(.a(gate247inter5), .b(gate247inter2), .O(gate247inter6));
  inv1  gate2864(.a(G251), .O(gate247inter7));
  inv1  gate2865(.a(G739), .O(gate247inter8));
  nand2 gate2866(.a(gate247inter8), .b(gate247inter7), .O(gate247inter9));
  nand2 gate2867(.a(s_331), .b(gate247inter3), .O(gate247inter10));
  nor2  gate2868(.a(gate247inter10), .b(gate247inter9), .O(gate247inter11));
  nor2  gate2869(.a(gate247inter11), .b(gate247inter6), .O(gate247inter12));
  nand2 gate2870(.a(gate247inter12), .b(gate247inter1), .O(G760));

  xor2  gate2255(.a(G739), .b(G727), .O(gate248inter0));
  nand2 gate2256(.a(gate248inter0), .b(s_244), .O(gate248inter1));
  and2  gate2257(.a(G739), .b(G727), .O(gate248inter2));
  inv1  gate2258(.a(s_244), .O(gate248inter3));
  inv1  gate2259(.a(s_245), .O(gate248inter4));
  nand2 gate2260(.a(gate248inter4), .b(gate248inter3), .O(gate248inter5));
  nor2  gate2261(.a(gate248inter5), .b(gate248inter2), .O(gate248inter6));
  inv1  gate2262(.a(G727), .O(gate248inter7));
  inv1  gate2263(.a(G739), .O(gate248inter8));
  nand2 gate2264(.a(gate248inter8), .b(gate248inter7), .O(gate248inter9));
  nand2 gate2265(.a(s_245), .b(gate248inter3), .O(gate248inter10));
  nor2  gate2266(.a(gate248inter10), .b(gate248inter9), .O(gate248inter11));
  nor2  gate2267(.a(gate248inter11), .b(gate248inter6), .O(gate248inter12));
  nand2 gate2268(.a(gate248inter12), .b(gate248inter1), .O(G761));

  xor2  gate1121(.a(G742), .b(G254), .O(gate249inter0));
  nand2 gate1122(.a(gate249inter0), .b(s_82), .O(gate249inter1));
  and2  gate1123(.a(G742), .b(G254), .O(gate249inter2));
  inv1  gate1124(.a(s_82), .O(gate249inter3));
  inv1  gate1125(.a(s_83), .O(gate249inter4));
  nand2 gate1126(.a(gate249inter4), .b(gate249inter3), .O(gate249inter5));
  nor2  gate1127(.a(gate249inter5), .b(gate249inter2), .O(gate249inter6));
  inv1  gate1128(.a(G254), .O(gate249inter7));
  inv1  gate1129(.a(G742), .O(gate249inter8));
  nand2 gate1130(.a(gate249inter8), .b(gate249inter7), .O(gate249inter9));
  nand2 gate1131(.a(s_83), .b(gate249inter3), .O(gate249inter10));
  nor2  gate1132(.a(gate249inter10), .b(gate249inter9), .O(gate249inter11));
  nor2  gate1133(.a(gate249inter11), .b(gate249inter6), .O(gate249inter12));
  nand2 gate1134(.a(gate249inter12), .b(gate249inter1), .O(G762));

  xor2  gate2493(.a(G742), .b(G706), .O(gate250inter0));
  nand2 gate2494(.a(gate250inter0), .b(s_278), .O(gate250inter1));
  and2  gate2495(.a(G742), .b(G706), .O(gate250inter2));
  inv1  gate2496(.a(s_278), .O(gate250inter3));
  inv1  gate2497(.a(s_279), .O(gate250inter4));
  nand2 gate2498(.a(gate250inter4), .b(gate250inter3), .O(gate250inter5));
  nor2  gate2499(.a(gate250inter5), .b(gate250inter2), .O(gate250inter6));
  inv1  gate2500(.a(G706), .O(gate250inter7));
  inv1  gate2501(.a(G742), .O(gate250inter8));
  nand2 gate2502(.a(gate250inter8), .b(gate250inter7), .O(gate250inter9));
  nand2 gate2503(.a(s_279), .b(gate250inter3), .O(gate250inter10));
  nor2  gate2504(.a(gate250inter10), .b(gate250inter9), .O(gate250inter11));
  nor2  gate2505(.a(gate250inter11), .b(gate250inter6), .O(gate250inter12));
  nand2 gate2506(.a(gate250inter12), .b(gate250inter1), .O(G763));

  xor2  gate1261(.a(G745), .b(G257), .O(gate251inter0));
  nand2 gate1262(.a(gate251inter0), .b(s_102), .O(gate251inter1));
  and2  gate1263(.a(G745), .b(G257), .O(gate251inter2));
  inv1  gate1264(.a(s_102), .O(gate251inter3));
  inv1  gate1265(.a(s_103), .O(gate251inter4));
  nand2 gate1266(.a(gate251inter4), .b(gate251inter3), .O(gate251inter5));
  nor2  gate1267(.a(gate251inter5), .b(gate251inter2), .O(gate251inter6));
  inv1  gate1268(.a(G257), .O(gate251inter7));
  inv1  gate1269(.a(G745), .O(gate251inter8));
  nand2 gate1270(.a(gate251inter8), .b(gate251inter7), .O(gate251inter9));
  nand2 gate1271(.a(s_103), .b(gate251inter3), .O(gate251inter10));
  nor2  gate1272(.a(gate251inter10), .b(gate251inter9), .O(gate251inter11));
  nor2  gate1273(.a(gate251inter11), .b(gate251inter6), .O(gate251inter12));
  nand2 gate1274(.a(gate251inter12), .b(gate251inter1), .O(G764));
nand2 gate252( .a(G709), .b(G745), .O(G765) );
nand2 gate253( .a(G260), .b(G748), .O(G766) );

  xor2  gate1233(.a(G748), .b(G712), .O(gate254inter0));
  nand2 gate1234(.a(gate254inter0), .b(s_98), .O(gate254inter1));
  and2  gate1235(.a(G748), .b(G712), .O(gate254inter2));
  inv1  gate1236(.a(s_98), .O(gate254inter3));
  inv1  gate1237(.a(s_99), .O(gate254inter4));
  nand2 gate1238(.a(gate254inter4), .b(gate254inter3), .O(gate254inter5));
  nor2  gate1239(.a(gate254inter5), .b(gate254inter2), .O(gate254inter6));
  inv1  gate1240(.a(G712), .O(gate254inter7));
  inv1  gate1241(.a(G748), .O(gate254inter8));
  nand2 gate1242(.a(gate254inter8), .b(gate254inter7), .O(gate254inter9));
  nand2 gate1243(.a(s_99), .b(gate254inter3), .O(gate254inter10));
  nor2  gate1244(.a(gate254inter10), .b(gate254inter9), .O(gate254inter11));
  nor2  gate1245(.a(gate254inter11), .b(gate254inter6), .O(gate254inter12));
  nand2 gate1246(.a(gate254inter12), .b(gate254inter1), .O(G767));
nand2 gate255( .a(G263), .b(G751), .O(G768) );
nand2 gate256( .a(G715), .b(G751), .O(G769) );
nand2 gate257( .a(G754), .b(G755), .O(G770) );
nand2 gate258( .a(G756), .b(G757), .O(G773) );
nand2 gate259( .a(G758), .b(G759), .O(G776) );
nand2 gate260( .a(G760), .b(G761), .O(G779) );

  xor2  gate1597(.a(G763), .b(G762), .O(gate261inter0));
  nand2 gate1598(.a(gate261inter0), .b(s_150), .O(gate261inter1));
  and2  gate1599(.a(G763), .b(G762), .O(gate261inter2));
  inv1  gate1600(.a(s_150), .O(gate261inter3));
  inv1  gate1601(.a(s_151), .O(gate261inter4));
  nand2 gate1602(.a(gate261inter4), .b(gate261inter3), .O(gate261inter5));
  nor2  gate1603(.a(gate261inter5), .b(gate261inter2), .O(gate261inter6));
  inv1  gate1604(.a(G762), .O(gate261inter7));
  inv1  gate1605(.a(G763), .O(gate261inter8));
  nand2 gate1606(.a(gate261inter8), .b(gate261inter7), .O(gate261inter9));
  nand2 gate1607(.a(s_151), .b(gate261inter3), .O(gate261inter10));
  nor2  gate1608(.a(gate261inter10), .b(gate261inter9), .O(gate261inter11));
  nor2  gate1609(.a(gate261inter11), .b(gate261inter6), .O(gate261inter12));
  nand2 gate1610(.a(gate261inter12), .b(gate261inter1), .O(G782));
nand2 gate262( .a(G764), .b(G765), .O(G785) );
nand2 gate263( .a(G766), .b(G767), .O(G788) );

  xor2  gate3025(.a(G769), .b(G768), .O(gate264inter0));
  nand2 gate3026(.a(gate264inter0), .b(s_354), .O(gate264inter1));
  and2  gate3027(.a(G769), .b(G768), .O(gate264inter2));
  inv1  gate3028(.a(s_354), .O(gate264inter3));
  inv1  gate3029(.a(s_355), .O(gate264inter4));
  nand2 gate3030(.a(gate264inter4), .b(gate264inter3), .O(gate264inter5));
  nor2  gate3031(.a(gate264inter5), .b(gate264inter2), .O(gate264inter6));
  inv1  gate3032(.a(G768), .O(gate264inter7));
  inv1  gate3033(.a(G769), .O(gate264inter8));
  nand2 gate3034(.a(gate264inter8), .b(gate264inter7), .O(gate264inter9));
  nand2 gate3035(.a(s_355), .b(gate264inter3), .O(gate264inter10));
  nor2  gate3036(.a(gate264inter10), .b(gate264inter9), .O(gate264inter11));
  nor2  gate3037(.a(gate264inter11), .b(gate264inter6), .O(gate264inter12));
  nand2 gate3038(.a(gate264inter12), .b(gate264inter1), .O(G791));
nand2 gate265( .a(G642), .b(G770), .O(G794) );

  xor2  gate1443(.a(G773), .b(G645), .O(gate266inter0));
  nand2 gate1444(.a(gate266inter0), .b(s_128), .O(gate266inter1));
  and2  gate1445(.a(G773), .b(G645), .O(gate266inter2));
  inv1  gate1446(.a(s_128), .O(gate266inter3));
  inv1  gate1447(.a(s_129), .O(gate266inter4));
  nand2 gate1448(.a(gate266inter4), .b(gate266inter3), .O(gate266inter5));
  nor2  gate1449(.a(gate266inter5), .b(gate266inter2), .O(gate266inter6));
  inv1  gate1450(.a(G645), .O(gate266inter7));
  inv1  gate1451(.a(G773), .O(gate266inter8));
  nand2 gate1452(.a(gate266inter8), .b(gate266inter7), .O(gate266inter9));
  nand2 gate1453(.a(s_129), .b(gate266inter3), .O(gate266inter10));
  nor2  gate1454(.a(gate266inter10), .b(gate266inter9), .O(gate266inter11));
  nor2  gate1455(.a(gate266inter11), .b(gate266inter6), .O(gate266inter12));
  nand2 gate1456(.a(gate266inter12), .b(gate266inter1), .O(G797));
nand2 gate267( .a(G648), .b(G776), .O(G800) );

  xor2  gate1373(.a(G779), .b(G651), .O(gate268inter0));
  nand2 gate1374(.a(gate268inter0), .b(s_118), .O(gate268inter1));
  and2  gate1375(.a(G779), .b(G651), .O(gate268inter2));
  inv1  gate1376(.a(s_118), .O(gate268inter3));
  inv1  gate1377(.a(s_119), .O(gate268inter4));
  nand2 gate1378(.a(gate268inter4), .b(gate268inter3), .O(gate268inter5));
  nor2  gate1379(.a(gate268inter5), .b(gate268inter2), .O(gate268inter6));
  inv1  gate1380(.a(G651), .O(gate268inter7));
  inv1  gate1381(.a(G779), .O(gate268inter8));
  nand2 gate1382(.a(gate268inter8), .b(gate268inter7), .O(gate268inter9));
  nand2 gate1383(.a(s_119), .b(gate268inter3), .O(gate268inter10));
  nor2  gate1384(.a(gate268inter10), .b(gate268inter9), .O(gate268inter11));
  nor2  gate1385(.a(gate268inter11), .b(gate268inter6), .O(gate268inter12));
  nand2 gate1386(.a(gate268inter12), .b(gate268inter1), .O(G803));

  xor2  gate2409(.a(G782), .b(G654), .O(gate269inter0));
  nand2 gate2410(.a(gate269inter0), .b(s_266), .O(gate269inter1));
  and2  gate2411(.a(G782), .b(G654), .O(gate269inter2));
  inv1  gate2412(.a(s_266), .O(gate269inter3));
  inv1  gate2413(.a(s_267), .O(gate269inter4));
  nand2 gate2414(.a(gate269inter4), .b(gate269inter3), .O(gate269inter5));
  nor2  gate2415(.a(gate269inter5), .b(gate269inter2), .O(gate269inter6));
  inv1  gate2416(.a(G654), .O(gate269inter7));
  inv1  gate2417(.a(G782), .O(gate269inter8));
  nand2 gate2418(.a(gate269inter8), .b(gate269inter7), .O(gate269inter9));
  nand2 gate2419(.a(s_267), .b(gate269inter3), .O(gate269inter10));
  nor2  gate2420(.a(gate269inter10), .b(gate269inter9), .O(gate269inter11));
  nor2  gate2421(.a(gate269inter11), .b(gate269inter6), .O(gate269inter12));
  nand2 gate2422(.a(gate269inter12), .b(gate269inter1), .O(G806));

  xor2  gate2731(.a(G785), .b(G657), .O(gate270inter0));
  nand2 gate2732(.a(gate270inter0), .b(s_312), .O(gate270inter1));
  and2  gate2733(.a(G785), .b(G657), .O(gate270inter2));
  inv1  gate2734(.a(s_312), .O(gate270inter3));
  inv1  gate2735(.a(s_313), .O(gate270inter4));
  nand2 gate2736(.a(gate270inter4), .b(gate270inter3), .O(gate270inter5));
  nor2  gate2737(.a(gate270inter5), .b(gate270inter2), .O(gate270inter6));
  inv1  gate2738(.a(G657), .O(gate270inter7));
  inv1  gate2739(.a(G785), .O(gate270inter8));
  nand2 gate2740(.a(gate270inter8), .b(gate270inter7), .O(gate270inter9));
  nand2 gate2741(.a(s_313), .b(gate270inter3), .O(gate270inter10));
  nor2  gate2742(.a(gate270inter10), .b(gate270inter9), .O(gate270inter11));
  nor2  gate2743(.a(gate270inter11), .b(gate270inter6), .O(gate270inter12));
  nand2 gate2744(.a(gate270inter12), .b(gate270inter1), .O(G809));

  xor2  gate2479(.a(G788), .b(G660), .O(gate271inter0));
  nand2 gate2480(.a(gate271inter0), .b(s_276), .O(gate271inter1));
  and2  gate2481(.a(G788), .b(G660), .O(gate271inter2));
  inv1  gate2482(.a(s_276), .O(gate271inter3));
  inv1  gate2483(.a(s_277), .O(gate271inter4));
  nand2 gate2484(.a(gate271inter4), .b(gate271inter3), .O(gate271inter5));
  nor2  gate2485(.a(gate271inter5), .b(gate271inter2), .O(gate271inter6));
  inv1  gate2486(.a(G660), .O(gate271inter7));
  inv1  gate2487(.a(G788), .O(gate271inter8));
  nand2 gate2488(.a(gate271inter8), .b(gate271inter7), .O(gate271inter9));
  nand2 gate2489(.a(s_277), .b(gate271inter3), .O(gate271inter10));
  nor2  gate2490(.a(gate271inter10), .b(gate271inter9), .O(gate271inter11));
  nor2  gate2491(.a(gate271inter11), .b(gate271inter6), .O(gate271inter12));
  nand2 gate2492(.a(gate271inter12), .b(gate271inter1), .O(G812));

  xor2  gate1639(.a(G791), .b(G663), .O(gate272inter0));
  nand2 gate1640(.a(gate272inter0), .b(s_156), .O(gate272inter1));
  and2  gate1641(.a(G791), .b(G663), .O(gate272inter2));
  inv1  gate1642(.a(s_156), .O(gate272inter3));
  inv1  gate1643(.a(s_157), .O(gate272inter4));
  nand2 gate1644(.a(gate272inter4), .b(gate272inter3), .O(gate272inter5));
  nor2  gate1645(.a(gate272inter5), .b(gate272inter2), .O(gate272inter6));
  inv1  gate1646(.a(G663), .O(gate272inter7));
  inv1  gate1647(.a(G791), .O(gate272inter8));
  nand2 gate1648(.a(gate272inter8), .b(gate272inter7), .O(gate272inter9));
  nand2 gate1649(.a(s_157), .b(gate272inter3), .O(gate272inter10));
  nor2  gate1650(.a(gate272inter10), .b(gate272inter9), .O(gate272inter11));
  nor2  gate1651(.a(gate272inter11), .b(gate272inter6), .O(gate272inter12));
  nand2 gate1652(.a(gate272inter12), .b(gate272inter1), .O(G815));
nand2 gate273( .a(G642), .b(G794), .O(G818) );
nand2 gate274( .a(G770), .b(G794), .O(G819) );
nand2 gate275( .a(G645), .b(G797), .O(G820) );
nand2 gate276( .a(G773), .b(G797), .O(G821) );
nand2 gate277( .a(G648), .b(G800), .O(G822) );

  xor2  gate1975(.a(G800), .b(G776), .O(gate278inter0));
  nand2 gate1976(.a(gate278inter0), .b(s_204), .O(gate278inter1));
  and2  gate1977(.a(G800), .b(G776), .O(gate278inter2));
  inv1  gate1978(.a(s_204), .O(gate278inter3));
  inv1  gate1979(.a(s_205), .O(gate278inter4));
  nand2 gate1980(.a(gate278inter4), .b(gate278inter3), .O(gate278inter5));
  nor2  gate1981(.a(gate278inter5), .b(gate278inter2), .O(gate278inter6));
  inv1  gate1982(.a(G776), .O(gate278inter7));
  inv1  gate1983(.a(G800), .O(gate278inter8));
  nand2 gate1984(.a(gate278inter8), .b(gate278inter7), .O(gate278inter9));
  nand2 gate1985(.a(s_205), .b(gate278inter3), .O(gate278inter10));
  nor2  gate1986(.a(gate278inter10), .b(gate278inter9), .O(gate278inter11));
  nor2  gate1987(.a(gate278inter11), .b(gate278inter6), .O(gate278inter12));
  nand2 gate1988(.a(gate278inter12), .b(gate278inter1), .O(G823));

  xor2  gate1863(.a(G803), .b(G651), .O(gate279inter0));
  nand2 gate1864(.a(gate279inter0), .b(s_188), .O(gate279inter1));
  and2  gate1865(.a(G803), .b(G651), .O(gate279inter2));
  inv1  gate1866(.a(s_188), .O(gate279inter3));
  inv1  gate1867(.a(s_189), .O(gate279inter4));
  nand2 gate1868(.a(gate279inter4), .b(gate279inter3), .O(gate279inter5));
  nor2  gate1869(.a(gate279inter5), .b(gate279inter2), .O(gate279inter6));
  inv1  gate1870(.a(G651), .O(gate279inter7));
  inv1  gate1871(.a(G803), .O(gate279inter8));
  nand2 gate1872(.a(gate279inter8), .b(gate279inter7), .O(gate279inter9));
  nand2 gate1873(.a(s_189), .b(gate279inter3), .O(gate279inter10));
  nor2  gate1874(.a(gate279inter10), .b(gate279inter9), .O(gate279inter11));
  nor2  gate1875(.a(gate279inter11), .b(gate279inter6), .O(gate279inter12));
  nand2 gate1876(.a(gate279inter12), .b(gate279inter1), .O(G824));
nand2 gate280( .a(G779), .b(G803), .O(G825) );

  xor2  gate855(.a(G806), .b(G654), .O(gate281inter0));
  nand2 gate856(.a(gate281inter0), .b(s_44), .O(gate281inter1));
  and2  gate857(.a(G806), .b(G654), .O(gate281inter2));
  inv1  gate858(.a(s_44), .O(gate281inter3));
  inv1  gate859(.a(s_45), .O(gate281inter4));
  nand2 gate860(.a(gate281inter4), .b(gate281inter3), .O(gate281inter5));
  nor2  gate861(.a(gate281inter5), .b(gate281inter2), .O(gate281inter6));
  inv1  gate862(.a(G654), .O(gate281inter7));
  inv1  gate863(.a(G806), .O(gate281inter8));
  nand2 gate864(.a(gate281inter8), .b(gate281inter7), .O(gate281inter9));
  nand2 gate865(.a(s_45), .b(gate281inter3), .O(gate281inter10));
  nor2  gate866(.a(gate281inter10), .b(gate281inter9), .O(gate281inter11));
  nor2  gate867(.a(gate281inter11), .b(gate281inter6), .O(gate281inter12));
  nand2 gate868(.a(gate281inter12), .b(gate281inter1), .O(G826));
nand2 gate282( .a(G782), .b(G806), .O(G827) );
nand2 gate283( .a(G657), .b(G809), .O(G828) );
nand2 gate284( .a(G785), .b(G809), .O(G829) );
nand2 gate285( .a(G660), .b(G812), .O(G830) );
nand2 gate286( .a(G788), .b(G812), .O(G831) );

  xor2  gate1905(.a(G815), .b(G663), .O(gate287inter0));
  nand2 gate1906(.a(gate287inter0), .b(s_194), .O(gate287inter1));
  and2  gate1907(.a(G815), .b(G663), .O(gate287inter2));
  inv1  gate1908(.a(s_194), .O(gate287inter3));
  inv1  gate1909(.a(s_195), .O(gate287inter4));
  nand2 gate1910(.a(gate287inter4), .b(gate287inter3), .O(gate287inter5));
  nor2  gate1911(.a(gate287inter5), .b(gate287inter2), .O(gate287inter6));
  inv1  gate1912(.a(G663), .O(gate287inter7));
  inv1  gate1913(.a(G815), .O(gate287inter8));
  nand2 gate1914(.a(gate287inter8), .b(gate287inter7), .O(gate287inter9));
  nand2 gate1915(.a(s_195), .b(gate287inter3), .O(gate287inter10));
  nor2  gate1916(.a(gate287inter10), .b(gate287inter9), .O(gate287inter11));
  nor2  gate1917(.a(gate287inter11), .b(gate287inter6), .O(gate287inter12));
  nand2 gate1918(.a(gate287inter12), .b(gate287inter1), .O(G832));
nand2 gate288( .a(G791), .b(G815), .O(G833) );

  xor2  gate911(.a(G819), .b(G818), .O(gate289inter0));
  nand2 gate912(.a(gate289inter0), .b(s_52), .O(gate289inter1));
  and2  gate913(.a(G819), .b(G818), .O(gate289inter2));
  inv1  gate914(.a(s_52), .O(gate289inter3));
  inv1  gate915(.a(s_53), .O(gate289inter4));
  nand2 gate916(.a(gate289inter4), .b(gate289inter3), .O(gate289inter5));
  nor2  gate917(.a(gate289inter5), .b(gate289inter2), .O(gate289inter6));
  inv1  gate918(.a(G818), .O(gate289inter7));
  inv1  gate919(.a(G819), .O(gate289inter8));
  nand2 gate920(.a(gate289inter8), .b(gate289inter7), .O(gate289inter9));
  nand2 gate921(.a(s_53), .b(gate289inter3), .O(gate289inter10));
  nor2  gate922(.a(gate289inter10), .b(gate289inter9), .O(gate289inter11));
  nor2  gate923(.a(gate289inter11), .b(gate289inter6), .O(gate289inter12));
  nand2 gate924(.a(gate289inter12), .b(gate289inter1), .O(G834));
nand2 gate290( .a(G820), .b(G821), .O(G847) );
nand2 gate291( .a(G822), .b(G823), .O(G860) );

  xor2  gate2633(.a(G825), .b(G824), .O(gate292inter0));
  nand2 gate2634(.a(gate292inter0), .b(s_298), .O(gate292inter1));
  and2  gate2635(.a(G825), .b(G824), .O(gate292inter2));
  inv1  gate2636(.a(s_298), .O(gate292inter3));
  inv1  gate2637(.a(s_299), .O(gate292inter4));
  nand2 gate2638(.a(gate292inter4), .b(gate292inter3), .O(gate292inter5));
  nor2  gate2639(.a(gate292inter5), .b(gate292inter2), .O(gate292inter6));
  inv1  gate2640(.a(G824), .O(gate292inter7));
  inv1  gate2641(.a(G825), .O(gate292inter8));
  nand2 gate2642(.a(gate292inter8), .b(gate292inter7), .O(gate292inter9));
  nand2 gate2643(.a(s_299), .b(gate292inter3), .O(gate292inter10));
  nor2  gate2644(.a(gate292inter10), .b(gate292inter9), .O(gate292inter11));
  nor2  gate2645(.a(gate292inter11), .b(gate292inter6), .O(gate292inter12));
  nand2 gate2646(.a(gate292inter12), .b(gate292inter1), .O(G873));
nand2 gate293( .a(G828), .b(G829), .O(G886) );
nand2 gate294( .a(G832), .b(G833), .O(G899) );

  xor2  gate1527(.a(G831), .b(G830), .O(gate295inter0));
  nand2 gate1528(.a(gate295inter0), .b(s_140), .O(gate295inter1));
  and2  gate1529(.a(G831), .b(G830), .O(gate295inter2));
  inv1  gate1530(.a(s_140), .O(gate295inter3));
  inv1  gate1531(.a(s_141), .O(gate295inter4));
  nand2 gate1532(.a(gate295inter4), .b(gate295inter3), .O(gate295inter5));
  nor2  gate1533(.a(gate295inter5), .b(gate295inter2), .O(gate295inter6));
  inv1  gate1534(.a(G830), .O(gate295inter7));
  inv1  gate1535(.a(G831), .O(gate295inter8));
  nand2 gate1536(.a(gate295inter8), .b(gate295inter7), .O(gate295inter9));
  nand2 gate1537(.a(s_141), .b(gate295inter3), .O(gate295inter10));
  nor2  gate1538(.a(gate295inter10), .b(gate295inter9), .O(gate295inter11));
  nor2  gate1539(.a(gate295inter11), .b(gate295inter6), .O(gate295inter12));
  nand2 gate1540(.a(gate295inter12), .b(gate295inter1), .O(G912));

  xor2  gate687(.a(G827), .b(G826), .O(gate296inter0));
  nand2 gate688(.a(gate296inter0), .b(s_20), .O(gate296inter1));
  and2  gate689(.a(G827), .b(G826), .O(gate296inter2));
  inv1  gate690(.a(s_20), .O(gate296inter3));
  inv1  gate691(.a(s_21), .O(gate296inter4));
  nand2 gate692(.a(gate296inter4), .b(gate296inter3), .O(gate296inter5));
  nor2  gate693(.a(gate296inter5), .b(gate296inter2), .O(gate296inter6));
  inv1  gate694(.a(G826), .O(gate296inter7));
  inv1  gate695(.a(G827), .O(gate296inter8));
  nand2 gate696(.a(gate296inter8), .b(gate296inter7), .O(gate296inter9));
  nand2 gate697(.a(s_21), .b(gate296inter3), .O(gate296inter10));
  nor2  gate698(.a(gate296inter10), .b(gate296inter9), .O(gate296inter11));
  nor2  gate699(.a(gate296inter11), .b(gate296inter6), .O(gate296inter12));
  nand2 gate700(.a(gate296inter12), .b(gate296inter1), .O(G925));
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );

  xor2  gate1583(.a(G1036), .b(G1), .O(gate387inter0));
  nand2 gate1584(.a(gate387inter0), .b(s_148), .O(gate387inter1));
  and2  gate1585(.a(G1036), .b(G1), .O(gate387inter2));
  inv1  gate1586(.a(s_148), .O(gate387inter3));
  inv1  gate1587(.a(s_149), .O(gate387inter4));
  nand2 gate1588(.a(gate387inter4), .b(gate387inter3), .O(gate387inter5));
  nor2  gate1589(.a(gate387inter5), .b(gate387inter2), .O(gate387inter6));
  inv1  gate1590(.a(G1), .O(gate387inter7));
  inv1  gate1591(.a(G1036), .O(gate387inter8));
  nand2 gate1592(.a(gate387inter8), .b(gate387inter7), .O(gate387inter9));
  nand2 gate1593(.a(s_149), .b(gate387inter3), .O(gate387inter10));
  nor2  gate1594(.a(gate387inter10), .b(gate387inter9), .O(gate387inter11));
  nor2  gate1595(.a(gate387inter11), .b(gate387inter6), .O(gate387inter12));
  nand2 gate1596(.a(gate387inter12), .b(gate387inter1), .O(G1132));
nand2 gate388( .a(G2), .b(G1039), .O(G1135) );
nand2 gate389( .a(G3), .b(G1042), .O(G1138) );
nand2 gate390( .a(G4), .b(G1045), .O(G1141) );

  xor2  gate1205(.a(G1048), .b(G5), .O(gate391inter0));
  nand2 gate1206(.a(gate391inter0), .b(s_94), .O(gate391inter1));
  and2  gate1207(.a(G1048), .b(G5), .O(gate391inter2));
  inv1  gate1208(.a(s_94), .O(gate391inter3));
  inv1  gate1209(.a(s_95), .O(gate391inter4));
  nand2 gate1210(.a(gate391inter4), .b(gate391inter3), .O(gate391inter5));
  nor2  gate1211(.a(gate391inter5), .b(gate391inter2), .O(gate391inter6));
  inv1  gate1212(.a(G5), .O(gate391inter7));
  inv1  gate1213(.a(G1048), .O(gate391inter8));
  nand2 gate1214(.a(gate391inter8), .b(gate391inter7), .O(gate391inter9));
  nand2 gate1215(.a(s_95), .b(gate391inter3), .O(gate391inter10));
  nor2  gate1216(.a(gate391inter10), .b(gate391inter9), .O(gate391inter11));
  nor2  gate1217(.a(gate391inter11), .b(gate391inter6), .O(gate391inter12));
  nand2 gate1218(.a(gate391inter12), .b(gate391inter1), .O(G1144));

  xor2  gate3137(.a(G1051), .b(G6), .O(gate392inter0));
  nand2 gate3138(.a(gate392inter0), .b(s_370), .O(gate392inter1));
  and2  gate3139(.a(G1051), .b(G6), .O(gate392inter2));
  inv1  gate3140(.a(s_370), .O(gate392inter3));
  inv1  gate3141(.a(s_371), .O(gate392inter4));
  nand2 gate3142(.a(gate392inter4), .b(gate392inter3), .O(gate392inter5));
  nor2  gate3143(.a(gate392inter5), .b(gate392inter2), .O(gate392inter6));
  inv1  gate3144(.a(G6), .O(gate392inter7));
  inv1  gate3145(.a(G1051), .O(gate392inter8));
  nand2 gate3146(.a(gate392inter8), .b(gate392inter7), .O(gate392inter9));
  nand2 gate3147(.a(s_371), .b(gate392inter3), .O(gate392inter10));
  nor2  gate3148(.a(gate392inter10), .b(gate392inter9), .O(gate392inter11));
  nor2  gate3149(.a(gate392inter11), .b(gate392inter6), .O(gate392inter12));
  nand2 gate3150(.a(gate392inter12), .b(gate392inter1), .O(G1147));
nand2 gate393( .a(G7), .b(G1054), .O(G1150) );

  xor2  gate2227(.a(G1057), .b(G8), .O(gate394inter0));
  nand2 gate2228(.a(gate394inter0), .b(s_240), .O(gate394inter1));
  and2  gate2229(.a(G1057), .b(G8), .O(gate394inter2));
  inv1  gate2230(.a(s_240), .O(gate394inter3));
  inv1  gate2231(.a(s_241), .O(gate394inter4));
  nand2 gate2232(.a(gate394inter4), .b(gate394inter3), .O(gate394inter5));
  nor2  gate2233(.a(gate394inter5), .b(gate394inter2), .O(gate394inter6));
  inv1  gate2234(.a(G8), .O(gate394inter7));
  inv1  gate2235(.a(G1057), .O(gate394inter8));
  nand2 gate2236(.a(gate394inter8), .b(gate394inter7), .O(gate394inter9));
  nand2 gate2237(.a(s_241), .b(gate394inter3), .O(gate394inter10));
  nor2  gate2238(.a(gate394inter10), .b(gate394inter9), .O(gate394inter11));
  nor2  gate2239(.a(gate394inter11), .b(gate394inter6), .O(gate394inter12));
  nand2 gate2240(.a(gate394inter12), .b(gate394inter1), .O(G1153));

  xor2  gate1569(.a(G1060), .b(G9), .O(gate395inter0));
  nand2 gate1570(.a(gate395inter0), .b(s_146), .O(gate395inter1));
  and2  gate1571(.a(G1060), .b(G9), .O(gate395inter2));
  inv1  gate1572(.a(s_146), .O(gate395inter3));
  inv1  gate1573(.a(s_147), .O(gate395inter4));
  nand2 gate1574(.a(gate395inter4), .b(gate395inter3), .O(gate395inter5));
  nor2  gate1575(.a(gate395inter5), .b(gate395inter2), .O(gate395inter6));
  inv1  gate1576(.a(G9), .O(gate395inter7));
  inv1  gate1577(.a(G1060), .O(gate395inter8));
  nand2 gate1578(.a(gate395inter8), .b(gate395inter7), .O(gate395inter9));
  nand2 gate1579(.a(s_147), .b(gate395inter3), .O(gate395inter10));
  nor2  gate1580(.a(gate395inter10), .b(gate395inter9), .O(gate395inter11));
  nor2  gate1581(.a(gate395inter11), .b(gate395inter6), .O(gate395inter12));
  nand2 gate1582(.a(gate395inter12), .b(gate395inter1), .O(G1156));

  xor2  gate1723(.a(G1063), .b(G10), .O(gate396inter0));
  nand2 gate1724(.a(gate396inter0), .b(s_168), .O(gate396inter1));
  and2  gate1725(.a(G1063), .b(G10), .O(gate396inter2));
  inv1  gate1726(.a(s_168), .O(gate396inter3));
  inv1  gate1727(.a(s_169), .O(gate396inter4));
  nand2 gate1728(.a(gate396inter4), .b(gate396inter3), .O(gate396inter5));
  nor2  gate1729(.a(gate396inter5), .b(gate396inter2), .O(gate396inter6));
  inv1  gate1730(.a(G10), .O(gate396inter7));
  inv1  gate1731(.a(G1063), .O(gate396inter8));
  nand2 gate1732(.a(gate396inter8), .b(gate396inter7), .O(gate396inter9));
  nand2 gate1733(.a(s_169), .b(gate396inter3), .O(gate396inter10));
  nor2  gate1734(.a(gate396inter10), .b(gate396inter9), .O(gate396inter11));
  nor2  gate1735(.a(gate396inter11), .b(gate396inter6), .O(gate396inter12));
  nand2 gate1736(.a(gate396inter12), .b(gate396inter1), .O(G1159));
nand2 gate397( .a(G11), .b(G1066), .O(G1162) );
nand2 gate398( .a(G12), .b(G1069), .O(G1165) );

  xor2  gate3123(.a(G1072), .b(G13), .O(gate399inter0));
  nand2 gate3124(.a(gate399inter0), .b(s_368), .O(gate399inter1));
  and2  gate3125(.a(G1072), .b(G13), .O(gate399inter2));
  inv1  gate3126(.a(s_368), .O(gate399inter3));
  inv1  gate3127(.a(s_369), .O(gate399inter4));
  nand2 gate3128(.a(gate399inter4), .b(gate399inter3), .O(gate399inter5));
  nor2  gate3129(.a(gate399inter5), .b(gate399inter2), .O(gate399inter6));
  inv1  gate3130(.a(G13), .O(gate399inter7));
  inv1  gate3131(.a(G1072), .O(gate399inter8));
  nand2 gate3132(.a(gate399inter8), .b(gate399inter7), .O(gate399inter9));
  nand2 gate3133(.a(s_369), .b(gate399inter3), .O(gate399inter10));
  nor2  gate3134(.a(gate399inter10), .b(gate399inter9), .O(gate399inter11));
  nor2  gate3135(.a(gate399inter11), .b(gate399inter6), .O(gate399inter12));
  nand2 gate3136(.a(gate399inter12), .b(gate399inter1), .O(G1168));

  xor2  gate2801(.a(G1075), .b(G14), .O(gate400inter0));
  nand2 gate2802(.a(gate400inter0), .b(s_322), .O(gate400inter1));
  and2  gate2803(.a(G1075), .b(G14), .O(gate400inter2));
  inv1  gate2804(.a(s_322), .O(gate400inter3));
  inv1  gate2805(.a(s_323), .O(gate400inter4));
  nand2 gate2806(.a(gate400inter4), .b(gate400inter3), .O(gate400inter5));
  nor2  gate2807(.a(gate400inter5), .b(gate400inter2), .O(gate400inter6));
  inv1  gate2808(.a(G14), .O(gate400inter7));
  inv1  gate2809(.a(G1075), .O(gate400inter8));
  nand2 gate2810(.a(gate400inter8), .b(gate400inter7), .O(gate400inter9));
  nand2 gate2811(.a(s_323), .b(gate400inter3), .O(gate400inter10));
  nor2  gate2812(.a(gate400inter10), .b(gate400inter9), .O(gate400inter11));
  nor2  gate2813(.a(gate400inter11), .b(gate400inter6), .O(gate400inter12));
  nand2 gate2814(.a(gate400inter12), .b(gate400inter1), .O(G1171));
nand2 gate401( .a(G15), .b(G1078), .O(G1174) );

  xor2  gate897(.a(G1081), .b(G16), .O(gate402inter0));
  nand2 gate898(.a(gate402inter0), .b(s_50), .O(gate402inter1));
  and2  gate899(.a(G1081), .b(G16), .O(gate402inter2));
  inv1  gate900(.a(s_50), .O(gate402inter3));
  inv1  gate901(.a(s_51), .O(gate402inter4));
  nand2 gate902(.a(gate402inter4), .b(gate402inter3), .O(gate402inter5));
  nor2  gate903(.a(gate402inter5), .b(gate402inter2), .O(gate402inter6));
  inv1  gate904(.a(G16), .O(gate402inter7));
  inv1  gate905(.a(G1081), .O(gate402inter8));
  nand2 gate906(.a(gate402inter8), .b(gate402inter7), .O(gate402inter9));
  nand2 gate907(.a(s_51), .b(gate402inter3), .O(gate402inter10));
  nor2  gate908(.a(gate402inter10), .b(gate402inter9), .O(gate402inter11));
  nor2  gate909(.a(gate402inter11), .b(gate402inter6), .O(gate402inter12));
  nand2 gate910(.a(gate402inter12), .b(gate402inter1), .O(G1177));
nand2 gate403( .a(G17), .b(G1084), .O(G1180) );

  xor2  gate2549(.a(G1087), .b(G18), .O(gate404inter0));
  nand2 gate2550(.a(gate404inter0), .b(s_286), .O(gate404inter1));
  and2  gate2551(.a(G1087), .b(G18), .O(gate404inter2));
  inv1  gate2552(.a(s_286), .O(gate404inter3));
  inv1  gate2553(.a(s_287), .O(gate404inter4));
  nand2 gate2554(.a(gate404inter4), .b(gate404inter3), .O(gate404inter5));
  nor2  gate2555(.a(gate404inter5), .b(gate404inter2), .O(gate404inter6));
  inv1  gate2556(.a(G18), .O(gate404inter7));
  inv1  gate2557(.a(G1087), .O(gate404inter8));
  nand2 gate2558(.a(gate404inter8), .b(gate404inter7), .O(gate404inter9));
  nand2 gate2559(.a(s_287), .b(gate404inter3), .O(gate404inter10));
  nor2  gate2560(.a(gate404inter10), .b(gate404inter9), .O(gate404inter11));
  nor2  gate2561(.a(gate404inter11), .b(gate404inter6), .O(gate404inter12));
  nand2 gate2562(.a(gate404inter12), .b(gate404inter1), .O(G1183));

  xor2  gate3081(.a(G1090), .b(G19), .O(gate405inter0));
  nand2 gate3082(.a(gate405inter0), .b(s_362), .O(gate405inter1));
  and2  gate3083(.a(G1090), .b(G19), .O(gate405inter2));
  inv1  gate3084(.a(s_362), .O(gate405inter3));
  inv1  gate3085(.a(s_363), .O(gate405inter4));
  nand2 gate3086(.a(gate405inter4), .b(gate405inter3), .O(gate405inter5));
  nor2  gate3087(.a(gate405inter5), .b(gate405inter2), .O(gate405inter6));
  inv1  gate3088(.a(G19), .O(gate405inter7));
  inv1  gate3089(.a(G1090), .O(gate405inter8));
  nand2 gate3090(.a(gate405inter8), .b(gate405inter7), .O(gate405inter9));
  nand2 gate3091(.a(s_363), .b(gate405inter3), .O(gate405inter10));
  nor2  gate3092(.a(gate405inter10), .b(gate405inter9), .O(gate405inter11));
  nor2  gate3093(.a(gate405inter11), .b(gate405inter6), .O(gate405inter12));
  nand2 gate3094(.a(gate405inter12), .b(gate405inter1), .O(G1186));
nand2 gate406( .a(G20), .b(G1093), .O(G1189) );

  xor2  gate757(.a(G1096), .b(G21), .O(gate407inter0));
  nand2 gate758(.a(gate407inter0), .b(s_30), .O(gate407inter1));
  and2  gate759(.a(G1096), .b(G21), .O(gate407inter2));
  inv1  gate760(.a(s_30), .O(gate407inter3));
  inv1  gate761(.a(s_31), .O(gate407inter4));
  nand2 gate762(.a(gate407inter4), .b(gate407inter3), .O(gate407inter5));
  nor2  gate763(.a(gate407inter5), .b(gate407inter2), .O(gate407inter6));
  inv1  gate764(.a(G21), .O(gate407inter7));
  inv1  gate765(.a(G1096), .O(gate407inter8));
  nand2 gate766(.a(gate407inter8), .b(gate407inter7), .O(gate407inter9));
  nand2 gate767(.a(s_31), .b(gate407inter3), .O(gate407inter10));
  nor2  gate768(.a(gate407inter10), .b(gate407inter9), .O(gate407inter11));
  nor2  gate769(.a(gate407inter11), .b(gate407inter6), .O(gate407inter12));
  nand2 gate770(.a(gate407inter12), .b(gate407inter1), .O(G1192));
nand2 gate408( .a(G22), .b(G1099), .O(G1195) );

  xor2  gate2451(.a(G1102), .b(G23), .O(gate409inter0));
  nand2 gate2452(.a(gate409inter0), .b(s_272), .O(gate409inter1));
  and2  gate2453(.a(G1102), .b(G23), .O(gate409inter2));
  inv1  gate2454(.a(s_272), .O(gate409inter3));
  inv1  gate2455(.a(s_273), .O(gate409inter4));
  nand2 gate2456(.a(gate409inter4), .b(gate409inter3), .O(gate409inter5));
  nor2  gate2457(.a(gate409inter5), .b(gate409inter2), .O(gate409inter6));
  inv1  gate2458(.a(G23), .O(gate409inter7));
  inv1  gate2459(.a(G1102), .O(gate409inter8));
  nand2 gate2460(.a(gate409inter8), .b(gate409inter7), .O(gate409inter9));
  nand2 gate2461(.a(s_273), .b(gate409inter3), .O(gate409inter10));
  nor2  gate2462(.a(gate409inter10), .b(gate409inter9), .O(gate409inter11));
  nor2  gate2463(.a(gate409inter11), .b(gate409inter6), .O(gate409inter12));
  nand2 gate2464(.a(gate409inter12), .b(gate409inter1), .O(G1198));

  xor2  gate2717(.a(G1105), .b(G24), .O(gate410inter0));
  nand2 gate2718(.a(gate410inter0), .b(s_310), .O(gate410inter1));
  and2  gate2719(.a(G1105), .b(G24), .O(gate410inter2));
  inv1  gate2720(.a(s_310), .O(gate410inter3));
  inv1  gate2721(.a(s_311), .O(gate410inter4));
  nand2 gate2722(.a(gate410inter4), .b(gate410inter3), .O(gate410inter5));
  nor2  gate2723(.a(gate410inter5), .b(gate410inter2), .O(gate410inter6));
  inv1  gate2724(.a(G24), .O(gate410inter7));
  inv1  gate2725(.a(G1105), .O(gate410inter8));
  nand2 gate2726(.a(gate410inter8), .b(gate410inter7), .O(gate410inter9));
  nand2 gate2727(.a(s_311), .b(gate410inter3), .O(gate410inter10));
  nor2  gate2728(.a(gate410inter10), .b(gate410inter9), .O(gate410inter11));
  nor2  gate2729(.a(gate410inter11), .b(gate410inter6), .O(gate410inter12));
  nand2 gate2730(.a(gate410inter12), .b(gate410inter1), .O(G1201));

  xor2  gate995(.a(G1108), .b(G25), .O(gate411inter0));
  nand2 gate996(.a(gate411inter0), .b(s_64), .O(gate411inter1));
  and2  gate997(.a(G1108), .b(G25), .O(gate411inter2));
  inv1  gate998(.a(s_64), .O(gate411inter3));
  inv1  gate999(.a(s_65), .O(gate411inter4));
  nand2 gate1000(.a(gate411inter4), .b(gate411inter3), .O(gate411inter5));
  nor2  gate1001(.a(gate411inter5), .b(gate411inter2), .O(gate411inter6));
  inv1  gate1002(.a(G25), .O(gate411inter7));
  inv1  gate1003(.a(G1108), .O(gate411inter8));
  nand2 gate1004(.a(gate411inter8), .b(gate411inter7), .O(gate411inter9));
  nand2 gate1005(.a(s_65), .b(gate411inter3), .O(gate411inter10));
  nor2  gate1006(.a(gate411inter10), .b(gate411inter9), .O(gate411inter11));
  nor2  gate1007(.a(gate411inter11), .b(gate411inter6), .O(gate411inter12));
  nand2 gate1008(.a(gate411inter12), .b(gate411inter1), .O(G1204));
nand2 gate412( .a(G26), .b(G1111), .O(G1207) );

  xor2  gate1107(.a(G1114), .b(G27), .O(gate413inter0));
  nand2 gate1108(.a(gate413inter0), .b(s_80), .O(gate413inter1));
  and2  gate1109(.a(G1114), .b(G27), .O(gate413inter2));
  inv1  gate1110(.a(s_80), .O(gate413inter3));
  inv1  gate1111(.a(s_81), .O(gate413inter4));
  nand2 gate1112(.a(gate413inter4), .b(gate413inter3), .O(gate413inter5));
  nor2  gate1113(.a(gate413inter5), .b(gate413inter2), .O(gate413inter6));
  inv1  gate1114(.a(G27), .O(gate413inter7));
  inv1  gate1115(.a(G1114), .O(gate413inter8));
  nand2 gate1116(.a(gate413inter8), .b(gate413inter7), .O(gate413inter9));
  nand2 gate1117(.a(s_81), .b(gate413inter3), .O(gate413inter10));
  nor2  gate1118(.a(gate413inter10), .b(gate413inter9), .O(gate413inter11));
  nor2  gate1119(.a(gate413inter11), .b(gate413inter6), .O(gate413inter12));
  nand2 gate1120(.a(gate413inter12), .b(gate413inter1), .O(G1210));
nand2 gate414( .a(G28), .b(G1117), .O(G1213) );

  xor2  gate1877(.a(G1120), .b(G29), .O(gate415inter0));
  nand2 gate1878(.a(gate415inter0), .b(s_190), .O(gate415inter1));
  and2  gate1879(.a(G1120), .b(G29), .O(gate415inter2));
  inv1  gate1880(.a(s_190), .O(gate415inter3));
  inv1  gate1881(.a(s_191), .O(gate415inter4));
  nand2 gate1882(.a(gate415inter4), .b(gate415inter3), .O(gate415inter5));
  nor2  gate1883(.a(gate415inter5), .b(gate415inter2), .O(gate415inter6));
  inv1  gate1884(.a(G29), .O(gate415inter7));
  inv1  gate1885(.a(G1120), .O(gate415inter8));
  nand2 gate1886(.a(gate415inter8), .b(gate415inter7), .O(gate415inter9));
  nand2 gate1887(.a(s_191), .b(gate415inter3), .O(gate415inter10));
  nor2  gate1888(.a(gate415inter10), .b(gate415inter9), .O(gate415inter11));
  nor2  gate1889(.a(gate415inter11), .b(gate415inter6), .O(gate415inter12));
  nand2 gate1890(.a(gate415inter12), .b(gate415inter1), .O(G1216));

  xor2  gate3053(.a(G1123), .b(G30), .O(gate416inter0));
  nand2 gate3054(.a(gate416inter0), .b(s_358), .O(gate416inter1));
  and2  gate3055(.a(G1123), .b(G30), .O(gate416inter2));
  inv1  gate3056(.a(s_358), .O(gate416inter3));
  inv1  gate3057(.a(s_359), .O(gate416inter4));
  nand2 gate3058(.a(gate416inter4), .b(gate416inter3), .O(gate416inter5));
  nor2  gate3059(.a(gate416inter5), .b(gate416inter2), .O(gate416inter6));
  inv1  gate3060(.a(G30), .O(gate416inter7));
  inv1  gate3061(.a(G1123), .O(gate416inter8));
  nand2 gate3062(.a(gate416inter8), .b(gate416inter7), .O(gate416inter9));
  nand2 gate3063(.a(s_359), .b(gate416inter3), .O(gate416inter10));
  nor2  gate3064(.a(gate416inter10), .b(gate416inter9), .O(gate416inter11));
  nor2  gate3065(.a(gate416inter11), .b(gate416inter6), .O(gate416inter12));
  nand2 gate3066(.a(gate416inter12), .b(gate416inter1), .O(G1219));

  xor2  gate813(.a(G1126), .b(G31), .O(gate417inter0));
  nand2 gate814(.a(gate417inter0), .b(s_38), .O(gate417inter1));
  and2  gate815(.a(G1126), .b(G31), .O(gate417inter2));
  inv1  gate816(.a(s_38), .O(gate417inter3));
  inv1  gate817(.a(s_39), .O(gate417inter4));
  nand2 gate818(.a(gate417inter4), .b(gate417inter3), .O(gate417inter5));
  nor2  gate819(.a(gate417inter5), .b(gate417inter2), .O(gate417inter6));
  inv1  gate820(.a(G31), .O(gate417inter7));
  inv1  gate821(.a(G1126), .O(gate417inter8));
  nand2 gate822(.a(gate417inter8), .b(gate417inter7), .O(gate417inter9));
  nand2 gate823(.a(s_39), .b(gate417inter3), .O(gate417inter10));
  nor2  gate824(.a(gate417inter10), .b(gate417inter9), .O(gate417inter11));
  nor2  gate825(.a(gate417inter11), .b(gate417inter6), .O(gate417inter12));
  nand2 gate826(.a(gate417inter12), .b(gate417inter1), .O(G1222));
nand2 gate418( .a(G32), .b(G1129), .O(G1225) );

  xor2  gate617(.a(G1132), .b(G1), .O(gate419inter0));
  nand2 gate618(.a(gate419inter0), .b(s_10), .O(gate419inter1));
  and2  gate619(.a(G1132), .b(G1), .O(gate419inter2));
  inv1  gate620(.a(s_10), .O(gate419inter3));
  inv1  gate621(.a(s_11), .O(gate419inter4));
  nand2 gate622(.a(gate419inter4), .b(gate419inter3), .O(gate419inter5));
  nor2  gate623(.a(gate419inter5), .b(gate419inter2), .O(gate419inter6));
  inv1  gate624(.a(G1), .O(gate419inter7));
  inv1  gate625(.a(G1132), .O(gate419inter8));
  nand2 gate626(.a(gate419inter8), .b(gate419inter7), .O(gate419inter9));
  nand2 gate627(.a(s_11), .b(gate419inter3), .O(gate419inter10));
  nor2  gate628(.a(gate419inter10), .b(gate419inter9), .O(gate419inter11));
  nor2  gate629(.a(gate419inter11), .b(gate419inter6), .O(gate419inter12));
  nand2 gate630(.a(gate419inter12), .b(gate419inter1), .O(G1228));
nand2 gate420( .a(G1036), .b(G1132), .O(G1229) );

  xor2  gate575(.a(G1135), .b(G2), .O(gate421inter0));
  nand2 gate576(.a(gate421inter0), .b(s_4), .O(gate421inter1));
  and2  gate577(.a(G1135), .b(G2), .O(gate421inter2));
  inv1  gate578(.a(s_4), .O(gate421inter3));
  inv1  gate579(.a(s_5), .O(gate421inter4));
  nand2 gate580(.a(gate421inter4), .b(gate421inter3), .O(gate421inter5));
  nor2  gate581(.a(gate421inter5), .b(gate421inter2), .O(gate421inter6));
  inv1  gate582(.a(G2), .O(gate421inter7));
  inv1  gate583(.a(G1135), .O(gate421inter8));
  nand2 gate584(.a(gate421inter8), .b(gate421inter7), .O(gate421inter9));
  nand2 gate585(.a(s_5), .b(gate421inter3), .O(gate421inter10));
  nor2  gate586(.a(gate421inter10), .b(gate421inter9), .O(gate421inter11));
  nor2  gate587(.a(gate421inter11), .b(gate421inter6), .O(gate421inter12));
  nand2 gate588(.a(gate421inter12), .b(gate421inter1), .O(G1230));

  xor2  gate2941(.a(G1135), .b(G1039), .O(gate422inter0));
  nand2 gate2942(.a(gate422inter0), .b(s_342), .O(gate422inter1));
  and2  gate2943(.a(G1135), .b(G1039), .O(gate422inter2));
  inv1  gate2944(.a(s_342), .O(gate422inter3));
  inv1  gate2945(.a(s_343), .O(gate422inter4));
  nand2 gate2946(.a(gate422inter4), .b(gate422inter3), .O(gate422inter5));
  nor2  gate2947(.a(gate422inter5), .b(gate422inter2), .O(gate422inter6));
  inv1  gate2948(.a(G1039), .O(gate422inter7));
  inv1  gate2949(.a(G1135), .O(gate422inter8));
  nand2 gate2950(.a(gate422inter8), .b(gate422inter7), .O(gate422inter9));
  nand2 gate2951(.a(s_343), .b(gate422inter3), .O(gate422inter10));
  nor2  gate2952(.a(gate422inter10), .b(gate422inter9), .O(gate422inter11));
  nor2  gate2953(.a(gate422inter11), .b(gate422inter6), .O(gate422inter12));
  nand2 gate2954(.a(gate422inter12), .b(gate422inter1), .O(G1231));
nand2 gate423( .a(G3), .b(G1138), .O(G1232) );
nand2 gate424( .a(G1042), .b(G1138), .O(G1233) );

  xor2  gate1219(.a(G1141), .b(G4), .O(gate425inter0));
  nand2 gate1220(.a(gate425inter0), .b(s_96), .O(gate425inter1));
  and2  gate1221(.a(G1141), .b(G4), .O(gate425inter2));
  inv1  gate1222(.a(s_96), .O(gate425inter3));
  inv1  gate1223(.a(s_97), .O(gate425inter4));
  nand2 gate1224(.a(gate425inter4), .b(gate425inter3), .O(gate425inter5));
  nor2  gate1225(.a(gate425inter5), .b(gate425inter2), .O(gate425inter6));
  inv1  gate1226(.a(G4), .O(gate425inter7));
  inv1  gate1227(.a(G1141), .O(gate425inter8));
  nand2 gate1228(.a(gate425inter8), .b(gate425inter7), .O(gate425inter9));
  nand2 gate1229(.a(s_97), .b(gate425inter3), .O(gate425inter10));
  nor2  gate1230(.a(gate425inter10), .b(gate425inter9), .O(gate425inter11));
  nor2  gate1231(.a(gate425inter11), .b(gate425inter6), .O(gate425inter12));
  nand2 gate1232(.a(gate425inter12), .b(gate425inter1), .O(G1234));

  xor2  gate2185(.a(G1141), .b(G1045), .O(gate426inter0));
  nand2 gate2186(.a(gate426inter0), .b(s_234), .O(gate426inter1));
  and2  gate2187(.a(G1141), .b(G1045), .O(gate426inter2));
  inv1  gate2188(.a(s_234), .O(gate426inter3));
  inv1  gate2189(.a(s_235), .O(gate426inter4));
  nand2 gate2190(.a(gate426inter4), .b(gate426inter3), .O(gate426inter5));
  nor2  gate2191(.a(gate426inter5), .b(gate426inter2), .O(gate426inter6));
  inv1  gate2192(.a(G1045), .O(gate426inter7));
  inv1  gate2193(.a(G1141), .O(gate426inter8));
  nand2 gate2194(.a(gate426inter8), .b(gate426inter7), .O(gate426inter9));
  nand2 gate2195(.a(s_235), .b(gate426inter3), .O(gate426inter10));
  nor2  gate2196(.a(gate426inter10), .b(gate426inter9), .O(gate426inter11));
  nor2  gate2197(.a(gate426inter11), .b(gate426inter6), .O(gate426inter12));
  nand2 gate2198(.a(gate426inter12), .b(gate426inter1), .O(G1235));
nand2 gate427( .a(G5), .b(G1144), .O(G1236) );

  xor2  gate589(.a(G1144), .b(G1048), .O(gate428inter0));
  nand2 gate590(.a(gate428inter0), .b(s_6), .O(gate428inter1));
  and2  gate591(.a(G1144), .b(G1048), .O(gate428inter2));
  inv1  gate592(.a(s_6), .O(gate428inter3));
  inv1  gate593(.a(s_7), .O(gate428inter4));
  nand2 gate594(.a(gate428inter4), .b(gate428inter3), .O(gate428inter5));
  nor2  gate595(.a(gate428inter5), .b(gate428inter2), .O(gate428inter6));
  inv1  gate596(.a(G1048), .O(gate428inter7));
  inv1  gate597(.a(G1144), .O(gate428inter8));
  nand2 gate598(.a(gate428inter8), .b(gate428inter7), .O(gate428inter9));
  nand2 gate599(.a(s_7), .b(gate428inter3), .O(gate428inter10));
  nor2  gate600(.a(gate428inter10), .b(gate428inter9), .O(gate428inter11));
  nor2  gate601(.a(gate428inter11), .b(gate428inter6), .O(gate428inter12));
  nand2 gate602(.a(gate428inter12), .b(gate428inter1), .O(G1237));
nand2 gate429( .a(G6), .b(G1147), .O(G1238) );

  xor2  gate2563(.a(G1147), .b(G1051), .O(gate430inter0));
  nand2 gate2564(.a(gate430inter0), .b(s_288), .O(gate430inter1));
  and2  gate2565(.a(G1147), .b(G1051), .O(gate430inter2));
  inv1  gate2566(.a(s_288), .O(gate430inter3));
  inv1  gate2567(.a(s_289), .O(gate430inter4));
  nand2 gate2568(.a(gate430inter4), .b(gate430inter3), .O(gate430inter5));
  nor2  gate2569(.a(gate430inter5), .b(gate430inter2), .O(gate430inter6));
  inv1  gate2570(.a(G1051), .O(gate430inter7));
  inv1  gate2571(.a(G1147), .O(gate430inter8));
  nand2 gate2572(.a(gate430inter8), .b(gate430inter7), .O(gate430inter9));
  nand2 gate2573(.a(s_289), .b(gate430inter3), .O(gate430inter10));
  nor2  gate2574(.a(gate430inter10), .b(gate430inter9), .O(gate430inter11));
  nor2  gate2575(.a(gate430inter11), .b(gate430inter6), .O(gate430inter12));
  nand2 gate2576(.a(gate430inter12), .b(gate430inter1), .O(G1239));
nand2 gate431( .a(G7), .b(G1150), .O(G1240) );
nand2 gate432( .a(G1054), .b(G1150), .O(G1241) );

  xor2  gate1667(.a(G1153), .b(G8), .O(gate433inter0));
  nand2 gate1668(.a(gate433inter0), .b(s_160), .O(gate433inter1));
  and2  gate1669(.a(G1153), .b(G8), .O(gate433inter2));
  inv1  gate1670(.a(s_160), .O(gate433inter3));
  inv1  gate1671(.a(s_161), .O(gate433inter4));
  nand2 gate1672(.a(gate433inter4), .b(gate433inter3), .O(gate433inter5));
  nor2  gate1673(.a(gate433inter5), .b(gate433inter2), .O(gate433inter6));
  inv1  gate1674(.a(G8), .O(gate433inter7));
  inv1  gate1675(.a(G1153), .O(gate433inter8));
  nand2 gate1676(.a(gate433inter8), .b(gate433inter7), .O(gate433inter9));
  nand2 gate1677(.a(s_161), .b(gate433inter3), .O(gate433inter10));
  nor2  gate1678(.a(gate433inter10), .b(gate433inter9), .O(gate433inter11));
  nor2  gate1679(.a(gate433inter11), .b(gate433inter6), .O(gate433inter12));
  nand2 gate1680(.a(gate433inter12), .b(gate433inter1), .O(G1242));

  xor2  gate1415(.a(G1153), .b(G1057), .O(gate434inter0));
  nand2 gate1416(.a(gate434inter0), .b(s_124), .O(gate434inter1));
  and2  gate1417(.a(G1153), .b(G1057), .O(gate434inter2));
  inv1  gate1418(.a(s_124), .O(gate434inter3));
  inv1  gate1419(.a(s_125), .O(gate434inter4));
  nand2 gate1420(.a(gate434inter4), .b(gate434inter3), .O(gate434inter5));
  nor2  gate1421(.a(gate434inter5), .b(gate434inter2), .O(gate434inter6));
  inv1  gate1422(.a(G1057), .O(gate434inter7));
  inv1  gate1423(.a(G1153), .O(gate434inter8));
  nand2 gate1424(.a(gate434inter8), .b(gate434inter7), .O(gate434inter9));
  nand2 gate1425(.a(s_125), .b(gate434inter3), .O(gate434inter10));
  nor2  gate1426(.a(gate434inter10), .b(gate434inter9), .O(gate434inter11));
  nor2  gate1427(.a(gate434inter11), .b(gate434inter6), .O(gate434inter12));
  nand2 gate1428(.a(gate434inter12), .b(gate434inter1), .O(G1243));

  xor2  gate2437(.a(G1156), .b(G9), .O(gate435inter0));
  nand2 gate2438(.a(gate435inter0), .b(s_270), .O(gate435inter1));
  and2  gate2439(.a(G1156), .b(G9), .O(gate435inter2));
  inv1  gate2440(.a(s_270), .O(gate435inter3));
  inv1  gate2441(.a(s_271), .O(gate435inter4));
  nand2 gate2442(.a(gate435inter4), .b(gate435inter3), .O(gate435inter5));
  nor2  gate2443(.a(gate435inter5), .b(gate435inter2), .O(gate435inter6));
  inv1  gate2444(.a(G9), .O(gate435inter7));
  inv1  gate2445(.a(G1156), .O(gate435inter8));
  nand2 gate2446(.a(gate435inter8), .b(gate435inter7), .O(gate435inter9));
  nand2 gate2447(.a(s_271), .b(gate435inter3), .O(gate435inter10));
  nor2  gate2448(.a(gate435inter10), .b(gate435inter9), .O(gate435inter11));
  nor2  gate2449(.a(gate435inter11), .b(gate435inter6), .O(gate435inter12));
  nand2 gate2450(.a(gate435inter12), .b(gate435inter1), .O(G1244));
nand2 gate436( .a(G1060), .b(G1156), .O(G1245) );
nand2 gate437( .a(G10), .b(G1159), .O(G1246) );

  xor2  gate3221(.a(G1159), .b(G1063), .O(gate438inter0));
  nand2 gate3222(.a(gate438inter0), .b(s_382), .O(gate438inter1));
  and2  gate3223(.a(G1159), .b(G1063), .O(gate438inter2));
  inv1  gate3224(.a(s_382), .O(gate438inter3));
  inv1  gate3225(.a(s_383), .O(gate438inter4));
  nand2 gate3226(.a(gate438inter4), .b(gate438inter3), .O(gate438inter5));
  nor2  gate3227(.a(gate438inter5), .b(gate438inter2), .O(gate438inter6));
  inv1  gate3228(.a(G1063), .O(gate438inter7));
  inv1  gate3229(.a(G1159), .O(gate438inter8));
  nand2 gate3230(.a(gate438inter8), .b(gate438inter7), .O(gate438inter9));
  nand2 gate3231(.a(s_383), .b(gate438inter3), .O(gate438inter10));
  nor2  gate3232(.a(gate438inter10), .b(gate438inter9), .O(gate438inter11));
  nor2  gate3233(.a(gate438inter11), .b(gate438inter6), .O(gate438inter12));
  nand2 gate3234(.a(gate438inter12), .b(gate438inter1), .O(G1247));
nand2 gate439( .a(G11), .b(G1162), .O(G1248) );
nand2 gate440( .a(G1066), .b(G1162), .O(G1249) );

  xor2  gate659(.a(G1165), .b(G12), .O(gate441inter0));
  nand2 gate660(.a(gate441inter0), .b(s_16), .O(gate441inter1));
  and2  gate661(.a(G1165), .b(G12), .O(gate441inter2));
  inv1  gate662(.a(s_16), .O(gate441inter3));
  inv1  gate663(.a(s_17), .O(gate441inter4));
  nand2 gate664(.a(gate441inter4), .b(gate441inter3), .O(gate441inter5));
  nor2  gate665(.a(gate441inter5), .b(gate441inter2), .O(gate441inter6));
  inv1  gate666(.a(G12), .O(gate441inter7));
  inv1  gate667(.a(G1165), .O(gate441inter8));
  nand2 gate668(.a(gate441inter8), .b(gate441inter7), .O(gate441inter9));
  nand2 gate669(.a(s_17), .b(gate441inter3), .O(gate441inter10));
  nor2  gate670(.a(gate441inter10), .b(gate441inter9), .O(gate441inter11));
  nor2  gate671(.a(gate441inter11), .b(gate441inter6), .O(gate441inter12));
  nand2 gate672(.a(gate441inter12), .b(gate441inter1), .O(G1250));
nand2 gate442( .a(G1069), .b(G1165), .O(G1251) );

  xor2  gate561(.a(G1168), .b(G13), .O(gate443inter0));
  nand2 gate562(.a(gate443inter0), .b(s_2), .O(gate443inter1));
  and2  gate563(.a(G1168), .b(G13), .O(gate443inter2));
  inv1  gate564(.a(s_2), .O(gate443inter3));
  inv1  gate565(.a(s_3), .O(gate443inter4));
  nand2 gate566(.a(gate443inter4), .b(gate443inter3), .O(gate443inter5));
  nor2  gate567(.a(gate443inter5), .b(gate443inter2), .O(gate443inter6));
  inv1  gate568(.a(G13), .O(gate443inter7));
  inv1  gate569(.a(G1168), .O(gate443inter8));
  nand2 gate570(.a(gate443inter8), .b(gate443inter7), .O(gate443inter9));
  nand2 gate571(.a(s_3), .b(gate443inter3), .O(gate443inter10));
  nor2  gate572(.a(gate443inter10), .b(gate443inter9), .O(gate443inter11));
  nor2  gate573(.a(gate443inter11), .b(gate443inter6), .O(gate443inter12));
  nand2 gate574(.a(gate443inter12), .b(gate443inter1), .O(G1252));

  xor2  gate2465(.a(G1168), .b(G1072), .O(gate444inter0));
  nand2 gate2466(.a(gate444inter0), .b(s_274), .O(gate444inter1));
  and2  gate2467(.a(G1168), .b(G1072), .O(gate444inter2));
  inv1  gate2468(.a(s_274), .O(gate444inter3));
  inv1  gate2469(.a(s_275), .O(gate444inter4));
  nand2 gate2470(.a(gate444inter4), .b(gate444inter3), .O(gate444inter5));
  nor2  gate2471(.a(gate444inter5), .b(gate444inter2), .O(gate444inter6));
  inv1  gate2472(.a(G1072), .O(gate444inter7));
  inv1  gate2473(.a(G1168), .O(gate444inter8));
  nand2 gate2474(.a(gate444inter8), .b(gate444inter7), .O(gate444inter9));
  nand2 gate2475(.a(s_275), .b(gate444inter3), .O(gate444inter10));
  nor2  gate2476(.a(gate444inter10), .b(gate444inter9), .O(gate444inter11));
  nor2  gate2477(.a(gate444inter11), .b(gate444inter6), .O(gate444inter12));
  nand2 gate2478(.a(gate444inter12), .b(gate444inter1), .O(G1253));

  xor2  gate1793(.a(G1171), .b(G14), .O(gate445inter0));
  nand2 gate1794(.a(gate445inter0), .b(s_178), .O(gate445inter1));
  and2  gate1795(.a(G1171), .b(G14), .O(gate445inter2));
  inv1  gate1796(.a(s_178), .O(gate445inter3));
  inv1  gate1797(.a(s_179), .O(gate445inter4));
  nand2 gate1798(.a(gate445inter4), .b(gate445inter3), .O(gate445inter5));
  nor2  gate1799(.a(gate445inter5), .b(gate445inter2), .O(gate445inter6));
  inv1  gate1800(.a(G14), .O(gate445inter7));
  inv1  gate1801(.a(G1171), .O(gate445inter8));
  nand2 gate1802(.a(gate445inter8), .b(gate445inter7), .O(gate445inter9));
  nand2 gate1803(.a(s_179), .b(gate445inter3), .O(gate445inter10));
  nor2  gate1804(.a(gate445inter10), .b(gate445inter9), .O(gate445inter11));
  nor2  gate1805(.a(gate445inter11), .b(gate445inter6), .O(gate445inter12));
  nand2 gate1806(.a(gate445inter12), .b(gate445inter1), .O(G1254));

  xor2  gate2899(.a(G1171), .b(G1075), .O(gate446inter0));
  nand2 gate2900(.a(gate446inter0), .b(s_336), .O(gate446inter1));
  and2  gate2901(.a(G1171), .b(G1075), .O(gate446inter2));
  inv1  gate2902(.a(s_336), .O(gate446inter3));
  inv1  gate2903(.a(s_337), .O(gate446inter4));
  nand2 gate2904(.a(gate446inter4), .b(gate446inter3), .O(gate446inter5));
  nor2  gate2905(.a(gate446inter5), .b(gate446inter2), .O(gate446inter6));
  inv1  gate2906(.a(G1075), .O(gate446inter7));
  inv1  gate2907(.a(G1171), .O(gate446inter8));
  nand2 gate2908(.a(gate446inter8), .b(gate446inter7), .O(gate446inter9));
  nand2 gate2909(.a(s_337), .b(gate446inter3), .O(gate446inter10));
  nor2  gate2910(.a(gate446inter10), .b(gate446inter9), .O(gate446inter11));
  nor2  gate2911(.a(gate446inter11), .b(gate446inter6), .O(gate446inter12));
  nand2 gate2912(.a(gate446inter12), .b(gate446inter1), .O(G1255));

  xor2  gate2997(.a(G1174), .b(G15), .O(gate447inter0));
  nand2 gate2998(.a(gate447inter0), .b(s_350), .O(gate447inter1));
  and2  gate2999(.a(G1174), .b(G15), .O(gate447inter2));
  inv1  gate3000(.a(s_350), .O(gate447inter3));
  inv1  gate3001(.a(s_351), .O(gate447inter4));
  nand2 gate3002(.a(gate447inter4), .b(gate447inter3), .O(gate447inter5));
  nor2  gate3003(.a(gate447inter5), .b(gate447inter2), .O(gate447inter6));
  inv1  gate3004(.a(G15), .O(gate447inter7));
  inv1  gate3005(.a(G1174), .O(gate447inter8));
  nand2 gate3006(.a(gate447inter8), .b(gate447inter7), .O(gate447inter9));
  nand2 gate3007(.a(s_351), .b(gate447inter3), .O(gate447inter10));
  nor2  gate3008(.a(gate447inter10), .b(gate447inter9), .O(gate447inter11));
  nor2  gate3009(.a(gate447inter11), .b(gate447inter6), .O(gate447inter12));
  nand2 gate3010(.a(gate447inter12), .b(gate447inter1), .O(G1256));
nand2 gate448( .a(G1078), .b(G1174), .O(G1257) );

  xor2  gate2675(.a(G1177), .b(G16), .O(gate449inter0));
  nand2 gate2676(.a(gate449inter0), .b(s_304), .O(gate449inter1));
  and2  gate2677(.a(G1177), .b(G16), .O(gate449inter2));
  inv1  gate2678(.a(s_304), .O(gate449inter3));
  inv1  gate2679(.a(s_305), .O(gate449inter4));
  nand2 gate2680(.a(gate449inter4), .b(gate449inter3), .O(gate449inter5));
  nor2  gate2681(.a(gate449inter5), .b(gate449inter2), .O(gate449inter6));
  inv1  gate2682(.a(G16), .O(gate449inter7));
  inv1  gate2683(.a(G1177), .O(gate449inter8));
  nand2 gate2684(.a(gate449inter8), .b(gate449inter7), .O(gate449inter9));
  nand2 gate2685(.a(s_305), .b(gate449inter3), .O(gate449inter10));
  nor2  gate2686(.a(gate449inter10), .b(gate449inter9), .O(gate449inter11));
  nor2  gate2687(.a(gate449inter11), .b(gate449inter6), .O(gate449inter12));
  nand2 gate2688(.a(gate449inter12), .b(gate449inter1), .O(G1258));
nand2 gate450( .a(G1081), .b(G1177), .O(G1259) );
nand2 gate451( .a(G17), .b(G1180), .O(G1260) );
nand2 gate452( .a(G1084), .b(G1180), .O(G1261) );

  xor2  gate2101(.a(G1183), .b(G18), .O(gate453inter0));
  nand2 gate2102(.a(gate453inter0), .b(s_222), .O(gate453inter1));
  and2  gate2103(.a(G1183), .b(G18), .O(gate453inter2));
  inv1  gate2104(.a(s_222), .O(gate453inter3));
  inv1  gate2105(.a(s_223), .O(gate453inter4));
  nand2 gate2106(.a(gate453inter4), .b(gate453inter3), .O(gate453inter5));
  nor2  gate2107(.a(gate453inter5), .b(gate453inter2), .O(gate453inter6));
  inv1  gate2108(.a(G18), .O(gate453inter7));
  inv1  gate2109(.a(G1183), .O(gate453inter8));
  nand2 gate2110(.a(gate453inter8), .b(gate453inter7), .O(gate453inter9));
  nand2 gate2111(.a(s_223), .b(gate453inter3), .O(gate453inter10));
  nor2  gate2112(.a(gate453inter10), .b(gate453inter9), .O(gate453inter11));
  nor2  gate2113(.a(gate453inter11), .b(gate453inter6), .O(gate453inter12));
  nand2 gate2114(.a(gate453inter12), .b(gate453inter1), .O(G1262));
nand2 gate454( .a(G1087), .b(G1183), .O(G1263) );
nand2 gate455( .a(G19), .b(G1186), .O(G1264) );
nand2 gate456( .a(G1090), .b(G1186), .O(G1265) );

  xor2  gate1499(.a(G1189), .b(G20), .O(gate457inter0));
  nand2 gate1500(.a(gate457inter0), .b(s_136), .O(gate457inter1));
  and2  gate1501(.a(G1189), .b(G20), .O(gate457inter2));
  inv1  gate1502(.a(s_136), .O(gate457inter3));
  inv1  gate1503(.a(s_137), .O(gate457inter4));
  nand2 gate1504(.a(gate457inter4), .b(gate457inter3), .O(gate457inter5));
  nor2  gate1505(.a(gate457inter5), .b(gate457inter2), .O(gate457inter6));
  inv1  gate1506(.a(G20), .O(gate457inter7));
  inv1  gate1507(.a(G1189), .O(gate457inter8));
  nand2 gate1508(.a(gate457inter8), .b(gate457inter7), .O(gate457inter9));
  nand2 gate1509(.a(s_137), .b(gate457inter3), .O(gate457inter10));
  nor2  gate1510(.a(gate457inter10), .b(gate457inter9), .O(gate457inter11));
  nor2  gate1511(.a(gate457inter11), .b(gate457inter6), .O(gate457inter12));
  nand2 gate1512(.a(gate457inter12), .b(gate457inter1), .O(G1266));

  xor2  gate981(.a(G1189), .b(G1093), .O(gate458inter0));
  nand2 gate982(.a(gate458inter0), .b(s_62), .O(gate458inter1));
  and2  gate983(.a(G1189), .b(G1093), .O(gate458inter2));
  inv1  gate984(.a(s_62), .O(gate458inter3));
  inv1  gate985(.a(s_63), .O(gate458inter4));
  nand2 gate986(.a(gate458inter4), .b(gate458inter3), .O(gate458inter5));
  nor2  gate987(.a(gate458inter5), .b(gate458inter2), .O(gate458inter6));
  inv1  gate988(.a(G1093), .O(gate458inter7));
  inv1  gate989(.a(G1189), .O(gate458inter8));
  nand2 gate990(.a(gate458inter8), .b(gate458inter7), .O(gate458inter9));
  nand2 gate991(.a(s_63), .b(gate458inter3), .O(gate458inter10));
  nor2  gate992(.a(gate458inter10), .b(gate458inter9), .O(gate458inter11));
  nor2  gate993(.a(gate458inter11), .b(gate458inter6), .O(gate458inter12));
  nand2 gate994(.a(gate458inter12), .b(gate458inter1), .O(G1267));

  xor2  gate827(.a(G1192), .b(G21), .O(gate459inter0));
  nand2 gate828(.a(gate459inter0), .b(s_40), .O(gate459inter1));
  and2  gate829(.a(G1192), .b(G21), .O(gate459inter2));
  inv1  gate830(.a(s_40), .O(gate459inter3));
  inv1  gate831(.a(s_41), .O(gate459inter4));
  nand2 gate832(.a(gate459inter4), .b(gate459inter3), .O(gate459inter5));
  nor2  gate833(.a(gate459inter5), .b(gate459inter2), .O(gate459inter6));
  inv1  gate834(.a(G21), .O(gate459inter7));
  inv1  gate835(.a(G1192), .O(gate459inter8));
  nand2 gate836(.a(gate459inter8), .b(gate459inter7), .O(gate459inter9));
  nand2 gate837(.a(s_41), .b(gate459inter3), .O(gate459inter10));
  nor2  gate838(.a(gate459inter10), .b(gate459inter9), .O(gate459inter11));
  nor2  gate839(.a(gate459inter11), .b(gate459inter6), .O(gate459inter12));
  nand2 gate840(.a(gate459inter12), .b(gate459inter1), .O(G1268));

  xor2  gate1163(.a(G1192), .b(G1096), .O(gate460inter0));
  nand2 gate1164(.a(gate460inter0), .b(s_88), .O(gate460inter1));
  and2  gate1165(.a(G1192), .b(G1096), .O(gate460inter2));
  inv1  gate1166(.a(s_88), .O(gate460inter3));
  inv1  gate1167(.a(s_89), .O(gate460inter4));
  nand2 gate1168(.a(gate460inter4), .b(gate460inter3), .O(gate460inter5));
  nor2  gate1169(.a(gate460inter5), .b(gate460inter2), .O(gate460inter6));
  inv1  gate1170(.a(G1096), .O(gate460inter7));
  inv1  gate1171(.a(G1192), .O(gate460inter8));
  nand2 gate1172(.a(gate460inter8), .b(gate460inter7), .O(gate460inter9));
  nand2 gate1173(.a(s_89), .b(gate460inter3), .O(gate460inter10));
  nor2  gate1174(.a(gate460inter10), .b(gate460inter9), .O(gate460inter11));
  nor2  gate1175(.a(gate460inter11), .b(gate460inter6), .O(gate460inter12));
  nand2 gate1176(.a(gate460inter12), .b(gate460inter1), .O(G1269));

  xor2  gate2871(.a(G1195), .b(G22), .O(gate461inter0));
  nand2 gate2872(.a(gate461inter0), .b(s_332), .O(gate461inter1));
  and2  gate2873(.a(G1195), .b(G22), .O(gate461inter2));
  inv1  gate2874(.a(s_332), .O(gate461inter3));
  inv1  gate2875(.a(s_333), .O(gate461inter4));
  nand2 gate2876(.a(gate461inter4), .b(gate461inter3), .O(gate461inter5));
  nor2  gate2877(.a(gate461inter5), .b(gate461inter2), .O(gate461inter6));
  inv1  gate2878(.a(G22), .O(gate461inter7));
  inv1  gate2879(.a(G1195), .O(gate461inter8));
  nand2 gate2880(.a(gate461inter8), .b(gate461inter7), .O(gate461inter9));
  nand2 gate2881(.a(s_333), .b(gate461inter3), .O(gate461inter10));
  nor2  gate2882(.a(gate461inter10), .b(gate461inter9), .O(gate461inter11));
  nor2  gate2883(.a(gate461inter11), .b(gate461inter6), .O(gate461inter12));
  nand2 gate2884(.a(gate461inter12), .b(gate461inter1), .O(G1270));

  xor2  gate1989(.a(G1195), .b(G1099), .O(gate462inter0));
  nand2 gate1990(.a(gate462inter0), .b(s_206), .O(gate462inter1));
  and2  gate1991(.a(G1195), .b(G1099), .O(gate462inter2));
  inv1  gate1992(.a(s_206), .O(gate462inter3));
  inv1  gate1993(.a(s_207), .O(gate462inter4));
  nand2 gate1994(.a(gate462inter4), .b(gate462inter3), .O(gate462inter5));
  nor2  gate1995(.a(gate462inter5), .b(gate462inter2), .O(gate462inter6));
  inv1  gate1996(.a(G1099), .O(gate462inter7));
  inv1  gate1997(.a(G1195), .O(gate462inter8));
  nand2 gate1998(.a(gate462inter8), .b(gate462inter7), .O(gate462inter9));
  nand2 gate1999(.a(s_207), .b(gate462inter3), .O(gate462inter10));
  nor2  gate2000(.a(gate462inter10), .b(gate462inter9), .O(gate462inter11));
  nor2  gate2001(.a(gate462inter11), .b(gate462inter6), .O(gate462inter12));
  nand2 gate2002(.a(gate462inter12), .b(gate462inter1), .O(G1271));

  xor2  gate2843(.a(G1198), .b(G23), .O(gate463inter0));
  nand2 gate2844(.a(gate463inter0), .b(s_328), .O(gate463inter1));
  and2  gate2845(.a(G1198), .b(G23), .O(gate463inter2));
  inv1  gate2846(.a(s_328), .O(gate463inter3));
  inv1  gate2847(.a(s_329), .O(gate463inter4));
  nand2 gate2848(.a(gate463inter4), .b(gate463inter3), .O(gate463inter5));
  nor2  gate2849(.a(gate463inter5), .b(gate463inter2), .O(gate463inter6));
  inv1  gate2850(.a(G23), .O(gate463inter7));
  inv1  gate2851(.a(G1198), .O(gate463inter8));
  nand2 gate2852(.a(gate463inter8), .b(gate463inter7), .O(gate463inter9));
  nand2 gate2853(.a(s_329), .b(gate463inter3), .O(gate463inter10));
  nor2  gate2854(.a(gate463inter10), .b(gate463inter9), .O(gate463inter11));
  nor2  gate2855(.a(gate463inter11), .b(gate463inter6), .O(gate463inter12));
  nand2 gate2856(.a(gate463inter12), .b(gate463inter1), .O(G1272));
nand2 gate464( .a(G1102), .b(G1198), .O(G1273) );
nand2 gate465( .a(G24), .b(G1201), .O(G1274) );
nand2 gate466( .a(G1105), .b(G1201), .O(G1275) );

  xor2  gate2339(.a(G1204), .b(G25), .O(gate467inter0));
  nand2 gate2340(.a(gate467inter0), .b(s_256), .O(gate467inter1));
  and2  gate2341(.a(G1204), .b(G25), .O(gate467inter2));
  inv1  gate2342(.a(s_256), .O(gate467inter3));
  inv1  gate2343(.a(s_257), .O(gate467inter4));
  nand2 gate2344(.a(gate467inter4), .b(gate467inter3), .O(gate467inter5));
  nor2  gate2345(.a(gate467inter5), .b(gate467inter2), .O(gate467inter6));
  inv1  gate2346(.a(G25), .O(gate467inter7));
  inv1  gate2347(.a(G1204), .O(gate467inter8));
  nand2 gate2348(.a(gate467inter8), .b(gate467inter7), .O(gate467inter9));
  nand2 gate2349(.a(s_257), .b(gate467inter3), .O(gate467inter10));
  nor2  gate2350(.a(gate467inter10), .b(gate467inter9), .O(gate467inter11));
  nor2  gate2351(.a(gate467inter11), .b(gate467inter6), .O(gate467inter12));
  nand2 gate2352(.a(gate467inter12), .b(gate467inter1), .O(G1276));

  xor2  gate3193(.a(G1204), .b(G1108), .O(gate468inter0));
  nand2 gate3194(.a(gate468inter0), .b(s_378), .O(gate468inter1));
  and2  gate3195(.a(G1204), .b(G1108), .O(gate468inter2));
  inv1  gate3196(.a(s_378), .O(gate468inter3));
  inv1  gate3197(.a(s_379), .O(gate468inter4));
  nand2 gate3198(.a(gate468inter4), .b(gate468inter3), .O(gate468inter5));
  nor2  gate3199(.a(gate468inter5), .b(gate468inter2), .O(gate468inter6));
  inv1  gate3200(.a(G1108), .O(gate468inter7));
  inv1  gate3201(.a(G1204), .O(gate468inter8));
  nand2 gate3202(.a(gate468inter8), .b(gate468inter7), .O(gate468inter9));
  nand2 gate3203(.a(s_379), .b(gate468inter3), .O(gate468inter10));
  nor2  gate3204(.a(gate468inter10), .b(gate468inter9), .O(gate468inter11));
  nor2  gate3205(.a(gate468inter11), .b(gate468inter6), .O(gate468inter12));
  nand2 gate3206(.a(gate468inter12), .b(gate468inter1), .O(G1277));
nand2 gate469( .a(G26), .b(G1207), .O(G1278) );

  xor2  gate743(.a(G1207), .b(G1111), .O(gate470inter0));
  nand2 gate744(.a(gate470inter0), .b(s_28), .O(gate470inter1));
  and2  gate745(.a(G1207), .b(G1111), .O(gate470inter2));
  inv1  gate746(.a(s_28), .O(gate470inter3));
  inv1  gate747(.a(s_29), .O(gate470inter4));
  nand2 gate748(.a(gate470inter4), .b(gate470inter3), .O(gate470inter5));
  nor2  gate749(.a(gate470inter5), .b(gate470inter2), .O(gate470inter6));
  inv1  gate750(.a(G1111), .O(gate470inter7));
  inv1  gate751(.a(G1207), .O(gate470inter8));
  nand2 gate752(.a(gate470inter8), .b(gate470inter7), .O(gate470inter9));
  nand2 gate753(.a(s_29), .b(gate470inter3), .O(gate470inter10));
  nor2  gate754(.a(gate470inter10), .b(gate470inter9), .O(gate470inter11));
  nor2  gate755(.a(gate470inter11), .b(gate470inter6), .O(gate470inter12));
  nand2 gate756(.a(gate470inter12), .b(gate470inter1), .O(G1279));
nand2 gate471( .a(G27), .b(G1210), .O(G1280) );
nand2 gate472( .a(G1114), .b(G1210), .O(G1281) );

  xor2  gate925(.a(G1213), .b(G28), .O(gate473inter0));
  nand2 gate926(.a(gate473inter0), .b(s_54), .O(gate473inter1));
  and2  gate927(.a(G1213), .b(G28), .O(gate473inter2));
  inv1  gate928(.a(s_54), .O(gate473inter3));
  inv1  gate929(.a(s_55), .O(gate473inter4));
  nand2 gate930(.a(gate473inter4), .b(gate473inter3), .O(gate473inter5));
  nor2  gate931(.a(gate473inter5), .b(gate473inter2), .O(gate473inter6));
  inv1  gate932(.a(G28), .O(gate473inter7));
  inv1  gate933(.a(G1213), .O(gate473inter8));
  nand2 gate934(.a(gate473inter8), .b(gate473inter7), .O(gate473inter9));
  nand2 gate935(.a(s_55), .b(gate473inter3), .O(gate473inter10));
  nor2  gate936(.a(gate473inter10), .b(gate473inter9), .O(gate473inter11));
  nor2  gate937(.a(gate473inter11), .b(gate473inter6), .O(gate473inter12));
  nand2 gate938(.a(gate473inter12), .b(gate473inter1), .O(G1282));
nand2 gate474( .a(G1117), .b(G1213), .O(G1283) );

  xor2  gate1093(.a(G1216), .b(G29), .O(gate475inter0));
  nand2 gate1094(.a(gate475inter0), .b(s_78), .O(gate475inter1));
  and2  gate1095(.a(G1216), .b(G29), .O(gate475inter2));
  inv1  gate1096(.a(s_78), .O(gate475inter3));
  inv1  gate1097(.a(s_79), .O(gate475inter4));
  nand2 gate1098(.a(gate475inter4), .b(gate475inter3), .O(gate475inter5));
  nor2  gate1099(.a(gate475inter5), .b(gate475inter2), .O(gate475inter6));
  inv1  gate1100(.a(G29), .O(gate475inter7));
  inv1  gate1101(.a(G1216), .O(gate475inter8));
  nand2 gate1102(.a(gate475inter8), .b(gate475inter7), .O(gate475inter9));
  nand2 gate1103(.a(s_79), .b(gate475inter3), .O(gate475inter10));
  nor2  gate1104(.a(gate475inter10), .b(gate475inter9), .O(gate475inter11));
  nor2  gate1105(.a(gate475inter11), .b(gate475inter6), .O(gate475inter12));
  nand2 gate1106(.a(gate475inter12), .b(gate475inter1), .O(G1284));
nand2 gate476( .a(G1120), .b(G1216), .O(G1285) );
nand2 gate477( .a(G30), .b(G1219), .O(G1286) );
nand2 gate478( .a(G1123), .b(G1219), .O(G1287) );
nand2 gate479( .a(G31), .b(G1222), .O(G1288) );
nand2 gate480( .a(G1126), .b(G1222), .O(G1289) );

  xor2  gate1457(.a(G1225), .b(G32), .O(gate481inter0));
  nand2 gate1458(.a(gate481inter0), .b(s_130), .O(gate481inter1));
  and2  gate1459(.a(G1225), .b(G32), .O(gate481inter2));
  inv1  gate1460(.a(s_130), .O(gate481inter3));
  inv1  gate1461(.a(s_131), .O(gate481inter4));
  nand2 gate1462(.a(gate481inter4), .b(gate481inter3), .O(gate481inter5));
  nor2  gate1463(.a(gate481inter5), .b(gate481inter2), .O(gate481inter6));
  inv1  gate1464(.a(G32), .O(gate481inter7));
  inv1  gate1465(.a(G1225), .O(gate481inter8));
  nand2 gate1466(.a(gate481inter8), .b(gate481inter7), .O(gate481inter9));
  nand2 gate1467(.a(s_131), .b(gate481inter3), .O(gate481inter10));
  nor2  gate1468(.a(gate481inter10), .b(gate481inter9), .O(gate481inter11));
  nor2  gate1469(.a(gate481inter11), .b(gate481inter6), .O(gate481inter12));
  nand2 gate1470(.a(gate481inter12), .b(gate481inter1), .O(G1290));

  xor2  gate1625(.a(G1225), .b(G1129), .O(gate482inter0));
  nand2 gate1626(.a(gate482inter0), .b(s_154), .O(gate482inter1));
  and2  gate1627(.a(G1225), .b(G1129), .O(gate482inter2));
  inv1  gate1628(.a(s_154), .O(gate482inter3));
  inv1  gate1629(.a(s_155), .O(gate482inter4));
  nand2 gate1630(.a(gate482inter4), .b(gate482inter3), .O(gate482inter5));
  nor2  gate1631(.a(gate482inter5), .b(gate482inter2), .O(gate482inter6));
  inv1  gate1632(.a(G1129), .O(gate482inter7));
  inv1  gate1633(.a(G1225), .O(gate482inter8));
  nand2 gate1634(.a(gate482inter8), .b(gate482inter7), .O(gate482inter9));
  nand2 gate1635(.a(s_155), .b(gate482inter3), .O(gate482inter10));
  nor2  gate1636(.a(gate482inter10), .b(gate482inter9), .O(gate482inter11));
  nor2  gate1637(.a(gate482inter11), .b(gate482inter6), .O(gate482inter12));
  nand2 gate1638(.a(gate482inter12), .b(gate482inter1), .O(G1291));

  xor2  gate1891(.a(G1229), .b(G1228), .O(gate483inter0));
  nand2 gate1892(.a(gate483inter0), .b(s_192), .O(gate483inter1));
  and2  gate1893(.a(G1229), .b(G1228), .O(gate483inter2));
  inv1  gate1894(.a(s_192), .O(gate483inter3));
  inv1  gate1895(.a(s_193), .O(gate483inter4));
  nand2 gate1896(.a(gate483inter4), .b(gate483inter3), .O(gate483inter5));
  nor2  gate1897(.a(gate483inter5), .b(gate483inter2), .O(gate483inter6));
  inv1  gate1898(.a(G1228), .O(gate483inter7));
  inv1  gate1899(.a(G1229), .O(gate483inter8));
  nand2 gate1900(.a(gate483inter8), .b(gate483inter7), .O(gate483inter9));
  nand2 gate1901(.a(s_193), .b(gate483inter3), .O(gate483inter10));
  nor2  gate1902(.a(gate483inter10), .b(gate483inter9), .O(gate483inter11));
  nor2  gate1903(.a(gate483inter11), .b(gate483inter6), .O(gate483inter12));
  nand2 gate1904(.a(gate483inter12), .b(gate483inter1), .O(G1292));
nand2 gate484( .a(G1230), .b(G1231), .O(G1293) );

  xor2  gate2689(.a(G1233), .b(G1232), .O(gate485inter0));
  nand2 gate2690(.a(gate485inter0), .b(s_306), .O(gate485inter1));
  and2  gate2691(.a(G1233), .b(G1232), .O(gate485inter2));
  inv1  gate2692(.a(s_306), .O(gate485inter3));
  inv1  gate2693(.a(s_307), .O(gate485inter4));
  nand2 gate2694(.a(gate485inter4), .b(gate485inter3), .O(gate485inter5));
  nor2  gate2695(.a(gate485inter5), .b(gate485inter2), .O(gate485inter6));
  inv1  gate2696(.a(G1232), .O(gate485inter7));
  inv1  gate2697(.a(G1233), .O(gate485inter8));
  nand2 gate2698(.a(gate485inter8), .b(gate485inter7), .O(gate485inter9));
  nand2 gate2699(.a(s_307), .b(gate485inter3), .O(gate485inter10));
  nor2  gate2700(.a(gate485inter10), .b(gate485inter9), .O(gate485inter11));
  nor2  gate2701(.a(gate485inter11), .b(gate485inter6), .O(gate485inter12));
  nand2 gate2702(.a(gate485inter12), .b(gate485inter1), .O(G1294));
nand2 gate486( .a(G1234), .b(G1235), .O(G1295) );
nand2 gate487( .a(G1236), .b(G1237), .O(G1296) );

  xor2  gate2325(.a(G1239), .b(G1238), .O(gate488inter0));
  nand2 gate2326(.a(gate488inter0), .b(s_254), .O(gate488inter1));
  and2  gate2327(.a(G1239), .b(G1238), .O(gate488inter2));
  inv1  gate2328(.a(s_254), .O(gate488inter3));
  inv1  gate2329(.a(s_255), .O(gate488inter4));
  nand2 gate2330(.a(gate488inter4), .b(gate488inter3), .O(gate488inter5));
  nor2  gate2331(.a(gate488inter5), .b(gate488inter2), .O(gate488inter6));
  inv1  gate2332(.a(G1238), .O(gate488inter7));
  inv1  gate2333(.a(G1239), .O(gate488inter8));
  nand2 gate2334(.a(gate488inter8), .b(gate488inter7), .O(gate488inter9));
  nand2 gate2335(.a(s_255), .b(gate488inter3), .O(gate488inter10));
  nor2  gate2336(.a(gate488inter10), .b(gate488inter9), .O(gate488inter11));
  nor2  gate2337(.a(gate488inter11), .b(gate488inter6), .O(gate488inter12));
  nand2 gate2338(.a(gate488inter12), .b(gate488inter1), .O(G1297));
nand2 gate489( .a(G1240), .b(G1241), .O(G1298) );
nand2 gate490( .a(G1242), .b(G1243), .O(G1299) );
nand2 gate491( .a(G1244), .b(G1245), .O(G1300) );

  xor2  gate1275(.a(G1247), .b(G1246), .O(gate492inter0));
  nand2 gate1276(.a(gate492inter0), .b(s_104), .O(gate492inter1));
  and2  gate1277(.a(G1247), .b(G1246), .O(gate492inter2));
  inv1  gate1278(.a(s_104), .O(gate492inter3));
  inv1  gate1279(.a(s_105), .O(gate492inter4));
  nand2 gate1280(.a(gate492inter4), .b(gate492inter3), .O(gate492inter5));
  nor2  gate1281(.a(gate492inter5), .b(gate492inter2), .O(gate492inter6));
  inv1  gate1282(.a(G1246), .O(gate492inter7));
  inv1  gate1283(.a(G1247), .O(gate492inter8));
  nand2 gate1284(.a(gate492inter8), .b(gate492inter7), .O(gate492inter9));
  nand2 gate1285(.a(s_105), .b(gate492inter3), .O(gate492inter10));
  nor2  gate1286(.a(gate492inter10), .b(gate492inter9), .O(gate492inter11));
  nor2  gate1287(.a(gate492inter11), .b(gate492inter6), .O(gate492inter12));
  nand2 gate1288(.a(gate492inter12), .b(gate492inter1), .O(G1301));

  xor2  gate2087(.a(G1249), .b(G1248), .O(gate493inter0));
  nand2 gate2088(.a(gate493inter0), .b(s_220), .O(gate493inter1));
  and2  gate2089(.a(G1249), .b(G1248), .O(gate493inter2));
  inv1  gate2090(.a(s_220), .O(gate493inter3));
  inv1  gate2091(.a(s_221), .O(gate493inter4));
  nand2 gate2092(.a(gate493inter4), .b(gate493inter3), .O(gate493inter5));
  nor2  gate2093(.a(gate493inter5), .b(gate493inter2), .O(gate493inter6));
  inv1  gate2094(.a(G1248), .O(gate493inter7));
  inv1  gate2095(.a(G1249), .O(gate493inter8));
  nand2 gate2096(.a(gate493inter8), .b(gate493inter7), .O(gate493inter9));
  nand2 gate2097(.a(s_221), .b(gate493inter3), .O(gate493inter10));
  nor2  gate2098(.a(gate493inter10), .b(gate493inter9), .O(gate493inter11));
  nor2  gate2099(.a(gate493inter11), .b(gate493inter6), .O(gate493inter12));
  nand2 gate2100(.a(gate493inter12), .b(gate493inter1), .O(G1302));

  xor2  gate547(.a(G1251), .b(G1250), .O(gate494inter0));
  nand2 gate548(.a(gate494inter0), .b(s_0), .O(gate494inter1));
  and2  gate549(.a(G1251), .b(G1250), .O(gate494inter2));
  inv1  gate550(.a(s_0), .O(gate494inter3));
  inv1  gate551(.a(s_1), .O(gate494inter4));
  nand2 gate552(.a(gate494inter4), .b(gate494inter3), .O(gate494inter5));
  nor2  gate553(.a(gate494inter5), .b(gate494inter2), .O(gate494inter6));
  inv1  gate554(.a(G1250), .O(gate494inter7));
  inv1  gate555(.a(G1251), .O(gate494inter8));
  nand2 gate556(.a(gate494inter8), .b(gate494inter7), .O(gate494inter9));
  nand2 gate557(.a(s_1), .b(gate494inter3), .O(gate494inter10));
  nor2  gate558(.a(gate494inter10), .b(gate494inter9), .O(gate494inter11));
  nor2  gate559(.a(gate494inter11), .b(gate494inter6), .O(gate494inter12));
  nand2 gate560(.a(gate494inter12), .b(gate494inter1), .O(G1303));
nand2 gate495( .a(G1252), .b(G1253), .O(G1304) );

  xor2  gate3207(.a(G1255), .b(G1254), .O(gate496inter0));
  nand2 gate3208(.a(gate496inter0), .b(s_380), .O(gate496inter1));
  and2  gate3209(.a(G1255), .b(G1254), .O(gate496inter2));
  inv1  gate3210(.a(s_380), .O(gate496inter3));
  inv1  gate3211(.a(s_381), .O(gate496inter4));
  nand2 gate3212(.a(gate496inter4), .b(gate496inter3), .O(gate496inter5));
  nor2  gate3213(.a(gate496inter5), .b(gate496inter2), .O(gate496inter6));
  inv1  gate3214(.a(G1254), .O(gate496inter7));
  inv1  gate3215(.a(G1255), .O(gate496inter8));
  nand2 gate3216(.a(gate496inter8), .b(gate496inter7), .O(gate496inter9));
  nand2 gate3217(.a(s_381), .b(gate496inter3), .O(gate496inter10));
  nor2  gate3218(.a(gate496inter10), .b(gate496inter9), .O(gate496inter11));
  nor2  gate3219(.a(gate496inter11), .b(gate496inter6), .O(gate496inter12));
  nand2 gate3220(.a(gate496inter12), .b(gate496inter1), .O(G1305));
nand2 gate497( .a(G1256), .b(G1257), .O(G1306) );
nand2 gate498( .a(G1258), .b(G1259), .O(G1307) );
nand2 gate499( .a(G1260), .b(G1261), .O(G1308) );
nand2 gate500( .a(G1262), .b(G1263), .O(G1309) );

  xor2  gate2059(.a(G1265), .b(G1264), .O(gate501inter0));
  nand2 gate2060(.a(gate501inter0), .b(s_216), .O(gate501inter1));
  and2  gate2061(.a(G1265), .b(G1264), .O(gate501inter2));
  inv1  gate2062(.a(s_216), .O(gate501inter3));
  inv1  gate2063(.a(s_217), .O(gate501inter4));
  nand2 gate2064(.a(gate501inter4), .b(gate501inter3), .O(gate501inter5));
  nor2  gate2065(.a(gate501inter5), .b(gate501inter2), .O(gate501inter6));
  inv1  gate2066(.a(G1264), .O(gate501inter7));
  inv1  gate2067(.a(G1265), .O(gate501inter8));
  nand2 gate2068(.a(gate501inter8), .b(gate501inter7), .O(gate501inter9));
  nand2 gate2069(.a(s_217), .b(gate501inter3), .O(gate501inter10));
  nor2  gate2070(.a(gate501inter10), .b(gate501inter9), .O(gate501inter11));
  nor2  gate2071(.a(gate501inter11), .b(gate501inter6), .O(gate501inter12));
  nand2 gate2072(.a(gate501inter12), .b(gate501inter1), .O(G1310));

  xor2  gate3109(.a(G1267), .b(G1266), .O(gate502inter0));
  nand2 gate3110(.a(gate502inter0), .b(s_366), .O(gate502inter1));
  and2  gate3111(.a(G1267), .b(G1266), .O(gate502inter2));
  inv1  gate3112(.a(s_366), .O(gate502inter3));
  inv1  gate3113(.a(s_367), .O(gate502inter4));
  nand2 gate3114(.a(gate502inter4), .b(gate502inter3), .O(gate502inter5));
  nor2  gate3115(.a(gate502inter5), .b(gate502inter2), .O(gate502inter6));
  inv1  gate3116(.a(G1266), .O(gate502inter7));
  inv1  gate3117(.a(G1267), .O(gate502inter8));
  nand2 gate3118(.a(gate502inter8), .b(gate502inter7), .O(gate502inter9));
  nand2 gate3119(.a(s_367), .b(gate502inter3), .O(gate502inter10));
  nor2  gate3120(.a(gate502inter10), .b(gate502inter9), .O(gate502inter11));
  nor2  gate3121(.a(gate502inter11), .b(gate502inter6), .O(gate502inter12));
  nand2 gate3122(.a(gate502inter12), .b(gate502inter1), .O(G1311));
nand2 gate503( .a(G1268), .b(G1269), .O(G1312) );
nand2 gate504( .a(G1270), .b(G1271), .O(G1313) );
nand2 gate505( .a(G1272), .b(G1273), .O(G1314) );

  xor2  gate2759(.a(G1275), .b(G1274), .O(gate506inter0));
  nand2 gate2760(.a(gate506inter0), .b(s_316), .O(gate506inter1));
  and2  gate2761(.a(G1275), .b(G1274), .O(gate506inter2));
  inv1  gate2762(.a(s_316), .O(gate506inter3));
  inv1  gate2763(.a(s_317), .O(gate506inter4));
  nand2 gate2764(.a(gate506inter4), .b(gate506inter3), .O(gate506inter5));
  nor2  gate2765(.a(gate506inter5), .b(gate506inter2), .O(gate506inter6));
  inv1  gate2766(.a(G1274), .O(gate506inter7));
  inv1  gate2767(.a(G1275), .O(gate506inter8));
  nand2 gate2768(.a(gate506inter8), .b(gate506inter7), .O(gate506inter9));
  nand2 gate2769(.a(s_317), .b(gate506inter3), .O(gate506inter10));
  nor2  gate2770(.a(gate506inter10), .b(gate506inter9), .O(gate506inter11));
  nor2  gate2771(.a(gate506inter11), .b(gate506inter6), .O(gate506inter12));
  nand2 gate2772(.a(gate506inter12), .b(gate506inter1), .O(G1315));

  xor2  gate3179(.a(G1277), .b(G1276), .O(gate507inter0));
  nand2 gate3180(.a(gate507inter0), .b(s_376), .O(gate507inter1));
  and2  gate3181(.a(G1277), .b(G1276), .O(gate507inter2));
  inv1  gate3182(.a(s_376), .O(gate507inter3));
  inv1  gate3183(.a(s_377), .O(gate507inter4));
  nand2 gate3184(.a(gate507inter4), .b(gate507inter3), .O(gate507inter5));
  nor2  gate3185(.a(gate507inter5), .b(gate507inter2), .O(gate507inter6));
  inv1  gate3186(.a(G1276), .O(gate507inter7));
  inv1  gate3187(.a(G1277), .O(gate507inter8));
  nand2 gate3188(.a(gate507inter8), .b(gate507inter7), .O(gate507inter9));
  nand2 gate3189(.a(s_377), .b(gate507inter3), .O(gate507inter10));
  nor2  gate3190(.a(gate507inter10), .b(gate507inter9), .O(gate507inter11));
  nor2  gate3191(.a(gate507inter11), .b(gate507inter6), .O(gate507inter12));
  nand2 gate3192(.a(gate507inter12), .b(gate507inter1), .O(G1316));
nand2 gate508( .a(G1278), .b(G1279), .O(G1317) );

  xor2  gate2171(.a(G1281), .b(G1280), .O(gate509inter0));
  nand2 gate2172(.a(gate509inter0), .b(s_232), .O(gate509inter1));
  and2  gate2173(.a(G1281), .b(G1280), .O(gate509inter2));
  inv1  gate2174(.a(s_232), .O(gate509inter3));
  inv1  gate2175(.a(s_233), .O(gate509inter4));
  nand2 gate2176(.a(gate509inter4), .b(gate509inter3), .O(gate509inter5));
  nor2  gate2177(.a(gate509inter5), .b(gate509inter2), .O(gate509inter6));
  inv1  gate2178(.a(G1280), .O(gate509inter7));
  inv1  gate2179(.a(G1281), .O(gate509inter8));
  nand2 gate2180(.a(gate509inter8), .b(gate509inter7), .O(gate509inter9));
  nand2 gate2181(.a(s_233), .b(gate509inter3), .O(gate509inter10));
  nor2  gate2182(.a(gate509inter10), .b(gate509inter9), .O(gate509inter11));
  nor2  gate2183(.a(gate509inter11), .b(gate509inter6), .O(gate509inter12));
  nand2 gate2184(.a(gate509inter12), .b(gate509inter1), .O(G1318));

  xor2  gate2521(.a(G1283), .b(G1282), .O(gate510inter0));
  nand2 gate2522(.a(gate510inter0), .b(s_282), .O(gate510inter1));
  and2  gate2523(.a(G1283), .b(G1282), .O(gate510inter2));
  inv1  gate2524(.a(s_282), .O(gate510inter3));
  inv1  gate2525(.a(s_283), .O(gate510inter4));
  nand2 gate2526(.a(gate510inter4), .b(gate510inter3), .O(gate510inter5));
  nor2  gate2527(.a(gate510inter5), .b(gate510inter2), .O(gate510inter6));
  inv1  gate2528(.a(G1282), .O(gate510inter7));
  inv1  gate2529(.a(G1283), .O(gate510inter8));
  nand2 gate2530(.a(gate510inter8), .b(gate510inter7), .O(gate510inter9));
  nand2 gate2531(.a(s_283), .b(gate510inter3), .O(gate510inter10));
  nor2  gate2532(.a(gate510inter10), .b(gate510inter9), .O(gate510inter11));
  nor2  gate2533(.a(gate510inter11), .b(gate510inter6), .O(gate510inter12));
  nand2 gate2534(.a(gate510inter12), .b(gate510inter1), .O(G1319));
nand2 gate511( .a(G1284), .b(G1285), .O(G1320) );

  xor2  gate771(.a(G1287), .b(G1286), .O(gate512inter0));
  nand2 gate772(.a(gate512inter0), .b(s_32), .O(gate512inter1));
  and2  gate773(.a(G1287), .b(G1286), .O(gate512inter2));
  inv1  gate774(.a(s_32), .O(gate512inter3));
  inv1  gate775(.a(s_33), .O(gate512inter4));
  nand2 gate776(.a(gate512inter4), .b(gate512inter3), .O(gate512inter5));
  nor2  gate777(.a(gate512inter5), .b(gate512inter2), .O(gate512inter6));
  inv1  gate778(.a(G1286), .O(gate512inter7));
  inv1  gate779(.a(G1287), .O(gate512inter8));
  nand2 gate780(.a(gate512inter8), .b(gate512inter7), .O(gate512inter9));
  nand2 gate781(.a(s_33), .b(gate512inter3), .O(gate512inter10));
  nor2  gate782(.a(gate512inter10), .b(gate512inter9), .O(gate512inter11));
  nor2  gate783(.a(gate512inter11), .b(gate512inter6), .O(gate512inter12));
  nand2 gate784(.a(gate512inter12), .b(gate512inter1), .O(G1321));

  xor2  gate701(.a(G1289), .b(G1288), .O(gate513inter0));
  nand2 gate702(.a(gate513inter0), .b(s_22), .O(gate513inter1));
  and2  gate703(.a(G1289), .b(G1288), .O(gate513inter2));
  inv1  gate704(.a(s_22), .O(gate513inter3));
  inv1  gate705(.a(s_23), .O(gate513inter4));
  nand2 gate706(.a(gate513inter4), .b(gate513inter3), .O(gate513inter5));
  nor2  gate707(.a(gate513inter5), .b(gate513inter2), .O(gate513inter6));
  inv1  gate708(.a(G1288), .O(gate513inter7));
  inv1  gate709(.a(G1289), .O(gate513inter8));
  nand2 gate710(.a(gate513inter8), .b(gate513inter7), .O(gate513inter9));
  nand2 gate711(.a(s_23), .b(gate513inter3), .O(gate513inter10));
  nor2  gate712(.a(gate513inter10), .b(gate513inter9), .O(gate513inter11));
  nor2  gate713(.a(gate513inter11), .b(gate513inter6), .O(gate513inter12));
  nand2 gate714(.a(gate513inter12), .b(gate513inter1), .O(G1322));

  xor2  gate1401(.a(G1291), .b(G1290), .O(gate514inter0));
  nand2 gate1402(.a(gate514inter0), .b(s_122), .O(gate514inter1));
  and2  gate1403(.a(G1291), .b(G1290), .O(gate514inter2));
  inv1  gate1404(.a(s_122), .O(gate514inter3));
  inv1  gate1405(.a(s_123), .O(gate514inter4));
  nand2 gate1406(.a(gate514inter4), .b(gate514inter3), .O(gate514inter5));
  nor2  gate1407(.a(gate514inter5), .b(gate514inter2), .O(gate514inter6));
  inv1  gate1408(.a(G1290), .O(gate514inter7));
  inv1  gate1409(.a(G1291), .O(gate514inter8));
  nand2 gate1410(.a(gate514inter8), .b(gate514inter7), .O(gate514inter9));
  nand2 gate1411(.a(s_123), .b(gate514inter3), .O(gate514inter10));
  nor2  gate1412(.a(gate514inter10), .b(gate514inter9), .O(gate514inter11));
  nor2  gate1413(.a(gate514inter11), .b(gate514inter6), .O(gate514inter12));
  nand2 gate1414(.a(gate514inter12), .b(gate514inter1), .O(G1323));
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule