module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);

input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;//RE__PI;

input s_0,s_1;//RE__ALLOW(00,01,10,11);
input s_2,s_3;//RE__ALLOW(00,01,10,11);
input s_4,s_5;//RE__ALLOW(00,01,10,11);
input s_6,s_7;//RE__ALLOW(00,01,10,11);
input s_8,s_9;//RE__ALLOW(00,01,10,11);
input s_10,s_11;//RE__ALLOW(00,01,10,11);
input s_12,s_13;//RE__ALLOW(00,01,10,11);
input s_14,s_15;//RE__ALLOW(00,01,10,11);
input s_16,s_17;//RE__ALLOW(00,01,10,11);
input s_18,s_19;//RE__ALLOW(00,01,10,11);
input s_20,s_21;//RE__ALLOW(00,01,10,11);
input s_22,s_23;//RE__ALLOW(00,01,10,11);
input s_24,s_25;//RE__ALLOW(00,01,10,11);
input s_26,s_27;//RE__ALLOW(00,01,10,11);
input s_28,s_29;//RE__ALLOW(00,01,10,11);
input s_30,s_31;//RE__ALLOW(00,01,10,11);
input s_32,s_33;//RE__ALLOW(00,01,10,11);
input s_34,s_35;//RE__ALLOW(00,01,10,11);
input s_36,s_37;//RE__ALLOW(00,01,10,11);
input s_38,s_39;//RE__ALLOW(00,01,10,11);
input s_40,s_41;//RE__ALLOW(00,01,10,11);
input s_42,s_43;//RE__ALLOW(00,01,10,11);
input s_44,s_45;//RE__ALLOW(00,01,10,11);
input s_46,s_47;//RE__ALLOW(00,01,10,11);
input s_48,s_49;//RE__ALLOW(00,01,10,11);
input s_50,s_51;//RE__ALLOW(00,01,10,11);
input s_52,s_53;//RE__ALLOW(00,01,10,11);
input s_54,s_55;//RE__ALLOW(00,01,10,11);
input s_56,s_57;//RE__ALLOW(00,01,10,11);
input s_58,s_59;//RE__ALLOW(00,01,10,11);
input s_60,s_61;//RE__ALLOW(00,01,10,11);
input s_62,s_63;//RE__ALLOW(00,01,10,11);
input s_64,s_65;//RE__ALLOW(00,01,10,11);
input s_66,s_67;//RE__ALLOW(00,01,10,11);
input s_68,s_69;//RE__ALLOW(00,01,10,11);
input s_70,s_71;//RE__ALLOW(00,01,10,11);
input s_72,s_73;//RE__ALLOW(00,01,10,11);
input s_74,s_75;//RE__ALLOW(00,01,10,11);
input s_76,s_77;//RE__ALLOW(00,01,10,11);
input s_78,s_79;//RE__ALLOW(00,01,10,11);
input s_80,s_81;//RE__ALLOW(00,01,10,11);
input s_82,s_83;//RE__ALLOW(00,01,10,11);
input s_84,s_85;//RE__ALLOW(00,01,10,11);
input s_86,s_87;//RE__ALLOW(00,01,10,11);
input s_88,s_89;//RE__ALLOW(00,01,10,11);
input s_90,s_91;//RE__ALLOW(00,01,10,11);
input s_92,s_93;//RE__ALLOW(00,01,10,11);
input s_94,s_95;//RE__ALLOW(00,01,10,11);
input s_96,s_97;//RE__ALLOW(00,01,10,11);
input s_98,s_99;//RE__ALLOW(00,01,10,11);
input s_100,s_101;//RE__ALLOW(00,01,10,11);
input s_102,s_103;//RE__ALLOW(00,01,10,11);
input s_104,s_105;//RE__ALLOW(00,01,10,11);
input s_106,s_107;//RE__ALLOW(00,01,10,11);
input s_108,s_109;//RE__ALLOW(00,01,10,11);
input s_110,s_111;//RE__ALLOW(00,01,10,11);
input s_112,s_113;//RE__ALLOW(00,01,10,11);
input s_114,s_115;//RE__ALLOW(00,01,10,11);
input s_116,s_117;//RE__ALLOW(00,01,10,11);
input s_118,s_119;//RE__ALLOW(00,01,10,11);
input s_120,s_121;//RE__ALLOW(00,01,10,11);
input s_122,s_123;//RE__ALLOW(00,01,10,11);
input s_124,s_125;//RE__ALLOW(00,01,10,11);
input s_126,s_127;//RE__ALLOW(00,01,10,11);
input s_128,s_129;//RE__ALLOW(00,01,10,11);
input s_130,s_131;//RE__ALLOW(00,01,10,11);
input s_132,s_133;//RE__ALLOW(00,01,10,11);
input s_134,s_135;//RE__ALLOW(00,01,10,11);
input s_136,s_137;//RE__ALLOW(00,01,10,11);
input s_138,s_139;//RE__ALLOW(00,01,10,11);
input s_140,s_141;//RE__ALLOW(00,01,10,11);
input s_142,s_143;//RE__ALLOW(00,01,10,11);
input s_144,s_145;//RE__ALLOW(00,01,10,11);
input s_146,s_147;//RE__ALLOW(00,01,10,11);
input s_148,s_149;//RE__ALLOW(00,01,10,11);
input s_150,s_151;//RE__ALLOW(00,01,10,11);
input s_152,s_153;//RE__ALLOW(00,01,10,11);
input s_154,s_155;//RE__ALLOW(00,01,10,11);
input s_156,s_157;//RE__ALLOW(00,01,10,11);
input s_158,s_159;//RE__ALLOW(00,01,10,11);
input s_160,s_161;//RE__ALLOW(00,01,10,11);
input s_162,s_163;//RE__ALLOW(00,01,10,11);
input s_164,s_165;//RE__ALLOW(00,01,10,11);
input s_166,s_167;//RE__ALLOW(00,01,10,11);
input s_168,s_169;//RE__ALLOW(00,01,10,11);
input s_170,s_171;//RE__ALLOW(00,01,10,11);
input s_172,s_173;//RE__ALLOW(00,01,10,11);
input s_174,s_175;//RE__ALLOW(00,01,10,11);
input s_176,s_177;//RE__ALLOW(00,01,10,11);
input s_178,s_179;//RE__ALLOW(00,01,10,11);
input s_180,s_181;//RE__ALLOW(00,01,10,11);
input s_182,s_183;//RE__ALLOW(00,01,10,11);
input s_184,s_185;//RE__ALLOW(00,01,10,11);
input s_186,s_187;//RE__ALLOW(00,01,10,11);
input s_188,s_189;//RE__ALLOW(00,01,10,11);
input s_190,s_191;//RE__ALLOW(00,01,10,11);
input s_192,s_193;//RE__ALLOW(00,01,10,11);
input s_194,s_195;//RE__ALLOW(00,01,10,11);
input s_196,s_197;//RE__ALLOW(00,01,10,11);
input s_198,s_199;//RE__ALLOW(00,01,10,11);
input s_200,s_201;//RE__ALLOW(00,01,10,11);
input s_202,s_203;//RE__ALLOW(00,01,10,11);
input s_204,s_205;//RE__ALLOW(00,01,10,11);
input s_206,s_207;//RE__ALLOW(00,01,10,11);
input s_208,s_209;//RE__ALLOW(00,01,10,11);
input s_210,s_211;//RE__ALLOW(00,01,10,11);
input s_212,s_213;//RE__ALLOW(00,01,10,11);
input s_214,s_215;//RE__ALLOW(00,01,10,11);
input s_216,s_217;//RE__ALLOW(00,01,10,11);
input s_218,s_219;//RE__ALLOW(00,01,10,11);
input s_220,s_221;//RE__ALLOW(00,01,10,11);
input s_222,s_223;//RE__ALLOW(00,01,10,11);
input s_224,s_225;//RE__ALLOW(00,01,10,11);
input s_226,s_227;//RE__ALLOW(00,01,10,11);
input s_228,s_229;//RE__ALLOW(00,01,10,11);
input s_230,s_231;//RE__ALLOW(00,01,10,11);
input s_232,s_233;//RE__ALLOW(00,01,10,11);
input s_234,s_235;//RE__ALLOW(00,01,10,11);
input s_236,s_237;//RE__ALLOW(00,01,10,11);
input s_238,s_239;//RE__ALLOW(00,01,10,11);
input s_240,s_241;//RE__ALLOW(00,01,10,11);
input s_242,s_243;//RE__ALLOW(00,01,10,11);
input s_244,s_245;//RE__ALLOW(00,01,10,11);
input s_246,s_247;//RE__ALLOW(00,01,10,11);
input s_248,s_249;//RE__ALLOW(00,01,10,11);
input s_250,s_251;//RE__ALLOW(00,01,10,11);
input s_252,s_253;//RE__ALLOW(00,01,10,11);
input s_254,s_255;//RE__ALLOW(00,01,10,11);
input s_256,s_257;//RE__ALLOW(00,01,10,11);
input s_258,s_259;//RE__ALLOW(00,01,10,11);
input s_260,s_261;//RE__ALLOW(00,01,10,11);
input s_262,s_263;//RE__ALLOW(00,01,10,11);
input s_264,s_265;//RE__ALLOW(00,01,10,11);
input s_266,s_267;//RE__ALLOW(00,01,10,11);
input s_268,s_269;//RE__ALLOW(00,01,10,11);
input s_270,s_271;//RE__ALLOW(00,01,10,11);
input s_272,s_273;//RE__ALLOW(00,01,10,11);
input s_274,s_275;//RE__ALLOW(00,01,10,11);
input s_276,s_277;//RE__ALLOW(00,01,10,11);
input s_278,s_279;//RE__ALLOW(00,01,10,11);
input s_280,s_281;//RE__ALLOW(00,01,10,11);
input s_282,s_283;//RE__ALLOW(00,01,10,11);
input s_284,s_285;//RE__ALLOW(00,01,10,11);
input s_286,s_287;//RE__ALLOW(00,01,10,11);
input s_288,s_289;//RE__ALLOW(00,01,10,11);
input s_290,s_291;//RE__ALLOW(00,01,10,11);
input s_292,s_293;//RE__ALLOW(00,01,10,11);
input s_294,s_295;//RE__ALLOW(00,01,10,11);
input s_296,s_297;//RE__ALLOW(00,01,10,11);
input s_298,s_299;//RE__ALLOW(00,01,10,11);
input s_300,s_301;//RE__ALLOW(00,01,10,11);
input s_302,s_303;//RE__ALLOW(00,01,10,11);
input s_304,s_305;//RE__ALLOW(00,01,10,11);
input s_306,s_307;//RE__ALLOW(00,01,10,11);
input s_308,s_309;//RE__ALLOW(00,01,10,11);
input s_310,s_311;//RE__ALLOW(00,01,10,11);
input s_312,s_313;//RE__ALLOW(00,01,10,11);
input s_314,s_315;//RE__ALLOW(00,01,10,11);
input s_316,s_317;//RE__ALLOW(00,01,10,11);
input s_318,s_319;//RE__ALLOW(00,01,10,11);
input s_320,s_321;//RE__ALLOW(00,01,10,11);
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;

  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate435inter0, gate435inter1, gate435inter2, gate435inter3, gate435inter4, gate435inter5, gate435inter6, gate435inter7, gate435inter8, gate435inter9, gate435inter10, gate435inter11, gate435inter12, gate450inter0, gate450inter1, gate450inter2, gate450inter3, gate450inter4, gate450inter5, gate450inter6, gate450inter7, gate450inter8, gate450inter9, gate450inter10, gate450inter11, gate450inter12, gate271inter0, gate271inter1, gate271inter2, gate271inter3, gate271inter4, gate271inter5, gate271inter6, gate271inter7, gate271inter8, gate271inter9, gate271inter10, gate271inter11, gate271inter12, gate257inter0, gate257inter1, gate257inter2, gate257inter3, gate257inter4, gate257inter5, gate257inter6, gate257inter7, gate257inter8, gate257inter9, gate257inter10, gate257inter11, gate257inter12, gate43inter0, gate43inter1, gate43inter2, gate43inter3, gate43inter4, gate43inter5, gate43inter6, gate43inter7, gate43inter8, gate43inter9, gate43inter10, gate43inter11, gate43inter12, gate393inter0, gate393inter1, gate393inter2, gate393inter3, gate393inter4, gate393inter5, gate393inter6, gate393inter7, gate393inter8, gate393inter9, gate393inter10, gate393inter11, gate393inter12, gate32inter0, gate32inter1, gate32inter2, gate32inter3, gate32inter4, gate32inter5, gate32inter6, gate32inter7, gate32inter8, gate32inter9, gate32inter10, gate32inter11, gate32inter12, gate104inter0, gate104inter1, gate104inter2, gate104inter3, gate104inter4, gate104inter5, gate104inter6, gate104inter7, gate104inter8, gate104inter9, gate104inter10, gate104inter11, gate104inter12, gate224inter0, gate224inter1, gate224inter2, gate224inter3, gate224inter4, gate224inter5, gate224inter6, gate224inter7, gate224inter8, gate224inter9, gate224inter10, gate224inter11, gate224inter12, gate227inter0, gate227inter1, gate227inter2, gate227inter3, gate227inter4, gate227inter5, gate227inter6, gate227inter7, gate227inter8, gate227inter9, gate227inter10, gate227inter11, gate227inter12, gate75inter0, gate75inter1, gate75inter2, gate75inter3, gate75inter4, gate75inter5, gate75inter6, gate75inter7, gate75inter8, gate75inter9, gate75inter10, gate75inter11, gate75inter12, gate426inter0, gate426inter1, gate426inter2, gate426inter3, gate426inter4, gate426inter5, gate426inter6, gate426inter7, gate426inter8, gate426inter9, gate426inter10, gate426inter11, gate426inter12, gate112inter0, gate112inter1, gate112inter2, gate112inter3, gate112inter4, gate112inter5, gate112inter6, gate112inter7, gate112inter8, gate112inter9, gate112inter10, gate112inter11, gate112inter12, gate136inter0, gate136inter1, gate136inter2, gate136inter3, gate136inter4, gate136inter5, gate136inter6, gate136inter7, gate136inter8, gate136inter9, gate136inter10, gate136inter11, gate136inter12, gate46inter0, gate46inter1, gate46inter2, gate46inter3, gate46inter4, gate46inter5, gate46inter6, gate46inter7, gate46inter8, gate46inter9, gate46inter10, gate46inter11, gate46inter12, gate248inter0, gate248inter1, gate248inter2, gate248inter3, gate248inter4, gate248inter5, gate248inter6, gate248inter7, gate248inter8, gate248inter9, gate248inter10, gate248inter11, gate248inter12, gate507inter0, gate507inter1, gate507inter2, gate507inter3, gate507inter4, gate507inter5, gate507inter6, gate507inter7, gate507inter8, gate507inter9, gate507inter10, gate507inter11, gate507inter12, gate137inter0, gate137inter1, gate137inter2, gate137inter3, gate137inter4, gate137inter5, gate137inter6, gate137inter7, gate137inter8, gate137inter9, gate137inter10, gate137inter11, gate137inter12, gate10inter0, gate10inter1, gate10inter2, gate10inter3, gate10inter4, gate10inter5, gate10inter6, gate10inter7, gate10inter8, gate10inter9, gate10inter10, gate10inter11, gate10inter12, gate229inter0, gate229inter1, gate229inter2, gate229inter3, gate229inter4, gate229inter5, gate229inter6, gate229inter7, gate229inter8, gate229inter9, gate229inter10, gate229inter11, gate229inter12, gate155inter0, gate155inter1, gate155inter2, gate155inter3, gate155inter4, gate155inter5, gate155inter6, gate155inter7, gate155inter8, gate155inter9, gate155inter10, gate155inter11, gate155inter12, gate171inter0, gate171inter1, gate171inter2, gate171inter3, gate171inter4, gate171inter5, gate171inter6, gate171inter7, gate171inter8, gate171inter9, gate171inter10, gate171inter11, gate171inter12, gate294inter0, gate294inter1, gate294inter2, gate294inter3, gate294inter4, gate294inter5, gate294inter6, gate294inter7, gate294inter8, gate294inter9, gate294inter10, gate294inter11, gate294inter12, gate151inter0, gate151inter1, gate151inter2, gate151inter3, gate151inter4, gate151inter5, gate151inter6, gate151inter7, gate151inter8, gate151inter9, gate151inter10, gate151inter11, gate151inter12, gate169inter0, gate169inter1, gate169inter2, gate169inter3, gate169inter4, gate169inter5, gate169inter6, gate169inter7, gate169inter8, gate169inter9, gate169inter10, gate169inter11, gate169inter12, gate133inter0, gate133inter1, gate133inter2, gate133inter3, gate133inter4, gate133inter5, gate133inter6, gate133inter7, gate133inter8, gate133inter9, gate133inter10, gate133inter11, gate133inter12, gate499inter0, gate499inter1, gate499inter2, gate499inter3, gate499inter4, gate499inter5, gate499inter6, gate499inter7, gate499inter8, gate499inter9, gate499inter10, gate499inter11, gate499inter12, gate85inter0, gate85inter1, gate85inter2, gate85inter3, gate85inter4, gate85inter5, gate85inter6, gate85inter7, gate85inter8, gate85inter9, gate85inter10, gate85inter11, gate85inter12, gate116inter0, gate116inter1, gate116inter2, gate116inter3, gate116inter4, gate116inter5, gate116inter6, gate116inter7, gate116inter8, gate116inter9, gate116inter10, gate116inter11, gate116inter12, gate486inter0, gate486inter1, gate486inter2, gate486inter3, gate486inter4, gate486inter5, gate486inter6, gate486inter7, gate486inter8, gate486inter9, gate486inter10, gate486inter11, gate486inter12, gate502inter0, gate502inter1, gate502inter2, gate502inter3, gate502inter4, gate502inter5, gate502inter6, gate502inter7, gate502inter8, gate502inter9, gate502inter10, gate502inter11, gate502inter12, gate401inter0, gate401inter1, gate401inter2, gate401inter3, gate401inter4, gate401inter5, gate401inter6, gate401inter7, gate401inter8, gate401inter9, gate401inter10, gate401inter11, gate401inter12, gate398inter0, gate398inter1, gate398inter2, gate398inter3, gate398inter4, gate398inter5, gate398inter6, gate398inter7, gate398inter8, gate398inter9, gate398inter10, gate398inter11, gate398inter12, gate418inter0, gate418inter1, gate418inter2, gate418inter3, gate418inter4, gate418inter5, gate418inter6, gate418inter7, gate418inter8, gate418inter9, gate418inter10, gate418inter11, gate418inter12, gate253inter0, gate253inter1, gate253inter2, gate253inter3, gate253inter4, gate253inter5, gate253inter6, gate253inter7, gate253inter8, gate253inter9, gate253inter10, gate253inter11, gate253inter12, gate49inter0, gate49inter1, gate49inter2, gate49inter3, gate49inter4, gate49inter5, gate49inter6, gate49inter7, gate49inter8, gate49inter9, gate49inter10, gate49inter11, gate49inter12, gate128inter0, gate128inter1, gate128inter2, gate128inter3, gate128inter4, gate128inter5, gate128inter6, gate128inter7, gate128inter8, gate128inter9, gate128inter10, gate128inter11, gate128inter12, gate437inter0, gate437inter1, gate437inter2, gate437inter3, gate437inter4, gate437inter5, gate437inter6, gate437inter7, gate437inter8, gate437inter9, gate437inter10, gate437inter11, gate437inter12, gate216inter0, gate216inter1, gate216inter2, gate216inter3, gate216inter4, gate216inter5, gate216inter6, gate216inter7, gate216inter8, gate216inter9, gate216inter10, gate216inter11, gate216inter12, gate183inter0, gate183inter1, gate183inter2, gate183inter3, gate183inter4, gate183inter5, gate183inter6, gate183inter7, gate183inter8, gate183inter9, gate183inter10, gate183inter11, gate183inter12, gate404inter0, gate404inter1, gate404inter2, gate404inter3, gate404inter4, gate404inter5, gate404inter6, gate404inter7, gate404inter8, gate404inter9, gate404inter10, gate404inter11, gate404inter12, gate124inter0, gate124inter1, gate124inter2, gate124inter3, gate124inter4, gate124inter5, gate124inter6, gate124inter7, gate124inter8, gate124inter9, gate124inter10, gate124inter11, gate124inter12, gate130inter0, gate130inter1, gate130inter2, gate130inter3, gate130inter4, gate130inter5, gate130inter6, gate130inter7, gate130inter8, gate130inter9, gate130inter10, gate130inter11, gate130inter12, gate479inter0, gate479inter1, gate479inter2, gate479inter3, gate479inter4, gate479inter5, gate479inter6, gate479inter7, gate479inter8, gate479inter9, gate479inter10, gate479inter11, gate479inter12, gate208inter0, gate208inter1, gate208inter2, gate208inter3, gate208inter4, gate208inter5, gate208inter6, gate208inter7, gate208inter8, gate208inter9, gate208inter10, gate208inter11, gate208inter12, gate44inter0, gate44inter1, gate44inter2, gate44inter3, gate44inter4, gate44inter5, gate44inter6, gate44inter7, gate44inter8, gate44inter9, gate44inter10, gate44inter11, gate44inter12, gate213inter0, gate213inter1, gate213inter2, gate213inter3, gate213inter4, gate213inter5, gate213inter6, gate213inter7, gate213inter8, gate213inter9, gate213inter10, gate213inter11, gate213inter12, gate115inter0, gate115inter1, gate115inter2, gate115inter3, gate115inter4, gate115inter5, gate115inter6, gate115inter7, gate115inter8, gate115inter9, gate115inter10, gate115inter11, gate115inter12, gate400inter0, gate400inter1, gate400inter2, gate400inter3, gate400inter4, gate400inter5, gate400inter6, gate400inter7, gate400inter8, gate400inter9, gate400inter10, gate400inter11, gate400inter12, gate94inter0, gate94inter1, gate94inter2, gate94inter3, gate94inter4, gate94inter5, gate94inter6, gate94inter7, gate94inter8, gate94inter9, gate94inter10, gate94inter11, gate94inter12, gate498inter0, gate498inter1, gate498inter2, gate498inter3, gate498inter4, gate498inter5, gate498inter6, gate498inter7, gate498inter8, gate498inter9, gate498inter10, gate498inter11, gate498inter12, gate191inter0, gate191inter1, gate191inter2, gate191inter3, gate191inter4, gate191inter5, gate191inter6, gate191inter7, gate191inter8, gate191inter9, gate191inter10, gate191inter11, gate191inter12, gate158inter0, gate158inter1, gate158inter2, gate158inter3, gate158inter4, gate158inter5, gate158inter6, gate158inter7, gate158inter8, gate158inter9, gate158inter10, gate158inter11, gate158inter12, gate496inter0, gate496inter1, gate496inter2, gate496inter3, gate496inter4, gate496inter5, gate496inter6, gate496inter7, gate496inter8, gate496inter9, gate496inter10, gate496inter11, gate496inter12, gate172inter0, gate172inter1, gate172inter2, gate172inter3, gate172inter4, gate172inter5, gate172inter6, gate172inter7, gate172inter8, gate172inter9, gate172inter10, gate172inter11, gate172inter12, gate165inter0, gate165inter1, gate165inter2, gate165inter3, gate165inter4, gate165inter5, gate165inter6, gate165inter7, gate165inter8, gate165inter9, gate165inter10, gate165inter11, gate165inter12, gate296inter0, gate296inter1, gate296inter2, gate296inter3, gate296inter4, gate296inter5, gate296inter6, gate296inter7, gate296inter8, gate296inter9, gate296inter10, gate296inter11, gate296inter12, gate63inter0, gate63inter1, gate63inter2, gate63inter3, gate63inter4, gate63inter5, gate63inter6, gate63inter7, gate63inter8, gate63inter9, gate63inter10, gate63inter11, gate63inter12, gate230inter0, gate230inter1, gate230inter2, gate230inter3, gate230inter4, gate230inter5, gate230inter6, gate230inter7, gate230inter8, gate230inter9, gate230inter10, gate230inter11, gate230inter12, gate184inter0, gate184inter1, gate184inter2, gate184inter3, gate184inter4, gate184inter5, gate184inter6, gate184inter7, gate184inter8, gate184inter9, gate184inter10, gate184inter11, gate184inter12, gate232inter0, gate232inter1, gate232inter2, gate232inter3, gate232inter4, gate232inter5, gate232inter6, gate232inter7, gate232inter8, gate232inter9, gate232inter10, gate232inter11, gate232inter12, gate396inter0, gate396inter1, gate396inter2, gate396inter3, gate396inter4, gate396inter5, gate396inter6, gate396inter7, gate396inter8, gate396inter9, gate396inter10, gate396inter11, gate396inter12, gate185inter0, gate185inter1, gate185inter2, gate185inter3, gate185inter4, gate185inter5, gate185inter6, gate185inter7, gate185inter8, gate185inter9, gate185inter10, gate185inter11, gate185inter12, gate449inter0, gate449inter1, gate449inter2, gate449inter3, gate449inter4, gate449inter5, gate449inter6, gate449inter7, gate449inter8, gate449inter9, gate449inter10, gate449inter11, gate449inter12, gate261inter0, gate261inter1, gate261inter2, gate261inter3, gate261inter4, gate261inter5, gate261inter6, gate261inter7, gate261inter8, gate261inter9, gate261inter10, gate261inter11, gate261inter12, gate119inter0, gate119inter1, gate119inter2, gate119inter3, gate119inter4, gate119inter5, gate119inter6, gate119inter7, gate119inter8, gate119inter9, gate119inter10, gate119inter11, gate119inter12, gate188inter0, gate188inter1, gate188inter2, gate188inter3, gate188inter4, gate188inter5, gate188inter6, gate188inter7, gate188inter8, gate188inter9, gate188inter10, gate188inter11, gate188inter12, gate233inter0, gate233inter1, gate233inter2, gate233inter3, gate233inter4, gate233inter5, gate233inter6, gate233inter7, gate233inter8, gate233inter9, gate233inter10, gate233inter11, gate233inter12, gate471inter0, gate471inter1, gate471inter2, gate471inter3, gate471inter4, gate471inter5, gate471inter6, gate471inter7, gate471inter8, gate471inter9, gate471inter10, gate471inter11, gate471inter12, gate387inter0, gate387inter1, gate387inter2, gate387inter3, gate387inter4, gate387inter5, gate387inter6, gate387inter7, gate387inter8, gate387inter9, gate387inter10, gate387inter11, gate387inter12, gate167inter0, gate167inter1, gate167inter2, gate167inter3, gate167inter4, gate167inter5, gate167inter6, gate167inter7, gate167inter8, gate167inter9, gate167inter10, gate167inter11, gate167inter12, gate495inter0, gate495inter1, gate495inter2, gate495inter3, gate495inter4, gate495inter5, gate495inter6, gate495inter7, gate495inter8, gate495inter9, gate495inter10, gate495inter11, gate495inter12, gate200inter0, gate200inter1, gate200inter2, gate200inter3, gate200inter4, gate200inter5, gate200inter6, gate200inter7, gate200inter8, gate200inter9, gate200inter10, gate200inter11, gate200inter12, gate407inter0, gate407inter1, gate407inter2, gate407inter3, gate407inter4, gate407inter5, gate407inter6, gate407inter7, gate407inter8, gate407inter9, gate407inter10, gate407inter11, gate407inter12, gate429inter0, gate429inter1, gate429inter2, gate429inter3, gate429inter4, gate429inter5, gate429inter6, gate429inter7, gate429inter8, gate429inter9, gate429inter10, gate429inter11, gate429inter12, gate226inter0, gate226inter1, gate226inter2, gate226inter3, gate226inter4, gate226inter5, gate226inter6, gate226inter7, gate226inter8, gate226inter9, gate226inter10, gate226inter11, gate226inter12, gate41inter0, gate41inter1, gate41inter2, gate41inter3, gate41inter4, gate41inter5, gate41inter6, gate41inter7, gate41inter8, gate41inter9, gate41inter10, gate41inter11, gate41inter12, gate219inter0, gate219inter1, gate219inter2, gate219inter3, gate219inter4, gate219inter5, gate219inter6, gate219inter7, gate219inter8, gate219inter9, gate219inter10, gate219inter11, gate219inter12, gate83inter0, gate83inter1, gate83inter2, gate83inter3, gate83inter4, gate83inter5, gate83inter6, gate83inter7, gate83inter8, gate83inter9, gate83inter10, gate83inter11, gate83inter12, gate107inter0, gate107inter1, gate107inter2, gate107inter3, gate107inter4, gate107inter5, gate107inter6, gate107inter7, gate107inter8, gate107inter9, gate107inter10, gate107inter11, gate107inter12, gate173inter0, gate173inter1, gate173inter2, gate173inter3, gate173inter4, gate173inter5, gate173inter6, gate173inter7, gate173inter8, gate173inter9, gate173inter10, gate173inter11, gate173inter12, gate289inter0, gate289inter1, gate289inter2, gate289inter3, gate289inter4, gate289inter5, gate289inter6, gate289inter7, gate289inter8, gate289inter9, gate289inter10, gate289inter11, gate289inter12, gate192inter0, gate192inter1, gate192inter2, gate192inter3, gate192inter4, gate192inter5, gate192inter6, gate192inter7, gate192inter8, gate192inter9, gate192inter10, gate192inter11, gate192inter12, gate174inter0, gate174inter1, gate174inter2, gate174inter3, gate174inter4, gate174inter5, gate174inter6, gate174inter7, gate174inter8, gate174inter9, gate174inter10, gate174inter11, gate174inter12, gate448inter0, gate448inter1, gate448inter2, gate448inter3, gate448inter4, gate448inter5, gate448inter6, gate448inter7, gate448inter8, gate448inter9, gate448inter10, gate448inter11, gate448inter12, gate170inter0, gate170inter1, gate170inter2, gate170inter3, gate170inter4, gate170inter5, gate170inter6, gate170inter7, gate170inter8, gate170inter9, gate170inter10, gate170inter11, gate170inter12, gate490inter0, gate490inter1, gate490inter2, gate490inter3, gate490inter4, gate490inter5, gate490inter6, gate490inter7, gate490inter8, gate490inter9, gate490inter10, gate490inter11, gate490inter12, gate18inter0, gate18inter1, gate18inter2, gate18inter3, gate18inter4, gate18inter5, gate18inter6, gate18inter7, gate18inter8, gate18inter9, gate18inter10, gate18inter11, gate18inter12, gate483inter0, gate483inter1, gate483inter2, gate483inter3, gate483inter4, gate483inter5, gate483inter6, gate483inter7, gate483inter8, gate483inter9, gate483inter10, gate483inter11, gate483inter12, gate64inter0, gate64inter1, gate64inter2, gate64inter3, gate64inter4, gate64inter5, gate64inter6, gate64inter7, gate64inter8, gate64inter9, gate64inter10, gate64inter11, gate64inter12, gate474inter0, gate474inter1, gate474inter2, gate474inter3, gate474inter4, gate474inter5, gate474inter6, gate474inter7, gate474inter8, gate474inter9, gate474inter10, gate474inter11, gate474inter12, gate93inter0, gate93inter1, gate93inter2, gate93inter3, gate93inter4, gate93inter5, gate93inter6, gate93inter7, gate93inter8, gate93inter9, gate93inter10, gate93inter11, gate93inter12, gate214inter0, gate214inter1, gate214inter2, gate214inter3, gate214inter4, gate214inter5, gate214inter6, gate214inter7, gate214inter8, gate214inter9, gate214inter10, gate214inter11, gate214inter12, gate117inter0, gate117inter1, gate117inter2, gate117inter3, gate117inter4, gate117inter5, gate117inter6, gate117inter7, gate117inter8, gate117inter9, gate117inter10, gate117inter11, gate117inter12, gate12inter0, gate12inter1, gate12inter2, gate12inter3, gate12inter4, gate12inter5, gate12inter6, gate12inter7, gate12inter8, gate12inter9, gate12inter10, gate12inter11, gate12inter12, gate228inter0, gate228inter1, gate228inter2, gate228inter3, gate228inter4, gate228inter5, gate228inter6, gate228inter7, gate228inter8, gate228inter9, gate228inter10, gate228inter11, gate228inter12, gate28inter0, gate28inter1, gate28inter2, gate28inter3, gate28inter4, gate28inter5, gate28inter6, gate28inter7, gate28inter8, gate28inter9, gate28inter10, gate28inter11, gate28inter12, gate488inter0, gate488inter1, gate488inter2, gate488inter3, gate488inter4, gate488inter5, gate488inter6, gate488inter7, gate488inter8, gate488inter9, gate488inter10, gate488inter11, gate488inter12, gate181inter0, gate181inter1, gate181inter2, gate181inter3, gate181inter4, gate181inter5, gate181inter6, gate181inter7, gate181inter8, gate181inter9, gate181inter10, gate181inter11, gate181inter12, gate60inter0, gate60inter1, gate60inter2, gate60inter3, gate60inter4, gate60inter5, gate60inter6, gate60inter7, gate60inter8, gate60inter9, gate60inter10, gate60inter11, gate60inter12, gate413inter0, gate413inter1, gate413inter2, gate413inter3, gate413inter4, gate413inter5, gate413inter6, gate413inter7, gate413inter8, gate413inter9, gate413inter10, gate413inter11, gate413inter12, gate102inter0, gate102inter1, gate102inter2, gate102inter3, gate102inter4, gate102inter5, gate102inter6, gate102inter7, gate102inter8, gate102inter9, gate102inter10, gate102inter11, gate102inter12, gate204inter0, gate204inter1, gate204inter2, gate204inter3, gate204inter4, gate204inter5, gate204inter6, gate204inter7, gate204inter8, gate204inter9, gate204inter10, gate204inter11, gate204inter12, gate36inter0, gate36inter1, gate36inter2, gate36inter3, gate36inter4, gate36inter5, gate36inter6, gate36inter7, gate36inter8, gate36inter9, gate36inter10, gate36inter11, gate36inter12, gate53inter0, gate53inter1, gate53inter2, gate53inter3, gate53inter4, gate53inter5, gate53inter6, gate53inter7, gate53inter8, gate53inter9, gate53inter10, gate53inter11, gate53inter12, gate39inter0, gate39inter1, gate39inter2, gate39inter3, gate39inter4, gate39inter5, gate39inter6, gate39inter7, gate39inter8, gate39inter9, gate39inter10, gate39inter11, gate39inter12, gate255inter0, gate255inter1, gate255inter2, gate255inter3, gate255inter4, gate255inter5, gate255inter6, gate255inter7, gate255inter8, gate255inter9, gate255inter10, gate255inter11, gate255inter12, gate247inter0, gate247inter1, gate247inter2, gate247inter3, gate247inter4, gate247inter5, gate247inter6, gate247inter7, gate247inter8, gate247inter9, gate247inter10, gate247inter11, gate247inter12, gate465inter0, gate465inter1, gate465inter2, gate465inter3, gate465inter4, gate465inter5, gate465inter6, gate465inter7, gate465inter8, gate465inter9, gate465inter10, gate465inter11, gate465inter12, gate275inter0, gate275inter1, gate275inter2, gate275inter3, gate275inter4, gate275inter5, gate275inter6, gate275inter7, gate275inter8, gate275inter9, gate275inter10, gate275inter11, gate275inter12, gate74inter0, gate74inter1, gate74inter2, gate74inter3, gate74inter4, gate74inter5, gate74inter6, gate74inter7, gate74inter8, gate74inter9, gate74inter10, gate74inter11, gate74inter12, gate290inter0, gate290inter1, gate290inter2, gate290inter3, gate290inter4, gate290inter5, gate290inter6, gate290inter7, gate290inter8, gate290inter9, gate290inter10, gate290inter11, gate290inter12, gate410inter0, gate410inter1, gate410inter2, gate410inter3, gate410inter4, gate410inter5, gate410inter6, gate410inter7, gate410inter8, gate410inter9, gate410inter10, gate410inter11, gate410inter12, gate239inter0, gate239inter1, gate239inter2, gate239inter3, gate239inter4, gate239inter5, gate239inter6, gate239inter7, gate239inter8, gate239inter9, gate239inter10, gate239inter11, gate239inter12, gate236inter0, gate236inter1, gate236inter2, gate236inter3, gate236inter4, gate236inter5, gate236inter6, gate236inter7, gate236inter8, gate236inter9, gate236inter10, gate236inter11, gate236inter12, gate21inter0, gate21inter1, gate21inter2, gate21inter3, gate21inter4, gate21inter5, gate21inter6, gate21inter7, gate21inter8, gate21inter9, gate21inter10, gate21inter11, gate21inter12, gate262inter0, gate262inter1, gate262inter2, gate262inter3, gate262inter4, gate262inter5, gate262inter6, gate262inter7, gate262inter8, gate262inter9, gate262inter10, gate262inter11, gate262inter12, gate238inter0, gate238inter1, gate238inter2, gate238inter3, gate238inter4, gate238inter5, gate238inter6, gate238inter7, gate238inter8, gate238inter9, gate238inter10, gate238inter11, gate238inter12, gate464inter0, gate464inter1, gate464inter2, gate464inter3, gate464inter4, gate464inter5, gate464inter6, gate464inter7, gate464inter8, gate464inter9, gate464inter10, gate464inter11, gate464inter12, gate154inter0, gate154inter1, gate154inter2, gate154inter3, gate154inter4, gate154inter5, gate154inter6, gate154inter7, gate154inter8, gate154inter9, gate154inter10, gate154inter11, gate154inter12, gate187inter0, gate187inter1, gate187inter2, gate187inter3, gate187inter4, gate187inter5, gate187inter6, gate187inter7, gate187inter8, gate187inter9, gate187inter10, gate187inter11, gate187inter12, gate251inter0, gate251inter1, gate251inter2, gate251inter3, gate251inter4, gate251inter5, gate251inter6, gate251inter7, gate251inter8, gate251inter9, gate251inter10, gate251inter11, gate251inter12, gate421inter0, gate421inter1, gate421inter2, gate421inter3, gate421inter4, gate421inter5, gate421inter6, gate421inter7, gate421inter8, gate421inter9, gate421inter10, gate421inter11, gate421inter12, gate503inter0, gate503inter1, gate503inter2, gate503inter3, gate503inter4, gate503inter5, gate503inter6, gate503inter7, gate503inter8, gate503inter9, gate503inter10, gate503inter11, gate503inter12, gate268inter0, gate268inter1, gate268inter2, gate268inter3, gate268inter4, gate268inter5, gate268inter6, gate268inter7, gate268inter8, gate268inter9, gate268inter10, gate268inter11, gate268inter12, gate121inter0, gate121inter1, gate121inter2, gate121inter3, gate121inter4, gate121inter5, gate121inter6, gate121inter7, gate121inter8, gate121inter9, gate121inter10, gate121inter11, gate121inter12, gate50inter0, gate50inter1, gate50inter2, gate50inter3, gate50inter4, gate50inter5, gate50inter6, gate50inter7, gate50inter8, gate50inter9, gate50inter10, gate50inter11, gate50inter12, gate114inter0, gate114inter1, gate114inter2, gate114inter3, gate114inter4, gate114inter5, gate114inter6, gate114inter7, gate114inter8, gate114inter9, gate114inter10, gate114inter11, gate114inter12, gate139inter0, gate139inter1, gate139inter2, gate139inter3, gate139inter4, gate139inter5, gate139inter6, gate139inter7, gate139inter8, gate139inter9, gate139inter10, gate139inter11, gate139inter12, gate202inter0, gate202inter1, gate202inter2, gate202inter3, gate202inter4, gate202inter5, gate202inter6, gate202inter7, gate202inter8, gate202inter9, gate202inter10, gate202inter11, gate202inter12, gate48inter0, gate48inter1, gate48inter2, gate48inter3, gate48inter4, gate48inter5, gate48inter6, gate48inter7, gate48inter8, gate48inter9, gate48inter10, gate48inter11, gate48inter12, gate220inter0, gate220inter1, gate220inter2, gate220inter3, gate220inter4, gate220inter5, gate220inter6, gate220inter7, gate220inter8, gate220inter9, gate220inter10, gate220inter11, gate220inter12, gate194inter0, gate194inter1, gate194inter2, gate194inter3, gate194inter4, gate194inter5, gate194inter6, gate194inter7, gate194inter8, gate194inter9, gate194inter10, gate194inter11, gate194inter12, gate453inter0, gate453inter1, gate453inter2, gate453inter3, gate453inter4, gate453inter5, gate453inter6, gate453inter7, gate453inter8, gate453inter9, gate453inter10, gate453inter11, gate453inter12, gate62inter0, gate62inter1, gate62inter2, gate62inter3, gate62inter4, gate62inter5, gate62inter6, gate62inter7, gate62inter8, gate62inter9, gate62inter10, gate62inter11, gate62inter12, gate89inter0, gate89inter1, gate89inter2, gate89inter3, gate89inter4, gate89inter5, gate89inter6, gate89inter7, gate89inter8, gate89inter9, gate89inter10, gate89inter11, gate89inter12, gate241inter0, gate241inter1, gate241inter2, gate241inter3, gate241inter4, gate241inter5, gate241inter6, gate241inter7, gate241inter8, gate241inter9, gate241inter10, gate241inter11, gate241inter12, gate110inter0, gate110inter1, gate110inter2, gate110inter3, gate110inter4, gate110inter5, gate110inter6, gate110inter7, gate110inter8, gate110inter9, gate110inter10, gate110inter11, gate110inter12, gate33inter0, gate33inter1, gate33inter2, gate33inter3, gate33inter4, gate33inter5, gate33inter6, gate33inter7, gate33inter8, gate33inter9, gate33inter10, gate33inter11, gate33inter12, gate286inter0, gate286inter1, gate286inter2, gate286inter3, gate286inter4, gate286inter5, gate286inter6, gate286inter7, gate286inter8, gate286inter9, gate286inter10, gate286inter11, gate286inter12, gate269inter0, gate269inter1, gate269inter2, gate269inter3, gate269inter4, gate269inter5, gate269inter6, gate269inter7, gate269inter8, gate269inter9, gate269inter10, gate269inter11, gate269inter12, gate467inter0, gate467inter1, gate467inter2, gate467inter3, gate467inter4, gate467inter5, gate467inter6, gate467inter7, gate467inter8, gate467inter9, gate467inter10, gate467inter11, gate467inter12, gate505inter0, gate505inter1, gate505inter2, gate505inter3, gate505inter4, gate505inter5, gate505inter6, gate505inter7, gate505inter8, gate505inter9, gate505inter10, gate505inter11, gate505inter12, gate178inter0, gate178inter1, gate178inter2, gate178inter3, gate178inter4, gate178inter5, gate178inter6, gate178inter7, gate178inter8, gate178inter9, gate178inter10, gate178inter11, gate178inter12, gate231inter0, gate231inter1, gate231inter2, gate231inter3, gate231inter4, gate231inter5, gate231inter6, gate231inter7, gate231inter8, gate231inter9, gate231inter10, gate231inter11, gate231inter12, gate245inter0, gate245inter1, gate245inter2, gate245inter3, gate245inter4, gate245inter5, gate245inter6, gate245inter7, gate245inter8, gate245inter9, gate245inter10, gate245inter11, gate245inter12, gate180inter0, gate180inter1, gate180inter2, gate180inter3, gate180inter4, gate180inter5, gate180inter6, gate180inter7, gate180inter8, gate180inter9, gate180inter10, gate180inter11, gate180inter12, gate389inter0, gate389inter1, gate389inter2, gate389inter3, gate389inter4, gate389inter5, gate389inter6, gate389inter7, gate389inter8, gate389inter9, gate389inter10, gate389inter11, gate389inter12, gate160inter0, gate160inter1, gate160inter2, gate160inter3, gate160inter4, gate160inter5, gate160inter6, gate160inter7, gate160inter8, gate160inter9, gate160inter10, gate160inter11, gate160inter12, gate478inter0, gate478inter1, gate478inter2, gate478inter3, gate478inter4, gate478inter5, gate478inter6, gate478inter7, gate478inter8, gate478inter9, gate478inter10, gate478inter11, gate478inter12, gate295inter0, gate295inter1, gate295inter2, gate295inter3, gate295inter4, gate295inter5, gate295inter6, gate295inter7, gate295inter8, gate295inter9, gate295inter10, gate295inter11, gate295inter12, gate218inter0, gate218inter1, gate218inter2, gate218inter3, gate218inter4, gate218inter5, gate218inter6, gate218inter7, gate218inter8, gate218inter9, gate218inter10, gate218inter11, gate218inter12, gate52inter0, gate52inter1, gate52inter2, gate52inter3, gate52inter4, gate52inter5, gate52inter6, gate52inter7, gate52inter8, gate52inter9, gate52inter10, gate52inter11, gate52inter12, gate484inter0, gate484inter1, gate484inter2, gate484inter3, gate484inter4, gate484inter5, gate484inter6, gate484inter7, gate484inter8, gate484inter9, gate484inter10, gate484inter11, gate484inter12, gate19inter0, gate19inter1, gate19inter2, gate19inter3, gate19inter4, gate19inter5, gate19inter6, gate19inter7, gate19inter8, gate19inter9, gate19inter10, gate19inter11, gate19inter12, gate71inter0, gate71inter1, gate71inter2, gate71inter3, gate71inter4, gate71inter5, gate71inter6, gate71inter7, gate71inter8, gate71inter9, gate71inter10, gate71inter11, gate71inter12, gate441inter0, gate441inter1, gate441inter2, gate441inter3, gate441inter4, gate441inter5, gate441inter6, gate441inter7, gate441inter8, gate441inter9, gate441inter10, gate441inter11, gate441inter12, gate182inter0, gate182inter1, gate182inter2, gate182inter3, gate182inter4, gate182inter5, gate182inter6, gate182inter7, gate182inter8, gate182inter9, gate182inter10, gate182inter11, gate182inter12, gate123inter0, gate123inter1, gate123inter2, gate123inter3, gate123inter4, gate123inter5, gate123inter6, gate123inter7, gate123inter8, gate123inter9, gate123inter10, gate123inter11, gate123inter12, gate451inter0, gate451inter1, gate451inter2, gate451inter3, gate451inter4, gate451inter5, gate451inter6, gate451inter7, gate451inter8, gate451inter9, gate451inter10, gate451inter11, gate451inter12, gate460inter0, gate460inter1, gate460inter2, gate460inter3, gate460inter4, gate460inter5, gate460inter6, gate460inter7, gate460inter8, gate460inter9, gate460inter10, gate460inter11, gate460inter12;



and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );
nand2 gate9( .a(G1), .b(G2), .O(G266) );

  xor2  gate799(.a(G4), .b(G3), .O(gate10inter0));
  nand2 gate800(.a(gate10inter0), .b(s_36), .O(gate10inter1));
  and2  gate801(.a(G4), .b(G3), .O(gate10inter2));
  inv1  gate802(.a(s_36), .O(gate10inter3));
  inv1  gate803(.a(s_37), .O(gate10inter4));
  nand2 gate804(.a(gate10inter4), .b(gate10inter3), .O(gate10inter5));
  nor2  gate805(.a(gate10inter5), .b(gate10inter2), .O(gate10inter6));
  inv1  gate806(.a(G3), .O(gate10inter7));
  inv1  gate807(.a(G4), .O(gate10inter8));
  nand2 gate808(.a(gate10inter8), .b(gate10inter7), .O(gate10inter9));
  nand2 gate809(.a(s_37), .b(gate10inter3), .O(gate10inter10));
  nor2  gate810(.a(gate10inter10), .b(gate10inter9), .O(gate10inter11));
  nor2  gate811(.a(gate10inter11), .b(gate10inter6), .O(gate10inter12));
  nand2 gate812(.a(gate10inter12), .b(gate10inter1), .O(G269));
nand2 gate11( .a(G5), .b(G6), .O(G272) );

  xor2  gate1863(.a(G8), .b(G7), .O(gate12inter0));
  nand2 gate1864(.a(gate12inter0), .b(s_188), .O(gate12inter1));
  and2  gate1865(.a(G8), .b(G7), .O(gate12inter2));
  inv1  gate1866(.a(s_188), .O(gate12inter3));
  inv1  gate1867(.a(s_189), .O(gate12inter4));
  nand2 gate1868(.a(gate12inter4), .b(gate12inter3), .O(gate12inter5));
  nor2  gate1869(.a(gate12inter5), .b(gate12inter2), .O(gate12inter6));
  inv1  gate1870(.a(G7), .O(gate12inter7));
  inv1  gate1871(.a(G8), .O(gate12inter8));
  nand2 gate1872(.a(gate12inter8), .b(gate12inter7), .O(gate12inter9));
  nand2 gate1873(.a(s_189), .b(gate12inter3), .O(gate12inter10));
  nor2  gate1874(.a(gate12inter10), .b(gate12inter9), .O(gate12inter11));
  nor2  gate1875(.a(gate12inter11), .b(gate12inter6), .O(gate12inter12));
  nand2 gate1876(.a(gate12inter12), .b(gate12inter1), .O(G275));
nand2 gate13( .a(G9), .b(G10), .O(G278) );
nand2 gate14( .a(G11), .b(G12), .O(G281) );
nand2 gate15( .a(G13), .b(G14), .O(G284) );
nand2 gate16( .a(G15), .b(G16), .O(G287) );
nand2 gate17( .a(G17), .b(G18), .O(G290) );

  xor2  gate1765(.a(G20), .b(G19), .O(gate18inter0));
  nand2 gate1766(.a(gate18inter0), .b(s_174), .O(gate18inter1));
  and2  gate1767(.a(G20), .b(G19), .O(gate18inter2));
  inv1  gate1768(.a(s_174), .O(gate18inter3));
  inv1  gate1769(.a(s_175), .O(gate18inter4));
  nand2 gate1770(.a(gate18inter4), .b(gate18inter3), .O(gate18inter5));
  nor2  gate1771(.a(gate18inter5), .b(gate18inter2), .O(gate18inter6));
  inv1  gate1772(.a(G19), .O(gate18inter7));
  inv1  gate1773(.a(G20), .O(gate18inter8));
  nand2 gate1774(.a(gate18inter8), .b(gate18inter7), .O(gate18inter9));
  nand2 gate1775(.a(s_175), .b(gate18inter3), .O(gate18inter10));
  nor2  gate1776(.a(gate18inter10), .b(gate18inter9), .O(gate18inter11));
  nor2  gate1777(.a(gate18inter11), .b(gate18inter6), .O(gate18inter12));
  nand2 gate1778(.a(gate18inter12), .b(gate18inter1), .O(G293));

  xor2  gate2703(.a(G22), .b(G21), .O(gate19inter0));
  nand2 gate2704(.a(gate19inter0), .b(s_308), .O(gate19inter1));
  and2  gate2705(.a(G22), .b(G21), .O(gate19inter2));
  inv1  gate2706(.a(s_308), .O(gate19inter3));
  inv1  gate2707(.a(s_309), .O(gate19inter4));
  nand2 gate2708(.a(gate19inter4), .b(gate19inter3), .O(gate19inter5));
  nor2  gate2709(.a(gate19inter5), .b(gate19inter2), .O(gate19inter6));
  inv1  gate2710(.a(G21), .O(gate19inter7));
  inv1  gate2711(.a(G22), .O(gate19inter8));
  nand2 gate2712(.a(gate19inter8), .b(gate19inter7), .O(gate19inter9));
  nand2 gate2713(.a(s_309), .b(gate19inter3), .O(gate19inter10));
  nor2  gate2714(.a(gate19inter10), .b(gate19inter9), .O(gate19inter11));
  nor2  gate2715(.a(gate19inter11), .b(gate19inter6), .O(gate19inter12));
  nand2 gate2716(.a(gate19inter12), .b(gate19inter1), .O(G296));
nand2 gate20( .a(G23), .b(G24), .O(G299) );

  xor2  gate2157(.a(G26), .b(G25), .O(gate21inter0));
  nand2 gate2158(.a(gate21inter0), .b(s_230), .O(gate21inter1));
  and2  gate2159(.a(G26), .b(G25), .O(gate21inter2));
  inv1  gate2160(.a(s_230), .O(gate21inter3));
  inv1  gate2161(.a(s_231), .O(gate21inter4));
  nand2 gate2162(.a(gate21inter4), .b(gate21inter3), .O(gate21inter5));
  nor2  gate2163(.a(gate21inter5), .b(gate21inter2), .O(gate21inter6));
  inv1  gate2164(.a(G25), .O(gate21inter7));
  inv1  gate2165(.a(G26), .O(gate21inter8));
  nand2 gate2166(.a(gate21inter8), .b(gate21inter7), .O(gate21inter9));
  nand2 gate2167(.a(s_231), .b(gate21inter3), .O(gate21inter10));
  nor2  gate2168(.a(gate21inter10), .b(gate21inter9), .O(gate21inter11));
  nor2  gate2169(.a(gate21inter11), .b(gate21inter6), .O(gate21inter12));
  nand2 gate2170(.a(gate21inter12), .b(gate21inter1), .O(G302));
nand2 gate22( .a(G27), .b(G28), .O(G305) );
nand2 gate23( .a(G29), .b(G30), .O(G308) );
nand2 gate24( .a(G31), .b(G32), .O(G311) );
nand2 gate25( .a(G1), .b(G5), .O(G314) );
nand2 gate26( .a(G9), .b(G13), .O(G317) );
nand2 gate27( .a(G2), .b(G6), .O(G320) );

  xor2  gate1891(.a(G14), .b(G10), .O(gate28inter0));
  nand2 gate1892(.a(gate28inter0), .b(s_192), .O(gate28inter1));
  and2  gate1893(.a(G14), .b(G10), .O(gate28inter2));
  inv1  gate1894(.a(s_192), .O(gate28inter3));
  inv1  gate1895(.a(s_193), .O(gate28inter4));
  nand2 gate1896(.a(gate28inter4), .b(gate28inter3), .O(gate28inter5));
  nor2  gate1897(.a(gate28inter5), .b(gate28inter2), .O(gate28inter6));
  inv1  gate1898(.a(G10), .O(gate28inter7));
  inv1  gate1899(.a(G14), .O(gate28inter8));
  nand2 gate1900(.a(gate28inter8), .b(gate28inter7), .O(gate28inter9));
  nand2 gate1901(.a(s_193), .b(gate28inter3), .O(gate28inter10));
  nor2  gate1902(.a(gate28inter10), .b(gate28inter9), .O(gate28inter11));
  nor2  gate1903(.a(gate28inter11), .b(gate28inter6), .O(gate28inter12));
  nand2 gate1904(.a(gate28inter12), .b(gate28inter1), .O(G323));
nand2 gate29( .a(G3), .b(G7), .O(G326) );
nand2 gate30( .a(G11), .b(G15), .O(G329) );
nand2 gate31( .a(G4), .b(G8), .O(G332) );

  xor2  gate631(.a(G16), .b(G12), .O(gate32inter0));
  nand2 gate632(.a(gate32inter0), .b(s_12), .O(gate32inter1));
  and2  gate633(.a(G16), .b(G12), .O(gate32inter2));
  inv1  gate634(.a(s_12), .O(gate32inter3));
  inv1  gate635(.a(s_13), .O(gate32inter4));
  nand2 gate636(.a(gate32inter4), .b(gate32inter3), .O(gate32inter5));
  nor2  gate637(.a(gate32inter5), .b(gate32inter2), .O(gate32inter6));
  inv1  gate638(.a(G12), .O(gate32inter7));
  inv1  gate639(.a(G16), .O(gate32inter8));
  nand2 gate640(.a(gate32inter8), .b(gate32inter7), .O(gate32inter9));
  nand2 gate641(.a(s_13), .b(gate32inter3), .O(gate32inter10));
  nor2  gate642(.a(gate32inter10), .b(gate32inter9), .O(gate32inter11));
  nor2  gate643(.a(gate32inter11), .b(gate32inter6), .O(gate32inter12));
  nand2 gate644(.a(gate32inter12), .b(gate32inter1), .O(G335));

  xor2  gate2479(.a(G21), .b(G17), .O(gate33inter0));
  nand2 gate2480(.a(gate33inter0), .b(s_276), .O(gate33inter1));
  and2  gate2481(.a(G21), .b(G17), .O(gate33inter2));
  inv1  gate2482(.a(s_276), .O(gate33inter3));
  inv1  gate2483(.a(s_277), .O(gate33inter4));
  nand2 gate2484(.a(gate33inter4), .b(gate33inter3), .O(gate33inter5));
  nor2  gate2485(.a(gate33inter5), .b(gate33inter2), .O(gate33inter6));
  inv1  gate2486(.a(G17), .O(gate33inter7));
  inv1  gate2487(.a(G21), .O(gate33inter8));
  nand2 gate2488(.a(gate33inter8), .b(gate33inter7), .O(gate33inter9));
  nand2 gate2489(.a(s_277), .b(gate33inter3), .O(gate33inter10));
  nor2  gate2490(.a(gate33inter10), .b(gate33inter9), .O(gate33inter11));
  nor2  gate2491(.a(gate33inter11), .b(gate33inter6), .O(gate33inter12));
  nand2 gate2492(.a(gate33inter12), .b(gate33inter1), .O(G338));
nand2 gate34( .a(G25), .b(G29), .O(G341) );
nand2 gate35( .a(G18), .b(G22), .O(G344) );

  xor2  gate1989(.a(G30), .b(G26), .O(gate36inter0));
  nand2 gate1990(.a(gate36inter0), .b(s_206), .O(gate36inter1));
  and2  gate1991(.a(G30), .b(G26), .O(gate36inter2));
  inv1  gate1992(.a(s_206), .O(gate36inter3));
  inv1  gate1993(.a(s_207), .O(gate36inter4));
  nand2 gate1994(.a(gate36inter4), .b(gate36inter3), .O(gate36inter5));
  nor2  gate1995(.a(gate36inter5), .b(gate36inter2), .O(gate36inter6));
  inv1  gate1996(.a(G26), .O(gate36inter7));
  inv1  gate1997(.a(G30), .O(gate36inter8));
  nand2 gate1998(.a(gate36inter8), .b(gate36inter7), .O(gate36inter9));
  nand2 gate1999(.a(s_207), .b(gate36inter3), .O(gate36inter10));
  nor2  gate2000(.a(gate36inter10), .b(gate36inter9), .O(gate36inter11));
  nor2  gate2001(.a(gate36inter11), .b(gate36inter6), .O(gate36inter12));
  nand2 gate2002(.a(gate36inter12), .b(gate36inter1), .O(G347));
nand2 gate37( .a(G19), .b(G23), .O(G350) );
nand2 gate38( .a(G27), .b(G31), .O(G353) );

  xor2  gate2017(.a(G24), .b(G20), .O(gate39inter0));
  nand2 gate2018(.a(gate39inter0), .b(s_210), .O(gate39inter1));
  and2  gate2019(.a(G24), .b(G20), .O(gate39inter2));
  inv1  gate2020(.a(s_210), .O(gate39inter3));
  inv1  gate2021(.a(s_211), .O(gate39inter4));
  nand2 gate2022(.a(gate39inter4), .b(gate39inter3), .O(gate39inter5));
  nor2  gate2023(.a(gate39inter5), .b(gate39inter2), .O(gate39inter6));
  inv1  gate2024(.a(G20), .O(gate39inter7));
  inv1  gate2025(.a(G24), .O(gate39inter8));
  nand2 gate2026(.a(gate39inter8), .b(gate39inter7), .O(gate39inter9));
  nand2 gate2027(.a(s_211), .b(gate39inter3), .O(gate39inter10));
  nor2  gate2028(.a(gate39inter10), .b(gate39inter9), .O(gate39inter11));
  nor2  gate2029(.a(gate39inter11), .b(gate39inter6), .O(gate39inter12));
  nand2 gate2030(.a(gate39inter12), .b(gate39inter1), .O(G356));
nand2 gate40( .a(G28), .b(G32), .O(G359) );

  xor2  gate1611(.a(G266), .b(G1), .O(gate41inter0));
  nand2 gate1612(.a(gate41inter0), .b(s_152), .O(gate41inter1));
  and2  gate1613(.a(G266), .b(G1), .O(gate41inter2));
  inv1  gate1614(.a(s_152), .O(gate41inter3));
  inv1  gate1615(.a(s_153), .O(gate41inter4));
  nand2 gate1616(.a(gate41inter4), .b(gate41inter3), .O(gate41inter5));
  nor2  gate1617(.a(gate41inter5), .b(gate41inter2), .O(gate41inter6));
  inv1  gate1618(.a(G1), .O(gate41inter7));
  inv1  gate1619(.a(G266), .O(gate41inter8));
  nand2 gate1620(.a(gate41inter8), .b(gate41inter7), .O(gate41inter9));
  nand2 gate1621(.a(s_153), .b(gate41inter3), .O(gate41inter10));
  nor2  gate1622(.a(gate41inter10), .b(gate41inter9), .O(gate41inter11));
  nor2  gate1623(.a(gate41inter11), .b(gate41inter6), .O(gate41inter12));
  nand2 gate1624(.a(gate41inter12), .b(gate41inter1), .O(G362));
nand2 gate42( .a(G2), .b(G266), .O(G363) );

  xor2  gate603(.a(G269), .b(G3), .O(gate43inter0));
  nand2 gate604(.a(gate43inter0), .b(s_8), .O(gate43inter1));
  and2  gate605(.a(G269), .b(G3), .O(gate43inter2));
  inv1  gate606(.a(s_8), .O(gate43inter3));
  inv1  gate607(.a(s_9), .O(gate43inter4));
  nand2 gate608(.a(gate43inter4), .b(gate43inter3), .O(gate43inter5));
  nor2  gate609(.a(gate43inter5), .b(gate43inter2), .O(gate43inter6));
  inv1  gate610(.a(G3), .O(gate43inter7));
  inv1  gate611(.a(G269), .O(gate43inter8));
  nand2 gate612(.a(gate43inter8), .b(gate43inter7), .O(gate43inter9));
  nand2 gate613(.a(s_9), .b(gate43inter3), .O(gate43inter10));
  nor2  gate614(.a(gate43inter10), .b(gate43inter9), .O(gate43inter11));
  nor2  gate615(.a(gate43inter11), .b(gate43inter6), .O(gate43inter12));
  nand2 gate616(.a(gate43inter12), .b(gate43inter1), .O(G364));

  xor2  gate1177(.a(G269), .b(G4), .O(gate44inter0));
  nand2 gate1178(.a(gate44inter0), .b(s_90), .O(gate44inter1));
  and2  gate1179(.a(G269), .b(G4), .O(gate44inter2));
  inv1  gate1180(.a(s_90), .O(gate44inter3));
  inv1  gate1181(.a(s_91), .O(gate44inter4));
  nand2 gate1182(.a(gate44inter4), .b(gate44inter3), .O(gate44inter5));
  nor2  gate1183(.a(gate44inter5), .b(gate44inter2), .O(gate44inter6));
  inv1  gate1184(.a(G4), .O(gate44inter7));
  inv1  gate1185(.a(G269), .O(gate44inter8));
  nand2 gate1186(.a(gate44inter8), .b(gate44inter7), .O(gate44inter9));
  nand2 gate1187(.a(s_91), .b(gate44inter3), .O(gate44inter10));
  nor2  gate1188(.a(gate44inter10), .b(gate44inter9), .O(gate44inter11));
  nor2  gate1189(.a(gate44inter11), .b(gate44inter6), .O(gate44inter12));
  nand2 gate1190(.a(gate44inter12), .b(gate44inter1), .O(G365));
nand2 gate45( .a(G5), .b(G272), .O(G366) );

  xor2  gate743(.a(G272), .b(G6), .O(gate46inter0));
  nand2 gate744(.a(gate46inter0), .b(s_28), .O(gate46inter1));
  and2  gate745(.a(G272), .b(G6), .O(gate46inter2));
  inv1  gate746(.a(s_28), .O(gate46inter3));
  inv1  gate747(.a(s_29), .O(gate46inter4));
  nand2 gate748(.a(gate46inter4), .b(gate46inter3), .O(gate46inter5));
  nor2  gate749(.a(gate46inter5), .b(gate46inter2), .O(gate46inter6));
  inv1  gate750(.a(G6), .O(gate46inter7));
  inv1  gate751(.a(G272), .O(gate46inter8));
  nand2 gate752(.a(gate46inter8), .b(gate46inter7), .O(gate46inter9));
  nand2 gate753(.a(s_29), .b(gate46inter3), .O(gate46inter10));
  nor2  gate754(.a(gate46inter10), .b(gate46inter9), .O(gate46inter11));
  nor2  gate755(.a(gate46inter11), .b(gate46inter6), .O(gate46inter12));
  nand2 gate756(.a(gate46inter12), .b(gate46inter1), .O(G367));
nand2 gate47( .a(G7), .b(G275), .O(G368) );

  xor2  gate2367(.a(G275), .b(G8), .O(gate48inter0));
  nand2 gate2368(.a(gate48inter0), .b(s_260), .O(gate48inter1));
  and2  gate2369(.a(G275), .b(G8), .O(gate48inter2));
  inv1  gate2370(.a(s_260), .O(gate48inter3));
  inv1  gate2371(.a(s_261), .O(gate48inter4));
  nand2 gate2372(.a(gate48inter4), .b(gate48inter3), .O(gate48inter5));
  nor2  gate2373(.a(gate48inter5), .b(gate48inter2), .O(gate48inter6));
  inv1  gate2374(.a(G8), .O(gate48inter7));
  inv1  gate2375(.a(G275), .O(gate48inter8));
  nand2 gate2376(.a(gate48inter8), .b(gate48inter7), .O(gate48inter9));
  nand2 gate2377(.a(s_261), .b(gate48inter3), .O(gate48inter10));
  nor2  gate2378(.a(gate48inter10), .b(gate48inter9), .O(gate48inter11));
  nor2  gate2379(.a(gate48inter11), .b(gate48inter6), .O(gate48inter12));
  nand2 gate2380(.a(gate48inter12), .b(gate48inter1), .O(G369));

  xor2  gate1037(.a(G278), .b(G9), .O(gate49inter0));
  nand2 gate1038(.a(gate49inter0), .b(s_70), .O(gate49inter1));
  and2  gate1039(.a(G278), .b(G9), .O(gate49inter2));
  inv1  gate1040(.a(s_70), .O(gate49inter3));
  inv1  gate1041(.a(s_71), .O(gate49inter4));
  nand2 gate1042(.a(gate49inter4), .b(gate49inter3), .O(gate49inter5));
  nor2  gate1043(.a(gate49inter5), .b(gate49inter2), .O(gate49inter6));
  inv1  gate1044(.a(G9), .O(gate49inter7));
  inv1  gate1045(.a(G278), .O(gate49inter8));
  nand2 gate1046(.a(gate49inter8), .b(gate49inter7), .O(gate49inter9));
  nand2 gate1047(.a(s_71), .b(gate49inter3), .O(gate49inter10));
  nor2  gate1048(.a(gate49inter10), .b(gate49inter9), .O(gate49inter11));
  nor2  gate1049(.a(gate49inter11), .b(gate49inter6), .O(gate49inter12));
  nand2 gate1050(.a(gate49inter12), .b(gate49inter1), .O(G370));

  xor2  gate2311(.a(G278), .b(G10), .O(gate50inter0));
  nand2 gate2312(.a(gate50inter0), .b(s_252), .O(gate50inter1));
  and2  gate2313(.a(G278), .b(G10), .O(gate50inter2));
  inv1  gate2314(.a(s_252), .O(gate50inter3));
  inv1  gate2315(.a(s_253), .O(gate50inter4));
  nand2 gate2316(.a(gate50inter4), .b(gate50inter3), .O(gate50inter5));
  nor2  gate2317(.a(gate50inter5), .b(gate50inter2), .O(gate50inter6));
  inv1  gate2318(.a(G10), .O(gate50inter7));
  inv1  gate2319(.a(G278), .O(gate50inter8));
  nand2 gate2320(.a(gate50inter8), .b(gate50inter7), .O(gate50inter9));
  nand2 gate2321(.a(s_253), .b(gate50inter3), .O(gate50inter10));
  nor2  gate2322(.a(gate50inter10), .b(gate50inter9), .O(gate50inter11));
  nor2  gate2323(.a(gate50inter11), .b(gate50inter6), .O(gate50inter12));
  nand2 gate2324(.a(gate50inter12), .b(gate50inter1), .O(G371));
nand2 gate51( .a(G11), .b(G281), .O(G372) );

  xor2  gate2675(.a(G281), .b(G12), .O(gate52inter0));
  nand2 gate2676(.a(gate52inter0), .b(s_304), .O(gate52inter1));
  and2  gate2677(.a(G281), .b(G12), .O(gate52inter2));
  inv1  gate2678(.a(s_304), .O(gate52inter3));
  inv1  gate2679(.a(s_305), .O(gate52inter4));
  nand2 gate2680(.a(gate52inter4), .b(gate52inter3), .O(gate52inter5));
  nor2  gate2681(.a(gate52inter5), .b(gate52inter2), .O(gate52inter6));
  inv1  gate2682(.a(G12), .O(gate52inter7));
  inv1  gate2683(.a(G281), .O(gate52inter8));
  nand2 gate2684(.a(gate52inter8), .b(gate52inter7), .O(gate52inter9));
  nand2 gate2685(.a(s_305), .b(gate52inter3), .O(gate52inter10));
  nor2  gate2686(.a(gate52inter10), .b(gate52inter9), .O(gate52inter11));
  nor2  gate2687(.a(gate52inter11), .b(gate52inter6), .O(gate52inter12));
  nand2 gate2688(.a(gate52inter12), .b(gate52inter1), .O(G373));

  xor2  gate2003(.a(G284), .b(G13), .O(gate53inter0));
  nand2 gate2004(.a(gate53inter0), .b(s_208), .O(gate53inter1));
  and2  gate2005(.a(G284), .b(G13), .O(gate53inter2));
  inv1  gate2006(.a(s_208), .O(gate53inter3));
  inv1  gate2007(.a(s_209), .O(gate53inter4));
  nand2 gate2008(.a(gate53inter4), .b(gate53inter3), .O(gate53inter5));
  nor2  gate2009(.a(gate53inter5), .b(gate53inter2), .O(gate53inter6));
  inv1  gate2010(.a(G13), .O(gate53inter7));
  inv1  gate2011(.a(G284), .O(gate53inter8));
  nand2 gate2012(.a(gate53inter8), .b(gate53inter7), .O(gate53inter9));
  nand2 gate2013(.a(s_209), .b(gate53inter3), .O(gate53inter10));
  nor2  gate2014(.a(gate53inter10), .b(gate53inter9), .O(gate53inter11));
  nor2  gate2015(.a(gate53inter11), .b(gate53inter6), .O(gate53inter12));
  nand2 gate2016(.a(gate53inter12), .b(gate53inter1), .O(G374));
nand2 gate54( .a(G14), .b(G284), .O(G375) );
nand2 gate55( .a(G15), .b(G287), .O(G376) );
nand2 gate56( .a(G16), .b(G287), .O(G377) );
nand2 gate57( .a(G17), .b(G290), .O(G378) );
nand2 gate58( .a(G18), .b(G290), .O(G379) );
nand2 gate59( .a(G19), .b(G293), .O(G380) );

  xor2  gate1933(.a(G293), .b(G20), .O(gate60inter0));
  nand2 gate1934(.a(gate60inter0), .b(s_198), .O(gate60inter1));
  and2  gate1935(.a(G293), .b(G20), .O(gate60inter2));
  inv1  gate1936(.a(s_198), .O(gate60inter3));
  inv1  gate1937(.a(s_199), .O(gate60inter4));
  nand2 gate1938(.a(gate60inter4), .b(gate60inter3), .O(gate60inter5));
  nor2  gate1939(.a(gate60inter5), .b(gate60inter2), .O(gate60inter6));
  inv1  gate1940(.a(G20), .O(gate60inter7));
  inv1  gate1941(.a(G293), .O(gate60inter8));
  nand2 gate1942(.a(gate60inter8), .b(gate60inter7), .O(gate60inter9));
  nand2 gate1943(.a(s_199), .b(gate60inter3), .O(gate60inter10));
  nor2  gate1944(.a(gate60inter10), .b(gate60inter9), .O(gate60inter11));
  nor2  gate1945(.a(gate60inter11), .b(gate60inter6), .O(gate60inter12));
  nand2 gate1946(.a(gate60inter12), .b(gate60inter1), .O(G381));
nand2 gate61( .a(G21), .b(G296), .O(G382) );

  xor2  gate2423(.a(G296), .b(G22), .O(gate62inter0));
  nand2 gate2424(.a(gate62inter0), .b(s_268), .O(gate62inter1));
  and2  gate2425(.a(G296), .b(G22), .O(gate62inter2));
  inv1  gate2426(.a(s_268), .O(gate62inter3));
  inv1  gate2427(.a(s_269), .O(gate62inter4));
  nand2 gate2428(.a(gate62inter4), .b(gate62inter3), .O(gate62inter5));
  nor2  gate2429(.a(gate62inter5), .b(gate62inter2), .O(gate62inter6));
  inv1  gate2430(.a(G22), .O(gate62inter7));
  inv1  gate2431(.a(G296), .O(gate62inter8));
  nand2 gate2432(.a(gate62inter8), .b(gate62inter7), .O(gate62inter9));
  nand2 gate2433(.a(s_269), .b(gate62inter3), .O(gate62inter10));
  nor2  gate2434(.a(gate62inter10), .b(gate62inter9), .O(gate62inter11));
  nor2  gate2435(.a(gate62inter11), .b(gate62inter6), .O(gate62inter12));
  nand2 gate2436(.a(gate62inter12), .b(gate62inter1), .O(G383));

  xor2  gate1345(.a(G299), .b(G23), .O(gate63inter0));
  nand2 gate1346(.a(gate63inter0), .b(s_114), .O(gate63inter1));
  and2  gate1347(.a(G299), .b(G23), .O(gate63inter2));
  inv1  gate1348(.a(s_114), .O(gate63inter3));
  inv1  gate1349(.a(s_115), .O(gate63inter4));
  nand2 gate1350(.a(gate63inter4), .b(gate63inter3), .O(gate63inter5));
  nor2  gate1351(.a(gate63inter5), .b(gate63inter2), .O(gate63inter6));
  inv1  gate1352(.a(G23), .O(gate63inter7));
  inv1  gate1353(.a(G299), .O(gate63inter8));
  nand2 gate1354(.a(gate63inter8), .b(gate63inter7), .O(gate63inter9));
  nand2 gate1355(.a(s_115), .b(gate63inter3), .O(gate63inter10));
  nor2  gate1356(.a(gate63inter10), .b(gate63inter9), .O(gate63inter11));
  nor2  gate1357(.a(gate63inter11), .b(gate63inter6), .O(gate63inter12));
  nand2 gate1358(.a(gate63inter12), .b(gate63inter1), .O(G384));

  xor2  gate1793(.a(G299), .b(G24), .O(gate64inter0));
  nand2 gate1794(.a(gate64inter0), .b(s_178), .O(gate64inter1));
  and2  gate1795(.a(G299), .b(G24), .O(gate64inter2));
  inv1  gate1796(.a(s_178), .O(gate64inter3));
  inv1  gate1797(.a(s_179), .O(gate64inter4));
  nand2 gate1798(.a(gate64inter4), .b(gate64inter3), .O(gate64inter5));
  nor2  gate1799(.a(gate64inter5), .b(gate64inter2), .O(gate64inter6));
  inv1  gate1800(.a(G24), .O(gate64inter7));
  inv1  gate1801(.a(G299), .O(gate64inter8));
  nand2 gate1802(.a(gate64inter8), .b(gate64inter7), .O(gate64inter9));
  nand2 gate1803(.a(s_179), .b(gate64inter3), .O(gate64inter10));
  nor2  gate1804(.a(gate64inter10), .b(gate64inter9), .O(gate64inter11));
  nor2  gate1805(.a(gate64inter11), .b(gate64inter6), .O(gate64inter12));
  nand2 gate1806(.a(gate64inter12), .b(gate64inter1), .O(G385));
nand2 gate65( .a(G25), .b(G302), .O(G386) );
nand2 gate66( .a(G26), .b(G302), .O(G387) );
nand2 gate67( .a(G27), .b(G305), .O(G388) );
nand2 gate68( .a(G28), .b(G305), .O(G389) );
nand2 gate69( .a(G29), .b(G308), .O(G390) );
nand2 gate70( .a(G30), .b(G308), .O(G391) );

  xor2  gate2717(.a(G311), .b(G31), .O(gate71inter0));
  nand2 gate2718(.a(gate71inter0), .b(s_310), .O(gate71inter1));
  and2  gate2719(.a(G311), .b(G31), .O(gate71inter2));
  inv1  gate2720(.a(s_310), .O(gate71inter3));
  inv1  gate2721(.a(s_311), .O(gate71inter4));
  nand2 gate2722(.a(gate71inter4), .b(gate71inter3), .O(gate71inter5));
  nor2  gate2723(.a(gate71inter5), .b(gate71inter2), .O(gate71inter6));
  inv1  gate2724(.a(G31), .O(gate71inter7));
  inv1  gate2725(.a(G311), .O(gate71inter8));
  nand2 gate2726(.a(gate71inter8), .b(gate71inter7), .O(gate71inter9));
  nand2 gate2727(.a(s_311), .b(gate71inter3), .O(gate71inter10));
  nor2  gate2728(.a(gate71inter10), .b(gate71inter9), .O(gate71inter11));
  nor2  gate2729(.a(gate71inter11), .b(gate71inter6), .O(gate71inter12));
  nand2 gate2730(.a(gate71inter12), .b(gate71inter1), .O(G392));
nand2 gate72( .a(G32), .b(G311), .O(G393) );
nand2 gate73( .a(G1), .b(G314), .O(G394) );

  xor2  gate2087(.a(G314), .b(G5), .O(gate74inter0));
  nand2 gate2088(.a(gate74inter0), .b(s_220), .O(gate74inter1));
  and2  gate2089(.a(G314), .b(G5), .O(gate74inter2));
  inv1  gate2090(.a(s_220), .O(gate74inter3));
  inv1  gate2091(.a(s_221), .O(gate74inter4));
  nand2 gate2092(.a(gate74inter4), .b(gate74inter3), .O(gate74inter5));
  nor2  gate2093(.a(gate74inter5), .b(gate74inter2), .O(gate74inter6));
  inv1  gate2094(.a(G5), .O(gate74inter7));
  inv1  gate2095(.a(G314), .O(gate74inter8));
  nand2 gate2096(.a(gate74inter8), .b(gate74inter7), .O(gate74inter9));
  nand2 gate2097(.a(s_221), .b(gate74inter3), .O(gate74inter10));
  nor2  gate2098(.a(gate74inter10), .b(gate74inter9), .O(gate74inter11));
  nor2  gate2099(.a(gate74inter11), .b(gate74inter6), .O(gate74inter12));
  nand2 gate2100(.a(gate74inter12), .b(gate74inter1), .O(G395));

  xor2  gate687(.a(G317), .b(G9), .O(gate75inter0));
  nand2 gate688(.a(gate75inter0), .b(s_20), .O(gate75inter1));
  and2  gate689(.a(G317), .b(G9), .O(gate75inter2));
  inv1  gate690(.a(s_20), .O(gate75inter3));
  inv1  gate691(.a(s_21), .O(gate75inter4));
  nand2 gate692(.a(gate75inter4), .b(gate75inter3), .O(gate75inter5));
  nor2  gate693(.a(gate75inter5), .b(gate75inter2), .O(gate75inter6));
  inv1  gate694(.a(G9), .O(gate75inter7));
  inv1  gate695(.a(G317), .O(gate75inter8));
  nand2 gate696(.a(gate75inter8), .b(gate75inter7), .O(gate75inter9));
  nand2 gate697(.a(s_21), .b(gate75inter3), .O(gate75inter10));
  nor2  gate698(.a(gate75inter10), .b(gate75inter9), .O(gate75inter11));
  nor2  gate699(.a(gate75inter11), .b(gate75inter6), .O(gate75inter12));
  nand2 gate700(.a(gate75inter12), .b(gate75inter1), .O(G396));
nand2 gate76( .a(G13), .b(G317), .O(G397) );
nand2 gate77( .a(G2), .b(G320), .O(G398) );
nand2 gate78( .a(G6), .b(G320), .O(G399) );
nand2 gate79( .a(G10), .b(G323), .O(G400) );
nand2 gate80( .a(G14), .b(G323), .O(G401) );
nand2 gate81( .a(G3), .b(G326), .O(G402) );
nand2 gate82( .a(G7), .b(G326), .O(G403) );

  xor2  gate1639(.a(G329), .b(G11), .O(gate83inter0));
  nand2 gate1640(.a(gate83inter0), .b(s_156), .O(gate83inter1));
  and2  gate1641(.a(G329), .b(G11), .O(gate83inter2));
  inv1  gate1642(.a(s_156), .O(gate83inter3));
  inv1  gate1643(.a(s_157), .O(gate83inter4));
  nand2 gate1644(.a(gate83inter4), .b(gate83inter3), .O(gate83inter5));
  nor2  gate1645(.a(gate83inter5), .b(gate83inter2), .O(gate83inter6));
  inv1  gate1646(.a(G11), .O(gate83inter7));
  inv1  gate1647(.a(G329), .O(gate83inter8));
  nand2 gate1648(.a(gate83inter8), .b(gate83inter7), .O(gate83inter9));
  nand2 gate1649(.a(s_157), .b(gate83inter3), .O(gate83inter10));
  nor2  gate1650(.a(gate83inter10), .b(gate83inter9), .O(gate83inter11));
  nor2  gate1651(.a(gate83inter11), .b(gate83inter6), .O(gate83inter12));
  nand2 gate1652(.a(gate83inter12), .b(gate83inter1), .O(G404));
nand2 gate84( .a(G15), .b(G329), .O(G405) );

  xor2  gate925(.a(G332), .b(G4), .O(gate85inter0));
  nand2 gate926(.a(gate85inter0), .b(s_54), .O(gate85inter1));
  and2  gate927(.a(G332), .b(G4), .O(gate85inter2));
  inv1  gate928(.a(s_54), .O(gate85inter3));
  inv1  gate929(.a(s_55), .O(gate85inter4));
  nand2 gate930(.a(gate85inter4), .b(gate85inter3), .O(gate85inter5));
  nor2  gate931(.a(gate85inter5), .b(gate85inter2), .O(gate85inter6));
  inv1  gate932(.a(G4), .O(gate85inter7));
  inv1  gate933(.a(G332), .O(gate85inter8));
  nand2 gate934(.a(gate85inter8), .b(gate85inter7), .O(gate85inter9));
  nand2 gate935(.a(s_55), .b(gate85inter3), .O(gate85inter10));
  nor2  gate936(.a(gate85inter10), .b(gate85inter9), .O(gate85inter11));
  nor2  gate937(.a(gate85inter11), .b(gate85inter6), .O(gate85inter12));
  nand2 gate938(.a(gate85inter12), .b(gate85inter1), .O(G406));
nand2 gate86( .a(G8), .b(G332), .O(G407) );
nand2 gate87( .a(G12), .b(G335), .O(G408) );
nand2 gate88( .a(G16), .b(G335), .O(G409) );

  xor2  gate2437(.a(G338), .b(G17), .O(gate89inter0));
  nand2 gate2438(.a(gate89inter0), .b(s_270), .O(gate89inter1));
  and2  gate2439(.a(G338), .b(G17), .O(gate89inter2));
  inv1  gate2440(.a(s_270), .O(gate89inter3));
  inv1  gate2441(.a(s_271), .O(gate89inter4));
  nand2 gate2442(.a(gate89inter4), .b(gate89inter3), .O(gate89inter5));
  nor2  gate2443(.a(gate89inter5), .b(gate89inter2), .O(gate89inter6));
  inv1  gate2444(.a(G17), .O(gate89inter7));
  inv1  gate2445(.a(G338), .O(gate89inter8));
  nand2 gate2446(.a(gate89inter8), .b(gate89inter7), .O(gate89inter9));
  nand2 gate2447(.a(s_271), .b(gate89inter3), .O(gate89inter10));
  nor2  gate2448(.a(gate89inter10), .b(gate89inter9), .O(gate89inter11));
  nor2  gate2449(.a(gate89inter11), .b(gate89inter6), .O(gate89inter12));
  nand2 gate2450(.a(gate89inter12), .b(gate89inter1), .O(G410));
nand2 gate90( .a(G21), .b(G338), .O(G411) );
nand2 gate91( .a(G25), .b(G341), .O(G412) );
nand2 gate92( .a(G29), .b(G341), .O(G413) );

  xor2  gate1821(.a(G344), .b(G18), .O(gate93inter0));
  nand2 gate1822(.a(gate93inter0), .b(s_182), .O(gate93inter1));
  and2  gate1823(.a(G344), .b(G18), .O(gate93inter2));
  inv1  gate1824(.a(s_182), .O(gate93inter3));
  inv1  gate1825(.a(s_183), .O(gate93inter4));
  nand2 gate1826(.a(gate93inter4), .b(gate93inter3), .O(gate93inter5));
  nor2  gate1827(.a(gate93inter5), .b(gate93inter2), .O(gate93inter6));
  inv1  gate1828(.a(G18), .O(gate93inter7));
  inv1  gate1829(.a(G344), .O(gate93inter8));
  nand2 gate1830(.a(gate93inter8), .b(gate93inter7), .O(gate93inter9));
  nand2 gate1831(.a(s_183), .b(gate93inter3), .O(gate93inter10));
  nor2  gate1832(.a(gate93inter10), .b(gate93inter9), .O(gate93inter11));
  nor2  gate1833(.a(gate93inter11), .b(gate93inter6), .O(gate93inter12));
  nand2 gate1834(.a(gate93inter12), .b(gate93inter1), .O(G414));

  xor2  gate1233(.a(G344), .b(G22), .O(gate94inter0));
  nand2 gate1234(.a(gate94inter0), .b(s_98), .O(gate94inter1));
  and2  gate1235(.a(G344), .b(G22), .O(gate94inter2));
  inv1  gate1236(.a(s_98), .O(gate94inter3));
  inv1  gate1237(.a(s_99), .O(gate94inter4));
  nand2 gate1238(.a(gate94inter4), .b(gate94inter3), .O(gate94inter5));
  nor2  gate1239(.a(gate94inter5), .b(gate94inter2), .O(gate94inter6));
  inv1  gate1240(.a(G22), .O(gate94inter7));
  inv1  gate1241(.a(G344), .O(gate94inter8));
  nand2 gate1242(.a(gate94inter8), .b(gate94inter7), .O(gate94inter9));
  nand2 gate1243(.a(s_99), .b(gate94inter3), .O(gate94inter10));
  nor2  gate1244(.a(gate94inter10), .b(gate94inter9), .O(gate94inter11));
  nor2  gate1245(.a(gate94inter11), .b(gate94inter6), .O(gate94inter12));
  nand2 gate1246(.a(gate94inter12), .b(gate94inter1), .O(G415));
nand2 gate95( .a(G26), .b(G347), .O(G416) );
nand2 gate96( .a(G30), .b(G347), .O(G417) );
nand2 gate97( .a(G19), .b(G350), .O(G418) );
nand2 gate98( .a(G23), .b(G350), .O(G419) );
nand2 gate99( .a(G27), .b(G353), .O(G420) );
nand2 gate100( .a(G31), .b(G353), .O(G421) );
nand2 gate101( .a(G20), .b(G356), .O(G422) );

  xor2  gate1961(.a(G356), .b(G24), .O(gate102inter0));
  nand2 gate1962(.a(gate102inter0), .b(s_202), .O(gate102inter1));
  and2  gate1963(.a(G356), .b(G24), .O(gate102inter2));
  inv1  gate1964(.a(s_202), .O(gate102inter3));
  inv1  gate1965(.a(s_203), .O(gate102inter4));
  nand2 gate1966(.a(gate102inter4), .b(gate102inter3), .O(gate102inter5));
  nor2  gate1967(.a(gate102inter5), .b(gate102inter2), .O(gate102inter6));
  inv1  gate1968(.a(G24), .O(gate102inter7));
  inv1  gate1969(.a(G356), .O(gate102inter8));
  nand2 gate1970(.a(gate102inter8), .b(gate102inter7), .O(gate102inter9));
  nand2 gate1971(.a(s_203), .b(gate102inter3), .O(gate102inter10));
  nor2  gate1972(.a(gate102inter10), .b(gate102inter9), .O(gate102inter11));
  nor2  gate1973(.a(gate102inter11), .b(gate102inter6), .O(gate102inter12));
  nand2 gate1974(.a(gate102inter12), .b(gate102inter1), .O(G423));
nand2 gate103( .a(G28), .b(G359), .O(G424) );

  xor2  gate645(.a(G359), .b(G32), .O(gate104inter0));
  nand2 gate646(.a(gate104inter0), .b(s_14), .O(gate104inter1));
  and2  gate647(.a(G359), .b(G32), .O(gate104inter2));
  inv1  gate648(.a(s_14), .O(gate104inter3));
  inv1  gate649(.a(s_15), .O(gate104inter4));
  nand2 gate650(.a(gate104inter4), .b(gate104inter3), .O(gate104inter5));
  nor2  gate651(.a(gate104inter5), .b(gate104inter2), .O(gate104inter6));
  inv1  gate652(.a(G32), .O(gate104inter7));
  inv1  gate653(.a(G359), .O(gate104inter8));
  nand2 gate654(.a(gate104inter8), .b(gate104inter7), .O(gate104inter9));
  nand2 gate655(.a(s_15), .b(gate104inter3), .O(gate104inter10));
  nor2  gate656(.a(gate104inter10), .b(gate104inter9), .O(gate104inter11));
  nor2  gate657(.a(gate104inter11), .b(gate104inter6), .O(gate104inter12));
  nand2 gate658(.a(gate104inter12), .b(gate104inter1), .O(G425));
nand2 gate105( .a(G362), .b(G363), .O(G426) );
nand2 gate106( .a(G364), .b(G365), .O(G429) );

  xor2  gate1653(.a(G367), .b(G366), .O(gate107inter0));
  nand2 gate1654(.a(gate107inter0), .b(s_158), .O(gate107inter1));
  and2  gate1655(.a(G367), .b(G366), .O(gate107inter2));
  inv1  gate1656(.a(s_158), .O(gate107inter3));
  inv1  gate1657(.a(s_159), .O(gate107inter4));
  nand2 gate1658(.a(gate107inter4), .b(gate107inter3), .O(gate107inter5));
  nor2  gate1659(.a(gate107inter5), .b(gate107inter2), .O(gate107inter6));
  inv1  gate1660(.a(G366), .O(gate107inter7));
  inv1  gate1661(.a(G367), .O(gate107inter8));
  nand2 gate1662(.a(gate107inter8), .b(gate107inter7), .O(gate107inter9));
  nand2 gate1663(.a(s_159), .b(gate107inter3), .O(gate107inter10));
  nor2  gate1664(.a(gate107inter10), .b(gate107inter9), .O(gate107inter11));
  nor2  gate1665(.a(gate107inter11), .b(gate107inter6), .O(gate107inter12));
  nand2 gate1666(.a(gate107inter12), .b(gate107inter1), .O(G432));
nand2 gate108( .a(G368), .b(G369), .O(G435) );
nand2 gate109( .a(G370), .b(G371), .O(G438) );

  xor2  gate2465(.a(G373), .b(G372), .O(gate110inter0));
  nand2 gate2466(.a(gate110inter0), .b(s_274), .O(gate110inter1));
  and2  gate2467(.a(G373), .b(G372), .O(gate110inter2));
  inv1  gate2468(.a(s_274), .O(gate110inter3));
  inv1  gate2469(.a(s_275), .O(gate110inter4));
  nand2 gate2470(.a(gate110inter4), .b(gate110inter3), .O(gate110inter5));
  nor2  gate2471(.a(gate110inter5), .b(gate110inter2), .O(gate110inter6));
  inv1  gate2472(.a(G372), .O(gate110inter7));
  inv1  gate2473(.a(G373), .O(gate110inter8));
  nand2 gate2474(.a(gate110inter8), .b(gate110inter7), .O(gate110inter9));
  nand2 gate2475(.a(s_275), .b(gate110inter3), .O(gate110inter10));
  nor2  gate2476(.a(gate110inter10), .b(gate110inter9), .O(gate110inter11));
  nor2  gate2477(.a(gate110inter11), .b(gate110inter6), .O(gate110inter12));
  nand2 gate2478(.a(gate110inter12), .b(gate110inter1), .O(G441));
nand2 gate111( .a(G374), .b(G375), .O(G444) );

  xor2  gate715(.a(G377), .b(G376), .O(gate112inter0));
  nand2 gate716(.a(gate112inter0), .b(s_24), .O(gate112inter1));
  and2  gate717(.a(G377), .b(G376), .O(gate112inter2));
  inv1  gate718(.a(s_24), .O(gate112inter3));
  inv1  gate719(.a(s_25), .O(gate112inter4));
  nand2 gate720(.a(gate112inter4), .b(gate112inter3), .O(gate112inter5));
  nor2  gate721(.a(gate112inter5), .b(gate112inter2), .O(gate112inter6));
  inv1  gate722(.a(G376), .O(gate112inter7));
  inv1  gate723(.a(G377), .O(gate112inter8));
  nand2 gate724(.a(gate112inter8), .b(gate112inter7), .O(gate112inter9));
  nand2 gate725(.a(s_25), .b(gate112inter3), .O(gate112inter10));
  nor2  gate726(.a(gate112inter10), .b(gate112inter9), .O(gate112inter11));
  nor2  gate727(.a(gate112inter11), .b(gate112inter6), .O(gate112inter12));
  nand2 gate728(.a(gate112inter12), .b(gate112inter1), .O(G447));
nand2 gate113( .a(G378), .b(G379), .O(G450) );

  xor2  gate2325(.a(G381), .b(G380), .O(gate114inter0));
  nand2 gate2326(.a(gate114inter0), .b(s_254), .O(gate114inter1));
  and2  gate2327(.a(G381), .b(G380), .O(gate114inter2));
  inv1  gate2328(.a(s_254), .O(gate114inter3));
  inv1  gate2329(.a(s_255), .O(gate114inter4));
  nand2 gate2330(.a(gate114inter4), .b(gate114inter3), .O(gate114inter5));
  nor2  gate2331(.a(gate114inter5), .b(gate114inter2), .O(gate114inter6));
  inv1  gate2332(.a(G380), .O(gate114inter7));
  inv1  gate2333(.a(G381), .O(gate114inter8));
  nand2 gate2334(.a(gate114inter8), .b(gate114inter7), .O(gate114inter9));
  nand2 gate2335(.a(s_255), .b(gate114inter3), .O(gate114inter10));
  nor2  gate2336(.a(gate114inter10), .b(gate114inter9), .O(gate114inter11));
  nor2  gate2337(.a(gate114inter11), .b(gate114inter6), .O(gate114inter12));
  nand2 gate2338(.a(gate114inter12), .b(gate114inter1), .O(G453));

  xor2  gate1205(.a(G383), .b(G382), .O(gate115inter0));
  nand2 gate1206(.a(gate115inter0), .b(s_94), .O(gate115inter1));
  and2  gate1207(.a(G383), .b(G382), .O(gate115inter2));
  inv1  gate1208(.a(s_94), .O(gate115inter3));
  inv1  gate1209(.a(s_95), .O(gate115inter4));
  nand2 gate1210(.a(gate115inter4), .b(gate115inter3), .O(gate115inter5));
  nor2  gate1211(.a(gate115inter5), .b(gate115inter2), .O(gate115inter6));
  inv1  gate1212(.a(G382), .O(gate115inter7));
  inv1  gate1213(.a(G383), .O(gate115inter8));
  nand2 gate1214(.a(gate115inter8), .b(gate115inter7), .O(gate115inter9));
  nand2 gate1215(.a(s_95), .b(gate115inter3), .O(gate115inter10));
  nor2  gate1216(.a(gate115inter10), .b(gate115inter9), .O(gate115inter11));
  nor2  gate1217(.a(gate115inter11), .b(gate115inter6), .O(gate115inter12));
  nand2 gate1218(.a(gate115inter12), .b(gate115inter1), .O(G456));

  xor2  gate939(.a(G385), .b(G384), .O(gate116inter0));
  nand2 gate940(.a(gate116inter0), .b(s_56), .O(gate116inter1));
  and2  gate941(.a(G385), .b(G384), .O(gate116inter2));
  inv1  gate942(.a(s_56), .O(gate116inter3));
  inv1  gate943(.a(s_57), .O(gate116inter4));
  nand2 gate944(.a(gate116inter4), .b(gate116inter3), .O(gate116inter5));
  nor2  gate945(.a(gate116inter5), .b(gate116inter2), .O(gate116inter6));
  inv1  gate946(.a(G384), .O(gate116inter7));
  inv1  gate947(.a(G385), .O(gate116inter8));
  nand2 gate948(.a(gate116inter8), .b(gate116inter7), .O(gate116inter9));
  nand2 gate949(.a(s_57), .b(gate116inter3), .O(gate116inter10));
  nor2  gate950(.a(gate116inter10), .b(gate116inter9), .O(gate116inter11));
  nor2  gate951(.a(gate116inter11), .b(gate116inter6), .O(gate116inter12));
  nand2 gate952(.a(gate116inter12), .b(gate116inter1), .O(G459));

  xor2  gate1849(.a(G387), .b(G386), .O(gate117inter0));
  nand2 gate1850(.a(gate117inter0), .b(s_186), .O(gate117inter1));
  and2  gate1851(.a(G387), .b(G386), .O(gate117inter2));
  inv1  gate1852(.a(s_186), .O(gate117inter3));
  inv1  gate1853(.a(s_187), .O(gate117inter4));
  nand2 gate1854(.a(gate117inter4), .b(gate117inter3), .O(gate117inter5));
  nor2  gate1855(.a(gate117inter5), .b(gate117inter2), .O(gate117inter6));
  inv1  gate1856(.a(G386), .O(gate117inter7));
  inv1  gate1857(.a(G387), .O(gate117inter8));
  nand2 gate1858(.a(gate117inter8), .b(gate117inter7), .O(gate117inter9));
  nand2 gate1859(.a(s_187), .b(gate117inter3), .O(gate117inter10));
  nor2  gate1860(.a(gate117inter10), .b(gate117inter9), .O(gate117inter11));
  nor2  gate1861(.a(gate117inter11), .b(gate117inter6), .O(gate117inter12));
  nand2 gate1862(.a(gate117inter12), .b(gate117inter1), .O(G462));
nand2 gate118( .a(G388), .b(G389), .O(G465) );

  xor2  gate1457(.a(G391), .b(G390), .O(gate119inter0));
  nand2 gate1458(.a(gate119inter0), .b(s_130), .O(gate119inter1));
  and2  gate1459(.a(G391), .b(G390), .O(gate119inter2));
  inv1  gate1460(.a(s_130), .O(gate119inter3));
  inv1  gate1461(.a(s_131), .O(gate119inter4));
  nand2 gate1462(.a(gate119inter4), .b(gate119inter3), .O(gate119inter5));
  nor2  gate1463(.a(gate119inter5), .b(gate119inter2), .O(gate119inter6));
  inv1  gate1464(.a(G390), .O(gate119inter7));
  inv1  gate1465(.a(G391), .O(gate119inter8));
  nand2 gate1466(.a(gate119inter8), .b(gate119inter7), .O(gate119inter9));
  nand2 gate1467(.a(s_131), .b(gate119inter3), .O(gate119inter10));
  nor2  gate1468(.a(gate119inter10), .b(gate119inter9), .O(gate119inter11));
  nor2  gate1469(.a(gate119inter11), .b(gate119inter6), .O(gate119inter12));
  nand2 gate1470(.a(gate119inter12), .b(gate119inter1), .O(G468));
nand2 gate120( .a(G392), .b(G393), .O(G471) );

  xor2  gate2297(.a(G395), .b(G394), .O(gate121inter0));
  nand2 gate2298(.a(gate121inter0), .b(s_250), .O(gate121inter1));
  and2  gate2299(.a(G395), .b(G394), .O(gate121inter2));
  inv1  gate2300(.a(s_250), .O(gate121inter3));
  inv1  gate2301(.a(s_251), .O(gate121inter4));
  nand2 gate2302(.a(gate121inter4), .b(gate121inter3), .O(gate121inter5));
  nor2  gate2303(.a(gate121inter5), .b(gate121inter2), .O(gate121inter6));
  inv1  gate2304(.a(G394), .O(gate121inter7));
  inv1  gate2305(.a(G395), .O(gate121inter8));
  nand2 gate2306(.a(gate121inter8), .b(gate121inter7), .O(gate121inter9));
  nand2 gate2307(.a(s_251), .b(gate121inter3), .O(gate121inter10));
  nor2  gate2308(.a(gate121inter10), .b(gate121inter9), .O(gate121inter11));
  nor2  gate2309(.a(gate121inter11), .b(gate121inter6), .O(gate121inter12));
  nand2 gate2310(.a(gate121inter12), .b(gate121inter1), .O(G474));
nand2 gate122( .a(G396), .b(G397), .O(G477) );

  xor2  gate2759(.a(G399), .b(G398), .O(gate123inter0));
  nand2 gate2760(.a(gate123inter0), .b(s_316), .O(gate123inter1));
  and2  gate2761(.a(G399), .b(G398), .O(gate123inter2));
  inv1  gate2762(.a(s_316), .O(gate123inter3));
  inv1  gate2763(.a(s_317), .O(gate123inter4));
  nand2 gate2764(.a(gate123inter4), .b(gate123inter3), .O(gate123inter5));
  nor2  gate2765(.a(gate123inter5), .b(gate123inter2), .O(gate123inter6));
  inv1  gate2766(.a(G398), .O(gate123inter7));
  inv1  gate2767(.a(G399), .O(gate123inter8));
  nand2 gate2768(.a(gate123inter8), .b(gate123inter7), .O(gate123inter9));
  nand2 gate2769(.a(s_317), .b(gate123inter3), .O(gate123inter10));
  nor2  gate2770(.a(gate123inter10), .b(gate123inter9), .O(gate123inter11));
  nor2  gate2771(.a(gate123inter11), .b(gate123inter6), .O(gate123inter12));
  nand2 gate2772(.a(gate123inter12), .b(gate123inter1), .O(G480));

  xor2  gate1121(.a(G401), .b(G400), .O(gate124inter0));
  nand2 gate1122(.a(gate124inter0), .b(s_82), .O(gate124inter1));
  and2  gate1123(.a(G401), .b(G400), .O(gate124inter2));
  inv1  gate1124(.a(s_82), .O(gate124inter3));
  inv1  gate1125(.a(s_83), .O(gate124inter4));
  nand2 gate1126(.a(gate124inter4), .b(gate124inter3), .O(gate124inter5));
  nor2  gate1127(.a(gate124inter5), .b(gate124inter2), .O(gate124inter6));
  inv1  gate1128(.a(G400), .O(gate124inter7));
  inv1  gate1129(.a(G401), .O(gate124inter8));
  nand2 gate1130(.a(gate124inter8), .b(gate124inter7), .O(gate124inter9));
  nand2 gate1131(.a(s_83), .b(gate124inter3), .O(gate124inter10));
  nor2  gate1132(.a(gate124inter10), .b(gate124inter9), .O(gate124inter11));
  nor2  gate1133(.a(gate124inter11), .b(gate124inter6), .O(gate124inter12));
  nand2 gate1134(.a(gate124inter12), .b(gate124inter1), .O(G483));
nand2 gate125( .a(G402), .b(G403), .O(G486) );
nand2 gate126( .a(G404), .b(G405), .O(G489) );
nand2 gate127( .a(G406), .b(G407), .O(G492) );

  xor2  gate1051(.a(G409), .b(G408), .O(gate128inter0));
  nand2 gate1052(.a(gate128inter0), .b(s_72), .O(gate128inter1));
  and2  gate1053(.a(G409), .b(G408), .O(gate128inter2));
  inv1  gate1054(.a(s_72), .O(gate128inter3));
  inv1  gate1055(.a(s_73), .O(gate128inter4));
  nand2 gate1056(.a(gate128inter4), .b(gate128inter3), .O(gate128inter5));
  nor2  gate1057(.a(gate128inter5), .b(gate128inter2), .O(gate128inter6));
  inv1  gate1058(.a(G408), .O(gate128inter7));
  inv1  gate1059(.a(G409), .O(gate128inter8));
  nand2 gate1060(.a(gate128inter8), .b(gate128inter7), .O(gate128inter9));
  nand2 gate1061(.a(s_73), .b(gate128inter3), .O(gate128inter10));
  nor2  gate1062(.a(gate128inter10), .b(gate128inter9), .O(gate128inter11));
  nor2  gate1063(.a(gate128inter11), .b(gate128inter6), .O(gate128inter12));
  nand2 gate1064(.a(gate128inter12), .b(gate128inter1), .O(G495));
nand2 gate129( .a(G410), .b(G411), .O(G498) );

  xor2  gate1135(.a(G413), .b(G412), .O(gate130inter0));
  nand2 gate1136(.a(gate130inter0), .b(s_84), .O(gate130inter1));
  and2  gate1137(.a(G413), .b(G412), .O(gate130inter2));
  inv1  gate1138(.a(s_84), .O(gate130inter3));
  inv1  gate1139(.a(s_85), .O(gate130inter4));
  nand2 gate1140(.a(gate130inter4), .b(gate130inter3), .O(gate130inter5));
  nor2  gate1141(.a(gate130inter5), .b(gate130inter2), .O(gate130inter6));
  inv1  gate1142(.a(G412), .O(gate130inter7));
  inv1  gate1143(.a(G413), .O(gate130inter8));
  nand2 gate1144(.a(gate130inter8), .b(gate130inter7), .O(gate130inter9));
  nand2 gate1145(.a(s_85), .b(gate130inter3), .O(gate130inter10));
  nor2  gate1146(.a(gate130inter10), .b(gate130inter9), .O(gate130inter11));
  nor2  gate1147(.a(gate130inter11), .b(gate130inter6), .O(gate130inter12));
  nand2 gate1148(.a(gate130inter12), .b(gate130inter1), .O(G501));
nand2 gate131( .a(G414), .b(G415), .O(G504) );
nand2 gate132( .a(G416), .b(G417), .O(G507) );

  xor2  gate897(.a(G419), .b(G418), .O(gate133inter0));
  nand2 gate898(.a(gate133inter0), .b(s_50), .O(gate133inter1));
  and2  gate899(.a(G419), .b(G418), .O(gate133inter2));
  inv1  gate900(.a(s_50), .O(gate133inter3));
  inv1  gate901(.a(s_51), .O(gate133inter4));
  nand2 gate902(.a(gate133inter4), .b(gate133inter3), .O(gate133inter5));
  nor2  gate903(.a(gate133inter5), .b(gate133inter2), .O(gate133inter6));
  inv1  gate904(.a(G418), .O(gate133inter7));
  inv1  gate905(.a(G419), .O(gate133inter8));
  nand2 gate906(.a(gate133inter8), .b(gate133inter7), .O(gate133inter9));
  nand2 gate907(.a(s_51), .b(gate133inter3), .O(gate133inter10));
  nor2  gate908(.a(gate133inter10), .b(gate133inter9), .O(gate133inter11));
  nor2  gate909(.a(gate133inter11), .b(gate133inter6), .O(gate133inter12));
  nand2 gate910(.a(gate133inter12), .b(gate133inter1), .O(G510));
nand2 gate134( .a(G420), .b(G421), .O(G513) );
nand2 gate135( .a(G422), .b(G423), .O(G516) );

  xor2  gate729(.a(G425), .b(G424), .O(gate136inter0));
  nand2 gate730(.a(gate136inter0), .b(s_26), .O(gate136inter1));
  and2  gate731(.a(G425), .b(G424), .O(gate136inter2));
  inv1  gate732(.a(s_26), .O(gate136inter3));
  inv1  gate733(.a(s_27), .O(gate136inter4));
  nand2 gate734(.a(gate136inter4), .b(gate136inter3), .O(gate136inter5));
  nor2  gate735(.a(gate136inter5), .b(gate136inter2), .O(gate136inter6));
  inv1  gate736(.a(G424), .O(gate136inter7));
  inv1  gate737(.a(G425), .O(gate136inter8));
  nand2 gate738(.a(gate136inter8), .b(gate136inter7), .O(gate136inter9));
  nand2 gate739(.a(s_27), .b(gate136inter3), .O(gate136inter10));
  nor2  gate740(.a(gate136inter10), .b(gate136inter9), .O(gate136inter11));
  nor2  gate741(.a(gate136inter11), .b(gate136inter6), .O(gate136inter12));
  nand2 gate742(.a(gate136inter12), .b(gate136inter1), .O(G519));

  xor2  gate785(.a(G429), .b(G426), .O(gate137inter0));
  nand2 gate786(.a(gate137inter0), .b(s_34), .O(gate137inter1));
  and2  gate787(.a(G429), .b(G426), .O(gate137inter2));
  inv1  gate788(.a(s_34), .O(gate137inter3));
  inv1  gate789(.a(s_35), .O(gate137inter4));
  nand2 gate790(.a(gate137inter4), .b(gate137inter3), .O(gate137inter5));
  nor2  gate791(.a(gate137inter5), .b(gate137inter2), .O(gate137inter6));
  inv1  gate792(.a(G426), .O(gate137inter7));
  inv1  gate793(.a(G429), .O(gate137inter8));
  nand2 gate794(.a(gate137inter8), .b(gate137inter7), .O(gate137inter9));
  nand2 gate795(.a(s_35), .b(gate137inter3), .O(gate137inter10));
  nor2  gate796(.a(gate137inter10), .b(gate137inter9), .O(gate137inter11));
  nor2  gate797(.a(gate137inter11), .b(gate137inter6), .O(gate137inter12));
  nand2 gate798(.a(gate137inter12), .b(gate137inter1), .O(G522));
nand2 gate138( .a(G432), .b(G435), .O(G525) );

  xor2  gate2339(.a(G441), .b(G438), .O(gate139inter0));
  nand2 gate2340(.a(gate139inter0), .b(s_256), .O(gate139inter1));
  and2  gate2341(.a(G441), .b(G438), .O(gate139inter2));
  inv1  gate2342(.a(s_256), .O(gate139inter3));
  inv1  gate2343(.a(s_257), .O(gate139inter4));
  nand2 gate2344(.a(gate139inter4), .b(gate139inter3), .O(gate139inter5));
  nor2  gate2345(.a(gate139inter5), .b(gate139inter2), .O(gate139inter6));
  inv1  gate2346(.a(G438), .O(gate139inter7));
  inv1  gate2347(.a(G441), .O(gate139inter8));
  nand2 gate2348(.a(gate139inter8), .b(gate139inter7), .O(gate139inter9));
  nand2 gate2349(.a(s_257), .b(gate139inter3), .O(gate139inter10));
  nor2  gate2350(.a(gate139inter10), .b(gate139inter9), .O(gate139inter11));
  nor2  gate2351(.a(gate139inter11), .b(gate139inter6), .O(gate139inter12));
  nand2 gate2352(.a(gate139inter12), .b(gate139inter1), .O(G528));
nand2 gate140( .a(G444), .b(G447), .O(G531) );
nand2 gate141( .a(G450), .b(G453), .O(G534) );
nand2 gate142( .a(G456), .b(G459), .O(G537) );
nand2 gate143( .a(G462), .b(G465), .O(G540) );
nand2 gate144( .a(G468), .b(G471), .O(G543) );
nand2 gate145( .a(G474), .b(G477), .O(G546) );
nand2 gate146( .a(G480), .b(G483), .O(G549) );
nand2 gate147( .a(G486), .b(G489), .O(G552) );
nand2 gate148( .a(G492), .b(G495), .O(G555) );
nand2 gate149( .a(G498), .b(G501), .O(G558) );
nand2 gate150( .a(G504), .b(G507), .O(G561) );

  xor2  gate869(.a(G513), .b(G510), .O(gate151inter0));
  nand2 gate870(.a(gate151inter0), .b(s_46), .O(gate151inter1));
  and2  gate871(.a(G513), .b(G510), .O(gate151inter2));
  inv1  gate872(.a(s_46), .O(gate151inter3));
  inv1  gate873(.a(s_47), .O(gate151inter4));
  nand2 gate874(.a(gate151inter4), .b(gate151inter3), .O(gate151inter5));
  nor2  gate875(.a(gate151inter5), .b(gate151inter2), .O(gate151inter6));
  inv1  gate876(.a(G510), .O(gate151inter7));
  inv1  gate877(.a(G513), .O(gate151inter8));
  nand2 gate878(.a(gate151inter8), .b(gate151inter7), .O(gate151inter9));
  nand2 gate879(.a(s_47), .b(gate151inter3), .O(gate151inter10));
  nor2  gate880(.a(gate151inter10), .b(gate151inter9), .O(gate151inter11));
  nor2  gate881(.a(gate151inter11), .b(gate151inter6), .O(gate151inter12));
  nand2 gate882(.a(gate151inter12), .b(gate151inter1), .O(G564));
nand2 gate152( .a(G516), .b(G519), .O(G567) );
nand2 gate153( .a(G426), .b(G522), .O(G570) );

  xor2  gate2213(.a(G522), .b(G429), .O(gate154inter0));
  nand2 gate2214(.a(gate154inter0), .b(s_238), .O(gate154inter1));
  and2  gate2215(.a(G522), .b(G429), .O(gate154inter2));
  inv1  gate2216(.a(s_238), .O(gate154inter3));
  inv1  gate2217(.a(s_239), .O(gate154inter4));
  nand2 gate2218(.a(gate154inter4), .b(gate154inter3), .O(gate154inter5));
  nor2  gate2219(.a(gate154inter5), .b(gate154inter2), .O(gate154inter6));
  inv1  gate2220(.a(G429), .O(gate154inter7));
  inv1  gate2221(.a(G522), .O(gate154inter8));
  nand2 gate2222(.a(gate154inter8), .b(gate154inter7), .O(gate154inter9));
  nand2 gate2223(.a(s_239), .b(gate154inter3), .O(gate154inter10));
  nor2  gate2224(.a(gate154inter10), .b(gate154inter9), .O(gate154inter11));
  nor2  gate2225(.a(gate154inter11), .b(gate154inter6), .O(gate154inter12));
  nand2 gate2226(.a(gate154inter12), .b(gate154inter1), .O(G571));

  xor2  gate827(.a(G525), .b(G432), .O(gate155inter0));
  nand2 gate828(.a(gate155inter0), .b(s_40), .O(gate155inter1));
  and2  gate829(.a(G525), .b(G432), .O(gate155inter2));
  inv1  gate830(.a(s_40), .O(gate155inter3));
  inv1  gate831(.a(s_41), .O(gate155inter4));
  nand2 gate832(.a(gate155inter4), .b(gate155inter3), .O(gate155inter5));
  nor2  gate833(.a(gate155inter5), .b(gate155inter2), .O(gate155inter6));
  inv1  gate834(.a(G432), .O(gate155inter7));
  inv1  gate835(.a(G525), .O(gate155inter8));
  nand2 gate836(.a(gate155inter8), .b(gate155inter7), .O(gate155inter9));
  nand2 gate837(.a(s_41), .b(gate155inter3), .O(gate155inter10));
  nor2  gate838(.a(gate155inter10), .b(gate155inter9), .O(gate155inter11));
  nor2  gate839(.a(gate155inter11), .b(gate155inter6), .O(gate155inter12));
  nand2 gate840(.a(gate155inter12), .b(gate155inter1), .O(G572));
nand2 gate156( .a(G435), .b(G525), .O(G573) );
nand2 gate157( .a(G438), .b(G528), .O(G574) );

  xor2  gate1275(.a(G528), .b(G441), .O(gate158inter0));
  nand2 gate1276(.a(gate158inter0), .b(s_104), .O(gate158inter1));
  and2  gate1277(.a(G528), .b(G441), .O(gate158inter2));
  inv1  gate1278(.a(s_104), .O(gate158inter3));
  inv1  gate1279(.a(s_105), .O(gate158inter4));
  nand2 gate1280(.a(gate158inter4), .b(gate158inter3), .O(gate158inter5));
  nor2  gate1281(.a(gate158inter5), .b(gate158inter2), .O(gate158inter6));
  inv1  gate1282(.a(G441), .O(gate158inter7));
  inv1  gate1283(.a(G528), .O(gate158inter8));
  nand2 gate1284(.a(gate158inter8), .b(gate158inter7), .O(gate158inter9));
  nand2 gate1285(.a(s_105), .b(gate158inter3), .O(gate158inter10));
  nor2  gate1286(.a(gate158inter10), .b(gate158inter9), .O(gate158inter11));
  nor2  gate1287(.a(gate158inter11), .b(gate158inter6), .O(gate158inter12));
  nand2 gate1288(.a(gate158inter12), .b(gate158inter1), .O(G575));
nand2 gate159( .a(G444), .b(G531), .O(G576) );

  xor2  gate2619(.a(G531), .b(G447), .O(gate160inter0));
  nand2 gate2620(.a(gate160inter0), .b(s_296), .O(gate160inter1));
  and2  gate2621(.a(G531), .b(G447), .O(gate160inter2));
  inv1  gate2622(.a(s_296), .O(gate160inter3));
  inv1  gate2623(.a(s_297), .O(gate160inter4));
  nand2 gate2624(.a(gate160inter4), .b(gate160inter3), .O(gate160inter5));
  nor2  gate2625(.a(gate160inter5), .b(gate160inter2), .O(gate160inter6));
  inv1  gate2626(.a(G447), .O(gate160inter7));
  inv1  gate2627(.a(G531), .O(gate160inter8));
  nand2 gate2628(.a(gate160inter8), .b(gate160inter7), .O(gate160inter9));
  nand2 gate2629(.a(s_297), .b(gate160inter3), .O(gate160inter10));
  nor2  gate2630(.a(gate160inter10), .b(gate160inter9), .O(gate160inter11));
  nor2  gate2631(.a(gate160inter11), .b(gate160inter6), .O(gate160inter12));
  nand2 gate2632(.a(gate160inter12), .b(gate160inter1), .O(G577));
nand2 gate161( .a(G450), .b(G534), .O(G578) );
nand2 gate162( .a(G453), .b(G534), .O(G579) );
nand2 gate163( .a(G456), .b(G537), .O(G580) );
nand2 gate164( .a(G459), .b(G537), .O(G581) );

  xor2  gate1317(.a(G540), .b(G462), .O(gate165inter0));
  nand2 gate1318(.a(gate165inter0), .b(s_110), .O(gate165inter1));
  and2  gate1319(.a(G540), .b(G462), .O(gate165inter2));
  inv1  gate1320(.a(s_110), .O(gate165inter3));
  inv1  gate1321(.a(s_111), .O(gate165inter4));
  nand2 gate1322(.a(gate165inter4), .b(gate165inter3), .O(gate165inter5));
  nor2  gate1323(.a(gate165inter5), .b(gate165inter2), .O(gate165inter6));
  inv1  gate1324(.a(G462), .O(gate165inter7));
  inv1  gate1325(.a(G540), .O(gate165inter8));
  nand2 gate1326(.a(gate165inter8), .b(gate165inter7), .O(gate165inter9));
  nand2 gate1327(.a(s_111), .b(gate165inter3), .O(gate165inter10));
  nor2  gate1328(.a(gate165inter10), .b(gate165inter9), .O(gate165inter11));
  nor2  gate1329(.a(gate165inter11), .b(gate165inter6), .O(gate165inter12));
  nand2 gate1330(.a(gate165inter12), .b(gate165inter1), .O(G582));
nand2 gate166( .a(G465), .b(G540), .O(G583) );

  xor2  gate1527(.a(G543), .b(G468), .O(gate167inter0));
  nand2 gate1528(.a(gate167inter0), .b(s_140), .O(gate167inter1));
  and2  gate1529(.a(G543), .b(G468), .O(gate167inter2));
  inv1  gate1530(.a(s_140), .O(gate167inter3));
  inv1  gate1531(.a(s_141), .O(gate167inter4));
  nand2 gate1532(.a(gate167inter4), .b(gate167inter3), .O(gate167inter5));
  nor2  gate1533(.a(gate167inter5), .b(gate167inter2), .O(gate167inter6));
  inv1  gate1534(.a(G468), .O(gate167inter7));
  inv1  gate1535(.a(G543), .O(gate167inter8));
  nand2 gate1536(.a(gate167inter8), .b(gate167inter7), .O(gate167inter9));
  nand2 gate1537(.a(s_141), .b(gate167inter3), .O(gate167inter10));
  nor2  gate1538(.a(gate167inter10), .b(gate167inter9), .O(gate167inter11));
  nor2  gate1539(.a(gate167inter11), .b(gate167inter6), .O(gate167inter12));
  nand2 gate1540(.a(gate167inter12), .b(gate167inter1), .O(G584));
nand2 gate168( .a(G471), .b(G543), .O(G585) );

  xor2  gate883(.a(G546), .b(G474), .O(gate169inter0));
  nand2 gate884(.a(gate169inter0), .b(s_48), .O(gate169inter1));
  and2  gate885(.a(G546), .b(G474), .O(gate169inter2));
  inv1  gate886(.a(s_48), .O(gate169inter3));
  inv1  gate887(.a(s_49), .O(gate169inter4));
  nand2 gate888(.a(gate169inter4), .b(gate169inter3), .O(gate169inter5));
  nor2  gate889(.a(gate169inter5), .b(gate169inter2), .O(gate169inter6));
  inv1  gate890(.a(G474), .O(gate169inter7));
  inv1  gate891(.a(G546), .O(gate169inter8));
  nand2 gate892(.a(gate169inter8), .b(gate169inter7), .O(gate169inter9));
  nand2 gate893(.a(s_49), .b(gate169inter3), .O(gate169inter10));
  nor2  gate894(.a(gate169inter10), .b(gate169inter9), .O(gate169inter11));
  nor2  gate895(.a(gate169inter11), .b(gate169inter6), .O(gate169inter12));
  nand2 gate896(.a(gate169inter12), .b(gate169inter1), .O(G586));

  xor2  gate1737(.a(G546), .b(G477), .O(gate170inter0));
  nand2 gate1738(.a(gate170inter0), .b(s_170), .O(gate170inter1));
  and2  gate1739(.a(G546), .b(G477), .O(gate170inter2));
  inv1  gate1740(.a(s_170), .O(gate170inter3));
  inv1  gate1741(.a(s_171), .O(gate170inter4));
  nand2 gate1742(.a(gate170inter4), .b(gate170inter3), .O(gate170inter5));
  nor2  gate1743(.a(gate170inter5), .b(gate170inter2), .O(gate170inter6));
  inv1  gate1744(.a(G477), .O(gate170inter7));
  inv1  gate1745(.a(G546), .O(gate170inter8));
  nand2 gate1746(.a(gate170inter8), .b(gate170inter7), .O(gate170inter9));
  nand2 gate1747(.a(s_171), .b(gate170inter3), .O(gate170inter10));
  nor2  gate1748(.a(gate170inter10), .b(gate170inter9), .O(gate170inter11));
  nor2  gate1749(.a(gate170inter11), .b(gate170inter6), .O(gate170inter12));
  nand2 gate1750(.a(gate170inter12), .b(gate170inter1), .O(G587));

  xor2  gate841(.a(G549), .b(G480), .O(gate171inter0));
  nand2 gate842(.a(gate171inter0), .b(s_42), .O(gate171inter1));
  and2  gate843(.a(G549), .b(G480), .O(gate171inter2));
  inv1  gate844(.a(s_42), .O(gate171inter3));
  inv1  gate845(.a(s_43), .O(gate171inter4));
  nand2 gate846(.a(gate171inter4), .b(gate171inter3), .O(gate171inter5));
  nor2  gate847(.a(gate171inter5), .b(gate171inter2), .O(gate171inter6));
  inv1  gate848(.a(G480), .O(gate171inter7));
  inv1  gate849(.a(G549), .O(gate171inter8));
  nand2 gate850(.a(gate171inter8), .b(gate171inter7), .O(gate171inter9));
  nand2 gate851(.a(s_43), .b(gate171inter3), .O(gate171inter10));
  nor2  gate852(.a(gate171inter10), .b(gate171inter9), .O(gate171inter11));
  nor2  gate853(.a(gate171inter11), .b(gate171inter6), .O(gate171inter12));
  nand2 gate854(.a(gate171inter12), .b(gate171inter1), .O(G588));

  xor2  gate1303(.a(G549), .b(G483), .O(gate172inter0));
  nand2 gate1304(.a(gate172inter0), .b(s_108), .O(gate172inter1));
  and2  gate1305(.a(G549), .b(G483), .O(gate172inter2));
  inv1  gate1306(.a(s_108), .O(gate172inter3));
  inv1  gate1307(.a(s_109), .O(gate172inter4));
  nand2 gate1308(.a(gate172inter4), .b(gate172inter3), .O(gate172inter5));
  nor2  gate1309(.a(gate172inter5), .b(gate172inter2), .O(gate172inter6));
  inv1  gate1310(.a(G483), .O(gate172inter7));
  inv1  gate1311(.a(G549), .O(gate172inter8));
  nand2 gate1312(.a(gate172inter8), .b(gate172inter7), .O(gate172inter9));
  nand2 gate1313(.a(s_109), .b(gate172inter3), .O(gate172inter10));
  nor2  gate1314(.a(gate172inter10), .b(gate172inter9), .O(gate172inter11));
  nor2  gate1315(.a(gate172inter11), .b(gate172inter6), .O(gate172inter12));
  nand2 gate1316(.a(gate172inter12), .b(gate172inter1), .O(G589));

  xor2  gate1667(.a(G552), .b(G486), .O(gate173inter0));
  nand2 gate1668(.a(gate173inter0), .b(s_160), .O(gate173inter1));
  and2  gate1669(.a(G552), .b(G486), .O(gate173inter2));
  inv1  gate1670(.a(s_160), .O(gate173inter3));
  inv1  gate1671(.a(s_161), .O(gate173inter4));
  nand2 gate1672(.a(gate173inter4), .b(gate173inter3), .O(gate173inter5));
  nor2  gate1673(.a(gate173inter5), .b(gate173inter2), .O(gate173inter6));
  inv1  gate1674(.a(G486), .O(gate173inter7));
  inv1  gate1675(.a(G552), .O(gate173inter8));
  nand2 gate1676(.a(gate173inter8), .b(gate173inter7), .O(gate173inter9));
  nand2 gate1677(.a(s_161), .b(gate173inter3), .O(gate173inter10));
  nor2  gate1678(.a(gate173inter10), .b(gate173inter9), .O(gate173inter11));
  nor2  gate1679(.a(gate173inter11), .b(gate173inter6), .O(gate173inter12));
  nand2 gate1680(.a(gate173inter12), .b(gate173inter1), .O(G590));

  xor2  gate1709(.a(G552), .b(G489), .O(gate174inter0));
  nand2 gate1710(.a(gate174inter0), .b(s_166), .O(gate174inter1));
  and2  gate1711(.a(G552), .b(G489), .O(gate174inter2));
  inv1  gate1712(.a(s_166), .O(gate174inter3));
  inv1  gate1713(.a(s_167), .O(gate174inter4));
  nand2 gate1714(.a(gate174inter4), .b(gate174inter3), .O(gate174inter5));
  nor2  gate1715(.a(gate174inter5), .b(gate174inter2), .O(gate174inter6));
  inv1  gate1716(.a(G489), .O(gate174inter7));
  inv1  gate1717(.a(G552), .O(gate174inter8));
  nand2 gate1718(.a(gate174inter8), .b(gate174inter7), .O(gate174inter9));
  nand2 gate1719(.a(s_167), .b(gate174inter3), .O(gate174inter10));
  nor2  gate1720(.a(gate174inter10), .b(gate174inter9), .O(gate174inter11));
  nor2  gate1721(.a(gate174inter11), .b(gate174inter6), .O(gate174inter12));
  nand2 gate1722(.a(gate174inter12), .b(gate174inter1), .O(G591));
nand2 gate175( .a(G492), .b(G555), .O(G592) );
nand2 gate176( .a(G495), .b(G555), .O(G593) );
nand2 gate177( .a(G498), .b(G558), .O(G594) );

  xor2  gate2549(.a(G558), .b(G501), .O(gate178inter0));
  nand2 gate2550(.a(gate178inter0), .b(s_286), .O(gate178inter1));
  and2  gate2551(.a(G558), .b(G501), .O(gate178inter2));
  inv1  gate2552(.a(s_286), .O(gate178inter3));
  inv1  gate2553(.a(s_287), .O(gate178inter4));
  nand2 gate2554(.a(gate178inter4), .b(gate178inter3), .O(gate178inter5));
  nor2  gate2555(.a(gate178inter5), .b(gate178inter2), .O(gate178inter6));
  inv1  gate2556(.a(G501), .O(gate178inter7));
  inv1  gate2557(.a(G558), .O(gate178inter8));
  nand2 gate2558(.a(gate178inter8), .b(gate178inter7), .O(gate178inter9));
  nand2 gate2559(.a(s_287), .b(gate178inter3), .O(gate178inter10));
  nor2  gate2560(.a(gate178inter10), .b(gate178inter9), .O(gate178inter11));
  nor2  gate2561(.a(gate178inter11), .b(gate178inter6), .O(gate178inter12));
  nand2 gate2562(.a(gate178inter12), .b(gate178inter1), .O(G595));
nand2 gate179( .a(G504), .b(G561), .O(G596) );

  xor2  gate2591(.a(G561), .b(G507), .O(gate180inter0));
  nand2 gate2592(.a(gate180inter0), .b(s_292), .O(gate180inter1));
  and2  gate2593(.a(G561), .b(G507), .O(gate180inter2));
  inv1  gate2594(.a(s_292), .O(gate180inter3));
  inv1  gate2595(.a(s_293), .O(gate180inter4));
  nand2 gate2596(.a(gate180inter4), .b(gate180inter3), .O(gate180inter5));
  nor2  gate2597(.a(gate180inter5), .b(gate180inter2), .O(gate180inter6));
  inv1  gate2598(.a(G507), .O(gate180inter7));
  inv1  gate2599(.a(G561), .O(gate180inter8));
  nand2 gate2600(.a(gate180inter8), .b(gate180inter7), .O(gate180inter9));
  nand2 gate2601(.a(s_293), .b(gate180inter3), .O(gate180inter10));
  nor2  gate2602(.a(gate180inter10), .b(gate180inter9), .O(gate180inter11));
  nor2  gate2603(.a(gate180inter11), .b(gate180inter6), .O(gate180inter12));
  nand2 gate2604(.a(gate180inter12), .b(gate180inter1), .O(G597));

  xor2  gate1919(.a(G564), .b(G510), .O(gate181inter0));
  nand2 gate1920(.a(gate181inter0), .b(s_196), .O(gate181inter1));
  and2  gate1921(.a(G564), .b(G510), .O(gate181inter2));
  inv1  gate1922(.a(s_196), .O(gate181inter3));
  inv1  gate1923(.a(s_197), .O(gate181inter4));
  nand2 gate1924(.a(gate181inter4), .b(gate181inter3), .O(gate181inter5));
  nor2  gate1925(.a(gate181inter5), .b(gate181inter2), .O(gate181inter6));
  inv1  gate1926(.a(G510), .O(gate181inter7));
  inv1  gate1927(.a(G564), .O(gate181inter8));
  nand2 gate1928(.a(gate181inter8), .b(gate181inter7), .O(gate181inter9));
  nand2 gate1929(.a(s_197), .b(gate181inter3), .O(gate181inter10));
  nor2  gate1930(.a(gate181inter10), .b(gate181inter9), .O(gate181inter11));
  nor2  gate1931(.a(gate181inter11), .b(gate181inter6), .O(gate181inter12));
  nand2 gate1932(.a(gate181inter12), .b(gate181inter1), .O(G598));

  xor2  gate2745(.a(G564), .b(G513), .O(gate182inter0));
  nand2 gate2746(.a(gate182inter0), .b(s_314), .O(gate182inter1));
  and2  gate2747(.a(G564), .b(G513), .O(gate182inter2));
  inv1  gate2748(.a(s_314), .O(gate182inter3));
  inv1  gate2749(.a(s_315), .O(gate182inter4));
  nand2 gate2750(.a(gate182inter4), .b(gate182inter3), .O(gate182inter5));
  nor2  gate2751(.a(gate182inter5), .b(gate182inter2), .O(gate182inter6));
  inv1  gate2752(.a(G513), .O(gate182inter7));
  inv1  gate2753(.a(G564), .O(gate182inter8));
  nand2 gate2754(.a(gate182inter8), .b(gate182inter7), .O(gate182inter9));
  nand2 gate2755(.a(s_315), .b(gate182inter3), .O(gate182inter10));
  nor2  gate2756(.a(gate182inter10), .b(gate182inter9), .O(gate182inter11));
  nor2  gate2757(.a(gate182inter11), .b(gate182inter6), .O(gate182inter12));
  nand2 gate2758(.a(gate182inter12), .b(gate182inter1), .O(G599));

  xor2  gate1093(.a(G567), .b(G516), .O(gate183inter0));
  nand2 gate1094(.a(gate183inter0), .b(s_78), .O(gate183inter1));
  and2  gate1095(.a(G567), .b(G516), .O(gate183inter2));
  inv1  gate1096(.a(s_78), .O(gate183inter3));
  inv1  gate1097(.a(s_79), .O(gate183inter4));
  nand2 gate1098(.a(gate183inter4), .b(gate183inter3), .O(gate183inter5));
  nor2  gate1099(.a(gate183inter5), .b(gate183inter2), .O(gate183inter6));
  inv1  gate1100(.a(G516), .O(gate183inter7));
  inv1  gate1101(.a(G567), .O(gate183inter8));
  nand2 gate1102(.a(gate183inter8), .b(gate183inter7), .O(gate183inter9));
  nand2 gate1103(.a(s_79), .b(gate183inter3), .O(gate183inter10));
  nor2  gate1104(.a(gate183inter10), .b(gate183inter9), .O(gate183inter11));
  nor2  gate1105(.a(gate183inter11), .b(gate183inter6), .O(gate183inter12));
  nand2 gate1106(.a(gate183inter12), .b(gate183inter1), .O(G600));

  xor2  gate1373(.a(G567), .b(G519), .O(gate184inter0));
  nand2 gate1374(.a(gate184inter0), .b(s_118), .O(gate184inter1));
  and2  gate1375(.a(G567), .b(G519), .O(gate184inter2));
  inv1  gate1376(.a(s_118), .O(gate184inter3));
  inv1  gate1377(.a(s_119), .O(gate184inter4));
  nand2 gate1378(.a(gate184inter4), .b(gate184inter3), .O(gate184inter5));
  nor2  gate1379(.a(gate184inter5), .b(gate184inter2), .O(gate184inter6));
  inv1  gate1380(.a(G519), .O(gate184inter7));
  inv1  gate1381(.a(G567), .O(gate184inter8));
  nand2 gate1382(.a(gate184inter8), .b(gate184inter7), .O(gate184inter9));
  nand2 gate1383(.a(s_119), .b(gate184inter3), .O(gate184inter10));
  nor2  gate1384(.a(gate184inter10), .b(gate184inter9), .O(gate184inter11));
  nor2  gate1385(.a(gate184inter11), .b(gate184inter6), .O(gate184inter12));
  nand2 gate1386(.a(gate184inter12), .b(gate184inter1), .O(G601));

  xor2  gate1415(.a(G571), .b(G570), .O(gate185inter0));
  nand2 gate1416(.a(gate185inter0), .b(s_124), .O(gate185inter1));
  and2  gate1417(.a(G571), .b(G570), .O(gate185inter2));
  inv1  gate1418(.a(s_124), .O(gate185inter3));
  inv1  gate1419(.a(s_125), .O(gate185inter4));
  nand2 gate1420(.a(gate185inter4), .b(gate185inter3), .O(gate185inter5));
  nor2  gate1421(.a(gate185inter5), .b(gate185inter2), .O(gate185inter6));
  inv1  gate1422(.a(G570), .O(gate185inter7));
  inv1  gate1423(.a(G571), .O(gate185inter8));
  nand2 gate1424(.a(gate185inter8), .b(gate185inter7), .O(gate185inter9));
  nand2 gate1425(.a(s_125), .b(gate185inter3), .O(gate185inter10));
  nor2  gate1426(.a(gate185inter10), .b(gate185inter9), .O(gate185inter11));
  nor2  gate1427(.a(gate185inter11), .b(gate185inter6), .O(gate185inter12));
  nand2 gate1428(.a(gate185inter12), .b(gate185inter1), .O(G602));
nand2 gate186( .a(G572), .b(G573), .O(G607) );

  xor2  gate2227(.a(G575), .b(G574), .O(gate187inter0));
  nand2 gate2228(.a(gate187inter0), .b(s_240), .O(gate187inter1));
  and2  gate2229(.a(G575), .b(G574), .O(gate187inter2));
  inv1  gate2230(.a(s_240), .O(gate187inter3));
  inv1  gate2231(.a(s_241), .O(gate187inter4));
  nand2 gate2232(.a(gate187inter4), .b(gate187inter3), .O(gate187inter5));
  nor2  gate2233(.a(gate187inter5), .b(gate187inter2), .O(gate187inter6));
  inv1  gate2234(.a(G574), .O(gate187inter7));
  inv1  gate2235(.a(G575), .O(gate187inter8));
  nand2 gate2236(.a(gate187inter8), .b(gate187inter7), .O(gate187inter9));
  nand2 gate2237(.a(s_241), .b(gate187inter3), .O(gate187inter10));
  nor2  gate2238(.a(gate187inter10), .b(gate187inter9), .O(gate187inter11));
  nor2  gate2239(.a(gate187inter11), .b(gate187inter6), .O(gate187inter12));
  nand2 gate2240(.a(gate187inter12), .b(gate187inter1), .O(G612));

  xor2  gate1471(.a(G577), .b(G576), .O(gate188inter0));
  nand2 gate1472(.a(gate188inter0), .b(s_132), .O(gate188inter1));
  and2  gate1473(.a(G577), .b(G576), .O(gate188inter2));
  inv1  gate1474(.a(s_132), .O(gate188inter3));
  inv1  gate1475(.a(s_133), .O(gate188inter4));
  nand2 gate1476(.a(gate188inter4), .b(gate188inter3), .O(gate188inter5));
  nor2  gate1477(.a(gate188inter5), .b(gate188inter2), .O(gate188inter6));
  inv1  gate1478(.a(G576), .O(gate188inter7));
  inv1  gate1479(.a(G577), .O(gate188inter8));
  nand2 gate1480(.a(gate188inter8), .b(gate188inter7), .O(gate188inter9));
  nand2 gate1481(.a(s_133), .b(gate188inter3), .O(gate188inter10));
  nor2  gate1482(.a(gate188inter10), .b(gate188inter9), .O(gate188inter11));
  nor2  gate1483(.a(gate188inter11), .b(gate188inter6), .O(gate188inter12));
  nand2 gate1484(.a(gate188inter12), .b(gate188inter1), .O(G617));
nand2 gate189( .a(G578), .b(G579), .O(G622) );
nand2 gate190( .a(G580), .b(G581), .O(G627) );

  xor2  gate1261(.a(G583), .b(G582), .O(gate191inter0));
  nand2 gate1262(.a(gate191inter0), .b(s_102), .O(gate191inter1));
  and2  gate1263(.a(G583), .b(G582), .O(gate191inter2));
  inv1  gate1264(.a(s_102), .O(gate191inter3));
  inv1  gate1265(.a(s_103), .O(gate191inter4));
  nand2 gate1266(.a(gate191inter4), .b(gate191inter3), .O(gate191inter5));
  nor2  gate1267(.a(gate191inter5), .b(gate191inter2), .O(gate191inter6));
  inv1  gate1268(.a(G582), .O(gate191inter7));
  inv1  gate1269(.a(G583), .O(gate191inter8));
  nand2 gate1270(.a(gate191inter8), .b(gate191inter7), .O(gate191inter9));
  nand2 gate1271(.a(s_103), .b(gate191inter3), .O(gate191inter10));
  nor2  gate1272(.a(gate191inter10), .b(gate191inter9), .O(gate191inter11));
  nor2  gate1273(.a(gate191inter11), .b(gate191inter6), .O(gate191inter12));
  nand2 gate1274(.a(gate191inter12), .b(gate191inter1), .O(G632));

  xor2  gate1695(.a(G585), .b(G584), .O(gate192inter0));
  nand2 gate1696(.a(gate192inter0), .b(s_164), .O(gate192inter1));
  and2  gate1697(.a(G585), .b(G584), .O(gate192inter2));
  inv1  gate1698(.a(s_164), .O(gate192inter3));
  inv1  gate1699(.a(s_165), .O(gate192inter4));
  nand2 gate1700(.a(gate192inter4), .b(gate192inter3), .O(gate192inter5));
  nor2  gate1701(.a(gate192inter5), .b(gate192inter2), .O(gate192inter6));
  inv1  gate1702(.a(G584), .O(gate192inter7));
  inv1  gate1703(.a(G585), .O(gate192inter8));
  nand2 gate1704(.a(gate192inter8), .b(gate192inter7), .O(gate192inter9));
  nand2 gate1705(.a(s_165), .b(gate192inter3), .O(gate192inter10));
  nor2  gate1706(.a(gate192inter10), .b(gate192inter9), .O(gate192inter11));
  nor2  gate1707(.a(gate192inter11), .b(gate192inter6), .O(gate192inter12));
  nand2 gate1708(.a(gate192inter12), .b(gate192inter1), .O(G637));
nand2 gate193( .a(G586), .b(G587), .O(G642) );

  xor2  gate2395(.a(G589), .b(G588), .O(gate194inter0));
  nand2 gate2396(.a(gate194inter0), .b(s_264), .O(gate194inter1));
  and2  gate2397(.a(G589), .b(G588), .O(gate194inter2));
  inv1  gate2398(.a(s_264), .O(gate194inter3));
  inv1  gate2399(.a(s_265), .O(gate194inter4));
  nand2 gate2400(.a(gate194inter4), .b(gate194inter3), .O(gate194inter5));
  nor2  gate2401(.a(gate194inter5), .b(gate194inter2), .O(gate194inter6));
  inv1  gate2402(.a(G588), .O(gate194inter7));
  inv1  gate2403(.a(G589), .O(gate194inter8));
  nand2 gate2404(.a(gate194inter8), .b(gate194inter7), .O(gate194inter9));
  nand2 gate2405(.a(s_265), .b(gate194inter3), .O(gate194inter10));
  nor2  gate2406(.a(gate194inter10), .b(gate194inter9), .O(gate194inter11));
  nor2  gate2407(.a(gate194inter11), .b(gate194inter6), .O(gate194inter12));
  nand2 gate2408(.a(gate194inter12), .b(gate194inter1), .O(G645));
nand2 gate195( .a(G590), .b(G591), .O(G648) );
nand2 gate196( .a(G592), .b(G593), .O(G651) );
nand2 gate197( .a(G594), .b(G595), .O(G654) );
nand2 gate198( .a(G596), .b(G597), .O(G657) );
nand2 gate199( .a(G598), .b(G599), .O(G660) );

  xor2  gate1555(.a(G601), .b(G600), .O(gate200inter0));
  nand2 gate1556(.a(gate200inter0), .b(s_144), .O(gate200inter1));
  and2  gate1557(.a(G601), .b(G600), .O(gate200inter2));
  inv1  gate1558(.a(s_144), .O(gate200inter3));
  inv1  gate1559(.a(s_145), .O(gate200inter4));
  nand2 gate1560(.a(gate200inter4), .b(gate200inter3), .O(gate200inter5));
  nor2  gate1561(.a(gate200inter5), .b(gate200inter2), .O(gate200inter6));
  inv1  gate1562(.a(G600), .O(gate200inter7));
  inv1  gate1563(.a(G601), .O(gate200inter8));
  nand2 gate1564(.a(gate200inter8), .b(gate200inter7), .O(gate200inter9));
  nand2 gate1565(.a(s_145), .b(gate200inter3), .O(gate200inter10));
  nor2  gate1566(.a(gate200inter10), .b(gate200inter9), .O(gate200inter11));
  nor2  gate1567(.a(gate200inter11), .b(gate200inter6), .O(gate200inter12));
  nand2 gate1568(.a(gate200inter12), .b(gate200inter1), .O(G663));
nand2 gate201( .a(G602), .b(G607), .O(G666) );

  xor2  gate2353(.a(G617), .b(G612), .O(gate202inter0));
  nand2 gate2354(.a(gate202inter0), .b(s_258), .O(gate202inter1));
  and2  gate2355(.a(G617), .b(G612), .O(gate202inter2));
  inv1  gate2356(.a(s_258), .O(gate202inter3));
  inv1  gate2357(.a(s_259), .O(gate202inter4));
  nand2 gate2358(.a(gate202inter4), .b(gate202inter3), .O(gate202inter5));
  nor2  gate2359(.a(gate202inter5), .b(gate202inter2), .O(gate202inter6));
  inv1  gate2360(.a(G612), .O(gate202inter7));
  inv1  gate2361(.a(G617), .O(gate202inter8));
  nand2 gate2362(.a(gate202inter8), .b(gate202inter7), .O(gate202inter9));
  nand2 gate2363(.a(s_259), .b(gate202inter3), .O(gate202inter10));
  nor2  gate2364(.a(gate202inter10), .b(gate202inter9), .O(gate202inter11));
  nor2  gate2365(.a(gate202inter11), .b(gate202inter6), .O(gate202inter12));
  nand2 gate2366(.a(gate202inter12), .b(gate202inter1), .O(G669));
nand2 gate203( .a(G602), .b(G612), .O(G672) );

  xor2  gate1975(.a(G617), .b(G607), .O(gate204inter0));
  nand2 gate1976(.a(gate204inter0), .b(s_204), .O(gate204inter1));
  and2  gate1977(.a(G617), .b(G607), .O(gate204inter2));
  inv1  gate1978(.a(s_204), .O(gate204inter3));
  inv1  gate1979(.a(s_205), .O(gate204inter4));
  nand2 gate1980(.a(gate204inter4), .b(gate204inter3), .O(gate204inter5));
  nor2  gate1981(.a(gate204inter5), .b(gate204inter2), .O(gate204inter6));
  inv1  gate1982(.a(G607), .O(gate204inter7));
  inv1  gate1983(.a(G617), .O(gate204inter8));
  nand2 gate1984(.a(gate204inter8), .b(gate204inter7), .O(gate204inter9));
  nand2 gate1985(.a(s_205), .b(gate204inter3), .O(gate204inter10));
  nor2  gate1986(.a(gate204inter10), .b(gate204inter9), .O(gate204inter11));
  nor2  gate1987(.a(gate204inter11), .b(gate204inter6), .O(gate204inter12));
  nand2 gate1988(.a(gate204inter12), .b(gate204inter1), .O(G675));
nand2 gate205( .a(G622), .b(G627), .O(G678) );
nand2 gate206( .a(G632), .b(G637), .O(G681) );
nand2 gate207( .a(G622), .b(G632), .O(G684) );

  xor2  gate1163(.a(G637), .b(G627), .O(gate208inter0));
  nand2 gate1164(.a(gate208inter0), .b(s_88), .O(gate208inter1));
  and2  gate1165(.a(G637), .b(G627), .O(gate208inter2));
  inv1  gate1166(.a(s_88), .O(gate208inter3));
  inv1  gate1167(.a(s_89), .O(gate208inter4));
  nand2 gate1168(.a(gate208inter4), .b(gate208inter3), .O(gate208inter5));
  nor2  gate1169(.a(gate208inter5), .b(gate208inter2), .O(gate208inter6));
  inv1  gate1170(.a(G627), .O(gate208inter7));
  inv1  gate1171(.a(G637), .O(gate208inter8));
  nand2 gate1172(.a(gate208inter8), .b(gate208inter7), .O(gate208inter9));
  nand2 gate1173(.a(s_89), .b(gate208inter3), .O(gate208inter10));
  nor2  gate1174(.a(gate208inter10), .b(gate208inter9), .O(gate208inter11));
  nor2  gate1175(.a(gate208inter11), .b(gate208inter6), .O(gate208inter12));
  nand2 gate1176(.a(gate208inter12), .b(gate208inter1), .O(G687));
nand2 gate209( .a(G602), .b(G666), .O(G690) );
nand2 gate210( .a(G607), .b(G666), .O(G691) );
nand2 gate211( .a(G612), .b(G669), .O(G692) );
nand2 gate212( .a(G617), .b(G669), .O(G693) );

  xor2  gate1191(.a(G672), .b(G602), .O(gate213inter0));
  nand2 gate1192(.a(gate213inter0), .b(s_92), .O(gate213inter1));
  and2  gate1193(.a(G672), .b(G602), .O(gate213inter2));
  inv1  gate1194(.a(s_92), .O(gate213inter3));
  inv1  gate1195(.a(s_93), .O(gate213inter4));
  nand2 gate1196(.a(gate213inter4), .b(gate213inter3), .O(gate213inter5));
  nor2  gate1197(.a(gate213inter5), .b(gate213inter2), .O(gate213inter6));
  inv1  gate1198(.a(G602), .O(gate213inter7));
  inv1  gate1199(.a(G672), .O(gate213inter8));
  nand2 gate1200(.a(gate213inter8), .b(gate213inter7), .O(gate213inter9));
  nand2 gate1201(.a(s_93), .b(gate213inter3), .O(gate213inter10));
  nor2  gate1202(.a(gate213inter10), .b(gate213inter9), .O(gate213inter11));
  nor2  gate1203(.a(gate213inter11), .b(gate213inter6), .O(gate213inter12));
  nand2 gate1204(.a(gate213inter12), .b(gate213inter1), .O(G694));

  xor2  gate1835(.a(G672), .b(G612), .O(gate214inter0));
  nand2 gate1836(.a(gate214inter0), .b(s_184), .O(gate214inter1));
  and2  gate1837(.a(G672), .b(G612), .O(gate214inter2));
  inv1  gate1838(.a(s_184), .O(gate214inter3));
  inv1  gate1839(.a(s_185), .O(gate214inter4));
  nand2 gate1840(.a(gate214inter4), .b(gate214inter3), .O(gate214inter5));
  nor2  gate1841(.a(gate214inter5), .b(gate214inter2), .O(gate214inter6));
  inv1  gate1842(.a(G612), .O(gate214inter7));
  inv1  gate1843(.a(G672), .O(gate214inter8));
  nand2 gate1844(.a(gate214inter8), .b(gate214inter7), .O(gate214inter9));
  nand2 gate1845(.a(s_185), .b(gate214inter3), .O(gate214inter10));
  nor2  gate1846(.a(gate214inter10), .b(gate214inter9), .O(gate214inter11));
  nor2  gate1847(.a(gate214inter11), .b(gate214inter6), .O(gate214inter12));
  nand2 gate1848(.a(gate214inter12), .b(gate214inter1), .O(G695));
nand2 gate215( .a(G607), .b(G675), .O(G696) );

  xor2  gate1079(.a(G675), .b(G617), .O(gate216inter0));
  nand2 gate1080(.a(gate216inter0), .b(s_76), .O(gate216inter1));
  and2  gate1081(.a(G675), .b(G617), .O(gate216inter2));
  inv1  gate1082(.a(s_76), .O(gate216inter3));
  inv1  gate1083(.a(s_77), .O(gate216inter4));
  nand2 gate1084(.a(gate216inter4), .b(gate216inter3), .O(gate216inter5));
  nor2  gate1085(.a(gate216inter5), .b(gate216inter2), .O(gate216inter6));
  inv1  gate1086(.a(G617), .O(gate216inter7));
  inv1  gate1087(.a(G675), .O(gate216inter8));
  nand2 gate1088(.a(gate216inter8), .b(gate216inter7), .O(gate216inter9));
  nand2 gate1089(.a(s_77), .b(gate216inter3), .O(gate216inter10));
  nor2  gate1090(.a(gate216inter10), .b(gate216inter9), .O(gate216inter11));
  nor2  gate1091(.a(gate216inter11), .b(gate216inter6), .O(gate216inter12));
  nand2 gate1092(.a(gate216inter12), .b(gate216inter1), .O(G697));
nand2 gate217( .a(G622), .b(G678), .O(G698) );

  xor2  gate2661(.a(G678), .b(G627), .O(gate218inter0));
  nand2 gate2662(.a(gate218inter0), .b(s_302), .O(gate218inter1));
  and2  gate2663(.a(G678), .b(G627), .O(gate218inter2));
  inv1  gate2664(.a(s_302), .O(gate218inter3));
  inv1  gate2665(.a(s_303), .O(gate218inter4));
  nand2 gate2666(.a(gate218inter4), .b(gate218inter3), .O(gate218inter5));
  nor2  gate2667(.a(gate218inter5), .b(gate218inter2), .O(gate218inter6));
  inv1  gate2668(.a(G627), .O(gate218inter7));
  inv1  gate2669(.a(G678), .O(gate218inter8));
  nand2 gate2670(.a(gate218inter8), .b(gate218inter7), .O(gate218inter9));
  nand2 gate2671(.a(s_303), .b(gate218inter3), .O(gate218inter10));
  nor2  gate2672(.a(gate218inter10), .b(gate218inter9), .O(gate218inter11));
  nor2  gate2673(.a(gate218inter11), .b(gate218inter6), .O(gate218inter12));
  nand2 gate2674(.a(gate218inter12), .b(gate218inter1), .O(G699));

  xor2  gate1625(.a(G681), .b(G632), .O(gate219inter0));
  nand2 gate1626(.a(gate219inter0), .b(s_154), .O(gate219inter1));
  and2  gate1627(.a(G681), .b(G632), .O(gate219inter2));
  inv1  gate1628(.a(s_154), .O(gate219inter3));
  inv1  gate1629(.a(s_155), .O(gate219inter4));
  nand2 gate1630(.a(gate219inter4), .b(gate219inter3), .O(gate219inter5));
  nor2  gate1631(.a(gate219inter5), .b(gate219inter2), .O(gate219inter6));
  inv1  gate1632(.a(G632), .O(gate219inter7));
  inv1  gate1633(.a(G681), .O(gate219inter8));
  nand2 gate1634(.a(gate219inter8), .b(gate219inter7), .O(gate219inter9));
  nand2 gate1635(.a(s_155), .b(gate219inter3), .O(gate219inter10));
  nor2  gate1636(.a(gate219inter10), .b(gate219inter9), .O(gate219inter11));
  nor2  gate1637(.a(gate219inter11), .b(gate219inter6), .O(gate219inter12));
  nand2 gate1638(.a(gate219inter12), .b(gate219inter1), .O(G700));

  xor2  gate2381(.a(G681), .b(G637), .O(gate220inter0));
  nand2 gate2382(.a(gate220inter0), .b(s_262), .O(gate220inter1));
  and2  gate2383(.a(G681), .b(G637), .O(gate220inter2));
  inv1  gate2384(.a(s_262), .O(gate220inter3));
  inv1  gate2385(.a(s_263), .O(gate220inter4));
  nand2 gate2386(.a(gate220inter4), .b(gate220inter3), .O(gate220inter5));
  nor2  gate2387(.a(gate220inter5), .b(gate220inter2), .O(gate220inter6));
  inv1  gate2388(.a(G637), .O(gate220inter7));
  inv1  gate2389(.a(G681), .O(gate220inter8));
  nand2 gate2390(.a(gate220inter8), .b(gate220inter7), .O(gate220inter9));
  nand2 gate2391(.a(s_263), .b(gate220inter3), .O(gate220inter10));
  nor2  gate2392(.a(gate220inter10), .b(gate220inter9), .O(gate220inter11));
  nor2  gate2393(.a(gate220inter11), .b(gate220inter6), .O(gate220inter12));
  nand2 gate2394(.a(gate220inter12), .b(gate220inter1), .O(G701));
nand2 gate221( .a(G622), .b(G684), .O(G702) );
nand2 gate222( .a(G632), .b(G684), .O(G703) );
nand2 gate223( .a(G627), .b(G687), .O(G704) );

  xor2  gate659(.a(G687), .b(G637), .O(gate224inter0));
  nand2 gate660(.a(gate224inter0), .b(s_16), .O(gate224inter1));
  and2  gate661(.a(G687), .b(G637), .O(gate224inter2));
  inv1  gate662(.a(s_16), .O(gate224inter3));
  inv1  gate663(.a(s_17), .O(gate224inter4));
  nand2 gate664(.a(gate224inter4), .b(gate224inter3), .O(gate224inter5));
  nor2  gate665(.a(gate224inter5), .b(gate224inter2), .O(gate224inter6));
  inv1  gate666(.a(G637), .O(gate224inter7));
  inv1  gate667(.a(G687), .O(gate224inter8));
  nand2 gate668(.a(gate224inter8), .b(gate224inter7), .O(gate224inter9));
  nand2 gate669(.a(s_17), .b(gate224inter3), .O(gate224inter10));
  nor2  gate670(.a(gate224inter10), .b(gate224inter9), .O(gate224inter11));
  nor2  gate671(.a(gate224inter11), .b(gate224inter6), .O(gate224inter12));
  nand2 gate672(.a(gate224inter12), .b(gate224inter1), .O(G705));
nand2 gate225( .a(G690), .b(G691), .O(G706) );

  xor2  gate1597(.a(G693), .b(G692), .O(gate226inter0));
  nand2 gate1598(.a(gate226inter0), .b(s_150), .O(gate226inter1));
  and2  gate1599(.a(G693), .b(G692), .O(gate226inter2));
  inv1  gate1600(.a(s_150), .O(gate226inter3));
  inv1  gate1601(.a(s_151), .O(gate226inter4));
  nand2 gate1602(.a(gate226inter4), .b(gate226inter3), .O(gate226inter5));
  nor2  gate1603(.a(gate226inter5), .b(gate226inter2), .O(gate226inter6));
  inv1  gate1604(.a(G692), .O(gate226inter7));
  inv1  gate1605(.a(G693), .O(gate226inter8));
  nand2 gate1606(.a(gate226inter8), .b(gate226inter7), .O(gate226inter9));
  nand2 gate1607(.a(s_151), .b(gate226inter3), .O(gate226inter10));
  nor2  gate1608(.a(gate226inter10), .b(gate226inter9), .O(gate226inter11));
  nor2  gate1609(.a(gate226inter11), .b(gate226inter6), .O(gate226inter12));
  nand2 gate1610(.a(gate226inter12), .b(gate226inter1), .O(G709));

  xor2  gate673(.a(G695), .b(G694), .O(gate227inter0));
  nand2 gate674(.a(gate227inter0), .b(s_18), .O(gate227inter1));
  and2  gate675(.a(G695), .b(G694), .O(gate227inter2));
  inv1  gate676(.a(s_18), .O(gate227inter3));
  inv1  gate677(.a(s_19), .O(gate227inter4));
  nand2 gate678(.a(gate227inter4), .b(gate227inter3), .O(gate227inter5));
  nor2  gate679(.a(gate227inter5), .b(gate227inter2), .O(gate227inter6));
  inv1  gate680(.a(G694), .O(gate227inter7));
  inv1  gate681(.a(G695), .O(gate227inter8));
  nand2 gate682(.a(gate227inter8), .b(gate227inter7), .O(gate227inter9));
  nand2 gate683(.a(s_19), .b(gate227inter3), .O(gate227inter10));
  nor2  gate684(.a(gate227inter10), .b(gate227inter9), .O(gate227inter11));
  nor2  gate685(.a(gate227inter11), .b(gate227inter6), .O(gate227inter12));
  nand2 gate686(.a(gate227inter12), .b(gate227inter1), .O(G712));

  xor2  gate1877(.a(G697), .b(G696), .O(gate228inter0));
  nand2 gate1878(.a(gate228inter0), .b(s_190), .O(gate228inter1));
  and2  gate1879(.a(G697), .b(G696), .O(gate228inter2));
  inv1  gate1880(.a(s_190), .O(gate228inter3));
  inv1  gate1881(.a(s_191), .O(gate228inter4));
  nand2 gate1882(.a(gate228inter4), .b(gate228inter3), .O(gate228inter5));
  nor2  gate1883(.a(gate228inter5), .b(gate228inter2), .O(gate228inter6));
  inv1  gate1884(.a(G696), .O(gate228inter7));
  inv1  gate1885(.a(G697), .O(gate228inter8));
  nand2 gate1886(.a(gate228inter8), .b(gate228inter7), .O(gate228inter9));
  nand2 gate1887(.a(s_191), .b(gate228inter3), .O(gate228inter10));
  nor2  gate1888(.a(gate228inter10), .b(gate228inter9), .O(gate228inter11));
  nor2  gate1889(.a(gate228inter11), .b(gate228inter6), .O(gate228inter12));
  nand2 gate1890(.a(gate228inter12), .b(gate228inter1), .O(G715));

  xor2  gate813(.a(G699), .b(G698), .O(gate229inter0));
  nand2 gate814(.a(gate229inter0), .b(s_38), .O(gate229inter1));
  and2  gate815(.a(G699), .b(G698), .O(gate229inter2));
  inv1  gate816(.a(s_38), .O(gate229inter3));
  inv1  gate817(.a(s_39), .O(gate229inter4));
  nand2 gate818(.a(gate229inter4), .b(gate229inter3), .O(gate229inter5));
  nor2  gate819(.a(gate229inter5), .b(gate229inter2), .O(gate229inter6));
  inv1  gate820(.a(G698), .O(gate229inter7));
  inv1  gate821(.a(G699), .O(gate229inter8));
  nand2 gate822(.a(gate229inter8), .b(gate229inter7), .O(gate229inter9));
  nand2 gate823(.a(s_39), .b(gate229inter3), .O(gate229inter10));
  nor2  gate824(.a(gate229inter10), .b(gate229inter9), .O(gate229inter11));
  nor2  gate825(.a(gate229inter11), .b(gate229inter6), .O(gate229inter12));
  nand2 gate826(.a(gate229inter12), .b(gate229inter1), .O(G718));

  xor2  gate1359(.a(G701), .b(G700), .O(gate230inter0));
  nand2 gate1360(.a(gate230inter0), .b(s_116), .O(gate230inter1));
  and2  gate1361(.a(G701), .b(G700), .O(gate230inter2));
  inv1  gate1362(.a(s_116), .O(gate230inter3));
  inv1  gate1363(.a(s_117), .O(gate230inter4));
  nand2 gate1364(.a(gate230inter4), .b(gate230inter3), .O(gate230inter5));
  nor2  gate1365(.a(gate230inter5), .b(gate230inter2), .O(gate230inter6));
  inv1  gate1366(.a(G700), .O(gate230inter7));
  inv1  gate1367(.a(G701), .O(gate230inter8));
  nand2 gate1368(.a(gate230inter8), .b(gate230inter7), .O(gate230inter9));
  nand2 gate1369(.a(s_117), .b(gate230inter3), .O(gate230inter10));
  nor2  gate1370(.a(gate230inter10), .b(gate230inter9), .O(gate230inter11));
  nor2  gate1371(.a(gate230inter11), .b(gate230inter6), .O(gate230inter12));
  nand2 gate1372(.a(gate230inter12), .b(gate230inter1), .O(G721));

  xor2  gate2563(.a(G703), .b(G702), .O(gate231inter0));
  nand2 gate2564(.a(gate231inter0), .b(s_288), .O(gate231inter1));
  and2  gate2565(.a(G703), .b(G702), .O(gate231inter2));
  inv1  gate2566(.a(s_288), .O(gate231inter3));
  inv1  gate2567(.a(s_289), .O(gate231inter4));
  nand2 gate2568(.a(gate231inter4), .b(gate231inter3), .O(gate231inter5));
  nor2  gate2569(.a(gate231inter5), .b(gate231inter2), .O(gate231inter6));
  inv1  gate2570(.a(G702), .O(gate231inter7));
  inv1  gate2571(.a(G703), .O(gate231inter8));
  nand2 gate2572(.a(gate231inter8), .b(gate231inter7), .O(gate231inter9));
  nand2 gate2573(.a(s_289), .b(gate231inter3), .O(gate231inter10));
  nor2  gate2574(.a(gate231inter10), .b(gate231inter9), .O(gate231inter11));
  nor2  gate2575(.a(gate231inter11), .b(gate231inter6), .O(gate231inter12));
  nand2 gate2576(.a(gate231inter12), .b(gate231inter1), .O(G724));

  xor2  gate1387(.a(G705), .b(G704), .O(gate232inter0));
  nand2 gate1388(.a(gate232inter0), .b(s_120), .O(gate232inter1));
  and2  gate1389(.a(G705), .b(G704), .O(gate232inter2));
  inv1  gate1390(.a(s_120), .O(gate232inter3));
  inv1  gate1391(.a(s_121), .O(gate232inter4));
  nand2 gate1392(.a(gate232inter4), .b(gate232inter3), .O(gate232inter5));
  nor2  gate1393(.a(gate232inter5), .b(gate232inter2), .O(gate232inter6));
  inv1  gate1394(.a(G704), .O(gate232inter7));
  inv1  gate1395(.a(G705), .O(gate232inter8));
  nand2 gate1396(.a(gate232inter8), .b(gate232inter7), .O(gate232inter9));
  nand2 gate1397(.a(s_121), .b(gate232inter3), .O(gate232inter10));
  nor2  gate1398(.a(gate232inter10), .b(gate232inter9), .O(gate232inter11));
  nor2  gate1399(.a(gate232inter11), .b(gate232inter6), .O(gate232inter12));
  nand2 gate1400(.a(gate232inter12), .b(gate232inter1), .O(G727));

  xor2  gate1485(.a(G718), .b(G242), .O(gate233inter0));
  nand2 gate1486(.a(gate233inter0), .b(s_134), .O(gate233inter1));
  and2  gate1487(.a(G718), .b(G242), .O(gate233inter2));
  inv1  gate1488(.a(s_134), .O(gate233inter3));
  inv1  gate1489(.a(s_135), .O(gate233inter4));
  nand2 gate1490(.a(gate233inter4), .b(gate233inter3), .O(gate233inter5));
  nor2  gate1491(.a(gate233inter5), .b(gate233inter2), .O(gate233inter6));
  inv1  gate1492(.a(G242), .O(gate233inter7));
  inv1  gate1493(.a(G718), .O(gate233inter8));
  nand2 gate1494(.a(gate233inter8), .b(gate233inter7), .O(gate233inter9));
  nand2 gate1495(.a(s_135), .b(gate233inter3), .O(gate233inter10));
  nor2  gate1496(.a(gate233inter10), .b(gate233inter9), .O(gate233inter11));
  nor2  gate1497(.a(gate233inter11), .b(gate233inter6), .O(gate233inter12));
  nand2 gate1498(.a(gate233inter12), .b(gate233inter1), .O(G730));
nand2 gate234( .a(G245), .b(G721), .O(G733) );
nand2 gate235( .a(G248), .b(G724), .O(G736) );

  xor2  gate2143(.a(G727), .b(G251), .O(gate236inter0));
  nand2 gate2144(.a(gate236inter0), .b(s_228), .O(gate236inter1));
  and2  gate2145(.a(G727), .b(G251), .O(gate236inter2));
  inv1  gate2146(.a(s_228), .O(gate236inter3));
  inv1  gate2147(.a(s_229), .O(gate236inter4));
  nand2 gate2148(.a(gate236inter4), .b(gate236inter3), .O(gate236inter5));
  nor2  gate2149(.a(gate236inter5), .b(gate236inter2), .O(gate236inter6));
  inv1  gate2150(.a(G251), .O(gate236inter7));
  inv1  gate2151(.a(G727), .O(gate236inter8));
  nand2 gate2152(.a(gate236inter8), .b(gate236inter7), .O(gate236inter9));
  nand2 gate2153(.a(s_229), .b(gate236inter3), .O(gate236inter10));
  nor2  gate2154(.a(gate236inter10), .b(gate236inter9), .O(gate236inter11));
  nor2  gate2155(.a(gate236inter11), .b(gate236inter6), .O(gate236inter12));
  nand2 gate2156(.a(gate236inter12), .b(gate236inter1), .O(G739));
nand2 gate237( .a(G254), .b(G706), .O(G742) );

  xor2  gate2185(.a(G709), .b(G257), .O(gate238inter0));
  nand2 gate2186(.a(gate238inter0), .b(s_234), .O(gate238inter1));
  and2  gate2187(.a(G709), .b(G257), .O(gate238inter2));
  inv1  gate2188(.a(s_234), .O(gate238inter3));
  inv1  gate2189(.a(s_235), .O(gate238inter4));
  nand2 gate2190(.a(gate238inter4), .b(gate238inter3), .O(gate238inter5));
  nor2  gate2191(.a(gate238inter5), .b(gate238inter2), .O(gate238inter6));
  inv1  gate2192(.a(G257), .O(gate238inter7));
  inv1  gate2193(.a(G709), .O(gate238inter8));
  nand2 gate2194(.a(gate238inter8), .b(gate238inter7), .O(gate238inter9));
  nand2 gate2195(.a(s_235), .b(gate238inter3), .O(gate238inter10));
  nor2  gate2196(.a(gate238inter10), .b(gate238inter9), .O(gate238inter11));
  nor2  gate2197(.a(gate238inter11), .b(gate238inter6), .O(gate238inter12));
  nand2 gate2198(.a(gate238inter12), .b(gate238inter1), .O(G745));

  xor2  gate2129(.a(G712), .b(G260), .O(gate239inter0));
  nand2 gate2130(.a(gate239inter0), .b(s_226), .O(gate239inter1));
  and2  gate2131(.a(G712), .b(G260), .O(gate239inter2));
  inv1  gate2132(.a(s_226), .O(gate239inter3));
  inv1  gate2133(.a(s_227), .O(gate239inter4));
  nand2 gate2134(.a(gate239inter4), .b(gate239inter3), .O(gate239inter5));
  nor2  gate2135(.a(gate239inter5), .b(gate239inter2), .O(gate239inter6));
  inv1  gate2136(.a(G260), .O(gate239inter7));
  inv1  gate2137(.a(G712), .O(gate239inter8));
  nand2 gate2138(.a(gate239inter8), .b(gate239inter7), .O(gate239inter9));
  nand2 gate2139(.a(s_227), .b(gate239inter3), .O(gate239inter10));
  nor2  gate2140(.a(gate239inter10), .b(gate239inter9), .O(gate239inter11));
  nor2  gate2141(.a(gate239inter11), .b(gate239inter6), .O(gate239inter12));
  nand2 gate2142(.a(gate239inter12), .b(gate239inter1), .O(G748));
nand2 gate240( .a(G263), .b(G715), .O(G751) );

  xor2  gate2451(.a(G730), .b(G242), .O(gate241inter0));
  nand2 gate2452(.a(gate241inter0), .b(s_272), .O(gate241inter1));
  and2  gate2453(.a(G730), .b(G242), .O(gate241inter2));
  inv1  gate2454(.a(s_272), .O(gate241inter3));
  inv1  gate2455(.a(s_273), .O(gate241inter4));
  nand2 gate2456(.a(gate241inter4), .b(gate241inter3), .O(gate241inter5));
  nor2  gate2457(.a(gate241inter5), .b(gate241inter2), .O(gate241inter6));
  inv1  gate2458(.a(G242), .O(gate241inter7));
  inv1  gate2459(.a(G730), .O(gate241inter8));
  nand2 gate2460(.a(gate241inter8), .b(gate241inter7), .O(gate241inter9));
  nand2 gate2461(.a(s_273), .b(gate241inter3), .O(gate241inter10));
  nor2  gate2462(.a(gate241inter10), .b(gate241inter9), .O(gate241inter11));
  nor2  gate2463(.a(gate241inter11), .b(gate241inter6), .O(gate241inter12));
  nand2 gate2464(.a(gate241inter12), .b(gate241inter1), .O(G754));
nand2 gate242( .a(G718), .b(G730), .O(G755) );
nand2 gate243( .a(G245), .b(G733), .O(G756) );
nand2 gate244( .a(G721), .b(G733), .O(G757) );

  xor2  gate2577(.a(G736), .b(G248), .O(gate245inter0));
  nand2 gate2578(.a(gate245inter0), .b(s_290), .O(gate245inter1));
  and2  gate2579(.a(G736), .b(G248), .O(gate245inter2));
  inv1  gate2580(.a(s_290), .O(gate245inter3));
  inv1  gate2581(.a(s_291), .O(gate245inter4));
  nand2 gate2582(.a(gate245inter4), .b(gate245inter3), .O(gate245inter5));
  nor2  gate2583(.a(gate245inter5), .b(gate245inter2), .O(gate245inter6));
  inv1  gate2584(.a(G248), .O(gate245inter7));
  inv1  gate2585(.a(G736), .O(gate245inter8));
  nand2 gate2586(.a(gate245inter8), .b(gate245inter7), .O(gate245inter9));
  nand2 gate2587(.a(s_291), .b(gate245inter3), .O(gate245inter10));
  nor2  gate2588(.a(gate245inter10), .b(gate245inter9), .O(gate245inter11));
  nor2  gate2589(.a(gate245inter11), .b(gate245inter6), .O(gate245inter12));
  nand2 gate2590(.a(gate245inter12), .b(gate245inter1), .O(G758));
nand2 gate246( .a(G724), .b(G736), .O(G759) );

  xor2  gate2045(.a(G739), .b(G251), .O(gate247inter0));
  nand2 gate2046(.a(gate247inter0), .b(s_214), .O(gate247inter1));
  and2  gate2047(.a(G739), .b(G251), .O(gate247inter2));
  inv1  gate2048(.a(s_214), .O(gate247inter3));
  inv1  gate2049(.a(s_215), .O(gate247inter4));
  nand2 gate2050(.a(gate247inter4), .b(gate247inter3), .O(gate247inter5));
  nor2  gate2051(.a(gate247inter5), .b(gate247inter2), .O(gate247inter6));
  inv1  gate2052(.a(G251), .O(gate247inter7));
  inv1  gate2053(.a(G739), .O(gate247inter8));
  nand2 gate2054(.a(gate247inter8), .b(gate247inter7), .O(gate247inter9));
  nand2 gate2055(.a(s_215), .b(gate247inter3), .O(gate247inter10));
  nor2  gate2056(.a(gate247inter10), .b(gate247inter9), .O(gate247inter11));
  nor2  gate2057(.a(gate247inter11), .b(gate247inter6), .O(gate247inter12));
  nand2 gate2058(.a(gate247inter12), .b(gate247inter1), .O(G760));

  xor2  gate757(.a(G739), .b(G727), .O(gate248inter0));
  nand2 gate758(.a(gate248inter0), .b(s_30), .O(gate248inter1));
  and2  gate759(.a(G739), .b(G727), .O(gate248inter2));
  inv1  gate760(.a(s_30), .O(gate248inter3));
  inv1  gate761(.a(s_31), .O(gate248inter4));
  nand2 gate762(.a(gate248inter4), .b(gate248inter3), .O(gate248inter5));
  nor2  gate763(.a(gate248inter5), .b(gate248inter2), .O(gate248inter6));
  inv1  gate764(.a(G727), .O(gate248inter7));
  inv1  gate765(.a(G739), .O(gate248inter8));
  nand2 gate766(.a(gate248inter8), .b(gate248inter7), .O(gate248inter9));
  nand2 gate767(.a(s_31), .b(gate248inter3), .O(gate248inter10));
  nor2  gate768(.a(gate248inter10), .b(gate248inter9), .O(gate248inter11));
  nor2  gate769(.a(gate248inter11), .b(gate248inter6), .O(gate248inter12));
  nand2 gate770(.a(gate248inter12), .b(gate248inter1), .O(G761));
nand2 gate249( .a(G254), .b(G742), .O(G762) );
nand2 gate250( .a(G706), .b(G742), .O(G763) );

  xor2  gate2241(.a(G745), .b(G257), .O(gate251inter0));
  nand2 gate2242(.a(gate251inter0), .b(s_242), .O(gate251inter1));
  and2  gate2243(.a(G745), .b(G257), .O(gate251inter2));
  inv1  gate2244(.a(s_242), .O(gate251inter3));
  inv1  gate2245(.a(s_243), .O(gate251inter4));
  nand2 gate2246(.a(gate251inter4), .b(gate251inter3), .O(gate251inter5));
  nor2  gate2247(.a(gate251inter5), .b(gate251inter2), .O(gate251inter6));
  inv1  gate2248(.a(G257), .O(gate251inter7));
  inv1  gate2249(.a(G745), .O(gate251inter8));
  nand2 gate2250(.a(gate251inter8), .b(gate251inter7), .O(gate251inter9));
  nand2 gate2251(.a(s_243), .b(gate251inter3), .O(gate251inter10));
  nor2  gate2252(.a(gate251inter10), .b(gate251inter9), .O(gate251inter11));
  nor2  gate2253(.a(gate251inter11), .b(gate251inter6), .O(gate251inter12));
  nand2 gate2254(.a(gate251inter12), .b(gate251inter1), .O(G764));
nand2 gate252( .a(G709), .b(G745), .O(G765) );

  xor2  gate1023(.a(G748), .b(G260), .O(gate253inter0));
  nand2 gate1024(.a(gate253inter0), .b(s_68), .O(gate253inter1));
  and2  gate1025(.a(G748), .b(G260), .O(gate253inter2));
  inv1  gate1026(.a(s_68), .O(gate253inter3));
  inv1  gate1027(.a(s_69), .O(gate253inter4));
  nand2 gate1028(.a(gate253inter4), .b(gate253inter3), .O(gate253inter5));
  nor2  gate1029(.a(gate253inter5), .b(gate253inter2), .O(gate253inter6));
  inv1  gate1030(.a(G260), .O(gate253inter7));
  inv1  gate1031(.a(G748), .O(gate253inter8));
  nand2 gate1032(.a(gate253inter8), .b(gate253inter7), .O(gate253inter9));
  nand2 gate1033(.a(s_69), .b(gate253inter3), .O(gate253inter10));
  nor2  gate1034(.a(gate253inter10), .b(gate253inter9), .O(gate253inter11));
  nor2  gate1035(.a(gate253inter11), .b(gate253inter6), .O(gate253inter12));
  nand2 gate1036(.a(gate253inter12), .b(gate253inter1), .O(G766));
nand2 gate254( .a(G712), .b(G748), .O(G767) );

  xor2  gate2031(.a(G751), .b(G263), .O(gate255inter0));
  nand2 gate2032(.a(gate255inter0), .b(s_212), .O(gate255inter1));
  and2  gate2033(.a(G751), .b(G263), .O(gate255inter2));
  inv1  gate2034(.a(s_212), .O(gate255inter3));
  inv1  gate2035(.a(s_213), .O(gate255inter4));
  nand2 gate2036(.a(gate255inter4), .b(gate255inter3), .O(gate255inter5));
  nor2  gate2037(.a(gate255inter5), .b(gate255inter2), .O(gate255inter6));
  inv1  gate2038(.a(G263), .O(gate255inter7));
  inv1  gate2039(.a(G751), .O(gate255inter8));
  nand2 gate2040(.a(gate255inter8), .b(gate255inter7), .O(gate255inter9));
  nand2 gate2041(.a(s_213), .b(gate255inter3), .O(gate255inter10));
  nor2  gate2042(.a(gate255inter10), .b(gate255inter9), .O(gate255inter11));
  nor2  gate2043(.a(gate255inter11), .b(gate255inter6), .O(gate255inter12));
  nand2 gate2044(.a(gate255inter12), .b(gate255inter1), .O(G768));
nand2 gate256( .a(G715), .b(G751), .O(G769) );

  xor2  gate589(.a(G755), .b(G754), .O(gate257inter0));
  nand2 gate590(.a(gate257inter0), .b(s_6), .O(gate257inter1));
  and2  gate591(.a(G755), .b(G754), .O(gate257inter2));
  inv1  gate592(.a(s_6), .O(gate257inter3));
  inv1  gate593(.a(s_7), .O(gate257inter4));
  nand2 gate594(.a(gate257inter4), .b(gate257inter3), .O(gate257inter5));
  nor2  gate595(.a(gate257inter5), .b(gate257inter2), .O(gate257inter6));
  inv1  gate596(.a(G754), .O(gate257inter7));
  inv1  gate597(.a(G755), .O(gate257inter8));
  nand2 gate598(.a(gate257inter8), .b(gate257inter7), .O(gate257inter9));
  nand2 gate599(.a(s_7), .b(gate257inter3), .O(gate257inter10));
  nor2  gate600(.a(gate257inter10), .b(gate257inter9), .O(gate257inter11));
  nor2  gate601(.a(gate257inter11), .b(gate257inter6), .O(gate257inter12));
  nand2 gate602(.a(gate257inter12), .b(gate257inter1), .O(G770));
nand2 gate258( .a(G756), .b(G757), .O(G773) );
nand2 gate259( .a(G758), .b(G759), .O(G776) );
nand2 gate260( .a(G760), .b(G761), .O(G779) );

  xor2  gate1443(.a(G763), .b(G762), .O(gate261inter0));
  nand2 gate1444(.a(gate261inter0), .b(s_128), .O(gate261inter1));
  and2  gate1445(.a(G763), .b(G762), .O(gate261inter2));
  inv1  gate1446(.a(s_128), .O(gate261inter3));
  inv1  gate1447(.a(s_129), .O(gate261inter4));
  nand2 gate1448(.a(gate261inter4), .b(gate261inter3), .O(gate261inter5));
  nor2  gate1449(.a(gate261inter5), .b(gate261inter2), .O(gate261inter6));
  inv1  gate1450(.a(G762), .O(gate261inter7));
  inv1  gate1451(.a(G763), .O(gate261inter8));
  nand2 gate1452(.a(gate261inter8), .b(gate261inter7), .O(gate261inter9));
  nand2 gate1453(.a(s_129), .b(gate261inter3), .O(gate261inter10));
  nor2  gate1454(.a(gate261inter10), .b(gate261inter9), .O(gate261inter11));
  nor2  gate1455(.a(gate261inter11), .b(gate261inter6), .O(gate261inter12));
  nand2 gate1456(.a(gate261inter12), .b(gate261inter1), .O(G782));

  xor2  gate2171(.a(G765), .b(G764), .O(gate262inter0));
  nand2 gate2172(.a(gate262inter0), .b(s_232), .O(gate262inter1));
  and2  gate2173(.a(G765), .b(G764), .O(gate262inter2));
  inv1  gate2174(.a(s_232), .O(gate262inter3));
  inv1  gate2175(.a(s_233), .O(gate262inter4));
  nand2 gate2176(.a(gate262inter4), .b(gate262inter3), .O(gate262inter5));
  nor2  gate2177(.a(gate262inter5), .b(gate262inter2), .O(gate262inter6));
  inv1  gate2178(.a(G764), .O(gate262inter7));
  inv1  gate2179(.a(G765), .O(gate262inter8));
  nand2 gate2180(.a(gate262inter8), .b(gate262inter7), .O(gate262inter9));
  nand2 gate2181(.a(s_233), .b(gate262inter3), .O(gate262inter10));
  nor2  gate2182(.a(gate262inter10), .b(gate262inter9), .O(gate262inter11));
  nor2  gate2183(.a(gate262inter11), .b(gate262inter6), .O(gate262inter12));
  nand2 gate2184(.a(gate262inter12), .b(gate262inter1), .O(G785));
nand2 gate263( .a(G766), .b(G767), .O(G788) );
nand2 gate264( .a(G768), .b(G769), .O(G791) );
nand2 gate265( .a(G642), .b(G770), .O(G794) );
nand2 gate266( .a(G645), .b(G773), .O(G797) );
nand2 gate267( .a(G648), .b(G776), .O(G800) );

  xor2  gate2283(.a(G779), .b(G651), .O(gate268inter0));
  nand2 gate2284(.a(gate268inter0), .b(s_248), .O(gate268inter1));
  and2  gate2285(.a(G779), .b(G651), .O(gate268inter2));
  inv1  gate2286(.a(s_248), .O(gate268inter3));
  inv1  gate2287(.a(s_249), .O(gate268inter4));
  nand2 gate2288(.a(gate268inter4), .b(gate268inter3), .O(gate268inter5));
  nor2  gate2289(.a(gate268inter5), .b(gate268inter2), .O(gate268inter6));
  inv1  gate2290(.a(G651), .O(gate268inter7));
  inv1  gate2291(.a(G779), .O(gate268inter8));
  nand2 gate2292(.a(gate268inter8), .b(gate268inter7), .O(gate268inter9));
  nand2 gate2293(.a(s_249), .b(gate268inter3), .O(gate268inter10));
  nor2  gate2294(.a(gate268inter10), .b(gate268inter9), .O(gate268inter11));
  nor2  gate2295(.a(gate268inter11), .b(gate268inter6), .O(gate268inter12));
  nand2 gate2296(.a(gate268inter12), .b(gate268inter1), .O(G803));

  xor2  gate2507(.a(G782), .b(G654), .O(gate269inter0));
  nand2 gate2508(.a(gate269inter0), .b(s_280), .O(gate269inter1));
  and2  gate2509(.a(G782), .b(G654), .O(gate269inter2));
  inv1  gate2510(.a(s_280), .O(gate269inter3));
  inv1  gate2511(.a(s_281), .O(gate269inter4));
  nand2 gate2512(.a(gate269inter4), .b(gate269inter3), .O(gate269inter5));
  nor2  gate2513(.a(gate269inter5), .b(gate269inter2), .O(gate269inter6));
  inv1  gate2514(.a(G654), .O(gate269inter7));
  inv1  gate2515(.a(G782), .O(gate269inter8));
  nand2 gate2516(.a(gate269inter8), .b(gate269inter7), .O(gate269inter9));
  nand2 gate2517(.a(s_281), .b(gate269inter3), .O(gate269inter10));
  nor2  gate2518(.a(gate269inter10), .b(gate269inter9), .O(gate269inter11));
  nor2  gate2519(.a(gate269inter11), .b(gate269inter6), .O(gate269inter12));
  nand2 gate2520(.a(gate269inter12), .b(gate269inter1), .O(G806));
nand2 gate270( .a(G657), .b(G785), .O(G809) );

  xor2  gate575(.a(G788), .b(G660), .O(gate271inter0));
  nand2 gate576(.a(gate271inter0), .b(s_4), .O(gate271inter1));
  and2  gate577(.a(G788), .b(G660), .O(gate271inter2));
  inv1  gate578(.a(s_4), .O(gate271inter3));
  inv1  gate579(.a(s_5), .O(gate271inter4));
  nand2 gate580(.a(gate271inter4), .b(gate271inter3), .O(gate271inter5));
  nor2  gate581(.a(gate271inter5), .b(gate271inter2), .O(gate271inter6));
  inv1  gate582(.a(G660), .O(gate271inter7));
  inv1  gate583(.a(G788), .O(gate271inter8));
  nand2 gate584(.a(gate271inter8), .b(gate271inter7), .O(gate271inter9));
  nand2 gate585(.a(s_5), .b(gate271inter3), .O(gate271inter10));
  nor2  gate586(.a(gate271inter10), .b(gate271inter9), .O(gate271inter11));
  nor2  gate587(.a(gate271inter11), .b(gate271inter6), .O(gate271inter12));
  nand2 gate588(.a(gate271inter12), .b(gate271inter1), .O(G812));
nand2 gate272( .a(G663), .b(G791), .O(G815) );
nand2 gate273( .a(G642), .b(G794), .O(G818) );
nand2 gate274( .a(G770), .b(G794), .O(G819) );

  xor2  gate2073(.a(G797), .b(G645), .O(gate275inter0));
  nand2 gate2074(.a(gate275inter0), .b(s_218), .O(gate275inter1));
  and2  gate2075(.a(G797), .b(G645), .O(gate275inter2));
  inv1  gate2076(.a(s_218), .O(gate275inter3));
  inv1  gate2077(.a(s_219), .O(gate275inter4));
  nand2 gate2078(.a(gate275inter4), .b(gate275inter3), .O(gate275inter5));
  nor2  gate2079(.a(gate275inter5), .b(gate275inter2), .O(gate275inter6));
  inv1  gate2080(.a(G645), .O(gate275inter7));
  inv1  gate2081(.a(G797), .O(gate275inter8));
  nand2 gate2082(.a(gate275inter8), .b(gate275inter7), .O(gate275inter9));
  nand2 gate2083(.a(s_219), .b(gate275inter3), .O(gate275inter10));
  nor2  gate2084(.a(gate275inter10), .b(gate275inter9), .O(gate275inter11));
  nor2  gate2085(.a(gate275inter11), .b(gate275inter6), .O(gate275inter12));
  nand2 gate2086(.a(gate275inter12), .b(gate275inter1), .O(G820));
nand2 gate276( .a(G773), .b(G797), .O(G821) );
nand2 gate277( .a(G648), .b(G800), .O(G822) );
nand2 gate278( .a(G776), .b(G800), .O(G823) );
nand2 gate279( .a(G651), .b(G803), .O(G824) );
nand2 gate280( .a(G779), .b(G803), .O(G825) );
nand2 gate281( .a(G654), .b(G806), .O(G826) );
nand2 gate282( .a(G782), .b(G806), .O(G827) );
nand2 gate283( .a(G657), .b(G809), .O(G828) );
nand2 gate284( .a(G785), .b(G809), .O(G829) );
nand2 gate285( .a(G660), .b(G812), .O(G830) );

  xor2  gate2493(.a(G812), .b(G788), .O(gate286inter0));
  nand2 gate2494(.a(gate286inter0), .b(s_278), .O(gate286inter1));
  and2  gate2495(.a(G812), .b(G788), .O(gate286inter2));
  inv1  gate2496(.a(s_278), .O(gate286inter3));
  inv1  gate2497(.a(s_279), .O(gate286inter4));
  nand2 gate2498(.a(gate286inter4), .b(gate286inter3), .O(gate286inter5));
  nor2  gate2499(.a(gate286inter5), .b(gate286inter2), .O(gate286inter6));
  inv1  gate2500(.a(G788), .O(gate286inter7));
  inv1  gate2501(.a(G812), .O(gate286inter8));
  nand2 gate2502(.a(gate286inter8), .b(gate286inter7), .O(gate286inter9));
  nand2 gate2503(.a(s_279), .b(gate286inter3), .O(gate286inter10));
  nor2  gate2504(.a(gate286inter10), .b(gate286inter9), .O(gate286inter11));
  nor2  gate2505(.a(gate286inter11), .b(gate286inter6), .O(gate286inter12));
  nand2 gate2506(.a(gate286inter12), .b(gate286inter1), .O(G831));
nand2 gate287( .a(G663), .b(G815), .O(G832) );
nand2 gate288( .a(G791), .b(G815), .O(G833) );

  xor2  gate1681(.a(G819), .b(G818), .O(gate289inter0));
  nand2 gate1682(.a(gate289inter0), .b(s_162), .O(gate289inter1));
  and2  gate1683(.a(G819), .b(G818), .O(gate289inter2));
  inv1  gate1684(.a(s_162), .O(gate289inter3));
  inv1  gate1685(.a(s_163), .O(gate289inter4));
  nand2 gate1686(.a(gate289inter4), .b(gate289inter3), .O(gate289inter5));
  nor2  gate1687(.a(gate289inter5), .b(gate289inter2), .O(gate289inter6));
  inv1  gate1688(.a(G818), .O(gate289inter7));
  inv1  gate1689(.a(G819), .O(gate289inter8));
  nand2 gate1690(.a(gate289inter8), .b(gate289inter7), .O(gate289inter9));
  nand2 gate1691(.a(s_163), .b(gate289inter3), .O(gate289inter10));
  nor2  gate1692(.a(gate289inter10), .b(gate289inter9), .O(gate289inter11));
  nor2  gate1693(.a(gate289inter11), .b(gate289inter6), .O(gate289inter12));
  nand2 gate1694(.a(gate289inter12), .b(gate289inter1), .O(G834));

  xor2  gate2101(.a(G821), .b(G820), .O(gate290inter0));
  nand2 gate2102(.a(gate290inter0), .b(s_222), .O(gate290inter1));
  and2  gate2103(.a(G821), .b(G820), .O(gate290inter2));
  inv1  gate2104(.a(s_222), .O(gate290inter3));
  inv1  gate2105(.a(s_223), .O(gate290inter4));
  nand2 gate2106(.a(gate290inter4), .b(gate290inter3), .O(gate290inter5));
  nor2  gate2107(.a(gate290inter5), .b(gate290inter2), .O(gate290inter6));
  inv1  gate2108(.a(G820), .O(gate290inter7));
  inv1  gate2109(.a(G821), .O(gate290inter8));
  nand2 gate2110(.a(gate290inter8), .b(gate290inter7), .O(gate290inter9));
  nand2 gate2111(.a(s_223), .b(gate290inter3), .O(gate290inter10));
  nor2  gate2112(.a(gate290inter10), .b(gate290inter9), .O(gate290inter11));
  nor2  gate2113(.a(gate290inter11), .b(gate290inter6), .O(gate290inter12));
  nand2 gate2114(.a(gate290inter12), .b(gate290inter1), .O(G847));
nand2 gate291( .a(G822), .b(G823), .O(G860) );
nand2 gate292( .a(G824), .b(G825), .O(G873) );
nand2 gate293( .a(G828), .b(G829), .O(G886) );

  xor2  gate855(.a(G833), .b(G832), .O(gate294inter0));
  nand2 gate856(.a(gate294inter0), .b(s_44), .O(gate294inter1));
  and2  gate857(.a(G833), .b(G832), .O(gate294inter2));
  inv1  gate858(.a(s_44), .O(gate294inter3));
  inv1  gate859(.a(s_45), .O(gate294inter4));
  nand2 gate860(.a(gate294inter4), .b(gate294inter3), .O(gate294inter5));
  nor2  gate861(.a(gate294inter5), .b(gate294inter2), .O(gate294inter6));
  inv1  gate862(.a(G832), .O(gate294inter7));
  inv1  gate863(.a(G833), .O(gate294inter8));
  nand2 gate864(.a(gate294inter8), .b(gate294inter7), .O(gate294inter9));
  nand2 gate865(.a(s_45), .b(gate294inter3), .O(gate294inter10));
  nor2  gate866(.a(gate294inter10), .b(gate294inter9), .O(gate294inter11));
  nor2  gate867(.a(gate294inter11), .b(gate294inter6), .O(gate294inter12));
  nand2 gate868(.a(gate294inter12), .b(gate294inter1), .O(G899));

  xor2  gate2647(.a(G831), .b(G830), .O(gate295inter0));
  nand2 gate2648(.a(gate295inter0), .b(s_300), .O(gate295inter1));
  and2  gate2649(.a(G831), .b(G830), .O(gate295inter2));
  inv1  gate2650(.a(s_300), .O(gate295inter3));
  inv1  gate2651(.a(s_301), .O(gate295inter4));
  nand2 gate2652(.a(gate295inter4), .b(gate295inter3), .O(gate295inter5));
  nor2  gate2653(.a(gate295inter5), .b(gate295inter2), .O(gate295inter6));
  inv1  gate2654(.a(G830), .O(gate295inter7));
  inv1  gate2655(.a(G831), .O(gate295inter8));
  nand2 gate2656(.a(gate295inter8), .b(gate295inter7), .O(gate295inter9));
  nand2 gate2657(.a(s_301), .b(gate295inter3), .O(gate295inter10));
  nor2  gate2658(.a(gate295inter10), .b(gate295inter9), .O(gate295inter11));
  nor2  gate2659(.a(gate295inter11), .b(gate295inter6), .O(gate295inter12));
  nand2 gate2660(.a(gate295inter12), .b(gate295inter1), .O(G912));

  xor2  gate1331(.a(G827), .b(G826), .O(gate296inter0));
  nand2 gate1332(.a(gate296inter0), .b(s_112), .O(gate296inter1));
  and2  gate1333(.a(G827), .b(G826), .O(gate296inter2));
  inv1  gate1334(.a(s_112), .O(gate296inter3));
  inv1  gate1335(.a(s_113), .O(gate296inter4));
  nand2 gate1336(.a(gate296inter4), .b(gate296inter3), .O(gate296inter5));
  nor2  gate1337(.a(gate296inter5), .b(gate296inter2), .O(gate296inter6));
  inv1  gate1338(.a(G826), .O(gate296inter7));
  inv1  gate1339(.a(G827), .O(gate296inter8));
  nand2 gate1340(.a(gate296inter8), .b(gate296inter7), .O(gate296inter9));
  nand2 gate1341(.a(s_113), .b(gate296inter3), .O(gate296inter10));
  nor2  gate1342(.a(gate296inter10), .b(gate296inter9), .O(gate296inter11));
  nor2  gate1343(.a(gate296inter11), .b(gate296inter6), .O(gate296inter12));
  nand2 gate1344(.a(gate296inter12), .b(gate296inter1), .O(G925));
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );

  xor2  gate1513(.a(G1036), .b(G1), .O(gate387inter0));
  nand2 gate1514(.a(gate387inter0), .b(s_138), .O(gate387inter1));
  and2  gate1515(.a(G1036), .b(G1), .O(gate387inter2));
  inv1  gate1516(.a(s_138), .O(gate387inter3));
  inv1  gate1517(.a(s_139), .O(gate387inter4));
  nand2 gate1518(.a(gate387inter4), .b(gate387inter3), .O(gate387inter5));
  nor2  gate1519(.a(gate387inter5), .b(gate387inter2), .O(gate387inter6));
  inv1  gate1520(.a(G1), .O(gate387inter7));
  inv1  gate1521(.a(G1036), .O(gate387inter8));
  nand2 gate1522(.a(gate387inter8), .b(gate387inter7), .O(gate387inter9));
  nand2 gate1523(.a(s_139), .b(gate387inter3), .O(gate387inter10));
  nor2  gate1524(.a(gate387inter10), .b(gate387inter9), .O(gate387inter11));
  nor2  gate1525(.a(gate387inter11), .b(gate387inter6), .O(gate387inter12));
  nand2 gate1526(.a(gate387inter12), .b(gate387inter1), .O(G1132));
nand2 gate388( .a(G2), .b(G1039), .O(G1135) );

  xor2  gate2605(.a(G1042), .b(G3), .O(gate389inter0));
  nand2 gate2606(.a(gate389inter0), .b(s_294), .O(gate389inter1));
  and2  gate2607(.a(G1042), .b(G3), .O(gate389inter2));
  inv1  gate2608(.a(s_294), .O(gate389inter3));
  inv1  gate2609(.a(s_295), .O(gate389inter4));
  nand2 gate2610(.a(gate389inter4), .b(gate389inter3), .O(gate389inter5));
  nor2  gate2611(.a(gate389inter5), .b(gate389inter2), .O(gate389inter6));
  inv1  gate2612(.a(G3), .O(gate389inter7));
  inv1  gate2613(.a(G1042), .O(gate389inter8));
  nand2 gate2614(.a(gate389inter8), .b(gate389inter7), .O(gate389inter9));
  nand2 gate2615(.a(s_295), .b(gate389inter3), .O(gate389inter10));
  nor2  gate2616(.a(gate389inter10), .b(gate389inter9), .O(gate389inter11));
  nor2  gate2617(.a(gate389inter11), .b(gate389inter6), .O(gate389inter12));
  nand2 gate2618(.a(gate389inter12), .b(gate389inter1), .O(G1138));
nand2 gate390( .a(G4), .b(G1045), .O(G1141) );
nand2 gate391( .a(G5), .b(G1048), .O(G1144) );
nand2 gate392( .a(G6), .b(G1051), .O(G1147) );

  xor2  gate617(.a(G1054), .b(G7), .O(gate393inter0));
  nand2 gate618(.a(gate393inter0), .b(s_10), .O(gate393inter1));
  and2  gate619(.a(G1054), .b(G7), .O(gate393inter2));
  inv1  gate620(.a(s_10), .O(gate393inter3));
  inv1  gate621(.a(s_11), .O(gate393inter4));
  nand2 gate622(.a(gate393inter4), .b(gate393inter3), .O(gate393inter5));
  nor2  gate623(.a(gate393inter5), .b(gate393inter2), .O(gate393inter6));
  inv1  gate624(.a(G7), .O(gate393inter7));
  inv1  gate625(.a(G1054), .O(gate393inter8));
  nand2 gate626(.a(gate393inter8), .b(gate393inter7), .O(gate393inter9));
  nand2 gate627(.a(s_11), .b(gate393inter3), .O(gate393inter10));
  nor2  gate628(.a(gate393inter10), .b(gate393inter9), .O(gate393inter11));
  nor2  gate629(.a(gate393inter11), .b(gate393inter6), .O(gate393inter12));
  nand2 gate630(.a(gate393inter12), .b(gate393inter1), .O(G1150));
nand2 gate394( .a(G8), .b(G1057), .O(G1153) );
nand2 gate395( .a(G9), .b(G1060), .O(G1156) );

  xor2  gate1401(.a(G1063), .b(G10), .O(gate396inter0));
  nand2 gate1402(.a(gate396inter0), .b(s_122), .O(gate396inter1));
  and2  gate1403(.a(G1063), .b(G10), .O(gate396inter2));
  inv1  gate1404(.a(s_122), .O(gate396inter3));
  inv1  gate1405(.a(s_123), .O(gate396inter4));
  nand2 gate1406(.a(gate396inter4), .b(gate396inter3), .O(gate396inter5));
  nor2  gate1407(.a(gate396inter5), .b(gate396inter2), .O(gate396inter6));
  inv1  gate1408(.a(G10), .O(gate396inter7));
  inv1  gate1409(.a(G1063), .O(gate396inter8));
  nand2 gate1410(.a(gate396inter8), .b(gate396inter7), .O(gate396inter9));
  nand2 gate1411(.a(s_123), .b(gate396inter3), .O(gate396inter10));
  nor2  gate1412(.a(gate396inter10), .b(gate396inter9), .O(gate396inter11));
  nor2  gate1413(.a(gate396inter11), .b(gate396inter6), .O(gate396inter12));
  nand2 gate1414(.a(gate396inter12), .b(gate396inter1), .O(G1159));
nand2 gate397( .a(G11), .b(G1066), .O(G1162) );

  xor2  gate995(.a(G1069), .b(G12), .O(gate398inter0));
  nand2 gate996(.a(gate398inter0), .b(s_64), .O(gate398inter1));
  and2  gate997(.a(G1069), .b(G12), .O(gate398inter2));
  inv1  gate998(.a(s_64), .O(gate398inter3));
  inv1  gate999(.a(s_65), .O(gate398inter4));
  nand2 gate1000(.a(gate398inter4), .b(gate398inter3), .O(gate398inter5));
  nor2  gate1001(.a(gate398inter5), .b(gate398inter2), .O(gate398inter6));
  inv1  gate1002(.a(G12), .O(gate398inter7));
  inv1  gate1003(.a(G1069), .O(gate398inter8));
  nand2 gate1004(.a(gate398inter8), .b(gate398inter7), .O(gate398inter9));
  nand2 gate1005(.a(s_65), .b(gate398inter3), .O(gate398inter10));
  nor2  gate1006(.a(gate398inter10), .b(gate398inter9), .O(gate398inter11));
  nor2  gate1007(.a(gate398inter11), .b(gate398inter6), .O(gate398inter12));
  nand2 gate1008(.a(gate398inter12), .b(gate398inter1), .O(G1165));
nand2 gate399( .a(G13), .b(G1072), .O(G1168) );

  xor2  gate1219(.a(G1075), .b(G14), .O(gate400inter0));
  nand2 gate1220(.a(gate400inter0), .b(s_96), .O(gate400inter1));
  and2  gate1221(.a(G1075), .b(G14), .O(gate400inter2));
  inv1  gate1222(.a(s_96), .O(gate400inter3));
  inv1  gate1223(.a(s_97), .O(gate400inter4));
  nand2 gate1224(.a(gate400inter4), .b(gate400inter3), .O(gate400inter5));
  nor2  gate1225(.a(gate400inter5), .b(gate400inter2), .O(gate400inter6));
  inv1  gate1226(.a(G14), .O(gate400inter7));
  inv1  gate1227(.a(G1075), .O(gate400inter8));
  nand2 gate1228(.a(gate400inter8), .b(gate400inter7), .O(gate400inter9));
  nand2 gate1229(.a(s_97), .b(gate400inter3), .O(gate400inter10));
  nor2  gate1230(.a(gate400inter10), .b(gate400inter9), .O(gate400inter11));
  nor2  gate1231(.a(gate400inter11), .b(gate400inter6), .O(gate400inter12));
  nand2 gate1232(.a(gate400inter12), .b(gate400inter1), .O(G1171));

  xor2  gate981(.a(G1078), .b(G15), .O(gate401inter0));
  nand2 gate982(.a(gate401inter0), .b(s_62), .O(gate401inter1));
  and2  gate983(.a(G1078), .b(G15), .O(gate401inter2));
  inv1  gate984(.a(s_62), .O(gate401inter3));
  inv1  gate985(.a(s_63), .O(gate401inter4));
  nand2 gate986(.a(gate401inter4), .b(gate401inter3), .O(gate401inter5));
  nor2  gate987(.a(gate401inter5), .b(gate401inter2), .O(gate401inter6));
  inv1  gate988(.a(G15), .O(gate401inter7));
  inv1  gate989(.a(G1078), .O(gate401inter8));
  nand2 gate990(.a(gate401inter8), .b(gate401inter7), .O(gate401inter9));
  nand2 gate991(.a(s_63), .b(gate401inter3), .O(gate401inter10));
  nor2  gate992(.a(gate401inter10), .b(gate401inter9), .O(gate401inter11));
  nor2  gate993(.a(gate401inter11), .b(gate401inter6), .O(gate401inter12));
  nand2 gate994(.a(gate401inter12), .b(gate401inter1), .O(G1174));
nand2 gate402( .a(G16), .b(G1081), .O(G1177) );
nand2 gate403( .a(G17), .b(G1084), .O(G1180) );

  xor2  gate1107(.a(G1087), .b(G18), .O(gate404inter0));
  nand2 gate1108(.a(gate404inter0), .b(s_80), .O(gate404inter1));
  and2  gate1109(.a(G1087), .b(G18), .O(gate404inter2));
  inv1  gate1110(.a(s_80), .O(gate404inter3));
  inv1  gate1111(.a(s_81), .O(gate404inter4));
  nand2 gate1112(.a(gate404inter4), .b(gate404inter3), .O(gate404inter5));
  nor2  gate1113(.a(gate404inter5), .b(gate404inter2), .O(gate404inter6));
  inv1  gate1114(.a(G18), .O(gate404inter7));
  inv1  gate1115(.a(G1087), .O(gate404inter8));
  nand2 gate1116(.a(gate404inter8), .b(gate404inter7), .O(gate404inter9));
  nand2 gate1117(.a(s_81), .b(gate404inter3), .O(gate404inter10));
  nor2  gate1118(.a(gate404inter10), .b(gate404inter9), .O(gate404inter11));
  nor2  gate1119(.a(gate404inter11), .b(gate404inter6), .O(gate404inter12));
  nand2 gate1120(.a(gate404inter12), .b(gate404inter1), .O(G1183));
nand2 gate405( .a(G19), .b(G1090), .O(G1186) );
nand2 gate406( .a(G20), .b(G1093), .O(G1189) );

  xor2  gate1569(.a(G1096), .b(G21), .O(gate407inter0));
  nand2 gate1570(.a(gate407inter0), .b(s_146), .O(gate407inter1));
  and2  gate1571(.a(G1096), .b(G21), .O(gate407inter2));
  inv1  gate1572(.a(s_146), .O(gate407inter3));
  inv1  gate1573(.a(s_147), .O(gate407inter4));
  nand2 gate1574(.a(gate407inter4), .b(gate407inter3), .O(gate407inter5));
  nor2  gate1575(.a(gate407inter5), .b(gate407inter2), .O(gate407inter6));
  inv1  gate1576(.a(G21), .O(gate407inter7));
  inv1  gate1577(.a(G1096), .O(gate407inter8));
  nand2 gate1578(.a(gate407inter8), .b(gate407inter7), .O(gate407inter9));
  nand2 gate1579(.a(s_147), .b(gate407inter3), .O(gate407inter10));
  nor2  gate1580(.a(gate407inter10), .b(gate407inter9), .O(gate407inter11));
  nor2  gate1581(.a(gate407inter11), .b(gate407inter6), .O(gate407inter12));
  nand2 gate1582(.a(gate407inter12), .b(gate407inter1), .O(G1192));
nand2 gate408( .a(G22), .b(G1099), .O(G1195) );
nand2 gate409( .a(G23), .b(G1102), .O(G1198) );

  xor2  gate2115(.a(G1105), .b(G24), .O(gate410inter0));
  nand2 gate2116(.a(gate410inter0), .b(s_224), .O(gate410inter1));
  and2  gate2117(.a(G1105), .b(G24), .O(gate410inter2));
  inv1  gate2118(.a(s_224), .O(gate410inter3));
  inv1  gate2119(.a(s_225), .O(gate410inter4));
  nand2 gate2120(.a(gate410inter4), .b(gate410inter3), .O(gate410inter5));
  nor2  gate2121(.a(gate410inter5), .b(gate410inter2), .O(gate410inter6));
  inv1  gate2122(.a(G24), .O(gate410inter7));
  inv1  gate2123(.a(G1105), .O(gate410inter8));
  nand2 gate2124(.a(gate410inter8), .b(gate410inter7), .O(gate410inter9));
  nand2 gate2125(.a(s_225), .b(gate410inter3), .O(gate410inter10));
  nor2  gate2126(.a(gate410inter10), .b(gate410inter9), .O(gate410inter11));
  nor2  gate2127(.a(gate410inter11), .b(gate410inter6), .O(gate410inter12));
  nand2 gate2128(.a(gate410inter12), .b(gate410inter1), .O(G1201));
nand2 gate411( .a(G25), .b(G1108), .O(G1204) );
nand2 gate412( .a(G26), .b(G1111), .O(G1207) );

  xor2  gate1947(.a(G1114), .b(G27), .O(gate413inter0));
  nand2 gate1948(.a(gate413inter0), .b(s_200), .O(gate413inter1));
  and2  gate1949(.a(G1114), .b(G27), .O(gate413inter2));
  inv1  gate1950(.a(s_200), .O(gate413inter3));
  inv1  gate1951(.a(s_201), .O(gate413inter4));
  nand2 gate1952(.a(gate413inter4), .b(gate413inter3), .O(gate413inter5));
  nor2  gate1953(.a(gate413inter5), .b(gate413inter2), .O(gate413inter6));
  inv1  gate1954(.a(G27), .O(gate413inter7));
  inv1  gate1955(.a(G1114), .O(gate413inter8));
  nand2 gate1956(.a(gate413inter8), .b(gate413inter7), .O(gate413inter9));
  nand2 gate1957(.a(s_201), .b(gate413inter3), .O(gate413inter10));
  nor2  gate1958(.a(gate413inter10), .b(gate413inter9), .O(gate413inter11));
  nor2  gate1959(.a(gate413inter11), .b(gate413inter6), .O(gate413inter12));
  nand2 gate1960(.a(gate413inter12), .b(gate413inter1), .O(G1210));
nand2 gate414( .a(G28), .b(G1117), .O(G1213) );
nand2 gate415( .a(G29), .b(G1120), .O(G1216) );
nand2 gate416( .a(G30), .b(G1123), .O(G1219) );
nand2 gate417( .a(G31), .b(G1126), .O(G1222) );

  xor2  gate1009(.a(G1129), .b(G32), .O(gate418inter0));
  nand2 gate1010(.a(gate418inter0), .b(s_66), .O(gate418inter1));
  and2  gate1011(.a(G1129), .b(G32), .O(gate418inter2));
  inv1  gate1012(.a(s_66), .O(gate418inter3));
  inv1  gate1013(.a(s_67), .O(gate418inter4));
  nand2 gate1014(.a(gate418inter4), .b(gate418inter3), .O(gate418inter5));
  nor2  gate1015(.a(gate418inter5), .b(gate418inter2), .O(gate418inter6));
  inv1  gate1016(.a(G32), .O(gate418inter7));
  inv1  gate1017(.a(G1129), .O(gate418inter8));
  nand2 gate1018(.a(gate418inter8), .b(gate418inter7), .O(gate418inter9));
  nand2 gate1019(.a(s_67), .b(gate418inter3), .O(gate418inter10));
  nor2  gate1020(.a(gate418inter10), .b(gate418inter9), .O(gate418inter11));
  nor2  gate1021(.a(gate418inter11), .b(gate418inter6), .O(gate418inter12));
  nand2 gate1022(.a(gate418inter12), .b(gate418inter1), .O(G1225));
nand2 gate419( .a(G1), .b(G1132), .O(G1228) );
nand2 gate420( .a(G1036), .b(G1132), .O(G1229) );

  xor2  gate2255(.a(G1135), .b(G2), .O(gate421inter0));
  nand2 gate2256(.a(gate421inter0), .b(s_244), .O(gate421inter1));
  and2  gate2257(.a(G1135), .b(G2), .O(gate421inter2));
  inv1  gate2258(.a(s_244), .O(gate421inter3));
  inv1  gate2259(.a(s_245), .O(gate421inter4));
  nand2 gate2260(.a(gate421inter4), .b(gate421inter3), .O(gate421inter5));
  nor2  gate2261(.a(gate421inter5), .b(gate421inter2), .O(gate421inter6));
  inv1  gate2262(.a(G2), .O(gate421inter7));
  inv1  gate2263(.a(G1135), .O(gate421inter8));
  nand2 gate2264(.a(gate421inter8), .b(gate421inter7), .O(gate421inter9));
  nand2 gate2265(.a(s_245), .b(gate421inter3), .O(gate421inter10));
  nor2  gate2266(.a(gate421inter10), .b(gate421inter9), .O(gate421inter11));
  nor2  gate2267(.a(gate421inter11), .b(gate421inter6), .O(gate421inter12));
  nand2 gate2268(.a(gate421inter12), .b(gate421inter1), .O(G1230));
nand2 gate422( .a(G1039), .b(G1135), .O(G1231) );
nand2 gate423( .a(G3), .b(G1138), .O(G1232) );
nand2 gate424( .a(G1042), .b(G1138), .O(G1233) );
nand2 gate425( .a(G4), .b(G1141), .O(G1234) );

  xor2  gate701(.a(G1141), .b(G1045), .O(gate426inter0));
  nand2 gate702(.a(gate426inter0), .b(s_22), .O(gate426inter1));
  and2  gate703(.a(G1141), .b(G1045), .O(gate426inter2));
  inv1  gate704(.a(s_22), .O(gate426inter3));
  inv1  gate705(.a(s_23), .O(gate426inter4));
  nand2 gate706(.a(gate426inter4), .b(gate426inter3), .O(gate426inter5));
  nor2  gate707(.a(gate426inter5), .b(gate426inter2), .O(gate426inter6));
  inv1  gate708(.a(G1045), .O(gate426inter7));
  inv1  gate709(.a(G1141), .O(gate426inter8));
  nand2 gate710(.a(gate426inter8), .b(gate426inter7), .O(gate426inter9));
  nand2 gate711(.a(s_23), .b(gate426inter3), .O(gate426inter10));
  nor2  gate712(.a(gate426inter10), .b(gate426inter9), .O(gate426inter11));
  nor2  gate713(.a(gate426inter11), .b(gate426inter6), .O(gate426inter12));
  nand2 gate714(.a(gate426inter12), .b(gate426inter1), .O(G1235));
nand2 gate427( .a(G5), .b(G1144), .O(G1236) );
nand2 gate428( .a(G1048), .b(G1144), .O(G1237) );

  xor2  gate1583(.a(G1147), .b(G6), .O(gate429inter0));
  nand2 gate1584(.a(gate429inter0), .b(s_148), .O(gate429inter1));
  and2  gate1585(.a(G1147), .b(G6), .O(gate429inter2));
  inv1  gate1586(.a(s_148), .O(gate429inter3));
  inv1  gate1587(.a(s_149), .O(gate429inter4));
  nand2 gate1588(.a(gate429inter4), .b(gate429inter3), .O(gate429inter5));
  nor2  gate1589(.a(gate429inter5), .b(gate429inter2), .O(gate429inter6));
  inv1  gate1590(.a(G6), .O(gate429inter7));
  inv1  gate1591(.a(G1147), .O(gate429inter8));
  nand2 gate1592(.a(gate429inter8), .b(gate429inter7), .O(gate429inter9));
  nand2 gate1593(.a(s_149), .b(gate429inter3), .O(gate429inter10));
  nor2  gate1594(.a(gate429inter10), .b(gate429inter9), .O(gate429inter11));
  nor2  gate1595(.a(gate429inter11), .b(gate429inter6), .O(gate429inter12));
  nand2 gate1596(.a(gate429inter12), .b(gate429inter1), .O(G1238));
nand2 gate430( .a(G1051), .b(G1147), .O(G1239) );
nand2 gate431( .a(G7), .b(G1150), .O(G1240) );
nand2 gate432( .a(G1054), .b(G1150), .O(G1241) );
nand2 gate433( .a(G8), .b(G1153), .O(G1242) );
nand2 gate434( .a(G1057), .b(G1153), .O(G1243) );

  xor2  gate547(.a(G1156), .b(G9), .O(gate435inter0));
  nand2 gate548(.a(gate435inter0), .b(s_0), .O(gate435inter1));
  and2  gate549(.a(G1156), .b(G9), .O(gate435inter2));
  inv1  gate550(.a(s_0), .O(gate435inter3));
  inv1  gate551(.a(s_1), .O(gate435inter4));
  nand2 gate552(.a(gate435inter4), .b(gate435inter3), .O(gate435inter5));
  nor2  gate553(.a(gate435inter5), .b(gate435inter2), .O(gate435inter6));
  inv1  gate554(.a(G9), .O(gate435inter7));
  inv1  gate555(.a(G1156), .O(gate435inter8));
  nand2 gate556(.a(gate435inter8), .b(gate435inter7), .O(gate435inter9));
  nand2 gate557(.a(s_1), .b(gate435inter3), .O(gate435inter10));
  nor2  gate558(.a(gate435inter10), .b(gate435inter9), .O(gate435inter11));
  nor2  gate559(.a(gate435inter11), .b(gate435inter6), .O(gate435inter12));
  nand2 gate560(.a(gate435inter12), .b(gate435inter1), .O(G1244));
nand2 gate436( .a(G1060), .b(G1156), .O(G1245) );

  xor2  gate1065(.a(G1159), .b(G10), .O(gate437inter0));
  nand2 gate1066(.a(gate437inter0), .b(s_74), .O(gate437inter1));
  and2  gate1067(.a(G1159), .b(G10), .O(gate437inter2));
  inv1  gate1068(.a(s_74), .O(gate437inter3));
  inv1  gate1069(.a(s_75), .O(gate437inter4));
  nand2 gate1070(.a(gate437inter4), .b(gate437inter3), .O(gate437inter5));
  nor2  gate1071(.a(gate437inter5), .b(gate437inter2), .O(gate437inter6));
  inv1  gate1072(.a(G10), .O(gate437inter7));
  inv1  gate1073(.a(G1159), .O(gate437inter8));
  nand2 gate1074(.a(gate437inter8), .b(gate437inter7), .O(gate437inter9));
  nand2 gate1075(.a(s_75), .b(gate437inter3), .O(gate437inter10));
  nor2  gate1076(.a(gate437inter10), .b(gate437inter9), .O(gate437inter11));
  nor2  gate1077(.a(gate437inter11), .b(gate437inter6), .O(gate437inter12));
  nand2 gate1078(.a(gate437inter12), .b(gate437inter1), .O(G1246));
nand2 gate438( .a(G1063), .b(G1159), .O(G1247) );
nand2 gate439( .a(G11), .b(G1162), .O(G1248) );
nand2 gate440( .a(G1066), .b(G1162), .O(G1249) );

  xor2  gate2731(.a(G1165), .b(G12), .O(gate441inter0));
  nand2 gate2732(.a(gate441inter0), .b(s_312), .O(gate441inter1));
  and2  gate2733(.a(G1165), .b(G12), .O(gate441inter2));
  inv1  gate2734(.a(s_312), .O(gate441inter3));
  inv1  gate2735(.a(s_313), .O(gate441inter4));
  nand2 gate2736(.a(gate441inter4), .b(gate441inter3), .O(gate441inter5));
  nor2  gate2737(.a(gate441inter5), .b(gate441inter2), .O(gate441inter6));
  inv1  gate2738(.a(G12), .O(gate441inter7));
  inv1  gate2739(.a(G1165), .O(gate441inter8));
  nand2 gate2740(.a(gate441inter8), .b(gate441inter7), .O(gate441inter9));
  nand2 gate2741(.a(s_313), .b(gate441inter3), .O(gate441inter10));
  nor2  gate2742(.a(gate441inter10), .b(gate441inter9), .O(gate441inter11));
  nor2  gate2743(.a(gate441inter11), .b(gate441inter6), .O(gate441inter12));
  nand2 gate2744(.a(gate441inter12), .b(gate441inter1), .O(G1250));
nand2 gate442( .a(G1069), .b(G1165), .O(G1251) );
nand2 gate443( .a(G13), .b(G1168), .O(G1252) );
nand2 gate444( .a(G1072), .b(G1168), .O(G1253) );
nand2 gate445( .a(G14), .b(G1171), .O(G1254) );
nand2 gate446( .a(G1075), .b(G1171), .O(G1255) );
nand2 gate447( .a(G15), .b(G1174), .O(G1256) );

  xor2  gate1723(.a(G1174), .b(G1078), .O(gate448inter0));
  nand2 gate1724(.a(gate448inter0), .b(s_168), .O(gate448inter1));
  and2  gate1725(.a(G1174), .b(G1078), .O(gate448inter2));
  inv1  gate1726(.a(s_168), .O(gate448inter3));
  inv1  gate1727(.a(s_169), .O(gate448inter4));
  nand2 gate1728(.a(gate448inter4), .b(gate448inter3), .O(gate448inter5));
  nor2  gate1729(.a(gate448inter5), .b(gate448inter2), .O(gate448inter6));
  inv1  gate1730(.a(G1078), .O(gate448inter7));
  inv1  gate1731(.a(G1174), .O(gate448inter8));
  nand2 gate1732(.a(gate448inter8), .b(gate448inter7), .O(gate448inter9));
  nand2 gate1733(.a(s_169), .b(gate448inter3), .O(gate448inter10));
  nor2  gate1734(.a(gate448inter10), .b(gate448inter9), .O(gate448inter11));
  nor2  gate1735(.a(gate448inter11), .b(gate448inter6), .O(gate448inter12));
  nand2 gate1736(.a(gate448inter12), .b(gate448inter1), .O(G1257));

  xor2  gate1429(.a(G1177), .b(G16), .O(gate449inter0));
  nand2 gate1430(.a(gate449inter0), .b(s_126), .O(gate449inter1));
  and2  gate1431(.a(G1177), .b(G16), .O(gate449inter2));
  inv1  gate1432(.a(s_126), .O(gate449inter3));
  inv1  gate1433(.a(s_127), .O(gate449inter4));
  nand2 gate1434(.a(gate449inter4), .b(gate449inter3), .O(gate449inter5));
  nor2  gate1435(.a(gate449inter5), .b(gate449inter2), .O(gate449inter6));
  inv1  gate1436(.a(G16), .O(gate449inter7));
  inv1  gate1437(.a(G1177), .O(gate449inter8));
  nand2 gate1438(.a(gate449inter8), .b(gate449inter7), .O(gate449inter9));
  nand2 gate1439(.a(s_127), .b(gate449inter3), .O(gate449inter10));
  nor2  gate1440(.a(gate449inter10), .b(gate449inter9), .O(gate449inter11));
  nor2  gate1441(.a(gate449inter11), .b(gate449inter6), .O(gate449inter12));
  nand2 gate1442(.a(gate449inter12), .b(gate449inter1), .O(G1258));

  xor2  gate561(.a(G1177), .b(G1081), .O(gate450inter0));
  nand2 gate562(.a(gate450inter0), .b(s_2), .O(gate450inter1));
  and2  gate563(.a(G1177), .b(G1081), .O(gate450inter2));
  inv1  gate564(.a(s_2), .O(gate450inter3));
  inv1  gate565(.a(s_3), .O(gate450inter4));
  nand2 gate566(.a(gate450inter4), .b(gate450inter3), .O(gate450inter5));
  nor2  gate567(.a(gate450inter5), .b(gate450inter2), .O(gate450inter6));
  inv1  gate568(.a(G1081), .O(gate450inter7));
  inv1  gate569(.a(G1177), .O(gate450inter8));
  nand2 gate570(.a(gate450inter8), .b(gate450inter7), .O(gate450inter9));
  nand2 gate571(.a(s_3), .b(gate450inter3), .O(gate450inter10));
  nor2  gate572(.a(gate450inter10), .b(gate450inter9), .O(gate450inter11));
  nor2  gate573(.a(gate450inter11), .b(gate450inter6), .O(gate450inter12));
  nand2 gate574(.a(gate450inter12), .b(gate450inter1), .O(G1259));

  xor2  gate2773(.a(G1180), .b(G17), .O(gate451inter0));
  nand2 gate2774(.a(gate451inter0), .b(s_318), .O(gate451inter1));
  and2  gate2775(.a(G1180), .b(G17), .O(gate451inter2));
  inv1  gate2776(.a(s_318), .O(gate451inter3));
  inv1  gate2777(.a(s_319), .O(gate451inter4));
  nand2 gate2778(.a(gate451inter4), .b(gate451inter3), .O(gate451inter5));
  nor2  gate2779(.a(gate451inter5), .b(gate451inter2), .O(gate451inter6));
  inv1  gate2780(.a(G17), .O(gate451inter7));
  inv1  gate2781(.a(G1180), .O(gate451inter8));
  nand2 gate2782(.a(gate451inter8), .b(gate451inter7), .O(gate451inter9));
  nand2 gate2783(.a(s_319), .b(gate451inter3), .O(gate451inter10));
  nor2  gate2784(.a(gate451inter10), .b(gate451inter9), .O(gate451inter11));
  nor2  gate2785(.a(gate451inter11), .b(gate451inter6), .O(gate451inter12));
  nand2 gate2786(.a(gate451inter12), .b(gate451inter1), .O(G1260));
nand2 gate452( .a(G1084), .b(G1180), .O(G1261) );

  xor2  gate2409(.a(G1183), .b(G18), .O(gate453inter0));
  nand2 gate2410(.a(gate453inter0), .b(s_266), .O(gate453inter1));
  and2  gate2411(.a(G1183), .b(G18), .O(gate453inter2));
  inv1  gate2412(.a(s_266), .O(gate453inter3));
  inv1  gate2413(.a(s_267), .O(gate453inter4));
  nand2 gate2414(.a(gate453inter4), .b(gate453inter3), .O(gate453inter5));
  nor2  gate2415(.a(gate453inter5), .b(gate453inter2), .O(gate453inter6));
  inv1  gate2416(.a(G18), .O(gate453inter7));
  inv1  gate2417(.a(G1183), .O(gate453inter8));
  nand2 gate2418(.a(gate453inter8), .b(gate453inter7), .O(gate453inter9));
  nand2 gate2419(.a(s_267), .b(gate453inter3), .O(gate453inter10));
  nor2  gate2420(.a(gate453inter10), .b(gate453inter9), .O(gate453inter11));
  nor2  gate2421(.a(gate453inter11), .b(gate453inter6), .O(gate453inter12));
  nand2 gate2422(.a(gate453inter12), .b(gate453inter1), .O(G1262));
nand2 gate454( .a(G1087), .b(G1183), .O(G1263) );
nand2 gate455( .a(G19), .b(G1186), .O(G1264) );
nand2 gate456( .a(G1090), .b(G1186), .O(G1265) );
nand2 gate457( .a(G20), .b(G1189), .O(G1266) );
nand2 gate458( .a(G1093), .b(G1189), .O(G1267) );
nand2 gate459( .a(G21), .b(G1192), .O(G1268) );

  xor2  gate2787(.a(G1192), .b(G1096), .O(gate460inter0));
  nand2 gate2788(.a(gate460inter0), .b(s_320), .O(gate460inter1));
  and2  gate2789(.a(G1192), .b(G1096), .O(gate460inter2));
  inv1  gate2790(.a(s_320), .O(gate460inter3));
  inv1  gate2791(.a(s_321), .O(gate460inter4));
  nand2 gate2792(.a(gate460inter4), .b(gate460inter3), .O(gate460inter5));
  nor2  gate2793(.a(gate460inter5), .b(gate460inter2), .O(gate460inter6));
  inv1  gate2794(.a(G1096), .O(gate460inter7));
  inv1  gate2795(.a(G1192), .O(gate460inter8));
  nand2 gate2796(.a(gate460inter8), .b(gate460inter7), .O(gate460inter9));
  nand2 gate2797(.a(s_321), .b(gate460inter3), .O(gate460inter10));
  nor2  gate2798(.a(gate460inter10), .b(gate460inter9), .O(gate460inter11));
  nor2  gate2799(.a(gate460inter11), .b(gate460inter6), .O(gate460inter12));
  nand2 gate2800(.a(gate460inter12), .b(gate460inter1), .O(G1269));
nand2 gate461( .a(G22), .b(G1195), .O(G1270) );
nand2 gate462( .a(G1099), .b(G1195), .O(G1271) );
nand2 gate463( .a(G23), .b(G1198), .O(G1272) );

  xor2  gate2199(.a(G1198), .b(G1102), .O(gate464inter0));
  nand2 gate2200(.a(gate464inter0), .b(s_236), .O(gate464inter1));
  and2  gate2201(.a(G1198), .b(G1102), .O(gate464inter2));
  inv1  gate2202(.a(s_236), .O(gate464inter3));
  inv1  gate2203(.a(s_237), .O(gate464inter4));
  nand2 gate2204(.a(gate464inter4), .b(gate464inter3), .O(gate464inter5));
  nor2  gate2205(.a(gate464inter5), .b(gate464inter2), .O(gate464inter6));
  inv1  gate2206(.a(G1102), .O(gate464inter7));
  inv1  gate2207(.a(G1198), .O(gate464inter8));
  nand2 gate2208(.a(gate464inter8), .b(gate464inter7), .O(gate464inter9));
  nand2 gate2209(.a(s_237), .b(gate464inter3), .O(gate464inter10));
  nor2  gate2210(.a(gate464inter10), .b(gate464inter9), .O(gate464inter11));
  nor2  gate2211(.a(gate464inter11), .b(gate464inter6), .O(gate464inter12));
  nand2 gate2212(.a(gate464inter12), .b(gate464inter1), .O(G1273));

  xor2  gate2059(.a(G1201), .b(G24), .O(gate465inter0));
  nand2 gate2060(.a(gate465inter0), .b(s_216), .O(gate465inter1));
  and2  gate2061(.a(G1201), .b(G24), .O(gate465inter2));
  inv1  gate2062(.a(s_216), .O(gate465inter3));
  inv1  gate2063(.a(s_217), .O(gate465inter4));
  nand2 gate2064(.a(gate465inter4), .b(gate465inter3), .O(gate465inter5));
  nor2  gate2065(.a(gate465inter5), .b(gate465inter2), .O(gate465inter6));
  inv1  gate2066(.a(G24), .O(gate465inter7));
  inv1  gate2067(.a(G1201), .O(gate465inter8));
  nand2 gate2068(.a(gate465inter8), .b(gate465inter7), .O(gate465inter9));
  nand2 gate2069(.a(s_217), .b(gate465inter3), .O(gate465inter10));
  nor2  gate2070(.a(gate465inter10), .b(gate465inter9), .O(gate465inter11));
  nor2  gate2071(.a(gate465inter11), .b(gate465inter6), .O(gate465inter12));
  nand2 gate2072(.a(gate465inter12), .b(gate465inter1), .O(G1274));
nand2 gate466( .a(G1105), .b(G1201), .O(G1275) );

  xor2  gate2521(.a(G1204), .b(G25), .O(gate467inter0));
  nand2 gate2522(.a(gate467inter0), .b(s_282), .O(gate467inter1));
  and2  gate2523(.a(G1204), .b(G25), .O(gate467inter2));
  inv1  gate2524(.a(s_282), .O(gate467inter3));
  inv1  gate2525(.a(s_283), .O(gate467inter4));
  nand2 gate2526(.a(gate467inter4), .b(gate467inter3), .O(gate467inter5));
  nor2  gate2527(.a(gate467inter5), .b(gate467inter2), .O(gate467inter6));
  inv1  gate2528(.a(G25), .O(gate467inter7));
  inv1  gate2529(.a(G1204), .O(gate467inter8));
  nand2 gate2530(.a(gate467inter8), .b(gate467inter7), .O(gate467inter9));
  nand2 gate2531(.a(s_283), .b(gate467inter3), .O(gate467inter10));
  nor2  gate2532(.a(gate467inter10), .b(gate467inter9), .O(gate467inter11));
  nor2  gate2533(.a(gate467inter11), .b(gate467inter6), .O(gate467inter12));
  nand2 gate2534(.a(gate467inter12), .b(gate467inter1), .O(G1276));
nand2 gate468( .a(G1108), .b(G1204), .O(G1277) );
nand2 gate469( .a(G26), .b(G1207), .O(G1278) );
nand2 gate470( .a(G1111), .b(G1207), .O(G1279) );

  xor2  gate1499(.a(G1210), .b(G27), .O(gate471inter0));
  nand2 gate1500(.a(gate471inter0), .b(s_136), .O(gate471inter1));
  and2  gate1501(.a(G1210), .b(G27), .O(gate471inter2));
  inv1  gate1502(.a(s_136), .O(gate471inter3));
  inv1  gate1503(.a(s_137), .O(gate471inter4));
  nand2 gate1504(.a(gate471inter4), .b(gate471inter3), .O(gate471inter5));
  nor2  gate1505(.a(gate471inter5), .b(gate471inter2), .O(gate471inter6));
  inv1  gate1506(.a(G27), .O(gate471inter7));
  inv1  gate1507(.a(G1210), .O(gate471inter8));
  nand2 gate1508(.a(gate471inter8), .b(gate471inter7), .O(gate471inter9));
  nand2 gate1509(.a(s_137), .b(gate471inter3), .O(gate471inter10));
  nor2  gate1510(.a(gate471inter10), .b(gate471inter9), .O(gate471inter11));
  nor2  gate1511(.a(gate471inter11), .b(gate471inter6), .O(gate471inter12));
  nand2 gate1512(.a(gate471inter12), .b(gate471inter1), .O(G1280));
nand2 gate472( .a(G1114), .b(G1210), .O(G1281) );
nand2 gate473( .a(G28), .b(G1213), .O(G1282) );

  xor2  gate1807(.a(G1213), .b(G1117), .O(gate474inter0));
  nand2 gate1808(.a(gate474inter0), .b(s_180), .O(gate474inter1));
  and2  gate1809(.a(G1213), .b(G1117), .O(gate474inter2));
  inv1  gate1810(.a(s_180), .O(gate474inter3));
  inv1  gate1811(.a(s_181), .O(gate474inter4));
  nand2 gate1812(.a(gate474inter4), .b(gate474inter3), .O(gate474inter5));
  nor2  gate1813(.a(gate474inter5), .b(gate474inter2), .O(gate474inter6));
  inv1  gate1814(.a(G1117), .O(gate474inter7));
  inv1  gate1815(.a(G1213), .O(gate474inter8));
  nand2 gate1816(.a(gate474inter8), .b(gate474inter7), .O(gate474inter9));
  nand2 gate1817(.a(s_181), .b(gate474inter3), .O(gate474inter10));
  nor2  gate1818(.a(gate474inter10), .b(gate474inter9), .O(gate474inter11));
  nor2  gate1819(.a(gate474inter11), .b(gate474inter6), .O(gate474inter12));
  nand2 gate1820(.a(gate474inter12), .b(gate474inter1), .O(G1283));
nand2 gate475( .a(G29), .b(G1216), .O(G1284) );
nand2 gate476( .a(G1120), .b(G1216), .O(G1285) );
nand2 gate477( .a(G30), .b(G1219), .O(G1286) );

  xor2  gate2633(.a(G1219), .b(G1123), .O(gate478inter0));
  nand2 gate2634(.a(gate478inter0), .b(s_298), .O(gate478inter1));
  and2  gate2635(.a(G1219), .b(G1123), .O(gate478inter2));
  inv1  gate2636(.a(s_298), .O(gate478inter3));
  inv1  gate2637(.a(s_299), .O(gate478inter4));
  nand2 gate2638(.a(gate478inter4), .b(gate478inter3), .O(gate478inter5));
  nor2  gate2639(.a(gate478inter5), .b(gate478inter2), .O(gate478inter6));
  inv1  gate2640(.a(G1123), .O(gate478inter7));
  inv1  gate2641(.a(G1219), .O(gate478inter8));
  nand2 gate2642(.a(gate478inter8), .b(gate478inter7), .O(gate478inter9));
  nand2 gate2643(.a(s_299), .b(gate478inter3), .O(gate478inter10));
  nor2  gate2644(.a(gate478inter10), .b(gate478inter9), .O(gate478inter11));
  nor2  gate2645(.a(gate478inter11), .b(gate478inter6), .O(gate478inter12));
  nand2 gate2646(.a(gate478inter12), .b(gate478inter1), .O(G1287));

  xor2  gate1149(.a(G1222), .b(G31), .O(gate479inter0));
  nand2 gate1150(.a(gate479inter0), .b(s_86), .O(gate479inter1));
  and2  gate1151(.a(G1222), .b(G31), .O(gate479inter2));
  inv1  gate1152(.a(s_86), .O(gate479inter3));
  inv1  gate1153(.a(s_87), .O(gate479inter4));
  nand2 gate1154(.a(gate479inter4), .b(gate479inter3), .O(gate479inter5));
  nor2  gate1155(.a(gate479inter5), .b(gate479inter2), .O(gate479inter6));
  inv1  gate1156(.a(G31), .O(gate479inter7));
  inv1  gate1157(.a(G1222), .O(gate479inter8));
  nand2 gate1158(.a(gate479inter8), .b(gate479inter7), .O(gate479inter9));
  nand2 gate1159(.a(s_87), .b(gate479inter3), .O(gate479inter10));
  nor2  gate1160(.a(gate479inter10), .b(gate479inter9), .O(gate479inter11));
  nor2  gate1161(.a(gate479inter11), .b(gate479inter6), .O(gate479inter12));
  nand2 gate1162(.a(gate479inter12), .b(gate479inter1), .O(G1288));
nand2 gate480( .a(G1126), .b(G1222), .O(G1289) );
nand2 gate481( .a(G32), .b(G1225), .O(G1290) );
nand2 gate482( .a(G1129), .b(G1225), .O(G1291) );

  xor2  gate1779(.a(G1229), .b(G1228), .O(gate483inter0));
  nand2 gate1780(.a(gate483inter0), .b(s_176), .O(gate483inter1));
  and2  gate1781(.a(G1229), .b(G1228), .O(gate483inter2));
  inv1  gate1782(.a(s_176), .O(gate483inter3));
  inv1  gate1783(.a(s_177), .O(gate483inter4));
  nand2 gate1784(.a(gate483inter4), .b(gate483inter3), .O(gate483inter5));
  nor2  gate1785(.a(gate483inter5), .b(gate483inter2), .O(gate483inter6));
  inv1  gate1786(.a(G1228), .O(gate483inter7));
  inv1  gate1787(.a(G1229), .O(gate483inter8));
  nand2 gate1788(.a(gate483inter8), .b(gate483inter7), .O(gate483inter9));
  nand2 gate1789(.a(s_177), .b(gate483inter3), .O(gate483inter10));
  nor2  gate1790(.a(gate483inter10), .b(gate483inter9), .O(gate483inter11));
  nor2  gate1791(.a(gate483inter11), .b(gate483inter6), .O(gate483inter12));
  nand2 gate1792(.a(gate483inter12), .b(gate483inter1), .O(G1292));

  xor2  gate2689(.a(G1231), .b(G1230), .O(gate484inter0));
  nand2 gate2690(.a(gate484inter0), .b(s_306), .O(gate484inter1));
  and2  gate2691(.a(G1231), .b(G1230), .O(gate484inter2));
  inv1  gate2692(.a(s_306), .O(gate484inter3));
  inv1  gate2693(.a(s_307), .O(gate484inter4));
  nand2 gate2694(.a(gate484inter4), .b(gate484inter3), .O(gate484inter5));
  nor2  gate2695(.a(gate484inter5), .b(gate484inter2), .O(gate484inter6));
  inv1  gate2696(.a(G1230), .O(gate484inter7));
  inv1  gate2697(.a(G1231), .O(gate484inter8));
  nand2 gate2698(.a(gate484inter8), .b(gate484inter7), .O(gate484inter9));
  nand2 gate2699(.a(s_307), .b(gate484inter3), .O(gate484inter10));
  nor2  gate2700(.a(gate484inter10), .b(gate484inter9), .O(gate484inter11));
  nor2  gate2701(.a(gate484inter11), .b(gate484inter6), .O(gate484inter12));
  nand2 gate2702(.a(gate484inter12), .b(gate484inter1), .O(G1293));
nand2 gate485( .a(G1232), .b(G1233), .O(G1294) );

  xor2  gate953(.a(G1235), .b(G1234), .O(gate486inter0));
  nand2 gate954(.a(gate486inter0), .b(s_58), .O(gate486inter1));
  and2  gate955(.a(G1235), .b(G1234), .O(gate486inter2));
  inv1  gate956(.a(s_58), .O(gate486inter3));
  inv1  gate957(.a(s_59), .O(gate486inter4));
  nand2 gate958(.a(gate486inter4), .b(gate486inter3), .O(gate486inter5));
  nor2  gate959(.a(gate486inter5), .b(gate486inter2), .O(gate486inter6));
  inv1  gate960(.a(G1234), .O(gate486inter7));
  inv1  gate961(.a(G1235), .O(gate486inter8));
  nand2 gate962(.a(gate486inter8), .b(gate486inter7), .O(gate486inter9));
  nand2 gate963(.a(s_59), .b(gate486inter3), .O(gate486inter10));
  nor2  gate964(.a(gate486inter10), .b(gate486inter9), .O(gate486inter11));
  nor2  gate965(.a(gate486inter11), .b(gate486inter6), .O(gate486inter12));
  nand2 gate966(.a(gate486inter12), .b(gate486inter1), .O(G1295));
nand2 gate487( .a(G1236), .b(G1237), .O(G1296) );

  xor2  gate1905(.a(G1239), .b(G1238), .O(gate488inter0));
  nand2 gate1906(.a(gate488inter0), .b(s_194), .O(gate488inter1));
  and2  gate1907(.a(G1239), .b(G1238), .O(gate488inter2));
  inv1  gate1908(.a(s_194), .O(gate488inter3));
  inv1  gate1909(.a(s_195), .O(gate488inter4));
  nand2 gate1910(.a(gate488inter4), .b(gate488inter3), .O(gate488inter5));
  nor2  gate1911(.a(gate488inter5), .b(gate488inter2), .O(gate488inter6));
  inv1  gate1912(.a(G1238), .O(gate488inter7));
  inv1  gate1913(.a(G1239), .O(gate488inter8));
  nand2 gate1914(.a(gate488inter8), .b(gate488inter7), .O(gate488inter9));
  nand2 gate1915(.a(s_195), .b(gate488inter3), .O(gate488inter10));
  nor2  gate1916(.a(gate488inter10), .b(gate488inter9), .O(gate488inter11));
  nor2  gate1917(.a(gate488inter11), .b(gate488inter6), .O(gate488inter12));
  nand2 gate1918(.a(gate488inter12), .b(gate488inter1), .O(G1297));
nand2 gate489( .a(G1240), .b(G1241), .O(G1298) );

  xor2  gate1751(.a(G1243), .b(G1242), .O(gate490inter0));
  nand2 gate1752(.a(gate490inter0), .b(s_172), .O(gate490inter1));
  and2  gate1753(.a(G1243), .b(G1242), .O(gate490inter2));
  inv1  gate1754(.a(s_172), .O(gate490inter3));
  inv1  gate1755(.a(s_173), .O(gate490inter4));
  nand2 gate1756(.a(gate490inter4), .b(gate490inter3), .O(gate490inter5));
  nor2  gate1757(.a(gate490inter5), .b(gate490inter2), .O(gate490inter6));
  inv1  gate1758(.a(G1242), .O(gate490inter7));
  inv1  gate1759(.a(G1243), .O(gate490inter8));
  nand2 gate1760(.a(gate490inter8), .b(gate490inter7), .O(gate490inter9));
  nand2 gate1761(.a(s_173), .b(gate490inter3), .O(gate490inter10));
  nor2  gate1762(.a(gate490inter10), .b(gate490inter9), .O(gate490inter11));
  nor2  gate1763(.a(gate490inter11), .b(gate490inter6), .O(gate490inter12));
  nand2 gate1764(.a(gate490inter12), .b(gate490inter1), .O(G1299));
nand2 gate491( .a(G1244), .b(G1245), .O(G1300) );
nand2 gate492( .a(G1246), .b(G1247), .O(G1301) );
nand2 gate493( .a(G1248), .b(G1249), .O(G1302) );
nand2 gate494( .a(G1250), .b(G1251), .O(G1303) );

  xor2  gate1541(.a(G1253), .b(G1252), .O(gate495inter0));
  nand2 gate1542(.a(gate495inter0), .b(s_142), .O(gate495inter1));
  and2  gate1543(.a(G1253), .b(G1252), .O(gate495inter2));
  inv1  gate1544(.a(s_142), .O(gate495inter3));
  inv1  gate1545(.a(s_143), .O(gate495inter4));
  nand2 gate1546(.a(gate495inter4), .b(gate495inter3), .O(gate495inter5));
  nor2  gate1547(.a(gate495inter5), .b(gate495inter2), .O(gate495inter6));
  inv1  gate1548(.a(G1252), .O(gate495inter7));
  inv1  gate1549(.a(G1253), .O(gate495inter8));
  nand2 gate1550(.a(gate495inter8), .b(gate495inter7), .O(gate495inter9));
  nand2 gate1551(.a(s_143), .b(gate495inter3), .O(gate495inter10));
  nor2  gate1552(.a(gate495inter10), .b(gate495inter9), .O(gate495inter11));
  nor2  gate1553(.a(gate495inter11), .b(gate495inter6), .O(gate495inter12));
  nand2 gate1554(.a(gate495inter12), .b(gate495inter1), .O(G1304));

  xor2  gate1289(.a(G1255), .b(G1254), .O(gate496inter0));
  nand2 gate1290(.a(gate496inter0), .b(s_106), .O(gate496inter1));
  and2  gate1291(.a(G1255), .b(G1254), .O(gate496inter2));
  inv1  gate1292(.a(s_106), .O(gate496inter3));
  inv1  gate1293(.a(s_107), .O(gate496inter4));
  nand2 gate1294(.a(gate496inter4), .b(gate496inter3), .O(gate496inter5));
  nor2  gate1295(.a(gate496inter5), .b(gate496inter2), .O(gate496inter6));
  inv1  gate1296(.a(G1254), .O(gate496inter7));
  inv1  gate1297(.a(G1255), .O(gate496inter8));
  nand2 gate1298(.a(gate496inter8), .b(gate496inter7), .O(gate496inter9));
  nand2 gate1299(.a(s_107), .b(gate496inter3), .O(gate496inter10));
  nor2  gate1300(.a(gate496inter10), .b(gate496inter9), .O(gate496inter11));
  nor2  gate1301(.a(gate496inter11), .b(gate496inter6), .O(gate496inter12));
  nand2 gate1302(.a(gate496inter12), .b(gate496inter1), .O(G1305));
nand2 gate497( .a(G1256), .b(G1257), .O(G1306) );

  xor2  gate1247(.a(G1259), .b(G1258), .O(gate498inter0));
  nand2 gate1248(.a(gate498inter0), .b(s_100), .O(gate498inter1));
  and2  gate1249(.a(G1259), .b(G1258), .O(gate498inter2));
  inv1  gate1250(.a(s_100), .O(gate498inter3));
  inv1  gate1251(.a(s_101), .O(gate498inter4));
  nand2 gate1252(.a(gate498inter4), .b(gate498inter3), .O(gate498inter5));
  nor2  gate1253(.a(gate498inter5), .b(gate498inter2), .O(gate498inter6));
  inv1  gate1254(.a(G1258), .O(gate498inter7));
  inv1  gate1255(.a(G1259), .O(gate498inter8));
  nand2 gate1256(.a(gate498inter8), .b(gate498inter7), .O(gate498inter9));
  nand2 gate1257(.a(s_101), .b(gate498inter3), .O(gate498inter10));
  nor2  gate1258(.a(gate498inter10), .b(gate498inter9), .O(gate498inter11));
  nor2  gate1259(.a(gate498inter11), .b(gate498inter6), .O(gate498inter12));
  nand2 gate1260(.a(gate498inter12), .b(gate498inter1), .O(G1307));

  xor2  gate911(.a(G1261), .b(G1260), .O(gate499inter0));
  nand2 gate912(.a(gate499inter0), .b(s_52), .O(gate499inter1));
  and2  gate913(.a(G1261), .b(G1260), .O(gate499inter2));
  inv1  gate914(.a(s_52), .O(gate499inter3));
  inv1  gate915(.a(s_53), .O(gate499inter4));
  nand2 gate916(.a(gate499inter4), .b(gate499inter3), .O(gate499inter5));
  nor2  gate917(.a(gate499inter5), .b(gate499inter2), .O(gate499inter6));
  inv1  gate918(.a(G1260), .O(gate499inter7));
  inv1  gate919(.a(G1261), .O(gate499inter8));
  nand2 gate920(.a(gate499inter8), .b(gate499inter7), .O(gate499inter9));
  nand2 gate921(.a(s_53), .b(gate499inter3), .O(gate499inter10));
  nor2  gate922(.a(gate499inter10), .b(gate499inter9), .O(gate499inter11));
  nor2  gate923(.a(gate499inter11), .b(gate499inter6), .O(gate499inter12));
  nand2 gate924(.a(gate499inter12), .b(gate499inter1), .O(G1308));
nand2 gate500( .a(G1262), .b(G1263), .O(G1309) );
nand2 gate501( .a(G1264), .b(G1265), .O(G1310) );

  xor2  gate967(.a(G1267), .b(G1266), .O(gate502inter0));
  nand2 gate968(.a(gate502inter0), .b(s_60), .O(gate502inter1));
  and2  gate969(.a(G1267), .b(G1266), .O(gate502inter2));
  inv1  gate970(.a(s_60), .O(gate502inter3));
  inv1  gate971(.a(s_61), .O(gate502inter4));
  nand2 gate972(.a(gate502inter4), .b(gate502inter3), .O(gate502inter5));
  nor2  gate973(.a(gate502inter5), .b(gate502inter2), .O(gate502inter6));
  inv1  gate974(.a(G1266), .O(gate502inter7));
  inv1  gate975(.a(G1267), .O(gate502inter8));
  nand2 gate976(.a(gate502inter8), .b(gate502inter7), .O(gate502inter9));
  nand2 gate977(.a(s_61), .b(gate502inter3), .O(gate502inter10));
  nor2  gate978(.a(gate502inter10), .b(gate502inter9), .O(gate502inter11));
  nor2  gate979(.a(gate502inter11), .b(gate502inter6), .O(gate502inter12));
  nand2 gate980(.a(gate502inter12), .b(gate502inter1), .O(G1311));

  xor2  gate2269(.a(G1269), .b(G1268), .O(gate503inter0));
  nand2 gate2270(.a(gate503inter0), .b(s_246), .O(gate503inter1));
  and2  gate2271(.a(G1269), .b(G1268), .O(gate503inter2));
  inv1  gate2272(.a(s_246), .O(gate503inter3));
  inv1  gate2273(.a(s_247), .O(gate503inter4));
  nand2 gate2274(.a(gate503inter4), .b(gate503inter3), .O(gate503inter5));
  nor2  gate2275(.a(gate503inter5), .b(gate503inter2), .O(gate503inter6));
  inv1  gate2276(.a(G1268), .O(gate503inter7));
  inv1  gate2277(.a(G1269), .O(gate503inter8));
  nand2 gate2278(.a(gate503inter8), .b(gate503inter7), .O(gate503inter9));
  nand2 gate2279(.a(s_247), .b(gate503inter3), .O(gate503inter10));
  nor2  gate2280(.a(gate503inter10), .b(gate503inter9), .O(gate503inter11));
  nor2  gate2281(.a(gate503inter11), .b(gate503inter6), .O(gate503inter12));
  nand2 gate2282(.a(gate503inter12), .b(gate503inter1), .O(G1312));
nand2 gate504( .a(G1270), .b(G1271), .O(G1313) );

  xor2  gate2535(.a(G1273), .b(G1272), .O(gate505inter0));
  nand2 gate2536(.a(gate505inter0), .b(s_284), .O(gate505inter1));
  and2  gate2537(.a(G1273), .b(G1272), .O(gate505inter2));
  inv1  gate2538(.a(s_284), .O(gate505inter3));
  inv1  gate2539(.a(s_285), .O(gate505inter4));
  nand2 gate2540(.a(gate505inter4), .b(gate505inter3), .O(gate505inter5));
  nor2  gate2541(.a(gate505inter5), .b(gate505inter2), .O(gate505inter6));
  inv1  gate2542(.a(G1272), .O(gate505inter7));
  inv1  gate2543(.a(G1273), .O(gate505inter8));
  nand2 gate2544(.a(gate505inter8), .b(gate505inter7), .O(gate505inter9));
  nand2 gate2545(.a(s_285), .b(gate505inter3), .O(gate505inter10));
  nor2  gate2546(.a(gate505inter10), .b(gate505inter9), .O(gate505inter11));
  nor2  gate2547(.a(gate505inter11), .b(gate505inter6), .O(gate505inter12));
  nand2 gate2548(.a(gate505inter12), .b(gate505inter1), .O(G1314));
nand2 gate506( .a(G1274), .b(G1275), .O(G1315) );

  xor2  gate771(.a(G1277), .b(G1276), .O(gate507inter0));
  nand2 gate772(.a(gate507inter0), .b(s_32), .O(gate507inter1));
  and2  gate773(.a(G1277), .b(G1276), .O(gate507inter2));
  inv1  gate774(.a(s_32), .O(gate507inter3));
  inv1  gate775(.a(s_33), .O(gate507inter4));
  nand2 gate776(.a(gate507inter4), .b(gate507inter3), .O(gate507inter5));
  nor2  gate777(.a(gate507inter5), .b(gate507inter2), .O(gate507inter6));
  inv1  gate778(.a(G1276), .O(gate507inter7));
  inv1  gate779(.a(G1277), .O(gate507inter8));
  nand2 gate780(.a(gate507inter8), .b(gate507inter7), .O(gate507inter9));
  nand2 gate781(.a(s_33), .b(gate507inter3), .O(gate507inter10));
  nor2  gate782(.a(gate507inter10), .b(gate507inter9), .O(gate507inter11));
  nor2  gate783(.a(gate507inter11), .b(gate507inter6), .O(gate507inter12));
  nand2 gate784(.a(gate507inter12), .b(gate507inter1), .O(G1316));
nand2 gate508( .a(G1278), .b(G1279), .O(G1317) );
nand2 gate509( .a(G1280), .b(G1281), .O(G1318) );
nand2 gate510( .a(G1282), .b(G1283), .O(G1319) );
nand2 gate511( .a(G1284), .b(G1285), .O(G1320) );
nand2 gate512( .a(G1286), .b(G1287), .O(G1321) );
nand2 gate513( .a(G1288), .b(G1289), .O(G1322) );
nand2 gate514( .a(G1290), .b(G1291), .O(G1323) );
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule