module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);

input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;//RE__PI;

input s_0,s_1;//RE__ALLOW(00,01,10,11);
input s_2,s_3;//RE__ALLOW(00,01,10,11);
input s_4,s_5;//RE__ALLOW(00,01,10,11);
input s_6,s_7;//RE__ALLOW(00,01,10,11);
input s_8,s_9;//RE__ALLOW(00,01,10,11);
input s_10,s_11;//RE__ALLOW(00,01,10,11);
input s_12,s_13;//RE__ALLOW(00,01,10,11);
input s_14,s_15;//RE__ALLOW(00,01,10,11);
input s_16,s_17;//RE__ALLOW(00,01,10,11);
input s_18,s_19;//RE__ALLOW(00,01,10,11);
input s_20,s_21;//RE__ALLOW(00,01,10,11);
input s_22,s_23;//RE__ALLOW(00,01,10,11);
input s_24,s_25;//RE__ALLOW(00,01,10,11);
input s_26,s_27;//RE__ALLOW(00,01,10,11);
input s_28,s_29;//RE__ALLOW(00,01,10,11);
input s_30,s_31;//RE__ALLOW(00,01,10,11);
input s_32,s_33;//RE__ALLOW(00,01,10,11);
input s_34,s_35;//RE__ALLOW(00,01,10,11);
input s_36,s_37;//RE__ALLOW(00,01,10,11);
input s_38,s_39;//RE__ALLOW(00,01,10,11);
input s_40,s_41;//RE__ALLOW(00,01,10,11);
input s_42,s_43;//RE__ALLOW(00,01,10,11);
input s_44,s_45;//RE__ALLOW(00,01,10,11);
input s_46,s_47;//RE__ALLOW(00,01,10,11);
input s_48,s_49;//RE__ALLOW(00,01,10,11);
input s_50,s_51;//RE__ALLOW(00,01,10,11);
input s_52,s_53;//RE__ALLOW(00,01,10,11);
input s_54,s_55;//RE__ALLOW(00,01,10,11);
input s_56,s_57;//RE__ALLOW(00,01,10,11);
input s_58,s_59;//RE__ALLOW(00,01,10,11);
input s_60,s_61;//RE__ALLOW(00,01,10,11);
input s_62,s_63;//RE__ALLOW(00,01,10,11);
input s_64,s_65;//RE__ALLOW(00,01,10,11);
input s_66,s_67;//RE__ALLOW(00,01,10,11);
input s_68,s_69;//RE__ALLOW(00,01,10,11);
input s_70,s_71;//RE__ALLOW(00,01,10,11);
input s_72,s_73;//RE__ALLOW(00,01,10,11);
input s_74,s_75;//RE__ALLOW(00,01,10,11);
input s_76,s_77;//RE__ALLOW(00,01,10,11);
input s_78,s_79;//RE__ALLOW(00,01,10,11);
input s_80,s_81;//RE__ALLOW(00,01,10,11);
input s_82,s_83;//RE__ALLOW(00,01,10,11);
input s_84,s_85;//RE__ALLOW(00,01,10,11);
input s_86,s_87;//RE__ALLOW(00,01,10,11);
input s_88,s_89;//RE__ALLOW(00,01,10,11);
input s_90,s_91;//RE__ALLOW(00,01,10,11);
input s_92,s_93;//RE__ALLOW(00,01,10,11);
input s_94,s_95;//RE__ALLOW(00,01,10,11);
input s_96,s_97;//RE__ALLOW(00,01,10,11);
input s_98,s_99;//RE__ALLOW(00,01,10,11);
input s_100,s_101;//RE__ALLOW(00,01,10,11);
input s_102,s_103;//RE__ALLOW(00,01,10,11);
input s_104,s_105;//RE__ALLOW(00,01,10,11);
input s_106,s_107;//RE__ALLOW(00,01,10,11);
input s_108,s_109;//RE__ALLOW(00,01,10,11);
input s_110,s_111;//RE__ALLOW(00,01,10,11);
input s_112,s_113;//RE__ALLOW(00,01,10,11);
input s_114,s_115;//RE__ALLOW(00,01,10,11);
input s_116,s_117;//RE__ALLOW(00,01,10,11);
input s_118,s_119;//RE__ALLOW(00,01,10,11);
input s_120,s_121;//RE__ALLOW(00,01,10,11);
input s_122,s_123;//RE__ALLOW(00,01,10,11);
input s_124,s_125;//RE__ALLOW(00,01,10,11);
input s_126,s_127;//RE__ALLOW(00,01,10,11);
input s_128,s_129;//RE__ALLOW(00,01,10,11);
input s_130,s_131;//RE__ALLOW(00,01,10,11);
input s_132,s_133;//RE__ALLOW(00,01,10,11);
input s_134,s_135;//RE__ALLOW(00,01,10,11);
input s_136,s_137;//RE__ALLOW(00,01,10,11);
input s_138,s_139;//RE__ALLOW(00,01,10,11);
input s_140,s_141;//RE__ALLOW(00,01,10,11);
input s_142,s_143;//RE__ALLOW(00,01,10,11);
input s_144,s_145;//RE__ALLOW(00,01,10,11);
input s_146,s_147;//RE__ALLOW(00,01,10,11);
input s_148,s_149;//RE__ALLOW(00,01,10,11);
input s_150,s_151;//RE__ALLOW(00,01,10,11);
input s_152,s_153;//RE__ALLOW(00,01,10,11);
input s_154,s_155;//RE__ALLOW(00,01,10,11);
input s_156,s_157;//RE__ALLOW(00,01,10,11);
input s_158,s_159;//RE__ALLOW(00,01,10,11);
input s_160,s_161;//RE__ALLOW(00,01,10,11);
input s_162,s_163;//RE__ALLOW(00,01,10,11);
input s_164,s_165;//RE__ALLOW(00,01,10,11);
input s_166,s_167;//RE__ALLOW(00,01,10,11);
input s_168,s_169;//RE__ALLOW(00,01,10,11);
input s_170,s_171;//RE__ALLOW(00,01,10,11);
input s_172,s_173;//RE__ALLOW(00,01,10,11);
input s_174,s_175;//RE__ALLOW(00,01,10,11);
input s_176,s_177;//RE__ALLOW(00,01,10,11);
input s_178,s_179;//RE__ALLOW(00,01,10,11);
input s_180,s_181;//RE__ALLOW(00,01,10,11);
input s_182,s_183;//RE__ALLOW(00,01,10,11);
input s_184,s_185;//RE__ALLOW(00,01,10,11);
input s_186,s_187;//RE__ALLOW(00,01,10,11);
input s_188,s_189;//RE__ALLOW(00,01,10,11);
input s_190,s_191;//RE__ALLOW(00,01,10,11);
input s_192,s_193;//RE__ALLOW(00,01,10,11);
input s_194,s_195;//RE__ALLOW(00,01,10,11);
input s_196,s_197;//RE__ALLOW(00,01,10,11);
input s_198,s_199;//RE__ALLOW(00,01,10,11);
input s_200,s_201;//RE__ALLOW(00,01,10,11);
input s_202,s_203;//RE__ALLOW(00,01,10,11);
input s_204,s_205;//RE__ALLOW(00,01,10,11);
input s_206,s_207;//RE__ALLOW(00,01,10,11);
input s_208,s_209;//RE__ALLOW(00,01,10,11);
input s_210,s_211;//RE__ALLOW(00,01,10,11);
input s_212,s_213;//RE__ALLOW(00,01,10,11);
input s_214,s_215;//RE__ALLOW(00,01,10,11);
input s_216,s_217;//RE__ALLOW(00,01,10,11);
input s_218,s_219;//RE__ALLOW(00,01,10,11);
input s_220,s_221;//RE__ALLOW(00,01,10,11);
input s_222,s_223;//RE__ALLOW(00,01,10,11);
input s_224,s_225;//RE__ALLOW(00,01,10,11);
input s_226,s_227;//RE__ALLOW(00,01,10,11);
input s_228,s_229;//RE__ALLOW(00,01,10,11);
input s_230,s_231;//RE__ALLOW(00,01,10,11);
input s_232,s_233;//RE__ALLOW(00,01,10,11);
input s_234,s_235;//RE__ALLOW(00,01,10,11);
input s_236,s_237;//RE__ALLOW(00,01,10,11);
input s_238,s_239;//RE__ALLOW(00,01,10,11);
input s_240,s_241;//RE__ALLOW(00,01,10,11);
input s_242,s_243;//RE__ALLOW(00,01,10,11);
input s_244,s_245;//RE__ALLOW(00,01,10,11);
input s_246,s_247;//RE__ALLOW(00,01,10,11);
input s_248,s_249;//RE__ALLOW(00,01,10,11);
input s_250,s_251;//RE__ALLOW(00,01,10,11);
input s_252,s_253;//RE__ALLOW(00,01,10,11);
input s_254,s_255;//RE__ALLOW(00,01,10,11);
input s_256,s_257;//RE__ALLOW(00,01,10,11);
input s_258,s_259;//RE__ALLOW(00,01,10,11);
input s_260,s_261;//RE__ALLOW(00,01,10,11);
input s_262,s_263;//RE__ALLOW(00,01,10,11);
input s_264,s_265;//RE__ALLOW(00,01,10,11);
input s_266,s_267;//RE__ALLOW(00,01,10,11);
input s_268,s_269;//RE__ALLOW(00,01,10,11);
input s_270,s_271;//RE__ALLOW(00,01,10,11);
input s_272,s_273;//RE__ALLOW(00,01,10,11);
input s_274,s_275;//RE__ALLOW(00,01,10,11);
input s_276,s_277;//RE__ALLOW(00,01,10,11);
input s_278,s_279;//RE__ALLOW(00,01,10,11);
input s_280,s_281;//RE__ALLOW(00,01,10,11);
input s_282,s_283;//RE__ALLOW(00,01,10,11);
input s_284,s_285;//RE__ALLOW(00,01,10,11);
input s_286,s_287;//RE__ALLOW(00,01,10,11);
input s_288,s_289;//RE__ALLOW(00,01,10,11);
input s_290,s_291;//RE__ALLOW(00,01,10,11);
input s_292,s_293;//RE__ALLOW(00,01,10,11);
input s_294,s_295;//RE__ALLOW(00,01,10,11);
input s_296,s_297;//RE__ALLOW(00,01,10,11);
input s_298,s_299;//RE__ALLOW(00,01,10,11);
input s_300,s_301;//RE__ALLOW(00,01,10,11);
input s_302,s_303;//RE__ALLOW(00,01,10,11);
input s_304,s_305;//RE__ALLOW(00,01,10,11);
input s_306,s_307;//RE__ALLOW(00,01,10,11);
input s_308,s_309;//RE__ALLOW(00,01,10,11);
input s_310,s_311;//RE__ALLOW(00,01,10,11);
input s_312,s_313;//RE__ALLOW(00,01,10,11);
input s_314,s_315;//RE__ALLOW(00,01,10,11);
input s_316,s_317;//RE__ALLOW(00,01,10,11);
input s_318,s_319;//RE__ALLOW(00,01,10,11);
input s_320,s_321;//RE__ALLOW(00,01,10,11);
input s_322,s_323;//RE__ALLOW(00,01,10,11);
input s_324,s_325;//RE__ALLOW(00,01,10,11);
input s_326,s_327;//RE__ALLOW(00,01,10,11);
input s_328,s_329;//RE__ALLOW(00,01,10,11);
input s_330,s_331;//RE__ALLOW(00,01,10,11);
input s_332,s_333;//RE__ALLOW(00,01,10,11);
input s_334,s_335;//RE__ALLOW(00,01,10,11);
input s_336,s_337;//RE__ALLOW(00,01,10,11);
input s_338,s_339;//RE__ALLOW(00,01,10,11);
input s_340,s_341;//RE__ALLOW(00,01,10,11);
input s_342,s_343;//RE__ALLOW(00,01,10,11);
input s_344,s_345;//RE__ALLOW(00,01,10,11);
input s_346,s_347;//RE__ALLOW(00,01,10,11);
input s_348,s_349;//RE__ALLOW(00,01,10,11);
input s_350,s_351;//RE__ALLOW(00,01,10,11);
input s_352,s_353;//RE__ALLOW(00,01,10,11);
input s_354,s_355;//RE__ALLOW(00,01,10,11);
input s_356,s_357;//RE__ALLOW(00,01,10,11);
input s_358,s_359;//RE__ALLOW(00,01,10,11);
input s_360,s_361;//RE__ALLOW(00,01,10,11);
input s_362,s_363;//RE__ALLOW(00,01,10,11);
input s_364,s_365;//RE__ALLOW(00,01,10,11);
input s_366,s_367;//RE__ALLOW(00,01,10,11);
input s_368,s_369;//RE__ALLOW(00,01,10,11);
input s_370,s_371;//RE__ALLOW(00,01,10,11);
input s_372,s_373;//RE__ALLOW(00,01,10,11);
input s_374,s_375;//RE__ALLOW(00,01,10,11);
input s_376,s_377;//RE__ALLOW(00,01,10,11);
input s_378,s_379;//RE__ALLOW(00,01,10,11);
input s_380,s_381;//RE__ALLOW(00,01,10,11);
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;

  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate253inter0, gate253inter1, gate253inter2, gate253inter3, gate253inter4, gate253inter5, gate253inter6, gate253inter7, gate253inter8, gate253inter9, gate253inter10, gate253inter11, gate253inter12, gate496inter0, gate496inter1, gate496inter2, gate496inter3, gate496inter4, gate496inter5, gate496inter6, gate496inter7, gate496inter8, gate496inter9, gate496inter10, gate496inter11, gate496inter12, gate85inter0, gate85inter1, gate85inter2, gate85inter3, gate85inter4, gate85inter5, gate85inter6, gate85inter7, gate85inter8, gate85inter9, gate85inter10, gate85inter11, gate85inter12, gate228inter0, gate228inter1, gate228inter2, gate228inter3, gate228inter4, gate228inter5, gate228inter6, gate228inter7, gate228inter8, gate228inter9, gate228inter10, gate228inter11, gate228inter12, gate84inter0, gate84inter1, gate84inter2, gate84inter3, gate84inter4, gate84inter5, gate84inter6, gate84inter7, gate84inter8, gate84inter9, gate84inter10, gate84inter11, gate84inter12, gate186inter0, gate186inter1, gate186inter2, gate186inter3, gate186inter4, gate186inter5, gate186inter6, gate186inter7, gate186inter8, gate186inter9, gate186inter10, gate186inter11, gate186inter12, gate154inter0, gate154inter1, gate154inter2, gate154inter3, gate154inter4, gate154inter5, gate154inter6, gate154inter7, gate154inter8, gate154inter9, gate154inter10, gate154inter11, gate154inter12, gate474inter0, gate474inter1, gate474inter2, gate474inter3, gate474inter4, gate474inter5, gate474inter6, gate474inter7, gate474inter8, gate474inter9, gate474inter10, gate474inter11, gate474inter12, gate129inter0, gate129inter1, gate129inter2, gate129inter3, gate129inter4, gate129inter5, gate129inter6, gate129inter7, gate129inter8, gate129inter9, gate129inter10, gate129inter11, gate129inter12, gate499inter0, gate499inter1, gate499inter2, gate499inter3, gate499inter4, gate499inter5, gate499inter6, gate499inter7, gate499inter8, gate499inter9, gate499inter10, gate499inter11, gate499inter12, gate225inter0, gate225inter1, gate225inter2, gate225inter3, gate225inter4, gate225inter5, gate225inter6, gate225inter7, gate225inter8, gate225inter9, gate225inter10, gate225inter11, gate225inter12, gate259inter0, gate259inter1, gate259inter2, gate259inter3, gate259inter4, gate259inter5, gate259inter6, gate259inter7, gate259inter8, gate259inter9, gate259inter10, gate259inter11, gate259inter12, gate189inter0, gate189inter1, gate189inter2, gate189inter3, gate189inter4, gate189inter5, gate189inter6, gate189inter7, gate189inter8, gate189inter9, gate189inter10, gate189inter11, gate189inter12, gate270inter0, gate270inter1, gate270inter2, gate270inter3, gate270inter4, gate270inter5, gate270inter6, gate270inter7, gate270inter8, gate270inter9, gate270inter10, gate270inter11, gate270inter12, gate292inter0, gate292inter1, gate292inter2, gate292inter3, gate292inter4, gate292inter5, gate292inter6, gate292inter7, gate292inter8, gate292inter9, gate292inter10, gate292inter11, gate292inter12, gate188inter0, gate188inter1, gate188inter2, gate188inter3, gate188inter4, gate188inter5, gate188inter6, gate188inter7, gate188inter8, gate188inter9, gate188inter10, gate188inter11, gate188inter12, gate512inter0, gate512inter1, gate512inter2, gate512inter3, gate512inter4, gate512inter5, gate512inter6, gate512inter7, gate512inter8, gate512inter9, gate512inter10, gate512inter11, gate512inter12, gate185inter0, gate185inter1, gate185inter2, gate185inter3, gate185inter4, gate185inter5, gate185inter6, gate185inter7, gate185inter8, gate185inter9, gate185inter10, gate185inter11, gate185inter12, gate424inter0, gate424inter1, gate424inter2, gate424inter3, gate424inter4, gate424inter5, gate424inter6, gate424inter7, gate424inter8, gate424inter9, gate424inter10, gate424inter11, gate424inter12, gate508inter0, gate508inter1, gate508inter2, gate508inter3, gate508inter4, gate508inter5, gate508inter6, gate508inter7, gate508inter8, gate508inter9, gate508inter10, gate508inter11, gate508inter12, gate427inter0, gate427inter1, gate427inter2, gate427inter3, gate427inter4, gate427inter5, gate427inter6, gate427inter7, gate427inter8, gate427inter9, gate427inter10, gate427inter11, gate427inter12, gate75inter0, gate75inter1, gate75inter2, gate75inter3, gate75inter4, gate75inter5, gate75inter6, gate75inter7, gate75inter8, gate75inter9, gate75inter10, gate75inter11, gate75inter12, gate231inter0, gate231inter1, gate231inter2, gate231inter3, gate231inter4, gate231inter5, gate231inter6, gate231inter7, gate231inter8, gate231inter9, gate231inter10, gate231inter11, gate231inter12, gate266inter0, gate266inter1, gate266inter2, gate266inter3, gate266inter4, gate266inter5, gate266inter6, gate266inter7, gate266inter8, gate266inter9, gate266inter10, gate266inter11, gate266inter12, gate490inter0, gate490inter1, gate490inter2, gate490inter3, gate490inter4, gate490inter5, gate490inter6, gate490inter7, gate490inter8, gate490inter9, gate490inter10, gate490inter11, gate490inter12, gate242inter0, gate242inter1, gate242inter2, gate242inter3, gate242inter4, gate242inter5, gate242inter6, gate242inter7, gate242inter8, gate242inter9, gate242inter10, gate242inter11, gate242inter12, gate83inter0, gate83inter1, gate83inter2, gate83inter3, gate83inter4, gate83inter5, gate83inter6, gate83inter7, gate83inter8, gate83inter9, gate83inter10, gate83inter11, gate83inter12, gate86inter0, gate86inter1, gate86inter2, gate86inter3, gate86inter4, gate86inter5, gate86inter6, gate86inter7, gate86inter8, gate86inter9, gate86inter10, gate86inter11, gate86inter12, gate466inter0, gate466inter1, gate466inter2, gate466inter3, gate466inter4, gate466inter5, gate466inter6, gate466inter7, gate466inter8, gate466inter9, gate466inter10, gate466inter11, gate466inter12, gate180inter0, gate180inter1, gate180inter2, gate180inter3, gate180inter4, gate180inter5, gate180inter6, gate180inter7, gate180inter8, gate180inter9, gate180inter10, gate180inter11, gate180inter12, gate182inter0, gate182inter1, gate182inter2, gate182inter3, gate182inter4, gate182inter5, gate182inter6, gate182inter7, gate182inter8, gate182inter9, gate182inter10, gate182inter11, gate182inter12, gate82inter0, gate82inter1, gate82inter2, gate82inter3, gate82inter4, gate82inter5, gate82inter6, gate82inter7, gate82inter8, gate82inter9, gate82inter10, gate82inter11, gate82inter12, gate124inter0, gate124inter1, gate124inter2, gate124inter3, gate124inter4, gate124inter5, gate124inter6, gate124inter7, gate124inter8, gate124inter9, gate124inter10, gate124inter11, gate124inter12, gate23inter0, gate23inter1, gate23inter2, gate23inter3, gate23inter4, gate23inter5, gate23inter6, gate23inter7, gate23inter8, gate23inter9, gate23inter10, gate23inter11, gate23inter12, gate422inter0, gate422inter1, gate422inter2, gate422inter3, gate422inter4, gate422inter5, gate422inter6, gate422inter7, gate422inter8, gate422inter9, gate422inter10, gate422inter11, gate422inter12, gate407inter0, gate407inter1, gate407inter2, gate407inter3, gate407inter4, gate407inter5, gate407inter6, gate407inter7, gate407inter8, gate407inter9, gate407inter10, gate407inter11, gate407inter12, gate200inter0, gate200inter1, gate200inter2, gate200inter3, gate200inter4, gate200inter5, gate200inter6, gate200inter7, gate200inter8, gate200inter9, gate200inter10, gate200inter11, gate200inter12, gate212inter0, gate212inter1, gate212inter2, gate212inter3, gate212inter4, gate212inter5, gate212inter6, gate212inter7, gate212inter8, gate212inter9, gate212inter10, gate212inter11, gate212inter12, gate435inter0, gate435inter1, gate435inter2, gate435inter3, gate435inter4, gate435inter5, gate435inter6, gate435inter7, gate435inter8, gate435inter9, gate435inter10, gate435inter11, gate435inter12, gate101inter0, gate101inter1, gate101inter2, gate101inter3, gate101inter4, gate101inter5, gate101inter6, gate101inter7, gate101inter8, gate101inter9, gate101inter10, gate101inter11, gate101inter12, gate110inter0, gate110inter1, gate110inter2, gate110inter3, gate110inter4, gate110inter5, gate110inter6, gate110inter7, gate110inter8, gate110inter9, gate110inter10, gate110inter11, gate110inter12, gate463inter0, gate463inter1, gate463inter2, gate463inter3, gate463inter4, gate463inter5, gate463inter6, gate463inter7, gate463inter8, gate463inter9, gate463inter10, gate463inter11, gate463inter12, gate462inter0, gate462inter1, gate462inter2, gate462inter3, gate462inter4, gate462inter5, gate462inter6, gate462inter7, gate462inter8, gate462inter9, gate462inter10, gate462inter11, gate462inter12, gate15inter0, gate15inter1, gate15inter2, gate15inter3, gate15inter4, gate15inter5, gate15inter6, gate15inter7, gate15inter8, gate15inter9, gate15inter10, gate15inter11, gate15inter12, gate414inter0, gate414inter1, gate414inter2, gate414inter3, gate414inter4, gate414inter5, gate414inter6, gate414inter7, gate414inter8, gate414inter9, gate414inter10, gate414inter11, gate414inter12, gate61inter0, gate61inter1, gate61inter2, gate61inter3, gate61inter4, gate61inter5, gate61inter6, gate61inter7, gate61inter8, gate61inter9, gate61inter10, gate61inter11, gate61inter12, gate433inter0, gate433inter1, gate433inter2, gate433inter3, gate433inter4, gate433inter5, gate433inter6, gate433inter7, gate433inter8, gate433inter9, gate433inter10, gate433inter11, gate433inter12, gate421inter0, gate421inter1, gate421inter2, gate421inter3, gate421inter4, gate421inter5, gate421inter6, gate421inter7, gate421inter8, gate421inter9, gate421inter10, gate421inter11, gate421inter12, gate254inter0, gate254inter1, gate254inter2, gate254inter3, gate254inter4, gate254inter5, gate254inter6, gate254inter7, gate254inter8, gate254inter9, gate254inter10, gate254inter11, gate254inter12, gate472inter0, gate472inter1, gate472inter2, gate472inter3, gate472inter4, gate472inter5, gate472inter6, gate472inter7, gate472inter8, gate472inter9, gate472inter10, gate472inter11, gate472inter12, gate509inter0, gate509inter1, gate509inter2, gate509inter3, gate509inter4, gate509inter5, gate509inter6, gate509inter7, gate509inter8, gate509inter9, gate509inter10, gate509inter11, gate509inter12, gate41inter0, gate41inter1, gate41inter2, gate41inter3, gate41inter4, gate41inter5, gate41inter6, gate41inter7, gate41inter8, gate41inter9, gate41inter10, gate41inter11, gate41inter12, gate208inter0, gate208inter1, gate208inter2, gate208inter3, gate208inter4, gate208inter5, gate208inter6, gate208inter7, gate208inter8, gate208inter9, gate208inter10, gate208inter11, gate208inter12, gate505inter0, gate505inter1, gate505inter2, gate505inter3, gate505inter4, gate505inter5, gate505inter6, gate505inter7, gate505inter8, gate505inter9, gate505inter10, gate505inter11, gate505inter12, gate88inter0, gate88inter1, gate88inter2, gate88inter3, gate88inter4, gate88inter5, gate88inter6, gate88inter7, gate88inter8, gate88inter9, gate88inter10, gate88inter11, gate88inter12, gate152inter0, gate152inter1, gate152inter2, gate152inter3, gate152inter4, gate152inter5, gate152inter6, gate152inter7, gate152inter8, gate152inter9, gate152inter10, gate152inter11, gate152inter12, gate477inter0, gate477inter1, gate477inter2, gate477inter3, gate477inter4, gate477inter5, gate477inter6, gate477inter7, gate477inter8, gate477inter9, gate477inter10, gate477inter11, gate477inter12, gate513inter0, gate513inter1, gate513inter2, gate513inter3, gate513inter4, gate513inter5, gate513inter6, gate513inter7, gate513inter8, gate513inter9, gate513inter10, gate513inter11, gate513inter12, gate222inter0, gate222inter1, gate222inter2, gate222inter3, gate222inter4, gate222inter5, gate222inter6, gate222inter7, gate222inter8, gate222inter9, gate222inter10, gate222inter11, gate222inter12, gate221inter0, gate221inter1, gate221inter2, gate221inter3, gate221inter4, gate221inter5, gate221inter6, gate221inter7, gate221inter8, gate221inter9, gate221inter10, gate221inter11, gate221inter12, gate166inter0, gate166inter1, gate166inter2, gate166inter3, gate166inter4, gate166inter5, gate166inter6, gate166inter7, gate166inter8, gate166inter9, gate166inter10, gate166inter11, gate166inter12, gate402inter0, gate402inter1, gate402inter2, gate402inter3, gate402inter4, gate402inter5, gate402inter6, gate402inter7, gate402inter8, gate402inter9, gate402inter10, gate402inter11, gate402inter12, gate149inter0, gate149inter1, gate149inter2, gate149inter3, gate149inter4, gate149inter5, gate149inter6, gate149inter7, gate149inter8, gate149inter9, gate149inter10, gate149inter11, gate149inter12, gate106inter0, gate106inter1, gate106inter2, gate106inter3, gate106inter4, gate106inter5, gate106inter6, gate106inter7, gate106inter8, gate106inter9, gate106inter10, gate106inter11, gate106inter12, gate159inter0, gate159inter1, gate159inter2, gate159inter3, gate159inter4, gate159inter5, gate159inter6, gate159inter7, gate159inter8, gate159inter9, gate159inter10, gate159inter11, gate159inter12, gate487inter0, gate487inter1, gate487inter2, gate487inter3, gate487inter4, gate487inter5, gate487inter6, gate487inter7, gate487inter8, gate487inter9, gate487inter10, gate487inter11, gate487inter12, gate249inter0, gate249inter1, gate249inter2, gate249inter3, gate249inter4, gate249inter5, gate249inter6, gate249inter7, gate249inter8, gate249inter9, gate249inter10, gate249inter11, gate249inter12, gate287inter0, gate287inter1, gate287inter2, gate287inter3, gate287inter4, gate287inter5, gate287inter6, gate287inter7, gate287inter8, gate287inter9, gate287inter10, gate287inter11, gate287inter12, gate125inter0, gate125inter1, gate125inter2, gate125inter3, gate125inter4, gate125inter5, gate125inter6, gate125inter7, gate125inter8, gate125inter9, gate125inter10, gate125inter11, gate125inter12, gate410inter0, gate410inter1, gate410inter2, gate410inter3, gate410inter4, gate410inter5, gate410inter6, gate410inter7, gate410inter8, gate410inter9, gate410inter10, gate410inter11, gate410inter12, gate54inter0, gate54inter1, gate54inter2, gate54inter3, gate54inter4, gate54inter5, gate54inter6, gate54inter7, gate54inter8, gate54inter9, gate54inter10, gate54inter11, gate54inter12, gate501inter0, gate501inter1, gate501inter2, gate501inter3, gate501inter4, gate501inter5, gate501inter6, gate501inter7, gate501inter8, gate501inter9, gate501inter10, gate501inter11, gate501inter12, gate139inter0, gate139inter1, gate139inter2, gate139inter3, gate139inter4, gate139inter5, gate139inter6, gate139inter7, gate139inter8, gate139inter9, gate139inter10, gate139inter11, gate139inter12, gate36inter0, gate36inter1, gate36inter2, gate36inter3, gate36inter4, gate36inter5, gate36inter6, gate36inter7, gate36inter8, gate36inter9, gate36inter10, gate36inter11, gate36inter12, gate449inter0, gate449inter1, gate449inter2, gate449inter3, gate449inter4, gate449inter5, gate449inter6, gate449inter7, gate449inter8, gate449inter9, gate449inter10, gate449inter11, gate449inter12, gate48inter0, gate48inter1, gate48inter2, gate48inter3, gate48inter4, gate48inter5, gate48inter6, gate48inter7, gate48inter8, gate48inter9, gate48inter10, gate48inter11, gate48inter12, gate406inter0, gate406inter1, gate406inter2, gate406inter3, gate406inter4, gate406inter5, gate406inter6, gate406inter7, gate406inter8, gate406inter9, gate406inter10, gate406inter11, gate406inter12, gate121inter0, gate121inter1, gate121inter2, gate121inter3, gate121inter4, gate121inter5, gate121inter6, gate121inter7, gate121inter8, gate121inter9, gate121inter10, gate121inter11, gate121inter12, gate243inter0, gate243inter1, gate243inter2, gate243inter3, gate243inter4, gate243inter5, gate243inter6, gate243inter7, gate243inter8, gate243inter9, gate243inter10, gate243inter11, gate243inter12, gate459inter0, gate459inter1, gate459inter2, gate459inter3, gate459inter4, gate459inter5, gate459inter6, gate459inter7, gate459inter8, gate459inter9, gate459inter10, gate459inter11, gate459inter12, gate90inter0, gate90inter1, gate90inter2, gate90inter3, gate90inter4, gate90inter5, gate90inter6, gate90inter7, gate90inter8, gate90inter9, gate90inter10, gate90inter11, gate90inter12, gate94inter0, gate94inter1, gate94inter2, gate94inter3, gate94inter4, gate94inter5, gate94inter6, gate94inter7, gate94inter8, gate94inter9, gate94inter10, gate94inter11, gate94inter12, gate290inter0, gate290inter1, gate290inter2, gate290inter3, gate290inter4, gate290inter5, gate290inter6, gate290inter7, gate290inter8, gate290inter9, gate290inter10, gate290inter11, gate290inter12, gate284inter0, gate284inter1, gate284inter2, gate284inter3, gate284inter4, gate284inter5, gate284inter6, gate284inter7, gate284inter8, gate284inter9, gate284inter10, gate284inter11, gate284inter12, gate268inter0, gate268inter1, gate268inter2, gate268inter3, gate268inter4, gate268inter5, gate268inter6, gate268inter7, gate268inter8, gate268inter9, gate268inter10, gate268inter11, gate268inter12, gate251inter0, gate251inter1, gate251inter2, gate251inter3, gate251inter4, gate251inter5, gate251inter6, gate251inter7, gate251inter8, gate251inter9, gate251inter10, gate251inter11, gate251inter12, gate409inter0, gate409inter1, gate409inter2, gate409inter3, gate409inter4, gate409inter5, gate409inter6, gate409inter7, gate409inter8, gate409inter9, gate409inter10, gate409inter11, gate409inter12, gate181inter0, gate181inter1, gate181inter2, gate181inter3, gate181inter4, gate181inter5, gate181inter6, gate181inter7, gate181inter8, gate181inter9, gate181inter10, gate181inter11, gate181inter12, gate190inter0, gate190inter1, gate190inter2, gate190inter3, gate190inter4, gate190inter5, gate190inter6, gate190inter7, gate190inter8, gate190inter9, gate190inter10, gate190inter11, gate190inter12, gate137inter0, gate137inter1, gate137inter2, gate137inter3, gate137inter4, gate137inter5, gate137inter6, gate137inter7, gate137inter8, gate137inter9, gate137inter10, gate137inter11, gate137inter12, gate436inter0, gate436inter1, gate436inter2, gate436inter3, gate436inter4, gate436inter5, gate436inter6, gate436inter7, gate436inter8, gate436inter9, gate436inter10, gate436inter11, gate436inter12, gate395inter0, gate395inter1, gate395inter2, gate395inter3, gate395inter4, gate395inter5, gate395inter6, gate395inter7, gate395inter8, gate395inter9, gate395inter10, gate395inter11, gate395inter12, gate145inter0, gate145inter1, gate145inter2, gate145inter3, gate145inter4, gate145inter5, gate145inter6, gate145inter7, gate145inter8, gate145inter9, gate145inter10, gate145inter11, gate145inter12, gate419inter0, gate419inter1, gate419inter2, gate419inter3, gate419inter4, gate419inter5, gate419inter6, gate419inter7, gate419inter8, gate419inter9, gate419inter10, gate419inter11, gate419inter12, gate162inter0, gate162inter1, gate162inter2, gate162inter3, gate162inter4, gate162inter5, gate162inter6, gate162inter7, gate162inter8, gate162inter9, gate162inter10, gate162inter11, gate162inter12, gate43inter0, gate43inter1, gate43inter2, gate43inter3, gate43inter4, gate43inter5, gate43inter6, gate43inter7, gate43inter8, gate43inter9, gate43inter10, gate43inter11, gate43inter12, gate482inter0, gate482inter1, gate482inter2, gate482inter3, gate482inter4, gate482inter5, gate482inter6, gate482inter7, gate482inter8, gate482inter9, gate482inter10, gate482inter11, gate482inter12, gate510inter0, gate510inter1, gate510inter2, gate510inter3, gate510inter4, gate510inter5, gate510inter6, gate510inter7, gate510inter8, gate510inter9, gate510inter10, gate510inter11, gate510inter12, gate46inter0, gate46inter1, gate46inter2, gate46inter3, gate46inter4, gate46inter5, gate46inter6, gate46inter7, gate46inter8, gate46inter9, gate46inter10, gate46inter11, gate46inter12, gate42inter0, gate42inter1, gate42inter2, gate42inter3, gate42inter4, gate42inter5, gate42inter6, gate42inter7, gate42inter8, gate42inter9, gate42inter10, gate42inter11, gate42inter12, gate64inter0, gate64inter1, gate64inter2, gate64inter3, gate64inter4, gate64inter5, gate64inter6, gate64inter7, gate64inter8, gate64inter9, gate64inter10, gate64inter11, gate64inter12, gate282inter0, gate282inter1, gate282inter2, gate282inter3, gate282inter4, gate282inter5, gate282inter6, gate282inter7, gate282inter8, gate282inter9, gate282inter10, gate282inter11, gate282inter12, gate485inter0, gate485inter1, gate485inter2, gate485inter3, gate485inter4, gate485inter5, gate485inter6, gate485inter7, gate485inter8, gate485inter9, gate485inter10, gate485inter11, gate485inter12, gate105inter0, gate105inter1, gate105inter2, gate105inter3, gate105inter4, gate105inter5, gate105inter6, gate105inter7, gate105inter8, gate105inter9, gate105inter10, gate105inter11, gate105inter12, gate398inter0, gate398inter1, gate398inter2, gate398inter3, gate398inter4, gate398inter5, gate398inter6, gate398inter7, gate398inter8, gate398inter9, gate398inter10, gate398inter11, gate398inter12, gate173inter0, gate173inter1, gate173inter2, gate173inter3, gate173inter4, gate173inter5, gate173inter6, gate173inter7, gate173inter8, gate173inter9, gate173inter10, gate173inter11, gate173inter12, gate263inter0, gate263inter1, gate263inter2, gate263inter3, gate263inter4, gate263inter5, gate263inter6, gate263inter7, gate263inter8, gate263inter9, gate263inter10, gate263inter11, gate263inter12, gate128inter0, gate128inter1, gate128inter2, gate128inter3, gate128inter4, gate128inter5, gate128inter6, gate128inter7, gate128inter8, gate128inter9, gate128inter10, gate128inter11, gate128inter12, gate63inter0, gate63inter1, gate63inter2, gate63inter3, gate63inter4, gate63inter5, gate63inter6, gate63inter7, gate63inter8, gate63inter9, gate63inter10, gate63inter11, gate63inter12, gate514inter0, gate514inter1, gate514inter2, gate514inter3, gate514inter4, gate514inter5, gate514inter6, gate514inter7, gate514inter8, gate514inter9, gate514inter10, gate514inter11, gate514inter12, gate469inter0, gate469inter1, gate469inter2, gate469inter3, gate469inter4, gate469inter5, gate469inter6, gate469inter7, gate469inter8, gate469inter9, gate469inter10, gate469inter11, gate469inter12, gate25inter0, gate25inter1, gate25inter2, gate25inter3, gate25inter4, gate25inter5, gate25inter6, gate25inter7, gate25inter8, gate25inter9, gate25inter10, gate25inter11, gate25inter12, gate39inter0, gate39inter1, gate39inter2, gate39inter3, gate39inter4, gate39inter5, gate39inter6, gate39inter7, gate39inter8, gate39inter9, gate39inter10, gate39inter11, gate39inter12, gate224inter0, gate224inter1, gate224inter2, gate224inter3, gate224inter4, gate224inter5, gate224inter6, gate224inter7, gate224inter8, gate224inter9, gate224inter10, gate224inter11, gate224inter12, gate118inter0, gate118inter1, gate118inter2, gate118inter3, gate118inter4, gate118inter5, gate118inter6, gate118inter7, gate118inter8, gate118inter9, gate118inter10, gate118inter11, gate118inter12, gate34inter0, gate34inter1, gate34inter2, gate34inter3, gate34inter4, gate34inter5, gate34inter6, gate34inter7, gate34inter8, gate34inter9, gate34inter10, gate34inter11, gate34inter12, gate50inter0, gate50inter1, gate50inter2, gate50inter3, gate50inter4, gate50inter5, gate50inter6, gate50inter7, gate50inter8, gate50inter9, gate50inter10, gate50inter11, gate50inter12, gate205inter0, gate205inter1, gate205inter2, gate205inter3, gate205inter4, gate205inter5, gate205inter6, gate205inter7, gate205inter8, gate205inter9, gate205inter10, gate205inter11, gate205inter12, gate471inter0, gate471inter1, gate471inter2, gate471inter3, gate471inter4, gate471inter5, gate471inter6, gate471inter7, gate471inter8, gate471inter9, gate471inter10, gate471inter11, gate471inter12, gate241inter0, gate241inter1, gate241inter2, gate241inter3, gate241inter4, gate241inter5, gate241inter6, gate241inter7, gate241inter8, gate241inter9, gate241inter10, gate241inter11, gate241inter12, gate28inter0, gate28inter1, gate28inter2, gate28inter3, gate28inter4, gate28inter5, gate28inter6, gate28inter7, gate28inter8, gate28inter9, gate28inter10, gate28inter11, gate28inter12, gate73inter0, gate73inter1, gate73inter2, gate73inter3, gate73inter4, gate73inter5, gate73inter6, gate73inter7, gate73inter8, gate73inter9, gate73inter10, gate73inter11, gate73inter12, gate47inter0, gate47inter1, gate47inter2, gate47inter3, gate47inter4, gate47inter5, gate47inter6, gate47inter7, gate47inter8, gate47inter9, gate47inter10, gate47inter11, gate47inter12, gate96inter0, gate96inter1, gate96inter2, gate96inter3, gate96inter4, gate96inter5, gate96inter6, gate96inter7, gate96inter8, gate96inter9, gate96inter10, gate96inter11, gate96inter12, gate440inter0, gate440inter1, gate440inter2, gate440inter3, gate440inter4, gate440inter5, gate440inter6, gate440inter7, gate440inter8, gate440inter9, gate440inter10, gate440inter11, gate440inter12, gate286inter0, gate286inter1, gate286inter2, gate286inter3, gate286inter4, gate286inter5, gate286inter6, gate286inter7, gate286inter8, gate286inter9, gate286inter10, gate286inter11, gate286inter12, gate156inter0, gate156inter1, gate156inter2, gate156inter3, gate156inter4, gate156inter5, gate156inter6, gate156inter7, gate156inter8, gate156inter9, gate156inter10, gate156inter11, gate156inter12, gate493inter0, gate493inter1, gate493inter2, gate493inter3, gate493inter4, gate493inter5, gate493inter6, gate493inter7, gate493inter8, gate493inter9, gate493inter10, gate493inter11, gate493inter12, gate445inter0, gate445inter1, gate445inter2, gate445inter3, gate445inter4, gate445inter5, gate445inter6, gate445inter7, gate445inter8, gate445inter9, gate445inter10, gate445inter11, gate445inter12, gate494inter0, gate494inter1, gate494inter2, gate494inter3, gate494inter4, gate494inter5, gate494inter6, gate494inter7, gate494inter8, gate494inter9, gate494inter10, gate494inter11, gate494inter12, gate148inter0, gate148inter1, gate148inter2, gate148inter3, gate148inter4, gate148inter5, gate148inter6, gate148inter7, gate148inter8, gate148inter9, gate148inter10, gate148inter11, gate148inter12, gate403inter0, gate403inter1, gate403inter2, gate403inter3, gate403inter4, gate403inter5, gate403inter6, gate403inter7, gate403inter8, gate403inter9, gate403inter10, gate403inter11, gate403inter12, gate206inter0, gate206inter1, gate206inter2, gate206inter3, gate206inter4, gate206inter5, gate206inter6, gate206inter7, gate206inter8, gate206inter9, gate206inter10, gate206inter11, gate206inter12, gate167inter0, gate167inter1, gate167inter2, gate167inter3, gate167inter4, gate167inter5, gate167inter6, gate167inter7, gate167inter8, gate167inter9, gate167inter10, gate167inter11, gate167inter12, gate453inter0, gate453inter1, gate453inter2, gate453inter3, gate453inter4, gate453inter5, gate453inter6, gate453inter7, gate453inter8, gate453inter9, gate453inter10, gate453inter11, gate453inter12, gate123inter0, gate123inter1, gate123inter2, gate123inter3, gate123inter4, gate123inter5, gate123inter6, gate123inter7, gate123inter8, gate123inter9, gate123inter10, gate123inter11, gate123inter12, gate232inter0, gate232inter1, gate232inter2, gate232inter3, gate232inter4, gate232inter5, gate232inter6, gate232inter7, gate232inter8, gate232inter9, gate232inter10, gate232inter11, gate232inter12, gate272inter0, gate272inter1, gate272inter2, gate272inter3, gate272inter4, gate272inter5, gate272inter6, gate272inter7, gate272inter8, gate272inter9, gate272inter10, gate272inter11, gate272inter12, gate500inter0, gate500inter1, gate500inter2, gate500inter3, gate500inter4, gate500inter5, gate500inter6, gate500inter7, gate500inter8, gate500inter9, gate500inter10, gate500inter11, gate500inter12, gate488inter0, gate488inter1, gate488inter2, gate488inter3, gate488inter4, gate488inter5, gate488inter6, gate488inter7, gate488inter8, gate488inter9, gate488inter10, gate488inter11, gate488inter12, gate476inter0, gate476inter1, gate476inter2, gate476inter3, gate476inter4, gate476inter5, gate476inter6, gate476inter7, gate476inter8, gate476inter9, gate476inter10, gate476inter11, gate476inter12, gate99inter0, gate99inter1, gate99inter2, gate99inter3, gate99inter4, gate99inter5, gate99inter6, gate99inter7, gate99inter8, gate99inter9, gate99inter10, gate99inter11, gate99inter12, gate498inter0, gate498inter1, gate498inter2, gate498inter3, gate498inter4, gate498inter5, gate498inter6, gate498inter7, gate498inter8, gate498inter9, gate498inter10, gate498inter11, gate498inter12, gate196inter0, gate196inter1, gate196inter2, gate196inter3, gate196inter4, gate196inter5, gate196inter6, gate196inter7, gate196inter8, gate196inter9, gate196inter10, gate196inter11, gate196inter12, gate247inter0, gate247inter1, gate247inter2, gate247inter3, gate247inter4, gate247inter5, gate247inter6, gate247inter7, gate247inter8, gate247inter9, gate247inter10, gate247inter11, gate247inter12, gate79inter0, gate79inter1, gate79inter2, gate79inter3, gate79inter4, gate79inter5, gate79inter6, gate79inter7, gate79inter8, gate79inter9, gate79inter10, gate79inter11, gate79inter12, gate443inter0, gate443inter1, gate443inter2, gate443inter3, gate443inter4, gate443inter5, gate443inter6, gate443inter7, gate443inter8, gate443inter9, gate443inter10, gate443inter11, gate443inter12, gate244inter0, gate244inter1, gate244inter2, gate244inter3, gate244inter4, gate244inter5, gate244inter6, gate244inter7, gate244inter8, gate244inter9, gate244inter10, gate244inter11, gate244inter12, gate455inter0, gate455inter1, gate455inter2, gate455inter3, gate455inter4, gate455inter5, gate455inter6, gate455inter7, gate455inter8, gate455inter9, gate455inter10, gate455inter11, gate455inter12, gate95inter0, gate95inter1, gate95inter2, gate95inter3, gate95inter4, gate95inter5, gate95inter6, gate95inter7, gate95inter8, gate95inter9, gate95inter10, gate95inter11, gate95inter12, gate216inter0, gate216inter1, gate216inter2, gate216inter3, gate216inter4, gate216inter5, gate216inter6, gate216inter7, gate216inter8, gate216inter9, gate216inter10, gate216inter11, gate216inter12, gate164inter0, gate164inter1, gate164inter2, gate164inter3, gate164inter4, gate164inter5, gate164inter6, gate164inter7, gate164inter8, gate164inter9, gate164inter10, gate164inter11, gate164inter12, gate16inter0, gate16inter1, gate16inter2, gate16inter3, gate16inter4, gate16inter5, gate16inter6, gate16inter7, gate16inter8, gate16inter9, gate16inter10, gate16inter11, gate16inter12, gate194inter0, gate194inter1, gate194inter2, gate194inter3, gate194inter4, gate194inter5, gate194inter6, gate194inter7, gate194inter8, gate194inter9, gate194inter10, gate194inter11, gate194inter12, gate179inter0, gate179inter1, gate179inter2, gate179inter3, gate179inter4, gate179inter5, gate179inter6, gate179inter7, gate179inter8, gate179inter9, gate179inter10, gate179inter11, gate179inter12, gate211inter0, gate211inter1, gate211inter2, gate211inter3, gate211inter4, gate211inter5, gate211inter6, gate211inter7, gate211inter8, gate211inter9, gate211inter10, gate211inter11, gate211inter12, gate465inter0, gate465inter1, gate465inter2, gate465inter3, gate465inter4, gate465inter5, gate465inter6, gate465inter7, gate465inter8, gate465inter9, gate465inter10, gate465inter11, gate465inter12, gate130inter0, gate130inter1, gate130inter2, gate130inter3, gate130inter4, gate130inter5, gate130inter6, gate130inter7, gate130inter8, gate130inter9, gate130inter10, gate130inter11, gate130inter12, gate136inter0, gate136inter1, gate136inter2, gate136inter3, gate136inter4, gate136inter5, gate136inter6, gate136inter7, gate136inter8, gate136inter9, gate136inter10, gate136inter11, gate136inter12, gate44inter0, gate44inter1, gate44inter2, gate44inter3, gate44inter4, gate44inter5, gate44inter6, gate44inter7, gate44inter8, gate44inter9, gate44inter10, gate44inter11, gate44inter12, gate131inter0, gate131inter1, gate131inter2, gate131inter3, gate131inter4, gate131inter5, gate131inter6, gate131inter7, gate131inter8, gate131inter9, gate131inter10, gate131inter11, gate131inter12, gate115inter0, gate115inter1, gate115inter2, gate115inter3, gate115inter4, gate115inter5, gate115inter6, gate115inter7, gate115inter8, gate115inter9, gate115inter10, gate115inter11, gate115inter12, gate174inter0, gate174inter1, gate174inter2, gate174inter3, gate174inter4, gate174inter5, gate174inter6, gate174inter7, gate174inter8, gate174inter9, gate174inter10, gate174inter11, gate174inter12, gate52inter0, gate52inter1, gate52inter2, gate52inter3, gate52inter4, gate52inter5, gate52inter6, gate52inter7, gate52inter8, gate52inter9, gate52inter10, gate52inter11, gate52inter12, gate458inter0, gate458inter1, gate458inter2, gate458inter3, gate458inter4, gate458inter5, gate458inter6, gate458inter7, gate458inter8, gate458inter9, gate458inter10, gate458inter11, gate458inter12, gate214inter0, gate214inter1, gate214inter2, gate214inter3, gate214inter4, gate214inter5, gate214inter6, gate214inter7, gate214inter8, gate214inter9, gate214inter10, gate214inter11, gate214inter12, gate171inter0, gate171inter1, gate171inter2, gate171inter3, gate171inter4, gate171inter5, gate171inter6, gate171inter7, gate171inter8, gate171inter9, gate171inter10, gate171inter11, gate171inter12, gate388inter0, gate388inter1, gate388inter2, gate388inter3, gate388inter4, gate388inter5, gate388inter6, gate388inter7, gate388inter8, gate388inter9, gate388inter10, gate388inter11, gate388inter12, gate274inter0, gate274inter1, gate274inter2, gate274inter3, gate274inter4, gate274inter5, gate274inter6, gate274inter7, gate274inter8, gate274inter9, gate274inter10, gate274inter11, gate274inter12, gate412inter0, gate412inter1, gate412inter2, gate412inter3, gate412inter4, gate412inter5, gate412inter6, gate412inter7, gate412inter8, gate412inter9, gate412inter10, gate412inter11, gate412inter12, gate69inter0, gate69inter1, gate69inter2, gate69inter3, gate69inter4, gate69inter5, gate69inter6, gate69inter7, gate69inter8, gate69inter9, gate69inter10, gate69inter11, gate69inter12, gate163inter0, gate163inter1, gate163inter2, gate163inter3, gate163inter4, gate163inter5, gate163inter6, gate163inter7, gate163inter8, gate163inter9, gate163inter10, gate163inter11, gate163inter12, gate235inter0, gate235inter1, gate235inter2, gate235inter3, gate235inter4, gate235inter5, gate235inter6, gate235inter7, gate235inter8, gate235inter9, gate235inter10, gate235inter11, gate235inter12, gate234inter0, gate234inter1, gate234inter2, gate234inter3, gate234inter4, gate234inter5, gate234inter6, gate234inter7, gate234inter8, gate234inter9, gate234inter10, gate234inter11, gate234inter12, gate17inter0, gate17inter1, gate17inter2, gate17inter3, gate17inter4, gate17inter5, gate17inter6, gate17inter7, gate17inter8, gate17inter9, gate17inter10, gate17inter11, gate17inter12, gate60inter0, gate60inter1, gate60inter2, gate60inter3, gate60inter4, gate60inter5, gate60inter6, gate60inter7, gate60inter8, gate60inter9, gate60inter10, gate60inter11, gate60inter12, gate256inter0, gate256inter1, gate256inter2, gate256inter3, gate256inter4, gate256inter5, gate256inter6, gate256inter7, gate256inter8, gate256inter9, gate256inter10, gate256inter11, gate256inter12, gate127inter0, gate127inter1, gate127inter2, gate127inter3, gate127inter4, gate127inter5, gate127inter6, gate127inter7, gate127inter8, gate127inter9, gate127inter10, gate127inter11, gate127inter12, gate223inter0, gate223inter1, gate223inter2, gate223inter3, gate223inter4, gate223inter5, gate223inter6, gate223inter7, gate223inter8, gate223inter9, gate223inter10, gate223inter11, gate223inter12, gate158inter0, gate158inter1, gate158inter2, gate158inter3, gate158inter4, gate158inter5, gate158inter6, gate158inter7, gate158inter8, gate158inter9, gate158inter10, gate158inter11, gate158inter12, gate192inter0, gate192inter1, gate192inter2, gate192inter3, gate192inter4, gate192inter5, gate192inter6, gate192inter7, gate192inter8, gate192inter9, gate192inter10, gate192inter11, gate192inter12, gate59inter0, gate59inter1, gate59inter2, gate59inter3, gate59inter4, gate59inter5, gate59inter6, gate59inter7, gate59inter8, gate59inter9, gate59inter10, gate59inter11, gate59inter12, gate239inter0, gate239inter1, gate239inter2, gate239inter3, gate239inter4, gate239inter5, gate239inter6, gate239inter7, gate239inter8, gate239inter9, gate239inter10, gate239inter11, gate239inter12, gate195inter0, gate195inter1, gate195inter2, gate195inter3, gate195inter4, gate195inter5, gate195inter6, gate195inter7, gate195inter8, gate195inter9, gate195inter10, gate195inter11, gate195inter12, gate108inter0, gate108inter1, gate108inter2, gate108inter3, gate108inter4, gate108inter5, gate108inter6, gate108inter7, gate108inter8, gate108inter9, gate108inter10, gate108inter11, gate108inter12, gate170inter0, gate170inter1, gate170inter2, gate170inter3, gate170inter4, gate170inter5, gate170inter6, gate170inter7, gate170inter8, gate170inter9, gate170inter10, gate170inter11, gate170inter12, gate489inter0, gate489inter1, gate489inter2, gate489inter3, gate489inter4, gate489inter5, gate489inter6, gate489inter7, gate489inter8, gate489inter9, gate489inter10, gate489inter11, gate489inter12, gate126inter0, gate126inter1, gate126inter2, gate126inter3, gate126inter4, gate126inter5, gate126inter6, gate126inter7, gate126inter8, gate126inter9, gate126inter10, gate126inter11, gate126inter12, gate296inter0, gate296inter1, gate296inter2, gate296inter3, gate296inter4, gate296inter5, gate296inter6, gate296inter7, gate296inter8, gate296inter9, gate296inter10, gate296inter11, gate296inter12, gate491inter0, gate491inter1, gate491inter2, gate491inter3, gate491inter4, gate491inter5, gate491inter6, gate491inter7, gate491inter8, gate491inter9, gate491inter10, gate491inter11, gate491inter12, gate213inter0, gate213inter1, gate213inter2, gate213inter3, gate213inter4, gate213inter5, gate213inter6, gate213inter7, gate213inter8, gate213inter9, gate213inter10, gate213inter11, gate213inter12;



and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );
nand2 gate9( .a(G1), .b(G2), .O(G266) );
nand2 gate10( .a(G3), .b(G4), .O(G269) );
nand2 gate11( .a(G5), .b(G6), .O(G272) );
nand2 gate12( .a(G7), .b(G8), .O(G275) );
nand2 gate13( .a(G9), .b(G10), .O(G278) );
nand2 gate14( .a(G11), .b(G12), .O(G281) );

  xor2  gate1149(.a(G14), .b(G13), .O(gate15inter0));
  nand2 gate1150(.a(gate15inter0), .b(s_86), .O(gate15inter1));
  and2  gate1151(.a(G14), .b(G13), .O(gate15inter2));
  inv1  gate1152(.a(s_86), .O(gate15inter3));
  inv1  gate1153(.a(s_87), .O(gate15inter4));
  nand2 gate1154(.a(gate15inter4), .b(gate15inter3), .O(gate15inter5));
  nor2  gate1155(.a(gate15inter5), .b(gate15inter2), .O(gate15inter6));
  inv1  gate1156(.a(G13), .O(gate15inter7));
  inv1  gate1157(.a(G14), .O(gate15inter8));
  nand2 gate1158(.a(gate15inter8), .b(gate15inter7), .O(gate15inter9));
  nand2 gate1159(.a(s_87), .b(gate15inter3), .O(gate15inter10));
  nor2  gate1160(.a(gate15inter10), .b(gate15inter9), .O(gate15inter11));
  nor2  gate1161(.a(gate15inter11), .b(gate15inter6), .O(gate15inter12));
  nand2 gate1162(.a(gate15inter12), .b(gate15inter1), .O(G284));

  xor2  gate2675(.a(G16), .b(G15), .O(gate16inter0));
  nand2 gate2676(.a(gate16inter0), .b(s_304), .O(gate16inter1));
  and2  gate2677(.a(G16), .b(G15), .O(gate16inter2));
  inv1  gate2678(.a(s_304), .O(gate16inter3));
  inv1  gate2679(.a(s_305), .O(gate16inter4));
  nand2 gate2680(.a(gate16inter4), .b(gate16inter3), .O(gate16inter5));
  nor2  gate2681(.a(gate16inter5), .b(gate16inter2), .O(gate16inter6));
  inv1  gate2682(.a(G15), .O(gate16inter7));
  inv1  gate2683(.a(G16), .O(gate16inter8));
  nand2 gate2684(.a(gate16inter8), .b(gate16inter7), .O(gate16inter9));
  nand2 gate2685(.a(s_305), .b(gate16inter3), .O(gate16inter10));
  nor2  gate2686(.a(gate16inter10), .b(gate16inter9), .O(gate16inter11));
  nor2  gate2687(.a(gate16inter11), .b(gate16inter6), .O(gate16inter12));
  nand2 gate2688(.a(gate16inter12), .b(gate16inter1), .O(G287));

  xor2  gate2983(.a(G18), .b(G17), .O(gate17inter0));
  nand2 gate2984(.a(gate17inter0), .b(s_348), .O(gate17inter1));
  and2  gate2985(.a(G18), .b(G17), .O(gate17inter2));
  inv1  gate2986(.a(s_348), .O(gate17inter3));
  inv1  gate2987(.a(s_349), .O(gate17inter4));
  nand2 gate2988(.a(gate17inter4), .b(gate17inter3), .O(gate17inter5));
  nor2  gate2989(.a(gate17inter5), .b(gate17inter2), .O(gate17inter6));
  inv1  gate2990(.a(G17), .O(gate17inter7));
  inv1  gate2991(.a(G18), .O(gate17inter8));
  nand2 gate2992(.a(gate17inter8), .b(gate17inter7), .O(gate17inter9));
  nand2 gate2993(.a(s_349), .b(gate17inter3), .O(gate17inter10));
  nor2  gate2994(.a(gate17inter10), .b(gate17inter9), .O(gate17inter11));
  nor2  gate2995(.a(gate17inter11), .b(gate17inter6), .O(gate17inter12));
  nand2 gate2996(.a(gate17inter12), .b(gate17inter1), .O(G290));
nand2 gate18( .a(G19), .b(G20), .O(G293) );
nand2 gate19( .a(G21), .b(G22), .O(G296) );
nand2 gate20( .a(G23), .b(G24), .O(G299) );
nand2 gate21( .a(G25), .b(G26), .O(G302) );
nand2 gate22( .a(G27), .b(G28), .O(G305) );

  xor2  gate1009(.a(G30), .b(G29), .O(gate23inter0));
  nand2 gate1010(.a(gate23inter0), .b(s_66), .O(gate23inter1));
  and2  gate1011(.a(G30), .b(G29), .O(gate23inter2));
  inv1  gate1012(.a(s_66), .O(gate23inter3));
  inv1  gate1013(.a(s_67), .O(gate23inter4));
  nand2 gate1014(.a(gate23inter4), .b(gate23inter3), .O(gate23inter5));
  nor2  gate1015(.a(gate23inter5), .b(gate23inter2), .O(gate23inter6));
  inv1  gate1016(.a(G29), .O(gate23inter7));
  inv1  gate1017(.a(G30), .O(gate23inter8));
  nand2 gate1018(.a(gate23inter8), .b(gate23inter7), .O(gate23inter9));
  nand2 gate1019(.a(s_67), .b(gate23inter3), .O(gate23inter10));
  nor2  gate1020(.a(gate23inter10), .b(gate23inter9), .O(gate23inter11));
  nor2  gate1021(.a(gate23inter11), .b(gate23inter6), .O(gate23inter12));
  nand2 gate1022(.a(gate23inter12), .b(gate23inter1), .O(G308));
nand2 gate24( .a(G31), .b(G32), .O(G311) );

  xor2  gate2101(.a(G5), .b(G1), .O(gate25inter0));
  nand2 gate2102(.a(gate25inter0), .b(s_222), .O(gate25inter1));
  and2  gate2103(.a(G5), .b(G1), .O(gate25inter2));
  inv1  gate2104(.a(s_222), .O(gate25inter3));
  inv1  gate2105(.a(s_223), .O(gate25inter4));
  nand2 gate2106(.a(gate25inter4), .b(gate25inter3), .O(gate25inter5));
  nor2  gate2107(.a(gate25inter5), .b(gate25inter2), .O(gate25inter6));
  inv1  gate2108(.a(G1), .O(gate25inter7));
  inv1  gate2109(.a(G5), .O(gate25inter8));
  nand2 gate2110(.a(gate25inter8), .b(gate25inter7), .O(gate25inter9));
  nand2 gate2111(.a(s_223), .b(gate25inter3), .O(gate25inter10));
  nor2  gate2112(.a(gate25inter10), .b(gate25inter9), .O(gate25inter11));
  nor2  gate2113(.a(gate25inter11), .b(gate25inter6), .O(gate25inter12));
  nand2 gate2114(.a(gate25inter12), .b(gate25inter1), .O(G314));
nand2 gate26( .a(G9), .b(G13), .O(G317) );
nand2 gate27( .a(G2), .b(G6), .O(G320) );

  xor2  gate2227(.a(G14), .b(G10), .O(gate28inter0));
  nand2 gate2228(.a(gate28inter0), .b(s_240), .O(gate28inter1));
  and2  gate2229(.a(G14), .b(G10), .O(gate28inter2));
  inv1  gate2230(.a(s_240), .O(gate28inter3));
  inv1  gate2231(.a(s_241), .O(gate28inter4));
  nand2 gate2232(.a(gate28inter4), .b(gate28inter3), .O(gate28inter5));
  nor2  gate2233(.a(gate28inter5), .b(gate28inter2), .O(gate28inter6));
  inv1  gate2234(.a(G10), .O(gate28inter7));
  inv1  gate2235(.a(G14), .O(gate28inter8));
  nand2 gate2236(.a(gate28inter8), .b(gate28inter7), .O(gate28inter9));
  nand2 gate2237(.a(s_241), .b(gate28inter3), .O(gate28inter10));
  nor2  gate2238(.a(gate28inter10), .b(gate28inter9), .O(gate28inter11));
  nor2  gate2239(.a(gate28inter11), .b(gate28inter6), .O(gate28inter12));
  nand2 gate2240(.a(gate28inter12), .b(gate28inter1), .O(G323));
nand2 gate29( .a(G3), .b(G7), .O(G326) );
nand2 gate30( .a(G11), .b(G15), .O(G329) );
nand2 gate31( .a(G4), .b(G8), .O(G332) );
nand2 gate32( .a(G12), .b(G16), .O(G335) );
nand2 gate33( .a(G17), .b(G21), .O(G338) );

  xor2  gate2157(.a(G29), .b(G25), .O(gate34inter0));
  nand2 gate2158(.a(gate34inter0), .b(s_230), .O(gate34inter1));
  and2  gate2159(.a(G29), .b(G25), .O(gate34inter2));
  inv1  gate2160(.a(s_230), .O(gate34inter3));
  inv1  gate2161(.a(s_231), .O(gate34inter4));
  nand2 gate2162(.a(gate34inter4), .b(gate34inter3), .O(gate34inter5));
  nor2  gate2163(.a(gate34inter5), .b(gate34inter2), .O(gate34inter6));
  inv1  gate2164(.a(G25), .O(gate34inter7));
  inv1  gate2165(.a(G29), .O(gate34inter8));
  nand2 gate2166(.a(gate34inter8), .b(gate34inter7), .O(gate34inter9));
  nand2 gate2167(.a(s_231), .b(gate34inter3), .O(gate34inter10));
  nor2  gate2168(.a(gate34inter10), .b(gate34inter9), .O(gate34inter11));
  nor2  gate2169(.a(gate34inter11), .b(gate34inter6), .O(gate34inter12));
  nand2 gate2170(.a(gate34inter12), .b(gate34inter1), .O(G341));
nand2 gate35( .a(G18), .b(G22), .O(G344) );

  xor2  gate1569(.a(G30), .b(G26), .O(gate36inter0));
  nand2 gate1570(.a(gate36inter0), .b(s_146), .O(gate36inter1));
  and2  gate1571(.a(G30), .b(G26), .O(gate36inter2));
  inv1  gate1572(.a(s_146), .O(gate36inter3));
  inv1  gate1573(.a(s_147), .O(gate36inter4));
  nand2 gate1574(.a(gate36inter4), .b(gate36inter3), .O(gate36inter5));
  nor2  gate1575(.a(gate36inter5), .b(gate36inter2), .O(gate36inter6));
  inv1  gate1576(.a(G26), .O(gate36inter7));
  inv1  gate1577(.a(G30), .O(gate36inter8));
  nand2 gate1578(.a(gate36inter8), .b(gate36inter7), .O(gate36inter9));
  nand2 gate1579(.a(s_147), .b(gate36inter3), .O(gate36inter10));
  nor2  gate1580(.a(gate36inter10), .b(gate36inter9), .O(gate36inter11));
  nor2  gate1581(.a(gate36inter11), .b(gate36inter6), .O(gate36inter12));
  nand2 gate1582(.a(gate36inter12), .b(gate36inter1), .O(G347));
nand2 gate37( .a(G19), .b(G23), .O(G350) );
nand2 gate38( .a(G27), .b(G31), .O(G353) );

  xor2  gate2115(.a(G24), .b(G20), .O(gate39inter0));
  nand2 gate2116(.a(gate39inter0), .b(s_224), .O(gate39inter1));
  and2  gate2117(.a(G24), .b(G20), .O(gate39inter2));
  inv1  gate2118(.a(s_224), .O(gate39inter3));
  inv1  gate2119(.a(s_225), .O(gate39inter4));
  nand2 gate2120(.a(gate39inter4), .b(gate39inter3), .O(gate39inter5));
  nor2  gate2121(.a(gate39inter5), .b(gate39inter2), .O(gate39inter6));
  inv1  gate2122(.a(G20), .O(gate39inter7));
  inv1  gate2123(.a(G24), .O(gate39inter8));
  nand2 gate2124(.a(gate39inter8), .b(gate39inter7), .O(gate39inter9));
  nand2 gate2125(.a(s_225), .b(gate39inter3), .O(gate39inter10));
  nor2  gate2126(.a(gate39inter10), .b(gate39inter9), .O(gate39inter11));
  nor2  gate2127(.a(gate39inter11), .b(gate39inter6), .O(gate39inter12));
  nand2 gate2128(.a(gate39inter12), .b(gate39inter1), .O(G356));
nand2 gate40( .a(G28), .b(G32), .O(G359) );

  xor2  gate1261(.a(G266), .b(G1), .O(gate41inter0));
  nand2 gate1262(.a(gate41inter0), .b(s_102), .O(gate41inter1));
  and2  gate1263(.a(G266), .b(G1), .O(gate41inter2));
  inv1  gate1264(.a(s_102), .O(gate41inter3));
  inv1  gate1265(.a(s_103), .O(gate41inter4));
  nand2 gate1266(.a(gate41inter4), .b(gate41inter3), .O(gate41inter5));
  nor2  gate1267(.a(gate41inter5), .b(gate41inter2), .O(gate41inter6));
  inv1  gate1268(.a(G1), .O(gate41inter7));
  inv1  gate1269(.a(G266), .O(gate41inter8));
  nand2 gate1270(.a(gate41inter8), .b(gate41inter7), .O(gate41inter9));
  nand2 gate1271(.a(s_103), .b(gate41inter3), .O(gate41inter10));
  nor2  gate1272(.a(gate41inter10), .b(gate41inter9), .O(gate41inter11));
  nor2  gate1273(.a(gate41inter11), .b(gate41inter6), .O(gate41inter12));
  nand2 gate1274(.a(gate41inter12), .b(gate41inter1), .O(G362));

  xor2  gate1933(.a(G266), .b(G2), .O(gate42inter0));
  nand2 gate1934(.a(gate42inter0), .b(s_198), .O(gate42inter1));
  and2  gate1935(.a(G266), .b(G2), .O(gate42inter2));
  inv1  gate1936(.a(s_198), .O(gate42inter3));
  inv1  gate1937(.a(s_199), .O(gate42inter4));
  nand2 gate1938(.a(gate42inter4), .b(gate42inter3), .O(gate42inter5));
  nor2  gate1939(.a(gate42inter5), .b(gate42inter2), .O(gate42inter6));
  inv1  gate1940(.a(G2), .O(gate42inter7));
  inv1  gate1941(.a(G266), .O(gate42inter8));
  nand2 gate1942(.a(gate42inter8), .b(gate42inter7), .O(gate42inter9));
  nand2 gate1943(.a(s_199), .b(gate42inter3), .O(gate42inter10));
  nor2  gate1944(.a(gate42inter10), .b(gate42inter9), .O(gate42inter11));
  nor2  gate1945(.a(gate42inter11), .b(gate42inter6), .O(gate42inter12));
  nand2 gate1946(.a(gate42inter12), .b(gate42inter1), .O(G363));

  xor2  gate1877(.a(G269), .b(G3), .O(gate43inter0));
  nand2 gate1878(.a(gate43inter0), .b(s_190), .O(gate43inter1));
  and2  gate1879(.a(G269), .b(G3), .O(gate43inter2));
  inv1  gate1880(.a(s_190), .O(gate43inter3));
  inv1  gate1881(.a(s_191), .O(gate43inter4));
  nand2 gate1882(.a(gate43inter4), .b(gate43inter3), .O(gate43inter5));
  nor2  gate1883(.a(gate43inter5), .b(gate43inter2), .O(gate43inter6));
  inv1  gate1884(.a(G3), .O(gate43inter7));
  inv1  gate1885(.a(G269), .O(gate43inter8));
  nand2 gate1886(.a(gate43inter8), .b(gate43inter7), .O(gate43inter9));
  nand2 gate1887(.a(s_191), .b(gate43inter3), .O(gate43inter10));
  nor2  gate1888(.a(gate43inter10), .b(gate43inter9), .O(gate43inter11));
  nor2  gate1889(.a(gate43inter11), .b(gate43inter6), .O(gate43inter12));
  nand2 gate1890(.a(gate43inter12), .b(gate43inter1), .O(G364));

  xor2  gate2773(.a(G269), .b(G4), .O(gate44inter0));
  nand2 gate2774(.a(gate44inter0), .b(s_318), .O(gate44inter1));
  and2  gate2775(.a(G269), .b(G4), .O(gate44inter2));
  inv1  gate2776(.a(s_318), .O(gate44inter3));
  inv1  gate2777(.a(s_319), .O(gate44inter4));
  nand2 gate2778(.a(gate44inter4), .b(gate44inter3), .O(gate44inter5));
  nor2  gate2779(.a(gate44inter5), .b(gate44inter2), .O(gate44inter6));
  inv1  gate2780(.a(G4), .O(gate44inter7));
  inv1  gate2781(.a(G269), .O(gate44inter8));
  nand2 gate2782(.a(gate44inter8), .b(gate44inter7), .O(gate44inter9));
  nand2 gate2783(.a(s_319), .b(gate44inter3), .O(gate44inter10));
  nor2  gate2784(.a(gate44inter10), .b(gate44inter9), .O(gate44inter11));
  nor2  gate2785(.a(gate44inter11), .b(gate44inter6), .O(gate44inter12));
  nand2 gate2786(.a(gate44inter12), .b(gate44inter1), .O(G365));
nand2 gate45( .a(G5), .b(G272), .O(G366) );

  xor2  gate1919(.a(G272), .b(G6), .O(gate46inter0));
  nand2 gate1920(.a(gate46inter0), .b(s_196), .O(gate46inter1));
  and2  gate1921(.a(G272), .b(G6), .O(gate46inter2));
  inv1  gate1922(.a(s_196), .O(gate46inter3));
  inv1  gate1923(.a(s_197), .O(gate46inter4));
  nand2 gate1924(.a(gate46inter4), .b(gate46inter3), .O(gate46inter5));
  nor2  gate1925(.a(gate46inter5), .b(gate46inter2), .O(gate46inter6));
  inv1  gate1926(.a(G6), .O(gate46inter7));
  inv1  gate1927(.a(G272), .O(gate46inter8));
  nand2 gate1928(.a(gate46inter8), .b(gate46inter7), .O(gate46inter9));
  nand2 gate1929(.a(s_197), .b(gate46inter3), .O(gate46inter10));
  nor2  gate1930(.a(gate46inter10), .b(gate46inter9), .O(gate46inter11));
  nor2  gate1931(.a(gate46inter11), .b(gate46inter6), .O(gate46inter12));
  nand2 gate1932(.a(gate46inter12), .b(gate46inter1), .O(G367));

  xor2  gate2255(.a(G275), .b(G7), .O(gate47inter0));
  nand2 gate2256(.a(gate47inter0), .b(s_244), .O(gate47inter1));
  and2  gate2257(.a(G275), .b(G7), .O(gate47inter2));
  inv1  gate2258(.a(s_244), .O(gate47inter3));
  inv1  gate2259(.a(s_245), .O(gate47inter4));
  nand2 gate2260(.a(gate47inter4), .b(gate47inter3), .O(gate47inter5));
  nor2  gate2261(.a(gate47inter5), .b(gate47inter2), .O(gate47inter6));
  inv1  gate2262(.a(G7), .O(gate47inter7));
  inv1  gate2263(.a(G275), .O(gate47inter8));
  nand2 gate2264(.a(gate47inter8), .b(gate47inter7), .O(gate47inter9));
  nand2 gate2265(.a(s_245), .b(gate47inter3), .O(gate47inter10));
  nor2  gate2266(.a(gate47inter10), .b(gate47inter9), .O(gate47inter11));
  nor2  gate2267(.a(gate47inter11), .b(gate47inter6), .O(gate47inter12));
  nand2 gate2268(.a(gate47inter12), .b(gate47inter1), .O(G368));

  xor2  gate1597(.a(G275), .b(G8), .O(gate48inter0));
  nand2 gate1598(.a(gate48inter0), .b(s_150), .O(gate48inter1));
  and2  gate1599(.a(G275), .b(G8), .O(gate48inter2));
  inv1  gate1600(.a(s_150), .O(gate48inter3));
  inv1  gate1601(.a(s_151), .O(gate48inter4));
  nand2 gate1602(.a(gate48inter4), .b(gate48inter3), .O(gate48inter5));
  nor2  gate1603(.a(gate48inter5), .b(gate48inter2), .O(gate48inter6));
  inv1  gate1604(.a(G8), .O(gate48inter7));
  inv1  gate1605(.a(G275), .O(gate48inter8));
  nand2 gate1606(.a(gate48inter8), .b(gate48inter7), .O(gate48inter9));
  nand2 gate1607(.a(s_151), .b(gate48inter3), .O(gate48inter10));
  nor2  gate1608(.a(gate48inter10), .b(gate48inter9), .O(gate48inter11));
  nor2  gate1609(.a(gate48inter11), .b(gate48inter6), .O(gate48inter12));
  nand2 gate1610(.a(gate48inter12), .b(gate48inter1), .O(G369));
nand2 gate49( .a(G9), .b(G278), .O(G370) );

  xor2  gate2171(.a(G278), .b(G10), .O(gate50inter0));
  nand2 gate2172(.a(gate50inter0), .b(s_232), .O(gate50inter1));
  and2  gate2173(.a(G278), .b(G10), .O(gate50inter2));
  inv1  gate2174(.a(s_232), .O(gate50inter3));
  inv1  gate2175(.a(s_233), .O(gate50inter4));
  nand2 gate2176(.a(gate50inter4), .b(gate50inter3), .O(gate50inter5));
  nor2  gate2177(.a(gate50inter5), .b(gate50inter2), .O(gate50inter6));
  inv1  gate2178(.a(G10), .O(gate50inter7));
  inv1  gate2179(.a(G278), .O(gate50inter8));
  nand2 gate2180(.a(gate50inter8), .b(gate50inter7), .O(gate50inter9));
  nand2 gate2181(.a(s_233), .b(gate50inter3), .O(gate50inter10));
  nor2  gate2182(.a(gate50inter10), .b(gate50inter9), .O(gate50inter11));
  nor2  gate2183(.a(gate50inter11), .b(gate50inter6), .O(gate50inter12));
  nand2 gate2184(.a(gate50inter12), .b(gate50inter1), .O(G371));
nand2 gate51( .a(G11), .b(G281), .O(G372) );

  xor2  gate2829(.a(G281), .b(G12), .O(gate52inter0));
  nand2 gate2830(.a(gate52inter0), .b(s_326), .O(gate52inter1));
  and2  gate2831(.a(G281), .b(G12), .O(gate52inter2));
  inv1  gate2832(.a(s_326), .O(gate52inter3));
  inv1  gate2833(.a(s_327), .O(gate52inter4));
  nand2 gate2834(.a(gate52inter4), .b(gate52inter3), .O(gate52inter5));
  nor2  gate2835(.a(gate52inter5), .b(gate52inter2), .O(gate52inter6));
  inv1  gate2836(.a(G12), .O(gate52inter7));
  inv1  gate2837(.a(G281), .O(gate52inter8));
  nand2 gate2838(.a(gate52inter8), .b(gate52inter7), .O(gate52inter9));
  nand2 gate2839(.a(s_327), .b(gate52inter3), .O(gate52inter10));
  nor2  gate2840(.a(gate52inter10), .b(gate52inter9), .O(gate52inter11));
  nor2  gate2841(.a(gate52inter11), .b(gate52inter6), .O(gate52inter12));
  nand2 gate2842(.a(gate52inter12), .b(gate52inter1), .O(G373));
nand2 gate53( .a(G13), .b(G284), .O(G374) );

  xor2  gate1527(.a(G284), .b(G14), .O(gate54inter0));
  nand2 gate1528(.a(gate54inter0), .b(s_140), .O(gate54inter1));
  and2  gate1529(.a(G284), .b(G14), .O(gate54inter2));
  inv1  gate1530(.a(s_140), .O(gate54inter3));
  inv1  gate1531(.a(s_141), .O(gate54inter4));
  nand2 gate1532(.a(gate54inter4), .b(gate54inter3), .O(gate54inter5));
  nor2  gate1533(.a(gate54inter5), .b(gate54inter2), .O(gate54inter6));
  inv1  gate1534(.a(G14), .O(gate54inter7));
  inv1  gate1535(.a(G284), .O(gate54inter8));
  nand2 gate1536(.a(gate54inter8), .b(gate54inter7), .O(gate54inter9));
  nand2 gate1537(.a(s_141), .b(gate54inter3), .O(gate54inter10));
  nor2  gate1538(.a(gate54inter10), .b(gate54inter9), .O(gate54inter11));
  nor2  gate1539(.a(gate54inter11), .b(gate54inter6), .O(gate54inter12));
  nand2 gate1540(.a(gate54inter12), .b(gate54inter1), .O(G375));
nand2 gate55( .a(G15), .b(G287), .O(G376) );
nand2 gate56( .a(G16), .b(G287), .O(G377) );
nand2 gate57( .a(G17), .b(G290), .O(G378) );
nand2 gate58( .a(G18), .b(G290), .O(G379) );

  xor2  gate3081(.a(G293), .b(G19), .O(gate59inter0));
  nand2 gate3082(.a(gate59inter0), .b(s_362), .O(gate59inter1));
  and2  gate3083(.a(G293), .b(G19), .O(gate59inter2));
  inv1  gate3084(.a(s_362), .O(gate59inter3));
  inv1  gate3085(.a(s_363), .O(gate59inter4));
  nand2 gate3086(.a(gate59inter4), .b(gate59inter3), .O(gate59inter5));
  nor2  gate3087(.a(gate59inter5), .b(gate59inter2), .O(gate59inter6));
  inv1  gate3088(.a(G19), .O(gate59inter7));
  inv1  gate3089(.a(G293), .O(gate59inter8));
  nand2 gate3090(.a(gate59inter8), .b(gate59inter7), .O(gate59inter9));
  nand2 gate3091(.a(s_363), .b(gate59inter3), .O(gate59inter10));
  nor2  gate3092(.a(gate59inter10), .b(gate59inter9), .O(gate59inter11));
  nor2  gate3093(.a(gate59inter11), .b(gate59inter6), .O(gate59inter12));
  nand2 gate3094(.a(gate59inter12), .b(gate59inter1), .O(G380));

  xor2  gate2997(.a(G293), .b(G20), .O(gate60inter0));
  nand2 gate2998(.a(gate60inter0), .b(s_350), .O(gate60inter1));
  and2  gate2999(.a(G293), .b(G20), .O(gate60inter2));
  inv1  gate3000(.a(s_350), .O(gate60inter3));
  inv1  gate3001(.a(s_351), .O(gate60inter4));
  nand2 gate3002(.a(gate60inter4), .b(gate60inter3), .O(gate60inter5));
  nor2  gate3003(.a(gate60inter5), .b(gate60inter2), .O(gate60inter6));
  inv1  gate3004(.a(G20), .O(gate60inter7));
  inv1  gate3005(.a(G293), .O(gate60inter8));
  nand2 gate3006(.a(gate60inter8), .b(gate60inter7), .O(gate60inter9));
  nand2 gate3007(.a(s_351), .b(gate60inter3), .O(gate60inter10));
  nor2  gate3008(.a(gate60inter10), .b(gate60inter9), .O(gate60inter11));
  nor2  gate3009(.a(gate60inter11), .b(gate60inter6), .O(gate60inter12));
  nand2 gate3010(.a(gate60inter12), .b(gate60inter1), .O(G381));

  xor2  gate1177(.a(G296), .b(G21), .O(gate61inter0));
  nand2 gate1178(.a(gate61inter0), .b(s_90), .O(gate61inter1));
  and2  gate1179(.a(G296), .b(G21), .O(gate61inter2));
  inv1  gate1180(.a(s_90), .O(gate61inter3));
  inv1  gate1181(.a(s_91), .O(gate61inter4));
  nand2 gate1182(.a(gate61inter4), .b(gate61inter3), .O(gate61inter5));
  nor2  gate1183(.a(gate61inter5), .b(gate61inter2), .O(gate61inter6));
  inv1  gate1184(.a(G21), .O(gate61inter7));
  inv1  gate1185(.a(G296), .O(gate61inter8));
  nand2 gate1186(.a(gate61inter8), .b(gate61inter7), .O(gate61inter9));
  nand2 gate1187(.a(s_91), .b(gate61inter3), .O(gate61inter10));
  nor2  gate1188(.a(gate61inter10), .b(gate61inter9), .O(gate61inter11));
  nor2  gate1189(.a(gate61inter11), .b(gate61inter6), .O(gate61inter12));
  nand2 gate1190(.a(gate61inter12), .b(gate61inter1), .O(G382));
nand2 gate62( .a(G22), .b(G296), .O(G383) );

  xor2  gate2059(.a(G299), .b(G23), .O(gate63inter0));
  nand2 gate2060(.a(gate63inter0), .b(s_216), .O(gate63inter1));
  and2  gate2061(.a(G299), .b(G23), .O(gate63inter2));
  inv1  gate2062(.a(s_216), .O(gate63inter3));
  inv1  gate2063(.a(s_217), .O(gate63inter4));
  nand2 gate2064(.a(gate63inter4), .b(gate63inter3), .O(gate63inter5));
  nor2  gate2065(.a(gate63inter5), .b(gate63inter2), .O(gate63inter6));
  inv1  gate2066(.a(G23), .O(gate63inter7));
  inv1  gate2067(.a(G299), .O(gate63inter8));
  nand2 gate2068(.a(gate63inter8), .b(gate63inter7), .O(gate63inter9));
  nand2 gate2069(.a(s_217), .b(gate63inter3), .O(gate63inter10));
  nor2  gate2070(.a(gate63inter10), .b(gate63inter9), .O(gate63inter11));
  nor2  gate2071(.a(gate63inter11), .b(gate63inter6), .O(gate63inter12));
  nand2 gate2072(.a(gate63inter12), .b(gate63inter1), .O(G384));

  xor2  gate1947(.a(G299), .b(G24), .O(gate64inter0));
  nand2 gate1948(.a(gate64inter0), .b(s_200), .O(gate64inter1));
  and2  gate1949(.a(G299), .b(G24), .O(gate64inter2));
  inv1  gate1950(.a(s_200), .O(gate64inter3));
  inv1  gate1951(.a(s_201), .O(gate64inter4));
  nand2 gate1952(.a(gate64inter4), .b(gate64inter3), .O(gate64inter5));
  nor2  gate1953(.a(gate64inter5), .b(gate64inter2), .O(gate64inter6));
  inv1  gate1954(.a(G24), .O(gate64inter7));
  inv1  gate1955(.a(G299), .O(gate64inter8));
  nand2 gate1956(.a(gate64inter8), .b(gate64inter7), .O(gate64inter9));
  nand2 gate1957(.a(s_201), .b(gate64inter3), .O(gate64inter10));
  nor2  gate1958(.a(gate64inter10), .b(gate64inter9), .O(gate64inter11));
  nor2  gate1959(.a(gate64inter11), .b(gate64inter6), .O(gate64inter12));
  nand2 gate1960(.a(gate64inter12), .b(gate64inter1), .O(G385));
nand2 gate65( .a(G25), .b(G302), .O(G386) );
nand2 gate66( .a(G26), .b(G302), .O(G387) );
nand2 gate67( .a(G27), .b(G305), .O(G388) );
nand2 gate68( .a(G28), .b(G305), .O(G389) );

  xor2  gate2927(.a(G308), .b(G29), .O(gate69inter0));
  nand2 gate2928(.a(gate69inter0), .b(s_340), .O(gate69inter1));
  and2  gate2929(.a(G308), .b(G29), .O(gate69inter2));
  inv1  gate2930(.a(s_340), .O(gate69inter3));
  inv1  gate2931(.a(s_341), .O(gate69inter4));
  nand2 gate2932(.a(gate69inter4), .b(gate69inter3), .O(gate69inter5));
  nor2  gate2933(.a(gate69inter5), .b(gate69inter2), .O(gate69inter6));
  inv1  gate2934(.a(G29), .O(gate69inter7));
  inv1  gate2935(.a(G308), .O(gate69inter8));
  nand2 gate2936(.a(gate69inter8), .b(gate69inter7), .O(gate69inter9));
  nand2 gate2937(.a(s_341), .b(gate69inter3), .O(gate69inter10));
  nor2  gate2938(.a(gate69inter10), .b(gate69inter9), .O(gate69inter11));
  nor2  gate2939(.a(gate69inter11), .b(gate69inter6), .O(gate69inter12));
  nand2 gate2940(.a(gate69inter12), .b(gate69inter1), .O(G390));
nand2 gate70( .a(G30), .b(G308), .O(G391) );
nand2 gate71( .a(G31), .b(G311), .O(G392) );
nand2 gate72( .a(G32), .b(G311), .O(G393) );

  xor2  gate2241(.a(G314), .b(G1), .O(gate73inter0));
  nand2 gate2242(.a(gate73inter0), .b(s_242), .O(gate73inter1));
  and2  gate2243(.a(G314), .b(G1), .O(gate73inter2));
  inv1  gate2244(.a(s_242), .O(gate73inter3));
  inv1  gate2245(.a(s_243), .O(gate73inter4));
  nand2 gate2246(.a(gate73inter4), .b(gate73inter3), .O(gate73inter5));
  nor2  gate2247(.a(gate73inter5), .b(gate73inter2), .O(gate73inter6));
  inv1  gate2248(.a(G1), .O(gate73inter7));
  inv1  gate2249(.a(G314), .O(gate73inter8));
  nand2 gate2250(.a(gate73inter8), .b(gate73inter7), .O(gate73inter9));
  nand2 gate2251(.a(s_243), .b(gate73inter3), .O(gate73inter10));
  nor2  gate2252(.a(gate73inter10), .b(gate73inter9), .O(gate73inter11));
  nor2  gate2253(.a(gate73inter11), .b(gate73inter6), .O(gate73inter12));
  nand2 gate2254(.a(gate73inter12), .b(gate73inter1), .O(G394));
nand2 gate74( .a(G5), .b(G314), .O(G395) );

  xor2  gate841(.a(G317), .b(G9), .O(gate75inter0));
  nand2 gate842(.a(gate75inter0), .b(s_42), .O(gate75inter1));
  and2  gate843(.a(G317), .b(G9), .O(gate75inter2));
  inv1  gate844(.a(s_42), .O(gate75inter3));
  inv1  gate845(.a(s_43), .O(gate75inter4));
  nand2 gate846(.a(gate75inter4), .b(gate75inter3), .O(gate75inter5));
  nor2  gate847(.a(gate75inter5), .b(gate75inter2), .O(gate75inter6));
  inv1  gate848(.a(G9), .O(gate75inter7));
  inv1  gate849(.a(G317), .O(gate75inter8));
  nand2 gate850(.a(gate75inter8), .b(gate75inter7), .O(gate75inter9));
  nand2 gate851(.a(s_43), .b(gate75inter3), .O(gate75inter10));
  nor2  gate852(.a(gate75inter10), .b(gate75inter9), .O(gate75inter11));
  nor2  gate853(.a(gate75inter11), .b(gate75inter6), .O(gate75inter12));
  nand2 gate854(.a(gate75inter12), .b(gate75inter1), .O(G396));
nand2 gate76( .a(G13), .b(G317), .O(G397) );
nand2 gate77( .a(G2), .b(G320), .O(G398) );
nand2 gate78( .a(G6), .b(G320), .O(G399) );

  xor2  gate2577(.a(G323), .b(G10), .O(gate79inter0));
  nand2 gate2578(.a(gate79inter0), .b(s_290), .O(gate79inter1));
  and2  gate2579(.a(G323), .b(G10), .O(gate79inter2));
  inv1  gate2580(.a(s_290), .O(gate79inter3));
  inv1  gate2581(.a(s_291), .O(gate79inter4));
  nand2 gate2582(.a(gate79inter4), .b(gate79inter3), .O(gate79inter5));
  nor2  gate2583(.a(gate79inter5), .b(gate79inter2), .O(gate79inter6));
  inv1  gate2584(.a(G10), .O(gate79inter7));
  inv1  gate2585(.a(G323), .O(gate79inter8));
  nand2 gate2586(.a(gate79inter8), .b(gate79inter7), .O(gate79inter9));
  nand2 gate2587(.a(s_291), .b(gate79inter3), .O(gate79inter10));
  nor2  gate2588(.a(gate79inter10), .b(gate79inter9), .O(gate79inter11));
  nor2  gate2589(.a(gate79inter11), .b(gate79inter6), .O(gate79inter12));
  nand2 gate2590(.a(gate79inter12), .b(gate79inter1), .O(G400));
nand2 gate80( .a(G14), .b(G323), .O(G401) );
nand2 gate81( .a(G3), .b(G326), .O(G402) );

  xor2  gate981(.a(G326), .b(G7), .O(gate82inter0));
  nand2 gate982(.a(gate82inter0), .b(s_62), .O(gate82inter1));
  and2  gate983(.a(G326), .b(G7), .O(gate82inter2));
  inv1  gate984(.a(s_62), .O(gate82inter3));
  inv1  gate985(.a(s_63), .O(gate82inter4));
  nand2 gate986(.a(gate82inter4), .b(gate82inter3), .O(gate82inter5));
  nor2  gate987(.a(gate82inter5), .b(gate82inter2), .O(gate82inter6));
  inv1  gate988(.a(G7), .O(gate82inter7));
  inv1  gate989(.a(G326), .O(gate82inter8));
  nand2 gate990(.a(gate82inter8), .b(gate82inter7), .O(gate82inter9));
  nand2 gate991(.a(s_63), .b(gate82inter3), .O(gate82inter10));
  nor2  gate992(.a(gate82inter10), .b(gate82inter9), .O(gate82inter11));
  nor2  gate993(.a(gate82inter11), .b(gate82inter6), .O(gate82inter12));
  nand2 gate994(.a(gate82inter12), .b(gate82inter1), .O(G403));

  xor2  gate911(.a(G329), .b(G11), .O(gate83inter0));
  nand2 gate912(.a(gate83inter0), .b(s_52), .O(gate83inter1));
  and2  gate913(.a(G329), .b(G11), .O(gate83inter2));
  inv1  gate914(.a(s_52), .O(gate83inter3));
  inv1  gate915(.a(s_53), .O(gate83inter4));
  nand2 gate916(.a(gate83inter4), .b(gate83inter3), .O(gate83inter5));
  nor2  gate917(.a(gate83inter5), .b(gate83inter2), .O(gate83inter6));
  inv1  gate918(.a(G11), .O(gate83inter7));
  inv1  gate919(.a(G329), .O(gate83inter8));
  nand2 gate920(.a(gate83inter8), .b(gate83inter7), .O(gate83inter9));
  nand2 gate921(.a(s_53), .b(gate83inter3), .O(gate83inter10));
  nor2  gate922(.a(gate83inter10), .b(gate83inter9), .O(gate83inter11));
  nor2  gate923(.a(gate83inter11), .b(gate83inter6), .O(gate83inter12));
  nand2 gate924(.a(gate83inter12), .b(gate83inter1), .O(G404));

  xor2  gate603(.a(G329), .b(G15), .O(gate84inter0));
  nand2 gate604(.a(gate84inter0), .b(s_8), .O(gate84inter1));
  and2  gate605(.a(G329), .b(G15), .O(gate84inter2));
  inv1  gate606(.a(s_8), .O(gate84inter3));
  inv1  gate607(.a(s_9), .O(gate84inter4));
  nand2 gate608(.a(gate84inter4), .b(gate84inter3), .O(gate84inter5));
  nor2  gate609(.a(gate84inter5), .b(gate84inter2), .O(gate84inter6));
  inv1  gate610(.a(G15), .O(gate84inter7));
  inv1  gate611(.a(G329), .O(gate84inter8));
  nand2 gate612(.a(gate84inter8), .b(gate84inter7), .O(gate84inter9));
  nand2 gate613(.a(s_9), .b(gate84inter3), .O(gate84inter10));
  nor2  gate614(.a(gate84inter10), .b(gate84inter9), .O(gate84inter11));
  nor2  gate615(.a(gate84inter11), .b(gate84inter6), .O(gate84inter12));
  nand2 gate616(.a(gate84inter12), .b(gate84inter1), .O(G405));

  xor2  gate575(.a(G332), .b(G4), .O(gate85inter0));
  nand2 gate576(.a(gate85inter0), .b(s_4), .O(gate85inter1));
  and2  gate577(.a(G332), .b(G4), .O(gate85inter2));
  inv1  gate578(.a(s_4), .O(gate85inter3));
  inv1  gate579(.a(s_5), .O(gate85inter4));
  nand2 gate580(.a(gate85inter4), .b(gate85inter3), .O(gate85inter5));
  nor2  gate581(.a(gate85inter5), .b(gate85inter2), .O(gate85inter6));
  inv1  gate582(.a(G4), .O(gate85inter7));
  inv1  gate583(.a(G332), .O(gate85inter8));
  nand2 gate584(.a(gate85inter8), .b(gate85inter7), .O(gate85inter9));
  nand2 gate585(.a(s_5), .b(gate85inter3), .O(gate85inter10));
  nor2  gate586(.a(gate85inter10), .b(gate85inter9), .O(gate85inter11));
  nor2  gate587(.a(gate85inter11), .b(gate85inter6), .O(gate85inter12));
  nand2 gate588(.a(gate85inter12), .b(gate85inter1), .O(G406));

  xor2  gate925(.a(G332), .b(G8), .O(gate86inter0));
  nand2 gate926(.a(gate86inter0), .b(s_54), .O(gate86inter1));
  and2  gate927(.a(G332), .b(G8), .O(gate86inter2));
  inv1  gate928(.a(s_54), .O(gate86inter3));
  inv1  gate929(.a(s_55), .O(gate86inter4));
  nand2 gate930(.a(gate86inter4), .b(gate86inter3), .O(gate86inter5));
  nor2  gate931(.a(gate86inter5), .b(gate86inter2), .O(gate86inter6));
  inv1  gate932(.a(G8), .O(gate86inter7));
  inv1  gate933(.a(G332), .O(gate86inter8));
  nand2 gate934(.a(gate86inter8), .b(gate86inter7), .O(gate86inter9));
  nand2 gate935(.a(s_55), .b(gate86inter3), .O(gate86inter10));
  nor2  gate936(.a(gate86inter10), .b(gate86inter9), .O(gate86inter11));
  nor2  gate937(.a(gate86inter11), .b(gate86inter6), .O(gate86inter12));
  nand2 gate938(.a(gate86inter12), .b(gate86inter1), .O(G407));
nand2 gate87( .a(G12), .b(G335), .O(G408) );

  xor2  gate1303(.a(G335), .b(G16), .O(gate88inter0));
  nand2 gate1304(.a(gate88inter0), .b(s_108), .O(gate88inter1));
  and2  gate1305(.a(G335), .b(G16), .O(gate88inter2));
  inv1  gate1306(.a(s_108), .O(gate88inter3));
  inv1  gate1307(.a(s_109), .O(gate88inter4));
  nand2 gate1308(.a(gate88inter4), .b(gate88inter3), .O(gate88inter5));
  nor2  gate1309(.a(gate88inter5), .b(gate88inter2), .O(gate88inter6));
  inv1  gate1310(.a(G16), .O(gate88inter7));
  inv1  gate1311(.a(G335), .O(gate88inter8));
  nand2 gate1312(.a(gate88inter8), .b(gate88inter7), .O(gate88inter9));
  nand2 gate1313(.a(s_109), .b(gate88inter3), .O(gate88inter10));
  nor2  gate1314(.a(gate88inter10), .b(gate88inter9), .O(gate88inter11));
  nor2  gate1315(.a(gate88inter11), .b(gate88inter6), .O(gate88inter12));
  nand2 gate1316(.a(gate88inter12), .b(gate88inter1), .O(G409));
nand2 gate89( .a(G17), .b(G338), .O(G410) );

  xor2  gate1667(.a(G338), .b(G21), .O(gate90inter0));
  nand2 gate1668(.a(gate90inter0), .b(s_160), .O(gate90inter1));
  and2  gate1669(.a(G338), .b(G21), .O(gate90inter2));
  inv1  gate1670(.a(s_160), .O(gate90inter3));
  inv1  gate1671(.a(s_161), .O(gate90inter4));
  nand2 gate1672(.a(gate90inter4), .b(gate90inter3), .O(gate90inter5));
  nor2  gate1673(.a(gate90inter5), .b(gate90inter2), .O(gate90inter6));
  inv1  gate1674(.a(G21), .O(gate90inter7));
  inv1  gate1675(.a(G338), .O(gate90inter8));
  nand2 gate1676(.a(gate90inter8), .b(gate90inter7), .O(gate90inter9));
  nand2 gate1677(.a(s_161), .b(gate90inter3), .O(gate90inter10));
  nor2  gate1678(.a(gate90inter10), .b(gate90inter9), .O(gate90inter11));
  nor2  gate1679(.a(gate90inter11), .b(gate90inter6), .O(gate90inter12));
  nand2 gate1680(.a(gate90inter12), .b(gate90inter1), .O(G411));
nand2 gate91( .a(G25), .b(G341), .O(G412) );
nand2 gate92( .a(G29), .b(G341), .O(G413) );
nand2 gate93( .a(G18), .b(G344), .O(G414) );

  xor2  gate1681(.a(G344), .b(G22), .O(gate94inter0));
  nand2 gate1682(.a(gate94inter0), .b(s_162), .O(gate94inter1));
  and2  gate1683(.a(G344), .b(G22), .O(gate94inter2));
  inv1  gate1684(.a(s_162), .O(gate94inter3));
  inv1  gate1685(.a(s_163), .O(gate94inter4));
  nand2 gate1686(.a(gate94inter4), .b(gate94inter3), .O(gate94inter5));
  nor2  gate1687(.a(gate94inter5), .b(gate94inter2), .O(gate94inter6));
  inv1  gate1688(.a(G22), .O(gate94inter7));
  inv1  gate1689(.a(G344), .O(gate94inter8));
  nand2 gate1690(.a(gate94inter8), .b(gate94inter7), .O(gate94inter9));
  nand2 gate1691(.a(s_163), .b(gate94inter3), .O(gate94inter10));
  nor2  gate1692(.a(gate94inter10), .b(gate94inter9), .O(gate94inter11));
  nor2  gate1693(.a(gate94inter11), .b(gate94inter6), .O(gate94inter12));
  nand2 gate1694(.a(gate94inter12), .b(gate94inter1), .O(G415));

  xor2  gate2633(.a(G347), .b(G26), .O(gate95inter0));
  nand2 gate2634(.a(gate95inter0), .b(s_298), .O(gate95inter1));
  and2  gate2635(.a(G347), .b(G26), .O(gate95inter2));
  inv1  gate2636(.a(s_298), .O(gate95inter3));
  inv1  gate2637(.a(s_299), .O(gate95inter4));
  nand2 gate2638(.a(gate95inter4), .b(gate95inter3), .O(gate95inter5));
  nor2  gate2639(.a(gate95inter5), .b(gate95inter2), .O(gate95inter6));
  inv1  gate2640(.a(G26), .O(gate95inter7));
  inv1  gate2641(.a(G347), .O(gate95inter8));
  nand2 gate2642(.a(gate95inter8), .b(gate95inter7), .O(gate95inter9));
  nand2 gate2643(.a(s_299), .b(gate95inter3), .O(gate95inter10));
  nor2  gate2644(.a(gate95inter10), .b(gate95inter9), .O(gate95inter11));
  nor2  gate2645(.a(gate95inter11), .b(gate95inter6), .O(gate95inter12));
  nand2 gate2646(.a(gate95inter12), .b(gate95inter1), .O(G416));

  xor2  gate2269(.a(G347), .b(G30), .O(gate96inter0));
  nand2 gate2270(.a(gate96inter0), .b(s_246), .O(gate96inter1));
  and2  gate2271(.a(G347), .b(G30), .O(gate96inter2));
  inv1  gate2272(.a(s_246), .O(gate96inter3));
  inv1  gate2273(.a(s_247), .O(gate96inter4));
  nand2 gate2274(.a(gate96inter4), .b(gate96inter3), .O(gate96inter5));
  nor2  gate2275(.a(gate96inter5), .b(gate96inter2), .O(gate96inter6));
  inv1  gate2276(.a(G30), .O(gate96inter7));
  inv1  gate2277(.a(G347), .O(gate96inter8));
  nand2 gate2278(.a(gate96inter8), .b(gate96inter7), .O(gate96inter9));
  nand2 gate2279(.a(s_247), .b(gate96inter3), .O(gate96inter10));
  nor2  gate2280(.a(gate96inter10), .b(gate96inter9), .O(gate96inter11));
  nor2  gate2281(.a(gate96inter11), .b(gate96inter6), .O(gate96inter12));
  nand2 gate2282(.a(gate96inter12), .b(gate96inter1), .O(G417));
nand2 gate97( .a(G19), .b(G350), .O(G418) );
nand2 gate98( .a(G23), .b(G350), .O(G419) );

  xor2  gate2521(.a(G353), .b(G27), .O(gate99inter0));
  nand2 gate2522(.a(gate99inter0), .b(s_282), .O(gate99inter1));
  and2  gate2523(.a(G353), .b(G27), .O(gate99inter2));
  inv1  gate2524(.a(s_282), .O(gate99inter3));
  inv1  gate2525(.a(s_283), .O(gate99inter4));
  nand2 gate2526(.a(gate99inter4), .b(gate99inter3), .O(gate99inter5));
  nor2  gate2527(.a(gate99inter5), .b(gate99inter2), .O(gate99inter6));
  inv1  gate2528(.a(G27), .O(gate99inter7));
  inv1  gate2529(.a(G353), .O(gate99inter8));
  nand2 gate2530(.a(gate99inter8), .b(gate99inter7), .O(gate99inter9));
  nand2 gate2531(.a(s_283), .b(gate99inter3), .O(gate99inter10));
  nor2  gate2532(.a(gate99inter10), .b(gate99inter9), .O(gate99inter11));
  nor2  gate2533(.a(gate99inter11), .b(gate99inter6), .O(gate99inter12));
  nand2 gate2534(.a(gate99inter12), .b(gate99inter1), .O(G420));
nand2 gate100( .a(G31), .b(G353), .O(G421) );

  xor2  gate1093(.a(G356), .b(G20), .O(gate101inter0));
  nand2 gate1094(.a(gate101inter0), .b(s_78), .O(gate101inter1));
  and2  gate1095(.a(G356), .b(G20), .O(gate101inter2));
  inv1  gate1096(.a(s_78), .O(gate101inter3));
  inv1  gate1097(.a(s_79), .O(gate101inter4));
  nand2 gate1098(.a(gate101inter4), .b(gate101inter3), .O(gate101inter5));
  nor2  gate1099(.a(gate101inter5), .b(gate101inter2), .O(gate101inter6));
  inv1  gate1100(.a(G20), .O(gate101inter7));
  inv1  gate1101(.a(G356), .O(gate101inter8));
  nand2 gate1102(.a(gate101inter8), .b(gate101inter7), .O(gate101inter9));
  nand2 gate1103(.a(s_79), .b(gate101inter3), .O(gate101inter10));
  nor2  gate1104(.a(gate101inter10), .b(gate101inter9), .O(gate101inter11));
  nor2  gate1105(.a(gate101inter11), .b(gate101inter6), .O(gate101inter12));
  nand2 gate1106(.a(gate101inter12), .b(gate101inter1), .O(G422));
nand2 gate102( .a(G24), .b(G356), .O(G423) );
nand2 gate103( .a(G28), .b(G359), .O(G424) );
nand2 gate104( .a(G32), .b(G359), .O(G425) );

  xor2  gate1989(.a(G363), .b(G362), .O(gate105inter0));
  nand2 gate1990(.a(gate105inter0), .b(s_206), .O(gate105inter1));
  and2  gate1991(.a(G363), .b(G362), .O(gate105inter2));
  inv1  gate1992(.a(s_206), .O(gate105inter3));
  inv1  gate1993(.a(s_207), .O(gate105inter4));
  nand2 gate1994(.a(gate105inter4), .b(gate105inter3), .O(gate105inter5));
  nor2  gate1995(.a(gate105inter5), .b(gate105inter2), .O(gate105inter6));
  inv1  gate1996(.a(G362), .O(gate105inter7));
  inv1  gate1997(.a(G363), .O(gate105inter8));
  nand2 gate1998(.a(gate105inter8), .b(gate105inter7), .O(gate105inter9));
  nand2 gate1999(.a(s_207), .b(gate105inter3), .O(gate105inter10));
  nor2  gate2000(.a(gate105inter10), .b(gate105inter9), .O(gate105inter11));
  nor2  gate2001(.a(gate105inter11), .b(gate105inter6), .O(gate105inter12));
  nand2 gate2002(.a(gate105inter12), .b(gate105inter1), .O(G426));

  xor2  gate1429(.a(G365), .b(G364), .O(gate106inter0));
  nand2 gate1430(.a(gate106inter0), .b(s_126), .O(gate106inter1));
  and2  gate1431(.a(G365), .b(G364), .O(gate106inter2));
  inv1  gate1432(.a(s_126), .O(gate106inter3));
  inv1  gate1433(.a(s_127), .O(gate106inter4));
  nand2 gate1434(.a(gate106inter4), .b(gate106inter3), .O(gate106inter5));
  nor2  gate1435(.a(gate106inter5), .b(gate106inter2), .O(gate106inter6));
  inv1  gate1436(.a(G364), .O(gate106inter7));
  inv1  gate1437(.a(G365), .O(gate106inter8));
  nand2 gate1438(.a(gate106inter8), .b(gate106inter7), .O(gate106inter9));
  nand2 gate1439(.a(s_127), .b(gate106inter3), .O(gate106inter10));
  nor2  gate1440(.a(gate106inter10), .b(gate106inter9), .O(gate106inter11));
  nor2  gate1441(.a(gate106inter11), .b(gate106inter6), .O(gate106inter12));
  nand2 gate1442(.a(gate106inter12), .b(gate106inter1), .O(G429));
nand2 gate107( .a(G366), .b(G367), .O(G432) );

  xor2  gate3123(.a(G369), .b(G368), .O(gate108inter0));
  nand2 gate3124(.a(gate108inter0), .b(s_368), .O(gate108inter1));
  and2  gate3125(.a(G369), .b(G368), .O(gate108inter2));
  inv1  gate3126(.a(s_368), .O(gate108inter3));
  inv1  gate3127(.a(s_369), .O(gate108inter4));
  nand2 gate3128(.a(gate108inter4), .b(gate108inter3), .O(gate108inter5));
  nor2  gate3129(.a(gate108inter5), .b(gate108inter2), .O(gate108inter6));
  inv1  gate3130(.a(G368), .O(gate108inter7));
  inv1  gate3131(.a(G369), .O(gate108inter8));
  nand2 gate3132(.a(gate108inter8), .b(gate108inter7), .O(gate108inter9));
  nand2 gate3133(.a(s_369), .b(gate108inter3), .O(gate108inter10));
  nor2  gate3134(.a(gate108inter10), .b(gate108inter9), .O(gate108inter11));
  nor2  gate3135(.a(gate108inter11), .b(gate108inter6), .O(gate108inter12));
  nand2 gate3136(.a(gate108inter12), .b(gate108inter1), .O(G435));
nand2 gate109( .a(G370), .b(G371), .O(G438) );

  xor2  gate1107(.a(G373), .b(G372), .O(gate110inter0));
  nand2 gate1108(.a(gate110inter0), .b(s_80), .O(gate110inter1));
  and2  gate1109(.a(G373), .b(G372), .O(gate110inter2));
  inv1  gate1110(.a(s_80), .O(gate110inter3));
  inv1  gate1111(.a(s_81), .O(gate110inter4));
  nand2 gate1112(.a(gate110inter4), .b(gate110inter3), .O(gate110inter5));
  nor2  gate1113(.a(gate110inter5), .b(gate110inter2), .O(gate110inter6));
  inv1  gate1114(.a(G372), .O(gate110inter7));
  inv1  gate1115(.a(G373), .O(gate110inter8));
  nand2 gate1116(.a(gate110inter8), .b(gate110inter7), .O(gate110inter9));
  nand2 gate1117(.a(s_81), .b(gate110inter3), .O(gate110inter10));
  nor2  gate1118(.a(gate110inter10), .b(gate110inter9), .O(gate110inter11));
  nor2  gate1119(.a(gate110inter11), .b(gate110inter6), .O(gate110inter12));
  nand2 gate1120(.a(gate110inter12), .b(gate110inter1), .O(G441));
nand2 gate111( .a(G374), .b(G375), .O(G444) );
nand2 gate112( .a(G376), .b(G377), .O(G447) );
nand2 gate113( .a(G378), .b(G379), .O(G450) );
nand2 gate114( .a(G380), .b(G381), .O(G453) );

  xor2  gate2801(.a(G383), .b(G382), .O(gate115inter0));
  nand2 gate2802(.a(gate115inter0), .b(s_322), .O(gate115inter1));
  and2  gate2803(.a(G383), .b(G382), .O(gate115inter2));
  inv1  gate2804(.a(s_322), .O(gate115inter3));
  inv1  gate2805(.a(s_323), .O(gate115inter4));
  nand2 gate2806(.a(gate115inter4), .b(gate115inter3), .O(gate115inter5));
  nor2  gate2807(.a(gate115inter5), .b(gate115inter2), .O(gate115inter6));
  inv1  gate2808(.a(G382), .O(gate115inter7));
  inv1  gate2809(.a(G383), .O(gate115inter8));
  nand2 gate2810(.a(gate115inter8), .b(gate115inter7), .O(gate115inter9));
  nand2 gate2811(.a(s_323), .b(gate115inter3), .O(gate115inter10));
  nor2  gate2812(.a(gate115inter10), .b(gate115inter9), .O(gate115inter11));
  nor2  gate2813(.a(gate115inter11), .b(gate115inter6), .O(gate115inter12));
  nand2 gate2814(.a(gate115inter12), .b(gate115inter1), .O(G456));
nand2 gate116( .a(G384), .b(G385), .O(G459) );
nand2 gate117( .a(G386), .b(G387), .O(G462) );

  xor2  gate2143(.a(G389), .b(G388), .O(gate118inter0));
  nand2 gate2144(.a(gate118inter0), .b(s_228), .O(gate118inter1));
  and2  gate2145(.a(G389), .b(G388), .O(gate118inter2));
  inv1  gate2146(.a(s_228), .O(gate118inter3));
  inv1  gate2147(.a(s_229), .O(gate118inter4));
  nand2 gate2148(.a(gate118inter4), .b(gate118inter3), .O(gate118inter5));
  nor2  gate2149(.a(gate118inter5), .b(gate118inter2), .O(gate118inter6));
  inv1  gate2150(.a(G388), .O(gate118inter7));
  inv1  gate2151(.a(G389), .O(gate118inter8));
  nand2 gate2152(.a(gate118inter8), .b(gate118inter7), .O(gate118inter9));
  nand2 gate2153(.a(s_229), .b(gate118inter3), .O(gate118inter10));
  nor2  gate2154(.a(gate118inter10), .b(gate118inter9), .O(gate118inter11));
  nor2  gate2155(.a(gate118inter11), .b(gate118inter6), .O(gate118inter12));
  nand2 gate2156(.a(gate118inter12), .b(gate118inter1), .O(G465));
nand2 gate119( .a(G390), .b(G391), .O(G468) );
nand2 gate120( .a(G392), .b(G393), .O(G471) );

  xor2  gate1625(.a(G395), .b(G394), .O(gate121inter0));
  nand2 gate1626(.a(gate121inter0), .b(s_154), .O(gate121inter1));
  and2  gate1627(.a(G395), .b(G394), .O(gate121inter2));
  inv1  gate1628(.a(s_154), .O(gate121inter3));
  inv1  gate1629(.a(s_155), .O(gate121inter4));
  nand2 gate1630(.a(gate121inter4), .b(gate121inter3), .O(gate121inter5));
  nor2  gate1631(.a(gate121inter5), .b(gate121inter2), .O(gate121inter6));
  inv1  gate1632(.a(G394), .O(gate121inter7));
  inv1  gate1633(.a(G395), .O(gate121inter8));
  nand2 gate1634(.a(gate121inter8), .b(gate121inter7), .O(gate121inter9));
  nand2 gate1635(.a(s_155), .b(gate121inter3), .O(gate121inter10));
  nor2  gate1636(.a(gate121inter10), .b(gate121inter9), .O(gate121inter11));
  nor2  gate1637(.a(gate121inter11), .b(gate121inter6), .O(gate121inter12));
  nand2 gate1638(.a(gate121inter12), .b(gate121inter1), .O(G474));
nand2 gate122( .a(G396), .b(G397), .O(G477) );

  xor2  gate2437(.a(G399), .b(G398), .O(gate123inter0));
  nand2 gate2438(.a(gate123inter0), .b(s_270), .O(gate123inter1));
  and2  gate2439(.a(G399), .b(G398), .O(gate123inter2));
  inv1  gate2440(.a(s_270), .O(gate123inter3));
  inv1  gate2441(.a(s_271), .O(gate123inter4));
  nand2 gate2442(.a(gate123inter4), .b(gate123inter3), .O(gate123inter5));
  nor2  gate2443(.a(gate123inter5), .b(gate123inter2), .O(gate123inter6));
  inv1  gate2444(.a(G398), .O(gate123inter7));
  inv1  gate2445(.a(G399), .O(gate123inter8));
  nand2 gate2446(.a(gate123inter8), .b(gate123inter7), .O(gate123inter9));
  nand2 gate2447(.a(s_271), .b(gate123inter3), .O(gate123inter10));
  nor2  gate2448(.a(gate123inter10), .b(gate123inter9), .O(gate123inter11));
  nor2  gate2449(.a(gate123inter11), .b(gate123inter6), .O(gate123inter12));
  nand2 gate2450(.a(gate123inter12), .b(gate123inter1), .O(G480));

  xor2  gate995(.a(G401), .b(G400), .O(gate124inter0));
  nand2 gate996(.a(gate124inter0), .b(s_64), .O(gate124inter1));
  and2  gate997(.a(G401), .b(G400), .O(gate124inter2));
  inv1  gate998(.a(s_64), .O(gate124inter3));
  inv1  gate999(.a(s_65), .O(gate124inter4));
  nand2 gate1000(.a(gate124inter4), .b(gate124inter3), .O(gate124inter5));
  nor2  gate1001(.a(gate124inter5), .b(gate124inter2), .O(gate124inter6));
  inv1  gate1002(.a(G400), .O(gate124inter7));
  inv1  gate1003(.a(G401), .O(gate124inter8));
  nand2 gate1004(.a(gate124inter8), .b(gate124inter7), .O(gate124inter9));
  nand2 gate1005(.a(s_65), .b(gate124inter3), .O(gate124inter10));
  nor2  gate1006(.a(gate124inter10), .b(gate124inter9), .O(gate124inter11));
  nor2  gate1007(.a(gate124inter11), .b(gate124inter6), .O(gate124inter12));
  nand2 gate1008(.a(gate124inter12), .b(gate124inter1), .O(G483));

  xor2  gate1499(.a(G403), .b(G402), .O(gate125inter0));
  nand2 gate1500(.a(gate125inter0), .b(s_136), .O(gate125inter1));
  and2  gate1501(.a(G403), .b(G402), .O(gate125inter2));
  inv1  gate1502(.a(s_136), .O(gate125inter3));
  inv1  gate1503(.a(s_137), .O(gate125inter4));
  nand2 gate1504(.a(gate125inter4), .b(gate125inter3), .O(gate125inter5));
  nor2  gate1505(.a(gate125inter5), .b(gate125inter2), .O(gate125inter6));
  inv1  gate1506(.a(G402), .O(gate125inter7));
  inv1  gate1507(.a(G403), .O(gate125inter8));
  nand2 gate1508(.a(gate125inter8), .b(gate125inter7), .O(gate125inter9));
  nand2 gate1509(.a(s_137), .b(gate125inter3), .O(gate125inter10));
  nor2  gate1510(.a(gate125inter10), .b(gate125inter9), .O(gate125inter11));
  nor2  gate1511(.a(gate125inter11), .b(gate125inter6), .O(gate125inter12));
  nand2 gate1512(.a(gate125inter12), .b(gate125inter1), .O(G486));

  xor2  gate3165(.a(G405), .b(G404), .O(gate126inter0));
  nand2 gate3166(.a(gate126inter0), .b(s_374), .O(gate126inter1));
  and2  gate3167(.a(G405), .b(G404), .O(gate126inter2));
  inv1  gate3168(.a(s_374), .O(gate126inter3));
  inv1  gate3169(.a(s_375), .O(gate126inter4));
  nand2 gate3170(.a(gate126inter4), .b(gate126inter3), .O(gate126inter5));
  nor2  gate3171(.a(gate126inter5), .b(gate126inter2), .O(gate126inter6));
  inv1  gate3172(.a(G404), .O(gate126inter7));
  inv1  gate3173(.a(G405), .O(gate126inter8));
  nand2 gate3174(.a(gate126inter8), .b(gate126inter7), .O(gate126inter9));
  nand2 gate3175(.a(s_375), .b(gate126inter3), .O(gate126inter10));
  nor2  gate3176(.a(gate126inter10), .b(gate126inter9), .O(gate126inter11));
  nor2  gate3177(.a(gate126inter11), .b(gate126inter6), .O(gate126inter12));
  nand2 gate3178(.a(gate126inter12), .b(gate126inter1), .O(G489));

  xor2  gate3025(.a(G407), .b(G406), .O(gate127inter0));
  nand2 gate3026(.a(gate127inter0), .b(s_354), .O(gate127inter1));
  and2  gate3027(.a(G407), .b(G406), .O(gate127inter2));
  inv1  gate3028(.a(s_354), .O(gate127inter3));
  inv1  gate3029(.a(s_355), .O(gate127inter4));
  nand2 gate3030(.a(gate127inter4), .b(gate127inter3), .O(gate127inter5));
  nor2  gate3031(.a(gate127inter5), .b(gate127inter2), .O(gate127inter6));
  inv1  gate3032(.a(G406), .O(gate127inter7));
  inv1  gate3033(.a(G407), .O(gate127inter8));
  nand2 gate3034(.a(gate127inter8), .b(gate127inter7), .O(gate127inter9));
  nand2 gate3035(.a(s_355), .b(gate127inter3), .O(gate127inter10));
  nor2  gate3036(.a(gate127inter10), .b(gate127inter9), .O(gate127inter11));
  nor2  gate3037(.a(gate127inter11), .b(gate127inter6), .O(gate127inter12));
  nand2 gate3038(.a(gate127inter12), .b(gate127inter1), .O(G492));

  xor2  gate2045(.a(G409), .b(G408), .O(gate128inter0));
  nand2 gate2046(.a(gate128inter0), .b(s_214), .O(gate128inter1));
  and2  gate2047(.a(G409), .b(G408), .O(gate128inter2));
  inv1  gate2048(.a(s_214), .O(gate128inter3));
  inv1  gate2049(.a(s_215), .O(gate128inter4));
  nand2 gate2050(.a(gate128inter4), .b(gate128inter3), .O(gate128inter5));
  nor2  gate2051(.a(gate128inter5), .b(gate128inter2), .O(gate128inter6));
  inv1  gate2052(.a(G408), .O(gate128inter7));
  inv1  gate2053(.a(G409), .O(gate128inter8));
  nand2 gate2054(.a(gate128inter8), .b(gate128inter7), .O(gate128inter9));
  nand2 gate2055(.a(s_215), .b(gate128inter3), .O(gate128inter10));
  nor2  gate2056(.a(gate128inter10), .b(gate128inter9), .O(gate128inter11));
  nor2  gate2057(.a(gate128inter11), .b(gate128inter6), .O(gate128inter12));
  nand2 gate2058(.a(gate128inter12), .b(gate128inter1), .O(G495));

  xor2  gate659(.a(G411), .b(G410), .O(gate129inter0));
  nand2 gate660(.a(gate129inter0), .b(s_16), .O(gate129inter1));
  and2  gate661(.a(G411), .b(G410), .O(gate129inter2));
  inv1  gate662(.a(s_16), .O(gate129inter3));
  inv1  gate663(.a(s_17), .O(gate129inter4));
  nand2 gate664(.a(gate129inter4), .b(gate129inter3), .O(gate129inter5));
  nor2  gate665(.a(gate129inter5), .b(gate129inter2), .O(gate129inter6));
  inv1  gate666(.a(G410), .O(gate129inter7));
  inv1  gate667(.a(G411), .O(gate129inter8));
  nand2 gate668(.a(gate129inter8), .b(gate129inter7), .O(gate129inter9));
  nand2 gate669(.a(s_17), .b(gate129inter3), .O(gate129inter10));
  nor2  gate670(.a(gate129inter10), .b(gate129inter9), .O(gate129inter11));
  nor2  gate671(.a(gate129inter11), .b(gate129inter6), .O(gate129inter12));
  nand2 gate672(.a(gate129inter12), .b(gate129inter1), .O(G498));

  xor2  gate2745(.a(G413), .b(G412), .O(gate130inter0));
  nand2 gate2746(.a(gate130inter0), .b(s_314), .O(gate130inter1));
  and2  gate2747(.a(G413), .b(G412), .O(gate130inter2));
  inv1  gate2748(.a(s_314), .O(gate130inter3));
  inv1  gate2749(.a(s_315), .O(gate130inter4));
  nand2 gate2750(.a(gate130inter4), .b(gate130inter3), .O(gate130inter5));
  nor2  gate2751(.a(gate130inter5), .b(gate130inter2), .O(gate130inter6));
  inv1  gate2752(.a(G412), .O(gate130inter7));
  inv1  gate2753(.a(G413), .O(gate130inter8));
  nand2 gate2754(.a(gate130inter8), .b(gate130inter7), .O(gate130inter9));
  nand2 gate2755(.a(s_315), .b(gate130inter3), .O(gate130inter10));
  nor2  gate2756(.a(gate130inter10), .b(gate130inter9), .O(gate130inter11));
  nor2  gate2757(.a(gate130inter11), .b(gate130inter6), .O(gate130inter12));
  nand2 gate2758(.a(gate130inter12), .b(gate130inter1), .O(G501));

  xor2  gate2787(.a(G415), .b(G414), .O(gate131inter0));
  nand2 gate2788(.a(gate131inter0), .b(s_320), .O(gate131inter1));
  and2  gate2789(.a(G415), .b(G414), .O(gate131inter2));
  inv1  gate2790(.a(s_320), .O(gate131inter3));
  inv1  gate2791(.a(s_321), .O(gate131inter4));
  nand2 gate2792(.a(gate131inter4), .b(gate131inter3), .O(gate131inter5));
  nor2  gate2793(.a(gate131inter5), .b(gate131inter2), .O(gate131inter6));
  inv1  gate2794(.a(G414), .O(gate131inter7));
  inv1  gate2795(.a(G415), .O(gate131inter8));
  nand2 gate2796(.a(gate131inter8), .b(gate131inter7), .O(gate131inter9));
  nand2 gate2797(.a(s_321), .b(gate131inter3), .O(gate131inter10));
  nor2  gate2798(.a(gate131inter10), .b(gate131inter9), .O(gate131inter11));
  nor2  gate2799(.a(gate131inter11), .b(gate131inter6), .O(gate131inter12));
  nand2 gate2800(.a(gate131inter12), .b(gate131inter1), .O(G504));
nand2 gate132( .a(G416), .b(G417), .O(G507) );
nand2 gate133( .a(G418), .b(G419), .O(G510) );
nand2 gate134( .a(G420), .b(G421), .O(G513) );
nand2 gate135( .a(G422), .b(G423), .O(G516) );

  xor2  gate2759(.a(G425), .b(G424), .O(gate136inter0));
  nand2 gate2760(.a(gate136inter0), .b(s_316), .O(gate136inter1));
  and2  gate2761(.a(G425), .b(G424), .O(gate136inter2));
  inv1  gate2762(.a(s_316), .O(gate136inter3));
  inv1  gate2763(.a(s_317), .O(gate136inter4));
  nand2 gate2764(.a(gate136inter4), .b(gate136inter3), .O(gate136inter5));
  nor2  gate2765(.a(gate136inter5), .b(gate136inter2), .O(gate136inter6));
  inv1  gate2766(.a(G424), .O(gate136inter7));
  inv1  gate2767(.a(G425), .O(gate136inter8));
  nand2 gate2768(.a(gate136inter8), .b(gate136inter7), .O(gate136inter9));
  nand2 gate2769(.a(s_317), .b(gate136inter3), .O(gate136inter10));
  nor2  gate2770(.a(gate136inter10), .b(gate136inter9), .O(gate136inter11));
  nor2  gate2771(.a(gate136inter11), .b(gate136inter6), .O(gate136inter12));
  nand2 gate2772(.a(gate136inter12), .b(gate136inter1), .O(G519));

  xor2  gate1793(.a(G429), .b(G426), .O(gate137inter0));
  nand2 gate1794(.a(gate137inter0), .b(s_178), .O(gate137inter1));
  and2  gate1795(.a(G429), .b(G426), .O(gate137inter2));
  inv1  gate1796(.a(s_178), .O(gate137inter3));
  inv1  gate1797(.a(s_179), .O(gate137inter4));
  nand2 gate1798(.a(gate137inter4), .b(gate137inter3), .O(gate137inter5));
  nor2  gate1799(.a(gate137inter5), .b(gate137inter2), .O(gate137inter6));
  inv1  gate1800(.a(G426), .O(gate137inter7));
  inv1  gate1801(.a(G429), .O(gate137inter8));
  nand2 gate1802(.a(gate137inter8), .b(gate137inter7), .O(gate137inter9));
  nand2 gate1803(.a(s_179), .b(gate137inter3), .O(gate137inter10));
  nor2  gate1804(.a(gate137inter10), .b(gate137inter9), .O(gate137inter11));
  nor2  gate1805(.a(gate137inter11), .b(gate137inter6), .O(gate137inter12));
  nand2 gate1806(.a(gate137inter12), .b(gate137inter1), .O(G522));
nand2 gate138( .a(G432), .b(G435), .O(G525) );

  xor2  gate1555(.a(G441), .b(G438), .O(gate139inter0));
  nand2 gate1556(.a(gate139inter0), .b(s_144), .O(gate139inter1));
  and2  gate1557(.a(G441), .b(G438), .O(gate139inter2));
  inv1  gate1558(.a(s_144), .O(gate139inter3));
  inv1  gate1559(.a(s_145), .O(gate139inter4));
  nand2 gate1560(.a(gate139inter4), .b(gate139inter3), .O(gate139inter5));
  nor2  gate1561(.a(gate139inter5), .b(gate139inter2), .O(gate139inter6));
  inv1  gate1562(.a(G438), .O(gate139inter7));
  inv1  gate1563(.a(G441), .O(gate139inter8));
  nand2 gate1564(.a(gate139inter8), .b(gate139inter7), .O(gate139inter9));
  nand2 gate1565(.a(s_145), .b(gate139inter3), .O(gate139inter10));
  nor2  gate1566(.a(gate139inter10), .b(gate139inter9), .O(gate139inter11));
  nor2  gate1567(.a(gate139inter11), .b(gate139inter6), .O(gate139inter12));
  nand2 gate1568(.a(gate139inter12), .b(gate139inter1), .O(G528));
nand2 gate140( .a(G444), .b(G447), .O(G531) );
nand2 gate141( .a(G450), .b(G453), .O(G534) );
nand2 gate142( .a(G456), .b(G459), .O(G537) );
nand2 gate143( .a(G462), .b(G465), .O(G540) );
nand2 gate144( .a(G468), .b(G471), .O(G543) );

  xor2  gate1835(.a(G477), .b(G474), .O(gate145inter0));
  nand2 gate1836(.a(gate145inter0), .b(s_184), .O(gate145inter1));
  and2  gate1837(.a(G477), .b(G474), .O(gate145inter2));
  inv1  gate1838(.a(s_184), .O(gate145inter3));
  inv1  gate1839(.a(s_185), .O(gate145inter4));
  nand2 gate1840(.a(gate145inter4), .b(gate145inter3), .O(gate145inter5));
  nor2  gate1841(.a(gate145inter5), .b(gate145inter2), .O(gate145inter6));
  inv1  gate1842(.a(G474), .O(gate145inter7));
  inv1  gate1843(.a(G477), .O(gate145inter8));
  nand2 gate1844(.a(gate145inter8), .b(gate145inter7), .O(gate145inter9));
  nand2 gate1845(.a(s_185), .b(gate145inter3), .O(gate145inter10));
  nor2  gate1846(.a(gate145inter10), .b(gate145inter9), .O(gate145inter11));
  nor2  gate1847(.a(gate145inter11), .b(gate145inter6), .O(gate145inter12));
  nand2 gate1848(.a(gate145inter12), .b(gate145inter1), .O(G546));
nand2 gate146( .a(G480), .b(G483), .O(G549) );
nand2 gate147( .a(G486), .b(G489), .O(G552) );

  xor2  gate2367(.a(G495), .b(G492), .O(gate148inter0));
  nand2 gate2368(.a(gate148inter0), .b(s_260), .O(gate148inter1));
  and2  gate2369(.a(G495), .b(G492), .O(gate148inter2));
  inv1  gate2370(.a(s_260), .O(gate148inter3));
  inv1  gate2371(.a(s_261), .O(gate148inter4));
  nand2 gate2372(.a(gate148inter4), .b(gate148inter3), .O(gate148inter5));
  nor2  gate2373(.a(gate148inter5), .b(gate148inter2), .O(gate148inter6));
  inv1  gate2374(.a(G492), .O(gate148inter7));
  inv1  gate2375(.a(G495), .O(gate148inter8));
  nand2 gate2376(.a(gate148inter8), .b(gate148inter7), .O(gate148inter9));
  nand2 gate2377(.a(s_261), .b(gate148inter3), .O(gate148inter10));
  nor2  gate2378(.a(gate148inter10), .b(gate148inter9), .O(gate148inter11));
  nor2  gate2379(.a(gate148inter11), .b(gate148inter6), .O(gate148inter12));
  nand2 gate2380(.a(gate148inter12), .b(gate148inter1), .O(G555));

  xor2  gate1415(.a(G501), .b(G498), .O(gate149inter0));
  nand2 gate1416(.a(gate149inter0), .b(s_124), .O(gate149inter1));
  and2  gate1417(.a(G501), .b(G498), .O(gate149inter2));
  inv1  gate1418(.a(s_124), .O(gate149inter3));
  inv1  gate1419(.a(s_125), .O(gate149inter4));
  nand2 gate1420(.a(gate149inter4), .b(gate149inter3), .O(gate149inter5));
  nor2  gate1421(.a(gate149inter5), .b(gate149inter2), .O(gate149inter6));
  inv1  gate1422(.a(G498), .O(gate149inter7));
  inv1  gate1423(.a(G501), .O(gate149inter8));
  nand2 gate1424(.a(gate149inter8), .b(gate149inter7), .O(gate149inter9));
  nand2 gate1425(.a(s_125), .b(gate149inter3), .O(gate149inter10));
  nor2  gate1426(.a(gate149inter10), .b(gate149inter9), .O(gate149inter11));
  nor2  gate1427(.a(gate149inter11), .b(gate149inter6), .O(gate149inter12));
  nand2 gate1428(.a(gate149inter12), .b(gate149inter1), .O(G558));
nand2 gate150( .a(G504), .b(G507), .O(G561) );
nand2 gate151( .a(G510), .b(G513), .O(G564) );

  xor2  gate1317(.a(G519), .b(G516), .O(gate152inter0));
  nand2 gate1318(.a(gate152inter0), .b(s_110), .O(gate152inter1));
  and2  gate1319(.a(G519), .b(G516), .O(gate152inter2));
  inv1  gate1320(.a(s_110), .O(gate152inter3));
  inv1  gate1321(.a(s_111), .O(gate152inter4));
  nand2 gate1322(.a(gate152inter4), .b(gate152inter3), .O(gate152inter5));
  nor2  gate1323(.a(gate152inter5), .b(gate152inter2), .O(gate152inter6));
  inv1  gate1324(.a(G516), .O(gate152inter7));
  inv1  gate1325(.a(G519), .O(gate152inter8));
  nand2 gate1326(.a(gate152inter8), .b(gate152inter7), .O(gate152inter9));
  nand2 gate1327(.a(s_111), .b(gate152inter3), .O(gate152inter10));
  nor2  gate1328(.a(gate152inter10), .b(gate152inter9), .O(gate152inter11));
  nor2  gate1329(.a(gate152inter11), .b(gate152inter6), .O(gate152inter12));
  nand2 gate1330(.a(gate152inter12), .b(gate152inter1), .O(G567));
nand2 gate153( .a(G426), .b(G522), .O(G570) );

  xor2  gate631(.a(G522), .b(G429), .O(gate154inter0));
  nand2 gate632(.a(gate154inter0), .b(s_12), .O(gate154inter1));
  and2  gate633(.a(G522), .b(G429), .O(gate154inter2));
  inv1  gate634(.a(s_12), .O(gate154inter3));
  inv1  gate635(.a(s_13), .O(gate154inter4));
  nand2 gate636(.a(gate154inter4), .b(gate154inter3), .O(gate154inter5));
  nor2  gate637(.a(gate154inter5), .b(gate154inter2), .O(gate154inter6));
  inv1  gate638(.a(G429), .O(gate154inter7));
  inv1  gate639(.a(G522), .O(gate154inter8));
  nand2 gate640(.a(gate154inter8), .b(gate154inter7), .O(gate154inter9));
  nand2 gate641(.a(s_13), .b(gate154inter3), .O(gate154inter10));
  nor2  gate642(.a(gate154inter10), .b(gate154inter9), .O(gate154inter11));
  nor2  gate643(.a(gate154inter11), .b(gate154inter6), .O(gate154inter12));
  nand2 gate644(.a(gate154inter12), .b(gate154inter1), .O(G571));
nand2 gate155( .a(G432), .b(G525), .O(G572) );

  xor2  gate2311(.a(G525), .b(G435), .O(gate156inter0));
  nand2 gate2312(.a(gate156inter0), .b(s_252), .O(gate156inter1));
  and2  gate2313(.a(G525), .b(G435), .O(gate156inter2));
  inv1  gate2314(.a(s_252), .O(gate156inter3));
  inv1  gate2315(.a(s_253), .O(gate156inter4));
  nand2 gate2316(.a(gate156inter4), .b(gate156inter3), .O(gate156inter5));
  nor2  gate2317(.a(gate156inter5), .b(gate156inter2), .O(gate156inter6));
  inv1  gate2318(.a(G435), .O(gate156inter7));
  inv1  gate2319(.a(G525), .O(gate156inter8));
  nand2 gate2320(.a(gate156inter8), .b(gate156inter7), .O(gate156inter9));
  nand2 gate2321(.a(s_253), .b(gate156inter3), .O(gate156inter10));
  nor2  gate2322(.a(gate156inter10), .b(gate156inter9), .O(gate156inter11));
  nor2  gate2323(.a(gate156inter11), .b(gate156inter6), .O(gate156inter12));
  nand2 gate2324(.a(gate156inter12), .b(gate156inter1), .O(G573));
nand2 gate157( .a(G438), .b(G528), .O(G574) );

  xor2  gate3053(.a(G528), .b(G441), .O(gate158inter0));
  nand2 gate3054(.a(gate158inter0), .b(s_358), .O(gate158inter1));
  and2  gate3055(.a(G528), .b(G441), .O(gate158inter2));
  inv1  gate3056(.a(s_358), .O(gate158inter3));
  inv1  gate3057(.a(s_359), .O(gate158inter4));
  nand2 gate3058(.a(gate158inter4), .b(gate158inter3), .O(gate158inter5));
  nor2  gate3059(.a(gate158inter5), .b(gate158inter2), .O(gate158inter6));
  inv1  gate3060(.a(G441), .O(gate158inter7));
  inv1  gate3061(.a(G528), .O(gate158inter8));
  nand2 gate3062(.a(gate158inter8), .b(gate158inter7), .O(gate158inter9));
  nand2 gate3063(.a(s_359), .b(gate158inter3), .O(gate158inter10));
  nor2  gate3064(.a(gate158inter10), .b(gate158inter9), .O(gate158inter11));
  nor2  gate3065(.a(gate158inter11), .b(gate158inter6), .O(gate158inter12));
  nand2 gate3066(.a(gate158inter12), .b(gate158inter1), .O(G575));

  xor2  gate1443(.a(G531), .b(G444), .O(gate159inter0));
  nand2 gate1444(.a(gate159inter0), .b(s_128), .O(gate159inter1));
  and2  gate1445(.a(G531), .b(G444), .O(gate159inter2));
  inv1  gate1446(.a(s_128), .O(gate159inter3));
  inv1  gate1447(.a(s_129), .O(gate159inter4));
  nand2 gate1448(.a(gate159inter4), .b(gate159inter3), .O(gate159inter5));
  nor2  gate1449(.a(gate159inter5), .b(gate159inter2), .O(gate159inter6));
  inv1  gate1450(.a(G444), .O(gate159inter7));
  inv1  gate1451(.a(G531), .O(gate159inter8));
  nand2 gate1452(.a(gate159inter8), .b(gate159inter7), .O(gate159inter9));
  nand2 gate1453(.a(s_129), .b(gate159inter3), .O(gate159inter10));
  nor2  gate1454(.a(gate159inter10), .b(gate159inter9), .O(gate159inter11));
  nor2  gate1455(.a(gate159inter11), .b(gate159inter6), .O(gate159inter12));
  nand2 gate1456(.a(gate159inter12), .b(gate159inter1), .O(G576));
nand2 gate160( .a(G447), .b(G531), .O(G577) );
nand2 gate161( .a(G450), .b(G534), .O(G578) );

  xor2  gate1863(.a(G534), .b(G453), .O(gate162inter0));
  nand2 gate1864(.a(gate162inter0), .b(s_188), .O(gate162inter1));
  and2  gate1865(.a(G534), .b(G453), .O(gate162inter2));
  inv1  gate1866(.a(s_188), .O(gate162inter3));
  inv1  gate1867(.a(s_189), .O(gate162inter4));
  nand2 gate1868(.a(gate162inter4), .b(gate162inter3), .O(gate162inter5));
  nor2  gate1869(.a(gate162inter5), .b(gate162inter2), .O(gate162inter6));
  inv1  gate1870(.a(G453), .O(gate162inter7));
  inv1  gate1871(.a(G534), .O(gate162inter8));
  nand2 gate1872(.a(gate162inter8), .b(gate162inter7), .O(gate162inter9));
  nand2 gate1873(.a(s_189), .b(gate162inter3), .O(gate162inter10));
  nor2  gate1874(.a(gate162inter10), .b(gate162inter9), .O(gate162inter11));
  nor2  gate1875(.a(gate162inter11), .b(gate162inter6), .O(gate162inter12));
  nand2 gate1876(.a(gate162inter12), .b(gate162inter1), .O(G579));

  xor2  gate2941(.a(G537), .b(G456), .O(gate163inter0));
  nand2 gate2942(.a(gate163inter0), .b(s_342), .O(gate163inter1));
  and2  gate2943(.a(G537), .b(G456), .O(gate163inter2));
  inv1  gate2944(.a(s_342), .O(gate163inter3));
  inv1  gate2945(.a(s_343), .O(gate163inter4));
  nand2 gate2946(.a(gate163inter4), .b(gate163inter3), .O(gate163inter5));
  nor2  gate2947(.a(gate163inter5), .b(gate163inter2), .O(gate163inter6));
  inv1  gate2948(.a(G456), .O(gate163inter7));
  inv1  gate2949(.a(G537), .O(gate163inter8));
  nand2 gate2950(.a(gate163inter8), .b(gate163inter7), .O(gate163inter9));
  nand2 gate2951(.a(s_343), .b(gate163inter3), .O(gate163inter10));
  nor2  gate2952(.a(gate163inter10), .b(gate163inter9), .O(gate163inter11));
  nor2  gate2953(.a(gate163inter11), .b(gate163inter6), .O(gate163inter12));
  nand2 gate2954(.a(gate163inter12), .b(gate163inter1), .O(G580));

  xor2  gate2661(.a(G537), .b(G459), .O(gate164inter0));
  nand2 gate2662(.a(gate164inter0), .b(s_302), .O(gate164inter1));
  and2  gate2663(.a(G537), .b(G459), .O(gate164inter2));
  inv1  gate2664(.a(s_302), .O(gate164inter3));
  inv1  gate2665(.a(s_303), .O(gate164inter4));
  nand2 gate2666(.a(gate164inter4), .b(gate164inter3), .O(gate164inter5));
  nor2  gate2667(.a(gate164inter5), .b(gate164inter2), .O(gate164inter6));
  inv1  gate2668(.a(G459), .O(gate164inter7));
  inv1  gate2669(.a(G537), .O(gate164inter8));
  nand2 gate2670(.a(gate164inter8), .b(gate164inter7), .O(gate164inter9));
  nand2 gate2671(.a(s_303), .b(gate164inter3), .O(gate164inter10));
  nor2  gate2672(.a(gate164inter10), .b(gate164inter9), .O(gate164inter11));
  nor2  gate2673(.a(gate164inter11), .b(gate164inter6), .O(gate164inter12));
  nand2 gate2674(.a(gate164inter12), .b(gate164inter1), .O(G581));
nand2 gate165( .a(G462), .b(G540), .O(G582) );

  xor2  gate1387(.a(G540), .b(G465), .O(gate166inter0));
  nand2 gate1388(.a(gate166inter0), .b(s_120), .O(gate166inter1));
  and2  gate1389(.a(G540), .b(G465), .O(gate166inter2));
  inv1  gate1390(.a(s_120), .O(gate166inter3));
  inv1  gate1391(.a(s_121), .O(gate166inter4));
  nand2 gate1392(.a(gate166inter4), .b(gate166inter3), .O(gate166inter5));
  nor2  gate1393(.a(gate166inter5), .b(gate166inter2), .O(gate166inter6));
  inv1  gate1394(.a(G465), .O(gate166inter7));
  inv1  gate1395(.a(G540), .O(gate166inter8));
  nand2 gate1396(.a(gate166inter8), .b(gate166inter7), .O(gate166inter9));
  nand2 gate1397(.a(s_121), .b(gate166inter3), .O(gate166inter10));
  nor2  gate1398(.a(gate166inter10), .b(gate166inter9), .O(gate166inter11));
  nor2  gate1399(.a(gate166inter11), .b(gate166inter6), .O(gate166inter12));
  nand2 gate1400(.a(gate166inter12), .b(gate166inter1), .O(G583));

  xor2  gate2409(.a(G543), .b(G468), .O(gate167inter0));
  nand2 gate2410(.a(gate167inter0), .b(s_266), .O(gate167inter1));
  and2  gate2411(.a(G543), .b(G468), .O(gate167inter2));
  inv1  gate2412(.a(s_266), .O(gate167inter3));
  inv1  gate2413(.a(s_267), .O(gate167inter4));
  nand2 gate2414(.a(gate167inter4), .b(gate167inter3), .O(gate167inter5));
  nor2  gate2415(.a(gate167inter5), .b(gate167inter2), .O(gate167inter6));
  inv1  gate2416(.a(G468), .O(gate167inter7));
  inv1  gate2417(.a(G543), .O(gate167inter8));
  nand2 gate2418(.a(gate167inter8), .b(gate167inter7), .O(gate167inter9));
  nand2 gate2419(.a(s_267), .b(gate167inter3), .O(gate167inter10));
  nor2  gate2420(.a(gate167inter10), .b(gate167inter9), .O(gate167inter11));
  nor2  gate2421(.a(gate167inter11), .b(gate167inter6), .O(gate167inter12));
  nand2 gate2422(.a(gate167inter12), .b(gate167inter1), .O(G584));
nand2 gate168( .a(G471), .b(G543), .O(G585) );
nand2 gate169( .a(G474), .b(G546), .O(G586) );

  xor2  gate3137(.a(G546), .b(G477), .O(gate170inter0));
  nand2 gate3138(.a(gate170inter0), .b(s_370), .O(gate170inter1));
  and2  gate3139(.a(G546), .b(G477), .O(gate170inter2));
  inv1  gate3140(.a(s_370), .O(gate170inter3));
  inv1  gate3141(.a(s_371), .O(gate170inter4));
  nand2 gate3142(.a(gate170inter4), .b(gate170inter3), .O(gate170inter5));
  nor2  gate3143(.a(gate170inter5), .b(gate170inter2), .O(gate170inter6));
  inv1  gate3144(.a(G477), .O(gate170inter7));
  inv1  gate3145(.a(G546), .O(gate170inter8));
  nand2 gate3146(.a(gate170inter8), .b(gate170inter7), .O(gate170inter9));
  nand2 gate3147(.a(s_371), .b(gate170inter3), .O(gate170inter10));
  nor2  gate3148(.a(gate170inter10), .b(gate170inter9), .O(gate170inter11));
  nor2  gate3149(.a(gate170inter11), .b(gate170inter6), .O(gate170inter12));
  nand2 gate3150(.a(gate170inter12), .b(gate170inter1), .O(G587));

  xor2  gate2871(.a(G549), .b(G480), .O(gate171inter0));
  nand2 gate2872(.a(gate171inter0), .b(s_332), .O(gate171inter1));
  and2  gate2873(.a(G549), .b(G480), .O(gate171inter2));
  inv1  gate2874(.a(s_332), .O(gate171inter3));
  inv1  gate2875(.a(s_333), .O(gate171inter4));
  nand2 gate2876(.a(gate171inter4), .b(gate171inter3), .O(gate171inter5));
  nor2  gate2877(.a(gate171inter5), .b(gate171inter2), .O(gate171inter6));
  inv1  gate2878(.a(G480), .O(gate171inter7));
  inv1  gate2879(.a(G549), .O(gate171inter8));
  nand2 gate2880(.a(gate171inter8), .b(gate171inter7), .O(gate171inter9));
  nand2 gate2881(.a(s_333), .b(gate171inter3), .O(gate171inter10));
  nor2  gate2882(.a(gate171inter10), .b(gate171inter9), .O(gate171inter11));
  nor2  gate2883(.a(gate171inter11), .b(gate171inter6), .O(gate171inter12));
  nand2 gate2884(.a(gate171inter12), .b(gate171inter1), .O(G588));
nand2 gate172( .a(G483), .b(G549), .O(G589) );

  xor2  gate2017(.a(G552), .b(G486), .O(gate173inter0));
  nand2 gate2018(.a(gate173inter0), .b(s_210), .O(gate173inter1));
  and2  gate2019(.a(G552), .b(G486), .O(gate173inter2));
  inv1  gate2020(.a(s_210), .O(gate173inter3));
  inv1  gate2021(.a(s_211), .O(gate173inter4));
  nand2 gate2022(.a(gate173inter4), .b(gate173inter3), .O(gate173inter5));
  nor2  gate2023(.a(gate173inter5), .b(gate173inter2), .O(gate173inter6));
  inv1  gate2024(.a(G486), .O(gate173inter7));
  inv1  gate2025(.a(G552), .O(gate173inter8));
  nand2 gate2026(.a(gate173inter8), .b(gate173inter7), .O(gate173inter9));
  nand2 gate2027(.a(s_211), .b(gate173inter3), .O(gate173inter10));
  nor2  gate2028(.a(gate173inter10), .b(gate173inter9), .O(gate173inter11));
  nor2  gate2029(.a(gate173inter11), .b(gate173inter6), .O(gate173inter12));
  nand2 gate2030(.a(gate173inter12), .b(gate173inter1), .O(G590));

  xor2  gate2815(.a(G552), .b(G489), .O(gate174inter0));
  nand2 gate2816(.a(gate174inter0), .b(s_324), .O(gate174inter1));
  and2  gate2817(.a(G552), .b(G489), .O(gate174inter2));
  inv1  gate2818(.a(s_324), .O(gate174inter3));
  inv1  gate2819(.a(s_325), .O(gate174inter4));
  nand2 gate2820(.a(gate174inter4), .b(gate174inter3), .O(gate174inter5));
  nor2  gate2821(.a(gate174inter5), .b(gate174inter2), .O(gate174inter6));
  inv1  gate2822(.a(G489), .O(gate174inter7));
  inv1  gate2823(.a(G552), .O(gate174inter8));
  nand2 gate2824(.a(gate174inter8), .b(gate174inter7), .O(gate174inter9));
  nand2 gate2825(.a(s_325), .b(gate174inter3), .O(gate174inter10));
  nor2  gate2826(.a(gate174inter10), .b(gate174inter9), .O(gate174inter11));
  nor2  gate2827(.a(gate174inter11), .b(gate174inter6), .O(gate174inter12));
  nand2 gate2828(.a(gate174inter12), .b(gate174inter1), .O(G591));
nand2 gate175( .a(G492), .b(G555), .O(G592) );
nand2 gate176( .a(G495), .b(G555), .O(G593) );
nand2 gate177( .a(G498), .b(G558), .O(G594) );
nand2 gate178( .a(G501), .b(G558), .O(G595) );

  xor2  gate2703(.a(G561), .b(G504), .O(gate179inter0));
  nand2 gate2704(.a(gate179inter0), .b(s_308), .O(gate179inter1));
  and2  gate2705(.a(G561), .b(G504), .O(gate179inter2));
  inv1  gate2706(.a(s_308), .O(gate179inter3));
  inv1  gate2707(.a(s_309), .O(gate179inter4));
  nand2 gate2708(.a(gate179inter4), .b(gate179inter3), .O(gate179inter5));
  nor2  gate2709(.a(gate179inter5), .b(gate179inter2), .O(gate179inter6));
  inv1  gate2710(.a(G504), .O(gate179inter7));
  inv1  gate2711(.a(G561), .O(gate179inter8));
  nand2 gate2712(.a(gate179inter8), .b(gate179inter7), .O(gate179inter9));
  nand2 gate2713(.a(s_309), .b(gate179inter3), .O(gate179inter10));
  nor2  gate2714(.a(gate179inter10), .b(gate179inter9), .O(gate179inter11));
  nor2  gate2715(.a(gate179inter11), .b(gate179inter6), .O(gate179inter12));
  nand2 gate2716(.a(gate179inter12), .b(gate179inter1), .O(G596));

  xor2  gate953(.a(G561), .b(G507), .O(gate180inter0));
  nand2 gate954(.a(gate180inter0), .b(s_58), .O(gate180inter1));
  and2  gate955(.a(G561), .b(G507), .O(gate180inter2));
  inv1  gate956(.a(s_58), .O(gate180inter3));
  inv1  gate957(.a(s_59), .O(gate180inter4));
  nand2 gate958(.a(gate180inter4), .b(gate180inter3), .O(gate180inter5));
  nor2  gate959(.a(gate180inter5), .b(gate180inter2), .O(gate180inter6));
  inv1  gate960(.a(G507), .O(gate180inter7));
  inv1  gate961(.a(G561), .O(gate180inter8));
  nand2 gate962(.a(gate180inter8), .b(gate180inter7), .O(gate180inter9));
  nand2 gate963(.a(s_59), .b(gate180inter3), .O(gate180inter10));
  nor2  gate964(.a(gate180inter10), .b(gate180inter9), .O(gate180inter11));
  nor2  gate965(.a(gate180inter11), .b(gate180inter6), .O(gate180inter12));
  nand2 gate966(.a(gate180inter12), .b(gate180inter1), .O(G597));

  xor2  gate1765(.a(G564), .b(G510), .O(gate181inter0));
  nand2 gate1766(.a(gate181inter0), .b(s_174), .O(gate181inter1));
  and2  gate1767(.a(G564), .b(G510), .O(gate181inter2));
  inv1  gate1768(.a(s_174), .O(gate181inter3));
  inv1  gate1769(.a(s_175), .O(gate181inter4));
  nand2 gate1770(.a(gate181inter4), .b(gate181inter3), .O(gate181inter5));
  nor2  gate1771(.a(gate181inter5), .b(gate181inter2), .O(gate181inter6));
  inv1  gate1772(.a(G510), .O(gate181inter7));
  inv1  gate1773(.a(G564), .O(gate181inter8));
  nand2 gate1774(.a(gate181inter8), .b(gate181inter7), .O(gate181inter9));
  nand2 gate1775(.a(s_175), .b(gate181inter3), .O(gate181inter10));
  nor2  gate1776(.a(gate181inter10), .b(gate181inter9), .O(gate181inter11));
  nor2  gate1777(.a(gate181inter11), .b(gate181inter6), .O(gate181inter12));
  nand2 gate1778(.a(gate181inter12), .b(gate181inter1), .O(G598));

  xor2  gate967(.a(G564), .b(G513), .O(gate182inter0));
  nand2 gate968(.a(gate182inter0), .b(s_60), .O(gate182inter1));
  and2  gate969(.a(G564), .b(G513), .O(gate182inter2));
  inv1  gate970(.a(s_60), .O(gate182inter3));
  inv1  gate971(.a(s_61), .O(gate182inter4));
  nand2 gate972(.a(gate182inter4), .b(gate182inter3), .O(gate182inter5));
  nor2  gate973(.a(gate182inter5), .b(gate182inter2), .O(gate182inter6));
  inv1  gate974(.a(G513), .O(gate182inter7));
  inv1  gate975(.a(G564), .O(gate182inter8));
  nand2 gate976(.a(gate182inter8), .b(gate182inter7), .O(gate182inter9));
  nand2 gate977(.a(s_61), .b(gate182inter3), .O(gate182inter10));
  nor2  gate978(.a(gate182inter10), .b(gate182inter9), .O(gate182inter11));
  nor2  gate979(.a(gate182inter11), .b(gate182inter6), .O(gate182inter12));
  nand2 gate980(.a(gate182inter12), .b(gate182inter1), .O(G599));
nand2 gate183( .a(G516), .b(G567), .O(G600) );
nand2 gate184( .a(G519), .b(G567), .O(G601) );

  xor2  gate785(.a(G571), .b(G570), .O(gate185inter0));
  nand2 gate786(.a(gate185inter0), .b(s_34), .O(gate185inter1));
  and2  gate787(.a(G571), .b(G570), .O(gate185inter2));
  inv1  gate788(.a(s_34), .O(gate185inter3));
  inv1  gate789(.a(s_35), .O(gate185inter4));
  nand2 gate790(.a(gate185inter4), .b(gate185inter3), .O(gate185inter5));
  nor2  gate791(.a(gate185inter5), .b(gate185inter2), .O(gate185inter6));
  inv1  gate792(.a(G570), .O(gate185inter7));
  inv1  gate793(.a(G571), .O(gate185inter8));
  nand2 gate794(.a(gate185inter8), .b(gate185inter7), .O(gate185inter9));
  nand2 gate795(.a(s_35), .b(gate185inter3), .O(gate185inter10));
  nor2  gate796(.a(gate185inter10), .b(gate185inter9), .O(gate185inter11));
  nor2  gate797(.a(gate185inter11), .b(gate185inter6), .O(gate185inter12));
  nand2 gate798(.a(gate185inter12), .b(gate185inter1), .O(G602));

  xor2  gate617(.a(G573), .b(G572), .O(gate186inter0));
  nand2 gate618(.a(gate186inter0), .b(s_10), .O(gate186inter1));
  and2  gate619(.a(G573), .b(G572), .O(gate186inter2));
  inv1  gate620(.a(s_10), .O(gate186inter3));
  inv1  gate621(.a(s_11), .O(gate186inter4));
  nand2 gate622(.a(gate186inter4), .b(gate186inter3), .O(gate186inter5));
  nor2  gate623(.a(gate186inter5), .b(gate186inter2), .O(gate186inter6));
  inv1  gate624(.a(G572), .O(gate186inter7));
  inv1  gate625(.a(G573), .O(gate186inter8));
  nand2 gate626(.a(gate186inter8), .b(gate186inter7), .O(gate186inter9));
  nand2 gate627(.a(s_11), .b(gate186inter3), .O(gate186inter10));
  nor2  gate628(.a(gate186inter10), .b(gate186inter9), .O(gate186inter11));
  nor2  gate629(.a(gate186inter11), .b(gate186inter6), .O(gate186inter12));
  nand2 gate630(.a(gate186inter12), .b(gate186inter1), .O(G607));
nand2 gate187( .a(G574), .b(G575), .O(G612) );

  xor2  gate757(.a(G577), .b(G576), .O(gate188inter0));
  nand2 gate758(.a(gate188inter0), .b(s_30), .O(gate188inter1));
  and2  gate759(.a(G577), .b(G576), .O(gate188inter2));
  inv1  gate760(.a(s_30), .O(gate188inter3));
  inv1  gate761(.a(s_31), .O(gate188inter4));
  nand2 gate762(.a(gate188inter4), .b(gate188inter3), .O(gate188inter5));
  nor2  gate763(.a(gate188inter5), .b(gate188inter2), .O(gate188inter6));
  inv1  gate764(.a(G576), .O(gate188inter7));
  inv1  gate765(.a(G577), .O(gate188inter8));
  nand2 gate766(.a(gate188inter8), .b(gate188inter7), .O(gate188inter9));
  nand2 gate767(.a(s_31), .b(gate188inter3), .O(gate188inter10));
  nor2  gate768(.a(gate188inter10), .b(gate188inter9), .O(gate188inter11));
  nor2  gate769(.a(gate188inter11), .b(gate188inter6), .O(gate188inter12));
  nand2 gate770(.a(gate188inter12), .b(gate188inter1), .O(G617));

  xor2  gate715(.a(G579), .b(G578), .O(gate189inter0));
  nand2 gate716(.a(gate189inter0), .b(s_24), .O(gate189inter1));
  and2  gate717(.a(G579), .b(G578), .O(gate189inter2));
  inv1  gate718(.a(s_24), .O(gate189inter3));
  inv1  gate719(.a(s_25), .O(gate189inter4));
  nand2 gate720(.a(gate189inter4), .b(gate189inter3), .O(gate189inter5));
  nor2  gate721(.a(gate189inter5), .b(gate189inter2), .O(gate189inter6));
  inv1  gate722(.a(G578), .O(gate189inter7));
  inv1  gate723(.a(G579), .O(gate189inter8));
  nand2 gate724(.a(gate189inter8), .b(gate189inter7), .O(gate189inter9));
  nand2 gate725(.a(s_25), .b(gate189inter3), .O(gate189inter10));
  nor2  gate726(.a(gate189inter10), .b(gate189inter9), .O(gate189inter11));
  nor2  gate727(.a(gate189inter11), .b(gate189inter6), .O(gate189inter12));
  nand2 gate728(.a(gate189inter12), .b(gate189inter1), .O(G622));

  xor2  gate1779(.a(G581), .b(G580), .O(gate190inter0));
  nand2 gate1780(.a(gate190inter0), .b(s_176), .O(gate190inter1));
  and2  gate1781(.a(G581), .b(G580), .O(gate190inter2));
  inv1  gate1782(.a(s_176), .O(gate190inter3));
  inv1  gate1783(.a(s_177), .O(gate190inter4));
  nand2 gate1784(.a(gate190inter4), .b(gate190inter3), .O(gate190inter5));
  nor2  gate1785(.a(gate190inter5), .b(gate190inter2), .O(gate190inter6));
  inv1  gate1786(.a(G580), .O(gate190inter7));
  inv1  gate1787(.a(G581), .O(gate190inter8));
  nand2 gate1788(.a(gate190inter8), .b(gate190inter7), .O(gate190inter9));
  nand2 gate1789(.a(s_177), .b(gate190inter3), .O(gate190inter10));
  nor2  gate1790(.a(gate190inter10), .b(gate190inter9), .O(gate190inter11));
  nor2  gate1791(.a(gate190inter11), .b(gate190inter6), .O(gate190inter12));
  nand2 gate1792(.a(gate190inter12), .b(gate190inter1), .O(G627));
nand2 gate191( .a(G582), .b(G583), .O(G632) );

  xor2  gate3067(.a(G585), .b(G584), .O(gate192inter0));
  nand2 gate3068(.a(gate192inter0), .b(s_360), .O(gate192inter1));
  and2  gate3069(.a(G585), .b(G584), .O(gate192inter2));
  inv1  gate3070(.a(s_360), .O(gate192inter3));
  inv1  gate3071(.a(s_361), .O(gate192inter4));
  nand2 gate3072(.a(gate192inter4), .b(gate192inter3), .O(gate192inter5));
  nor2  gate3073(.a(gate192inter5), .b(gate192inter2), .O(gate192inter6));
  inv1  gate3074(.a(G584), .O(gate192inter7));
  inv1  gate3075(.a(G585), .O(gate192inter8));
  nand2 gate3076(.a(gate192inter8), .b(gate192inter7), .O(gate192inter9));
  nand2 gate3077(.a(s_361), .b(gate192inter3), .O(gate192inter10));
  nor2  gate3078(.a(gate192inter10), .b(gate192inter9), .O(gate192inter11));
  nor2  gate3079(.a(gate192inter11), .b(gate192inter6), .O(gate192inter12));
  nand2 gate3080(.a(gate192inter12), .b(gate192inter1), .O(G637));
nand2 gate193( .a(G586), .b(G587), .O(G642) );

  xor2  gate2689(.a(G589), .b(G588), .O(gate194inter0));
  nand2 gate2690(.a(gate194inter0), .b(s_306), .O(gate194inter1));
  and2  gate2691(.a(G589), .b(G588), .O(gate194inter2));
  inv1  gate2692(.a(s_306), .O(gate194inter3));
  inv1  gate2693(.a(s_307), .O(gate194inter4));
  nand2 gate2694(.a(gate194inter4), .b(gate194inter3), .O(gate194inter5));
  nor2  gate2695(.a(gate194inter5), .b(gate194inter2), .O(gate194inter6));
  inv1  gate2696(.a(G588), .O(gate194inter7));
  inv1  gate2697(.a(G589), .O(gate194inter8));
  nand2 gate2698(.a(gate194inter8), .b(gate194inter7), .O(gate194inter9));
  nand2 gate2699(.a(s_307), .b(gate194inter3), .O(gate194inter10));
  nor2  gate2700(.a(gate194inter10), .b(gate194inter9), .O(gate194inter11));
  nor2  gate2701(.a(gate194inter11), .b(gate194inter6), .O(gate194inter12));
  nand2 gate2702(.a(gate194inter12), .b(gate194inter1), .O(G645));

  xor2  gate3109(.a(G591), .b(G590), .O(gate195inter0));
  nand2 gate3110(.a(gate195inter0), .b(s_366), .O(gate195inter1));
  and2  gate3111(.a(G591), .b(G590), .O(gate195inter2));
  inv1  gate3112(.a(s_366), .O(gate195inter3));
  inv1  gate3113(.a(s_367), .O(gate195inter4));
  nand2 gate3114(.a(gate195inter4), .b(gate195inter3), .O(gate195inter5));
  nor2  gate3115(.a(gate195inter5), .b(gate195inter2), .O(gate195inter6));
  inv1  gate3116(.a(G590), .O(gate195inter7));
  inv1  gate3117(.a(G591), .O(gate195inter8));
  nand2 gate3118(.a(gate195inter8), .b(gate195inter7), .O(gate195inter9));
  nand2 gate3119(.a(s_367), .b(gate195inter3), .O(gate195inter10));
  nor2  gate3120(.a(gate195inter10), .b(gate195inter9), .O(gate195inter11));
  nor2  gate3121(.a(gate195inter11), .b(gate195inter6), .O(gate195inter12));
  nand2 gate3122(.a(gate195inter12), .b(gate195inter1), .O(G648));

  xor2  gate2549(.a(G593), .b(G592), .O(gate196inter0));
  nand2 gate2550(.a(gate196inter0), .b(s_286), .O(gate196inter1));
  and2  gate2551(.a(G593), .b(G592), .O(gate196inter2));
  inv1  gate2552(.a(s_286), .O(gate196inter3));
  inv1  gate2553(.a(s_287), .O(gate196inter4));
  nand2 gate2554(.a(gate196inter4), .b(gate196inter3), .O(gate196inter5));
  nor2  gate2555(.a(gate196inter5), .b(gate196inter2), .O(gate196inter6));
  inv1  gate2556(.a(G592), .O(gate196inter7));
  inv1  gate2557(.a(G593), .O(gate196inter8));
  nand2 gate2558(.a(gate196inter8), .b(gate196inter7), .O(gate196inter9));
  nand2 gate2559(.a(s_287), .b(gate196inter3), .O(gate196inter10));
  nor2  gate2560(.a(gate196inter10), .b(gate196inter9), .O(gate196inter11));
  nor2  gate2561(.a(gate196inter11), .b(gate196inter6), .O(gate196inter12));
  nand2 gate2562(.a(gate196inter12), .b(gate196inter1), .O(G651));
nand2 gate197( .a(G594), .b(G595), .O(G654) );
nand2 gate198( .a(G596), .b(G597), .O(G657) );
nand2 gate199( .a(G598), .b(G599), .O(G660) );

  xor2  gate1051(.a(G601), .b(G600), .O(gate200inter0));
  nand2 gate1052(.a(gate200inter0), .b(s_72), .O(gate200inter1));
  and2  gate1053(.a(G601), .b(G600), .O(gate200inter2));
  inv1  gate1054(.a(s_72), .O(gate200inter3));
  inv1  gate1055(.a(s_73), .O(gate200inter4));
  nand2 gate1056(.a(gate200inter4), .b(gate200inter3), .O(gate200inter5));
  nor2  gate1057(.a(gate200inter5), .b(gate200inter2), .O(gate200inter6));
  inv1  gate1058(.a(G600), .O(gate200inter7));
  inv1  gate1059(.a(G601), .O(gate200inter8));
  nand2 gate1060(.a(gate200inter8), .b(gate200inter7), .O(gate200inter9));
  nand2 gate1061(.a(s_73), .b(gate200inter3), .O(gate200inter10));
  nor2  gate1062(.a(gate200inter10), .b(gate200inter9), .O(gate200inter11));
  nor2  gate1063(.a(gate200inter11), .b(gate200inter6), .O(gate200inter12));
  nand2 gate1064(.a(gate200inter12), .b(gate200inter1), .O(G663));
nand2 gate201( .a(G602), .b(G607), .O(G666) );
nand2 gate202( .a(G612), .b(G617), .O(G669) );
nand2 gate203( .a(G602), .b(G612), .O(G672) );
nand2 gate204( .a(G607), .b(G617), .O(G675) );

  xor2  gate2185(.a(G627), .b(G622), .O(gate205inter0));
  nand2 gate2186(.a(gate205inter0), .b(s_234), .O(gate205inter1));
  and2  gate2187(.a(G627), .b(G622), .O(gate205inter2));
  inv1  gate2188(.a(s_234), .O(gate205inter3));
  inv1  gate2189(.a(s_235), .O(gate205inter4));
  nand2 gate2190(.a(gate205inter4), .b(gate205inter3), .O(gate205inter5));
  nor2  gate2191(.a(gate205inter5), .b(gate205inter2), .O(gate205inter6));
  inv1  gate2192(.a(G622), .O(gate205inter7));
  inv1  gate2193(.a(G627), .O(gate205inter8));
  nand2 gate2194(.a(gate205inter8), .b(gate205inter7), .O(gate205inter9));
  nand2 gate2195(.a(s_235), .b(gate205inter3), .O(gate205inter10));
  nor2  gate2196(.a(gate205inter10), .b(gate205inter9), .O(gate205inter11));
  nor2  gate2197(.a(gate205inter11), .b(gate205inter6), .O(gate205inter12));
  nand2 gate2198(.a(gate205inter12), .b(gate205inter1), .O(G678));

  xor2  gate2395(.a(G637), .b(G632), .O(gate206inter0));
  nand2 gate2396(.a(gate206inter0), .b(s_264), .O(gate206inter1));
  and2  gate2397(.a(G637), .b(G632), .O(gate206inter2));
  inv1  gate2398(.a(s_264), .O(gate206inter3));
  inv1  gate2399(.a(s_265), .O(gate206inter4));
  nand2 gate2400(.a(gate206inter4), .b(gate206inter3), .O(gate206inter5));
  nor2  gate2401(.a(gate206inter5), .b(gate206inter2), .O(gate206inter6));
  inv1  gate2402(.a(G632), .O(gate206inter7));
  inv1  gate2403(.a(G637), .O(gate206inter8));
  nand2 gate2404(.a(gate206inter8), .b(gate206inter7), .O(gate206inter9));
  nand2 gate2405(.a(s_265), .b(gate206inter3), .O(gate206inter10));
  nor2  gate2406(.a(gate206inter10), .b(gate206inter9), .O(gate206inter11));
  nor2  gate2407(.a(gate206inter11), .b(gate206inter6), .O(gate206inter12));
  nand2 gate2408(.a(gate206inter12), .b(gate206inter1), .O(G681));
nand2 gate207( .a(G622), .b(G632), .O(G684) );

  xor2  gate1275(.a(G637), .b(G627), .O(gate208inter0));
  nand2 gate1276(.a(gate208inter0), .b(s_104), .O(gate208inter1));
  and2  gate1277(.a(G637), .b(G627), .O(gate208inter2));
  inv1  gate1278(.a(s_104), .O(gate208inter3));
  inv1  gate1279(.a(s_105), .O(gate208inter4));
  nand2 gate1280(.a(gate208inter4), .b(gate208inter3), .O(gate208inter5));
  nor2  gate1281(.a(gate208inter5), .b(gate208inter2), .O(gate208inter6));
  inv1  gate1282(.a(G627), .O(gate208inter7));
  inv1  gate1283(.a(G637), .O(gate208inter8));
  nand2 gate1284(.a(gate208inter8), .b(gate208inter7), .O(gate208inter9));
  nand2 gate1285(.a(s_105), .b(gate208inter3), .O(gate208inter10));
  nor2  gate1286(.a(gate208inter10), .b(gate208inter9), .O(gate208inter11));
  nor2  gate1287(.a(gate208inter11), .b(gate208inter6), .O(gate208inter12));
  nand2 gate1288(.a(gate208inter12), .b(gate208inter1), .O(G687));
nand2 gate209( .a(G602), .b(G666), .O(G690) );
nand2 gate210( .a(G607), .b(G666), .O(G691) );

  xor2  gate2717(.a(G669), .b(G612), .O(gate211inter0));
  nand2 gate2718(.a(gate211inter0), .b(s_310), .O(gate211inter1));
  and2  gate2719(.a(G669), .b(G612), .O(gate211inter2));
  inv1  gate2720(.a(s_310), .O(gate211inter3));
  inv1  gate2721(.a(s_311), .O(gate211inter4));
  nand2 gate2722(.a(gate211inter4), .b(gate211inter3), .O(gate211inter5));
  nor2  gate2723(.a(gate211inter5), .b(gate211inter2), .O(gate211inter6));
  inv1  gate2724(.a(G612), .O(gate211inter7));
  inv1  gate2725(.a(G669), .O(gate211inter8));
  nand2 gate2726(.a(gate211inter8), .b(gate211inter7), .O(gate211inter9));
  nand2 gate2727(.a(s_311), .b(gate211inter3), .O(gate211inter10));
  nor2  gate2728(.a(gate211inter10), .b(gate211inter9), .O(gate211inter11));
  nor2  gate2729(.a(gate211inter11), .b(gate211inter6), .O(gate211inter12));
  nand2 gate2730(.a(gate211inter12), .b(gate211inter1), .O(G692));

  xor2  gate1065(.a(G669), .b(G617), .O(gate212inter0));
  nand2 gate1066(.a(gate212inter0), .b(s_74), .O(gate212inter1));
  and2  gate1067(.a(G669), .b(G617), .O(gate212inter2));
  inv1  gate1068(.a(s_74), .O(gate212inter3));
  inv1  gate1069(.a(s_75), .O(gate212inter4));
  nand2 gate1070(.a(gate212inter4), .b(gate212inter3), .O(gate212inter5));
  nor2  gate1071(.a(gate212inter5), .b(gate212inter2), .O(gate212inter6));
  inv1  gate1072(.a(G617), .O(gate212inter7));
  inv1  gate1073(.a(G669), .O(gate212inter8));
  nand2 gate1074(.a(gate212inter8), .b(gate212inter7), .O(gate212inter9));
  nand2 gate1075(.a(s_75), .b(gate212inter3), .O(gate212inter10));
  nor2  gate1076(.a(gate212inter10), .b(gate212inter9), .O(gate212inter11));
  nor2  gate1077(.a(gate212inter11), .b(gate212inter6), .O(gate212inter12));
  nand2 gate1078(.a(gate212inter12), .b(gate212inter1), .O(G693));

  xor2  gate3207(.a(G672), .b(G602), .O(gate213inter0));
  nand2 gate3208(.a(gate213inter0), .b(s_380), .O(gate213inter1));
  and2  gate3209(.a(G672), .b(G602), .O(gate213inter2));
  inv1  gate3210(.a(s_380), .O(gate213inter3));
  inv1  gate3211(.a(s_381), .O(gate213inter4));
  nand2 gate3212(.a(gate213inter4), .b(gate213inter3), .O(gate213inter5));
  nor2  gate3213(.a(gate213inter5), .b(gate213inter2), .O(gate213inter6));
  inv1  gate3214(.a(G602), .O(gate213inter7));
  inv1  gate3215(.a(G672), .O(gate213inter8));
  nand2 gate3216(.a(gate213inter8), .b(gate213inter7), .O(gate213inter9));
  nand2 gate3217(.a(s_381), .b(gate213inter3), .O(gate213inter10));
  nor2  gate3218(.a(gate213inter10), .b(gate213inter9), .O(gate213inter11));
  nor2  gate3219(.a(gate213inter11), .b(gate213inter6), .O(gate213inter12));
  nand2 gate3220(.a(gate213inter12), .b(gate213inter1), .O(G694));

  xor2  gate2857(.a(G672), .b(G612), .O(gate214inter0));
  nand2 gate2858(.a(gate214inter0), .b(s_330), .O(gate214inter1));
  and2  gate2859(.a(G672), .b(G612), .O(gate214inter2));
  inv1  gate2860(.a(s_330), .O(gate214inter3));
  inv1  gate2861(.a(s_331), .O(gate214inter4));
  nand2 gate2862(.a(gate214inter4), .b(gate214inter3), .O(gate214inter5));
  nor2  gate2863(.a(gate214inter5), .b(gate214inter2), .O(gate214inter6));
  inv1  gate2864(.a(G612), .O(gate214inter7));
  inv1  gate2865(.a(G672), .O(gate214inter8));
  nand2 gate2866(.a(gate214inter8), .b(gate214inter7), .O(gate214inter9));
  nand2 gate2867(.a(s_331), .b(gate214inter3), .O(gate214inter10));
  nor2  gate2868(.a(gate214inter10), .b(gate214inter9), .O(gate214inter11));
  nor2  gate2869(.a(gate214inter11), .b(gate214inter6), .O(gate214inter12));
  nand2 gate2870(.a(gate214inter12), .b(gate214inter1), .O(G695));
nand2 gate215( .a(G607), .b(G675), .O(G696) );

  xor2  gate2647(.a(G675), .b(G617), .O(gate216inter0));
  nand2 gate2648(.a(gate216inter0), .b(s_300), .O(gate216inter1));
  and2  gate2649(.a(G675), .b(G617), .O(gate216inter2));
  inv1  gate2650(.a(s_300), .O(gate216inter3));
  inv1  gate2651(.a(s_301), .O(gate216inter4));
  nand2 gate2652(.a(gate216inter4), .b(gate216inter3), .O(gate216inter5));
  nor2  gate2653(.a(gate216inter5), .b(gate216inter2), .O(gate216inter6));
  inv1  gate2654(.a(G617), .O(gate216inter7));
  inv1  gate2655(.a(G675), .O(gate216inter8));
  nand2 gate2656(.a(gate216inter8), .b(gate216inter7), .O(gate216inter9));
  nand2 gate2657(.a(s_301), .b(gate216inter3), .O(gate216inter10));
  nor2  gate2658(.a(gate216inter10), .b(gate216inter9), .O(gate216inter11));
  nor2  gate2659(.a(gate216inter11), .b(gate216inter6), .O(gate216inter12));
  nand2 gate2660(.a(gate216inter12), .b(gate216inter1), .O(G697));
nand2 gate217( .a(G622), .b(G678), .O(G698) );
nand2 gate218( .a(G627), .b(G678), .O(G699) );
nand2 gate219( .a(G632), .b(G681), .O(G700) );
nand2 gate220( .a(G637), .b(G681), .O(G701) );

  xor2  gate1373(.a(G684), .b(G622), .O(gate221inter0));
  nand2 gate1374(.a(gate221inter0), .b(s_118), .O(gate221inter1));
  and2  gate1375(.a(G684), .b(G622), .O(gate221inter2));
  inv1  gate1376(.a(s_118), .O(gate221inter3));
  inv1  gate1377(.a(s_119), .O(gate221inter4));
  nand2 gate1378(.a(gate221inter4), .b(gate221inter3), .O(gate221inter5));
  nor2  gate1379(.a(gate221inter5), .b(gate221inter2), .O(gate221inter6));
  inv1  gate1380(.a(G622), .O(gate221inter7));
  inv1  gate1381(.a(G684), .O(gate221inter8));
  nand2 gate1382(.a(gate221inter8), .b(gate221inter7), .O(gate221inter9));
  nand2 gate1383(.a(s_119), .b(gate221inter3), .O(gate221inter10));
  nor2  gate1384(.a(gate221inter10), .b(gate221inter9), .O(gate221inter11));
  nor2  gate1385(.a(gate221inter11), .b(gate221inter6), .O(gate221inter12));
  nand2 gate1386(.a(gate221inter12), .b(gate221inter1), .O(G702));

  xor2  gate1359(.a(G684), .b(G632), .O(gate222inter0));
  nand2 gate1360(.a(gate222inter0), .b(s_116), .O(gate222inter1));
  and2  gate1361(.a(G684), .b(G632), .O(gate222inter2));
  inv1  gate1362(.a(s_116), .O(gate222inter3));
  inv1  gate1363(.a(s_117), .O(gate222inter4));
  nand2 gate1364(.a(gate222inter4), .b(gate222inter3), .O(gate222inter5));
  nor2  gate1365(.a(gate222inter5), .b(gate222inter2), .O(gate222inter6));
  inv1  gate1366(.a(G632), .O(gate222inter7));
  inv1  gate1367(.a(G684), .O(gate222inter8));
  nand2 gate1368(.a(gate222inter8), .b(gate222inter7), .O(gate222inter9));
  nand2 gate1369(.a(s_117), .b(gate222inter3), .O(gate222inter10));
  nor2  gate1370(.a(gate222inter10), .b(gate222inter9), .O(gate222inter11));
  nor2  gate1371(.a(gate222inter11), .b(gate222inter6), .O(gate222inter12));
  nand2 gate1372(.a(gate222inter12), .b(gate222inter1), .O(G703));

  xor2  gate3039(.a(G687), .b(G627), .O(gate223inter0));
  nand2 gate3040(.a(gate223inter0), .b(s_356), .O(gate223inter1));
  and2  gate3041(.a(G687), .b(G627), .O(gate223inter2));
  inv1  gate3042(.a(s_356), .O(gate223inter3));
  inv1  gate3043(.a(s_357), .O(gate223inter4));
  nand2 gate3044(.a(gate223inter4), .b(gate223inter3), .O(gate223inter5));
  nor2  gate3045(.a(gate223inter5), .b(gate223inter2), .O(gate223inter6));
  inv1  gate3046(.a(G627), .O(gate223inter7));
  inv1  gate3047(.a(G687), .O(gate223inter8));
  nand2 gate3048(.a(gate223inter8), .b(gate223inter7), .O(gate223inter9));
  nand2 gate3049(.a(s_357), .b(gate223inter3), .O(gate223inter10));
  nor2  gate3050(.a(gate223inter10), .b(gate223inter9), .O(gate223inter11));
  nor2  gate3051(.a(gate223inter11), .b(gate223inter6), .O(gate223inter12));
  nand2 gate3052(.a(gate223inter12), .b(gate223inter1), .O(G704));

  xor2  gate2129(.a(G687), .b(G637), .O(gate224inter0));
  nand2 gate2130(.a(gate224inter0), .b(s_226), .O(gate224inter1));
  and2  gate2131(.a(G687), .b(G637), .O(gate224inter2));
  inv1  gate2132(.a(s_226), .O(gate224inter3));
  inv1  gate2133(.a(s_227), .O(gate224inter4));
  nand2 gate2134(.a(gate224inter4), .b(gate224inter3), .O(gate224inter5));
  nor2  gate2135(.a(gate224inter5), .b(gate224inter2), .O(gate224inter6));
  inv1  gate2136(.a(G637), .O(gate224inter7));
  inv1  gate2137(.a(G687), .O(gate224inter8));
  nand2 gate2138(.a(gate224inter8), .b(gate224inter7), .O(gate224inter9));
  nand2 gate2139(.a(s_227), .b(gate224inter3), .O(gate224inter10));
  nor2  gate2140(.a(gate224inter10), .b(gate224inter9), .O(gate224inter11));
  nor2  gate2141(.a(gate224inter11), .b(gate224inter6), .O(gate224inter12));
  nand2 gate2142(.a(gate224inter12), .b(gate224inter1), .O(G705));

  xor2  gate687(.a(G691), .b(G690), .O(gate225inter0));
  nand2 gate688(.a(gate225inter0), .b(s_20), .O(gate225inter1));
  and2  gate689(.a(G691), .b(G690), .O(gate225inter2));
  inv1  gate690(.a(s_20), .O(gate225inter3));
  inv1  gate691(.a(s_21), .O(gate225inter4));
  nand2 gate692(.a(gate225inter4), .b(gate225inter3), .O(gate225inter5));
  nor2  gate693(.a(gate225inter5), .b(gate225inter2), .O(gate225inter6));
  inv1  gate694(.a(G690), .O(gate225inter7));
  inv1  gate695(.a(G691), .O(gate225inter8));
  nand2 gate696(.a(gate225inter8), .b(gate225inter7), .O(gate225inter9));
  nand2 gate697(.a(s_21), .b(gate225inter3), .O(gate225inter10));
  nor2  gate698(.a(gate225inter10), .b(gate225inter9), .O(gate225inter11));
  nor2  gate699(.a(gate225inter11), .b(gate225inter6), .O(gate225inter12));
  nand2 gate700(.a(gate225inter12), .b(gate225inter1), .O(G706));
nand2 gate226( .a(G692), .b(G693), .O(G709) );
nand2 gate227( .a(G694), .b(G695), .O(G712) );

  xor2  gate589(.a(G697), .b(G696), .O(gate228inter0));
  nand2 gate590(.a(gate228inter0), .b(s_6), .O(gate228inter1));
  and2  gate591(.a(G697), .b(G696), .O(gate228inter2));
  inv1  gate592(.a(s_6), .O(gate228inter3));
  inv1  gate593(.a(s_7), .O(gate228inter4));
  nand2 gate594(.a(gate228inter4), .b(gate228inter3), .O(gate228inter5));
  nor2  gate595(.a(gate228inter5), .b(gate228inter2), .O(gate228inter6));
  inv1  gate596(.a(G696), .O(gate228inter7));
  inv1  gate597(.a(G697), .O(gate228inter8));
  nand2 gate598(.a(gate228inter8), .b(gate228inter7), .O(gate228inter9));
  nand2 gate599(.a(s_7), .b(gate228inter3), .O(gate228inter10));
  nor2  gate600(.a(gate228inter10), .b(gate228inter9), .O(gate228inter11));
  nor2  gate601(.a(gate228inter11), .b(gate228inter6), .O(gate228inter12));
  nand2 gate602(.a(gate228inter12), .b(gate228inter1), .O(G715));
nand2 gate229( .a(G698), .b(G699), .O(G718) );
nand2 gate230( .a(G700), .b(G701), .O(G721) );

  xor2  gate855(.a(G703), .b(G702), .O(gate231inter0));
  nand2 gate856(.a(gate231inter0), .b(s_44), .O(gate231inter1));
  and2  gate857(.a(G703), .b(G702), .O(gate231inter2));
  inv1  gate858(.a(s_44), .O(gate231inter3));
  inv1  gate859(.a(s_45), .O(gate231inter4));
  nand2 gate860(.a(gate231inter4), .b(gate231inter3), .O(gate231inter5));
  nor2  gate861(.a(gate231inter5), .b(gate231inter2), .O(gate231inter6));
  inv1  gate862(.a(G702), .O(gate231inter7));
  inv1  gate863(.a(G703), .O(gate231inter8));
  nand2 gate864(.a(gate231inter8), .b(gate231inter7), .O(gate231inter9));
  nand2 gate865(.a(s_45), .b(gate231inter3), .O(gate231inter10));
  nor2  gate866(.a(gate231inter10), .b(gate231inter9), .O(gate231inter11));
  nor2  gate867(.a(gate231inter11), .b(gate231inter6), .O(gate231inter12));
  nand2 gate868(.a(gate231inter12), .b(gate231inter1), .O(G724));

  xor2  gate2451(.a(G705), .b(G704), .O(gate232inter0));
  nand2 gate2452(.a(gate232inter0), .b(s_272), .O(gate232inter1));
  and2  gate2453(.a(G705), .b(G704), .O(gate232inter2));
  inv1  gate2454(.a(s_272), .O(gate232inter3));
  inv1  gate2455(.a(s_273), .O(gate232inter4));
  nand2 gate2456(.a(gate232inter4), .b(gate232inter3), .O(gate232inter5));
  nor2  gate2457(.a(gate232inter5), .b(gate232inter2), .O(gate232inter6));
  inv1  gate2458(.a(G704), .O(gate232inter7));
  inv1  gate2459(.a(G705), .O(gate232inter8));
  nand2 gate2460(.a(gate232inter8), .b(gate232inter7), .O(gate232inter9));
  nand2 gate2461(.a(s_273), .b(gate232inter3), .O(gate232inter10));
  nor2  gate2462(.a(gate232inter10), .b(gate232inter9), .O(gate232inter11));
  nor2  gate2463(.a(gate232inter11), .b(gate232inter6), .O(gate232inter12));
  nand2 gate2464(.a(gate232inter12), .b(gate232inter1), .O(G727));
nand2 gate233( .a(G242), .b(G718), .O(G730) );

  xor2  gate2969(.a(G721), .b(G245), .O(gate234inter0));
  nand2 gate2970(.a(gate234inter0), .b(s_346), .O(gate234inter1));
  and2  gate2971(.a(G721), .b(G245), .O(gate234inter2));
  inv1  gate2972(.a(s_346), .O(gate234inter3));
  inv1  gate2973(.a(s_347), .O(gate234inter4));
  nand2 gate2974(.a(gate234inter4), .b(gate234inter3), .O(gate234inter5));
  nor2  gate2975(.a(gate234inter5), .b(gate234inter2), .O(gate234inter6));
  inv1  gate2976(.a(G245), .O(gate234inter7));
  inv1  gate2977(.a(G721), .O(gate234inter8));
  nand2 gate2978(.a(gate234inter8), .b(gate234inter7), .O(gate234inter9));
  nand2 gate2979(.a(s_347), .b(gate234inter3), .O(gate234inter10));
  nor2  gate2980(.a(gate234inter10), .b(gate234inter9), .O(gate234inter11));
  nor2  gate2981(.a(gate234inter11), .b(gate234inter6), .O(gate234inter12));
  nand2 gate2982(.a(gate234inter12), .b(gate234inter1), .O(G733));

  xor2  gate2955(.a(G724), .b(G248), .O(gate235inter0));
  nand2 gate2956(.a(gate235inter0), .b(s_344), .O(gate235inter1));
  and2  gate2957(.a(G724), .b(G248), .O(gate235inter2));
  inv1  gate2958(.a(s_344), .O(gate235inter3));
  inv1  gate2959(.a(s_345), .O(gate235inter4));
  nand2 gate2960(.a(gate235inter4), .b(gate235inter3), .O(gate235inter5));
  nor2  gate2961(.a(gate235inter5), .b(gate235inter2), .O(gate235inter6));
  inv1  gate2962(.a(G248), .O(gate235inter7));
  inv1  gate2963(.a(G724), .O(gate235inter8));
  nand2 gate2964(.a(gate235inter8), .b(gate235inter7), .O(gate235inter9));
  nand2 gate2965(.a(s_345), .b(gate235inter3), .O(gate235inter10));
  nor2  gate2966(.a(gate235inter10), .b(gate235inter9), .O(gate235inter11));
  nor2  gate2967(.a(gate235inter11), .b(gate235inter6), .O(gate235inter12));
  nand2 gate2968(.a(gate235inter12), .b(gate235inter1), .O(G736));
nand2 gate236( .a(G251), .b(G727), .O(G739) );
nand2 gate237( .a(G254), .b(G706), .O(G742) );
nand2 gate238( .a(G257), .b(G709), .O(G745) );

  xor2  gate3095(.a(G712), .b(G260), .O(gate239inter0));
  nand2 gate3096(.a(gate239inter0), .b(s_364), .O(gate239inter1));
  and2  gate3097(.a(G712), .b(G260), .O(gate239inter2));
  inv1  gate3098(.a(s_364), .O(gate239inter3));
  inv1  gate3099(.a(s_365), .O(gate239inter4));
  nand2 gate3100(.a(gate239inter4), .b(gate239inter3), .O(gate239inter5));
  nor2  gate3101(.a(gate239inter5), .b(gate239inter2), .O(gate239inter6));
  inv1  gate3102(.a(G260), .O(gate239inter7));
  inv1  gate3103(.a(G712), .O(gate239inter8));
  nand2 gate3104(.a(gate239inter8), .b(gate239inter7), .O(gate239inter9));
  nand2 gate3105(.a(s_365), .b(gate239inter3), .O(gate239inter10));
  nor2  gate3106(.a(gate239inter10), .b(gate239inter9), .O(gate239inter11));
  nor2  gate3107(.a(gate239inter11), .b(gate239inter6), .O(gate239inter12));
  nand2 gate3108(.a(gate239inter12), .b(gate239inter1), .O(G748));
nand2 gate240( .a(G263), .b(G715), .O(G751) );

  xor2  gate2213(.a(G730), .b(G242), .O(gate241inter0));
  nand2 gate2214(.a(gate241inter0), .b(s_238), .O(gate241inter1));
  and2  gate2215(.a(G730), .b(G242), .O(gate241inter2));
  inv1  gate2216(.a(s_238), .O(gate241inter3));
  inv1  gate2217(.a(s_239), .O(gate241inter4));
  nand2 gate2218(.a(gate241inter4), .b(gate241inter3), .O(gate241inter5));
  nor2  gate2219(.a(gate241inter5), .b(gate241inter2), .O(gate241inter6));
  inv1  gate2220(.a(G242), .O(gate241inter7));
  inv1  gate2221(.a(G730), .O(gate241inter8));
  nand2 gate2222(.a(gate241inter8), .b(gate241inter7), .O(gate241inter9));
  nand2 gate2223(.a(s_239), .b(gate241inter3), .O(gate241inter10));
  nor2  gate2224(.a(gate241inter10), .b(gate241inter9), .O(gate241inter11));
  nor2  gate2225(.a(gate241inter11), .b(gate241inter6), .O(gate241inter12));
  nand2 gate2226(.a(gate241inter12), .b(gate241inter1), .O(G754));

  xor2  gate897(.a(G730), .b(G718), .O(gate242inter0));
  nand2 gate898(.a(gate242inter0), .b(s_50), .O(gate242inter1));
  and2  gate899(.a(G730), .b(G718), .O(gate242inter2));
  inv1  gate900(.a(s_50), .O(gate242inter3));
  inv1  gate901(.a(s_51), .O(gate242inter4));
  nand2 gate902(.a(gate242inter4), .b(gate242inter3), .O(gate242inter5));
  nor2  gate903(.a(gate242inter5), .b(gate242inter2), .O(gate242inter6));
  inv1  gate904(.a(G718), .O(gate242inter7));
  inv1  gate905(.a(G730), .O(gate242inter8));
  nand2 gate906(.a(gate242inter8), .b(gate242inter7), .O(gate242inter9));
  nand2 gate907(.a(s_51), .b(gate242inter3), .O(gate242inter10));
  nor2  gate908(.a(gate242inter10), .b(gate242inter9), .O(gate242inter11));
  nor2  gate909(.a(gate242inter11), .b(gate242inter6), .O(gate242inter12));
  nand2 gate910(.a(gate242inter12), .b(gate242inter1), .O(G755));

  xor2  gate1639(.a(G733), .b(G245), .O(gate243inter0));
  nand2 gate1640(.a(gate243inter0), .b(s_156), .O(gate243inter1));
  and2  gate1641(.a(G733), .b(G245), .O(gate243inter2));
  inv1  gate1642(.a(s_156), .O(gate243inter3));
  inv1  gate1643(.a(s_157), .O(gate243inter4));
  nand2 gate1644(.a(gate243inter4), .b(gate243inter3), .O(gate243inter5));
  nor2  gate1645(.a(gate243inter5), .b(gate243inter2), .O(gate243inter6));
  inv1  gate1646(.a(G245), .O(gate243inter7));
  inv1  gate1647(.a(G733), .O(gate243inter8));
  nand2 gate1648(.a(gate243inter8), .b(gate243inter7), .O(gate243inter9));
  nand2 gate1649(.a(s_157), .b(gate243inter3), .O(gate243inter10));
  nor2  gate1650(.a(gate243inter10), .b(gate243inter9), .O(gate243inter11));
  nor2  gate1651(.a(gate243inter11), .b(gate243inter6), .O(gate243inter12));
  nand2 gate1652(.a(gate243inter12), .b(gate243inter1), .O(G756));

  xor2  gate2605(.a(G733), .b(G721), .O(gate244inter0));
  nand2 gate2606(.a(gate244inter0), .b(s_294), .O(gate244inter1));
  and2  gate2607(.a(G733), .b(G721), .O(gate244inter2));
  inv1  gate2608(.a(s_294), .O(gate244inter3));
  inv1  gate2609(.a(s_295), .O(gate244inter4));
  nand2 gate2610(.a(gate244inter4), .b(gate244inter3), .O(gate244inter5));
  nor2  gate2611(.a(gate244inter5), .b(gate244inter2), .O(gate244inter6));
  inv1  gate2612(.a(G721), .O(gate244inter7));
  inv1  gate2613(.a(G733), .O(gate244inter8));
  nand2 gate2614(.a(gate244inter8), .b(gate244inter7), .O(gate244inter9));
  nand2 gate2615(.a(s_295), .b(gate244inter3), .O(gate244inter10));
  nor2  gate2616(.a(gate244inter10), .b(gate244inter9), .O(gate244inter11));
  nor2  gate2617(.a(gate244inter11), .b(gate244inter6), .O(gate244inter12));
  nand2 gate2618(.a(gate244inter12), .b(gate244inter1), .O(G757));
nand2 gate245( .a(G248), .b(G736), .O(G758) );
nand2 gate246( .a(G724), .b(G736), .O(G759) );

  xor2  gate2563(.a(G739), .b(G251), .O(gate247inter0));
  nand2 gate2564(.a(gate247inter0), .b(s_288), .O(gate247inter1));
  and2  gate2565(.a(G739), .b(G251), .O(gate247inter2));
  inv1  gate2566(.a(s_288), .O(gate247inter3));
  inv1  gate2567(.a(s_289), .O(gate247inter4));
  nand2 gate2568(.a(gate247inter4), .b(gate247inter3), .O(gate247inter5));
  nor2  gate2569(.a(gate247inter5), .b(gate247inter2), .O(gate247inter6));
  inv1  gate2570(.a(G251), .O(gate247inter7));
  inv1  gate2571(.a(G739), .O(gate247inter8));
  nand2 gate2572(.a(gate247inter8), .b(gate247inter7), .O(gate247inter9));
  nand2 gate2573(.a(s_289), .b(gate247inter3), .O(gate247inter10));
  nor2  gate2574(.a(gate247inter10), .b(gate247inter9), .O(gate247inter11));
  nor2  gate2575(.a(gate247inter11), .b(gate247inter6), .O(gate247inter12));
  nand2 gate2576(.a(gate247inter12), .b(gate247inter1), .O(G760));
nand2 gate248( .a(G727), .b(G739), .O(G761) );

  xor2  gate1471(.a(G742), .b(G254), .O(gate249inter0));
  nand2 gate1472(.a(gate249inter0), .b(s_132), .O(gate249inter1));
  and2  gate1473(.a(G742), .b(G254), .O(gate249inter2));
  inv1  gate1474(.a(s_132), .O(gate249inter3));
  inv1  gate1475(.a(s_133), .O(gate249inter4));
  nand2 gate1476(.a(gate249inter4), .b(gate249inter3), .O(gate249inter5));
  nor2  gate1477(.a(gate249inter5), .b(gate249inter2), .O(gate249inter6));
  inv1  gate1478(.a(G254), .O(gate249inter7));
  inv1  gate1479(.a(G742), .O(gate249inter8));
  nand2 gate1480(.a(gate249inter8), .b(gate249inter7), .O(gate249inter9));
  nand2 gate1481(.a(s_133), .b(gate249inter3), .O(gate249inter10));
  nor2  gate1482(.a(gate249inter10), .b(gate249inter9), .O(gate249inter11));
  nor2  gate1483(.a(gate249inter11), .b(gate249inter6), .O(gate249inter12));
  nand2 gate1484(.a(gate249inter12), .b(gate249inter1), .O(G762));
nand2 gate250( .a(G706), .b(G742), .O(G763) );

  xor2  gate1737(.a(G745), .b(G257), .O(gate251inter0));
  nand2 gate1738(.a(gate251inter0), .b(s_170), .O(gate251inter1));
  and2  gate1739(.a(G745), .b(G257), .O(gate251inter2));
  inv1  gate1740(.a(s_170), .O(gate251inter3));
  inv1  gate1741(.a(s_171), .O(gate251inter4));
  nand2 gate1742(.a(gate251inter4), .b(gate251inter3), .O(gate251inter5));
  nor2  gate1743(.a(gate251inter5), .b(gate251inter2), .O(gate251inter6));
  inv1  gate1744(.a(G257), .O(gate251inter7));
  inv1  gate1745(.a(G745), .O(gate251inter8));
  nand2 gate1746(.a(gate251inter8), .b(gate251inter7), .O(gate251inter9));
  nand2 gate1747(.a(s_171), .b(gate251inter3), .O(gate251inter10));
  nor2  gate1748(.a(gate251inter10), .b(gate251inter9), .O(gate251inter11));
  nor2  gate1749(.a(gate251inter11), .b(gate251inter6), .O(gate251inter12));
  nand2 gate1750(.a(gate251inter12), .b(gate251inter1), .O(G764));
nand2 gate252( .a(G709), .b(G745), .O(G765) );

  xor2  gate547(.a(G748), .b(G260), .O(gate253inter0));
  nand2 gate548(.a(gate253inter0), .b(s_0), .O(gate253inter1));
  and2  gate549(.a(G748), .b(G260), .O(gate253inter2));
  inv1  gate550(.a(s_0), .O(gate253inter3));
  inv1  gate551(.a(s_1), .O(gate253inter4));
  nand2 gate552(.a(gate253inter4), .b(gate253inter3), .O(gate253inter5));
  nor2  gate553(.a(gate253inter5), .b(gate253inter2), .O(gate253inter6));
  inv1  gate554(.a(G260), .O(gate253inter7));
  inv1  gate555(.a(G748), .O(gate253inter8));
  nand2 gate556(.a(gate253inter8), .b(gate253inter7), .O(gate253inter9));
  nand2 gate557(.a(s_1), .b(gate253inter3), .O(gate253inter10));
  nor2  gate558(.a(gate253inter10), .b(gate253inter9), .O(gate253inter11));
  nor2  gate559(.a(gate253inter11), .b(gate253inter6), .O(gate253inter12));
  nand2 gate560(.a(gate253inter12), .b(gate253inter1), .O(G766));

  xor2  gate1219(.a(G748), .b(G712), .O(gate254inter0));
  nand2 gate1220(.a(gate254inter0), .b(s_96), .O(gate254inter1));
  and2  gate1221(.a(G748), .b(G712), .O(gate254inter2));
  inv1  gate1222(.a(s_96), .O(gate254inter3));
  inv1  gate1223(.a(s_97), .O(gate254inter4));
  nand2 gate1224(.a(gate254inter4), .b(gate254inter3), .O(gate254inter5));
  nor2  gate1225(.a(gate254inter5), .b(gate254inter2), .O(gate254inter6));
  inv1  gate1226(.a(G712), .O(gate254inter7));
  inv1  gate1227(.a(G748), .O(gate254inter8));
  nand2 gate1228(.a(gate254inter8), .b(gate254inter7), .O(gate254inter9));
  nand2 gate1229(.a(s_97), .b(gate254inter3), .O(gate254inter10));
  nor2  gate1230(.a(gate254inter10), .b(gate254inter9), .O(gate254inter11));
  nor2  gate1231(.a(gate254inter11), .b(gate254inter6), .O(gate254inter12));
  nand2 gate1232(.a(gate254inter12), .b(gate254inter1), .O(G767));
nand2 gate255( .a(G263), .b(G751), .O(G768) );

  xor2  gate3011(.a(G751), .b(G715), .O(gate256inter0));
  nand2 gate3012(.a(gate256inter0), .b(s_352), .O(gate256inter1));
  and2  gate3013(.a(G751), .b(G715), .O(gate256inter2));
  inv1  gate3014(.a(s_352), .O(gate256inter3));
  inv1  gate3015(.a(s_353), .O(gate256inter4));
  nand2 gate3016(.a(gate256inter4), .b(gate256inter3), .O(gate256inter5));
  nor2  gate3017(.a(gate256inter5), .b(gate256inter2), .O(gate256inter6));
  inv1  gate3018(.a(G715), .O(gate256inter7));
  inv1  gate3019(.a(G751), .O(gate256inter8));
  nand2 gate3020(.a(gate256inter8), .b(gate256inter7), .O(gate256inter9));
  nand2 gate3021(.a(s_353), .b(gate256inter3), .O(gate256inter10));
  nor2  gate3022(.a(gate256inter10), .b(gate256inter9), .O(gate256inter11));
  nor2  gate3023(.a(gate256inter11), .b(gate256inter6), .O(gate256inter12));
  nand2 gate3024(.a(gate256inter12), .b(gate256inter1), .O(G769));
nand2 gate257( .a(G754), .b(G755), .O(G770) );
nand2 gate258( .a(G756), .b(G757), .O(G773) );

  xor2  gate701(.a(G759), .b(G758), .O(gate259inter0));
  nand2 gate702(.a(gate259inter0), .b(s_22), .O(gate259inter1));
  and2  gate703(.a(G759), .b(G758), .O(gate259inter2));
  inv1  gate704(.a(s_22), .O(gate259inter3));
  inv1  gate705(.a(s_23), .O(gate259inter4));
  nand2 gate706(.a(gate259inter4), .b(gate259inter3), .O(gate259inter5));
  nor2  gate707(.a(gate259inter5), .b(gate259inter2), .O(gate259inter6));
  inv1  gate708(.a(G758), .O(gate259inter7));
  inv1  gate709(.a(G759), .O(gate259inter8));
  nand2 gate710(.a(gate259inter8), .b(gate259inter7), .O(gate259inter9));
  nand2 gate711(.a(s_23), .b(gate259inter3), .O(gate259inter10));
  nor2  gate712(.a(gate259inter10), .b(gate259inter9), .O(gate259inter11));
  nor2  gate713(.a(gate259inter11), .b(gate259inter6), .O(gate259inter12));
  nand2 gate714(.a(gate259inter12), .b(gate259inter1), .O(G776));
nand2 gate260( .a(G760), .b(G761), .O(G779) );
nand2 gate261( .a(G762), .b(G763), .O(G782) );
nand2 gate262( .a(G764), .b(G765), .O(G785) );

  xor2  gate2031(.a(G767), .b(G766), .O(gate263inter0));
  nand2 gate2032(.a(gate263inter0), .b(s_212), .O(gate263inter1));
  and2  gate2033(.a(G767), .b(G766), .O(gate263inter2));
  inv1  gate2034(.a(s_212), .O(gate263inter3));
  inv1  gate2035(.a(s_213), .O(gate263inter4));
  nand2 gate2036(.a(gate263inter4), .b(gate263inter3), .O(gate263inter5));
  nor2  gate2037(.a(gate263inter5), .b(gate263inter2), .O(gate263inter6));
  inv1  gate2038(.a(G766), .O(gate263inter7));
  inv1  gate2039(.a(G767), .O(gate263inter8));
  nand2 gate2040(.a(gate263inter8), .b(gate263inter7), .O(gate263inter9));
  nand2 gate2041(.a(s_213), .b(gate263inter3), .O(gate263inter10));
  nor2  gate2042(.a(gate263inter10), .b(gate263inter9), .O(gate263inter11));
  nor2  gate2043(.a(gate263inter11), .b(gate263inter6), .O(gate263inter12));
  nand2 gate2044(.a(gate263inter12), .b(gate263inter1), .O(G788));
nand2 gate264( .a(G768), .b(G769), .O(G791) );
nand2 gate265( .a(G642), .b(G770), .O(G794) );

  xor2  gate869(.a(G773), .b(G645), .O(gate266inter0));
  nand2 gate870(.a(gate266inter0), .b(s_46), .O(gate266inter1));
  and2  gate871(.a(G773), .b(G645), .O(gate266inter2));
  inv1  gate872(.a(s_46), .O(gate266inter3));
  inv1  gate873(.a(s_47), .O(gate266inter4));
  nand2 gate874(.a(gate266inter4), .b(gate266inter3), .O(gate266inter5));
  nor2  gate875(.a(gate266inter5), .b(gate266inter2), .O(gate266inter6));
  inv1  gate876(.a(G645), .O(gate266inter7));
  inv1  gate877(.a(G773), .O(gate266inter8));
  nand2 gate878(.a(gate266inter8), .b(gate266inter7), .O(gate266inter9));
  nand2 gate879(.a(s_47), .b(gate266inter3), .O(gate266inter10));
  nor2  gate880(.a(gate266inter10), .b(gate266inter9), .O(gate266inter11));
  nor2  gate881(.a(gate266inter11), .b(gate266inter6), .O(gate266inter12));
  nand2 gate882(.a(gate266inter12), .b(gate266inter1), .O(G797));
nand2 gate267( .a(G648), .b(G776), .O(G800) );

  xor2  gate1723(.a(G779), .b(G651), .O(gate268inter0));
  nand2 gate1724(.a(gate268inter0), .b(s_168), .O(gate268inter1));
  and2  gate1725(.a(G779), .b(G651), .O(gate268inter2));
  inv1  gate1726(.a(s_168), .O(gate268inter3));
  inv1  gate1727(.a(s_169), .O(gate268inter4));
  nand2 gate1728(.a(gate268inter4), .b(gate268inter3), .O(gate268inter5));
  nor2  gate1729(.a(gate268inter5), .b(gate268inter2), .O(gate268inter6));
  inv1  gate1730(.a(G651), .O(gate268inter7));
  inv1  gate1731(.a(G779), .O(gate268inter8));
  nand2 gate1732(.a(gate268inter8), .b(gate268inter7), .O(gate268inter9));
  nand2 gate1733(.a(s_169), .b(gate268inter3), .O(gate268inter10));
  nor2  gate1734(.a(gate268inter10), .b(gate268inter9), .O(gate268inter11));
  nor2  gate1735(.a(gate268inter11), .b(gate268inter6), .O(gate268inter12));
  nand2 gate1736(.a(gate268inter12), .b(gate268inter1), .O(G803));
nand2 gate269( .a(G654), .b(G782), .O(G806) );

  xor2  gate729(.a(G785), .b(G657), .O(gate270inter0));
  nand2 gate730(.a(gate270inter0), .b(s_26), .O(gate270inter1));
  and2  gate731(.a(G785), .b(G657), .O(gate270inter2));
  inv1  gate732(.a(s_26), .O(gate270inter3));
  inv1  gate733(.a(s_27), .O(gate270inter4));
  nand2 gate734(.a(gate270inter4), .b(gate270inter3), .O(gate270inter5));
  nor2  gate735(.a(gate270inter5), .b(gate270inter2), .O(gate270inter6));
  inv1  gate736(.a(G657), .O(gate270inter7));
  inv1  gate737(.a(G785), .O(gate270inter8));
  nand2 gate738(.a(gate270inter8), .b(gate270inter7), .O(gate270inter9));
  nand2 gate739(.a(s_27), .b(gate270inter3), .O(gate270inter10));
  nor2  gate740(.a(gate270inter10), .b(gate270inter9), .O(gate270inter11));
  nor2  gate741(.a(gate270inter11), .b(gate270inter6), .O(gate270inter12));
  nand2 gate742(.a(gate270inter12), .b(gate270inter1), .O(G809));
nand2 gate271( .a(G660), .b(G788), .O(G812) );

  xor2  gate2465(.a(G791), .b(G663), .O(gate272inter0));
  nand2 gate2466(.a(gate272inter0), .b(s_274), .O(gate272inter1));
  and2  gate2467(.a(G791), .b(G663), .O(gate272inter2));
  inv1  gate2468(.a(s_274), .O(gate272inter3));
  inv1  gate2469(.a(s_275), .O(gate272inter4));
  nand2 gate2470(.a(gate272inter4), .b(gate272inter3), .O(gate272inter5));
  nor2  gate2471(.a(gate272inter5), .b(gate272inter2), .O(gate272inter6));
  inv1  gate2472(.a(G663), .O(gate272inter7));
  inv1  gate2473(.a(G791), .O(gate272inter8));
  nand2 gate2474(.a(gate272inter8), .b(gate272inter7), .O(gate272inter9));
  nand2 gate2475(.a(s_275), .b(gate272inter3), .O(gate272inter10));
  nor2  gate2476(.a(gate272inter10), .b(gate272inter9), .O(gate272inter11));
  nor2  gate2477(.a(gate272inter11), .b(gate272inter6), .O(gate272inter12));
  nand2 gate2478(.a(gate272inter12), .b(gate272inter1), .O(G815));
nand2 gate273( .a(G642), .b(G794), .O(G818) );

  xor2  gate2899(.a(G794), .b(G770), .O(gate274inter0));
  nand2 gate2900(.a(gate274inter0), .b(s_336), .O(gate274inter1));
  and2  gate2901(.a(G794), .b(G770), .O(gate274inter2));
  inv1  gate2902(.a(s_336), .O(gate274inter3));
  inv1  gate2903(.a(s_337), .O(gate274inter4));
  nand2 gate2904(.a(gate274inter4), .b(gate274inter3), .O(gate274inter5));
  nor2  gate2905(.a(gate274inter5), .b(gate274inter2), .O(gate274inter6));
  inv1  gate2906(.a(G770), .O(gate274inter7));
  inv1  gate2907(.a(G794), .O(gate274inter8));
  nand2 gate2908(.a(gate274inter8), .b(gate274inter7), .O(gate274inter9));
  nand2 gate2909(.a(s_337), .b(gate274inter3), .O(gate274inter10));
  nor2  gate2910(.a(gate274inter10), .b(gate274inter9), .O(gate274inter11));
  nor2  gate2911(.a(gate274inter11), .b(gate274inter6), .O(gate274inter12));
  nand2 gate2912(.a(gate274inter12), .b(gate274inter1), .O(G819));
nand2 gate275( .a(G645), .b(G797), .O(G820) );
nand2 gate276( .a(G773), .b(G797), .O(G821) );
nand2 gate277( .a(G648), .b(G800), .O(G822) );
nand2 gate278( .a(G776), .b(G800), .O(G823) );
nand2 gate279( .a(G651), .b(G803), .O(G824) );
nand2 gate280( .a(G779), .b(G803), .O(G825) );
nand2 gate281( .a(G654), .b(G806), .O(G826) );

  xor2  gate1961(.a(G806), .b(G782), .O(gate282inter0));
  nand2 gate1962(.a(gate282inter0), .b(s_202), .O(gate282inter1));
  and2  gate1963(.a(G806), .b(G782), .O(gate282inter2));
  inv1  gate1964(.a(s_202), .O(gate282inter3));
  inv1  gate1965(.a(s_203), .O(gate282inter4));
  nand2 gate1966(.a(gate282inter4), .b(gate282inter3), .O(gate282inter5));
  nor2  gate1967(.a(gate282inter5), .b(gate282inter2), .O(gate282inter6));
  inv1  gate1968(.a(G782), .O(gate282inter7));
  inv1  gate1969(.a(G806), .O(gate282inter8));
  nand2 gate1970(.a(gate282inter8), .b(gate282inter7), .O(gate282inter9));
  nand2 gate1971(.a(s_203), .b(gate282inter3), .O(gate282inter10));
  nor2  gate1972(.a(gate282inter10), .b(gate282inter9), .O(gate282inter11));
  nor2  gate1973(.a(gate282inter11), .b(gate282inter6), .O(gate282inter12));
  nand2 gate1974(.a(gate282inter12), .b(gate282inter1), .O(G827));
nand2 gate283( .a(G657), .b(G809), .O(G828) );

  xor2  gate1709(.a(G809), .b(G785), .O(gate284inter0));
  nand2 gate1710(.a(gate284inter0), .b(s_166), .O(gate284inter1));
  and2  gate1711(.a(G809), .b(G785), .O(gate284inter2));
  inv1  gate1712(.a(s_166), .O(gate284inter3));
  inv1  gate1713(.a(s_167), .O(gate284inter4));
  nand2 gate1714(.a(gate284inter4), .b(gate284inter3), .O(gate284inter5));
  nor2  gate1715(.a(gate284inter5), .b(gate284inter2), .O(gate284inter6));
  inv1  gate1716(.a(G785), .O(gate284inter7));
  inv1  gate1717(.a(G809), .O(gate284inter8));
  nand2 gate1718(.a(gate284inter8), .b(gate284inter7), .O(gate284inter9));
  nand2 gate1719(.a(s_167), .b(gate284inter3), .O(gate284inter10));
  nor2  gate1720(.a(gate284inter10), .b(gate284inter9), .O(gate284inter11));
  nor2  gate1721(.a(gate284inter11), .b(gate284inter6), .O(gate284inter12));
  nand2 gate1722(.a(gate284inter12), .b(gate284inter1), .O(G829));
nand2 gate285( .a(G660), .b(G812), .O(G830) );

  xor2  gate2297(.a(G812), .b(G788), .O(gate286inter0));
  nand2 gate2298(.a(gate286inter0), .b(s_250), .O(gate286inter1));
  and2  gate2299(.a(G812), .b(G788), .O(gate286inter2));
  inv1  gate2300(.a(s_250), .O(gate286inter3));
  inv1  gate2301(.a(s_251), .O(gate286inter4));
  nand2 gate2302(.a(gate286inter4), .b(gate286inter3), .O(gate286inter5));
  nor2  gate2303(.a(gate286inter5), .b(gate286inter2), .O(gate286inter6));
  inv1  gate2304(.a(G788), .O(gate286inter7));
  inv1  gate2305(.a(G812), .O(gate286inter8));
  nand2 gate2306(.a(gate286inter8), .b(gate286inter7), .O(gate286inter9));
  nand2 gate2307(.a(s_251), .b(gate286inter3), .O(gate286inter10));
  nor2  gate2308(.a(gate286inter10), .b(gate286inter9), .O(gate286inter11));
  nor2  gate2309(.a(gate286inter11), .b(gate286inter6), .O(gate286inter12));
  nand2 gate2310(.a(gate286inter12), .b(gate286inter1), .O(G831));

  xor2  gate1485(.a(G815), .b(G663), .O(gate287inter0));
  nand2 gate1486(.a(gate287inter0), .b(s_134), .O(gate287inter1));
  and2  gate1487(.a(G815), .b(G663), .O(gate287inter2));
  inv1  gate1488(.a(s_134), .O(gate287inter3));
  inv1  gate1489(.a(s_135), .O(gate287inter4));
  nand2 gate1490(.a(gate287inter4), .b(gate287inter3), .O(gate287inter5));
  nor2  gate1491(.a(gate287inter5), .b(gate287inter2), .O(gate287inter6));
  inv1  gate1492(.a(G663), .O(gate287inter7));
  inv1  gate1493(.a(G815), .O(gate287inter8));
  nand2 gate1494(.a(gate287inter8), .b(gate287inter7), .O(gate287inter9));
  nand2 gate1495(.a(s_135), .b(gate287inter3), .O(gate287inter10));
  nor2  gate1496(.a(gate287inter10), .b(gate287inter9), .O(gate287inter11));
  nor2  gate1497(.a(gate287inter11), .b(gate287inter6), .O(gate287inter12));
  nand2 gate1498(.a(gate287inter12), .b(gate287inter1), .O(G832));
nand2 gate288( .a(G791), .b(G815), .O(G833) );
nand2 gate289( .a(G818), .b(G819), .O(G834) );

  xor2  gate1695(.a(G821), .b(G820), .O(gate290inter0));
  nand2 gate1696(.a(gate290inter0), .b(s_164), .O(gate290inter1));
  and2  gate1697(.a(G821), .b(G820), .O(gate290inter2));
  inv1  gate1698(.a(s_164), .O(gate290inter3));
  inv1  gate1699(.a(s_165), .O(gate290inter4));
  nand2 gate1700(.a(gate290inter4), .b(gate290inter3), .O(gate290inter5));
  nor2  gate1701(.a(gate290inter5), .b(gate290inter2), .O(gate290inter6));
  inv1  gate1702(.a(G820), .O(gate290inter7));
  inv1  gate1703(.a(G821), .O(gate290inter8));
  nand2 gate1704(.a(gate290inter8), .b(gate290inter7), .O(gate290inter9));
  nand2 gate1705(.a(s_165), .b(gate290inter3), .O(gate290inter10));
  nor2  gate1706(.a(gate290inter10), .b(gate290inter9), .O(gate290inter11));
  nor2  gate1707(.a(gate290inter11), .b(gate290inter6), .O(gate290inter12));
  nand2 gate1708(.a(gate290inter12), .b(gate290inter1), .O(G847));
nand2 gate291( .a(G822), .b(G823), .O(G860) );

  xor2  gate743(.a(G825), .b(G824), .O(gate292inter0));
  nand2 gate744(.a(gate292inter0), .b(s_28), .O(gate292inter1));
  and2  gate745(.a(G825), .b(G824), .O(gate292inter2));
  inv1  gate746(.a(s_28), .O(gate292inter3));
  inv1  gate747(.a(s_29), .O(gate292inter4));
  nand2 gate748(.a(gate292inter4), .b(gate292inter3), .O(gate292inter5));
  nor2  gate749(.a(gate292inter5), .b(gate292inter2), .O(gate292inter6));
  inv1  gate750(.a(G824), .O(gate292inter7));
  inv1  gate751(.a(G825), .O(gate292inter8));
  nand2 gate752(.a(gate292inter8), .b(gate292inter7), .O(gate292inter9));
  nand2 gate753(.a(s_29), .b(gate292inter3), .O(gate292inter10));
  nor2  gate754(.a(gate292inter10), .b(gate292inter9), .O(gate292inter11));
  nor2  gate755(.a(gate292inter11), .b(gate292inter6), .O(gate292inter12));
  nand2 gate756(.a(gate292inter12), .b(gate292inter1), .O(G873));
nand2 gate293( .a(G828), .b(G829), .O(G886) );
nand2 gate294( .a(G832), .b(G833), .O(G899) );
nand2 gate295( .a(G830), .b(G831), .O(G912) );

  xor2  gate3179(.a(G827), .b(G826), .O(gate296inter0));
  nand2 gate3180(.a(gate296inter0), .b(s_376), .O(gate296inter1));
  and2  gate3181(.a(G827), .b(G826), .O(gate296inter2));
  inv1  gate3182(.a(s_376), .O(gate296inter3));
  inv1  gate3183(.a(s_377), .O(gate296inter4));
  nand2 gate3184(.a(gate296inter4), .b(gate296inter3), .O(gate296inter5));
  nor2  gate3185(.a(gate296inter5), .b(gate296inter2), .O(gate296inter6));
  inv1  gate3186(.a(G826), .O(gate296inter7));
  inv1  gate3187(.a(G827), .O(gate296inter8));
  nand2 gate3188(.a(gate296inter8), .b(gate296inter7), .O(gate296inter9));
  nand2 gate3189(.a(s_377), .b(gate296inter3), .O(gate296inter10));
  nor2  gate3190(.a(gate296inter10), .b(gate296inter9), .O(gate296inter11));
  nor2  gate3191(.a(gate296inter11), .b(gate296inter6), .O(gate296inter12));
  nand2 gate3192(.a(gate296inter12), .b(gate296inter1), .O(G925));
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );
nand2 gate387( .a(G1), .b(G1036), .O(G1132) );

  xor2  gate2885(.a(G1039), .b(G2), .O(gate388inter0));
  nand2 gate2886(.a(gate388inter0), .b(s_334), .O(gate388inter1));
  and2  gate2887(.a(G1039), .b(G2), .O(gate388inter2));
  inv1  gate2888(.a(s_334), .O(gate388inter3));
  inv1  gate2889(.a(s_335), .O(gate388inter4));
  nand2 gate2890(.a(gate388inter4), .b(gate388inter3), .O(gate388inter5));
  nor2  gate2891(.a(gate388inter5), .b(gate388inter2), .O(gate388inter6));
  inv1  gate2892(.a(G2), .O(gate388inter7));
  inv1  gate2893(.a(G1039), .O(gate388inter8));
  nand2 gate2894(.a(gate388inter8), .b(gate388inter7), .O(gate388inter9));
  nand2 gate2895(.a(s_335), .b(gate388inter3), .O(gate388inter10));
  nor2  gate2896(.a(gate388inter10), .b(gate388inter9), .O(gate388inter11));
  nor2  gate2897(.a(gate388inter11), .b(gate388inter6), .O(gate388inter12));
  nand2 gate2898(.a(gate388inter12), .b(gate388inter1), .O(G1135));
nand2 gate389( .a(G3), .b(G1042), .O(G1138) );
nand2 gate390( .a(G4), .b(G1045), .O(G1141) );
nand2 gate391( .a(G5), .b(G1048), .O(G1144) );
nand2 gate392( .a(G6), .b(G1051), .O(G1147) );
nand2 gate393( .a(G7), .b(G1054), .O(G1150) );
nand2 gate394( .a(G8), .b(G1057), .O(G1153) );

  xor2  gate1821(.a(G1060), .b(G9), .O(gate395inter0));
  nand2 gate1822(.a(gate395inter0), .b(s_182), .O(gate395inter1));
  and2  gate1823(.a(G1060), .b(G9), .O(gate395inter2));
  inv1  gate1824(.a(s_182), .O(gate395inter3));
  inv1  gate1825(.a(s_183), .O(gate395inter4));
  nand2 gate1826(.a(gate395inter4), .b(gate395inter3), .O(gate395inter5));
  nor2  gate1827(.a(gate395inter5), .b(gate395inter2), .O(gate395inter6));
  inv1  gate1828(.a(G9), .O(gate395inter7));
  inv1  gate1829(.a(G1060), .O(gate395inter8));
  nand2 gate1830(.a(gate395inter8), .b(gate395inter7), .O(gate395inter9));
  nand2 gate1831(.a(s_183), .b(gate395inter3), .O(gate395inter10));
  nor2  gate1832(.a(gate395inter10), .b(gate395inter9), .O(gate395inter11));
  nor2  gate1833(.a(gate395inter11), .b(gate395inter6), .O(gate395inter12));
  nand2 gate1834(.a(gate395inter12), .b(gate395inter1), .O(G1156));
nand2 gate396( .a(G10), .b(G1063), .O(G1159) );
nand2 gate397( .a(G11), .b(G1066), .O(G1162) );

  xor2  gate2003(.a(G1069), .b(G12), .O(gate398inter0));
  nand2 gate2004(.a(gate398inter0), .b(s_208), .O(gate398inter1));
  and2  gate2005(.a(G1069), .b(G12), .O(gate398inter2));
  inv1  gate2006(.a(s_208), .O(gate398inter3));
  inv1  gate2007(.a(s_209), .O(gate398inter4));
  nand2 gate2008(.a(gate398inter4), .b(gate398inter3), .O(gate398inter5));
  nor2  gate2009(.a(gate398inter5), .b(gate398inter2), .O(gate398inter6));
  inv1  gate2010(.a(G12), .O(gate398inter7));
  inv1  gate2011(.a(G1069), .O(gate398inter8));
  nand2 gate2012(.a(gate398inter8), .b(gate398inter7), .O(gate398inter9));
  nand2 gate2013(.a(s_209), .b(gate398inter3), .O(gate398inter10));
  nor2  gate2014(.a(gate398inter10), .b(gate398inter9), .O(gate398inter11));
  nor2  gate2015(.a(gate398inter11), .b(gate398inter6), .O(gate398inter12));
  nand2 gate2016(.a(gate398inter12), .b(gate398inter1), .O(G1165));
nand2 gate399( .a(G13), .b(G1072), .O(G1168) );
nand2 gate400( .a(G14), .b(G1075), .O(G1171) );
nand2 gate401( .a(G15), .b(G1078), .O(G1174) );

  xor2  gate1401(.a(G1081), .b(G16), .O(gate402inter0));
  nand2 gate1402(.a(gate402inter0), .b(s_122), .O(gate402inter1));
  and2  gate1403(.a(G1081), .b(G16), .O(gate402inter2));
  inv1  gate1404(.a(s_122), .O(gate402inter3));
  inv1  gate1405(.a(s_123), .O(gate402inter4));
  nand2 gate1406(.a(gate402inter4), .b(gate402inter3), .O(gate402inter5));
  nor2  gate1407(.a(gate402inter5), .b(gate402inter2), .O(gate402inter6));
  inv1  gate1408(.a(G16), .O(gate402inter7));
  inv1  gate1409(.a(G1081), .O(gate402inter8));
  nand2 gate1410(.a(gate402inter8), .b(gate402inter7), .O(gate402inter9));
  nand2 gate1411(.a(s_123), .b(gate402inter3), .O(gate402inter10));
  nor2  gate1412(.a(gate402inter10), .b(gate402inter9), .O(gate402inter11));
  nor2  gate1413(.a(gate402inter11), .b(gate402inter6), .O(gate402inter12));
  nand2 gate1414(.a(gate402inter12), .b(gate402inter1), .O(G1177));

  xor2  gate2381(.a(G1084), .b(G17), .O(gate403inter0));
  nand2 gate2382(.a(gate403inter0), .b(s_262), .O(gate403inter1));
  and2  gate2383(.a(G1084), .b(G17), .O(gate403inter2));
  inv1  gate2384(.a(s_262), .O(gate403inter3));
  inv1  gate2385(.a(s_263), .O(gate403inter4));
  nand2 gate2386(.a(gate403inter4), .b(gate403inter3), .O(gate403inter5));
  nor2  gate2387(.a(gate403inter5), .b(gate403inter2), .O(gate403inter6));
  inv1  gate2388(.a(G17), .O(gate403inter7));
  inv1  gate2389(.a(G1084), .O(gate403inter8));
  nand2 gate2390(.a(gate403inter8), .b(gate403inter7), .O(gate403inter9));
  nand2 gate2391(.a(s_263), .b(gate403inter3), .O(gate403inter10));
  nor2  gate2392(.a(gate403inter10), .b(gate403inter9), .O(gate403inter11));
  nor2  gate2393(.a(gate403inter11), .b(gate403inter6), .O(gate403inter12));
  nand2 gate2394(.a(gate403inter12), .b(gate403inter1), .O(G1180));
nand2 gate404( .a(G18), .b(G1087), .O(G1183) );
nand2 gate405( .a(G19), .b(G1090), .O(G1186) );

  xor2  gate1611(.a(G1093), .b(G20), .O(gate406inter0));
  nand2 gate1612(.a(gate406inter0), .b(s_152), .O(gate406inter1));
  and2  gate1613(.a(G1093), .b(G20), .O(gate406inter2));
  inv1  gate1614(.a(s_152), .O(gate406inter3));
  inv1  gate1615(.a(s_153), .O(gate406inter4));
  nand2 gate1616(.a(gate406inter4), .b(gate406inter3), .O(gate406inter5));
  nor2  gate1617(.a(gate406inter5), .b(gate406inter2), .O(gate406inter6));
  inv1  gate1618(.a(G20), .O(gate406inter7));
  inv1  gate1619(.a(G1093), .O(gate406inter8));
  nand2 gate1620(.a(gate406inter8), .b(gate406inter7), .O(gate406inter9));
  nand2 gate1621(.a(s_153), .b(gate406inter3), .O(gate406inter10));
  nor2  gate1622(.a(gate406inter10), .b(gate406inter9), .O(gate406inter11));
  nor2  gate1623(.a(gate406inter11), .b(gate406inter6), .O(gate406inter12));
  nand2 gate1624(.a(gate406inter12), .b(gate406inter1), .O(G1189));

  xor2  gate1037(.a(G1096), .b(G21), .O(gate407inter0));
  nand2 gate1038(.a(gate407inter0), .b(s_70), .O(gate407inter1));
  and2  gate1039(.a(G1096), .b(G21), .O(gate407inter2));
  inv1  gate1040(.a(s_70), .O(gate407inter3));
  inv1  gate1041(.a(s_71), .O(gate407inter4));
  nand2 gate1042(.a(gate407inter4), .b(gate407inter3), .O(gate407inter5));
  nor2  gate1043(.a(gate407inter5), .b(gate407inter2), .O(gate407inter6));
  inv1  gate1044(.a(G21), .O(gate407inter7));
  inv1  gate1045(.a(G1096), .O(gate407inter8));
  nand2 gate1046(.a(gate407inter8), .b(gate407inter7), .O(gate407inter9));
  nand2 gate1047(.a(s_71), .b(gate407inter3), .O(gate407inter10));
  nor2  gate1048(.a(gate407inter10), .b(gate407inter9), .O(gate407inter11));
  nor2  gate1049(.a(gate407inter11), .b(gate407inter6), .O(gate407inter12));
  nand2 gate1050(.a(gate407inter12), .b(gate407inter1), .O(G1192));
nand2 gate408( .a(G22), .b(G1099), .O(G1195) );

  xor2  gate1751(.a(G1102), .b(G23), .O(gate409inter0));
  nand2 gate1752(.a(gate409inter0), .b(s_172), .O(gate409inter1));
  and2  gate1753(.a(G1102), .b(G23), .O(gate409inter2));
  inv1  gate1754(.a(s_172), .O(gate409inter3));
  inv1  gate1755(.a(s_173), .O(gate409inter4));
  nand2 gate1756(.a(gate409inter4), .b(gate409inter3), .O(gate409inter5));
  nor2  gate1757(.a(gate409inter5), .b(gate409inter2), .O(gate409inter6));
  inv1  gate1758(.a(G23), .O(gate409inter7));
  inv1  gate1759(.a(G1102), .O(gate409inter8));
  nand2 gate1760(.a(gate409inter8), .b(gate409inter7), .O(gate409inter9));
  nand2 gate1761(.a(s_173), .b(gate409inter3), .O(gate409inter10));
  nor2  gate1762(.a(gate409inter10), .b(gate409inter9), .O(gate409inter11));
  nor2  gate1763(.a(gate409inter11), .b(gate409inter6), .O(gate409inter12));
  nand2 gate1764(.a(gate409inter12), .b(gate409inter1), .O(G1198));

  xor2  gate1513(.a(G1105), .b(G24), .O(gate410inter0));
  nand2 gate1514(.a(gate410inter0), .b(s_138), .O(gate410inter1));
  and2  gate1515(.a(G1105), .b(G24), .O(gate410inter2));
  inv1  gate1516(.a(s_138), .O(gate410inter3));
  inv1  gate1517(.a(s_139), .O(gate410inter4));
  nand2 gate1518(.a(gate410inter4), .b(gate410inter3), .O(gate410inter5));
  nor2  gate1519(.a(gate410inter5), .b(gate410inter2), .O(gate410inter6));
  inv1  gate1520(.a(G24), .O(gate410inter7));
  inv1  gate1521(.a(G1105), .O(gate410inter8));
  nand2 gate1522(.a(gate410inter8), .b(gate410inter7), .O(gate410inter9));
  nand2 gate1523(.a(s_139), .b(gate410inter3), .O(gate410inter10));
  nor2  gate1524(.a(gate410inter10), .b(gate410inter9), .O(gate410inter11));
  nor2  gate1525(.a(gate410inter11), .b(gate410inter6), .O(gate410inter12));
  nand2 gate1526(.a(gate410inter12), .b(gate410inter1), .O(G1201));
nand2 gate411( .a(G25), .b(G1108), .O(G1204) );

  xor2  gate2913(.a(G1111), .b(G26), .O(gate412inter0));
  nand2 gate2914(.a(gate412inter0), .b(s_338), .O(gate412inter1));
  and2  gate2915(.a(G1111), .b(G26), .O(gate412inter2));
  inv1  gate2916(.a(s_338), .O(gate412inter3));
  inv1  gate2917(.a(s_339), .O(gate412inter4));
  nand2 gate2918(.a(gate412inter4), .b(gate412inter3), .O(gate412inter5));
  nor2  gate2919(.a(gate412inter5), .b(gate412inter2), .O(gate412inter6));
  inv1  gate2920(.a(G26), .O(gate412inter7));
  inv1  gate2921(.a(G1111), .O(gate412inter8));
  nand2 gate2922(.a(gate412inter8), .b(gate412inter7), .O(gate412inter9));
  nand2 gate2923(.a(s_339), .b(gate412inter3), .O(gate412inter10));
  nor2  gate2924(.a(gate412inter10), .b(gate412inter9), .O(gate412inter11));
  nor2  gate2925(.a(gate412inter11), .b(gate412inter6), .O(gate412inter12));
  nand2 gate2926(.a(gate412inter12), .b(gate412inter1), .O(G1207));
nand2 gate413( .a(G27), .b(G1114), .O(G1210) );

  xor2  gate1163(.a(G1117), .b(G28), .O(gate414inter0));
  nand2 gate1164(.a(gate414inter0), .b(s_88), .O(gate414inter1));
  and2  gate1165(.a(G1117), .b(G28), .O(gate414inter2));
  inv1  gate1166(.a(s_88), .O(gate414inter3));
  inv1  gate1167(.a(s_89), .O(gate414inter4));
  nand2 gate1168(.a(gate414inter4), .b(gate414inter3), .O(gate414inter5));
  nor2  gate1169(.a(gate414inter5), .b(gate414inter2), .O(gate414inter6));
  inv1  gate1170(.a(G28), .O(gate414inter7));
  inv1  gate1171(.a(G1117), .O(gate414inter8));
  nand2 gate1172(.a(gate414inter8), .b(gate414inter7), .O(gate414inter9));
  nand2 gate1173(.a(s_89), .b(gate414inter3), .O(gate414inter10));
  nor2  gate1174(.a(gate414inter10), .b(gate414inter9), .O(gate414inter11));
  nor2  gate1175(.a(gate414inter11), .b(gate414inter6), .O(gate414inter12));
  nand2 gate1176(.a(gate414inter12), .b(gate414inter1), .O(G1213));
nand2 gate415( .a(G29), .b(G1120), .O(G1216) );
nand2 gate416( .a(G30), .b(G1123), .O(G1219) );
nand2 gate417( .a(G31), .b(G1126), .O(G1222) );
nand2 gate418( .a(G32), .b(G1129), .O(G1225) );

  xor2  gate1849(.a(G1132), .b(G1), .O(gate419inter0));
  nand2 gate1850(.a(gate419inter0), .b(s_186), .O(gate419inter1));
  and2  gate1851(.a(G1132), .b(G1), .O(gate419inter2));
  inv1  gate1852(.a(s_186), .O(gate419inter3));
  inv1  gate1853(.a(s_187), .O(gate419inter4));
  nand2 gate1854(.a(gate419inter4), .b(gate419inter3), .O(gate419inter5));
  nor2  gate1855(.a(gate419inter5), .b(gate419inter2), .O(gate419inter6));
  inv1  gate1856(.a(G1), .O(gate419inter7));
  inv1  gate1857(.a(G1132), .O(gate419inter8));
  nand2 gate1858(.a(gate419inter8), .b(gate419inter7), .O(gate419inter9));
  nand2 gate1859(.a(s_187), .b(gate419inter3), .O(gate419inter10));
  nor2  gate1860(.a(gate419inter10), .b(gate419inter9), .O(gate419inter11));
  nor2  gate1861(.a(gate419inter11), .b(gate419inter6), .O(gate419inter12));
  nand2 gate1862(.a(gate419inter12), .b(gate419inter1), .O(G1228));
nand2 gate420( .a(G1036), .b(G1132), .O(G1229) );

  xor2  gate1205(.a(G1135), .b(G2), .O(gate421inter0));
  nand2 gate1206(.a(gate421inter0), .b(s_94), .O(gate421inter1));
  and2  gate1207(.a(G1135), .b(G2), .O(gate421inter2));
  inv1  gate1208(.a(s_94), .O(gate421inter3));
  inv1  gate1209(.a(s_95), .O(gate421inter4));
  nand2 gate1210(.a(gate421inter4), .b(gate421inter3), .O(gate421inter5));
  nor2  gate1211(.a(gate421inter5), .b(gate421inter2), .O(gate421inter6));
  inv1  gate1212(.a(G2), .O(gate421inter7));
  inv1  gate1213(.a(G1135), .O(gate421inter8));
  nand2 gate1214(.a(gate421inter8), .b(gate421inter7), .O(gate421inter9));
  nand2 gate1215(.a(s_95), .b(gate421inter3), .O(gate421inter10));
  nor2  gate1216(.a(gate421inter10), .b(gate421inter9), .O(gate421inter11));
  nor2  gate1217(.a(gate421inter11), .b(gate421inter6), .O(gate421inter12));
  nand2 gate1218(.a(gate421inter12), .b(gate421inter1), .O(G1230));

  xor2  gate1023(.a(G1135), .b(G1039), .O(gate422inter0));
  nand2 gate1024(.a(gate422inter0), .b(s_68), .O(gate422inter1));
  and2  gate1025(.a(G1135), .b(G1039), .O(gate422inter2));
  inv1  gate1026(.a(s_68), .O(gate422inter3));
  inv1  gate1027(.a(s_69), .O(gate422inter4));
  nand2 gate1028(.a(gate422inter4), .b(gate422inter3), .O(gate422inter5));
  nor2  gate1029(.a(gate422inter5), .b(gate422inter2), .O(gate422inter6));
  inv1  gate1030(.a(G1039), .O(gate422inter7));
  inv1  gate1031(.a(G1135), .O(gate422inter8));
  nand2 gate1032(.a(gate422inter8), .b(gate422inter7), .O(gate422inter9));
  nand2 gate1033(.a(s_69), .b(gate422inter3), .O(gate422inter10));
  nor2  gate1034(.a(gate422inter10), .b(gate422inter9), .O(gate422inter11));
  nor2  gate1035(.a(gate422inter11), .b(gate422inter6), .O(gate422inter12));
  nand2 gate1036(.a(gate422inter12), .b(gate422inter1), .O(G1231));
nand2 gate423( .a(G3), .b(G1138), .O(G1232) );

  xor2  gate799(.a(G1138), .b(G1042), .O(gate424inter0));
  nand2 gate800(.a(gate424inter0), .b(s_36), .O(gate424inter1));
  and2  gate801(.a(G1138), .b(G1042), .O(gate424inter2));
  inv1  gate802(.a(s_36), .O(gate424inter3));
  inv1  gate803(.a(s_37), .O(gate424inter4));
  nand2 gate804(.a(gate424inter4), .b(gate424inter3), .O(gate424inter5));
  nor2  gate805(.a(gate424inter5), .b(gate424inter2), .O(gate424inter6));
  inv1  gate806(.a(G1042), .O(gate424inter7));
  inv1  gate807(.a(G1138), .O(gate424inter8));
  nand2 gate808(.a(gate424inter8), .b(gate424inter7), .O(gate424inter9));
  nand2 gate809(.a(s_37), .b(gate424inter3), .O(gate424inter10));
  nor2  gate810(.a(gate424inter10), .b(gate424inter9), .O(gate424inter11));
  nor2  gate811(.a(gate424inter11), .b(gate424inter6), .O(gate424inter12));
  nand2 gate812(.a(gate424inter12), .b(gate424inter1), .O(G1233));
nand2 gate425( .a(G4), .b(G1141), .O(G1234) );
nand2 gate426( .a(G1045), .b(G1141), .O(G1235) );

  xor2  gate827(.a(G1144), .b(G5), .O(gate427inter0));
  nand2 gate828(.a(gate427inter0), .b(s_40), .O(gate427inter1));
  and2  gate829(.a(G1144), .b(G5), .O(gate427inter2));
  inv1  gate830(.a(s_40), .O(gate427inter3));
  inv1  gate831(.a(s_41), .O(gate427inter4));
  nand2 gate832(.a(gate427inter4), .b(gate427inter3), .O(gate427inter5));
  nor2  gate833(.a(gate427inter5), .b(gate427inter2), .O(gate427inter6));
  inv1  gate834(.a(G5), .O(gate427inter7));
  inv1  gate835(.a(G1144), .O(gate427inter8));
  nand2 gate836(.a(gate427inter8), .b(gate427inter7), .O(gate427inter9));
  nand2 gate837(.a(s_41), .b(gate427inter3), .O(gate427inter10));
  nor2  gate838(.a(gate427inter10), .b(gate427inter9), .O(gate427inter11));
  nor2  gate839(.a(gate427inter11), .b(gate427inter6), .O(gate427inter12));
  nand2 gate840(.a(gate427inter12), .b(gate427inter1), .O(G1236));
nand2 gate428( .a(G1048), .b(G1144), .O(G1237) );
nand2 gate429( .a(G6), .b(G1147), .O(G1238) );
nand2 gate430( .a(G1051), .b(G1147), .O(G1239) );
nand2 gate431( .a(G7), .b(G1150), .O(G1240) );
nand2 gate432( .a(G1054), .b(G1150), .O(G1241) );

  xor2  gate1191(.a(G1153), .b(G8), .O(gate433inter0));
  nand2 gate1192(.a(gate433inter0), .b(s_92), .O(gate433inter1));
  and2  gate1193(.a(G1153), .b(G8), .O(gate433inter2));
  inv1  gate1194(.a(s_92), .O(gate433inter3));
  inv1  gate1195(.a(s_93), .O(gate433inter4));
  nand2 gate1196(.a(gate433inter4), .b(gate433inter3), .O(gate433inter5));
  nor2  gate1197(.a(gate433inter5), .b(gate433inter2), .O(gate433inter6));
  inv1  gate1198(.a(G8), .O(gate433inter7));
  inv1  gate1199(.a(G1153), .O(gate433inter8));
  nand2 gate1200(.a(gate433inter8), .b(gate433inter7), .O(gate433inter9));
  nand2 gate1201(.a(s_93), .b(gate433inter3), .O(gate433inter10));
  nor2  gate1202(.a(gate433inter10), .b(gate433inter9), .O(gate433inter11));
  nor2  gate1203(.a(gate433inter11), .b(gate433inter6), .O(gate433inter12));
  nand2 gate1204(.a(gate433inter12), .b(gate433inter1), .O(G1242));
nand2 gate434( .a(G1057), .b(G1153), .O(G1243) );

  xor2  gate1079(.a(G1156), .b(G9), .O(gate435inter0));
  nand2 gate1080(.a(gate435inter0), .b(s_76), .O(gate435inter1));
  and2  gate1081(.a(G1156), .b(G9), .O(gate435inter2));
  inv1  gate1082(.a(s_76), .O(gate435inter3));
  inv1  gate1083(.a(s_77), .O(gate435inter4));
  nand2 gate1084(.a(gate435inter4), .b(gate435inter3), .O(gate435inter5));
  nor2  gate1085(.a(gate435inter5), .b(gate435inter2), .O(gate435inter6));
  inv1  gate1086(.a(G9), .O(gate435inter7));
  inv1  gate1087(.a(G1156), .O(gate435inter8));
  nand2 gate1088(.a(gate435inter8), .b(gate435inter7), .O(gate435inter9));
  nand2 gate1089(.a(s_77), .b(gate435inter3), .O(gate435inter10));
  nor2  gate1090(.a(gate435inter10), .b(gate435inter9), .O(gate435inter11));
  nor2  gate1091(.a(gate435inter11), .b(gate435inter6), .O(gate435inter12));
  nand2 gate1092(.a(gate435inter12), .b(gate435inter1), .O(G1244));

  xor2  gate1807(.a(G1156), .b(G1060), .O(gate436inter0));
  nand2 gate1808(.a(gate436inter0), .b(s_180), .O(gate436inter1));
  and2  gate1809(.a(G1156), .b(G1060), .O(gate436inter2));
  inv1  gate1810(.a(s_180), .O(gate436inter3));
  inv1  gate1811(.a(s_181), .O(gate436inter4));
  nand2 gate1812(.a(gate436inter4), .b(gate436inter3), .O(gate436inter5));
  nor2  gate1813(.a(gate436inter5), .b(gate436inter2), .O(gate436inter6));
  inv1  gate1814(.a(G1060), .O(gate436inter7));
  inv1  gate1815(.a(G1156), .O(gate436inter8));
  nand2 gate1816(.a(gate436inter8), .b(gate436inter7), .O(gate436inter9));
  nand2 gate1817(.a(s_181), .b(gate436inter3), .O(gate436inter10));
  nor2  gate1818(.a(gate436inter10), .b(gate436inter9), .O(gate436inter11));
  nor2  gate1819(.a(gate436inter11), .b(gate436inter6), .O(gate436inter12));
  nand2 gate1820(.a(gate436inter12), .b(gate436inter1), .O(G1245));
nand2 gate437( .a(G10), .b(G1159), .O(G1246) );
nand2 gate438( .a(G1063), .b(G1159), .O(G1247) );
nand2 gate439( .a(G11), .b(G1162), .O(G1248) );

  xor2  gate2283(.a(G1162), .b(G1066), .O(gate440inter0));
  nand2 gate2284(.a(gate440inter0), .b(s_248), .O(gate440inter1));
  and2  gate2285(.a(G1162), .b(G1066), .O(gate440inter2));
  inv1  gate2286(.a(s_248), .O(gate440inter3));
  inv1  gate2287(.a(s_249), .O(gate440inter4));
  nand2 gate2288(.a(gate440inter4), .b(gate440inter3), .O(gate440inter5));
  nor2  gate2289(.a(gate440inter5), .b(gate440inter2), .O(gate440inter6));
  inv1  gate2290(.a(G1066), .O(gate440inter7));
  inv1  gate2291(.a(G1162), .O(gate440inter8));
  nand2 gate2292(.a(gate440inter8), .b(gate440inter7), .O(gate440inter9));
  nand2 gate2293(.a(s_249), .b(gate440inter3), .O(gate440inter10));
  nor2  gate2294(.a(gate440inter10), .b(gate440inter9), .O(gate440inter11));
  nor2  gate2295(.a(gate440inter11), .b(gate440inter6), .O(gate440inter12));
  nand2 gate2296(.a(gate440inter12), .b(gate440inter1), .O(G1249));
nand2 gate441( .a(G12), .b(G1165), .O(G1250) );
nand2 gate442( .a(G1069), .b(G1165), .O(G1251) );

  xor2  gate2591(.a(G1168), .b(G13), .O(gate443inter0));
  nand2 gate2592(.a(gate443inter0), .b(s_292), .O(gate443inter1));
  and2  gate2593(.a(G1168), .b(G13), .O(gate443inter2));
  inv1  gate2594(.a(s_292), .O(gate443inter3));
  inv1  gate2595(.a(s_293), .O(gate443inter4));
  nand2 gate2596(.a(gate443inter4), .b(gate443inter3), .O(gate443inter5));
  nor2  gate2597(.a(gate443inter5), .b(gate443inter2), .O(gate443inter6));
  inv1  gate2598(.a(G13), .O(gate443inter7));
  inv1  gate2599(.a(G1168), .O(gate443inter8));
  nand2 gate2600(.a(gate443inter8), .b(gate443inter7), .O(gate443inter9));
  nand2 gate2601(.a(s_293), .b(gate443inter3), .O(gate443inter10));
  nor2  gate2602(.a(gate443inter10), .b(gate443inter9), .O(gate443inter11));
  nor2  gate2603(.a(gate443inter11), .b(gate443inter6), .O(gate443inter12));
  nand2 gate2604(.a(gate443inter12), .b(gate443inter1), .O(G1252));
nand2 gate444( .a(G1072), .b(G1168), .O(G1253) );

  xor2  gate2339(.a(G1171), .b(G14), .O(gate445inter0));
  nand2 gate2340(.a(gate445inter0), .b(s_256), .O(gate445inter1));
  and2  gate2341(.a(G1171), .b(G14), .O(gate445inter2));
  inv1  gate2342(.a(s_256), .O(gate445inter3));
  inv1  gate2343(.a(s_257), .O(gate445inter4));
  nand2 gate2344(.a(gate445inter4), .b(gate445inter3), .O(gate445inter5));
  nor2  gate2345(.a(gate445inter5), .b(gate445inter2), .O(gate445inter6));
  inv1  gate2346(.a(G14), .O(gate445inter7));
  inv1  gate2347(.a(G1171), .O(gate445inter8));
  nand2 gate2348(.a(gate445inter8), .b(gate445inter7), .O(gate445inter9));
  nand2 gate2349(.a(s_257), .b(gate445inter3), .O(gate445inter10));
  nor2  gate2350(.a(gate445inter10), .b(gate445inter9), .O(gate445inter11));
  nor2  gate2351(.a(gate445inter11), .b(gate445inter6), .O(gate445inter12));
  nand2 gate2352(.a(gate445inter12), .b(gate445inter1), .O(G1254));
nand2 gate446( .a(G1075), .b(G1171), .O(G1255) );
nand2 gate447( .a(G15), .b(G1174), .O(G1256) );
nand2 gate448( .a(G1078), .b(G1174), .O(G1257) );

  xor2  gate1583(.a(G1177), .b(G16), .O(gate449inter0));
  nand2 gate1584(.a(gate449inter0), .b(s_148), .O(gate449inter1));
  and2  gate1585(.a(G1177), .b(G16), .O(gate449inter2));
  inv1  gate1586(.a(s_148), .O(gate449inter3));
  inv1  gate1587(.a(s_149), .O(gate449inter4));
  nand2 gate1588(.a(gate449inter4), .b(gate449inter3), .O(gate449inter5));
  nor2  gate1589(.a(gate449inter5), .b(gate449inter2), .O(gate449inter6));
  inv1  gate1590(.a(G16), .O(gate449inter7));
  inv1  gate1591(.a(G1177), .O(gate449inter8));
  nand2 gate1592(.a(gate449inter8), .b(gate449inter7), .O(gate449inter9));
  nand2 gate1593(.a(s_149), .b(gate449inter3), .O(gate449inter10));
  nor2  gate1594(.a(gate449inter10), .b(gate449inter9), .O(gate449inter11));
  nor2  gate1595(.a(gate449inter11), .b(gate449inter6), .O(gate449inter12));
  nand2 gate1596(.a(gate449inter12), .b(gate449inter1), .O(G1258));
nand2 gate450( .a(G1081), .b(G1177), .O(G1259) );
nand2 gate451( .a(G17), .b(G1180), .O(G1260) );
nand2 gate452( .a(G1084), .b(G1180), .O(G1261) );

  xor2  gate2423(.a(G1183), .b(G18), .O(gate453inter0));
  nand2 gate2424(.a(gate453inter0), .b(s_268), .O(gate453inter1));
  and2  gate2425(.a(G1183), .b(G18), .O(gate453inter2));
  inv1  gate2426(.a(s_268), .O(gate453inter3));
  inv1  gate2427(.a(s_269), .O(gate453inter4));
  nand2 gate2428(.a(gate453inter4), .b(gate453inter3), .O(gate453inter5));
  nor2  gate2429(.a(gate453inter5), .b(gate453inter2), .O(gate453inter6));
  inv1  gate2430(.a(G18), .O(gate453inter7));
  inv1  gate2431(.a(G1183), .O(gate453inter8));
  nand2 gate2432(.a(gate453inter8), .b(gate453inter7), .O(gate453inter9));
  nand2 gate2433(.a(s_269), .b(gate453inter3), .O(gate453inter10));
  nor2  gate2434(.a(gate453inter10), .b(gate453inter9), .O(gate453inter11));
  nor2  gate2435(.a(gate453inter11), .b(gate453inter6), .O(gate453inter12));
  nand2 gate2436(.a(gate453inter12), .b(gate453inter1), .O(G1262));
nand2 gate454( .a(G1087), .b(G1183), .O(G1263) );

  xor2  gate2619(.a(G1186), .b(G19), .O(gate455inter0));
  nand2 gate2620(.a(gate455inter0), .b(s_296), .O(gate455inter1));
  and2  gate2621(.a(G1186), .b(G19), .O(gate455inter2));
  inv1  gate2622(.a(s_296), .O(gate455inter3));
  inv1  gate2623(.a(s_297), .O(gate455inter4));
  nand2 gate2624(.a(gate455inter4), .b(gate455inter3), .O(gate455inter5));
  nor2  gate2625(.a(gate455inter5), .b(gate455inter2), .O(gate455inter6));
  inv1  gate2626(.a(G19), .O(gate455inter7));
  inv1  gate2627(.a(G1186), .O(gate455inter8));
  nand2 gate2628(.a(gate455inter8), .b(gate455inter7), .O(gate455inter9));
  nand2 gate2629(.a(s_297), .b(gate455inter3), .O(gate455inter10));
  nor2  gate2630(.a(gate455inter10), .b(gate455inter9), .O(gate455inter11));
  nor2  gate2631(.a(gate455inter11), .b(gate455inter6), .O(gate455inter12));
  nand2 gate2632(.a(gate455inter12), .b(gate455inter1), .O(G1264));
nand2 gate456( .a(G1090), .b(G1186), .O(G1265) );
nand2 gate457( .a(G20), .b(G1189), .O(G1266) );

  xor2  gate2843(.a(G1189), .b(G1093), .O(gate458inter0));
  nand2 gate2844(.a(gate458inter0), .b(s_328), .O(gate458inter1));
  and2  gate2845(.a(G1189), .b(G1093), .O(gate458inter2));
  inv1  gate2846(.a(s_328), .O(gate458inter3));
  inv1  gate2847(.a(s_329), .O(gate458inter4));
  nand2 gate2848(.a(gate458inter4), .b(gate458inter3), .O(gate458inter5));
  nor2  gate2849(.a(gate458inter5), .b(gate458inter2), .O(gate458inter6));
  inv1  gate2850(.a(G1093), .O(gate458inter7));
  inv1  gate2851(.a(G1189), .O(gate458inter8));
  nand2 gate2852(.a(gate458inter8), .b(gate458inter7), .O(gate458inter9));
  nand2 gate2853(.a(s_329), .b(gate458inter3), .O(gate458inter10));
  nor2  gate2854(.a(gate458inter10), .b(gate458inter9), .O(gate458inter11));
  nor2  gate2855(.a(gate458inter11), .b(gate458inter6), .O(gate458inter12));
  nand2 gate2856(.a(gate458inter12), .b(gate458inter1), .O(G1267));

  xor2  gate1653(.a(G1192), .b(G21), .O(gate459inter0));
  nand2 gate1654(.a(gate459inter0), .b(s_158), .O(gate459inter1));
  and2  gate1655(.a(G1192), .b(G21), .O(gate459inter2));
  inv1  gate1656(.a(s_158), .O(gate459inter3));
  inv1  gate1657(.a(s_159), .O(gate459inter4));
  nand2 gate1658(.a(gate459inter4), .b(gate459inter3), .O(gate459inter5));
  nor2  gate1659(.a(gate459inter5), .b(gate459inter2), .O(gate459inter6));
  inv1  gate1660(.a(G21), .O(gate459inter7));
  inv1  gate1661(.a(G1192), .O(gate459inter8));
  nand2 gate1662(.a(gate459inter8), .b(gate459inter7), .O(gate459inter9));
  nand2 gate1663(.a(s_159), .b(gate459inter3), .O(gate459inter10));
  nor2  gate1664(.a(gate459inter10), .b(gate459inter9), .O(gate459inter11));
  nor2  gate1665(.a(gate459inter11), .b(gate459inter6), .O(gate459inter12));
  nand2 gate1666(.a(gate459inter12), .b(gate459inter1), .O(G1268));
nand2 gate460( .a(G1096), .b(G1192), .O(G1269) );
nand2 gate461( .a(G22), .b(G1195), .O(G1270) );

  xor2  gate1135(.a(G1195), .b(G1099), .O(gate462inter0));
  nand2 gate1136(.a(gate462inter0), .b(s_84), .O(gate462inter1));
  and2  gate1137(.a(G1195), .b(G1099), .O(gate462inter2));
  inv1  gate1138(.a(s_84), .O(gate462inter3));
  inv1  gate1139(.a(s_85), .O(gate462inter4));
  nand2 gate1140(.a(gate462inter4), .b(gate462inter3), .O(gate462inter5));
  nor2  gate1141(.a(gate462inter5), .b(gate462inter2), .O(gate462inter6));
  inv1  gate1142(.a(G1099), .O(gate462inter7));
  inv1  gate1143(.a(G1195), .O(gate462inter8));
  nand2 gate1144(.a(gate462inter8), .b(gate462inter7), .O(gate462inter9));
  nand2 gate1145(.a(s_85), .b(gate462inter3), .O(gate462inter10));
  nor2  gate1146(.a(gate462inter10), .b(gate462inter9), .O(gate462inter11));
  nor2  gate1147(.a(gate462inter11), .b(gate462inter6), .O(gate462inter12));
  nand2 gate1148(.a(gate462inter12), .b(gate462inter1), .O(G1271));

  xor2  gate1121(.a(G1198), .b(G23), .O(gate463inter0));
  nand2 gate1122(.a(gate463inter0), .b(s_82), .O(gate463inter1));
  and2  gate1123(.a(G1198), .b(G23), .O(gate463inter2));
  inv1  gate1124(.a(s_82), .O(gate463inter3));
  inv1  gate1125(.a(s_83), .O(gate463inter4));
  nand2 gate1126(.a(gate463inter4), .b(gate463inter3), .O(gate463inter5));
  nor2  gate1127(.a(gate463inter5), .b(gate463inter2), .O(gate463inter6));
  inv1  gate1128(.a(G23), .O(gate463inter7));
  inv1  gate1129(.a(G1198), .O(gate463inter8));
  nand2 gate1130(.a(gate463inter8), .b(gate463inter7), .O(gate463inter9));
  nand2 gate1131(.a(s_83), .b(gate463inter3), .O(gate463inter10));
  nor2  gate1132(.a(gate463inter10), .b(gate463inter9), .O(gate463inter11));
  nor2  gate1133(.a(gate463inter11), .b(gate463inter6), .O(gate463inter12));
  nand2 gate1134(.a(gate463inter12), .b(gate463inter1), .O(G1272));
nand2 gate464( .a(G1102), .b(G1198), .O(G1273) );

  xor2  gate2731(.a(G1201), .b(G24), .O(gate465inter0));
  nand2 gate2732(.a(gate465inter0), .b(s_312), .O(gate465inter1));
  and2  gate2733(.a(G1201), .b(G24), .O(gate465inter2));
  inv1  gate2734(.a(s_312), .O(gate465inter3));
  inv1  gate2735(.a(s_313), .O(gate465inter4));
  nand2 gate2736(.a(gate465inter4), .b(gate465inter3), .O(gate465inter5));
  nor2  gate2737(.a(gate465inter5), .b(gate465inter2), .O(gate465inter6));
  inv1  gate2738(.a(G24), .O(gate465inter7));
  inv1  gate2739(.a(G1201), .O(gate465inter8));
  nand2 gate2740(.a(gate465inter8), .b(gate465inter7), .O(gate465inter9));
  nand2 gate2741(.a(s_313), .b(gate465inter3), .O(gate465inter10));
  nor2  gate2742(.a(gate465inter10), .b(gate465inter9), .O(gate465inter11));
  nor2  gate2743(.a(gate465inter11), .b(gate465inter6), .O(gate465inter12));
  nand2 gate2744(.a(gate465inter12), .b(gate465inter1), .O(G1274));

  xor2  gate939(.a(G1201), .b(G1105), .O(gate466inter0));
  nand2 gate940(.a(gate466inter0), .b(s_56), .O(gate466inter1));
  and2  gate941(.a(G1201), .b(G1105), .O(gate466inter2));
  inv1  gate942(.a(s_56), .O(gate466inter3));
  inv1  gate943(.a(s_57), .O(gate466inter4));
  nand2 gate944(.a(gate466inter4), .b(gate466inter3), .O(gate466inter5));
  nor2  gate945(.a(gate466inter5), .b(gate466inter2), .O(gate466inter6));
  inv1  gate946(.a(G1105), .O(gate466inter7));
  inv1  gate947(.a(G1201), .O(gate466inter8));
  nand2 gate948(.a(gate466inter8), .b(gate466inter7), .O(gate466inter9));
  nand2 gate949(.a(s_57), .b(gate466inter3), .O(gate466inter10));
  nor2  gate950(.a(gate466inter10), .b(gate466inter9), .O(gate466inter11));
  nor2  gate951(.a(gate466inter11), .b(gate466inter6), .O(gate466inter12));
  nand2 gate952(.a(gate466inter12), .b(gate466inter1), .O(G1275));
nand2 gate467( .a(G25), .b(G1204), .O(G1276) );
nand2 gate468( .a(G1108), .b(G1204), .O(G1277) );

  xor2  gate2087(.a(G1207), .b(G26), .O(gate469inter0));
  nand2 gate2088(.a(gate469inter0), .b(s_220), .O(gate469inter1));
  and2  gate2089(.a(G1207), .b(G26), .O(gate469inter2));
  inv1  gate2090(.a(s_220), .O(gate469inter3));
  inv1  gate2091(.a(s_221), .O(gate469inter4));
  nand2 gate2092(.a(gate469inter4), .b(gate469inter3), .O(gate469inter5));
  nor2  gate2093(.a(gate469inter5), .b(gate469inter2), .O(gate469inter6));
  inv1  gate2094(.a(G26), .O(gate469inter7));
  inv1  gate2095(.a(G1207), .O(gate469inter8));
  nand2 gate2096(.a(gate469inter8), .b(gate469inter7), .O(gate469inter9));
  nand2 gate2097(.a(s_221), .b(gate469inter3), .O(gate469inter10));
  nor2  gate2098(.a(gate469inter10), .b(gate469inter9), .O(gate469inter11));
  nor2  gate2099(.a(gate469inter11), .b(gate469inter6), .O(gate469inter12));
  nand2 gate2100(.a(gate469inter12), .b(gate469inter1), .O(G1278));
nand2 gate470( .a(G1111), .b(G1207), .O(G1279) );

  xor2  gate2199(.a(G1210), .b(G27), .O(gate471inter0));
  nand2 gate2200(.a(gate471inter0), .b(s_236), .O(gate471inter1));
  and2  gate2201(.a(G1210), .b(G27), .O(gate471inter2));
  inv1  gate2202(.a(s_236), .O(gate471inter3));
  inv1  gate2203(.a(s_237), .O(gate471inter4));
  nand2 gate2204(.a(gate471inter4), .b(gate471inter3), .O(gate471inter5));
  nor2  gate2205(.a(gate471inter5), .b(gate471inter2), .O(gate471inter6));
  inv1  gate2206(.a(G27), .O(gate471inter7));
  inv1  gate2207(.a(G1210), .O(gate471inter8));
  nand2 gate2208(.a(gate471inter8), .b(gate471inter7), .O(gate471inter9));
  nand2 gate2209(.a(s_237), .b(gate471inter3), .O(gate471inter10));
  nor2  gate2210(.a(gate471inter10), .b(gate471inter9), .O(gate471inter11));
  nor2  gate2211(.a(gate471inter11), .b(gate471inter6), .O(gate471inter12));
  nand2 gate2212(.a(gate471inter12), .b(gate471inter1), .O(G1280));

  xor2  gate1233(.a(G1210), .b(G1114), .O(gate472inter0));
  nand2 gate1234(.a(gate472inter0), .b(s_98), .O(gate472inter1));
  and2  gate1235(.a(G1210), .b(G1114), .O(gate472inter2));
  inv1  gate1236(.a(s_98), .O(gate472inter3));
  inv1  gate1237(.a(s_99), .O(gate472inter4));
  nand2 gate1238(.a(gate472inter4), .b(gate472inter3), .O(gate472inter5));
  nor2  gate1239(.a(gate472inter5), .b(gate472inter2), .O(gate472inter6));
  inv1  gate1240(.a(G1114), .O(gate472inter7));
  inv1  gate1241(.a(G1210), .O(gate472inter8));
  nand2 gate1242(.a(gate472inter8), .b(gate472inter7), .O(gate472inter9));
  nand2 gate1243(.a(s_99), .b(gate472inter3), .O(gate472inter10));
  nor2  gate1244(.a(gate472inter10), .b(gate472inter9), .O(gate472inter11));
  nor2  gate1245(.a(gate472inter11), .b(gate472inter6), .O(gate472inter12));
  nand2 gate1246(.a(gate472inter12), .b(gate472inter1), .O(G1281));
nand2 gate473( .a(G28), .b(G1213), .O(G1282) );

  xor2  gate645(.a(G1213), .b(G1117), .O(gate474inter0));
  nand2 gate646(.a(gate474inter0), .b(s_14), .O(gate474inter1));
  and2  gate647(.a(G1213), .b(G1117), .O(gate474inter2));
  inv1  gate648(.a(s_14), .O(gate474inter3));
  inv1  gate649(.a(s_15), .O(gate474inter4));
  nand2 gate650(.a(gate474inter4), .b(gate474inter3), .O(gate474inter5));
  nor2  gate651(.a(gate474inter5), .b(gate474inter2), .O(gate474inter6));
  inv1  gate652(.a(G1117), .O(gate474inter7));
  inv1  gate653(.a(G1213), .O(gate474inter8));
  nand2 gate654(.a(gate474inter8), .b(gate474inter7), .O(gate474inter9));
  nand2 gate655(.a(s_15), .b(gate474inter3), .O(gate474inter10));
  nor2  gate656(.a(gate474inter10), .b(gate474inter9), .O(gate474inter11));
  nor2  gate657(.a(gate474inter11), .b(gate474inter6), .O(gate474inter12));
  nand2 gate658(.a(gate474inter12), .b(gate474inter1), .O(G1283));
nand2 gate475( .a(G29), .b(G1216), .O(G1284) );

  xor2  gate2507(.a(G1216), .b(G1120), .O(gate476inter0));
  nand2 gate2508(.a(gate476inter0), .b(s_280), .O(gate476inter1));
  and2  gate2509(.a(G1216), .b(G1120), .O(gate476inter2));
  inv1  gate2510(.a(s_280), .O(gate476inter3));
  inv1  gate2511(.a(s_281), .O(gate476inter4));
  nand2 gate2512(.a(gate476inter4), .b(gate476inter3), .O(gate476inter5));
  nor2  gate2513(.a(gate476inter5), .b(gate476inter2), .O(gate476inter6));
  inv1  gate2514(.a(G1120), .O(gate476inter7));
  inv1  gate2515(.a(G1216), .O(gate476inter8));
  nand2 gate2516(.a(gate476inter8), .b(gate476inter7), .O(gate476inter9));
  nand2 gate2517(.a(s_281), .b(gate476inter3), .O(gate476inter10));
  nor2  gate2518(.a(gate476inter10), .b(gate476inter9), .O(gate476inter11));
  nor2  gate2519(.a(gate476inter11), .b(gate476inter6), .O(gate476inter12));
  nand2 gate2520(.a(gate476inter12), .b(gate476inter1), .O(G1285));

  xor2  gate1331(.a(G1219), .b(G30), .O(gate477inter0));
  nand2 gate1332(.a(gate477inter0), .b(s_112), .O(gate477inter1));
  and2  gate1333(.a(G1219), .b(G30), .O(gate477inter2));
  inv1  gate1334(.a(s_112), .O(gate477inter3));
  inv1  gate1335(.a(s_113), .O(gate477inter4));
  nand2 gate1336(.a(gate477inter4), .b(gate477inter3), .O(gate477inter5));
  nor2  gate1337(.a(gate477inter5), .b(gate477inter2), .O(gate477inter6));
  inv1  gate1338(.a(G30), .O(gate477inter7));
  inv1  gate1339(.a(G1219), .O(gate477inter8));
  nand2 gate1340(.a(gate477inter8), .b(gate477inter7), .O(gate477inter9));
  nand2 gate1341(.a(s_113), .b(gate477inter3), .O(gate477inter10));
  nor2  gate1342(.a(gate477inter10), .b(gate477inter9), .O(gate477inter11));
  nor2  gate1343(.a(gate477inter11), .b(gate477inter6), .O(gate477inter12));
  nand2 gate1344(.a(gate477inter12), .b(gate477inter1), .O(G1286));
nand2 gate478( .a(G1123), .b(G1219), .O(G1287) );
nand2 gate479( .a(G31), .b(G1222), .O(G1288) );
nand2 gate480( .a(G1126), .b(G1222), .O(G1289) );
nand2 gate481( .a(G32), .b(G1225), .O(G1290) );

  xor2  gate1891(.a(G1225), .b(G1129), .O(gate482inter0));
  nand2 gate1892(.a(gate482inter0), .b(s_192), .O(gate482inter1));
  and2  gate1893(.a(G1225), .b(G1129), .O(gate482inter2));
  inv1  gate1894(.a(s_192), .O(gate482inter3));
  inv1  gate1895(.a(s_193), .O(gate482inter4));
  nand2 gate1896(.a(gate482inter4), .b(gate482inter3), .O(gate482inter5));
  nor2  gate1897(.a(gate482inter5), .b(gate482inter2), .O(gate482inter6));
  inv1  gate1898(.a(G1129), .O(gate482inter7));
  inv1  gate1899(.a(G1225), .O(gate482inter8));
  nand2 gate1900(.a(gate482inter8), .b(gate482inter7), .O(gate482inter9));
  nand2 gate1901(.a(s_193), .b(gate482inter3), .O(gate482inter10));
  nor2  gate1902(.a(gate482inter10), .b(gate482inter9), .O(gate482inter11));
  nor2  gate1903(.a(gate482inter11), .b(gate482inter6), .O(gate482inter12));
  nand2 gate1904(.a(gate482inter12), .b(gate482inter1), .O(G1291));
nand2 gate483( .a(G1228), .b(G1229), .O(G1292) );
nand2 gate484( .a(G1230), .b(G1231), .O(G1293) );

  xor2  gate1975(.a(G1233), .b(G1232), .O(gate485inter0));
  nand2 gate1976(.a(gate485inter0), .b(s_204), .O(gate485inter1));
  and2  gate1977(.a(G1233), .b(G1232), .O(gate485inter2));
  inv1  gate1978(.a(s_204), .O(gate485inter3));
  inv1  gate1979(.a(s_205), .O(gate485inter4));
  nand2 gate1980(.a(gate485inter4), .b(gate485inter3), .O(gate485inter5));
  nor2  gate1981(.a(gate485inter5), .b(gate485inter2), .O(gate485inter6));
  inv1  gate1982(.a(G1232), .O(gate485inter7));
  inv1  gate1983(.a(G1233), .O(gate485inter8));
  nand2 gate1984(.a(gate485inter8), .b(gate485inter7), .O(gate485inter9));
  nand2 gate1985(.a(s_205), .b(gate485inter3), .O(gate485inter10));
  nor2  gate1986(.a(gate485inter10), .b(gate485inter9), .O(gate485inter11));
  nor2  gate1987(.a(gate485inter11), .b(gate485inter6), .O(gate485inter12));
  nand2 gate1988(.a(gate485inter12), .b(gate485inter1), .O(G1294));
nand2 gate486( .a(G1234), .b(G1235), .O(G1295) );

  xor2  gate1457(.a(G1237), .b(G1236), .O(gate487inter0));
  nand2 gate1458(.a(gate487inter0), .b(s_130), .O(gate487inter1));
  and2  gate1459(.a(G1237), .b(G1236), .O(gate487inter2));
  inv1  gate1460(.a(s_130), .O(gate487inter3));
  inv1  gate1461(.a(s_131), .O(gate487inter4));
  nand2 gate1462(.a(gate487inter4), .b(gate487inter3), .O(gate487inter5));
  nor2  gate1463(.a(gate487inter5), .b(gate487inter2), .O(gate487inter6));
  inv1  gate1464(.a(G1236), .O(gate487inter7));
  inv1  gate1465(.a(G1237), .O(gate487inter8));
  nand2 gate1466(.a(gate487inter8), .b(gate487inter7), .O(gate487inter9));
  nand2 gate1467(.a(s_131), .b(gate487inter3), .O(gate487inter10));
  nor2  gate1468(.a(gate487inter10), .b(gate487inter9), .O(gate487inter11));
  nor2  gate1469(.a(gate487inter11), .b(gate487inter6), .O(gate487inter12));
  nand2 gate1470(.a(gate487inter12), .b(gate487inter1), .O(G1296));

  xor2  gate2493(.a(G1239), .b(G1238), .O(gate488inter0));
  nand2 gate2494(.a(gate488inter0), .b(s_278), .O(gate488inter1));
  and2  gate2495(.a(G1239), .b(G1238), .O(gate488inter2));
  inv1  gate2496(.a(s_278), .O(gate488inter3));
  inv1  gate2497(.a(s_279), .O(gate488inter4));
  nand2 gate2498(.a(gate488inter4), .b(gate488inter3), .O(gate488inter5));
  nor2  gate2499(.a(gate488inter5), .b(gate488inter2), .O(gate488inter6));
  inv1  gate2500(.a(G1238), .O(gate488inter7));
  inv1  gate2501(.a(G1239), .O(gate488inter8));
  nand2 gate2502(.a(gate488inter8), .b(gate488inter7), .O(gate488inter9));
  nand2 gate2503(.a(s_279), .b(gate488inter3), .O(gate488inter10));
  nor2  gate2504(.a(gate488inter10), .b(gate488inter9), .O(gate488inter11));
  nor2  gate2505(.a(gate488inter11), .b(gate488inter6), .O(gate488inter12));
  nand2 gate2506(.a(gate488inter12), .b(gate488inter1), .O(G1297));

  xor2  gate3151(.a(G1241), .b(G1240), .O(gate489inter0));
  nand2 gate3152(.a(gate489inter0), .b(s_372), .O(gate489inter1));
  and2  gate3153(.a(G1241), .b(G1240), .O(gate489inter2));
  inv1  gate3154(.a(s_372), .O(gate489inter3));
  inv1  gate3155(.a(s_373), .O(gate489inter4));
  nand2 gate3156(.a(gate489inter4), .b(gate489inter3), .O(gate489inter5));
  nor2  gate3157(.a(gate489inter5), .b(gate489inter2), .O(gate489inter6));
  inv1  gate3158(.a(G1240), .O(gate489inter7));
  inv1  gate3159(.a(G1241), .O(gate489inter8));
  nand2 gate3160(.a(gate489inter8), .b(gate489inter7), .O(gate489inter9));
  nand2 gate3161(.a(s_373), .b(gate489inter3), .O(gate489inter10));
  nor2  gate3162(.a(gate489inter10), .b(gate489inter9), .O(gate489inter11));
  nor2  gate3163(.a(gate489inter11), .b(gate489inter6), .O(gate489inter12));
  nand2 gate3164(.a(gate489inter12), .b(gate489inter1), .O(G1298));

  xor2  gate883(.a(G1243), .b(G1242), .O(gate490inter0));
  nand2 gate884(.a(gate490inter0), .b(s_48), .O(gate490inter1));
  and2  gate885(.a(G1243), .b(G1242), .O(gate490inter2));
  inv1  gate886(.a(s_48), .O(gate490inter3));
  inv1  gate887(.a(s_49), .O(gate490inter4));
  nand2 gate888(.a(gate490inter4), .b(gate490inter3), .O(gate490inter5));
  nor2  gate889(.a(gate490inter5), .b(gate490inter2), .O(gate490inter6));
  inv1  gate890(.a(G1242), .O(gate490inter7));
  inv1  gate891(.a(G1243), .O(gate490inter8));
  nand2 gate892(.a(gate490inter8), .b(gate490inter7), .O(gate490inter9));
  nand2 gate893(.a(s_49), .b(gate490inter3), .O(gate490inter10));
  nor2  gate894(.a(gate490inter10), .b(gate490inter9), .O(gate490inter11));
  nor2  gate895(.a(gate490inter11), .b(gate490inter6), .O(gate490inter12));
  nand2 gate896(.a(gate490inter12), .b(gate490inter1), .O(G1299));

  xor2  gate3193(.a(G1245), .b(G1244), .O(gate491inter0));
  nand2 gate3194(.a(gate491inter0), .b(s_378), .O(gate491inter1));
  and2  gate3195(.a(G1245), .b(G1244), .O(gate491inter2));
  inv1  gate3196(.a(s_378), .O(gate491inter3));
  inv1  gate3197(.a(s_379), .O(gate491inter4));
  nand2 gate3198(.a(gate491inter4), .b(gate491inter3), .O(gate491inter5));
  nor2  gate3199(.a(gate491inter5), .b(gate491inter2), .O(gate491inter6));
  inv1  gate3200(.a(G1244), .O(gate491inter7));
  inv1  gate3201(.a(G1245), .O(gate491inter8));
  nand2 gate3202(.a(gate491inter8), .b(gate491inter7), .O(gate491inter9));
  nand2 gate3203(.a(s_379), .b(gate491inter3), .O(gate491inter10));
  nor2  gate3204(.a(gate491inter10), .b(gate491inter9), .O(gate491inter11));
  nor2  gate3205(.a(gate491inter11), .b(gate491inter6), .O(gate491inter12));
  nand2 gate3206(.a(gate491inter12), .b(gate491inter1), .O(G1300));
nand2 gate492( .a(G1246), .b(G1247), .O(G1301) );

  xor2  gate2325(.a(G1249), .b(G1248), .O(gate493inter0));
  nand2 gate2326(.a(gate493inter0), .b(s_254), .O(gate493inter1));
  and2  gate2327(.a(G1249), .b(G1248), .O(gate493inter2));
  inv1  gate2328(.a(s_254), .O(gate493inter3));
  inv1  gate2329(.a(s_255), .O(gate493inter4));
  nand2 gate2330(.a(gate493inter4), .b(gate493inter3), .O(gate493inter5));
  nor2  gate2331(.a(gate493inter5), .b(gate493inter2), .O(gate493inter6));
  inv1  gate2332(.a(G1248), .O(gate493inter7));
  inv1  gate2333(.a(G1249), .O(gate493inter8));
  nand2 gate2334(.a(gate493inter8), .b(gate493inter7), .O(gate493inter9));
  nand2 gate2335(.a(s_255), .b(gate493inter3), .O(gate493inter10));
  nor2  gate2336(.a(gate493inter10), .b(gate493inter9), .O(gate493inter11));
  nor2  gate2337(.a(gate493inter11), .b(gate493inter6), .O(gate493inter12));
  nand2 gate2338(.a(gate493inter12), .b(gate493inter1), .O(G1302));

  xor2  gate2353(.a(G1251), .b(G1250), .O(gate494inter0));
  nand2 gate2354(.a(gate494inter0), .b(s_258), .O(gate494inter1));
  and2  gate2355(.a(G1251), .b(G1250), .O(gate494inter2));
  inv1  gate2356(.a(s_258), .O(gate494inter3));
  inv1  gate2357(.a(s_259), .O(gate494inter4));
  nand2 gate2358(.a(gate494inter4), .b(gate494inter3), .O(gate494inter5));
  nor2  gate2359(.a(gate494inter5), .b(gate494inter2), .O(gate494inter6));
  inv1  gate2360(.a(G1250), .O(gate494inter7));
  inv1  gate2361(.a(G1251), .O(gate494inter8));
  nand2 gate2362(.a(gate494inter8), .b(gate494inter7), .O(gate494inter9));
  nand2 gate2363(.a(s_259), .b(gate494inter3), .O(gate494inter10));
  nor2  gate2364(.a(gate494inter10), .b(gate494inter9), .O(gate494inter11));
  nor2  gate2365(.a(gate494inter11), .b(gate494inter6), .O(gate494inter12));
  nand2 gate2366(.a(gate494inter12), .b(gate494inter1), .O(G1303));
nand2 gate495( .a(G1252), .b(G1253), .O(G1304) );

  xor2  gate561(.a(G1255), .b(G1254), .O(gate496inter0));
  nand2 gate562(.a(gate496inter0), .b(s_2), .O(gate496inter1));
  and2  gate563(.a(G1255), .b(G1254), .O(gate496inter2));
  inv1  gate564(.a(s_2), .O(gate496inter3));
  inv1  gate565(.a(s_3), .O(gate496inter4));
  nand2 gate566(.a(gate496inter4), .b(gate496inter3), .O(gate496inter5));
  nor2  gate567(.a(gate496inter5), .b(gate496inter2), .O(gate496inter6));
  inv1  gate568(.a(G1254), .O(gate496inter7));
  inv1  gate569(.a(G1255), .O(gate496inter8));
  nand2 gate570(.a(gate496inter8), .b(gate496inter7), .O(gate496inter9));
  nand2 gate571(.a(s_3), .b(gate496inter3), .O(gate496inter10));
  nor2  gate572(.a(gate496inter10), .b(gate496inter9), .O(gate496inter11));
  nor2  gate573(.a(gate496inter11), .b(gate496inter6), .O(gate496inter12));
  nand2 gate574(.a(gate496inter12), .b(gate496inter1), .O(G1305));
nand2 gate497( .a(G1256), .b(G1257), .O(G1306) );

  xor2  gate2535(.a(G1259), .b(G1258), .O(gate498inter0));
  nand2 gate2536(.a(gate498inter0), .b(s_284), .O(gate498inter1));
  and2  gate2537(.a(G1259), .b(G1258), .O(gate498inter2));
  inv1  gate2538(.a(s_284), .O(gate498inter3));
  inv1  gate2539(.a(s_285), .O(gate498inter4));
  nand2 gate2540(.a(gate498inter4), .b(gate498inter3), .O(gate498inter5));
  nor2  gate2541(.a(gate498inter5), .b(gate498inter2), .O(gate498inter6));
  inv1  gate2542(.a(G1258), .O(gate498inter7));
  inv1  gate2543(.a(G1259), .O(gate498inter8));
  nand2 gate2544(.a(gate498inter8), .b(gate498inter7), .O(gate498inter9));
  nand2 gate2545(.a(s_285), .b(gate498inter3), .O(gate498inter10));
  nor2  gate2546(.a(gate498inter10), .b(gate498inter9), .O(gate498inter11));
  nor2  gate2547(.a(gate498inter11), .b(gate498inter6), .O(gate498inter12));
  nand2 gate2548(.a(gate498inter12), .b(gate498inter1), .O(G1307));

  xor2  gate673(.a(G1261), .b(G1260), .O(gate499inter0));
  nand2 gate674(.a(gate499inter0), .b(s_18), .O(gate499inter1));
  and2  gate675(.a(G1261), .b(G1260), .O(gate499inter2));
  inv1  gate676(.a(s_18), .O(gate499inter3));
  inv1  gate677(.a(s_19), .O(gate499inter4));
  nand2 gate678(.a(gate499inter4), .b(gate499inter3), .O(gate499inter5));
  nor2  gate679(.a(gate499inter5), .b(gate499inter2), .O(gate499inter6));
  inv1  gate680(.a(G1260), .O(gate499inter7));
  inv1  gate681(.a(G1261), .O(gate499inter8));
  nand2 gate682(.a(gate499inter8), .b(gate499inter7), .O(gate499inter9));
  nand2 gate683(.a(s_19), .b(gate499inter3), .O(gate499inter10));
  nor2  gate684(.a(gate499inter10), .b(gate499inter9), .O(gate499inter11));
  nor2  gate685(.a(gate499inter11), .b(gate499inter6), .O(gate499inter12));
  nand2 gate686(.a(gate499inter12), .b(gate499inter1), .O(G1308));

  xor2  gate2479(.a(G1263), .b(G1262), .O(gate500inter0));
  nand2 gate2480(.a(gate500inter0), .b(s_276), .O(gate500inter1));
  and2  gate2481(.a(G1263), .b(G1262), .O(gate500inter2));
  inv1  gate2482(.a(s_276), .O(gate500inter3));
  inv1  gate2483(.a(s_277), .O(gate500inter4));
  nand2 gate2484(.a(gate500inter4), .b(gate500inter3), .O(gate500inter5));
  nor2  gate2485(.a(gate500inter5), .b(gate500inter2), .O(gate500inter6));
  inv1  gate2486(.a(G1262), .O(gate500inter7));
  inv1  gate2487(.a(G1263), .O(gate500inter8));
  nand2 gate2488(.a(gate500inter8), .b(gate500inter7), .O(gate500inter9));
  nand2 gate2489(.a(s_277), .b(gate500inter3), .O(gate500inter10));
  nor2  gate2490(.a(gate500inter10), .b(gate500inter9), .O(gate500inter11));
  nor2  gate2491(.a(gate500inter11), .b(gate500inter6), .O(gate500inter12));
  nand2 gate2492(.a(gate500inter12), .b(gate500inter1), .O(G1309));

  xor2  gate1541(.a(G1265), .b(G1264), .O(gate501inter0));
  nand2 gate1542(.a(gate501inter0), .b(s_142), .O(gate501inter1));
  and2  gate1543(.a(G1265), .b(G1264), .O(gate501inter2));
  inv1  gate1544(.a(s_142), .O(gate501inter3));
  inv1  gate1545(.a(s_143), .O(gate501inter4));
  nand2 gate1546(.a(gate501inter4), .b(gate501inter3), .O(gate501inter5));
  nor2  gate1547(.a(gate501inter5), .b(gate501inter2), .O(gate501inter6));
  inv1  gate1548(.a(G1264), .O(gate501inter7));
  inv1  gate1549(.a(G1265), .O(gate501inter8));
  nand2 gate1550(.a(gate501inter8), .b(gate501inter7), .O(gate501inter9));
  nand2 gate1551(.a(s_143), .b(gate501inter3), .O(gate501inter10));
  nor2  gate1552(.a(gate501inter10), .b(gate501inter9), .O(gate501inter11));
  nor2  gate1553(.a(gate501inter11), .b(gate501inter6), .O(gate501inter12));
  nand2 gate1554(.a(gate501inter12), .b(gate501inter1), .O(G1310));
nand2 gate502( .a(G1266), .b(G1267), .O(G1311) );
nand2 gate503( .a(G1268), .b(G1269), .O(G1312) );
nand2 gate504( .a(G1270), .b(G1271), .O(G1313) );

  xor2  gate1289(.a(G1273), .b(G1272), .O(gate505inter0));
  nand2 gate1290(.a(gate505inter0), .b(s_106), .O(gate505inter1));
  and2  gate1291(.a(G1273), .b(G1272), .O(gate505inter2));
  inv1  gate1292(.a(s_106), .O(gate505inter3));
  inv1  gate1293(.a(s_107), .O(gate505inter4));
  nand2 gate1294(.a(gate505inter4), .b(gate505inter3), .O(gate505inter5));
  nor2  gate1295(.a(gate505inter5), .b(gate505inter2), .O(gate505inter6));
  inv1  gate1296(.a(G1272), .O(gate505inter7));
  inv1  gate1297(.a(G1273), .O(gate505inter8));
  nand2 gate1298(.a(gate505inter8), .b(gate505inter7), .O(gate505inter9));
  nand2 gate1299(.a(s_107), .b(gate505inter3), .O(gate505inter10));
  nor2  gate1300(.a(gate505inter10), .b(gate505inter9), .O(gate505inter11));
  nor2  gate1301(.a(gate505inter11), .b(gate505inter6), .O(gate505inter12));
  nand2 gate1302(.a(gate505inter12), .b(gate505inter1), .O(G1314));
nand2 gate506( .a(G1274), .b(G1275), .O(G1315) );
nand2 gate507( .a(G1276), .b(G1277), .O(G1316) );

  xor2  gate813(.a(G1279), .b(G1278), .O(gate508inter0));
  nand2 gate814(.a(gate508inter0), .b(s_38), .O(gate508inter1));
  and2  gate815(.a(G1279), .b(G1278), .O(gate508inter2));
  inv1  gate816(.a(s_38), .O(gate508inter3));
  inv1  gate817(.a(s_39), .O(gate508inter4));
  nand2 gate818(.a(gate508inter4), .b(gate508inter3), .O(gate508inter5));
  nor2  gate819(.a(gate508inter5), .b(gate508inter2), .O(gate508inter6));
  inv1  gate820(.a(G1278), .O(gate508inter7));
  inv1  gate821(.a(G1279), .O(gate508inter8));
  nand2 gate822(.a(gate508inter8), .b(gate508inter7), .O(gate508inter9));
  nand2 gate823(.a(s_39), .b(gate508inter3), .O(gate508inter10));
  nor2  gate824(.a(gate508inter10), .b(gate508inter9), .O(gate508inter11));
  nor2  gate825(.a(gate508inter11), .b(gate508inter6), .O(gate508inter12));
  nand2 gate826(.a(gate508inter12), .b(gate508inter1), .O(G1317));

  xor2  gate1247(.a(G1281), .b(G1280), .O(gate509inter0));
  nand2 gate1248(.a(gate509inter0), .b(s_100), .O(gate509inter1));
  and2  gate1249(.a(G1281), .b(G1280), .O(gate509inter2));
  inv1  gate1250(.a(s_100), .O(gate509inter3));
  inv1  gate1251(.a(s_101), .O(gate509inter4));
  nand2 gate1252(.a(gate509inter4), .b(gate509inter3), .O(gate509inter5));
  nor2  gate1253(.a(gate509inter5), .b(gate509inter2), .O(gate509inter6));
  inv1  gate1254(.a(G1280), .O(gate509inter7));
  inv1  gate1255(.a(G1281), .O(gate509inter8));
  nand2 gate1256(.a(gate509inter8), .b(gate509inter7), .O(gate509inter9));
  nand2 gate1257(.a(s_101), .b(gate509inter3), .O(gate509inter10));
  nor2  gate1258(.a(gate509inter10), .b(gate509inter9), .O(gate509inter11));
  nor2  gate1259(.a(gate509inter11), .b(gate509inter6), .O(gate509inter12));
  nand2 gate1260(.a(gate509inter12), .b(gate509inter1), .O(G1318));

  xor2  gate1905(.a(G1283), .b(G1282), .O(gate510inter0));
  nand2 gate1906(.a(gate510inter0), .b(s_194), .O(gate510inter1));
  and2  gate1907(.a(G1283), .b(G1282), .O(gate510inter2));
  inv1  gate1908(.a(s_194), .O(gate510inter3));
  inv1  gate1909(.a(s_195), .O(gate510inter4));
  nand2 gate1910(.a(gate510inter4), .b(gate510inter3), .O(gate510inter5));
  nor2  gate1911(.a(gate510inter5), .b(gate510inter2), .O(gate510inter6));
  inv1  gate1912(.a(G1282), .O(gate510inter7));
  inv1  gate1913(.a(G1283), .O(gate510inter8));
  nand2 gate1914(.a(gate510inter8), .b(gate510inter7), .O(gate510inter9));
  nand2 gate1915(.a(s_195), .b(gate510inter3), .O(gate510inter10));
  nor2  gate1916(.a(gate510inter10), .b(gate510inter9), .O(gate510inter11));
  nor2  gate1917(.a(gate510inter11), .b(gate510inter6), .O(gate510inter12));
  nand2 gate1918(.a(gate510inter12), .b(gate510inter1), .O(G1319));
nand2 gate511( .a(G1284), .b(G1285), .O(G1320) );

  xor2  gate771(.a(G1287), .b(G1286), .O(gate512inter0));
  nand2 gate772(.a(gate512inter0), .b(s_32), .O(gate512inter1));
  and2  gate773(.a(G1287), .b(G1286), .O(gate512inter2));
  inv1  gate774(.a(s_32), .O(gate512inter3));
  inv1  gate775(.a(s_33), .O(gate512inter4));
  nand2 gate776(.a(gate512inter4), .b(gate512inter3), .O(gate512inter5));
  nor2  gate777(.a(gate512inter5), .b(gate512inter2), .O(gate512inter6));
  inv1  gate778(.a(G1286), .O(gate512inter7));
  inv1  gate779(.a(G1287), .O(gate512inter8));
  nand2 gate780(.a(gate512inter8), .b(gate512inter7), .O(gate512inter9));
  nand2 gate781(.a(s_33), .b(gate512inter3), .O(gate512inter10));
  nor2  gate782(.a(gate512inter10), .b(gate512inter9), .O(gate512inter11));
  nor2  gate783(.a(gate512inter11), .b(gate512inter6), .O(gate512inter12));
  nand2 gate784(.a(gate512inter12), .b(gate512inter1), .O(G1321));

  xor2  gate1345(.a(G1289), .b(G1288), .O(gate513inter0));
  nand2 gate1346(.a(gate513inter0), .b(s_114), .O(gate513inter1));
  and2  gate1347(.a(G1289), .b(G1288), .O(gate513inter2));
  inv1  gate1348(.a(s_114), .O(gate513inter3));
  inv1  gate1349(.a(s_115), .O(gate513inter4));
  nand2 gate1350(.a(gate513inter4), .b(gate513inter3), .O(gate513inter5));
  nor2  gate1351(.a(gate513inter5), .b(gate513inter2), .O(gate513inter6));
  inv1  gate1352(.a(G1288), .O(gate513inter7));
  inv1  gate1353(.a(G1289), .O(gate513inter8));
  nand2 gate1354(.a(gate513inter8), .b(gate513inter7), .O(gate513inter9));
  nand2 gate1355(.a(s_115), .b(gate513inter3), .O(gate513inter10));
  nor2  gate1356(.a(gate513inter10), .b(gate513inter9), .O(gate513inter11));
  nor2  gate1357(.a(gate513inter11), .b(gate513inter6), .O(gate513inter12));
  nand2 gate1358(.a(gate513inter12), .b(gate513inter1), .O(G1322));

  xor2  gate2073(.a(G1291), .b(G1290), .O(gate514inter0));
  nand2 gate2074(.a(gate514inter0), .b(s_218), .O(gate514inter1));
  and2  gate2075(.a(G1291), .b(G1290), .O(gate514inter2));
  inv1  gate2076(.a(s_218), .O(gate514inter3));
  inv1  gate2077(.a(s_219), .O(gate514inter4));
  nand2 gate2078(.a(gate514inter4), .b(gate514inter3), .O(gate514inter5));
  nor2  gate2079(.a(gate514inter5), .b(gate514inter2), .O(gate514inter6));
  inv1  gate2080(.a(G1290), .O(gate514inter7));
  inv1  gate2081(.a(G1291), .O(gate514inter8));
  nand2 gate2082(.a(gate514inter8), .b(gate514inter7), .O(gate514inter9));
  nand2 gate2083(.a(s_219), .b(gate514inter3), .O(gate514inter10));
  nor2  gate2084(.a(gate514inter10), .b(gate514inter9), .O(gate514inter11));
  nor2  gate2085(.a(gate514inter11), .b(gate514inter6), .O(gate514inter12));
  nand2 gate2086(.a(gate514inter12), .b(gate514inter1), .O(G1323));
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule