module c880 (N1,N8,N13,N17,N26,N29,N36,N42,N51,N55,
             N59,N68,N72,N73,N74,N75,N80,N85,N86,N87,
             N88,N89,N90,N91,N96,N101,N106,N111,N116,N121,
             N126,N130,N135,N138,N143,N146,N149,N152,N153,N156,
             N159,N165,N171,N177,N183,N189,N195,N201,N207,N210,
             N219,N228,N237,N246,N255,N259,N260,N261,N267,N268,
             N388,N389,N390,N391,N418,N419,N420,N421,N422,N423,
             N446,N447,N448,N449,N450,N767,N768,N850,N863,N864,
             N865,N866,N874,N878,N879,N880);

input N1,N8,N13,N17,N26,N29,N36,N42,N51,N55,
      N59,N68,N72,N73,N74,N75,N80,N85,N86,N87,
      N88,N89,N90,N91,N96,N101,N106,N111,N116,N121,
      N126,N130,N135,N138,N143,N146,N149,N152,N153,N156,
      N159,N165,N171,N177,N183,N189,N195,N201,N207,N210,
      N219,N228,N237,N246,N255,N259,N260,N261,N267,N268;//RE__PI;

input s_0,s_1;//RE__ALLOW(00,01,10,11);
input s_2,s_3;//RE__ALLOW(00,01,10,11);
input s_4,s_5;//RE__ALLOW(00,01,10,11);
input s_6,s_7;//RE__ALLOW(00,01,10,11);
input s_8,s_9;//RE__ALLOW(00,01,10,11);
input s_10,s_11;//RE__ALLOW(00,01,10,11);
input s_12,s_13;//RE__ALLOW(00,01,10,11);
input s_14,s_15;//RE__ALLOW(00,01,10,11);
input s_16,s_17;//RE__ALLOW(00,01,10,11);
input s_18,s_19;//RE__ALLOW(00,01,10,11);
input s_20,s_21;//RE__ALLOW(00,01,10,11);
input s_22,s_23;//RE__ALLOW(00,01,10,11);
input s_24,s_25;//RE__ALLOW(00,01,10,11);
input s_26,s_27;//RE__ALLOW(00,01,10,11);
input s_28,s_29;//RE__ALLOW(00,01,10,11);
input s_30,s_31;//RE__ALLOW(00,01,10,11);
input s_32,s_33;//RE__ALLOW(00,01,10,11);
input s_34,s_35;//RE__ALLOW(00,01,10,11);
input s_36,s_37;//RE__ALLOW(00,01,10,11);
input s_38,s_39;//RE__ALLOW(00,01,10,11);
input s_40,s_41;//RE__ALLOW(00,01,10,11);
input s_42,s_43;//RE__ALLOW(00,01,10,11);
input s_44,s_45;//RE__ALLOW(00,01,10,11);
input s_46,s_47;//RE__ALLOW(00,01,10,11);
input s_48,s_49;//RE__ALLOW(00,01,10,11);
input s_50,s_51;//RE__ALLOW(00,01,10,11);
input s_52,s_53;//RE__ALLOW(00,01,10,11);
input s_54,s_55;//RE__ALLOW(00,01,10,11);
input s_56,s_57;//RE__ALLOW(00,01,10,11);
input s_58,s_59;//RE__ALLOW(00,01,10,11);
input s_60,s_61;//RE__ALLOW(00,01,10,11);
input s_62,s_63;//RE__ALLOW(00,01,10,11);
input s_64,s_65;//RE__ALLOW(00,01,10,11);
input s_66,s_67;//RE__ALLOW(00,01,10,11);
input s_68,s_69;//RE__ALLOW(00,01,10,11);
input s_70,s_71;//RE__ALLOW(00,01,10,11);
output N388,N389,N390,N391,N418,N419,N420,N421,N422,N423,
       N446,N447,N448,N449,N450,N767,N768,N850,N863,N864,
       N865,N866,N874,N878,N879,N880;

wire N269,N270,N273,N276,N279,N280,N284,N285,N286,N287,
     N290,N291,N292,N293,N294,N295,N296,N297,N298,N301,
     N302,N303,N304,N305,N306,N307,N308,N309,N310,N316,
     N317,N318,N319,N322,N323,N324,N325,N326,N327,N328,
     N329,N330,N331,N332,N333,N334,N335,N336,N337,N338,
     N339,N340,N341,N342,N343,N344,N345,N346,N347,N348,
     N349,N350,N351,N352,N353,N354,N355,N356,N357,N360,
     N363,N366,N369,N375,N376,N379,N382,N385,N392,N393,
     N399,N400,N401,N402,N403,N404,N405,N406,N407,N408,
     N409,N410,N411,N412,N413,N414,N415,N416,N417,N424,
     N425,N426,N427,N432,N437,N442,N443,N444,N445,N451,
     N460,N463,N466,N475,N476,N477,N478,N479,N480,N481,
     N482,N483,N488,N489,N490,N491,N492,N495,N498,N499,
     N500,N501,N502,N503,N504,N505,N506,N507,N508,N509,
     N510,N511,N512,N513,N514,N515,N516,N517,N518,N519,
     N520,N521,N522,N523,N524,N525,N526,N527,N528,N529,
     N530,N533,N536,N537,N538,N539,N540,N541,N542,N543,
     N544,N547,N550,N551,N552,N553,N557,N561,N565,N569,
     N573,N577,N581,N585,N586,N587,N588,N589,N590,N593,
     N596,N597,N600,N605,N606,N609,N615,N616,N619,N624,
     N625,N628,N631,N632,N635,N640,N641,N644,N650,N651,
     N654,N659,N660,N661,N662,N665,N669,N670,N673,N677,
     N678,N682,N686,N687,N692,N696,N697,N700,N704,N705,
     N708,N712,N713,N717,N721,N722,N727,N731,N732,N733,
     N734,N735,N736,N737,N738,N739,N740,N741,N742,N743,
     N744,N745,N746,N747,N748,N749,N750,N751,N752,N753,
     N754,N755,N756,N757,N758,N759,N760,N761,N762,N763,
     N764,N765,N766,N769,N770,N771,N772,N773,N777,N778,
     N781,N782,N785,N786,N787,N788,N789,N790,N791,N792,
     N793,N794,N795,N796,N802,N803,N804,N805,N806,N807,
     N808,N809,N810,N811,N812,N813,N814,N815,N819,N822,
     N825,N826,N827,N828,N829,N830,N831,N832,N833,N834,
     N835,N836,N837,N838,N839,N840,N841,N842,N843,N844,
     N845,N846,N847,N848,N849,N851,N852,N853,N854,N855,
     N856,N857,N858,N859,N860,N861,N862,N867,N868,N869,
     N870,N871,N872,N873,N875,N876,N877, gate335inter0, gate335inter1, gate335inter2, gate335inter3, gate335inter4, gate335inter5, gate335inter6, gate335inter7, gate335inter8, gate335inter9, gate335inter10, gate335inter11, gate335inter12, gate346inter0, gate346inter1, gate346inter2, gate346inter3, gate346inter4, gate346inter5, gate346inter6, gate346inter7, gate346inter8, gate346inter9, gate346inter10, gate346inter11, gate346inter12, gate244inter0, gate244inter1, gate244inter2, gate244inter3, gate244inter4, gate244inter5, gate244inter6, gate244inter7, gate244inter8, gate244inter9, gate244inter10, gate244inter11, gate244inter12, gate40inter0, gate40inter1, gate40inter2, gate40inter3, gate40inter4, gate40inter5, gate40inter6, gate40inter7, gate40inter8, gate40inter9, gate40inter10, gate40inter11, gate40inter12, gate67inter0, gate67inter1, gate67inter2, gate67inter3, gate67inter4, gate67inter5, gate67inter6, gate67inter7, gate67inter8, gate67inter9, gate67inter10, gate67inter11, gate67inter12, gate196inter0, gate196inter1, gate196inter2, gate196inter3, gate196inter4, gate196inter5, gate196inter6, gate196inter7, gate196inter8, gate196inter9, gate196inter10, gate196inter11, gate196inter12, gate347inter0, gate347inter1, gate347inter2, gate347inter3, gate347inter4, gate347inter5, gate347inter6, gate347inter7, gate347inter8, gate347inter9, gate347inter10, gate347inter11, gate347inter12, gate193inter0, gate193inter1, gate193inter2, gate193inter3, gate193inter4, gate193inter5, gate193inter6, gate193inter7, gate193inter8, gate193inter9, gate193inter10, gate193inter11, gate193inter12, gate312inter0, gate312inter1, gate312inter2, gate312inter3, gate312inter4, gate312inter5, gate312inter6, gate312inter7, gate312inter8, gate312inter9, gate312inter10, gate312inter11, gate312inter12, gate192inter0, gate192inter1, gate192inter2, gate192inter3, gate192inter4, gate192inter5, gate192inter6, gate192inter7, gate192inter8, gate192inter9, gate192inter10, gate192inter11, gate192inter12, gate69inter0, gate69inter1, gate69inter2, gate69inter3, gate69inter4, gate69inter5, gate69inter6, gate69inter7, gate69inter8, gate69inter9, gate69inter10, gate69inter11, gate69inter12, gate313inter0, gate313inter1, gate313inter2, gate313inter3, gate313inter4, gate313inter5, gate313inter6, gate313inter7, gate313inter8, gate313inter9, gate313inter10, gate313inter11, gate313inter12, gate299inter0, gate299inter1, gate299inter2, gate299inter3, gate299inter4, gate299inter5, gate299inter6, gate299inter7, gate299inter8, gate299inter9, gate299inter10, gate299inter11, gate299inter12, gate247inter0, gate247inter1, gate247inter2, gate247inter3, gate247inter4, gate247inter5, gate247inter6, gate247inter7, gate247inter8, gate247inter9, gate247inter10, gate247inter11, gate247inter12, gate182inter0, gate182inter1, gate182inter2, gate182inter3, gate182inter4, gate182inter5, gate182inter6, gate182inter7, gate182inter8, gate182inter9, gate182inter10, gate182inter11, gate182inter12, gate222inter0, gate222inter1, gate222inter2, gate222inter3, gate222inter4, gate222inter5, gate222inter6, gate222inter7, gate222inter8, gate222inter9, gate222inter10, gate222inter11, gate222inter12, gate173inter0, gate173inter1, gate173inter2, gate173inter3, gate173inter4, gate173inter5, gate173inter6, gate173inter7, gate173inter8, gate173inter9, gate173inter10, gate173inter11, gate173inter12, gate219inter0, gate219inter1, gate219inter2, gate219inter3, gate219inter4, gate219inter5, gate219inter6, gate219inter7, gate219inter8, gate219inter9, gate219inter10, gate219inter11, gate219inter12, gate164inter0, gate164inter1, gate164inter2, gate164inter3, gate164inter4, gate164inter5, gate164inter6, gate164inter7, gate164inter8, gate164inter9, gate164inter10, gate164inter11, gate164inter12, gate364inter0, gate364inter1, gate364inter2, gate364inter3, gate364inter4, gate364inter5, gate364inter6, gate364inter7, gate364inter8, gate364inter9, gate364inter10, gate364inter11, gate364inter12, gate70inter0, gate70inter1, gate70inter2, gate70inter3, gate70inter4, gate70inter5, gate70inter6, gate70inter7, gate70inter8, gate70inter9, gate70inter10, gate70inter11, gate70inter12, gate26inter0, gate26inter1, gate26inter2, gate26inter3, gate26inter4, gate26inter5, gate26inter6, gate26inter7, gate26inter8, gate26inter9, gate26inter10, gate26inter11, gate26inter12, gate72inter0, gate72inter1, gate72inter2, gate72inter3, gate72inter4, gate72inter5, gate72inter6, gate72inter7, gate72inter8, gate72inter9, gate72inter10, gate72inter11, gate72inter12, gate293inter0, gate293inter1, gate293inter2, gate293inter3, gate293inter4, gate293inter5, gate293inter6, gate293inter7, gate293inter8, gate293inter9, gate293inter10, gate293inter11, gate293inter12, gate337inter0, gate337inter1, gate337inter2, gate337inter3, gate337inter4, gate337inter5, gate337inter6, gate337inter7, gate337inter8, gate337inter9, gate337inter10, gate337inter11, gate337inter12, gate175inter0, gate175inter1, gate175inter2, gate175inter3, gate175inter4, gate175inter5, gate175inter6, gate175inter7, gate175inter8, gate175inter9, gate175inter10, gate175inter11, gate175inter12, gate191inter0, gate191inter1, gate191inter2, gate191inter3, gate191inter4, gate191inter5, gate191inter6, gate191inter7, gate191inter8, gate191inter9, gate191inter10, gate191inter11, gate191inter12, gate144inter0, gate144inter1, gate144inter2, gate144inter3, gate144inter4, gate144inter5, gate144inter6, gate144inter7, gate144inter8, gate144inter9, gate144inter10, gate144inter11, gate144inter12, gate36inter0, gate36inter1, gate36inter2, gate36inter3, gate36inter4, gate36inter5, gate36inter6, gate36inter7, gate36inter8, gate36inter9, gate36inter10, gate36inter11, gate36inter12, gate153inter0, gate153inter1, gate153inter2, gate153inter3, gate153inter4, gate153inter5, gate153inter6, gate153inter7, gate153inter8, gate153inter9, gate153inter10, gate153inter11, gate153inter12, gate207inter0, gate207inter1, gate207inter2, gate207inter3, gate207inter4, gate207inter5, gate207inter6, gate207inter7, gate207inter8, gate207inter9, gate207inter10, gate207inter11, gate207inter12, gate22inter0, gate22inter1, gate22inter2, gate22inter3, gate22inter4, gate22inter5, gate22inter6, gate22inter7, gate22inter8, gate22inter9, gate22inter10, gate22inter11, gate22inter12, gate78inter0, gate78inter1, gate78inter2, gate78inter3, gate78inter4, gate78inter5, gate78inter6, gate78inter7, gate78inter8, gate78inter9, gate78inter10, gate78inter11, gate78inter12, gate137inter0, gate137inter1, gate137inter2, gate137inter3, gate137inter4, gate137inter5, gate137inter6, gate137inter7, gate137inter8, gate137inter9, gate137inter10, gate137inter11, gate137inter12, gate310inter0, gate310inter1, gate310inter2, gate310inter3, gate310inter4, gate310inter5, gate310inter6, gate310inter7, gate310inter8, gate310inter9, gate310inter10, gate310inter11, gate310inter12, gate254inter0, gate254inter1, gate254inter2, gate254inter3, gate254inter4, gate254inter5, gate254inter6, gate254inter7, gate254inter8, gate254inter9, gate254inter10, gate254inter11, gate254inter12;



nand4 gate1( .a(N1), .b(N8), .c(N13), .d(N17), .O(N269) );
nand4 gate2( .a(N1), .b(N26), .c(N13), .d(N17), .O(N270) );
and3 gate3( .a(N29), .b(N36), .c(N42), .O(N273) );
and3 gate4( .a(N1), .b(N26), .c(N51), .O(N276) );
nand4 gate5( .a(N1), .b(N8), .c(N51), .d(N17), .O(N279) );
nand4 gate6( .a(N1), .b(N8), .c(N13), .d(N55), .O(N280) );
nand4 gate7( .a(N59), .b(N42), .c(N68), .d(N72), .O(N284) );
nand2 gate8( .a(N29), .b(N68), .O(N285) );
nand3 gate9( .a(N59), .b(N68), .c(N74), .O(N286) );
and3 gate10( .a(N29), .b(N75), .c(N80), .O(N287) );
and3 gate11( .a(N29), .b(N75), .c(N42), .O(N290) );
and3 gate12( .a(N29), .b(N36), .c(N80), .O(N291) );
and3 gate13( .a(N29), .b(N36), .c(N42), .O(N292) );
and3 gate14( .a(N59), .b(N75), .c(N80), .O(N293) );
and3 gate15( .a(N59), .b(N75), .c(N42), .O(N294) );
and3 gate16( .a(N59), .b(N36), .c(N80), .O(N295) );
and3 gate17( .a(N59), .b(N36), .c(N42), .O(N296) );
and2 gate18( .a(N85), .b(N86), .O(N297) );
or2 gate19( .a(N87), .b(N88), .O(N298) );
nand2 gate20( .a(N91), .b(N96), .O(N301) );
or2 gate21( .a(N91), .b(N96), .O(N302) );

  xor2  gate818(.a(N106), .b(N101), .O(gate22inter0));
  nand2 gate819(.a(gate22inter0), .b(s_62), .O(gate22inter1));
  and2  gate820(.a(N106), .b(N101), .O(gate22inter2));
  inv1  gate821(.a(s_62), .O(gate22inter3));
  inv1  gate822(.a(s_63), .O(gate22inter4));
  nand2 gate823(.a(gate22inter4), .b(gate22inter3), .O(gate22inter5));
  nor2  gate824(.a(gate22inter5), .b(gate22inter2), .O(gate22inter6));
  inv1  gate825(.a(N101), .O(gate22inter7));
  inv1  gate826(.a(N106), .O(gate22inter8));
  nand2 gate827(.a(gate22inter8), .b(gate22inter7), .O(gate22inter9));
  nand2 gate828(.a(s_63), .b(gate22inter3), .O(gate22inter10));
  nor2  gate829(.a(gate22inter10), .b(gate22inter9), .O(gate22inter11));
  nor2  gate830(.a(gate22inter11), .b(gate22inter6), .O(gate22inter12));
  nand2 gate831(.a(gate22inter12), .b(gate22inter1), .O(N303));
or2 gate23( .a(N101), .b(N106), .O(N304) );
nand2 gate24( .a(N111), .b(N116), .O(N305) );
or2 gate25( .a(N111), .b(N116), .O(N306) );

  xor2  gate678(.a(N126), .b(N121), .O(gate26inter0));
  nand2 gate679(.a(gate26inter0), .b(s_42), .O(gate26inter1));
  and2  gate680(.a(N126), .b(N121), .O(gate26inter2));
  inv1  gate681(.a(s_42), .O(gate26inter3));
  inv1  gate682(.a(s_43), .O(gate26inter4));
  nand2 gate683(.a(gate26inter4), .b(gate26inter3), .O(gate26inter5));
  nor2  gate684(.a(gate26inter5), .b(gate26inter2), .O(gate26inter6));
  inv1  gate685(.a(N121), .O(gate26inter7));
  inv1  gate686(.a(N126), .O(gate26inter8));
  nand2 gate687(.a(gate26inter8), .b(gate26inter7), .O(gate26inter9));
  nand2 gate688(.a(s_43), .b(gate26inter3), .O(gate26inter10));
  nor2  gate689(.a(gate26inter10), .b(gate26inter9), .O(gate26inter11));
  nor2  gate690(.a(gate26inter11), .b(gate26inter6), .O(gate26inter12));
  nand2 gate691(.a(gate26inter12), .b(gate26inter1), .O(N307));
or2 gate27( .a(N121), .b(N126), .O(N308) );
and2 gate28( .a(N8), .b(N138), .O(N309) );
inv1 gate29( .a(N268), .O(N310) );
and2 gate30( .a(N51), .b(N138), .O(N316) );
and2 gate31( .a(N17), .b(N138), .O(N317) );
and2 gate32( .a(N152), .b(N138), .O(N318) );
nand2 gate33( .a(N59), .b(N156), .O(N319) );
nor2 gate34( .a(N17), .b(N42), .O(N322) );
and2 gate35( .a(N17), .b(N42), .O(N323) );

  xor2  gate776(.a(N165), .b(N159), .O(gate36inter0));
  nand2 gate777(.a(gate36inter0), .b(s_56), .O(gate36inter1));
  and2  gate778(.a(N165), .b(N159), .O(gate36inter2));
  inv1  gate779(.a(s_56), .O(gate36inter3));
  inv1  gate780(.a(s_57), .O(gate36inter4));
  nand2 gate781(.a(gate36inter4), .b(gate36inter3), .O(gate36inter5));
  nor2  gate782(.a(gate36inter5), .b(gate36inter2), .O(gate36inter6));
  inv1  gate783(.a(N159), .O(gate36inter7));
  inv1  gate784(.a(N165), .O(gate36inter8));
  nand2 gate785(.a(gate36inter8), .b(gate36inter7), .O(gate36inter9));
  nand2 gate786(.a(s_57), .b(gate36inter3), .O(gate36inter10));
  nor2  gate787(.a(gate36inter10), .b(gate36inter9), .O(gate36inter11));
  nor2  gate788(.a(gate36inter11), .b(gate36inter6), .O(gate36inter12));
  nand2 gate789(.a(gate36inter12), .b(gate36inter1), .O(N324));
or2 gate37( .a(N159), .b(N165), .O(N325) );
nand2 gate38( .a(N171), .b(N177), .O(N326) );
or2 gate39( .a(N171), .b(N177), .O(N327) );

  xor2  gate426(.a(N189), .b(N183), .O(gate40inter0));
  nand2 gate427(.a(gate40inter0), .b(s_6), .O(gate40inter1));
  and2  gate428(.a(N189), .b(N183), .O(gate40inter2));
  inv1  gate429(.a(s_6), .O(gate40inter3));
  inv1  gate430(.a(s_7), .O(gate40inter4));
  nand2 gate431(.a(gate40inter4), .b(gate40inter3), .O(gate40inter5));
  nor2  gate432(.a(gate40inter5), .b(gate40inter2), .O(gate40inter6));
  inv1  gate433(.a(N183), .O(gate40inter7));
  inv1  gate434(.a(N189), .O(gate40inter8));
  nand2 gate435(.a(gate40inter8), .b(gate40inter7), .O(gate40inter9));
  nand2 gate436(.a(s_7), .b(gate40inter3), .O(gate40inter10));
  nor2  gate437(.a(gate40inter10), .b(gate40inter9), .O(gate40inter11));
  nor2  gate438(.a(gate40inter11), .b(gate40inter6), .O(gate40inter12));
  nand2 gate439(.a(gate40inter12), .b(gate40inter1), .O(N328));
or2 gate41( .a(N183), .b(N189), .O(N329) );
nand2 gate42( .a(N195), .b(N201), .O(N330) );
or2 gate43( .a(N195), .b(N201), .O(N331) );
and2 gate44( .a(N210), .b(N91), .O(N332) );
and2 gate45( .a(N210), .b(N96), .O(N333) );
and2 gate46( .a(N210), .b(N101), .O(N334) );
and2 gate47( .a(N210), .b(N106), .O(N335) );
and2 gate48( .a(N210), .b(N111), .O(N336) );
and2 gate49( .a(N255), .b(N259), .O(N337) );
and2 gate50( .a(N210), .b(N116), .O(N338) );
and2 gate51( .a(N255), .b(N260), .O(N339) );
and2 gate52( .a(N210), .b(N121), .O(N340) );
and2 gate53( .a(N255), .b(N267), .O(N341) );
inv1 gate54( .a(N269), .O(N342) );
inv1 gate55( .a(N273), .O(N343) );
or2 gate56( .a(N270), .b(N273), .O(N344) );
inv1 gate57( .a(N276), .O(N345) );
inv1 gate58( .a(N276), .O(N346) );
inv1 gate59( .a(N279), .O(N347) );
nor2 gate60( .a(N280), .b(N284), .O(N348) );
or2 gate61( .a(N280), .b(N285), .O(N349) );
or2 gate62( .a(N280), .b(N286), .O(N350) );
inv1 gate63( .a(N293), .O(N351) );
inv1 gate64( .a(N294), .O(N352) );
inv1 gate65( .a(N295), .O(N353) );
inv1 gate66( .a(N296), .O(N354) );

  xor2  gate440(.a(N298), .b(N89), .O(gate67inter0));
  nand2 gate441(.a(gate67inter0), .b(s_8), .O(gate67inter1));
  and2  gate442(.a(N298), .b(N89), .O(gate67inter2));
  inv1  gate443(.a(s_8), .O(gate67inter3));
  inv1  gate444(.a(s_9), .O(gate67inter4));
  nand2 gate445(.a(gate67inter4), .b(gate67inter3), .O(gate67inter5));
  nor2  gate446(.a(gate67inter5), .b(gate67inter2), .O(gate67inter6));
  inv1  gate447(.a(N89), .O(gate67inter7));
  inv1  gate448(.a(N298), .O(gate67inter8));
  nand2 gate449(.a(gate67inter8), .b(gate67inter7), .O(gate67inter9));
  nand2 gate450(.a(s_9), .b(gate67inter3), .O(gate67inter10));
  nor2  gate451(.a(gate67inter10), .b(gate67inter9), .O(gate67inter11));
  nor2  gate452(.a(gate67inter11), .b(gate67inter6), .O(gate67inter12));
  nand2 gate453(.a(gate67inter12), .b(gate67inter1), .O(N355));
and2 gate68( .a(N90), .b(N298), .O(N356) );

  xor2  gate524(.a(N302), .b(N301), .O(gate69inter0));
  nand2 gate525(.a(gate69inter0), .b(s_20), .O(gate69inter1));
  and2  gate526(.a(N302), .b(N301), .O(gate69inter2));
  inv1  gate527(.a(s_20), .O(gate69inter3));
  inv1  gate528(.a(s_21), .O(gate69inter4));
  nand2 gate529(.a(gate69inter4), .b(gate69inter3), .O(gate69inter5));
  nor2  gate530(.a(gate69inter5), .b(gate69inter2), .O(gate69inter6));
  inv1  gate531(.a(N301), .O(gate69inter7));
  inv1  gate532(.a(N302), .O(gate69inter8));
  nand2 gate533(.a(gate69inter8), .b(gate69inter7), .O(gate69inter9));
  nand2 gate534(.a(s_21), .b(gate69inter3), .O(gate69inter10));
  nor2  gate535(.a(gate69inter10), .b(gate69inter9), .O(gate69inter11));
  nor2  gate536(.a(gate69inter11), .b(gate69inter6), .O(gate69inter12));
  nand2 gate537(.a(gate69inter12), .b(gate69inter1), .O(N357));

  xor2  gate664(.a(N304), .b(N303), .O(gate70inter0));
  nand2 gate665(.a(gate70inter0), .b(s_40), .O(gate70inter1));
  and2  gate666(.a(N304), .b(N303), .O(gate70inter2));
  inv1  gate667(.a(s_40), .O(gate70inter3));
  inv1  gate668(.a(s_41), .O(gate70inter4));
  nand2 gate669(.a(gate70inter4), .b(gate70inter3), .O(gate70inter5));
  nor2  gate670(.a(gate70inter5), .b(gate70inter2), .O(gate70inter6));
  inv1  gate671(.a(N303), .O(gate70inter7));
  inv1  gate672(.a(N304), .O(gate70inter8));
  nand2 gate673(.a(gate70inter8), .b(gate70inter7), .O(gate70inter9));
  nand2 gate674(.a(s_41), .b(gate70inter3), .O(gate70inter10));
  nor2  gate675(.a(gate70inter10), .b(gate70inter9), .O(gate70inter11));
  nor2  gate676(.a(gate70inter11), .b(gate70inter6), .O(gate70inter12));
  nand2 gate677(.a(gate70inter12), .b(gate70inter1), .O(N360));
nand2 gate71( .a(N305), .b(N306), .O(N363) );

  xor2  gate692(.a(N308), .b(N307), .O(gate72inter0));
  nand2 gate693(.a(gate72inter0), .b(s_44), .O(gate72inter1));
  and2  gate694(.a(N308), .b(N307), .O(gate72inter2));
  inv1  gate695(.a(s_44), .O(gate72inter3));
  inv1  gate696(.a(s_45), .O(gate72inter4));
  nand2 gate697(.a(gate72inter4), .b(gate72inter3), .O(gate72inter5));
  nor2  gate698(.a(gate72inter5), .b(gate72inter2), .O(gate72inter6));
  inv1  gate699(.a(N307), .O(gate72inter7));
  inv1  gate700(.a(N308), .O(gate72inter8));
  nand2 gate701(.a(gate72inter8), .b(gate72inter7), .O(gate72inter9));
  nand2 gate702(.a(s_45), .b(gate72inter3), .O(gate72inter10));
  nor2  gate703(.a(gate72inter10), .b(gate72inter9), .O(gate72inter11));
  nor2  gate704(.a(gate72inter11), .b(gate72inter6), .O(gate72inter12));
  nand2 gate705(.a(gate72inter12), .b(gate72inter1), .O(N366));
inv1 gate73( .a(N310), .O(N369) );
nor2 gate74( .a(N322), .b(N323), .O(N375) );
nand2 gate75( .a(N324), .b(N325), .O(N376) );
nand2 gate76( .a(N326), .b(N327), .O(N379) );
nand2 gate77( .a(N328), .b(N329), .O(N382) );

  xor2  gate832(.a(N331), .b(N330), .O(gate78inter0));
  nand2 gate833(.a(gate78inter0), .b(s_64), .O(gate78inter1));
  and2  gate834(.a(N331), .b(N330), .O(gate78inter2));
  inv1  gate835(.a(s_64), .O(gate78inter3));
  inv1  gate836(.a(s_65), .O(gate78inter4));
  nand2 gate837(.a(gate78inter4), .b(gate78inter3), .O(gate78inter5));
  nor2  gate838(.a(gate78inter5), .b(gate78inter2), .O(gate78inter6));
  inv1  gate839(.a(N330), .O(gate78inter7));
  inv1  gate840(.a(N331), .O(gate78inter8));
  nand2 gate841(.a(gate78inter8), .b(gate78inter7), .O(gate78inter9));
  nand2 gate842(.a(s_65), .b(gate78inter3), .O(gate78inter10));
  nor2  gate843(.a(gate78inter10), .b(gate78inter9), .O(gate78inter11));
  nor2  gate844(.a(gate78inter11), .b(gate78inter6), .O(gate78inter12));
  nand2 gate845(.a(gate78inter12), .b(gate78inter1), .O(N385));
buf1 gate79( .a(N290), .O(N388) );
buf1 gate80( .a(N291), .O(N389) );
buf1 gate81( .a(N292), .O(N390) );
buf1 gate82( .a(N297), .O(N391) );
or2 gate83( .a(N270), .b(N343), .O(N392) );
inv1 gate84( .a(N345), .O(N393) );
inv1 gate85( .a(N346), .O(N399) );
and2 gate86( .a(N348), .b(N73), .O(N400) );
inv1 gate87( .a(N349), .O(N401) );
inv1 gate88( .a(N350), .O(N402) );
inv1 gate89( .a(N355), .O(N403) );
inv1 gate90( .a(N357), .O(N404) );
inv1 gate91( .a(N360), .O(N405) );
and2 gate92( .a(N357), .b(N360), .O(N406) );
inv1 gate93( .a(N363), .O(N407) );
inv1 gate94( .a(N366), .O(N408) );
and2 gate95( .a(N363), .b(N366), .O(N409) );
nand2 gate96( .a(N347), .b(N352), .O(N410) );
inv1 gate97( .a(N376), .O(N411) );
inv1 gate98( .a(N379), .O(N412) );
and2 gate99( .a(N376), .b(N379), .O(N413) );
inv1 gate100( .a(N382), .O(N414) );
inv1 gate101( .a(N385), .O(N415) );
and2 gate102( .a(N382), .b(N385), .O(N416) );
and2 gate103( .a(N210), .b(N369), .O(N417) );
buf1 gate104( .a(N342), .O(N418) );
buf1 gate105( .a(N344), .O(N419) );
buf1 gate106( .a(N351), .O(N420) );
buf1 gate107( .a(N353), .O(N421) );
buf1 gate108( .a(N354), .O(N422) );
buf1 gate109( .a(N356), .O(N423) );
inv1 gate110( .a(N400), .O(N424) );
and2 gate111( .a(N404), .b(N405), .O(N425) );
and2 gate112( .a(N407), .b(N408), .O(N426) );
and3 gate113( .a(N319), .b(N393), .c(N55), .O(N427) );
and3 gate114( .a(N393), .b(N17), .c(N287), .O(N432) );
nand3 gate115( .a(N393), .b(N287), .c(N55), .O(N437) );
nand4 gate116( .a(N375), .b(N59), .c(N156), .d(N393), .O(N442) );
nand3 gate117( .a(N393), .b(N319), .c(N17), .O(N443) );
and2 gate118( .a(N411), .b(N412), .O(N444) );
and2 gate119( .a(N414), .b(N415), .O(N445) );
buf1 gate120( .a(N392), .O(N446) );
buf1 gate121( .a(N399), .O(N447) );
buf1 gate122( .a(N401), .O(N448) );
buf1 gate123( .a(N402), .O(N449) );
buf1 gate124( .a(N403), .O(N450) );
inv1 gate125( .a(N424), .O(N451) );
nor2 gate126( .a(N406), .b(N425), .O(N460) );
nor2 gate127( .a(N409), .b(N426), .O(N463) );
nand2 gate128( .a(N442), .b(N410), .O(N466) );
and2 gate129( .a(N143), .b(N427), .O(N475) );
and2 gate130( .a(N310), .b(N432), .O(N476) );
and2 gate131( .a(N146), .b(N427), .O(N477) );
and2 gate132( .a(N310), .b(N432), .O(N478) );
and2 gate133( .a(N149), .b(N427), .O(N479) );
and2 gate134( .a(N310), .b(N432), .O(N480) );
and2 gate135( .a(N153), .b(N427), .O(N481) );
and2 gate136( .a(N310), .b(N432), .O(N482) );

  xor2  gate846(.a(N1), .b(N443), .O(gate137inter0));
  nand2 gate847(.a(gate137inter0), .b(s_66), .O(gate137inter1));
  and2  gate848(.a(N1), .b(N443), .O(gate137inter2));
  inv1  gate849(.a(s_66), .O(gate137inter3));
  inv1  gate850(.a(s_67), .O(gate137inter4));
  nand2 gate851(.a(gate137inter4), .b(gate137inter3), .O(gate137inter5));
  nor2  gate852(.a(gate137inter5), .b(gate137inter2), .O(gate137inter6));
  inv1  gate853(.a(N443), .O(gate137inter7));
  inv1  gate854(.a(N1), .O(gate137inter8));
  nand2 gate855(.a(gate137inter8), .b(gate137inter7), .O(gate137inter9));
  nand2 gate856(.a(s_67), .b(gate137inter3), .O(gate137inter10));
  nor2  gate857(.a(gate137inter10), .b(gate137inter9), .O(gate137inter11));
  nor2  gate858(.a(gate137inter11), .b(gate137inter6), .O(gate137inter12));
  nand2 gate859(.a(gate137inter12), .b(gate137inter1), .O(N483));
or2 gate138( .a(N369), .b(N437), .O(N488) );
or2 gate139( .a(N369), .b(N437), .O(N489) );
or2 gate140( .a(N369), .b(N437), .O(N490) );
or2 gate141( .a(N369), .b(N437), .O(N491) );
nor2 gate142( .a(N413), .b(N444), .O(N492) );
nor2 gate143( .a(N416), .b(N445), .O(N495) );

  xor2  gate762(.a(N460), .b(N130), .O(gate144inter0));
  nand2 gate763(.a(gate144inter0), .b(s_54), .O(gate144inter1));
  and2  gate764(.a(N460), .b(N130), .O(gate144inter2));
  inv1  gate765(.a(s_54), .O(gate144inter3));
  inv1  gate766(.a(s_55), .O(gate144inter4));
  nand2 gate767(.a(gate144inter4), .b(gate144inter3), .O(gate144inter5));
  nor2  gate768(.a(gate144inter5), .b(gate144inter2), .O(gate144inter6));
  inv1  gate769(.a(N130), .O(gate144inter7));
  inv1  gate770(.a(N460), .O(gate144inter8));
  nand2 gate771(.a(gate144inter8), .b(gate144inter7), .O(gate144inter9));
  nand2 gate772(.a(s_55), .b(gate144inter3), .O(gate144inter10));
  nor2  gate773(.a(gate144inter10), .b(gate144inter9), .O(gate144inter11));
  nor2  gate774(.a(gate144inter11), .b(gate144inter6), .O(gate144inter12));
  nand2 gate775(.a(gate144inter12), .b(gate144inter1), .O(N498));
or2 gate145( .a(N130), .b(N460), .O(N499) );
nand2 gate146( .a(N463), .b(N135), .O(N500) );
or2 gate147( .a(N463), .b(N135), .O(N501) );
and2 gate148( .a(N91), .b(N466), .O(N502) );
nor2 gate149( .a(N475), .b(N476), .O(N503) );
and2 gate150( .a(N96), .b(N466), .O(N504) );
nor2 gate151( .a(N477), .b(N478), .O(N505) );
and2 gate152( .a(N101), .b(N466), .O(N506) );

  xor2  gate790(.a(N480), .b(N479), .O(gate153inter0));
  nand2 gate791(.a(gate153inter0), .b(s_58), .O(gate153inter1));
  and2  gate792(.a(N480), .b(N479), .O(gate153inter2));
  inv1  gate793(.a(s_58), .O(gate153inter3));
  inv1  gate794(.a(s_59), .O(gate153inter4));
  nand2 gate795(.a(gate153inter4), .b(gate153inter3), .O(gate153inter5));
  nor2  gate796(.a(gate153inter5), .b(gate153inter2), .O(gate153inter6));
  inv1  gate797(.a(N479), .O(gate153inter7));
  inv1  gate798(.a(N480), .O(gate153inter8));
  nand2 gate799(.a(gate153inter8), .b(gate153inter7), .O(gate153inter9));
  nand2 gate800(.a(s_59), .b(gate153inter3), .O(gate153inter10));
  nor2  gate801(.a(gate153inter10), .b(gate153inter9), .O(gate153inter11));
  nor2  gate802(.a(gate153inter11), .b(gate153inter6), .O(gate153inter12));
  nand2 gate803(.a(gate153inter12), .b(gate153inter1), .O(N507));
and2 gate154( .a(N106), .b(N466), .O(N508) );
nor2 gate155( .a(N481), .b(N482), .O(N509) );
and2 gate156( .a(N143), .b(N483), .O(N510) );
and2 gate157( .a(N111), .b(N466), .O(N511) );
and2 gate158( .a(N146), .b(N483), .O(N512) );
and2 gate159( .a(N116), .b(N466), .O(N513) );
and2 gate160( .a(N149), .b(N483), .O(N514) );
and2 gate161( .a(N121), .b(N466), .O(N515) );
and2 gate162( .a(N153), .b(N483), .O(N516) );
and2 gate163( .a(N126), .b(N466), .O(N517) );

  xor2  gate636(.a(N492), .b(N130), .O(gate164inter0));
  nand2 gate637(.a(gate164inter0), .b(s_36), .O(gate164inter1));
  and2  gate638(.a(N492), .b(N130), .O(gate164inter2));
  inv1  gate639(.a(s_36), .O(gate164inter3));
  inv1  gate640(.a(s_37), .O(gate164inter4));
  nand2 gate641(.a(gate164inter4), .b(gate164inter3), .O(gate164inter5));
  nor2  gate642(.a(gate164inter5), .b(gate164inter2), .O(gate164inter6));
  inv1  gate643(.a(N130), .O(gate164inter7));
  inv1  gate644(.a(N492), .O(gate164inter8));
  nand2 gate645(.a(gate164inter8), .b(gate164inter7), .O(gate164inter9));
  nand2 gate646(.a(s_37), .b(gate164inter3), .O(gate164inter10));
  nor2  gate647(.a(gate164inter10), .b(gate164inter9), .O(gate164inter11));
  nor2  gate648(.a(gate164inter11), .b(gate164inter6), .O(gate164inter12));
  nand2 gate649(.a(gate164inter12), .b(gate164inter1), .O(N518));
or2 gate165( .a(N130), .b(N492), .O(N519) );
nand2 gate166( .a(N495), .b(N207), .O(N520) );
or2 gate167( .a(N495), .b(N207), .O(N521) );
and2 gate168( .a(N451), .b(N159), .O(N522) );
and2 gate169( .a(N451), .b(N165), .O(N523) );
and2 gate170( .a(N451), .b(N171), .O(N524) );
and2 gate171( .a(N451), .b(N177), .O(N525) );
and2 gate172( .a(N451), .b(N183), .O(N526) );

  xor2  gate608(.a(N189), .b(N451), .O(gate173inter0));
  nand2 gate609(.a(gate173inter0), .b(s_32), .O(gate173inter1));
  and2  gate610(.a(N189), .b(N451), .O(gate173inter2));
  inv1  gate611(.a(s_32), .O(gate173inter3));
  inv1  gate612(.a(s_33), .O(gate173inter4));
  nand2 gate613(.a(gate173inter4), .b(gate173inter3), .O(gate173inter5));
  nor2  gate614(.a(gate173inter5), .b(gate173inter2), .O(gate173inter6));
  inv1  gate615(.a(N451), .O(gate173inter7));
  inv1  gate616(.a(N189), .O(gate173inter8));
  nand2 gate617(.a(gate173inter8), .b(gate173inter7), .O(gate173inter9));
  nand2 gate618(.a(s_33), .b(gate173inter3), .O(gate173inter10));
  nor2  gate619(.a(gate173inter10), .b(gate173inter9), .O(gate173inter11));
  nor2  gate620(.a(gate173inter11), .b(gate173inter6), .O(gate173inter12));
  nand2 gate621(.a(gate173inter12), .b(gate173inter1), .O(N527));
nand2 gate174( .a(N451), .b(N195), .O(N528) );

  xor2  gate734(.a(N201), .b(N451), .O(gate175inter0));
  nand2 gate735(.a(gate175inter0), .b(s_50), .O(gate175inter1));
  and2  gate736(.a(N201), .b(N451), .O(gate175inter2));
  inv1  gate737(.a(s_50), .O(gate175inter3));
  inv1  gate738(.a(s_51), .O(gate175inter4));
  nand2 gate739(.a(gate175inter4), .b(gate175inter3), .O(gate175inter5));
  nor2  gate740(.a(gate175inter5), .b(gate175inter2), .O(gate175inter6));
  inv1  gate741(.a(N451), .O(gate175inter7));
  inv1  gate742(.a(N201), .O(gate175inter8));
  nand2 gate743(.a(gate175inter8), .b(gate175inter7), .O(gate175inter9));
  nand2 gate744(.a(s_51), .b(gate175inter3), .O(gate175inter10));
  nor2  gate745(.a(gate175inter10), .b(gate175inter9), .O(gate175inter11));
  nor2  gate746(.a(gate175inter11), .b(gate175inter6), .O(gate175inter12));
  nand2 gate747(.a(gate175inter12), .b(gate175inter1), .O(N529));
nand2 gate176( .a(N498), .b(N499), .O(N530) );
nand2 gate177( .a(N500), .b(N501), .O(N533) );
nor2 gate178( .a(N309), .b(N502), .O(N536) );
nor2 gate179( .a(N316), .b(N504), .O(N537) );
nor2 gate180( .a(N317), .b(N506), .O(N538) );
nor2 gate181( .a(N318), .b(N508), .O(N539) );

  xor2  gate580(.a(N511), .b(N510), .O(gate182inter0));
  nand2 gate581(.a(gate182inter0), .b(s_28), .O(gate182inter1));
  and2  gate582(.a(N511), .b(N510), .O(gate182inter2));
  inv1  gate583(.a(s_28), .O(gate182inter3));
  inv1  gate584(.a(s_29), .O(gate182inter4));
  nand2 gate585(.a(gate182inter4), .b(gate182inter3), .O(gate182inter5));
  nor2  gate586(.a(gate182inter5), .b(gate182inter2), .O(gate182inter6));
  inv1  gate587(.a(N510), .O(gate182inter7));
  inv1  gate588(.a(N511), .O(gate182inter8));
  nand2 gate589(.a(gate182inter8), .b(gate182inter7), .O(gate182inter9));
  nand2 gate590(.a(s_29), .b(gate182inter3), .O(gate182inter10));
  nor2  gate591(.a(gate182inter10), .b(gate182inter9), .O(gate182inter11));
  nor2  gate592(.a(gate182inter11), .b(gate182inter6), .O(gate182inter12));
  nand2 gate593(.a(gate182inter12), .b(gate182inter1), .O(N540));
nor2 gate183( .a(N512), .b(N513), .O(N541) );
nor2 gate184( .a(N514), .b(N515), .O(N542) );
nor2 gate185( .a(N516), .b(N517), .O(N543) );
nand2 gate186( .a(N518), .b(N519), .O(N544) );
nand2 gate187( .a(N520), .b(N521), .O(N547) );
inv1 gate188( .a(N530), .O(N550) );
inv1 gate189( .a(N533), .O(N551) );
and2 gate190( .a(N530), .b(N533), .O(N552) );

  xor2  gate748(.a(N503), .b(N536), .O(gate191inter0));
  nand2 gate749(.a(gate191inter0), .b(s_52), .O(gate191inter1));
  and2  gate750(.a(N503), .b(N536), .O(gate191inter2));
  inv1  gate751(.a(s_52), .O(gate191inter3));
  inv1  gate752(.a(s_53), .O(gate191inter4));
  nand2 gate753(.a(gate191inter4), .b(gate191inter3), .O(gate191inter5));
  nor2  gate754(.a(gate191inter5), .b(gate191inter2), .O(gate191inter6));
  inv1  gate755(.a(N536), .O(gate191inter7));
  inv1  gate756(.a(N503), .O(gate191inter8));
  nand2 gate757(.a(gate191inter8), .b(gate191inter7), .O(gate191inter9));
  nand2 gate758(.a(s_53), .b(gate191inter3), .O(gate191inter10));
  nor2  gate759(.a(gate191inter10), .b(gate191inter9), .O(gate191inter11));
  nor2  gate760(.a(gate191inter11), .b(gate191inter6), .O(gate191inter12));
  nand2 gate761(.a(gate191inter12), .b(gate191inter1), .O(N553));

  xor2  gate510(.a(N505), .b(N537), .O(gate192inter0));
  nand2 gate511(.a(gate192inter0), .b(s_18), .O(gate192inter1));
  and2  gate512(.a(N505), .b(N537), .O(gate192inter2));
  inv1  gate513(.a(s_18), .O(gate192inter3));
  inv1  gate514(.a(s_19), .O(gate192inter4));
  nand2 gate515(.a(gate192inter4), .b(gate192inter3), .O(gate192inter5));
  nor2  gate516(.a(gate192inter5), .b(gate192inter2), .O(gate192inter6));
  inv1  gate517(.a(N537), .O(gate192inter7));
  inv1  gate518(.a(N505), .O(gate192inter8));
  nand2 gate519(.a(gate192inter8), .b(gate192inter7), .O(gate192inter9));
  nand2 gate520(.a(s_19), .b(gate192inter3), .O(gate192inter10));
  nor2  gate521(.a(gate192inter10), .b(gate192inter9), .O(gate192inter11));
  nor2  gate522(.a(gate192inter11), .b(gate192inter6), .O(gate192inter12));
  nand2 gate523(.a(gate192inter12), .b(gate192inter1), .O(N557));

  xor2  gate482(.a(N507), .b(N538), .O(gate193inter0));
  nand2 gate483(.a(gate193inter0), .b(s_14), .O(gate193inter1));
  and2  gate484(.a(N507), .b(N538), .O(gate193inter2));
  inv1  gate485(.a(s_14), .O(gate193inter3));
  inv1  gate486(.a(s_15), .O(gate193inter4));
  nand2 gate487(.a(gate193inter4), .b(gate193inter3), .O(gate193inter5));
  nor2  gate488(.a(gate193inter5), .b(gate193inter2), .O(gate193inter6));
  inv1  gate489(.a(N538), .O(gate193inter7));
  inv1  gate490(.a(N507), .O(gate193inter8));
  nand2 gate491(.a(gate193inter8), .b(gate193inter7), .O(gate193inter9));
  nand2 gate492(.a(s_15), .b(gate193inter3), .O(gate193inter10));
  nor2  gate493(.a(gate193inter10), .b(gate193inter9), .O(gate193inter11));
  nor2  gate494(.a(gate193inter11), .b(gate193inter6), .O(gate193inter12));
  nand2 gate495(.a(gate193inter12), .b(gate193inter1), .O(N561));
nand2 gate194( .a(N539), .b(N509), .O(N565) );
nand2 gate195( .a(N488), .b(N540), .O(N569) );

  xor2  gate454(.a(N541), .b(N489), .O(gate196inter0));
  nand2 gate455(.a(gate196inter0), .b(s_10), .O(gate196inter1));
  and2  gate456(.a(N541), .b(N489), .O(gate196inter2));
  inv1  gate457(.a(s_10), .O(gate196inter3));
  inv1  gate458(.a(s_11), .O(gate196inter4));
  nand2 gate459(.a(gate196inter4), .b(gate196inter3), .O(gate196inter5));
  nor2  gate460(.a(gate196inter5), .b(gate196inter2), .O(gate196inter6));
  inv1  gate461(.a(N489), .O(gate196inter7));
  inv1  gate462(.a(N541), .O(gate196inter8));
  nand2 gate463(.a(gate196inter8), .b(gate196inter7), .O(gate196inter9));
  nand2 gate464(.a(s_11), .b(gate196inter3), .O(gate196inter10));
  nor2  gate465(.a(gate196inter10), .b(gate196inter9), .O(gate196inter11));
  nor2  gate466(.a(gate196inter11), .b(gate196inter6), .O(gate196inter12));
  nand2 gate467(.a(gate196inter12), .b(gate196inter1), .O(N573));
nand2 gate197( .a(N490), .b(N542), .O(N577) );
nand2 gate198( .a(N491), .b(N543), .O(N581) );
inv1 gate199( .a(N544), .O(N585) );
inv1 gate200( .a(N547), .O(N586) );
and2 gate201( .a(N544), .b(N547), .O(N587) );
and2 gate202( .a(N550), .b(N551), .O(N588) );
and2 gate203( .a(N585), .b(N586), .O(N589) );
nand2 gate204( .a(N553), .b(N159), .O(N590) );
or2 gate205( .a(N553), .b(N159), .O(N593) );
and2 gate206( .a(N246), .b(N553), .O(N596) );

  xor2  gate804(.a(N165), .b(N557), .O(gate207inter0));
  nand2 gate805(.a(gate207inter0), .b(s_60), .O(gate207inter1));
  and2  gate806(.a(N165), .b(N557), .O(gate207inter2));
  inv1  gate807(.a(s_60), .O(gate207inter3));
  inv1  gate808(.a(s_61), .O(gate207inter4));
  nand2 gate809(.a(gate207inter4), .b(gate207inter3), .O(gate207inter5));
  nor2  gate810(.a(gate207inter5), .b(gate207inter2), .O(gate207inter6));
  inv1  gate811(.a(N557), .O(gate207inter7));
  inv1  gate812(.a(N165), .O(gate207inter8));
  nand2 gate813(.a(gate207inter8), .b(gate207inter7), .O(gate207inter9));
  nand2 gate814(.a(s_61), .b(gate207inter3), .O(gate207inter10));
  nor2  gate815(.a(gate207inter10), .b(gate207inter9), .O(gate207inter11));
  nor2  gate816(.a(gate207inter11), .b(gate207inter6), .O(gate207inter12));
  nand2 gate817(.a(gate207inter12), .b(gate207inter1), .O(N597));
or2 gate208( .a(N557), .b(N165), .O(N600) );
and2 gate209( .a(N246), .b(N557), .O(N605) );
nand2 gate210( .a(N561), .b(N171), .O(N606) );
or2 gate211( .a(N561), .b(N171), .O(N609) );
and2 gate212( .a(N246), .b(N561), .O(N615) );
nand2 gate213( .a(N565), .b(N177), .O(N616) );
or2 gate214( .a(N565), .b(N177), .O(N619) );
and2 gate215( .a(N246), .b(N565), .O(N624) );
nand2 gate216( .a(N569), .b(N183), .O(N625) );
or2 gate217( .a(N569), .b(N183), .O(N628) );
and2 gate218( .a(N246), .b(N569), .O(N631) );

  xor2  gate622(.a(N189), .b(N573), .O(gate219inter0));
  nand2 gate623(.a(gate219inter0), .b(s_34), .O(gate219inter1));
  and2  gate624(.a(N189), .b(N573), .O(gate219inter2));
  inv1  gate625(.a(s_34), .O(gate219inter3));
  inv1  gate626(.a(s_35), .O(gate219inter4));
  nand2 gate627(.a(gate219inter4), .b(gate219inter3), .O(gate219inter5));
  nor2  gate628(.a(gate219inter5), .b(gate219inter2), .O(gate219inter6));
  inv1  gate629(.a(N573), .O(gate219inter7));
  inv1  gate630(.a(N189), .O(gate219inter8));
  nand2 gate631(.a(gate219inter8), .b(gate219inter7), .O(gate219inter9));
  nand2 gate632(.a(s_35), .b(gate219inter3), .O(gate219inter10));
  nor2  gate633(.a(gate219inter10), .b(gate219inter9), .O(gate219inter11));
  nor2  gate634(.a(gate219inter11), .b(gate219inter6), .O(gate219inter12));
  nand2 gate635(.a(gate219inter12), .b(gate219inter1), .O(N632));
or2 gate220( .a(N573), .b(N189), .O(N635) );
and2 gate221( .a(N246), .b(N573), .O(N640) );

  xor2  gate594(.a(N195), .b(N577), .O(gate222inter0));
  nand2 gate595(.a(gate222inter0), .b(s_30), .O(gate222inter1));
  and2  gate596(.a(N195), .b(N577), .O(gate222inter2));
  inv1  gate597(.a(s_30), .O(gate222inter3));
  inv1  gate598(.a(s_31), .O(gate222inter4));
  nand2 gate599(.a(gate222inter4), .b(gate222inter3), .O(gate222inter5));
  nor2  gate600(.a(gate222inter5), .b(gate222inter2), .O(gate222inter6));
  inv1  gate601(.a(N577), .O(gate222inter7));
  inv1  gate602(.a(N195), .O(gate222inter8));
  nand2 gate603(.a(gate222inter8), .b(gate222inter7), .O(gate222inter9));
  nand2 gate604(.a(s_31), .b(gate222inter3), .O(gate222inter10));
  nor2  gate605(.a(gate222inter10), .b(gate222inter9), .O(gate222inter11));
  nor2  gate606(.a(gate222inter11), .b(gate222inter6), .O(gate222inter12));
  nand2 gate607(.a(gate222inter12), .b(gate222inter1), .O(N641));
or2 gate223( .a(N577), .b(N195), .O(N644) );
and2 gate224( .a(N246), .b(N577), .O(N650) );
nand2 gate225( .a(N581), .b(N201), .O(N651) );
or2 gate226( .a(N581), .b(N201), .O(N654) );
and2 gate227( .a(N246), .b(N581), .O(N659) );
nor2 gate228( .a(N552), .b(N588), .O(N660) );
nor2 gate229( .a(N587), .b(N589), .O(N661) );
inv1 gate230( .a(N590), .O(N662) );
and2 gate231( .a(N593), .b(N590), .O(N665) );
nor2 gate232( .a(N596), .b(N522), .O(N669) );
inv1 gate233( .a(N597), .O(N670) );
and2 gate234( .a(N600), .b(N597), .O(N673) );
nor2 gate235( .a(N605), .b(N523), .O(N677) );
inv1 gate236( .a(N606), .O(N678) );
and2 gate237( .a(N609), .b(N606), .O(N682) );
nor2 gate238( .a(N615), .b(N524), .O(N686) );
inv1 gate239( .a(N616), .O(N687) );
and2 gate240( .a(N619), .b(N616), .O(N692) );
nor2 gate241( .a(N624), .b(N525), .O(N696) );
inv1 gate242( .a(N625), .O(N697) );
and2 gate243( .a(N628), .b(N625), .O(N700) );

  xor2  gate412(.a(N526), .b(N631), .O(gate244inter0));
  nand2 gate413(.a(gate244inter0), .b(s_4), .O(gate244inter1));
  and2  gate414(.a(N526), .b(N631), .O(gate244inter2));
  inv1  gate415(.a(s_4), .O(gate244inter3));
  inv1  gate416(.a(s_5), .O(gate244inter4));
  nand2 gate417(.a(gate244inter4), .b(gate244inter3), .O(gate244inter5));
  nor2  gate418(.a(gate244inter5), .b(gate244inter2), .O(gate244inter6));
  inv1  gate419(.a(N631), .O(gate244inter7));
  inv1  gate420(.a(N526), .O(gate244inter8));
  nand2 gate421(.a(gate244inter8), .b(gate244inter7), .O(gate244inter9));
  nand2 gate422(.a(s_5), .b(gate244inter3), .O(gate244inter10));
  nor2  gate423(.a(gate244inter10), .b(gate244inter9), .O(gate244inter11));
  nor2  gate424(.a(gate244inter11), .b(gate244inter6), .O(gate244inter12));
  nand2 gate425(.a(gate244inter12), .b(gate244inter1), .O(N704));
inv1 gate245( .a(N632), .O(N705) );
and2 gate246( .a(N635), .b(N632), .O(N708) );

  xor2  gate566(.a(N640), .b(N337), .O(gate247inter0));
  nand2 gate567(.a(gate247inter0), .b(s_26), .O(gate247inter1));
  and2  gate568(.a(N640), .b(N337), .O(gate247inter2));
  inv1  gate569(.a(s_26), .O(gate247inter3));
  inv1  gate570(.a(s_27), .O(gate247inter4));
  nand2 gate571(.a(gate247inter4), .b(gate247inter3), .O(gate247inter5));
  nor2  gate572(.a(gate247inter5), .b(gate247inter2), .O(gate247inter6));
  inv1  gate573(.a(N337), .O(gate247inter7));
  inv1  gate574(.a(N640), .O(gate247inter8));
  nand2 gate575(.a(gate247inter8), .b(gate247inter7), .O(gate247inter9));
  nand2 gate576(.a(s_27), .b(gate247inter3), .O(gate247inter10));
  nor2  gate577(.a(gate247inter10), .b(gate247inter9), .O(gate247inter11));
  nor2  gate578(.a(gate247inter11), .b(gate247inter6), .O(gate247inter12));
  nand2 gate579(.a(gate247inter12), .b(gate247inter1), .O(N712));
inv1 gate248( .a(N641), .O(N713) );
and2 gate249( .a(N644), .b(N641), .O(N717) );
nor2 gate250( .a(N339), .b(N650), .O(N721) );
inv1 gate251( .a(N651), .O(N722) );
and2 gate252( .a(N654), .b(N651), .O(N727) );
nor2 gate253( .a(N341), .b(N659), .O(N731) );

  xor2  gate874(.a(N261), .b(N654), .O(gate254inter0));
  nand2 gate875(.a(gate254inter0), .b(s_70), .O(gate254inter1));
  and2  gate876(.a(N261), .b(N654), .O(gate254inter2));
  inv1  gate877(.a(s_70), .O(gate254inter3));
  inv1  gate878(.a(s_71), .O(gate254inter4));
  nand2 gate879(.a(gate254inter4), .b(gate254inter3), .O(gate254inter5));
  nor2  gate880(.a(gate254inter5), .b(gate254inter2), .O(gate254inter6));
  inv1  gate881(.a(N654), .O(gate254inter7));
  inv1  gate882(.a(N261), .O(gate254inter8));
  nand2 gate883(.a(gate254inter8), .b(gate254inter7), .O(gate254inter9));
  nand2 gate884(.a(s_71), .b(gate254inter3), .O(gate254inter10));
  nor2  gate885(.a(gate254inter10), .b(gate254inter9), .O(gate254inter11));
  nor2  gate886(.a(gate254inter11), .b(gate254inter6), .O(gate254inter12));
  nand2 gate887(.a(gate254inter12), .b(gate254inter1), .O(N732));
nand3 gate255( .a(N644), .b(N654), .c(N261), .O(N733) );
nand4 gate256( .a(N635), .b(N644), .c(N654), .d(N261), .O(N734) );
inv1 gate257( .a(N662), .O(N735) );
and2 gate258( .a(N228), .b(N665), .O(N736) );
and2 gate259( .a(N237), .b(N662), .O(N737) );
inv1 gate260( .a(N670), .O(N738) );
and2 gate261( .a(N228), .b(N673), .O(N739) );
and2 gate262( .a(N237), .b(N670), .O(N740) );
inv1 gate263( .a(N678), .O(N741) );
and2 gate264( .a(N228), .b(N682), .O(N742) );
and2 gate265( .a(N237), .b(N678), .O(N743) );
inv1 gate266( .a(N687), .O(N744) );
and2 gate267( .a(N228), .b(N692), .O(N745) );
and2 gate268( .a(N237), .b(N687), .O(N746) );
inv1 gate269( .a(N697), .O(N747) );
and2 gate270( .a(N228), .b(N700), .O(N748) );
and2 gate271( .a(N237), .b(N697), .O(N749) );
inv1 gate272( .a(N705), .O(N750) );
and2 gate273( .a(N228), .b(N708), .O(N751) );
and2 gate274( .a(N237), .b(N705), .O(N752) );
inv1 gate275( .a(N713), .O(N753) );
and2 gate276( .a(N228), .b(N717), .O(N754) );
and2 gate277( .a(N237), .b(N713), .O(N755) );
inv1 gate278( .a(N722), .O(N756) );
nor2 gate279( .a(N727), .b(N261), .O(N757) );
and2 gate280( .a(N727), .b(N261), .O(N758) );
and2 gate281( .a(N228), .b(N727), .O(N759) );
and2 gate282( .a(N237), .b(N722), .O(N760) );
nand2 gate283( .a(N644), .b(N722), .O(N761) );
nand2 gate284( .a(N635), .b(N713), .O(N762) );
nand3 gate285( .a(N635), .b(N644), .c(N722), .O(N763) );
nand2 gate286( .a(N609), .b(N687), .O(N764) );
nand2 gate287( .a(N600), .b(N678), .O(N765) );
nand3 gate288( .a(N600), .b(N609), .c(N687), .O(N766) );
buf1 gate289( .a(N660), .O(N767) );
buf1 gate290( .a(N661), .O(N768) );
nor2 gate291( .a(N736), .b(N737), .O(N769) );
nor2 gate292( .a(N739), .b(N740), .O(N770) );

  xor2  gate706(.a(N743), .b(N742), .O(gate293inter0));
  nand2 gate707(.a(gate293inter0), .b(s_46), .O(gate293inter1));
  and2  gate708(.a(N743), .b(N742), .O(gate293inter2));
  inv1  gate709(.a(s_46), .O(gate293inter3));
  inv1  gate710(.a(s_47), .O(gate293inter4));
  nand2 gate711(.a(gate293inter4), .b(gate293inter3), .O(gate293inter5));
  nor2  gate712(.a(gate293inter5), .b(gate293inter2), .O(gate293inter6));
  inv1  gate713(.a(N742), .O(gate293inter7));
  inv1  gate714(.a(N743), .O(gate293inter8));
  nand2 gate715(.a(gate293inter8), .b(gate293inter7), .O(gate293inter9));
  nand2 gate716(.a(s_47), .b(gate293inter3), .O(gate293inter10));
  nor2  gate717(.a(gate293inter10), .b(gate293inter9), .O(gate293inter11));
  nor2  gate718(.a(gate293inter11), .b(gate293inter6), .O(gate293inter12));
  nand2 gate719(.a(gate293inter12), .b(gate293inter1), .O(N771));
nor2 gate294( .a(N745), .b(N746), .O(N772) );
nand4 gate295( .a(N750), .b(N762), .c(N763), .d(N734), .O(N773) );
nor2 gate296( .a(N748), .b(N749), .O(N777) );
nand3 gate297( .a(N753), .b(N761), .c(N733), .O(N778) );
nor2 gate298( .a(N751), .b(N752), .O(N781) );

  xor2  gate552(.a(N732), .b(N756), .O(gate299inter0));
  nand2 gate553(.a(gate299inter0), .b(s_24), .O(gate299inter1));
  and2  gate554(.a(N732), .b(N756), .O(gate299inter2));
  inv1  gate555(.a(s_24), .O(gate299inter3));
  inv1  gate556(.a(s_25), .O(gate299inter4));
  nand2 gate557(.a(gate299inter4), .b(gate299inter3), .O(gate299inter5));
  nor2  gate558(.a(gate299inter5), .b(gate299inter2), .O(gate299inter6));
  inv1  gate559(.a(N756), .O(gate299inter7));
  inv1  gate560(.a(N732), .O(gate299inter8));
  nand2 gate561(.a(gate299inter8), .b(gate299inter7), .O(gate299inter9));
  nand2 gate562(.a(s_25), .b(gate299inter3), .O(gate299inter10));
  nor2  gate563(.a(gate299inter10), .b(gate299inter9), .O(gate299inter11));
  nor2  gate564(.a(gate299inter11), .b(gate299inter6), .O(gate299inter12));
  nand2 gate565(.a(gate299inter12), .b(gate299inter1), .O(N782));
nor2 gate300( .a(N754), .b(N755), .O(N785) );
nor2 gate301( .a(N757), .b(N758), .O(N786) );
nor2 gate302( .a(N759), .b(N760), .O(N787) );
nor2 gate303( .a(N700), .b(N773), .O(N788) );
and2 gate304( .a(N700), .b(N773), .O(N789) );
nor2 gate305( .a(N708), .b(N778), .O(N790) );
and2 gate306( .a(N708), .b(N778), .O(N791) );
nor2 gate307( .a(N717), .b(N782), .O(N792) );
and2 gate308( .a(N717), .b(N782), .O(N793) );
and2 gate309( .a(N219), .b(N786), .O(N794) );

  xor2  gate860(.a(N773), .b(N628), .O(gate310inter0));
  nand2 gate861(.a(gate310inter0), .b(s_68), .O(gate310inter1));
  and2  gate862(.a(N773), .b(N628), .O(gate310inter2));
  inv1  gate863(.a(s_68), .O(gate310inter3));
  inv1  gate864(.a(s_69), .O(gate310inter4));
  nand2 gate865(.a(gate310inter4), .b(gate310inter3), .O(gate310inter5));
  nor2  gate866(.a(gate310inter5), .b(gate310inter2), .O(gate310inter6));
  inv1  gate867(.a(N628), .O(gate310inter7));
  inv1  gate868(.a(N773), .O(gate310inter8));
  nand2 gate869(.a(gate310inter8), .b(gate310inter7), .O(gate310inter9));
  nand2 gate870(.a(s_69), .b(gate310inter3), .O(gate310inter10));
  nor2  gate871(.a(gate310inter10), .b(gate310inter9), .O(gate310inter11));
  nor2  gate872(.a(gate310inter11), .b(gate310inter6), .O(gate310inter12));
  nand2 gate873(.a(gate310inter12), .b(gate310inter1), .O(N795));
nand2 gate311( .a(N795), .b(N747), .O(N796) );

  xor2  gate496(.a(N789), .b(N788), .O(gate312inter0));
  nand2 gate497(.a(gate312inter0), .b(s_16), .O(gate312inter1));
  and2  gate498(.a(N789), .b(N788), .O(gate312inter2));
  inv1  gate499(.a(s_16), .O(gate312inter3));
  inv1  gate500(.a(s_17), .O(gate312inter4));
  nand2 gate501(.a(gate312inter4), .b(gate312inter3), .O(gate312inter5));
  nor2  gate502(.a(gate312inter5), .b(gate312inter2), .O(gate312inter6));
  inv1  gate503(.a(N788), .O(gate312inter7));
  inv1  gate504(.a(N789), .O(gate312inter8));
  nand2 gate505(.a(gate312inter8), .b(gate312inter7), .O(gate312inter9));
  nand2 gate506(.a(s_17), .b(gate312inter3), .O(gate312inter10));
  nor2  gate507(.a(gate312inter10), .b(gate312inter9), .O(gate312inter11));
  nor2  gate508(.a(gate312inter11), .b(gate312inter6), .O(gate312inter12));
  nand2 gate509(.a(gate312inter12), .b(gate312inter1), .O(N802));

  xor2  gate538(.a(N791), .b(N790), .O(gate313inter0));
  nand2 gate539(.a(gate313inter0), .b(s_22), .O(gate313inter1));
  and2  gate540(.a(N791), .b(N790), .O(gate313inter2));
  inv1  gate541(.a(s_22), .O(gate313inter3));
  inv1  gate542(.a(s_23), .O(gate313inter4));
  nand2 gate543(.a(gate313inter4), .b(gate313inter3), .O(gate313inter5));
  nor2  gate544(.a(gate313inter5), .b(gate313inter2), .O(gate313inter6));
  inv1  gate545(.a(N790), .O(gate313inter7));
  inv1  gate546(.a(N791), .O(gate313inter8));
  nand2 gate547(.a(gate313inter8), .b(gate313inter7), .O(gate313inter9));
  nand2 gate548(.a(s_23), .b(gate313inter3), .O(gate313inter10));
  nor2  gate549(.a(gate313inter10), .b(gate313inter9), .O(gate313inter11));
  nor2  gate550(.a(gate313inter11), .b(gate313inter6), .O(gate313inter12));
  nand2 gate551(.a(gate313inter12), .b(gate313inter1), .O(N803));
nor2 gate314( .a(N792), .b(N793), .O(N804) );
nor2 gate315( .a(N340), .b(N794), .O(N805) );
nor2 gate316( .a(N692), .b(N796), .O(N806) );
and2 gate317( .a(N692), .b(N796), .O(N807) );
and2 gate318( .a(N219), .b(N802), .O(N808) );
and2 gate319( .a(N219), .b(N803), .O(N809) );
and2 gate320( .a(N219), .b(N804), .O(N810) );
nand4 gate321( .a(N805), .b(N787), .c(N731), .d(N529), .O(N811) );
nand2 gate322( .a(N619), .b(N796), .O(N812) );
nand3 gate323( .a(N609), .b(N619), .c(N796), .O(N813) );
nand4 gate324( .a(N600), .b(N609), .c(N619), .d(N796), .O(N814) );
nand4 gate325( .a(N738), .b(N765), .c(N766), .d(N814), .O(N815) );
nand3 gate326( .a(N741), .b(N764), .c(N813), .O(N819) );
nand2 gate327( .a(N744), .b(N812), .O(N822) );
nor2 gate328( .a(N806), .b(N807), .O(N825) );
nor2 gate329( .a(N335), .b(N808), .O(N826) );
nor2 gate330( .a(N336), .b(N809), .O(N827) );
nor2 gate331( .a(N338), .b(N810), .O(N828) );
inv1 gate332( .a(N811), .O(N829) );
nor2 gate333( .a(N665), .b(N815), .O(N830) );
and2 gate334( .a(N665), .b(N815), .O(N831) );

  xor2  gate384(.a(N819), .b(N673), .O(gate335inter0));
  nand2 gate385(.a(gate335inter0), .b(s_0), .O(gate335inter1));
  and2  gate386(.a(N819), .b(N673), .O(gate335inter2));
  inv1  gate387(.a(s_0), .O(gate335inter3));
  inv1  gate388(.a(s_1), .O(gate335inter4));
  nand2 gate389(.a(gate335inter4), .b(gate335inter3), .O(gate335inter5));
  nor2  gate390(.a(gate335inter5), .b(gate335inter2), .O(gate335inter6));
  inv1  gate391(.a(N673), .O(gate335inter7));
  inv1  gate392(.a(N819), .O(gate335inter8));
  nand2 gate393(.a(gate335inter8), .b(gate335inter7), .O(gate335inter9));
  nand2 gate394(.a(s_1), .b(gate335inter3), .O(gate335inter10));
  nor2  gate395(.a(gate335inter10), .b(gate335inter9), .O(gate335inter11));
  nor2  gate396(.a(gate335inter11), .b(gate335inter6), .O(gate335inter12));
  nand2 gate397(.a(gate335inter12), .b(gate335inter1), .O(N832));
and2 gate336( .a(N673), .b(N819), .O(N833) );

  xor2  gate720(.a(N822), .b(N682), .O(gate337inter0));
  nand2 gate721(.a(gate337inter0), .b(s_48), .O(gate337inter1));
  and2  gate722(.a(N822), .b(N682), .O(gate337inter2));
  inv1  gate723(.a(s_48), .O(gate337inter3));
  inv1  gate724(.a(s_49), .O(gate337inter4));
  nand2 gate725(.a(gate337inter4), .b(gate337inter3), .O(gate337inter5));
  nor2  gate726(.a(gate337inter5), .b(gate337inter2), .O(gate337inter6));
  inv1  gate727(.a(N682), .O(gate337inter7));
  inv1  gate728(.a(N822), .O(gate337inter8));
  nand2 gate729(.a(gate337inter8), .b(gate337inter7), .O(gate337inter9));
  nand2 gate730(.a(s_49), .b(gate337inter3), .O(gate337inter10));
  nor2  gate731(.a(gate337inter10), .b(gate337inter9), .O(gate337inter11));
  nor2  gate732(.a(gate337inter11), .b(gate337inter6), .O(gate337inter12));
  nand2 gate733(.a(gate337inter12), .b(gate337inter1), .O(N834));
and2 gate338( .a(N682), .b(N822), .O(N835) );
and2 gate339( .a(N219), .b(N825), .O(N836) );
nand3 gate340( .a(N826), .b(N777), .c(N704), .O(N837) );
nand4 gate341( .a(N827), .b(N781), .c(N712), .d(N527), .O(N838) );
nand4 gate342( .a(N828), .b(N785), .c(N721), .d(N528), .O(N839) );
inv1 gate343( .a(N829), .O(N840) );
nand2 gate344( .a(N815), .b(N593), .O(N841) );
nor2 gate345( .a(N830), .b(N831), .O(N842) );

  xor2  gate398(.a(N833), .b(N832), .O(gate346inter0));
  nand2 gate399(.a(gate346inter0), .b(s_2), .O(gate346inter1));
  and2  gate400(.a(N833), .b(N832), .O(gate346inter2));
  inv1  gate401(.a(s_2), .O(gate346inter3));
  inv1  gate402(.a(s_3), .O(gate346inter4));
  nand2 gate403(.a(gate346inter4), .b(gate346inter3), .O(gate346inter5));
  nor2  gate404(.a(gate346inter5), .b(gate346inter2), .O(gate346inter6));
  inv1  gate405(.a(N832), .O(gate346inter7));
  inv1  gate406(.a(N833), .O(gate346inter8));
  nand2 gate407(.a(gate346inter8), .b(gate346inter7), .O(gate346inter9));
  nand2 gate408(.a(s_3), .b(gate346inter3), .O(gate346inter10));
  nor2  gate409(.a(gate346inter10), .b(gate346inter9), .O(gate346inter11));
  nor2  gate410(.a(gate346inter11), .b(gate346inter6), .O(gate346inter12));
  nand2 gate411(.a(gate346inter12), .b(gate346inter1), .O(N843));

  xor2  gate468(.a(N835), .b(N834), .O(gate347inter0));
  nand2 gate469(.a(gate347inter0), .b(s_12), .O(gate347inter1));
  and2  gate470(.a(N835), .b(N834), .O(gate347inter2));
  inv1  gate471(.a(s_12), .O(gate347inter3));
  inv1  gate472(.a(s_13), .O(gate347inter4));
  nand2 gate473(.a(gate347inter4), .b(gate347inter3), .O(gate347inter5));
  nor2  gate474(.a(gate347inter5), .b(gate347inter2), .O(gate347inter6));
  inv1  gate475(.a(N834), .O(gate347inter7));
  inv1  gate476(.a(N835), .O(gate347inter8));
  nand2 gate477(.a(gate347inter8), .b(gate347inter7), .O(gate347inter9));
  nand2 gate478(.a(s_13), .b(gate347inter3), .O(gate347inter10));
  nor2  gate479(.a(gate347inter10), .b(gate347inter9), .O(gate347inter11));
  nor2  gate480(.a(gate347inter11), .b(gate347inter6), .O(gate347inter12));
  nand2 gate481(.a(gate347inter12), .b(gate347inter1), .O(N844));
nor2 gate348( .a(N334), .b(N836), .O(N845) );
inv1 gate349( .a(N837), .O(N846) );
inv1 gate350( .a(N838), .O(N847) );
inv1 gate351( .a(N839), .O(N848) );
and2 gate352( .a(N735), .b(N841), .O(N849) );
buf1 gate353( .a(N840), .O(N850) );
and2 gate354( .a(N219), .b(N842), .O(N851) );
and2 gate355( .a(N219), .b(N843), .O(N852) );
and2 gate356( .a(N219), .b(N844), .O(N853) );
nand3 gate357( .a(N845), .b(N772), .c(N696), .O(N854) );
inv1 gate358( .a(N846), .O(N855) );
inv1 gate359( .a(N847), .O(N856) );
inv1 gate360( .a(N848), .O(N857) );
inv1 gate361( .a(N849), .O(N858) );
nor2 gate362( .a(N417), .b(N851), .O(N859) );
nor2 gate363( .a(N332), .b(N852), .O(N860) );

  xor2  gate650(.a(N853), .b(N333), .O(gate364inter0));
  nand2 gate651(.a(gate364inter0), .b(s_38), .O(gate364inter1));
  and2  gate652(.a(N853), .b(N333), .O(gate364inter2));
  inv1  gate653(.a(s_38), .O(gate364inter3));
  inv1  gate654(.a(s_39), .O(gate364inter4));
  nand2 gate655(.a(gate364inter4), .b(gate364inter3), .O(gate364inter5));
  nor2  gate656(.a(gate364inter5), .b(gate364inter2), .O(gate364inter6));
  inv1  gate657(.a(N333), .O(gate364inter7));
  inv1  gate658(.a(N853), .O(gate364inter8));
  nand2 gate659(.a(gate364inter8), .b(gate364inter7), .O(gate364inter9));
  nand2 gate660(.a(s_39), .b(gate364inter3), .O(gate364inter10));
  nor2  gate661(.a(gate364inter10), .b(gate364inter9), .O(gate364inter11));
  nor2  gate662(.a(gate364inter11), .b(gate364inter6), .O(gate364inter12));
  nand2 gate663(.a(gate364inter12), .b(gate364inter1), .O(N861));
inv1 gate365( .a(N854), .O(N862) );
buf1 gate366( .a(N855), .O(N863) );
buf1 gate367( .a(N856), .O(N864) );
buf1 gate368( .a(N857), .O(N865) );
buf1 gate369( .a(N858), .O(N866) );
nand3 gate370( .a(N859), .b(N769), .c(N669), .O(N867) );
nand3 gate371( .a(N860), .b(N770), .c(N677), .O(N868) );
nand3 gate372( .a(N861), .b(N771), .c(N686), .O(N869) );
inv1 gate373( .a(N862), .O(N870) );
inv1 gate374( .a(N867), .O(N871) );
inv1 gate375( .a(N868), .O(N872) );
inv1 gate376( .a(N869), .O(N873) );
buf1 gate377( .a(N870), .O(N874) );
inv1 gate378( .a(N871), .O(N875) );
inv1 gate379( .a(N872), .O(N876) );
inv1 gate380( .a(N873), .O(N877) );
buf1 gate381( .a(N875), .O(N878) );
buf1 gate382( .a(N876), .O(N879) );
buf1 gate383( .a(N877), .O(N880) );

endmodule