module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);

input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;//RE__PI;

input s_0,s_1;//RE__ALLOW(00,01,10,11);
input s_2,s_3;//RE__ALLOW(00,01,10,11);
input s_4,s_5;//RE__ALLOW(00,01,10,11);
input s_6,s_7;//RE__ALLOW(00,01,10,11);
input s_8,s_9;//RE__ALLOW(00,01,10,11);
input s_10,s_11;//RE__ALLOW(00,01,10,11);
input s_12,s_13;//RE__ALLOW(00,01,10,11);
input s_14,s_15;//RE__ALLOW(00,01,10,11);
input s_16,s_17;//RE__ALLOW(00,01,10,11);
input s_18,s_19;//RE__ALLOW(00,01,10,11);
input s_20,s_21;//RE__ALLOW(00,01,10,11);
input s_22,s_23;//RE__ALLOW(00,01,10,11);
input s_24,s_25;//RE__ALLOW(00,01,10,11);
input s_26,s_27;//RE__ALLOW(00,01,10,11);
input s_28,s_29;//RE__ALLOW(00,01,10,11);
input s_30,s_31;//RE__ALLOW(00,01,10,11);
input s_32,s_33;//RE__ALLOW(00,01,10,11);
input s_34,s_35;//RE__ALLOW(00,01,10,11);
input s_36,s_37;//RE__ALLOW(00,01,10,11);
input s_38,s_39;//RE__ALLOW(00,01,10,11);
input s_40,s_41;//RE__ALLOW(00,01,10,11);
input s_42,s_43;//RE__ALLOW(00,01,10,11);
input s_44,s_45;//RE__ALLOW(00,01,10,11);
input s_46,s_47;//RE__ALLOW(00,01,10,11);
input s_48,s_49;//RE__ALLOW(00,01,10,11);
input s_50,s_51;//RE__ALLOW(00,01,10,11);
input s_52,s_53;//RE__ALLOW(00,01,10,11);
input s_54,s_55;//RE__ALLOW(00,01,10,11);
input s_56,s_57;//RE__ALLOW(00,01,10,11);
input s_58,s_59;//RE__ALLOW(00,01,10,11);
input s_60,s_61;//RE__ALLOW(00,01,10,11);
input s_62,s_63;//RE__ALLOW(00,01,10,11);
input s_64,s_65;//RE__ALLOW(00,01,10,11);
input s_66,s_67;//RE__ALLOW(00,01,10,11);
input s_68,s_69;//RE__ALLOW(00,01,10,11);
input s_70,s_71;//RE__ALLOW(00,01,10,11);
input s_72,s_73;//RE__ALLOW(00,01,10,11);
input s_74,s_75;//RE__ALLOW(00,01,10,11);
input s_76,s_77;//RE__ALLOW(00,01,10,11);
input s_78,s_79;//RE__ALLOW(00,01,10,11);
input s_80,s_81;//RE__ALLOW(00,01,10,11);
input s_82,s_83;//RE__ALLOW(00,01,10,11);
input s_84,s_85;//RE__ALLOW(00,01,10,11);
input s_86,s_87;//RE__ALLOW(00,01,10,11);
input s_88,s_89;//RE__ALLOW(00,01,10,11);
input s_90,s_91;//RE__ALLOW(00,01,10,11);
input s_92,s_93;//RE__ALLOW(00,01,10,11);
input s_94,s_95;//RE__ALLOW(00,01,10,11);
input s_96,s_97;//RE__ALLOW(00,01,10,11);
input s_98,s_99;//RE__ALLOW(00,01,10,11);
input s_100,s_101;//RE__ALLOW(00,01,10,11);
input s_102,s_103;//RE__ALLOW(00,01,10,11);
input s_104,s_105;//RE__ALLOW(00,01,10,11);
input s_106,s_107;//RE__ALLOW(00,01,10,11);
input s_108,s_109;//RE__ALLOW(00,01,10,11);
input s_110,s_111;//RE__ALLOW(00,01,10,11);
input s_112,s_113;//RE__ALLOW(00,01,10,11);
input s_114,s_115;//RE__ALLOW(00,01,10,11);
input s_116,s_117;//RE__ALLOW(00,01,10,11);
input s_118,s_119;//RE__ALLOW(00,01,10,11);
input s_120,s_121;//RE__ALLOW(00,01,10,11);
input s_122,s_123;//RE__ALLOW(00,01,10,11);
input s_124,s_125;//RE__ALLOW(00,01,10,11);
input s_126,s_127;//RE__ALLOW(00,01,10,11);
input s_128,s_129;//RE__ALLOW(00,01,10,11);
input s_130,s_131;//RE__ALLOW(00,01,10,11);
input s_132,s_133;//RE__ALLOW(00,01,10,11);
input s_134,s_135;//RE__ALLOW(00,01,10,11);
input s_136,s_137;//RE__ALLOW(00,01,10,11);
input s_138,s_139;//RE__ALLOW(00,01,10,11);
input s_140,s_141;//RE__ALLOW(00,01,10,11);
input s_142,s_143;//RE__ALLOW(00,01,10,11);
input s_144,s_145;//RE__ALLOW(00,01,10,11);
input s_146,s_147;//RE__ALLOW(00,01,10,11);
input s_148,s_149;//RE__ALLOW(00,01,10,11);
input s_150,s_151;//RE__ALLOW(00,01,10,11);
input s_152,s_153;//RE__ALLOW(00,01,10,11);
input s_154,s_155;//RE__ALLOW(00,01,10,11);
input s_156,s_157;//RE__ALLOW(00,01,10,11);
input s_158,s_159;//RE__ALLOW(00,01,10,11);
input s_160,s_161;//RE__ALLOW(00,01,10,11);
input s_162,s_163;//RE__ALLOW(00,01,10,11);
input s_164,s_165;//RE__ALLOW(00,01,10,11);
input s_166,s_167;//RE__ALLOW(00,01,10,11);
input s_168,s_169;//RE__ALLOW(00,01,10,11);
input s_170,s_171;//RE__ALLOW(00,01,10,11);
input s_172,s_173;//RE__ALLOW(00,01,10,11);
input s_174,s_175;//RE__ALLOW(00,01,10,11);
input s_176,s_177;//RE__ALLOW(00,01,10,11);
input s_178,s_179;//RE__ALLOW(00,01,10,11);
input s_180,s_181;//RE__ALLOW(00,01,10,11);
input s_182,s_183;//RE__ALLOW(00,01,10,11);
input s_184,s_185;//RE__ALLOW(00,01,10,11);
input s_186,s_187;//RE__ALLOW(00,01,10,11);
input s_188,s_189;//RE__ALLOW(00,01,10,11);
input s_190,s_191;//RE__ALLOW(00,01,10,11);
input s_192,s_193;//RE__ALLOW(00,01,10,11);
input s_194,s_195;//RE__ALLOW(00,01,10,11);
input s_196,s_197;//RE__ALLOW(00,01,10,11);
input s_198,s_199;//RE__ALLOW(00,01,10,11);
input s_200,s_201;//RE__ALLOW(00,01,10,11);
input s_202,s_203;//RE__ALLOW(00,01,10,11);
input s_204,s_205;//RE__ALLOW(00,01,10,11);
input s_206,s_207;//RE__ALLOW(00,01,10,11);
input s_208,s_209;//RE__ALLOW(00,01,10,11);
input s_210,s_211;//RE__ALLOW(00,01,10,11);
input s_212,s_213;//RE__ALLOW(00,01,10,11);
input s_214,s_215;//RE__ALLOW(00,01,10,11);
input s_216,s_217;//RE__ALLOW(00,01,10,11);
input s_218,s_219;//RE__ALLOW(00,01,10,11);
input s_220,s_221;//RE__ALLOW(00,01,10,11);
input s_222,s_223;//RE__ALLOW(00,01,10,11);
input s_224,s_225;//RE__ALLOW(00,01,10,11);
input s_226,s_227;//RE__ALLOW(00,01,10,11);
input s_228,s_229;//RE__ALLOW(00,01,10,11);
input s_230,s_231;//RE__ALLOW(00,01,10,11);
input s_232,s_233;//RE__ALLOW(00,01,10,11);
input s_234,s_235;//RE__ALLOW(00,01,10,11);
input s_236,s_237;//RE__ALLOW(00,01,10,11);
input s_238,s_239;//RE__ALLOW(00,01,10,11);
input s_240,s_241;//RE__ALLOW(00,01,10,11);
input s_242,s_243;//RE__ALLOW(00,01,10,11);
input s_244,s_245;//RE__ALLOW(00,01,10,11);
input s_246,s_247;//RE__ALLOW(00,01,10,11);
input s_248,s_249;//RE__ALLOW(00,01,10,11);
input s_250,s_251;//RE__ALLOW(00,01,10,11);
input s_252,s_253;//RE__ALLOW(00,01,10,11);
input s_254,s_255;//RE__ALLOW(00,01,10,11);
input s_256,s_257;//RE__ALLOW(00,01,10,11);
input s_258,s_259;//RE__ALLOW(00,01,10,11);
input s_260,s_261;//RE__ALLOW(00,01,10,11);
input s_262,s_263;//RE__ALLOW(00,01,10,11);
input s_264,s_265;//RE__ALLOW(00,01,10,11);
input s_266,s_267;//RE__ALLOW(00,01,10,11);
input s_268,s_269;//RE__ALLOW(00,01,10,11);
input s_270,s_271;//RE__ALLOW(00,01,10,11);
input s_272,s_273;//RE__ALLOW(00,01,10,11);
input s_274,s_275;//RE__ALLOW(00,01,10,11);
input s_276,s_277;//RE__ALLOW(00,01,10,11);
input s_278,s_279;//RE__ALLOW(00,01,10,11);
input s_280,s_281;//RE__ALLOW(00,01,10,11);
input s_282,s_283;//RE__ALLOW(00,01,10,11);
input s_284,s_285;//RE__ALLOW(00,01,10,11);
input s_286,s_287;//RE__ALLOW(00,01,10,11);
input s_288,s_289;//RE__ALLOW(00,01,10,11);
input s_290,s_291;//RE__ALLOW(00,01,10,11);
input s_292,s_293;//RE__ALLOW(00,01,10,11);
input s_294,s_295;//RE__ALLOW(00,01,10,11);
input s_296,s_297;//RE__ALLOW(00,01,10,11);
input s_298,s_299;//RE__ALLOW(00,01,10,11);
input s_300,s_301;//RE__ALLOW(00,01,10,11);
input s_302,s_303;//RE__ALLOW(00,01,10,11);
input s_304,s_305;//RE__ALLOW(00,01,10,11);
input s_306,s_307;//RE__ALLOW(00,01,10,11);
input s_308,s_309;//RE__ALLOW(00,01,10,11);
input s_310,s_311;//RE__ALLOW(00,01,10,11);
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;

  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate405inter0, gate405inter1, gate405inter2, gate405inter3, gate405inter4, gate405inter5, gate405inter6, gate405inter7, gate405inter8, gate405inter9, gate405inter10, gate405inter11, gate405inter12, gate403inter0, gate403inter1, gate403inter2, gate403inter3, gate403inter4, gate403inter5, gate403inter6, gate403inter7, gate403inter8, gate403inter9, gate403inter10, gate403inter11, gate403inter12, gate439inter0, gate439inter1, gate439inter2, gate439inter3, gate439inter4, gate439inter5, gate439inter6, gate439inter7, gate439inter8, gate439inter9, gate439inter10, gate439inter11, gate439inter12, gate270inter0, gate270inter1, gate270inter2, gate270inter3, gate270inter4, gate270inter5, gate270inter6, gate270inter7, gate270inter8, gate270inter9, gate270inter10, gate270inter11, gate270inter12, gate59inter0, gate59inter1, gate59inter2, gate59inter3, gate59inter4, gate59inter5, gate59inter6, gate59inter7, gate59inter8, gate59inter9, gate59inter10, gate59inter11, gate59inter12, gate13inter0, gate13inter1, gate13inter2, gate13inter3, gate13inter4, gate13inter5, gate13inter6, gate13inter7, gate13inter8, gate13inter9, gate13inter10, gate13inter11, gate13inter12, gate490inter0, gate490inter1, gate490inter2, gate490inter3, gate490inter4, gate490inter5, gate490inter6, gate490inter7, gate490inter8, gate490inter9, gate490inter10, gate490inter11, gate490inter12, gate157inter0, gate157inter1, gate157inter2, gate157inter3, gate157inter4, gate157inter5, gate157inter6, gate157inter7, gate157inter8, gate157inter9, gate157inter10, gate157inter11, gate157inter12, gate263inter0, gate263inter1, gate263inter2, gate263inter3, gate263inter4, gate263inter5, gate263inter6, gate263inter7, gate263inter8, gate263inter9, gate263inter10, gate263inter11, gate263inter12, gate22inter0, gate22inter1, gate22inter2, gate22inter3, gate22inter4, gate22inter5, gate22inter6, gate22inter7, gate22inter8, gate22inter9, gate22inter10, gate22inter11, gate22inter12, gate65inter0, gate65inter1, gate65inter2, gate65inter3, gate65inter4, gate65inter5, gate65inter6, gate65inter7, gate65inter8, gate65inter9, gate65inter10, gate65inter11, gate65inter12, gate119inter0, gate119inter1, gate119inter2, gate119inter3, gate119inter4, gate119inter5, gate119inter6, gate119inter7, gate119inter8, gate119inter9, gate119inter10, gate119inter11, gate119inter12, gate52inter0, gate52inter1, gate52inter2, gate52inter3, gate52inter4, gate52inter5, gate52inter6, gate52inter7, gate52inter8, gate52inter9, gate52inter10, gate52inter11, gate52inter12, gate253inter0, gate253inter1, gate253inter2, gate253inter3, gate253inter4, gate253inter5, gate253inter6, gate253inter7, gate253inter8, gate253inter9, gate253inter10, gate253inter11, gate253inter12, gate396inter0, gate396inter1, gate396inter2, gate396inter3, gate396inter4, gate396inter5, gate396inter6, gate396inter7, gate396inter8, gate396inter9, gate396inter10, gate396inter11, gate396inter12, gate41inter0, gate41inter1, gate41inter2, gate41inter3, gate41inter4, gate41inter5, gate41inter6, gate41inter7, gate41inter8, gate41inter9, gate41inter10, gate41inter11, gate41inter12, gate282inter0, gate282inter1, gate282inter2, gate282inter3, gate282inter4, gate282inter5, gate282inter6, gate282inter7, gate282inter8, gate282inter9, gate282inter10, gate282inter11, gate282inter12, gate444inter0, gate444inter1, gate444inter2, gate444inter3, gate444inter4, gate444inter5, gate444inter6, gate444inter7, gate444inter8, gate444inter9, gate444inter10, gate444inter11, gate444inter12, gate25inter0, gate25inter1, gate25inter2, gate25inter3, gate25inter4, gate25inter5, gate25inter6, gate25inter7, gate25inter8, gate25inter9, gate25inter10, gate25inter11, gate25inter12, gate438inter0, gate438inter1, gate438inter2, gate438inter3, gate438inter4, gate438inter5, gate438inter6, gate438inter7, gate438inter8, gate438inter9, gate438inter10, gate438inter11, gate438inter12, gate295inter0, gate295inter1, gate295inter2, gate295inter3, gate295inter4, gate295inter5, gate295inter6, gate295inter7, gate295inter8, gate295inter9, gate295inter10, gate295inter11, gate295inter12, gate461inter0, gate461inter1, gate461inter2, gate461inter3, gate461inter4, gate461inter5, gate461inter6, gate461inter7, gate461inter8, gate461inter9, gate461inter10, gate461inter11, gate461inter12, gate274inter0, gate274inter1, gate274inter2, gate274inter3, gate274inter4, gate274inter5, gate274inter6, gate274inter7, gate274inter8, gate274inter9, gate274inter10, gate274inter11, gate274inter12, gate26inter0, gate26inter1, gate26inter2, gate26inter3, gate26inter4, gate26inter5, gate26inter6, gate26inter7, gate26inter8, gate26inter9, gate26inter10, gate26inter11, gate26inter12, gate85inter0, gate85inter1, gate85inter2, gate85inter3, gate85inter4, gate85inter5, gate85inter6, gate85inter7, gate85inter8, gate85inter9, gate85inter10, gate85inter11, gate85inter12, gate195inter0, gate195inter1, gate195inter2, gate195inter3, gate195inter4, gate195inter5, gate195inter6, gate195inter7, gate195inter8, gate195inter9, gate195inter10, gate195inter11, gate195inter12, gate249inter0, gate249inter1, gate249inter2, gate249inter3, gate249inter4, gate249inter5, gate249inter6, gate249inter7, gate249inter8, gate249inter9, gate249inter10, gate249inter11, gate249inter12, gate163inter0, gate163inter1, gate163inter2, gate163inter3, gate163inter4, gate163inter5, gate163inter6, gate163inter7, gate163inter8, gate163inter9, gate163inter10, gate163inter11, gate163inter12, gate109inter0, gate109inter1, gate109inter2, gate109inter3, gate109inter4, gate109inter5, gate109inter6, gate109inter7, gate109inter8, gate109inter9, gate109inter10, gate109inter11, gate109inter12, gate426inter0, gate426inter1, gate426inter2, gate426inter3, gate426inter4, gate426inter5, gate426inter6, gate426inter7, gate426inter8, gate426inter9, gate426inter10, gate426inter11, gate426inter12, gate55inter0, gate55inter1, gate55inter2, gate55inter3, gate55inter4, gate55inter5, gate55inter6, gate55inter7, gate55inter8, gate55inter9, gate55inter10, gate55inter11, gate55inter12, gate201inter0, gate201inter1, gate201inter2, gate201inter3, gate201inter4, gate201inter5, gate201inter6, gate201inter7, gate201inter8, gate201inter9, gate201inter10, gate201inter11, gate201inter12, gate144inter0, gate144inter1, gate144inter2, gate144inter3, gate144inter4, gate144inter5, gate144inter6, gate144inter7, gate144inter8, gate144inter9, gate144inter10, gate144inter11, gate144inter12, gate472inter0, gate472inter1, gate472inter2, gate472inter3, gate472inter4, gate472inter5, gate472inter6, gate472inter7, gate472inter8, gate472inter9, gate472inter10, gate472inter11, gate472inter12, gate88inter0, gate88inter1, gate88inter2, gate88inter3, gate88inter4, gate88inter5, gate88inter6, gate88inter7, gate88inter8, gate88inter9, gate88inter10, gate88inter11, gate88inter12, gate468inter0, gate468inter1, gate468inter2, gate468inter3, gate468inter4, gate468inter5, gate468inter6, gate468inter7, gate468inter8, gate468inter9, gate468inter10, gate468inter11, gate468inter12, gate235inter0, gate235inter1, gate235inter2, gate235inter3, gate235inter4, gate235inter5, gate235inter6, gate235inter7, gate235inter8, gate235inter9, gate235inter10, gate235inter11, gate235inter12, gate430inter0, gate430inter1, gate430inter2, gate430inter3, gate430inter4, gate430inter5, gate430inter6, gate430inter7, gate430inter8, gate430inter9, gate430inter10, gate430inter11, gate430inter12, gate167inter0, gate167inter1, gate167inter2, gate167inter3, gate167inter4, gate167inter5, gate167inter6, gate167inter7, gate167inter8, gate167inter9, gate167inter10, gate167inter11, gate167inter12, gate57inter0, gate57inter1, gate57inter2, gate57inter3, gate57inter4, gate57inter5, gate57inter6, gate57inter7, gate57inter8, gate57inter9, gate57inter10, gate57inter11, gate57inter12, gate82inter0, gate82inter1, gate82inter2, gate82inter3, gate82inter4, gate82inter5, gate82inter6, gate82inter7, gate82inter8, gate82inter9, gate82inter10, gate82inter11, gate82inter12, gate36inter0, gate36inter1, gate36inter2, gate36inter3, gate36inter4, gate36inter5, gate36inter6, gate36inter7, gate36inter8, gate36inter9, gate36inter10, gate36inter11, gate36inter12, gate402inter0, gate402inter1, gate402inter2, gate402inter3, gate402inter4, gate402inter5, gate402inter6, gate402inter7, gate402inter8, gate402inter9, gate402inter10, gate402inter11, gate402inter12, gate69inter0, gate69inter1, gate69inter2, gate69inter3, gate69inter4, gate69inter5, gate69inter6, gate69inter7, gate69inter8, gate69inter9, gate69inter10, gate69inter11, gate69inter12, gate268inter0, gate268inter1, gate268inter2, gate268inter3, gate268inter4, gate268inter5, gate268inter6, gate268inter7, gate268inter8, gate268inter9, gate268inter10, gate268inter11, gate268inter12, gate392inter0, gate392inter1, gate392inter2, gate392inter3, gate392inter4, gate392inter5, gate392inter6, gate392inter7, gate392inter8, gate392inter9, gate392inter10, gate392inter11, gate392inter12, gate454inter0, gate454inter1, gate454inter2, gate454inter3, gate454inter4, gate454inter5, gate454inter6, gate454inter7, gate454inter8, gate454inter9, gate454inter10, gate454inter11, gate454inter12, gate100inter0, gate100inter1, gate100inter2, gate100inter3, gate100inter4, gate100inter5, gate100inter6, gate100inter7, gate100inter8, gate100inter9, gate100inter10, gate100inter11, gate100inter12, gate64inter0, gate64inter1, gate64inter2, gate64inter3, gate64inter4, gate64inter5, gate64inter6, gate64inter7, gate64inter8, gate64inter9, gate64inter10, gate64inter11, gate64inter12, gate228inter0, gate228inter1, gate228inter2, gate228inter3, gate228inter4, gate228inter5, gate228inter6, gate228inter7, gate228inter8, gate228inter9, gate228inter10, gate228inter11, gate228inter12, gate31inter0, gate31inter1, gate31inter2, gate31inter3, gate31inter4, gate31inter5, gate31inter6, gate31inter7, gate31inter8, gate31inter9, gate31inter10, gate31inter11, gate31inter12, gate111inter0, gate111inter1, gate111inter2, gate111inter3, gate111inter4, gate111inter5, gate111inter6, gate111inter7, gate111inter8, gate111inter9, gate111inter10, gate111inter11, gate111inter12, gate418inter0, gate418inter1, gate418inter2, gate418inter3, gate418inter4, gate418inter5, gate418inter6, gate418inter7, gate418inter8, gate418inter9, gate418inter10, gate418inter11, gate418inter12, gate204inter0, gate204inter1, gate204inter2, gate204inter3, gate204inter4, gate204inter5, gate204inter6, gate204inter7, gate204inter8, gate204inter9, gate204inter10, gate204inter11, gate204inter12, gate446inter0, gate446inter1, gate446inter2, gate446inter3, gate446inter4, gate446inter5, gate446inter6, gate446inter7, gate446inter8, gate446inter9, gate446inter10, gate446inter11, gate446inter12, gate47inter0, gate47inter1, gate47inter2, gate47inter3, gate47inter4, gate47inter5, gate47inter6, gate47inter7, gate47inter8, gate47inter9, gate47inter10, gate47inter11, gate47inter12, gate96inter0, gate96inter1, gate96inter2, gate96inter3, gate96inter4, gate96inter5, gate96inter6, gate96inter7, gate96inter8, gate96inter9, gate96inter10, gate96inter11, gate96inter12, gate512inter0, gate512inter1, gate512inter2, gate512inter3, gate512inter4, gate512inter5, gate512inter6, gate512inter7, gate512inter8, gate512inter9, gate512inter10, gate512inter11, gate512inter12, gate178inter0, gate178inter1, gate178inter2, gate178inter3, gate178inter4, gate178inter5, gate178inter6, gate178inter7, gate178inter8, gate178inter9, gate178inter10, gate178inter11, gate178inter12, gate488inter0, gate488inter1, gate488inter2, gate488inter3, gate488inter4, gate488inter5, gate488inter6, gate488inter7, gate488inter8, gate488inter9, gate488inter10, gate488inter11, gate488inter12, gate129inter0, gate129inter1, gate129inter2, gate129inter3, gate129inter4, gate129inter5, gate129inter6, gate129inter7, gate129inter8, gate129inter9, gate129inter10, gate129inter11, gate129inter12, gate89inter0, gate89inter1, gate89inter2, gate89inter3, gate89inter4, gate89inter5, gate89inter6, gate89inter7, gate89inter8, gate89inter9, gate89inter10, gate89inter11, gate89inter12, gate480inter0, gate480inter1, gate480inter2, gate480inter3, gate480inter4, gate480inter5, gate480inter6, gate480inter7, gate480inter8, gate480inter9, gate480inter10, gate480inter11, gate480inter12, gate237inter0, gate237inter1, gate237inter2, gate237inter3, gate237inter4, gate237inter5, gate237inter6, gate237inter7, gate237inter8, gate237inter9, gate237inter10, gate237inter11, gate237inter12, gate264inter0, gate264inter1, gate264inter2, gate264inter3, gate264inter4, gate264inter5, gate264inter6, gate264inter7, gate264inter8, gate264inter9, gate264inter10, gate264inter11, gate264inter12, gate259inter0, gate259inter1, gate259inter2, gate259inter3, gate259inter4, gate259inter5, gate259inter6, gate259inter7, gate259inter8, gate259inter9, gate259inter10, gate259inter11, gate259inter12, gate72inter0, gate72inter1, gate72inter2, gate72inter3, gate72inter4, gate72inter5, gate72inter6, gate72inter7, gate72inter8, gate72inter9, gate72inter10, gate72inter11, gate72inter12, gate81inter0, gate81inter1, gate81inter2, gate81inter3, gate81inter4, gate81inter5, gate81inter6, gate81inter7, gate81inter8, gate81inter9, gate81inter10, gate81inter11, gate81inter12, gate208inter0, gate208inter1, gate208inter2, gate208inter3, gate208inter4, gate208inter5, gate208inter6, gate208inter7, gate208inter8, gate208inter9, gate208inter10, gate208inter11, gate208inter12, gate165inter0, gate165inter1, gate165inter2, gate165inter3, gate165inter4, gate165inter5, gate165inter6, gate165inter7, gate165inter8, gate165inter9, gate165inter10, gate165inter11, gate165inter12, gate113inter0, gate113inter1, gate113inter2, gate113inter3, gate113inter4, gate113inter5, gate113inter6, gate113inter7, gate113inter8, gate113inter9, gate113inter10, gate113inter11, gate113inter12, gate469inter0, gate469inter1, gate469inter2, gate469inter3, gate469inter4, gate469inter5, gate469inter6, gate469inter7, gate469inter8, gate469inter9, gate469inter10, gate469inter11, gate469inter12, gate283inter0, gate283inter1, gate283inter2, gate283inter3, gate283inter4, gate283inter5, gate283inter6, gate283inter7, gate283inter8, gate283inter9, gate283inter10, gate283inter11, gate283inter12, gate441inter0, gate441inter1, gate441inter2, gate441inter3, gate441inter4, gate441inter5, gate441inter6, gate441inter7, gate441inter8, gate441inter9, gate441inter10, gate441inter11, gate441inter12, gate118inter0, gate118inter1, gate118inter2, gate118inter3, gate118inter4, gate118inter5, gate118inter6, gate118inter7, gate118inter8, gate118inter9, gate118inter10, gate118inter11, gate118inter12, gate388inter0, gate388inter1, gate388inter2, gate388inter3, gate388inter4, gate388inter5, gate388inter6, gate388inter7, gate388inter8, gate388inter9, gate388inter10, gate388inter11, gate388inter12, gate436inter0, gate436inter1, gate436inter2, gate436inter3, gate436inter4, gate436inter5, gate436inter6, gate436inter7, gate436inter8, gate436inter9, gate436inter10, gate436inter11, gate436inter12, gate507inter0, gate507inter1, gate507inter2, gate507inter3, gate507inter4, gate507inter5, gate507inter6, gate507inter7, gate507inter8, gate507inter9, gate507inter10, gate507inter11, gate507inter12, gate255inter0, gate255inter1, gate255inter2, gate255inter3, gate255inter4, gate255inter5, gate255inter6, gate255inter7, gate255inter8, gate255inter9, gate255inter10, gate255inter11, gate255inter12, gate261inter0, gate261inter1, gate261inter2, gate261inter3, gate261inter4, gate261inter5, gate261inter6, gate261inter7, gate261inter8, gate261inter9, gate261inter10, gate261inter11, gate261inter12, gate500inter0, gate500inter1, gate500inter2, gate500inter3, gate500inter4, gate500inter5, gate500inter6, gate500inter7, gate500inter8, gate500inter9, gate500inter10, gate500inter11, gate500inter12, gate38inter0, gate38inter1, gate38inter2, gate38inter3, gate38inter4, gate38inter5, gate38inter6, gate38inter7, gate38inter8, gate38inter9, gate38inter10, gate38inter11, gate38inter12, gate275inter0, gate275inter1, gate275inter2, gate275inter3, gate275inter4, gate275inter5, gate275inter6, gate275inter7, gate275inter8, gate275inter9, gate275inter10, gate275inter11, gate275inter12, gate258inter0, gate258inter1, gate258inter2, gate258inter3, gate258inter4, gate258inter5, gate258inter6, gate258inter7, gate258inter8, gate258inter9, gate258inter10, gate258inter11, gate258inter12, gate481inter0, gate481inter1, gate481inter2, gate481inter3, gate481inter4, gate481inter5, gate481inter6, gate481inter7, gate481inter8, gate481inter9, gate481inter10, gate481inter11, gate481inter12, gate254inter0, gate254inter1, gate254inter2, gate254inter3, gate254inter4, gate254inter5, gate254inter6, gate254inter7, gate254inter8, gate254inter9, gate254inter10, gate254inter11, gate254inter12, gate460inter0, gate460inter1, gate460inter2, gate460inter3, gate460inter4, gate460inter5, gate460inter6, gate460inter7, gate460inter8, gate460inter9, gate460inter10, gate460inter11, gate460inter12, gate28inter0, gate28inter1, gate28inter2, gate28inter3, gate28inter4, gate28inter5, gate28inter6, gate28inter7, gate28inter8, gate28inter9, gate28inter10, gate28inter11, gate28inter12, gate143inter0, gate143inter1, gate143inter2, gate143inter3, gate143inter4, gate143inter5, gate143inter6, gate143inter7, gate143inter8, gate143inter9, gate143inter10, gate143inter11, gate143inter12, gate410inter0, gate410inter1, gate410inter2, gate410inter3, gate410inter4, gate410inter5, gate410inter6, gate410inter7, gate410inter8, gate410inter9, gate410inter10, gate410inter11, gate410inter12, gate287inter0, gate287inter1, gate287inter2, gate287inter3, gate287inter4, gate287inter5, gate287inter6, gate287inter7, gate287inter8, gate287inter9, gate287inter10, gate287inter11, gate287inter12, gate93inter0, gate93inter1, gate93inter2, gate93inter3, gate93inter4, gate93inter5, gate93inter6, gate93inter7, gate93inter8, gate93inter9, gate93inter10, gate93inter11, gate93inter12, gate149inter0, gate149inter1, gate149inter2, gate149inter3, gate149inter4, gate149inter5, gate149inter6, gate149inter7, gate149inter8, gate149inter9, gate149inter10, gate149inter11, gate149inter12, gate98inter0, gate98inter1, gate98inter2, gate98inter3, gate98inter4, gate98inter5, gate98inter6, gate98inter7, gate98inter8, gate98inter9, gate98inter10, gate98inter11, gate98inter12, gate16inter0, gate16inter1, gate16inter2, gate16inter3, gate16inter4, gate16inter5, gate16inter6, gate16inter7, gate16inter8, gate16inter9, gate16inter10, gate16inter11, gate16inter12, gate241inter0, gate241inter1, gate241inter2, gate241inter3, gate241inter4, gate241inter5, gate241inter6, gate241inter7, gate241inter8, gate241inter9, gate241inter10, gate241inter11, gate241inter12, gate497inter0, gate497inter1, gate497inter2, gate497inter3, gate497inter4, gate497inter5, gate497inter6, gate497inter7, gate497inter8, gate497inter9, gate497inter10, gate497inter11, gate497inter12, gate485inter0, gate485inter1, gate485inter2, gate485inter3, gate485inter4, gate485inter5, gate485inter6, gate485inter7, gate485inter8, gate485inter9, gate485inter10, gate485inter11, gate485inter12, gate226inter0, gate226inter1, gate226inter2, gate226inter3, gate226inter4, gate226inter5, gate226inter6, gate226inter7, gate226inter8, gate226inter9, gate226inter10, gate226inter11, gate226inter12, gate186inter0, gate186inter1, gate186inter2, gate186inter3, gate186inter4, gate186inter5, gate186inter6, gate186inter7, gate186inter8, gate186inter9, gate186inter10, gate186inter11, gate186inter12, gate133inter0, gate133inter1, gate133inter2, gate133inter3, gate133inter4, gate133inter5, gate133inter6, gate133inter7, gate133inter8, gate133inter9, gate133inter10, gate133inter11, gate133inter12, gate285inter0, gate285inter1, gate285inter2, gate285inter3, gate285inter4, gate285inter5, gate285inter6, gate285inter7, gate285inter8, gate285inter9, gate285inter10, gate285inter11, gate285inter12, gate220inter0, gate220inter1, gate220inter2, gate220inter3, gate220inter4, gate220inter5, gate220inter6, gate220inter7, gate220inter8, gate220inter9, gate220inter10, gate220inter11, gate220inter12, gate244inter0, gate244inter1, gate244inter2, gate244inter3, gate244inter4, gate244inter5, gate244inter6, gate244inter7, gate244inter8, gate244inter9, gate244inter10, gate244inter11, gate244inter12, gate389inter0, gate389inter1, gate389inter2, gate389inter3, gate389inter4, gate389inter5, gate389inter6, gate389inter7, gate389inter8, gate389inter9, gate389inter10, gate389inter11, gate389inter12, gate420inter0, gate420inter1, gate420inter2, gate420inter3, gate420inter4, gate420inter5, gate420inter6, gate420inter7, gate420inter8, gate420inter9, gate420inter10, gate420inter11, gate420inter12, gate508inter0, gate508inter1, gate508inter2, gate508inter3, gate508inter4, gate508inter5, gate508inter6, gate508inter7, gate508inter8, gate508inter9, gate508inter10, gate508inter11, gate508inter12, gate74inter0, gate74inter1, gate74inter2, gate74inter3, gate74inter4, gate74inter5, gate74inter6, gate74inter7, gate74inter8, gate74inter9, gate74inter10, gate74inter11, gate74inter12, gate457inter0, gate457inter1, gate457inter2, gate457inter3, gate457inter4, gate457inter5, gate457inter6, gate457inter7, gate457inter8, gate457inter9, gate457inter10, gate457inter11, gate457inter12, gate265inter0, gate265inter1, gate265inter2, gate265inter3, gate265inter4, gate265inter5, gate265inter6, gate265inter7, gate265inter8, gate265inter9, gate265inter10, gate265inter11, gate265inter12, gate137inter0, gate137inter1, gate137inter2, gate137inter3, gate137inter4, gate137inter5, gate137inter6, gate137inter7, gate137inter8, gate137inter9, gate137inter10, gate137inter11, gate137inter12, gate207inter0, gate207inter1, gate207inter2, gate207inter3, gate207inter4, gate207inter5, gate207inter6, gate207inter7, gate207inter8, gate207inter9, gate207inter10, gate207inter11, gate207inter12, gate151inter0, gate151inter1, gate151inter2, gate151inter3, gate151inter4, gate151inter5, gate151inter6, gate151inter7, gate151inter8, gate151inter9, gate151inter10, gate151inter11, gate151inter12, gate210inter0, gate210inter1, gate210inter2, gate210inter3, gate210inter4, gate210inter5, gate210inter6, gate210inter7, gate210inter8, gate210inter9, gate210inter10, gate210inter11, gate210inter12, gate279inter0, gate279inter1, gate279inter2, gate279inter3, gate279inter4, gate279inter5, gate279inter6, gate279inter7, gate279inter8, gate279inter9, gate279inter10, gate279inter11, gate279inter12, gate182inter0, gate182inter1, gate182inter2, gate182inter3, gate182inter4, gate182inter5, gate182inter6, gate182inter7, gate182inter8, gate182inter9, gate182inter10, gate182inter11, gate182inter12, gate391inter0, gate391inter1, gate391inter2, gate391inter3, gate391inter4, gate391inter5, gate391inter6, gate391inter7, gate391inter8, gate391inter9, gate391inter10, gate391inter11, gate391inter12, gate294inter0, gate294inter1, gate294inter2, gate294inter3, gate294inter4, gate294inter5, gate294inter6, gate294inter7, gate294inter8, gate294inter9, gate294inter10, gate294inter11, gate294inter12, gate193inter0, gate193inter1, gate193inter2, gate193inter3, gate193inter4, gate193inter5, gate193inter6, gate193inter7, gate193inter8, gate193inter9, gate193inter10, gate193inter11, gate193inter12, gate46inter0, gate46inter1, gate46inter2, gate46inter3, gate46inter4, gate46inter5, gate46inter6, gate46inter7, gate46inter8, gate46inter9, gate46inter10, gate46inter11, gate46inter12, gate415inter0, gate415inter1, gate415inter2, gate415inter3, gate415inter4, gate415inter5, gate415inter6, gate415inter7, gate415inter8, gate415inter9, gate415inter10, gate415inter11, gate415inter12, gate476inter0, gate476inter1, gate476inter2, gate476inter3, gate476inter4, gate476inter5, gate476inter6, gate476inter7, gate476inter8, gate476inter9, gate476inter10, gate476inter11, gate476inter12, gate284inter0, gate284inter1, gate284inter2, gate284inter3, gate284inter4, gate284inter5, gate284inter6, gate284inter7, gate284inter8, gate284inter9, gate284inter10, gate284inter11, gate284inter12, gate245inter0, gate245inter1, gate245inter2, gate245inter3, gate245inter4, gate245inter5, gate245inter6, gate245inter7, gate245inter8, gate245inter9, gate245inter10, gate245inter11, gate245inter12, gate23inter0, gate23inter1, gate23inter2, gate23inter3, gate23inter4, gate23inter5, gate23inter6, gate23inter7, gate23inter8, gate23inter9, gate23inter10, gate23inter11, gate23inter12, gate60inter0, gate60inter1, gate60inter2, gate60inter3, gate60inter4, gate60inter5, gate60inter6, gate60inter7, gate60inter8, gate60inter9, gate60inter10, gate60inter11, gate60inter12, gate409inter0, gate409inter1, gate409inter2, gate409inter3, gate409inter4, gate409inter5, gate409inter6, gate409inter7, gate409inter8, gate409inter9, gate409inter10, gate409inter11, gate409inter12, gate243inter0, gate243inter1, gate243inter2, gate243inter3, gate243inter4, gate243inter5, gate243inter6, gate243inter7, gate243inter8, gate243inter9, gate243inter10, gate243inter11, gate243inter12, gate106inter0, gate106inter1, gate106inter2, gate106inter3, gate106inter4, gate106inter5, gate106inter6, gate106inter7, gate106inter8, gate106inter9, gate106inter10, gate106inter11, gate106inter12, gate171inter0, gate171inter1, gate171inter2, gate171inter3, gate171inter4, gate171inter5, gate171inter6, gate171inter7, gate171inter8, gate171inter9, gate171inter10, gate171inter11, gate171inter12, gate401inter0, gate401inter1, gate401inter2, gate401inter3, gate401inter4, gate401inter5, gate401inter6, gate401inter7, gate401inter8, gate401inter9, gate401inter10, gate401inter11, gate401inter12, gate292inter0, gate292inter1, gate292inter2, gate292inter3, gate292inter4, gate292inter5, gate292inter6, gate292inter7, gate292inter8, gate292inter9, gate292inter10, gate292inter11, gate292inter12, gate127inter0, gate127inter1, gate127inter2, gate127inter3, gate127inter4, gate127inter5, gate127inter6, gate127inter7, gate127inter8, gate127inter9, gate127inter10, gate127inter11, gate127inter12, gate185inter0, gate185inter1, gate185inter2, gate185inter3, gate185inter4, gate185inter5, gate185inter6, gate185inter7, gate185inter8, gate185inter9, gate185inter10, gate185inter11, gate185inter12, gate123inter0, gate123inter1, gate123inter2, gate123inter3, gate123inter4, gate123inter5, gate123inter6, gate123inter7, gate123inter8, gate123inter9, gate123inter10, gate123inter11, gate123inter12, gate273inter0, gate273inter1, gate273inter2, gate273inter3, gate273inter4, gate273inter5, gate273inter6, gate273inter7, gate273inter8, gate273inter9, gate273inter10, gate273inter11, gate273inter12, gate453inter0, gate453inter1, gate453inter2, gate453inter3, gate453inter4, gate453inter5, gate453inter6, gate453inter7, gate453inter8, gate453inter9, gate453inter10, gate453inter11, gate453inter12, gate257inter0, gate257inter1, gate257inter2, gate257inter3, gate257inter4, gate257inter5, gate257inter6, gate257inter7, gate257inter8, gate257inter9, gate257inter10, gate257inter11, gate257inter12, gate71inter0, gate71inter1, gate71inter2, gate71inter3, gate71inter4, gate71inter5, gate71inter6, gate71inter7, gate71inter8, gate71inter9, gate71inter10, gate71inter11, gate71inter12, gate205inter0, gate205inter1, gate205inter2, gate205inter3, gate205inter4, gate205inter5, gate205inter6, gate205inter7, gate205inter8, gate205inter9, gate205inter10, gate205inter11, gate205inter12, gate450inter0, gate450inter1, gate450inter2, gate450inter3, gate450inter4, gate450inter5, gate450inter6, gate450inter7, gate450inter8, gate450inter9, gate450inter10, gate450inter11, gate450inter12, gate90inter0, gate90inter1, gate90inter2, gate90inter3, gate90inter4, gate90inter5, gate90inter6, gate90inter7, gate90inter8, gate90inter9, gate90inter10, gate90inter11, gate90inter12, gate502inter0, gate502inter1, gate502inter2, gate502inter3, gate502inter4, gate502inter5, gate502inter6, gate502inter7, gate502inter8, gate502inter9, gate502inter10, gate502inter11, gate502inter12, gate162inter0, gate162inter1, gate162inter2, gate162inter3, gate162inter4, gate162inter5, gate162inter6, gate162inter7, gate162inter8, gate162inter9, gate162inter10, gate162inter11, gate162inter12, gate79inter0, gate79inter1, gate79inter2, gate79inter3, gate79inter4, gate79inter5, gate79inter6, gate79inter7, gate79inter8, gate79inter9, gate79inter10, gate79inter11, gate79inter12, gate173inter0, gate173inter1, gate173inter2, gate173inter3, gate173inter4, gate173inter5, gate173inter6, gate173inter7, gate173inter8, gate173inter9, gate173inter10, gate173inter11, gate173inter12, gate102inter0, gate102inter1, gate102inter2, gate102inter3, gate102inter4, gate102inter5, gate102inter6, gate102inter7, gate102inter8, gate102inter9, gate102inter10, gate102inter11, gate102inter12, gate471inter0, gate471inter1, gate471inter2, gate471inter3, gate471inter4, gate471inter5, gate471inter6, gate471inter7, gate471inter8, gate471inter9, gate471inter10, gate471inter11, gate471inter12, gate404inter0, gate404inter1, gate404inter2, gate404inter3, gate404inter4, gate404inter5, gate404inter6, gate404inter7, gate404inter8, gate404inter9, gate404inter10, gate404inter11, gate404inter12, gate252inter0, gate252inter1, gate252inter2, gate252inter3, gate252inter4, gate252inter5, gate252inter6, gate252inter7, gate252inter8, gate252inter9, gate252inter10, gate252inter11, gate252inter12, gate451inter0, gate451inter1, gate451inter2, gate451inter3, gate451inter4, gate451inter5, gate451inter6, gate451inter7, gate451inter8, gate451inter9, gate451inter10, gate451inter11, gate451inter12, gate189inter0, gate189inter1, gate189inter2, gate189inter3, gate189inter4, gate189inter5, gate189inter6, gate189inter7, gate189inter8, gate189inter9, gate189inter10, gate189inter11, gate189inter12, gate492inter0, gate492inter1, gate492inter2, gate492inter3, gate492inter4, gate492inter5, gate492inter6, gate492inter7, gate492inter8, gate492inter9, gate492inter10, gate492inter11, gate492inter12, gate424inter0, gate424inter1, gate424inter2, gate424inter3, gate424inter4, gate424inter5, gate424inter6, gate424inter7, gate424inter8, gate424inter9, gate424inter10, gate424inter11, gate424inter12, gate225inter0, gate225inter1, gate225inter2, gate225inter3, gate225inter4, gate225inter5, gate225inter6, gate225inter7, gate225inter8, gate225inter9, gate225inter10, gate225inter11, gate225inter12, gate49inter0, gate49inter1, gate49inter2, gate49inter3, gate49inter4, gate49inter5, gate49inter6, gate49inter7, gate49inter8, gate49inter9, gate49inter10, gate49inter11, gate49inter12;



and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );
nand2 gate9( .a(G1), .b(G2), .O(G266) );
nand2 gate10( .a(G3), .b(G4), .O(G269) );
nand2 gate11( .a(G5), .b(G6), .O(G272) );
nand2 gate12( .a(G7), .b(G8), .O(G275) );

  xor2  gate617(.a(G10), .b(G9), .O(gate13inter0));
  nand2 gate618(.a(gate13inter0), .b(s_10), .O(gate13inter1));
  and2  gate619(.a(G10), .b(G9), .O(gate13inter2));
  inv1  gate620(.a(s_10), .O(gate13inter3));
  inv1  gate621(.a(s_11), .O(gate13inter4));
  nand2 gate622(.a(gate13inter4), .b(gate13inter3), .O(gate13inter5));
  nor2  gate623(.a(gate13inter5), .b(gate13inter2), .O(gate13inter6));
  inv1  gate624(.a(G9), .O(gate13inter7));
  inv1  gate625(.a(G10), .O(gate13inter8));
  nand2 gate626(.a(gate13inter8), .b(gate13inter7), .O(gate13inter9));
  nand2 gate627(.a(s_11), .b(gate13inter3), .O(gate13inter10));
  nor2  gate628(.a(gate13inter10), .b(gate13inter9), .O(gate13inter11));
  nor2  gate629(.a(gate13inter11), .b(gate13inter6), .O(gate13inter12));
  nand2 gate630(.a(gate13inter12), .b(gate13inter1), .O(G278));
nand2 gate14( .a(G11), .b(G12), .O(G281) );
nand2 gate15( .a(G13), .b(G14), .O(G284) );

  xor2  gate1863(.a(G16), .b(G15), .O(gate16inter0));
  nand2 gate1864(.a(gate16inter0), .b(s_188), .O(gate16inter1));
  and2  gate1865(.a(G16), .b(G15), .O(gate16inter2));
  inv1  gate1866(.a(s_188), .O(gate16inter3));
  inv1  gate1867(.a(s_189), .O(gate16inter4));
  nand2 gate1868(.a(gate16inter4), .b(gate16inter3), .O(gate16inter5));
  nor2  gate1869(.a(gate16inter5), .b(gate16inter2), .O(gate16inter6));
  inv1  gate1870(.a(G15), .O(gate16inter7));
  inv1  gate1871(.a(G16), .O(gate16inter8));
  nand2 gate1872(.a(gate16inter8), .b(gate16inter7), .O(gate16inter9));
  nand2 gate1873(.a(s_189), .b(gate16inter3), .O(gate16inter10));
  nor2  gate1874(.a(gate16inter10), .b(gate16inter9), .O(gate16inter11));
  nor2  gate1875(.a(gate16inter11), .b(gate16inter6), .O(gate16inter12));
  nand2 gate1876(.a(gate16inter12), .b(gate16inter1), .O(G287));
nand2 gate17( .a(G17), .b(G18), .O(G290) );
nand2 gate18( .a(G19), .b(G20), .O(G293) );
nand2 gate19( .a(G21), .b(G22), .O(G296) );
nand2 gate20( .a(G23), .b(G24), .O(G299) );
nand2 gate21( .a(G25), .b(G26), .O(G302) );

  xor2  gate673(.a(G28), .b(G27), .O(gate22inter0));
  nand2 gate674(.a(gate22inter0), .b(s_18), .O(gate22inter1));
  and2  gate675(.a(G28), .b(G27), .O(gate22inter2));
  inv1  gate676(.a(s_18), .O(gate22inter3));
  inv1  gate677(.a(s_19), .O(gate22inter4));
  nand2 gate678(.a(gate22inter4), .b(gate22inter3), .O(gate22inter5));
  nor2  gate679(.a(gate22inter5), .b(gate22inter2), .O(gate22inter6));
  inv1  gate680(.a(G27), .O(gate22inter7));
  inv1  gate681(.a(G28), .O(gate22inter8));
  nand2 gate682(.a(gate22inter8), .b(gate22inter7), .O(gate22inter9));
  nand2 gate683(.a(s_19), .b(gate22inter3), .O(gate22inter10));
  nor2  gate684(.a(gate22inter10), .b(gate22inter9), .O(gate22inter11));
  nor2  gate685(.a(gate22inter11), .b(gate22inter6), .O(gate22inter12));
  nand2 gate686(.a(gate22inter12), .b(gate22inter1), .O(G305));

  xor2  gate2283(.a(G30), .b(G29), .O(gate23inter0));
  nand2 gate2284(.a(gate23inter0), .b(s_248), .O(gate23inter1));
  and2  gate2285(.a(G30), .b(G29), .O(gate23inter2));
  inv1  gate2286(.a(s_248), .O(gate23inter3));
  inv1  gate2287(.a(s_249), .O(gate23inter4));
  nand2 gate2288(.a(gate23inter4), .b(gate23inter3), .O(gate23inter5));
  nor2  gate2289(.a(gate23inter5), .b(gate23inter2), .O(gate23inter6));
  inv1  gate2290(.a(G29), .O(gate23inter7));
  inv1  gate2291(.a(G30), .O(gate23inter8));
  nand2 gate2292(.a(gate23inter8), .b(gate23inter7), .O(gate23inter9));
  nand2 gate2293(.a(s_249), .b(gate23inter3), .O(gate23inter10));
  nor2  gate2294(.a(gate23inter10), .b(gate23inter9), .O(gate23inter11));
  nor2  gate2295(.a(gate23inter11), .b(gate23inter6), .O(gate23inter12));
  nand2 gate2296(.a(gate23inter12), .b(gate23inter1), .O(G308));
nand2 gate24( .a(G31), .b(G32), .O(G311) );

  xor2  gate799(.a(G5), .b(G1), .O(gate25inter0));
  nand2 gate800(.a(gate25inter0), .b(s_36), .O(gate25inter1));
  and2  gate801(.a(G5), .b(G1), .O(gate25inter2));
  inv1  gate802(.a(s_36), .O(gate25inter3));
  inv1  gate803(.a(s_37), .O(gate25inter4));
  nand2 gate804(.a(gate25inter4), .b(gate25inter3), .O(gate25inter5));
  nor2  gate805(.a(gate25inter5), .b(gate25inter2), .O(gate25inter6));
  inv1  gate806(.a(G1), .O(gate25inter7));
  inv1  gate807(.a(G5), .O(gate25inter8));
  nand2 gate808(.a(gate25inter8), .b(gate25inter7), .O(gate25inter9));
  nand2 gate809(.a(s_37), .b(gate25inter3), .O(gate25inter10));
  nor2  gate810(.a(gate25inter10), .b(gate25inter9), .O(gate25inter11));
  nor2  gate811(.a(gate25inter11), .b(gate25inter6), .O(gate25inter12));
  nand2 gate812(.a(gate25inter12), .b(gate25inter1), .O(G314));

  xor2  gate869(.a(G13), .b(G9), .O(gate26inter0));
  nand2 gate870(.a(gate26inter0), .b(s_46), .O(gate26inter1));
  and2  gate871(.a(G13), .b(G9), .O(gate26inter2));
  inv1  gate872(.a(s_46), .O(gate26inter3));
  inv1  gate873(.a(s_47), .O(gate26inter4));
  nand2 gate874(.a(gate26inter4), .b(gate26inter3), .O(gate26inter5));
  nor2  gate875(.a(gate26inter5), .b(gate26inter2), .O(gate26inter6));
  inv1  gate876(.a(G9), .O(gate26inter7));
  inv1  gate877(.a(G13), .O(gate26inter8));
  nand2 gate878(.a(gate26inter8), .b(gate26inter7), .O(gate26inter9));
  nand2 gate879(.a(s_47), .b(gate26inter3), .O(gate26inter10));
  nor2  gate880(.a(gate26inter10), .b(gate26inter9), .O(gate26inter11));
  nor2  gate881(.a(gate26inter11), .b(gate26inter6), .O(gate26inter12));
  nand2 gate882(.a(gate26inter12), .b(gate26inter1), .O(G317));
nand2 gate27( .a(G2), .b(G6), .O(G320) );

  xor2  gate1765(.a(G14), .b(G10), .O(gate28inter0));
  nand2 gate1766(.a(gate28inter0), .b(s_174), .O(gate28inter1));
  and2  gate1767(.a(G14), .b(G10), .O(gate28inter2));
  inv1  gate1768(.a(s_174), .O(gate28inter3));
  inv1  gate1769(.a(s_175), .O(gate28inter4));
  nand2 gate1770(.a(gate28inter4), .b(gate28inter3), .O(gate28inter5));
  nor2  gate1771(.a(gate28inter5), .b(gate28inter2), .O(gate28inter6));
  inv1  gate1772(.a(G10), .O(gate28inter7));
  inv1  gate1773(.a(G14), .O(gate28inter8));
  nand2 gate1774(.a(gate28inter8), .b(gate28inter7), .O(gate28inter9));
  nand2 gate1775(.a(s_175), .b(gate28inter3), .O(gate28inter10));
  nor2  gate1776(.a(gate28inter10), .b(gate28inter9), .O(gate28inter11));
  nor2  gate1777(.a(gate28inter11), .b(gate28inter6), .O(gate28inter12));
  nand2 gate1778(.a(gate28inter12), .b(gate28inter1), .O(G323));
nand2 gate29( .a(G3), .b(G7), .O(G326) );
nand2 gate30( .a(G11), .b(G15), .O(G329) );

  xor2  gate1247(.a(G8), .b(G4), .O(gate31inter0));
  nand2 gate1248(.a(gate31inter0), .b(s_100), .O(gate31inter1));
  and2  gate1249(.a(G8), .b(G4), .O(gate31inter2));
  inv1  gate1250(.a(s_100), .O(gate31inter3));
  inv1  gate1251(.a(s_101), .O(gate31inter4));
  nand2 gate1252(.a(gate31inter4), .b(gate31inter3), .O(gate31inter5));
  nor2  gate1253(.a(gate31inter5), .b(gate31inter2), .O(gate31inter6));
  inv1  gate1254(.a(G4), .O(gate31inter7));
  inv1  gate1255(.a(G8), .O(gate31inter8));
  nand2 gate1256(.a(gate31inter8), .b(gate31inter7), .O(gate31inter9));
  nand2 gate1257(.a(s_101), .b(gate31inter3), .O(gate31inter10));
  nor2  gate1258(.a(gate31inter10), .b(gate31inter9), .O(gate31inter11));
  nor2  gate1259(.a(gate31inter11), .b(gate31inter6), .O(gate31inter12));
  nand2 gate1260(.a(gate31inter12), .b(gate31inter1), .O(G332));
nand2 gate32( .a(G12), .b(G16), .O(G335) );
nand2 gate33( .a(G17), .b(G21), .O(G338) );
nand2 gate34( .a(G25), .b(G29), .O(G341) );
nand2 gate35( .a(G18), .b(G22), .O(G344) );

  xor2  gate1121(.a(G30), .b(G26), .O(gate36inter0));
  nand2 gate1122(.a(gate36inter0), .b(s_82), .O(gate36inter1));
  and2  gate1123(.a(G30), .b(G26), .O(gate36inter2));
  inv1  gate1124(.a(s_82), .O(gate36inter3));
  inv1  gate1125(.a(s_83), .O(gate36inter4));
  nand2 gate1126(.a(gate36inter4), .b(gate36inter3), .O(gate36inter5));
  nor2  gate1127(.a(gate36inter5), .b(gate36inter2), .O(gate36inter6));
  inv1  gate1128(.a(G26), .O(gate36inter7));
  inv1  gate1129(.a(G30), .O(gate36inter8));
  nand2 gate1130(.a(gate36inter8), .b(gate36inter7), .O(gate36inter9));
  nand2 gate1131(.a(s_83), .b(gate36inter3), .O(gate36inter10));
  nor2  gate1132(.a(gate36inter10), .b(gate36inter9), .O(gate36inter11));
  nor2  gate1133(.a(gate36inter11), .b(gate36inter6), .O(gate36inter12));
  nand2 gate1134(.a(gate36inter12), .b(gate36inter1), .O(G347));
nand2 gate37( .a(G19), .b(G23), .O(G350) );

  xor2  gate1681(.a(G31), .b(G27), .O(gate38inter0));
  nand2 gate1682(.a(gate38inter0), .b(s_162), .O(gate38inter1));
  and2  gate1683(.a(G31), .b(G27), .O(gate38inter2));
  inv1  gate1684(.a(s_162), .O(gate38inter3));
  inv1  gate1685(.a(s_163), .O(gate38inter4));
  nand2 gate1686(.a(gate38inter4), .b(gate38inter3), .O(gate38inter5));
  nor2  gate1687(.a(gate38inter5), .b(gate38inter2), .O(gate38inter6));
  inv1  gate1688(.a(G27), .O(gate38inter7));
  inv1  gate1689(.a(G31), .O(gate38inter8));
  nand2 gate1690(.a(gate38inter8), .b(gate38inter7), .O(gate38inter9));
  nand2 gate1691(.a(s_163), .b(gate38inter3), .O(gate38inter10));
  nor2  gate1692(.a(gate38inter10), .b(gate38inter9), .O(gate38inter11));
  nor2  gate1693(.a(gate38inter11), .b(gate38inter6), .O(gate38inter12));
  nand2 gate1694(.a(gate38inter12), .b(gate38inter1), .O(G353));
nand2 gate39( .a(G20), .b(G24), .O(G356) );
nand2 gate40( .a(G28), .b(G32), .O(G359) );

  xor2  gate757(.a(G266), .b(G1), .O(gate41inter0));
  nand2 gate758(.a(gate41inter0), .b(s_30), .O(gate41inter1));
  and2  gate759(.a(G266), .b(G1), .O(gate41inter2));
  inv1  gate760(.a(s_30), .O(gate41inter3));
  inv1  gate761(.a(s_31), .O(gate41inter4));
  nand2 gate762(.a(gate41inter4), .b(gate41inter3), .O(gate41inter5));
  nor2  gate763(.a(gate41inter5), .b(gate41inter2), .O(gate41inter6));
  inv1  gate764(.a(G1), .O(gate41inter7));
  inv1  gate765(.a(G266), .O(gate41inter8));
  nand2 gate766(.a(gate41inter8), .b(gate41inter7), .O(gate41inter9));
  nand2 gate767(.a(s_31), .b(gate41inter3), .O(gate41inter10));
  nor2  gate768(.a(gate41inter10), .b(gate41inter9), .O(gate41inter11));
  nor2  gate769(.a(gate41inter11), .b(gate41inter6), .O(gate41inter12));
  nand2 gate770(.a(gate41inter12), .b(gate41inter1), .O(G362));
nand2 gate42( .a(G2), .b(G266), .O(G363) );
nand2 gate43( .a(G3), .b(G269), .O(G364) );
nand2 gate44( .a(G4), .b(G269), .O(G365) );
nand2 gate45( .a(G5), .b(G272), .O(G366) );

  xor2  gate2213(.a(G272), .b(G6), .O(gate46inter0));
  nand2 gate2214(.a(gate46inter0), .b(s_238), .O(gate46inter1));
  and2  gate2215(.a(G272), .b(G6), .O(gate46inter2));
  inv1  gate2216(.a(s_238), .O(gate46inter3));
  inv1  gate2217(.a(s_239), .O(gate46inter4));
  nand2 gate2218(.a(gate46inter4), .b(gate46inter3), .O(gate46inter5));
  nor2  gate2219(.a(gate46inter5), .b(gate46inter2), .O(gate46inter6));
  inv1  gate2220(.a(G6), .O(gate46inter7));
  inv1  gate2221(.a(G272), .O(gate46inter8));
  nand2 gate2222(.a(gate46inter8), .b(gate46inter7), .O(gate46inter9));
  nand2 gate2223(.a(s_239), .b(gate46inter3), .O(gate46inter10));
  nor2  gate2224(.a(gate46inter10), .b(gate46inter9), .O(gate46inter11));
  nor2  gate2225(.a(gate46inter11), .b(gate46inter6), .O(gate46inter12));
  nand2 gate2226(.a(gate46inter12), .b(gate46inter1), .O(G367));

  xor2  gate1317(.a(G275), .b(G7), .O(gate47inter0));
  nand2 gate1318(.a(gate47inter0), .b(s_110), .O(gate47inter1));
  and2  gate1319(.a(G275), .b(G7), .O(gate47inter2));
  inv1  gate1320(.a(s_110), .O(gate47inter3));
  inv1  gate1321(.a(s_111), .O(gate47inter4));
  nand2 gate1322(.a(gate47inter4), .b(gate47inter3), .O(gate47inter5));
  nor2  gate1323(.a(gate47inter5), .b(gate47inter2), .O(gate47inter6));
  inv1  gate1324(.a(G7), .O(gate47inter7));
  inv1  gate1325(.a(G275), .O(gate47inter8));
  nand2 gate1326(.a(gate47inter8), .b(gate47inter7), .O(gate47inter9));
  nand2 gate1327(.a(s_111), .b(gate47inter3), .O(gate47inter10));
  nor2  gate1328(.a(gate47inter10), .b(gate47inter9), .O(gate47inter11));
  nor2  gate1329(.a(gate47inter11), .b(gate47inter6), .O(gate47inter12));
  nand2 gate1330(.a(gate47inter12), .b(gate47inter1), .O(G368));
nand2 gate48( .a(G8), .b(G275), .O(G369) );

  xor2  gate2717(.a(G278), .b(G9), .O(gate49inter0));
  nand2 gate2718(.a(gate49inter0), .b(s_310), .O(gate49inter1));
  and2  gate2719(.a(G278), .b(G9), .O(gate49inter2));
  inv1  gate2720(.a(s_310), .O(gate49inter3));
  inv1  gate2721(.a(s_311), .O(gate49inter4));
  nand2 gate2722(.a(gate49inter4), .b(gate49inter3), .O(gate49inter5));
  nor2  gate2723(.a(gate49inter5), .b(gate49inter2), .O(gate49inter6));
  inv1  gate2724(.a(G9), .O(gate49inter7));
  inv1  gate2725(.a(G278), .O(gate49inter8));
  nand2 gate2726(.a(gate49inter8), .b(gate49inter7), .O(gate49inter9));
  nand2 gate2727(.a(s_311), .b(gate49inter3), .O(gate49inter10));
  nor2  gate2728(.a(gate49inter10), .b(gate49inter9), .O(gate49inter11));
  nor2  gate2729(.a(gate49inter11), .b(gate49inter6), .O(gate49inter12));
  nand2 gate2730(.a(gate49inter12), .b(gate49inter1), .O(G370));
nand2 gate50( .a(G10), .b(G278), .O(G371) );
nand2 gate51( .a(G11), .b(G281), .O(G372) );

  xor2  gate715(.a(G281), .b(G12), .O(gate52inter0));
  nand2 gate716(.a(gate52inter0), .b(s_24), .O(gate52inter1));
  and2  gate717(.a(G281), .b(G12), .O(gate52inter2));
  inv1  gate718(.a(s_24), .O(gate52inter3));
  inv1  gate719(.a(s_25), .O(gate52inter4));
  nand2 gate720(.a(gate52inter4), .b(gate52inter3), .O(gate52inter5));
  nor2  gate721(.a(gate52inter5), .b(gate52inter2), .O(gate52inter6));
  inv1  gate722(.a(G12), .O(gate52inter7));
  inv1  gate723(.a(G281), .O(gate52inter8));
  nand2 gate724(.a(gate52inter8), .b(gate52inter7), .O(gate52inter9));
  nand2 gate725(.a(s_25), .b(gate52inter3), .O(gate52inter10));
  nor2  gate726(.a(gate52inter10), .b(gate52inter9), .O(gate52inter11));
  nor2  gate727(.a(gate52inter11), .b(gate52inter6), .O(gate52inter12));
  nand2 gate728(.a(gate52inter12), .b(gate52inter1), .O(G373));
nand2 gate53( .a(G13), .b(G284), .O(G374) );
nand2 gate54( .a(G14), .b(G284), .O(G375) );

  xor2  gate967(.a(G287), .b(G15), .O(gate55inter0));
  nand2 gate968(.a(gate55inter0), .b(s_60), .O(gate55inter1));
  and2  gate969(.a(G287), .b(G15), .O(gate55inter2));
  inv1  gate970(.a(s_60), .O(gate55inter3));
  inv1  gate971(.a(s_61), .O(gate55inter4));
  nand2 gate972(.a(gate55inter4), .b(gate55inter3), .O(gate55inter5));
  nor2  gate973(.a(gate55inter5), .b(gate55inter2), .O(gate55inter6));
  inv1  gate974(.a(G15), .O(gate55inter7));
  inv1  gate975(.a(G287), .O(gate55inter8));
  nand2 gate976(.a(gate55inter8), .b(gate55inter7), .O(gate55inter9));
  nand2 gate977(.a(s_61), .b(gate55inter3), .O(gate55inter10));
  nor2  gate978(.a(gate55inter10), .b(gate55inter9), .O(gate55inter11));
  nor2  gate979(.a(gate55inter11), .b(gate55inter6), .O(gate55inter12));
  nand2 gate980(.a(gate55inter12), .b(gate55inter1), .O(G376));
nand2 gate56( .a(G16), .b(G287), .O(G377) );

  xor2  gate1093(.a(G290), .b(G17), .O(gate57inter0));
  nand2 gate1094(.a(gate57inter0), .b(s_78), .O(gate57inter1));
  and2  gate1095(.a(G290), .b(G17), .O(gate57inter2));
  inv1  gate1096(.a(s_78), .O(gate57inter3));
  inv1  gate1097(.a(s_79), .O(gate57inter4));
  nand2 gate1098(.a(gate57inter4), .b(gate57inter3), .O(gate57inter5));
  nor2  gate1099(.a(gate57inter5), .b(gate57inter2), .O(gate57inter6));
  inv1  gate1100(.a(G17), .O(gate57inter7));
  inv1  gate1101(.a(G290), .O(gate57inter8));
  nand2 gate1102(.a(gate57inter8), .b(gate57inter7), .O(gate57inter9));
  nand2 gate1103(.a(s_79), .b(gate57inter3), .O(gate57inter10));
  nor2  gate1104(.a(gate57inter10), .b(gate57inter9), .O(gate57inter11));
  nor2  gate1105(.a(gate57inter11), .b(gate57inter6), .O(gate57inter12));
  nand2 gate1106(.a(gate57inter12), .b(gate57inter1), .O(G378));
nand2 gate58( .a(G18), .b(G290), .O(G379) );

  xor2  gate603(.a(G293), .b(G19), .O(gate59inter0));
  nand2 gate604(.a(gate59inter0), .b(s_8), .O(gate59inter1));
  and2  gate605(.a(G293), .b(G19), .O(gate59inter2));
  inv1  gate606(.a(s_8), .O(gate59inter3));
  inv1  gate607(.a(s_9), .O(gate59inter4));
  nand2 gate608(.a(gate59inter4), .b(gate59inter3), .O(gate59inter5));
  nor2  gate609(.a(gate59inter5), .b(gate59inter2), .O(gate59inter6));
  inv1  gate610(.a(G19), .O(gate59inter7));
  inv1  gate611(.a(G293), .O(gate59inter8));
  nand2 gate612(.a(gate59inter8), .b(gate59inter7), .O(gate59inter9));
  nand2 gate613(.a(s_9), .b(gate59inter3), .O(gate59inter10));
  nor2  gate614(.a(gate59inter10), .b(gate59inter9), .O(gate59inter11));
  nor2  gate615(.a(gate59inter11), .b(gate59inter6), .O(gate59inter12));
  nand2 gate616(.a(gate59inter12), .b(gate59inter1), .O(G380));

  xor2  gate2297(.a(G293), .b(G20), .O(gate60inter0));
  nand2 gate2298(.a(gate60inter0), .b(s_250), .O(gate60inter1));
  and2  gate2299(.a(G293), .b(G20), .O(gate60inter2));
  inv1  gate2300(.a(s_250), .O(gate60inter3));
  inv1  gate2301(.a(s_251), .O(gate60inter4));
  nand2 gate2302(.a(gate60inter4), .b(gate60inter3), .O(gate60inter5));
  nor2  gate2303(.a(gate60inter5), .b(gate60inter2), .O(gate60inter6));
  inv1  gate2304(.a(G20), .O(gate60inter7));
  inv1  gate2305(.a(G293), .O(gate60inter8));
  nand2 gate2306(.a(gate60inter8), .b(gate60inter7), .O(gate60inter9));
  nand2 gate2307(.a(s_251), .b(gate60inter3), .O(gate60inter10));
  nor2  gate2308(.a(gate60inter10), .b(gate60inter9), .O(gate60inter11));
  nor2  gate2309(.a(gate60inter11), .b(gate60inter6), .O(gate60inter12));
  nand2 gate2310(.a(gate60inter12), .b(gate60inter1), .O(G381));
nand2 gate61( .a(G21), .b(G296), .O(G382) );
nand2 gate62( .a(G22), .b(G296), .O(G383) );
nand2 gate63( .a(G23), .b(G299), .O(G384) );

  xor2  gate1219(.a(G299), .b(G24), .O(gate64inter0));
  nand2 gate1220(.a(gate64inter0), .b(s_96), .O(gate64inter1));
  and2  gate1221(.a(G299), .b(G24), .O(gate64inter2));
  inv1  gate1222(.a(s_96), .O(gate64inter3));
  inv1  gate1223(.a(s_97), .O(gate64inter4));
  nand2 gate1224(.a(gate64inter4), .b(gate64inter3), .O(gate64inter5));
  nor2  gate1225(.a(gate64inter5), .b(gate64inter2), .O(gate64inter6));
  inv1  gate1226(.a(G24), .O(gate64inter7));
  inv1  gate1227(.a(G299), .O(gate64inter8));
  nand2 gate1228(.a(gate64inter8), .b(gate64inter7), .O(gate64inter9));
  nand2 gate1229(.a(s_97), .b(gate64inter3), .O(gate64inter10));
  nor2  gate1230(.a(gate64inter10), .b(gate64inter9), .O(gate64inter11));
  nor2  gate1231(.a(gate64inter11), .b(gate64inter6), .O(gate64inter12));
  nand2 gate1232(.a(gate64inter12), .b(gate64inter1), .O(G385));

  xor2  gate687(.a(G302), .b(G25), .O(gate65inter0));
  nand2 gate688(.a(gate65inter0), .b(s_20), .O(gate65inter1));
  and2  gate689(.a(G302), .b(G25), .O(gate65inter2));
  inv1  gate690(.a(s_20), .O(gate65inter3));
  inv1  gate691(.a(s_21), .O(gate65inter4));
  nand2 gate692(.a(gate65inter4), .b(gate65inter3), .O(gate65inter5));
  nor2  gate693(.a(gate65inter5), .b(gate65inter2), .O(gate65inter6));
  inv1  gate694(.a(G25), .O(gate65inter7));
  inv1  gate695(.a(G302), .O(gate65inter8));
  nand2 gate696(.a(gate65inter8), .b(gate65inter7), .O(gate65inter9));
  nand2 gate697(.a(s_21), .b(gate65inter3), .O(gate65inter10));
  nor2  gate698(.a(gate65inter10), .b(gate65inter9), .O(gate65inter11));
  nor2  gate699(.a(gate65inter11), .b(gate65inter6), .O(gate65inter12));
  nand2 gate700(.a(gate65inter12), .b(gate65inter1), .O(G386));
nand2 gate66( .a(G26), .b(G302), .O(G387) );
nand2 gate67( .a(G27), .b(G305), .O(G388) );
nand2 gate68( .a(G28), .b(G305), .O(G389) );

  xor2  gate1149(.a(G308), .b(G29), .O(gate69inter0));
  nand2 gate1150(.a(gate69inter0), .b(s_86), .O(gate69inter1));
  and2  gate1151(.a(G308), .b(G29), .O(gate69inter2));
  inv1  gate1152(.a(s_86), .O(gate69inter3));
  inv1  gate1153(.a(s_87), .O(gate69inter4));
  nand2 gate1154(.a(gate69inter4), .b(gate69inter3), .O(gate69inter5));
  nor2  gate1155(.a(gate69inter5), .b(gate69inter2), .O(gate69inter6));
  inv1  gate1156(.a(G29), .O(gate69inter7));
  inv1  gate1157(.a(G308), .O(gate69inter8));
  nand2 gate1158(.a(gate69inter8), .b(gate69inter7), .O(gate69inter9));
  nand2 gate1159(.a(s_87), .b(gate69inter3), .O(gate69inter10));
  nor2  gate1160(.a(gate69inter10), .b(gate69inter9), .O(gate69inter11));
  nor2  gate1161(.a(gate69inter11), .b(gate69inter6), .O(gate69inter12));
  nand2 gate1162(.a(gate69inter12), .b(gate69inter1), .O(G390));
nand2 gate70( .a(G30), .b(G308), .O(G391) );

  xor2  gate2479(.a(G311), .b(G31), .O(gate71inter0));
  nand2 gate2480(.a(gate71inter0), .b(s_276), .O(gate71inter1));
  and2  gate2481(.a(G311), .b(G31), .O(gate71inter2));
  inv1  gate2482(.a(s_276), .O(gate71inter3));
  inv1  gate2483(.a(s_277), .O(gate71inter4));
  nand2 gate2484(.a(gate71inter4), .b(gate71inter3), .O(gate71inter5));
  nor2  gate2485(.a(gate71inter5), .b(gate71inter2), .O(gate71inter6));
  inv1  gate2486(.a(G31), .O(gate71inter7));
  inv1  gate2487(.a(G311), .O(gate71inter8));
  nand2 gate2488(.a(gate71inter8), .b(gate71inter7), .O(gate71inter9));
  nand2 gate2489(.a(s_277), .b(gate71inter3), .O(gate71inter10));
  nor2  gate2490(.a(gate71inter10), .b(gate71inter9), .O(gate71inter11));
  nor2  gate2491(.a(gate71inter11), .b(gate71inter6), .O(gate71inter12));
  nand2 gate2492(.a(gate71inter12), .b(gate71inter1), .O(G392));

  xor2  gate1471(.a(G311), .b(G32), .O(gate72inter0));
  nand2 gate1472(.a(gate72inter0), .b(s_132), .O(gate72inter1));
  and2  gate1473(.a(G311), .b(G32), .O(gate72inter2));
  inv1  gate1474(.a(s_132), .O(gate72inter3));
  inv1  gate1475(.a(s_133), .O(gate72inter4));
  nand2 gate1476(.a(gate72inter4), .b(gate72inter3), .O(gate72inter5));
  nor2  gate1477(.a(gate72inter5), .b(gate72inter2), .O(gate72inter6));
  inv1  gate1478(.a(G32), .O(gate72inter7));
  inv1  gate1479(.a(G311), .O(gate72inter8));
  nand2 gate1480(.a(gate72inter8), .b(gate72inter7), .O(gate72inter9));
  nand2 gate1481(.a(s_133), .b(gate72inter3), .O(gate72inter10));
  nor2  gate1482(.a(gate72inter10), .b(gate72inter9), .O(gate72inter11));
  nor2  gate1483(.a(gate72inter11), .b(gate72inter6), .O(gate72inter12));
  nand2 gate1484(.a(gate72inter12), .b(gate72inter1), .O(G393));
nand2 gate73( .a(G1), .b(G314), .O(G394) );

  xor2  gate2045(.a(G314), .b(G5), .O(gate74inter0));
  nand2 gate2046(.a(gate74inter0), .b(s_214), .O(gate74inter1));
  and2  gate2047(.a(G314), .b(G5), .O(gate74inter2));
  inv1  gate2048(.a(s_214), .O(gate74inter3));
  inv1  gate2049(.a(s_215), .O(gate74inter4));
  nand2 gate2050(.a(gate74inter4), .b(gate74inter3), .O(gate74inter5));
  nor2  gate2051(.a(gate74inter5), .b(gate74inter2), .O(gate74inter6));
  inv1  gate2052(.a(G5), .O(gate74inter7));
  inv1  gate2053(.a(G314), .O(gate74inter8));
  nand2 gate2054(.a(gate74inter8), .b(gate74inter7), .O(gate74inter9));
  nand2 gate2055(.a(s_215), .b(gate74inter3), .O(gate74inter10));
  nor2  gate2056(.a(gate74inter10), .b(gate74inter9), .O(gate74inter11));
  nor2  gate2057(.a(gate74inter11), .b(gate74inter6), .O(gate74inter12));
  nand2 gate2058(.a(gate74inter12), .b(gate74inter1), .O(G395));
nand2 gate75( .a(G9), .b(G317), .O(G396) );
nand2 gate76( .a(G13), .b(G317), .O(G397) );
nand2 gate77( .a(G2), .b(G320), .O(G398) );
nand2 gate78( .a(G6), .b(G320), .O(G399) );

  xor2  gate2563(.a(G323), .b(G10), .O(gate79inter0));
  nand2 gate2564(.a(gate79inter0), .b(s_288), .O(gate79inter1));
  and2  gate2565(.a(G323), .b(G10), .O(gate79inter2));
  inv1  gate2566(.a(s_288), .O(gate79inter3));
  inv1  gate2567(.a(s_289), .O(gate79inter4));
  nand2 gate2568(.a(gate79inter4), .b(gate79inter3), .O(gate79inter5));
  nor2  gate2569(.a(gate79inter5), .b(gate79inter2), .O(gate79inter6));
  inv1  gate2570(.a(G10), .O(gate79inter7));
  inv1  gate2571(.a(G323), .O(gate79inter8));
  nand2 gate2572(.a(gate79inter8), .b(gate79inter7), .O(gate79inter9));
  nand2 gate2573(.a(s_289), .b(gate79inter3), .O(gate79inter10));
  nor2  gate2574(.a(gate79inter10), .b(gate79inter9), .O(gate79inter11));
  nor2  gate2575(.a(gate79inter11), .b(gate79inter6), .O(gate79inter12));
  nand2 gate2576(.a(gate79inter12), .b(gate79inter1), .O(G400));
nand2 gate80( .a(G14), .b(G323), .O(G401) );

  xor2  gate1485(.a(G326), .b(G3), .O(gate81inter0));
  nand2 gate1486(.a(gate81inter0), .b(s_134), .O(gate81inter1));
  and2  gate1487(.a(G326), .b(G3), .O(gate81inter2));
  inv1  gate1488(.a(s_134), .O(gate81inter3));
  inv1  gate1489(.a(s_135), .O(gate81inter4));
  nand2 gate1490(.a(gate81inter4), .b(gate81inter3), .O(gate81inter5));
  nor2  gate1491(.a(gate81inter5), .b(gate81inter2), .O(gate81inter6));
  inv1  gate1492(.a(G3), .O(gate81inter7));
  inv1  gate1493(.a(G326), .O(gate81inter8));
  nand2 gate1494(.a(gate81inter8), .b(gate81inter7), .O(gate81inter9));
  nand2 gate1495(.a(s_135), .b(gate81inter3), .O(gate81inter10));
  nor2  gate1496(.a(gate81inter10), .b(gate81inter9), .O(gate81inter11));
  nor2  gate1497(.a(gate81inter11), .b(gate81inter6), .O(gate81inter12));
  nand2 gate1498(.a(gate81inter12), .b(gate81inter1), .O(G402));

  xor2  gate1107(.a(G326), .b(G7), .O(gate82inter0));
  nand2 gate1108(.a(gate82inter0), .b(s_80), .O(gate82inter1));
  and2  gate1109(.a(G326), .b(G7), .O(gate82inter2));
  inv1  gate1110(.a(s_80), .O(gate82inter3));
  inv1  gate1111(.a(s_81), .O(gate82inter4));
  nand2 gate1112(.a(gate82inter4), .b(gate82inter3), .O(gate82inter5));
  nor2  gate1113(.a(gate82inter5), .b(gate82inter2), .O(gate82inter6));
  inv1  gate1114(.a(G7), .O(gate82inter7));
  inv1  gate1115(.a(G326), .O(gate82inter8));
  nand2 gate1116(.a(gate82inter8), .b(gate82inter7), .O(gate82inter9));
  nand2 gate1117(.a(s_81), .b(gate82inter3), .O(gate82inter10));
  nor2  gate1118(.a(gate82inter10), .b(gate82inter9), .O(gate82inter11));
  nor2  gate1119(.a(gate82inter11), .b(gate82inter6), .O(gate82inter12));
  nand2 gate1120(.a(gate82inter12), .b(gate82inter1), .O(G403));
nand2 gate83( .a(G11), .b(G329), .O(G404) );
nand2 gate84( .a(G15), .b(G329), .O(G405) );

  xor2  gate883(.a(G332), .b(G4), .O(gate85inter0));
  nand2 gate884(.a(gate85inter0), .b(s_48), .O(gate85inter1));
  and2  gate885(.a(G332), .b(G4), .O(gate85inter2));
  inv1  gate886(.a(s_48), .O(gate85inter3));
  inv1  gate887(.a(s_49), .O(gate85inter4));
  nand2 gate888(.a(gate85inter4), .b(gate85inter3), .O(gate85inter5));
  nor2  gate889(.a(gate85inter5), .b(gate85inter2), .O(gate85inter6));
  inv1  gate890(.a(G4), .O(gate85inter7));
  inv1  gate891(.a(G332), .O(gate85inter8));
  nand2 gate892(.a(gate85inter8), .b(gate85inter7), .O(gate85inter9));
  nand2 gate893(.a(s_49), .b(gate85inter3), .O(gate85inter10));
  nor2  gate894(.a(gate85inter10), .b(gate85inter9), .O(gate85inter11));
  nor2  gate895(.a(gate85inter11), .b(gate85inter6), .O(gate85inter12));
  nand2 gate896(.a(gate85inter12), .b(gate85inter1), .O(G406));
nand2 gate86( .a(G8), .b(G332), .O(G407) );
nand2 gate87( .a(G12), .b(G335), .O(G408) );

  xor2  gate1023(.a(G335), .b(G16), .O(gate88inter0));
  nand2 gate1024(.a(gate88inter0), .b(s_68), .O(gate88inter1));
  and2  gate1025(.a(G335), .b(G16), .O(gate88inter2));
  inv1  gate1026(.a(s_68), .O(gate88inter3));
  inv1  gate1027(.a(s_69), .O(gate88inter4));
  nand2 gate1028(.a(gate88inter4), .b(gate88inter3), .O(gate88inter5));
  nor2  gate1029(.a(gate88inter5), .b(gate88inter2), .O(gate88inter6));
  inv1  gate1030(.a(G16), .O(gate88inter7));
  inv1  gate1031(.a(G335), .O(gate88inter8));
  nand2 gate1032(.a(gate88inter8), .b(gate88inter7), .O(gate88inter9));
  nand2 gate1033(.a(s_69), .b(gate88inter3), .O(gate88inter10));
  nor2  gate1034(.a(gate88inter10), .b(gate88inter9), .O(gate88inter11));
  nor2  gate1035(.a(gate88inter11), .b(gate88inter6), .O(gate88inter12));
  nand2 gate1036(.a(gate88inter12), .b(gate88inter1), .O(G409));

  xor2  gate1401(.a(G338), .b(G17), .O(gate89inter0));
  nand2 gate1402(.a(gate89inter0), .b(s_122), .O(gate89inter1));
  and2  gate1403(.a(G338), .b(G17), .O(gate89inter2));
  inv1  gate1404(.a(s_122), .O(gate89inter3));
  inv1  gate1405(.a(s_123), .O(gate89inter4));
  nand2 gate1406(.a(gate89inter4), .b(gate89inter3), .O(gate89inter5));
  nor2  gate1407(.a(gate89inter5), .b(gate89inter2), .O(gate89inter6));
  inv1  gate1408(.a(G17), .O(gate89inter7));
  inv1  gate1409(.a(G338), .O(gate89inter8));
  nand2 gate1410(.a(gate89inter8), .b(gate89inter7), .O(gate89inter9));
  nand2 gate1411(.a(s_123), .b(gate89inter3), .O(gate89inter10));
  nor2  gate1412(.a(gate89inter10), .b(gate89inter9), .O(gate89inter11));
  nor2  gate1413(.a(gate89inter11), .b(gate89inter6), .O(gate89inter12));
  nand2 gate1414(.a(gate89inter12), .b(gate89inter1), .O(G410));

  xor2  gate2521(.a(G338), .b(G21), .O(gate90inter0));
  nand2 gate2522(.a(gate90inter0), .b(s_282), .O(gate90inter1));
  and2  gate2523(.a(G338), .b(G21), .O(gate90inter2));
  inv1  gate2524(.a(s_282), .O(gate90inter3));
  inv1  gate2525(.a(s_283), .O(gate90inter4));
  nand2 gate2526(.a(gate90inter4), .b(gate90inter3), .O(gate90inter5));
  nor2  gate2527(.a(gate90inter5), .b(gate90inter2), .O(gate90inter6));
  inv1  gate2528(.a(G21), .O(gate90inter7));
  inv1  gate2529(.a(G338), .O(gate90inter8));
  nand2 gate2530(.a(gate90inter8), .b(gate90inter7), .O(gate90inter9));
  nand2 gate2531(.a(s_283), .b(gate90inter3), .O(gate90inter10));
  nor2  gate2532(.a(gate90inter10), .b(gate90inter9), .O(gate90inter11));
  nor2  gate2533(.a(gate90inter11), .b(gate90inter6), .O(gate90inter12));
  nand2 gate2534(.a(gate90inter12), .b(gate90inter1), .O(G411));
nand2 gate91( .a(G25), .b(G341), .O(G412) );
nand2 gate92( .a(G29), .b(G341), .O(G413) );

  xor2  gate1821(.a(G344), .b(G18), .O(gate93inter0));
  nand2 gate1822(.a(gate93inter0), .b(s_182), .O(gate93inter1));
  and2  gate1823(.a(G344), .b(G18), .O(gate93inter2));
  inv1  gate1824(.a(s_182), .O(gate93inter3));
  inv1  gate1825(.a(s_183), .O(gate93inter4));
  nand2 gate1826(.a(gate93inter4), .b(gate93inter3), .O(gate93inter5));
  nor2  gate1827(.a(gate93inter5), .b(gate93inter2), .O(gate93inter6));
  inv1  gate1828(.a(G18), .O(gate93inter7));
  inv1  gate1829(.a(G344), .O(gate93inter8));
  nand2 gate1830(.a(gate93inter8), .b(gate93inter7), .O(gate93inter9));
  nand2 gate1831(.a(s_183), .b(gate93inter3), .O(gate93inter10));
  nor2  gate1832(.a(gate93inter10), .b(gate93inter9), .O(gate93inter11));
  nor2  gate1833(.a(gate93inter11), .b(gate93inter6), .O(gate93inter12));
  nand2 gate1834(.a(gate93inter12), .b(gate93inter1), .O(G414));
nand2 gate94( .a(G22), .b(G344), .O(G415) );
nand2 gate95( .a(G26), .b(G347), .O(G416) );

  xor2  gate1331(.a(G347), .b(G30), .O(gate96inter0));
  nand2 gate1332(.a(gate96inter0), .b(s_112), .O(gate96inter1));
  and2  gate1333(.a(G347), .b(G30), .O(gate96inter2));
  inv1  gate1334(.a(s_112), .O(gate96inter3));
  inv1  gate1335(.a(s_113), .O(gate96inter4));
  nand2 gate1336(.a(gate96inter4), .b(gate96inter3), .O(gate96inter5));
  nor2  gate1337(.a(gate96inter5), .b(gate96inter2), .O(gate96inter6));
  inv1  gate1338(.a(G30), .O(gate96inter7));
  inv1  gate1339(.a(G347), .O(gate96inter8));
  nand2 gate1340(.a(gate96inter8), .b(gate96inter7), .O(gate96inter9));
  nand2 gate1341(.a(s_113), .b(gate96inter3), .O(gate96inter10));
  nor2  gate1342(.a(gate96inter10), .b(gate96inter9), .O(gate96inter11));
  nor2  gate1343(.a(gate96inter11), .b(gate96inter6), .O(gate96inter12));
  nand2 gate1344(.a(gate96inter12), .b(gate96inter1), .O(G417));
nand2 gate97( .a(G19), .b(G350), .O(G418) );

  xor2  gate1849(.a(G350), .b(G23), .O(gate98inter0));
  nand2 gate1850(.a(gate98inter0), .b(s_186), .O(gate98inter1));
  and2  gate1851(.a(G350), .b(G23), .O(gate98inter2));
  inv1  gate1852(.a(s_186), .O(gate98inter3));
  inv1  gate1853(.a(s_187), .O(gate98inter4));
  nand2 gate1854(.a(gate98inter4), .b(gate98inter3), .O(gate98inter5));
  nor2  gate1855(.a(gate98inter5), .b(gate98inter2), .O(gate98inter6));
  inv1  gate1856(.a(G23), .O(gate98inter7));
  inv1  gate1857(.a(G350), .O(gate98inter8));
  nand2 gate1858(.a(gate98inter8), .b(gate98inter7), .O(gate98inter9));
  nand2 gate1859(.a(s_187), .b(gate98inter3), .O(gate98inter10));
  nor2  gate1860(.a(gate98inter10), .b(gate98inter9), .O(gate98inter11));
  nor2  gate1861(.a(gate98inter11), .b(gate98inter6), .O(gate98inter12));
  nand2 gate1862(.a(gate98inter12), .b(gate98inter1), .O(G419));
nand2 gate99( .a(G27), .b(G353), .O(G420) );

  xor2  gate1205(.a(G353), .b(G31), .O(gate100inter0));
  nand2 gate1206(.a(gate100inter0), .b(s_94), .O(gate100inter1));
  and2  gate1207(.a(G353), .b(G31), .O(gate100inter2));
  inv1  gate1208(.a(s_94), .O(gate100inter3));
  inv1  gate1209(.a(s_95), .O(gate100inter4));
  nand2 gate1210(.a(gate100inter4), .b(gate100inter3), .O(gate100inter5));
  nor2  gate1211(.a(gate100inter5), .b(gate100inter2), .O(gate100inter6));
  inv1  gate1212(.a(G31), .O(gate100inter7));
  inv1  gate1213(.a(G353), .O(gate100inter8));
  nand2 gate1214(.a(gate100inter8), .b(gate100inter7), .O(gate100inter9));
  nand2 gate1215(.a(s_95), .b(gate100inter3), .O(gate100inter10));
  nor2  gate1216(.a(gate100inter10), .b(gate100inter9), .O(gate100inter11));
  nor2  gate1217(.a(gate100inter11), .b(gate100inter6), .O(gate100inter12));
  nand2 gate1218(.a(gate100inter12), .b(gate100inter1), .O(G421));
nand2 gate101( .a(G20), .b(G356), .O(G422) );

  xor2  gate2591(.a(G356), .b(G24), .O(gate102inter0));
  nand2 gate2592(.a(gate102inter0), .b(s_292), .O(gate102inter1));
  and2  gate2593(.a(G356), .b(G24), .O(gate102inter2));
  inv1  gate2594(.a(s_292), .O(gate102inter3));
  inv1  gate2595(.a(s_293), .O(gate102inter4));
  nand2 gate2596(.a(gate102inter4), .b(gate102inter3), .O(gate102inter5));
  nor2  gate2597(.a(gate102inter5), .b(gate102inter2), .O(gate102inter6));
  inv1  gate2598(.a(G24), .O(gate102inter7));
  inv1  gate2599(.a(G356), .O(gate102inter8));
  nand2 gate2600(.a(gate102inter8), .b(gate102inter7), .O(gate102inter9));
  nand2 gate2601(.a(s_293), .b(gate102inter3), .O(gate102inter10));
  nor2  gate2602(.a(gate102inter10), .b(gate102inter9), .O(gate102inter11));
  nor2  gate2603(.a(gate102inter11), .b(gate102inter6), .O(gate102inter12));
  nand2 gate2604(.a(gate102inter12), .b(gate102inter1), .O(G423));
nand2 gate103( .a(G28), .b(G359), .O(G424) );
nand2 gate104( .a(G32), .b(G359), .O(G425) );
nand2 gate105( .a(G362), .b(G363), .O(G426) );

  xor2  gate2339(.a(G365), .b(G364), .O(gate106inter0));
  nand2 gate2340(.a(gate106inter0), .b(s_256), .O(gate106inter1));
  and2  gate2341(.a(G365), .b(G364), .O(gate106inter2));
  inv1  gate2342(.a(s_256), .O(gate106inter3));
  inv1  gate2343(.a(s_257), .O(gate106inter4));
  nand2 gate2344(.a(gate106inter4), .b(gate106inter3), .O(gate106inter5));
  nor2  gate2345(.a(gate106inter5), .b(gate106inter2), .O(gate106inter6));
  inv1  gate2346(.a(G364), .O(gate106inter7));
  inv1  gate2347(.a(G365), .O(gate106inter8));
  nand2 gate2348(.a(gate106inter8), .b(gate106inter7), .O(gate106inter9));
  nand2 gate2349(.a(s_257), .b(gate106inter3), .O(gate106inter10));
  nor2  gate2350(.a(gate106inter10), .b(gate106inter9), .O(gate106inter11));
  nor2  gate2351(.a(gate106inter11), .b(gate106inter6), .O(gate106inter12));
  nand2 gate2352(.a(gate106inter12), .b(gate106inter1), .O(G429));
nand2 gate107( .a(G366), .b(G367), .O(G432) );
nand2 gate108( .a(G368), .b(G369), .O(G435) );

  xor2  gate939(.a(G371), .b(G370), .O(gate109inter0));
  nand2 gate940(.a(gate109inter0), .b(s_56), .O(gate109inter1));
  and2  gate941(.a(G371), .b(G370), .O(gate109inter2));
  inv1  gate942(.a(s_56), .O(gate109inter3));
  inv1  gate943(.a(s_57), .O(gate109inter4));
  nand2 gate944(.a(gate109inter4), .b(gate109inter3), .O(gate109inter5));
  nor2  gate945(.a(gate109inter5), .b(gate109inter2), .O(gate109inter6));
  inv1  gate946(.a(G370), .O(gate109inter7));
  inv1  gate947(.a(G371), .O(gate109inter8));
  nand2 gate948(.a(gate109inter8), .b(gate109inter7), .O(gate109inter9));
  nand2 gate949(.a(s_57), .b(gate109inter3), .O(gate109inter10));
  nor2  gate950(.a(gate109inter10), .b(gate109inter9), .O(gate109inter11));
  nor2  gate951(.a(gate109inter11), .b(gate109inter6), .O(gate109inter12));
  nand2 gate952(.a(gate109inter12), .b(gate109inter1), .O(G438));
nand2 gate110( .a(G372), .b(G373), .O(G441) );

  xor2  gate1261(.a(G375), .b(G374), .O(gate111inter0));
  nand2 gate1262(.a(gate111inter0), .b(s_102), .O(gate111inter1));
  and2  gate1263(.a(G375), .b(G374), .O(gate111inter2));
  inv1  gate1264(.a(s_102), .O(gate111inter3));
  inv1  gate1265(.a(s_103), .O(gate111inter4));
  nand2 gate1266(.a(gate111inter4), .b(gate111inter3), .O(gate111inter5));
  nor2  gate1267(.a(gate111inter5), .b(gate111inter2), .O(gate111inter6));
  inv1  gate1268(.a(G374), .O(gate111inter7));
  inv1  gate1269(.a(G375), .O(gate111inter8));
  nand2 gate1270(.a(gate111inter8), .b(gate111inter7), .O(gate111inter9));
  nand2 gate1271(.a(s_103), .b(gate111inter3), .O(gate111inter10));
  nor2  gate1272(.a(gate111inter10), .b(gate111inter9), .O(gate111inter11));
  nor2  gate1273(.a(gate111inter11), .b(gate111inter6), .O(gate111inter12));
  nand2 gate1274(.a(gate111inter12), .b(gate111inter1), .O(G444));
nand2 gate112( .a(G376), .b(G377), .O(G447) );

  xor2  gate1527(.a(G379), .b(G378), .O(gate113inter0));
  nand2 gate1528(.a(gate113inter0), .b(s_140), .O(gate113inter1));
  and2  gate1529(.a(G379), .b(G378), .O(gate113inter2));
  inv1  gate1530(.a(s_140), .O(gate113inter3));
  inv1  gate1531(.a(s_141), .O(gate113inter4));
  nand2 gate1532(.a(gate113inter4), .b(gate113inter3), .O(gate113inter5));
  nor2  gate1533(.a(gate113inter5), .b(gate113inter2), .O(gate113inter6));
  inv1  gate1534(.a(G378), .O(gate113inter7));
  inv1  gate1535(.a(G379), .O(gate113inter8));
  nand2 gate1536(.a(gate113inter8), .b(gate113inter7), .O(gate113inter9));
  nand2 gate1537(.a(s_141), .b(gate113inter3), .O(gate113inter10));
  nor2  gate1538(.a(gate113inter10), .b(gate113inter9), .O(gate113inter11));
  nor2  gate1539(.a(gate113inter11), .b(gate113inter6), .O(gate113inter12));
  nand2 gate1540(.a(gate113inter12), .b(gate113inter1), .O(G450));
nand2 gate114( .a(G380), .b(G381), .O(G453) );
nand2 gate115( .a(G382), .b(G383), .O(G456) );
nand2 gate116( .a(G384), .b(G385), .O(G459) );
nand2 gate117( .a(G386), .b(G387), .O(G462) );

  xor2  gate1583(.a(G389), .b(G388), .O(gate118inter0));
  nand2 gate1584(.a(gate118inter0), .b(s_148), .O(gate118inter1));
  and2  gate1585(.a(G389), .b(G388), .O(gate118inter2));
  inv1  gate1586(.a(s_148), .O(gate118inter3));
  inv1  gate1587(.a(s_149), .O(gate118inter4));
  nand2 gate1588(.a(gate118inter4), .b(gate118inter3), .O(gate118inter5));
  nor2  gate1589(.a(gate118inter5), .b(gate118inter2), .O(gate118inter6));
  inv1  gate1590(.a(G388), .O(gate118inter7));
  inv1  gate1591(.a(G389), .O(gate118inter8));
  nand2 gate1592(.a(gate118inter8), .b(gate118inter7), .O(gate118inter9));
  nand2 gate1593(.a(s_149), .b(gate118inter3), .O(gate118inter10));
  nor2  gate1594(.a(gate118inter10), .b(gate118inter9), .O(gate118inter11));
  nor2  gate1595(.a(gate118inter11), .b(gate118inter6), .O(gate118inter12));
  nand2 gate1596(.a(gate118inter12), .b(gate118inter1), .O(G465));

  xor2  gate701(.a(G391), .b(G390), .O(gate119inter0));
  nand2 gate702(.a(gate119inter0), .b(s_22), .O(gate119inter1));
  and2  gate703(.a(G391), .b(G390), .O(gate119inter2));
  inv1  gate704(.a(s_22), .O(gate119inter3));
  inv1  gate705(.a(s_23), .O(gate119inter4));
  nand2 gate706(.a(gate119inter4), .b(gate119inter3), .O(gate119inter5));
  nor2  gate707(.a(gate119inter5), .b(gate119inter2), .O(gate119inter6));
  inv1  gate708(.a(G390), .O(gate119inter7));
  inv1  gate709(.a(G391), .O(gate119inter8));
  nand2 gate710(.a(gate119inter8), .b(gate119inter7), .O(gate119inter9));
  nand2 gate711(.a(s_23), .b(gate119inter3), .O(gate119inter10));
  nor2  gate712(.a(gate119inter10), .b(gate119inter9), .O(gate119inter11));
  nor2  gate713(.a(gate119inter11), .b(gate119inter6), .O(gate119inter12));
  nand2 gate714(.a(gate119inter12), .b(gate119inter1), .O(G468));
nand2 gate120( .a(G392), .b(G393), .O(G471) );
nand2 gate121( .a(G394), .b(G395), .O(G474) );
nand2 gate122( .a(G396), .b(G397), .O(G477) );

  xor2  gate2423(.a(G399), .b(G398), .O(gate123inter0));
  nand2 gate2424(.a(gate123inter0), .b(s_268), .O(gate123inter1));
  and2  gate2425(.a(G399), .b(G398), .O(gate123inter2));
  inv1  gate2426(.a(s_268), .O(gate123inter3));
  inv1  gate2427(.a(s_269), .O(gate123inter4));
  nand2 gate2428(.a(gate123inter4), .b(gate123inter3), .O(gate123inter5));
  nor2  gate2429(.a(gate123inter5), .b(gate123inter2), .O(gate123inter6));
  inv1  gate2430(.a(G398), .O(gate123inter7));
  inv1  gate2431(.a(G399), .O(gate123inter8));
  nand2 gate2432(.a(gate123inter8), .b(gate123inter7), .O(gate123inter9));
  nand2 gate2433(.a(s_269), .b(gate123inter3), .O(gate123inter10));
  nor2  gate2434(.a(gate123inter10), .b(gate123inter9), .O(gate123inter11));
  nor2  gate2435(.a(gate123inter11), .b(gate123inter6), .O(gate123inter12));
  nand2 gate2436(.a(gate123inter12), .b(gate123inter1), .O(G480));
nand2 gate124( .a(G400), .b(G401), .O(G483) );
nand2 gate125( .a(G402), .b(G403), .O(G486) );
nand2 gate126( .a(G404), .b(G405), .O(G489) );

  xor2  gate2395(.a(G407), .b(G406), .O(gate127inter0));
  nand2 gate2396(.a(gate127inter0), .b(s_264), .O(gate127inter1));
  and2  gate2397(.a(G407), .b(G406), .O(gate127inter2));
  inv1  gate2398(.a(s_264), .O(gate127inter3));
  inv1  gate2399(.a(s_265), .O(gate127inter4));
  nand2 gate2400(.a(gate127inter4), .b(gate127inter3), .O(gate127inter5));
  nor2  gate2401(.a(gate127inter5), .b(gate127inter2), .O(gate127inter6));
  inv1  gate2402(.a(G406), .O(gate127inter7));
  inv1  gate2403(.a(G407), .O(gate127inter8));
  nand2 gate2404(.a(gate127inter8), .b(gate127inter7), .O(gate127inter9));
  nand2 gate2405(.a(s_265), .b(gate127inter3), .O(gate127inter10));
  nor2  gate2406(.a(gate127inter10), .b(gate127inter9), .O(gate127inter11));
  nor2  gate2407(.a(gate127inter11), .b(gate127inter6), .O(gate127inter12));
  nand2 gate2408(.a(gate127inter12), .b(gate127inter1), .O(G492));
nand2 gate128( .a(G408), .b(G409), .O(G495) );

  xor2  gate1387(.a(G411), .b(G410), .O(gate129inter0));
  nand2 gate1388(.a(gate129inter0), .b(s_120), .O(gate129inter1));
  and2  gate1389(.a(G411), .b(G410), .O(gate129inter2));
  inv1  gate1390(.a(s_120), .O(gate129inter3));
  inv1  gate1391(.a(s_121), .O(gate129inter4));
  nand2 gate1392(.a(gate129inter4), .b(gate129inter3), .O(gate129inter5));
  nor2  gate1393(.a(gate129inter5), .b(gate129inter2), .O(gate129inter6));
  inv1  gate1394(.a(G410), .O(gate129inter7));
  inv1  gate1395(.a(G411), .O(gate129inter8));
  nand2 gate1396(.a(gate129inter8), .b(gate129inter7), .O(gate129inter9));
  nand2 gate1397(.a(s_121), .b(gate129inter3), .O(gate129inter10));
  nor2  gate1398(.a(gate129inter10), .b(gate129inter9), .O(gate129inter11));
  nor2  gate1399(.a(gate129inter11), .b(gate129inter6), .O(gate129inter12));
  nand2 gate1400(.a(gate129inter12), .b(gate129inter1), .O(G498));
nand2 gate130( .a(G412), .b(G413), .O(G501) );
nand2 gate131( .a(G414), .b(G415), .O(G504) );
nand2 gate132( .a(G416), .b(G417), .O(G507) );

  xor2  gate1947(.a(G419), .b(G418), .O(gate133inter0));
  nand2 gate1948(.a(gate133inter0), .b(s_200), .O(gate133inter1));
  and2  gate1949(.a(G419), .b(G418), .O(gate133inter2));
  inv1  gate1950(.a(s_200), .O(gate133inter3));
  inv1  gate1951(.a(s_201), .O(gate133inter4));
  nand2 gate1952(.a(gate133inter4), .b(gate133inter3), .O(gate133inter5));
  nor2  gate1953(.a(gate133inter5), .b(gate133inter2), .O(gate133inter6));
  inv1  gate1954(.a(G418), .O(gate133inter7));
  inv1  gate1955(.a(G419), .O(gate133inter8));
  nand2 gate1956(.a(gate133inter8), .b(gate133inter7), .O(gate133inter9));
  nand2 gate1957(.a(s_201), .b(gate133inter3), .O(gate133inter10));
  nor2  gate1958(.a(gate133inter10), .b(gate133inter9), .O(gate133inter11));
  nor2  gate1959(.a(gate133inter11), .b(gate133inter6), .O(gate133inter12));
  nand2 gate1960(.a(gate133inter12), .b(gate133inter1), .O(G510));
nand2 gate134( .a(G420), .b(G421), .O(G513) );
nand2 gate135( .a(G422), .b(G423), .O(G516) );
nand2 gate136( .a(G424), .b(G425), .O(G519) );

  xor2  gate2087(.a(G429), .b(G426), .O(gate137inter0));
  nand2 gate2088(.a(gate137inter0), .b(s_220), .O(gate137inter1));
  and2  gate2089(.a(G429), .b(G426), .O(gate137inter2));
  inv1  gate2090(.a(s_220), .O(gate137inter3));
  inv1  gate2091(.a(s_221), .O(gate137inter4));
  nand2 gate2092(.a(gate137inter4), .b(gate137inter3), .O(gate137inter5));
  nor2  gate2093(.a(gate137inter5), .b(gate137inter2), .O(gate137inter6));
  inv1  gate2094(.a(G426), .O(gate137inter7));
  inv1  gate2095(.a(G429), .O(gate137inter8));
  nand2 gate2096(.a(gate137inter8), .b(gate137inter7), .O(gate137inter9));
  nand2 gate2097(.a(s_221), .b(gate137inter3), .O(gate137inter10));
  nor2  gate2098(.a(gate137inter10), .b(gate137inter9), .O(gate137inter11));
  nor2  gate2099(.a(gate137inter11), .b(gate137inter6), .O(gate137inter12));
  nand2 gate2100(.a(gate137inter12), .b(gate137inter1), .O(G522));
nand2 gate138( .a(G432), .b(G435), .O(G525) );
nand2 gate139( .a(G438), .b(G441), .O(G528) );
nand2 gate140( .a(G444), .b(G447), .O(G531) );
nand2 gate141( .a(G450), .b(G453), .O(G534) );
nand2 gate142( .a(G456), .b(G459), .O(G537) );

  xor2  gate1779(.a(G465), .b(G462), .O(gate143inter0));
  nand2 gate1780(.a(gate143inter0), .b(s_176), .O(gate143inter1));
  and2  gate1781(.a(G465), .b(G462), .O(gate143inter2));
  inv1  gate1782(.a(s_176), .O(gate143inter3));
  inv1  gate1783(.a(s_177), .O(gate143inter4));
  nand2 gate1784(.a(gate143inter4), .b(gate143inter3), .O(gate143inter5));
  nor2  gate1785(.a(gate143inter5), .b(gate143inter2), .O(gate143inter6));
  inv1  gate1786(.a(G462), .O(gate143inter7));
  inv1  gate1787(.a(G465), .O(gate143inter8));
  nand2 gate1788(.a(gate143inter8), .b(gate143inter7), .O(gate143inter9));
  nand2 gate1789(.a(s_177), .b(gate143inter3), .O(gate143inter10));
  nor2  gate1790(.a(gate143inter10), .b(gate143inter9), .O(gate143inter11));
  nor2  gate1791(.a(gate143inter11), .b(gate143inter6), .O(gate143inter12));
  nand2 gate1792(.a(gate143inter12), .b(gate143inter1), .O(G540));

  xor2  gate995(.a(G471), .b(G468), .O(gate144inter0));
  nand2 gate996(.a(gate144inter0), .b(s_64), .O(gate144inter1));
  and2  gate997(.a(G471), .b(G468), .O(gate144inter2));
  inv1  gate998(.a(s_64), .O(gate144inter3));
  inv1  gate999(.a(s_65), .O(gate144inter4));
  nand2 gate1000(.a(gate144inter4), .b(gate144inter3), .O(gate144inter5));
  nor2  gate1001(.a(gate144inter5), .b(gate144inter2), .O(gate144inter6));
  inv1  gate1002(.a(G468), .O(gate144inter7));
  inv1  gate1003(.a(G471), .O(gate144inter8));
  nand2 gate1004(.a(gate144inter8), .b(gate144inter7), .O(gate144inter9));
  nand2 gate1005(.a(s_65), .b(gate144inter3), .O(gate144inter10));
  nor2  gate1006(.a(gate144inter10), .b(gate144inter9), .O(gate144inter11));
  nor2  gate1007(.a(gate144inter11), .b(gate144inter6), .O(gate144inter12));
  nand2 gate1008(.a(gate144inter12), .b(gate144inter1), .O(G543));
nand2 gate145( .a(G474), .b(G477), .O(G546) );
nand2 gate146( .a(G480), .b(G483), .O(G549) );
nand2 gate147( .a(G486), .b(G489), .O(G552) );
nand2 gate148( .a(G492), .b(G495), .O(G555) );

  xor2  gate1835(.a(G501), .b(G498), .O(gate149inter0));
  nand2 gate1836(.a(gate149inter0), .b(s_184), .O(gate149inter1));
  and2  gate1837(.a(G501), .b(G498), .O(gate149inter2));
  inv1  gate1838(.a(s_184), .O(gate149inter3));
  inv1  gate1839(.a(s_185), .O(gate149inter4));
  nand2 gate1840(.a(gate149inter4), .b(gate149inter3), .O(gate149inter5));
  nor2  gate1841(.a(gate149inter5), .b(gate149inter2), .O(gate149inter6));
  inv1  gate1842(.a(G498), .O(gate149inter7));
  inv1  gate1843(.a(G501), .O(gate149inter8));
  nand2 gate1844(.a(gate149inter8), .b(gate149inter7), .O(gate149inter9));
  nand2 gate1845(.a(s_185), .b(gate149inter3), .O(gate149inter10));
  nor2  gate1846(.a(gate149inter10), .b(gate149inter9), .O(gate149inter11));
  nor2  gate1847(.a(gate149inter11), .b(gate149inter6), .O(gate149inter12));
  nand2 gate1848(.a(gate149inter12), .b(gate149inter1), .O(G558));
nand2 gate150( .a(G504), .b(G507), .O(G561) );

  xor2  gate2115(.a(G513), .b(G510), .O(gate151inter0));
  nand2 gate2116(.a(gate151inter0), .b(s_224), .O(gate151inter1));
  and2  gate2117(.a(G513), .b(G510), .O(gate151inter2));
  inv1  gate2118(.a(s_224), .O(gate151inter3));
  inv1  gate2119(.a(s_225), .O(gate151inter4));
  nand2 gate2120(.a(gate151inter4), .b(gate151inter3), .O(gate151inter5));
  nor2  gate2121(.a(gate151inter5), .b(gate151inter2), .O(gate151inter6));
  inv1  gate2122(.a(G510), .O(gate151inter7));
  inv1  gate2123(.a(G513), .O(gate151inter8));
  nand2 gate2124(.a(gate151inter8), .b(gate151inter7), .O(gate151inter9));
  nand2 gate2125(.a(s_225), .b(gate151inter3), .O(gate151inter10));
  nor2  gate2126(.a(gate151inter10), .b(gate151inter9), .O(gate151inter11));
  nor2  gate2127(.a(gate151inter11), .b(gate151inter6), .O(gate151inter12));
  nand2 gate2128(.a(gate151inter12), .b(gate151inter1), .O(G564));
nand2 gate152( .a(G516), .b(G519), .O(G567) );
nand2 gate153( .a(G426), .b(G522), .O(G570) );
nand2 gate154( .a(G429), .b(G522), .O(G571) );
nand2 gate155( .a(G432), .b(G525), .O(G572) );
nand2 gate156( .a(G435), .b(G525), .O(G573) );

  xor2  gate645(.a(G528), .b(G438), .O(gate157inter0));
  nand2 gate646(.a(gate157inter0), .b(s_14), .O(gate157inter1));
  and2  gate647(.a(G528), .b(G438), .O(gate157inter2));
  inv1  gate648(.a(s_14), .O(gate157inter3));
  inv1  gate649(.a(s_15), .O(gate157inter4));
  nand2 gate650(.a(gate157inter4), .b(gate157inter3), .O(gate157inter5));
  nor2  gate651(.a(gate157inter5), .b(gate157inter2), .O(gate157inter6));
  inv1  gate652(.a(G438), .O(gate157inter7));
  inv1  gate653(.a(G528), .O(gate157inter8));
  nand2 gate654(.a(gate157inter8), .b(gate157inter7), .O(gate157inter9));
  nand2 gate655(.a(s_15), .b(gate157inter3), .O(gate157inter10));
  nor2  gate656(.a(gate157inter10), .b(gate157inter9), .O(gate157inter11));
  nor2  gate657(.a(gate157inter11), .b(gate157inter6), .O(gate157inter12));
  nand2 gate658(.a(gate157inter12), .b(gate157inter1), .O(G574));
nand2 gate158( .a(G441), .b(G528), .O(G575) );
nand2 gate159( .a(G444), .b(G531), .O(G576) );
nand2 gate160( .a(G447), .b(G531), .O(G577) );
nand2 gate161( .a(G450), .b(G534), .O(G578) );

  xor2  gate2549(.a(G534), .b(G453), .O(gate162inter0));
  nand2 gate2550(.a(gate162inter0), .b(s_286), .O(gate162inter1));
  and2  gate2551(.a(G534), .b(G453), .O(gate162inter2));
  inv1  gate2552(.a(s_286), .O(gate162inter3));
  inv1  gate2553(.a(s_287), .O(gate162inter4));
  nand2 gate2554(.a(gate162inter4), .b(gate162inter3), .O(gate162inter5));
  nor2  gate2555(.a(gate162inter5), .b(gate162inter2), .O(gate162inter6));
  inv1  gate2556(.a(G453), .O(gate162inter7));
  inv1  gate2557(.a(G534), .O(gate162inter8));
  nand2 gate2558(.a(gate162inter8), .b(gate162inter7), .O(gate162inter9));
  nand2 gate2559(.a(s_287), .b(gate162inter3), .O(gate162inter10));
  nor2  gate2560(.a(gate162inter10), .b(gate162inter9), .O(gate162inter11));
  nor2  gate2561(.a(gate162inter11), .b(gate162inter6), .O(gate162inter12));
  nand2 gate2562(.a(gate162inter12), .b(gate162inter1), .O(G579));

  xor2  gate925(.a(G537), .b(G456), .O(gate163inter0));
  nand2 gate926(.a(gate163inter0), .b(s_54), .O(gate163inter1));
  and2  gate927(.a(G537), .b(G456), .O(gate163inter2));
  inv1  gate928(.a(s_54), .O(gate163inter3));
  inv1  gate929(.a(s_55), .O(gate163inter4));
  nand2 gate930(.a(gate163inter4), .b(gate163inter3), .O(gate163inter5));
  nor2  gate931(.a(gate163inter5), .b(gate163inter2), .O(gate163inter6));
  inv1  gate932(.a(G456), .O(gate163inter7));
  inv1  gate933(.a(G537), .O(gate163inter8));
  nand2 gate934(.a(gate163inter8), .b(gate163inter7), .O(gate163inter9));
  nand2 gate935(.a(s_55), .b(gate163inter3), .O(gate163inter10));
  nor2  gate936(.a(gate163inter10), .b(gate163inter9), .O(gate163inter11));
  nor2  gate937(.a(gate163inter11), .b(gate163inter6), .O(gate163inter12));
  nand2 gate938(.a(gate163inter12), .b(gate163inter1), .O(G580));
nand2 gate164( .a(G459), .b(G537), .O(G581) );

  xor2  gate1513(.a(G540), .b(G462), .O(gate165inter0));
  nand2 gate1514(.a(gate165inter0), .b(s_138), .O(gate165inter1));
  and2  gate1515(.a(G540), .b(G462), .O(gate165inter2));
  inv1  gate1516(.a(s_138), .O(gate165inter3));
  inv1  gate1517(.a(s_139), .O(gate165inter4));
  nand2 gate1518(.a(gate165inter4), .b(gate165inter3), .O(gate165inter5));
  nor2  gate1519(.a(gate165inter5), .b(gate165inter2), .O(gate165inter6));
  inv1  gate1520(.a(G462), .O(gate165inter7));
  inv1  gate1521(.a(G540), .O(gate165inter8));
  nand2 gate1522(.a(gate165inter8), .b(gate165inter7), .O(gate165inter9));
  nand2 gate1523(.a(s_139), .b(gate165inter3), .O(gate165inter10));
  nor2  gate1524(.a(gate165inter10), .b(gate165inter9), .O(gate165inter11));
  nor2  gate1525(.a(gate165inter11), .b(gate165inter6), .O(gate165inter12));
  nand2 gate1526(.a(gate165inter12), .b(gate165inter1), .O(G582));
nand2 gate166( .a(G465), .b(G540), .O(G583) );

  xor2  gate1079(.a(G543), .b(G468), .O(gate167inter0));
  nand2 gate1080(.a(gate167inter0), .b(s_76), .O(gate167inter1));
  and2  gate1081(.a(G543), .b(G468), .O(gate167inter2));
  inv1  gate1082(.a(s_76), .O(gate167inter3));
  inv1  gate1083(.a(s_77), .O(gate167inter4));
  nand2 gate1084(.a(gate167inter4), .b(gate167inter3), .O(gate167inter5));
  nor2  gate1085(.a(gate167inter5), .b(gate167inter2), .O(gate167inter6));
  inv1  gate1086(.a(G468), .O(gate167inter7));
  inv1  gate1087(.a(G543), .O(gate167inter8));
  nand2 gate1088(.a(gate167inter8), .b(gate167inter7), .O(gate167inter9));
  nand2 gate1089(.a(s_77), .b(gate167inter3), .O(gate167inter10));
  nor2  gate1090(.a(gate167inter10), .b(gate167inter9), .O(gate167inter11));
  nor2  gate1091(.a(gate167inter11), .b(gate167inter6), .O(gate167inter12));
  nand2 gate1092(.a(gate167inter12), .b(gate167inter1), .O(G584));
nand2 gate168( .a(G471), .b(G543), .O(G585) );
nand2 gate169( .a(G474), .b(G546), .O(G586) );
nand2 gate170( .a(G477), .b(G546), .O(G587) );

  xor2  gate2353(.a(G549), .b(G480), .O(gate171inter0));
  nand2 gate2354(.a(gate171inter0), .b(s_258), .O(gate171inter1));
  and2  gate2355(.a(G549), .b(G480), .O(gate171inter2));
  inv1  gate2356(.a(s_258), .O(gate171inter3));
  inv1  gate2357(.a(s_259), .O(gate171inter4));
  nand2 gate2358(.a(gate171inter4), .b(gate171inter3), .O(gate171inter5));
  nor2  gate2359(.a(gate171inter5), .b(gate171inter2), .O(gate171inter6));
  inv1  gate2360(.a(G480), .O(gate171inter7));
  inv1  gate2361(.a(G549), .O(gate171inter8));
  nand2 gate2362(.a(gate171inter8), .b(gate171inter7), .O(gate171inter9));
  nand2 gate2363(.a(s_259), .b(gate171inter3), .O(gate171inter10));
  nor2  gate2364(.a(gate171inter10), .b(gate171inter9), .O(gate171inter11));
  nor2  gate2365(.a(gate171inter11), .b(gate171inter6), .O(gate171inter12));
  nand2 gate2366(.a(gate171inter12), .b(gate171inter1), .O(G588));
nand2 gate172( .a(G483), .b(G549), .O(G589) );

  xor2  gate2577(.a(G552), .b(G486), .O(gate173inter0));
  nand2 gate2578(.a(gate173inter0), .b(s_290), .O(gate173inter1));
  and2  gate2579(.a(G552), .b(G486), .O(gate173inter2));
  inv1  gate2580(.a(s_290), .O(gate173inter3));
  inv1  gate2581(.a(s_291), .O(gate173inter4));
  nand2 gate2582(.a(gate173inter4), .b(gate173inter3), .O(gate173inter5));
  nor2  gate2583(.a(gate173inter5), .b(gate173inter2), .O(gate173inter6));
  inv1  gate2584(.a(G486), .O(gate173inter7));
  inv1  gate2585(.a(G552), .O(gate173inter8));
  nand2 gate2586(.a(gate173inter8), .b(gate173inter7), .O(gate173inter9));
  nand2 gate2587(.a(s_291), .b(gate173inter3), .O(gate173inter10));
  nor2  gate2588(.a(gate173inter10), .b(gate173inter9), .O(gate173inter11));
  nor2  gate2589(.a(gate173inter11), .b(gate173inter6), .O(gate173inter12));
  nand2 gate2590(.a(gate173inter12), .b(gate173inter1), .O(G590));
nand2 gate174( .a(G489), .b(G552), .O(G591) );
nand2 gate175( .a(G492), .b(G555), .O(G592) );
nand2 gate176( .a(G495), .b(G555), .O(G593) );
nand2 gate177( .a(G498), .b(G558), .O(G594) );

  xor2  gate1359(.a(G558), .b(G501), .O(gate178inter0));
  nand2 gate1360(.a(gate178inter0), .b(s_116), .O(gate178inter1));
  and2  gate1361(.a(G558), .b(G501), .O(gate178inter2));
  inv1  gate1362(.a(s_116), .O(gate178inter3));
  inv1  gate1363(.a(s_117), .O(gate178inter4));
  nand2 gate1364(.a(gate178inter4), .b(gate178inter3), .O(gate178inter5));
  nor2  gate1365(.a(gate178inter5), .b(gate178inter2), .O(gate178inter6));
  inv1  gate1366(.a(G501), .O(gate178inter7));
  inv1  gate1367(.a(G558), .O(gate178inter8));
  nand2 gate1368(.a(gate178inter8), .b(gate178inter7), .O(gate178inter9));
  nand2 gate1369(.a(s_117), .b(gate178inter3), .O(gate178inter10));
  nor2  gate1370(.a(gate178inter10), .b(gate178inter9), .O(gate178inter11));
  nor2  gate1371(.a(gate178inter11), .b(gate178inter6), .O(gate178inter12));
  nand2 gate1372(.a(gate178inter12), .b(gate178inter1), .O(G595));
nand2 gate179( .a(G504), .b(G561), .O(G596) );
nand2 gate180( .a(G507), .b(G561), .O(G597) );
nand2 gate181( .a(G510), .b(G564), .O(G598) );

  xor2  gate2157(.a(G564), .b(G513), .O(gate182inter0));
  nand2 gate2158(.a(gate182inter0), .b(s_230), .O(gate182inter1));
  and2  gate2159(.a(G564), .b(G513), .O(gate182inter2));
  inv1  gate2160(.a(s_230), .O(gate182inter3));
  inv1  gate2161(.a(s_231), .O(gate182inter4));
  nand2 gate2162(.a(gate182inter4), .b(gate182inter3), .O(gate182inter5));
  nor2  gate2163(.a(gate182inter5), .b(gate182inter2), .O(gate182inter6));
  inv1  gate2164(.a(G513), .O(gate182inter7));
  inv1  gate2165(.a(G564), .O(gate182inter8));
  nand2 gate2166(.a(gate182inter8), .b(gate182inter7), .O(gate182inter9));
  nand2 gate2167(.a(s_231), .b(gate182inter3), .O(gate182inter10));
  nor2  gate2168(.a(gate182inter10), .b(gate182inter9), .O(gate182inter11));
  nor2  gate2169(.a(gate182inter11), .b(gate182inter6), .O(gate182inter12));
  nand2 gate2170(.a(gate182inter12), .b(gate182inter1), .O(G599));
nand2 gate183( .a(G516), .b(G567), .O(G600) );
nand2 gate184( .a(G519), .b(G567), .O(G601) );

  xor2  gate2409(.a(G571), .b(G570), .O(gate185inter0));
  nand2 gate2410(.a(gate185inter0), .b(s_266), .O(gate185inter1));
  and2  gate2411(.a(G571), .b(G570), .O(gate185inter2));
  inv1  gate2412(.a(s_266), .O(gate185inter3));
  inv1  gate2413(.a(s_267), .O(gate185inter4));
  nand2 gate2414(.a(gate185inter4), .b(gate185inter3), .O(gate185inter5));
  nor2  gate2415(.a(gate185inter5), .b(gate185inter2), .O(gate185inter6));
  inv1  gate2416(.a(G570), .O(gate185inter7));
  inv1  gate2417(.a(G571), .O(gate185inter8));
  nand2 gate2418(.a(gate185inter8), .b(gate185inter7), .O(gate185inter9));
  nand2 gate2419(.a(s_267), .b(gate185inter3), .O(gate185inter10));
  nor2  gate2420(.a(gate185inter10), .b(gate185inter9), .O(gate185inter11));
  nor2  gate2421(.a(gate185inter11), .b(gate185inter6), .O(gate185inter12));
  nand2 gate2422(.a(gate185inter12), .b(gate185inter1), .O(G602));

  xor2  gate1933(.a(G573), .b(G572), .O(gate186inter0));
  nand2 gate1934(.a(gate186inter0), .b(s_198), .O(gate186inter1));
  and2  gate1935(.a(G573), .b(G572), .O(gate186inter2));
  inv1  gate1936(.a(s_198), .O(gate186inter3));
  inv1  gate1937(.a(s_199), .O(gate186inter4));
  nand2 gate1938(.a(gate186inter4), .b(gate186inter3), .O(gate186inter5));
  nor2  gate1939(.a(gate186inter5), .b(gate186inter2), .O(gate186inter6));
  inv1  gate1940(.a(G572), .O(gate186inter7));
  inv1  gate1941(.a(G573), .O(gate186inter8));
  nand2 gate1942(.a(gate186inter8), .b(gate186inter7), .O(gate186inter9));
  nand2 gate1943(.a(s_199), .b(gate186inter3), .O(gate186inter10));
  nor2  gate1944(.a(gate186inter10), .b(gate186inter9), .O(gate186inter11));
  nor2  gate1945(.a(gate186inter11), .b(gate186inter6), .O(gate186inter12));
  nand2 gate1946(.a(gate186inter12), .b(gate186inter1), .O(G607));
nand2 gate187( .a(G574), .b(G575), .O(G612) );
nand2 gate188( .a(G576), .b(G577), .O(G617) );

  xor2  gate2661(.a(G579), .b(G578), .O(gate189inter0));
  nand2 gate2662(.a(gate189inter0), .b(s_302), .O(gate189inter1));
  and2  gate2663(.a(G579), .b(G578), .O(gate189inter2));
  inv1  gate2664(.a(s_302), .O(gate189inter3));
  inv1  gate2665(.a(s_303), .O(gate189inter4));
  nand2 gate2666(.a(gate189inter4), .b(gate189inter3), .O(gate189inter5));
  nor2  gate2667(.a(gate189inter5), .b(gate189inter2), .O(gate189inter6));
  inv1  gate2668(.a(G578), .O(gate189inter7));
  inv1  gate2669(.a(G579), .O(gate189inter8));
  nand2 gate2670(.a(gate189inter8), .b(gate189inter7), .O(gate189inter9));
  nand2 gate2671(.a(s_303), .b(gate189inter3), .O(gate189inter10));
  nor2  gate2672(.a(gate189inter10), .b(gate189inter9), .O(gate189inter11));
  nor2  gate2673(.a(gate189inter11), .b(gate189inter6), .O(gate189inter12));
  nand2 gate2674(.a(gate189inter12), .b(gate189inter1), .O(G622));
nand2 gate190( .a(G580), .b(G581), .O(G627) );
nand2 gate191( .a(G582), .b(G583), .O(G632) );
nand2 gate192( .a(G584), .b(G585), .O(G637) );

  xor2  gate2199(.a(G587), .b(G586), .O(gate193inter0));
  nand2 gate2200(.a(gate193inter0), .b(s_236), .O(gate193inter1));
  and2  gate2201(.a(G587), .b(G586), .O(gate193inter2));
  inv1  gate2202(.a(s_236), .O(gate193inter3));
  inv1  gate2203(.a(s_237), .O(gate193inter4));
  nand2 gate2204(.a(gate193inter4), .b(gate193inter3), .O(gate193inter5));
  nor2  gate2205(.a(gate193inter5), .b(gate193inter2), .O(gate193inter6));
  inv1  gate2206(.a(G586), .O(gate193inter7));
  inv1  gate2207(.a(G587), .O(gate193inter8));
  nand2 gate2208(.a(gate193inter8), .b(gate193inter7), .O(gate193inter9));
  nand2 gate2209(.a(s_237), .b(gate193inter3), .O(gate193inter10));
  nor2  gate2210(.a(gate193inter10), .b(gate193inter9), .O(gate193inter11));
  nor2  gate2211(.a(gate193inter11), .b(gate193inter6), .O(gate193inter12));
  nand2 gate2212(.a(gate193inter12), .b(gate193inter1), .O(G642));
nand2 gate194( .a(G588), .b(G589), .O(G645) );

  xor2  gate897(.a(G591), .b(G590), .O(gate195inter0));
  nand2 gate898(.a(gate195inter0), .b(s_50), .O(gate195inter1));
  and2  gate899(.a(G591), .b(G590), .O(gate195inter2));
  inv1  gate900(.a(s_50), .O(gate195inter3));
  inv1  gate901(.a(s_51), .O(gate195inter4));
  nand2 gate902(.a(gate195inter4), .b(gate195inter3), .O(gate195inter5));
  nor2  gate903(.a(gate195inter5), .b(gate195inter2), .O(gate195inter6));
  inv1  gate904(.a(G590), .O(gate195inter7));
  inv1  gate905(.a(G591), .O(gate195inter8));
  nand2 gate906(.a(gate195inter8), .b(gate195inter7), .O(gate195inter9));
  nand2 gate907(.a(s_51), .b(gate195inter3), .O(gate195inter10));
  nor2  gate908(.a(gate195inter10), .b(gate195inter9), .O(gate195inter11));
  nor2  gate909(.a(gate195inter11), .b(gate195inter6), .O(gate195inter12));
  nand2 gate910(.a(gate195inter12), .b(gate195inter1), .O(G648));
nand2 gate196( .a(G592), .b(G593), .O(G651) );
nand2 gate197( .a(G594), .b(G595), .O(G654) );
nand2 gate198( .a(G596), .b(G597), .O(G657) );
nand2 gate199( .a(G598), .b(G599), .O(G660) );
nand2 gate200( .a(G600), .b(G601), .O(G663) );

  xor2  gate981(.a(G607), .b(G602), .O(gate201inter0));
  nand2 gate982(.a(gate201inter0), .b(s_62), .O(gate201inter1));
  and2  gate983(.a(G607), .b(G602), .O(gate201inter2));
  inv1  gate984(.a(s_62), .O(gate201inter3));
  inv1  gate985(.a(s_63), .O(gate201inter4));
  nand2 gate986(.a(gate201inter4), .b(gate201inter3), .O(gate201inter5));
  nor2  gate987(.a(gate201inter5), .b(gate201inter2), .O(gate201inter6));
  inv1  gate988(.a(G602), .O(gate201inter7));
  inv1  gate989(.a(G607), .O(gate201inter8));
  nand2 gate990(.a(gate201inter8), .b(gate201inter7), .O(gate201inter9));
  nand2 gate991(.a(s_63), .b(gate201inter3), .O(gate201inter10));
  nor2  gate992(.a(gate201inter10), .b(gate201inter9), .O(gate201inter11));
  nor2  gate993(.a(gate201inter11), .b(gate201inter6), .O(gate201inter12));
  nand2 gate994(.a(gate201inter12), .b(gate201inter1), .O(G666));
nand2 gate202( .a(G612), .b(G617), .O(G669) );
nand2 gate203( .a(G602), .b(G612), .O(G672) );

  xor2  gate1289(.a(G617), .b(G607), .O(gate204inter0));
  nand2 gate1290(.a(gate204inter0), .b(s_106), .O(gate204inter1));
  and2  gate1291(.a(G617), .b(G607), .O(gate204inter2));
  inv1  gate1292(.a(s_106), .O(gate204inter3));
  inv1  gate1293(.a(s_107), .O(gate204inter4));
  nand2 gate1294(.a(gate204inter4), .b(gate204inter3), .O(gate204inter5));
  nor2  gate1295(.a(gate204inter5), .b(gate204inter2), .O(gate204inter6));
  inv1  gate1296(.a(G607), .O(gate204inter7));
  inv1  gate1297(.a(G617), .O(gate204inter8));
  nand2 gate1298(.a(gate204inter8), .b(gate204inter7), .O(gate204inter9));
  nand2 gate1299(.a(s_107), .b(gate204inter3), .O(gate204inter10));
  nor2  gate1300(.a(gate204inter10), .b(gate204inter9), .O(gate204inter11));
  nor2  gate1301(.a(gate204inter11), .b(gate204inter6), .O(gate204inter12));
  nand2 gate1302(.a(gate204inter12), .b(gate204inter1), .O(G675));

  xor2  gate2493(.a(G627), .b(G622), .O(gate205inter0));
  nand2 gate2494(.a(gate205inter0), .b(s_278), .O(gate205inter1));
  and2  gate2495(.a(G627), .b(G622), .O(gate205inter2));
  inv1  gate2496(.a(s_278), .O(gate205inter3));
  inv1  gate2497(.a(s_279), .O(gate205inter4));
  nand2 gate2498(.a(gate205inter4), .b(gate205inter3), .O(gate205inter5));
  nor2  gate2499(.a(gate205inter5), .b(gate205inter2), .O(gate205inter6));
  inv1  gate2500(.a(G622), .O(gate205inter7));
  inv1  gate2501(.a(G627), .O(gate205inter8));
  nand2 gate2502(.a(gate205inter8), .b(gate205inter7), .O(gate205inter9));
  nand2 gate2503(.a(s_279), .b(gate205inter3), .O(gate205inter10));
  nor2  gate2504(.a(gate205inter10), .b(gate205inter9), .O(gate205inter11));
  nor2  gate2505(.a(gate205inter11), .b(gate205inter6), .O(gate205inter12));
  nand2 gate2506(.a(gate205inter12), .b(gate205inter1), .O(G678));
nand2 gate206( .a(G632), .b(G637), .O(G681) );

  xor2  gate2101(.a(G632), .b(G622), .O(gate207inter0));
  nand2 gate2102(.a(gate207inter0), .b(s_222), .O(gate207inter1));
  and2  gate2103(.a(G632), .b(G622), .O(gate207inter2));
  inv1  gate2104(.a(s_222), .O(gate207inter3));
  inv1  gate2105(.a(s_223), .O(gate207inter4));
  nand2 gate2106(.a(gate207inter4), .b(gate207inter3), .O(gate207inter5));
  nor2  gate2107(.a(gate207inter5), .b(gate207inter2), .O(gate207inter6));
  inv1  gate2108(.a(G622), .O(gate207inter7));
  inv1  gate2109(.a(G632), .O(gate207inter8));
  nand2 gate2110(.a(gate207inter8), .b(gate207inter7), .O(gate207inter9));
  nand2 gate2111(.a(s_223), .b(gate207inter3), .O(gate207inter10));
  nor2  gate2112(.a(gate207inter10), .b(gate207inter9), .O(gate207inter11));
  nor2  gate2113(.a(gate207inter11), .b(gate207inter6), .O(gate207inter12));
  nand2 gate2114(.a(gate207inter12), .b(gate207inter1), .O(G684));

  xor2  gate1499(.a(G637), .b(G627), .O(gate208inter0));
  nand2 gate1500(.a(gate208inter0), .b(s_136), .O(gate208inter1));
  and2  gate1501(.a(G637), .b(G627), .O(gate208inter2));
  inv1  gate1502(.a(s_136), .O(gate208inter3));
  inv1  gate1503(.a(s_137), .O(gate208inter4));
  nand2 gate1504(.a(gate208inter4), .b(gate208inter3), .O(gate208inter5));
  nor2  gate1505(.a(gate208inter5), .b(gate208inter2), .O(gate208inter6));
  inv1  gate1506(.a(G627), .O(gate208inter7));
  inv1  gate1507(.a(G637), .O(gate208inter8));
  nand2 gate1508(.a(gate208inter8), .b(gate208inter7), .O(gate208inter9));
  nand2 gate1509(.a(s_137), .b(gate208inter3), .O(gate208inter10));
  nor2  gate1510(.a(gate208inter10), .b(gate208inter9), .O(gate208inter11));
  nor2  gate1511(.a(gate208inter11), .b(gate208inter6), .O(gate208inter12));
  nand2 gate1512(.a(gate208inter12), .b(gate208inter1), .O(G687));
nand2 gate209( .a(G602), .b(G666), .O(G690) );

  xor2  gate2129(.a(G666), .b(G607), .O(gate210inter0));
  nand2 gate2130(.a(gate210inter0), .b(s_226), .O(gate210inter1));
  and2  gate2131(.a(G666), .b(G607), .O(gate210inter2));
  inv1  gate2132(.a(s_226), .O(gate210inter3));
  inv1  gate2133(.a(s_227), .O(gate210inter4));
  nand2 gate2134(.a(gate210inter4), .b(gate210inter3), .O(gate210inter5));
  nor2  gate2135(.a(gate210inter5), .b(gate210inter2), .O(gate210inter6));
  inv1  gate2136(.a(G607), .O(gate210inter7));
  inv1  gate2137(.a(G666), .O(gate210inter8));
  nand2 gate2138(.a(gate210inter8), .b(gate210inter7), .O(gate210inter9));
  nand2 gate2139(.a(s_227), .b(gate210inter3), .O(gate210inter10));
  nor2  gate2140(.a(gate210inter10), .b(gate210inter9), .O(gate210inter11));
  nor2  gate2141(.a(gate210inter11), .b(gate210inter6), .O(gate210inter12));
  nand2 gate2142(.a(gate210inter12), .b(gate210inter1), .O(G691));
nand2 gate211( .a(G612), .b(G669), .O(G692) );
nand2 gate212( .a(G617), .b(G669), .O(G693) );
nand2 gate213( .a(G602), .b(G672), .O(G694) );
nand2 gate214( .a(G612), .b(G672), .O(G695) );
nand2 gate215( .a(G607), .b(G675), .O(G696) );
nand2 gate216( .a(G617), .b(G675), .O(G697) );
nand2 gate217( .a(G622), .b(G678), .O(G698) );
nand2 gate218( .a(G627), .b(G678), .O(G699) );
nand2 gate219( .a(G632), .b(G681), .O(G700) );

  xor2  gate1975(.a(G681), .b(G637), .O(gate220inter0));
  nand2 gate1976(.a(gate220inter0), .b(s_204), .O(gate220inter1));
  and2  gate1977(.a(G681), .b(G637), .O(gate220inter2));
  inv1  gate1978(.a(s_204), .O(gate220inter3));
  inv1  gate1979(.a(s_205), .O(gate220inter4));
  nand2 gate1980(.a(gate220inter4), .b(gate220inter3), .O(gate220inter5));
  nor2  gate1981(.a(gate220inter5), .b(gate220inter2), .O(gate220inter6));
  inv1  gate1982(.a(G637), .O(gate220inter7));
  inv1  gate1983(.a(G681), .O(gate220inter8));
  nand2 gate1984(.a(gate220inter8), .b(gate220inter7), .O(gate220inter9));
  nand2 gate1985(.a(s_205), .b(gate220inter3), .O(gate220inter10));
  nor2  gate1986(.a(gate220inter10), .b(gate220inter9), .O(gate220inter11));
  nor2  gate1987(.a(gate220inter11), .b(gate220inter6), .O(gate220inter12));
  nand2 gate1988(.a(gate220inter12), .b(gate220inter1), .O(G701));
nand2 gate221( .a(G622), .b(G684), .O(G702) );
nand2 gate222( .a(G632), .b(G684), .O(G703) );
nand2 gate223( .a(G627), .b(G687), .O(G704) );
nand2 gate224( .a(G637), .b(G687), .O(G705) );

  xor2  gate2703(.a(G691), .b(G690), .O(gate225inter0));
  nand2 gate2704(.a(gate225inter0), .b(s_308), .O(gate225inter1));
  and2  gate2705(.a(G691), .b(G690), .O(gate225inter2));
  inv1  gate2706(.a(s_308), .O(gate225inter3));
  inv1  gate2707(.a(s_309), .O(gate225inter4));
  nand2 gate2708(.a(gate225inter4), .b(gate225inter3), .O(gate225inter5));
  nor2  gate2709(.a(gate225inter5), .b(gate225inter2), .O(gate225inter6));
  inv1  gate2710(.a(G690), .O(gate225inter7));
  inv1  gate2711(.a(G691), .O(gate225inter8));
  nand2 gate2712(.a(gate225inter8), .b(gate225inter7), .O(gate225inter9));
  nand2 gate2713(.a(s_309), .b(gate225inter3), .O(gate225inter10));
  nor2  gate2714(.a(gate225inter10), .b(gate225inter9), .O(gate225inter11));
  nor2  gate2715(.a(gate225inter11), .b(gate225inter6), .O(gate225inter12));
  nand2 gate2716(.a(gate225inter12), .b(gate225inter1), .O(G706));

  xor2  gate1919(.a(G693), .b(G692), .O(gate226inter0));
  nand2 gate1920(.a(gate226inter0), .b(s_196), .O(gate226inter1));
  and2  gate1921(.a(G693), .b(G692), .O(gate226inter2));
  inv1  gate1922(.a(s_196), .O(gate226inter3));
  inv1  gate1923(.a(s_197), .O(gate226inter4));
  nand2 gate1924(.a(gate226inter4), .b(gate226inter3), .O(gate226inter5));
  nor2  gate1925(.a(gate226inter5), .b(gate226inter2), .O(gate226inter6));
  inv1  gate1926(.a(G692), .O(gate226inter7));
  inv1  gate1927(.a(G693), .O(gate226inter8));
  nand2 gate1928(.a(gate226inter8), .b(gate226inter7), .O(gate226inter9));
  nand2 gate1929(.a(s_197), .b(gate226inter3), .O(gate226inter10));
  nor2  gate1930(.a(gate226inter10), .b(gate226inter9), .O(gate226inter11));
  nor2  gate1931(.a(gate226inter11), .b(gate226inter6), .O(gate226inter12));
  nand2 gate1932(.a(gate226inter12), .b(gate226inter1), .O(G709));
nand2 gate227( .a(G694), .b(G695), .O(G712) );

  xor2  gate1233(.a(G697), .b(G696), .O(gate228inter0));
  nand2 gate1234(.a(gate228inter0), .b(s_98), .O(gate228inter1));
  and2  gate1235(.a(G697), .b(G696), .O(gate228inter2));
  inv1  gate1236(.a(s_98), .O(gate228inter3));
  inv1  gate1237(.a(s_99), .O(gate228inter4));
  nand2 gate1238(.a(gate228inter4), .b(gate228inter3), .O(gate228inter5));
  nor2  gate1239(.a(gate228inter5), .b(gate228inter2), .O(gate228inter6));
  inv1  gate1240(.a(G696), .O(gate228inter7));
  inv1  gate1241(.a(G697), .O(gate228inter8));
  nand2 gate1242(.a(gate228inter8), .b(gate228inter7), .O(gate228inter9));
  nand2 gate1243(.a(s_99), .b(gate228inter3), .O(gate228inter10));
  nor2  gate1244(.a(gate228inter10), .b(gate228inter9), .O(gate228inter11));
  nor2  gate1245(.a(gate228inter11), .b(gate228inter6), .O(gate228inter12));
  nand2 gate1246(.a(gate228inter12), .b(gate228inter1), .O(G715));
nand2 gate229( .a(G698), .b(G699), .O(G718) );
nand2 gate230( .a(G700), .b(G701), .O(G721) );
nand2 gate231( .a(G702), .b(G703), .O(G724) );
nand2 gate232( .a(G704), .b(G705), .O(G727) );
nand2 gate233( .a(G242), .b(G718), .O(G730) );
nand2 gate234( .a(G245), .b(G721), .O(G733) );

  xor2  gate1051(.a(G724), .b(G248), .O(gate235inter0));
  nand2 gate1052(.a(gate235inter0), .b(s_72), .O(gate235inter1));
  and2  gate1053(.a(G724), .b(G248), .O(gate235inter2));
  inv1  gate1054(.a(s_72), .O(gate235inter3));
  inv1  gate1055(.a(s_73), .O(gate235inter4));
  nand2 gate1056(.a(gate235inter4), .b(gate235inter3), .O(gate235inter5));
  nor2  gate1057(.a(gate235inter5), .b(gate235inter2), .O(gate235inter6));
  inv1  gate1058(.a(G248), .O(gate235inter7));
  inv1  gate1059(.a(G724), .O(gate235inter8));
  nand2 gate1060(.a(gate235inter8), .b(gate235inter7), .O(gate235inter9));
  nand2 gate1061(.a(s_73), .b(gate235inter3), .O(gate235inter10));
  nor2  gate1062(.a(gate235inter10), .b(gate235inter9), .O(gate235inter11));
  nor2  gate1063(.a(gate235inter11), .b(gate235inter6), .O(gate235inter12));
  nand2 gate1064(.a(gate235inter12), .b(gate235inter1), .O(G736));
nand2 gate236( .a(G251), .b(G727), .O(G739) );

  xor2  gate1429(.a(G706), .b(G254), .O(gate237inter0));
  nand2 gate1430(.a(gate237inter0), .b(s_126), .O(gate237inter1));
  and2  gate1431(.a(G706), .b(G254), .O(gate237inter2));
  inv1  gate1432(.a(s_126), .O(gate237inter3));
  inv1  gate1433(.a(s_127), .O(gate237inter4));
  nand2 gate1434(.a(gate237inter4), .b(gate237inter3), .O(gate237inter5));
  nor2  gate1435(.a(gate237inter5), .b(gate237inter2), .O(gate237inter6));
  inv1  gate1436(.a(G254), .O(gate237inter7));
  inv1  gate1437(.a(G706), .O(gate237inter8));
  nand2 gate1438(.a(gate237inter8), .b(gate237inter7), .O(gate237inter9));
  nand2 gate1439(.a(s_127), .b(gate237inter3), .O(gate237inter10));
  nor2  gate1440(.a(gate237inter10), .b(gate237inter9), .O(gate237inter11));
  nor2  gate1441(.a(gate237inter11), .b(gate237inter6), .O(gate237inter12));
  nand2 gate1442(.a(gate237inter12), .b(gate237inter1), .O(G742));
nand2 gate238( .a(G257), .b(G709), .O(G745) );
nand2 gate239( .a(G260), .b(G712), .O(G748) );
nand2 gate240( .a(G263), .b(G715), .O(G751) );

  xor2  gate1877(.a(G730), .b(G242), .O(gate241inter0));
  nand2 gate1878(.a(gate241inter0), .b(s_190), .O(gate241inter1));
  and2  gate1879(.a(G730), .b(G242), .O(gate241inter2));
  inv1  gate1880(.a(s_190), .O(gate241inter3));
  inv1  gate1881(.a(s_191), .O(gate241inter4));
  nand2 gate1882(.a(gate241inter4), .b(gate241inter3), .O(gate241inter5));
  nor2  gate1883(.a(gate241inter5), .b(gate241inter2), .O(gate241inter6));
  inv1  gate1884(.a(G242), .O(gate241inter7));
  inv1  gate1885(.a(G730), .O(gate241inter8));
  nand2 gate1886(.a(gate241inter8), .b(gate241inter7), .O(gate241inter9));
  nand2 gate1887(.a(s_191), .b(gate241inter3), .O(gate241inter10));
  nor2  gate1888(.a(gate241inter10), .b(gate241inter9), .O(gate241inter11));
  nor2  gate1889(.a(gate241inter11), .b(gate241inter6), .O(gate241inter12));
  nand2 gate1890(.a(gate241inter12), .b(gate241inter1), .O(G754));
nand2 gate242( .a(G718), .b(G730), .O(G755) );

  xor2  gate2325(.a(G733), .b(G245), .O(gate243inter0));
  nand2 gate2326(.a(gate243inter0), .b(s_254), .O(gate243inter1));
  and2  gate2327(.a(G733), .b(G245), .O(gate243inter2));
  inv1  gate2328(.a(s_254), .O(gate243inter3));
  inv1  gate2329(.a(s_255), .O(gate243inter4));
  nand2 gate2330(.a(gate243inter4), .b(gate243inter3), .O(gate243inter5));
  nor2  gate2331(.a(gate243inter5), .b(gate243inter2), .O(gate243inter6));
  inv1  gate2332(.a(G245), .O(gate243inter7));
  inv1  gate2333(.a(G733), .O(gate243inter8));
  nand2 gate2334(.a(gate243inter8), .b(gate243inter7), .O(gate243inter9));
  nand2 gate2335(.a(s_255), .b(gate243inter3), .O(gate243inter10));
  nor2  gate2336(.a(gate243inter10), .b(gate243inter9), .O(gate243inter11));
  nor2  gate2337(.a(gate243inter11), .b(gate243inter6), .O(gate243inter12));
  nand2 gate2338(.a(gate243inter12), .b(gate243inter1), .O(G756));

  xor2  gate1989(.a(G733), .b(G721), .O(gate244inter0));
  nand2 gate1990(.a(gate244inter0), .b(s_206), .O(gate244inter1));
  and2  gate1991(.a(G733), .b(G721), .O(gate244inter2));
  inv1  gate1992(.a(s_206), .O(gate244inter3));
  inv1  gate1993(.a(s_207), .O(gate244inter4));
  nand2 gate1994(.a(gate244inter4), .b(gate244inter3), .O(gate244inter5));
  nor2  gate1995(.a(gate244inter5), .b(gate244inter2), .O(gate244inter6));
  inv1  gate1996(.a(G721), .O(gate244inter7));
  inv1  gate1997(.a(G733), .O(gate244inter8));
  nand2 gate1998(.a(gate244inter8), .b(gate244inter7), .O(gate244inter9));
  nand2 gate1999(.a(s_207), .b(gate244inter3), .O(gate244inter10));
  nor2  gate2000(.a(gate244inter10), .b(gate244inter9), .O(gate244inter11));
  nor2  gate2001(.a(gate244inter11), .b(gate244inter6), .O(gate244inter12));
  nand2 gate2002(.a(gate244inter12), .b(gate244inter1), .O(G757));

  xor2  gate2269(.a(G736), .b(G248), .O(gate245inter0));
  nand2 gate2270(.a(gate245inter0), .b(s_246), .O(gate245inter1));
  and2  gate2271(.a(G736), .b(G248), .O(gate245inter2));
  inv1  gate2272(.a(s_246), .O(gate245inter3));
  inv1  gate2273(.a(s_247), .O(gate245inter4));
  nand2 gate2274(.a(gate245inter4), .b(gate245inter3), .O(gate245inter5));
  nor2  gate2275(.a(gate245inter5), .b(gate245inter2), .O(gate245inter6));
  inv1  gate2276(.a(G248), .O(gate245inter7));
  inv1  gate2277(.a(G736), .O(gate245inter8));
  nand2 gate2278(.a(gate245inter8), .b(gate245inter7), .O(gate245inter9));
  nand2 gate2279(.a(s_247), .b(gate245inter3), .O(gate245inter10));
  nor2  gate2280(.a(gate245inter10), .b(gate245inter9), .O(gate245inter11));
  nor2  gate2281(.a(gate245inter11), .b(gate245inter6), .O(gate245inter12));
  nand2 gate2282(.a(gate245inter12), .b(gate245inter1), .O(G758));
nand2 gate246( .a(G724), .b(G736), .O(G759) );
nand2 gate247( .a(G251), .b(G739), .O(G760) );
nand2 gate248( .a(G727), .b(G739), .O(G761) );

  xor2  gate911(.a(G742), .b(G254), .O(gate249inter0));
  nand2 gate912(.a(gate249inter0), .b(s_52), .O(gate249inter1));
  and2  gate913(.a(G742), .b(G254), .O(gate249inter2));
  inv1  gate914(.a(s_52), .O(gate249inter3));
  inv1  gate915(.a(s_53), .O(gate249inter4));
  nand2 gate916(.a(gate249inter4), .b(gate249inter3), .O(gate249inter5));
  nor2  gate917(.a(gate249inter5), .b(gate249inter2), .O(gate249inter6));
  inv1  gate918(.a(G254), .O(gate249inter7));
  inv1  gate919(.a(G742), .O(gate249inter8));
  nand2 gate920(.a(gate249inter8), .b(gate249inter7), .O(gate249inter9));
  nand2 gate921(.a(s_53), .b(gate249inter3), .O(gate249inter10));
  nor2  gate922(.a(gate249inter10), .b(gate249inter9), .O(gate249inter11));
  nor2  gate923(.a(gate249inter11), .b(gate249inter6), .O(gate249inter12));
  nand2 gate924(.a(gate249inter12), .b(gate249inter1), .O(G762));
nand2 gate250( .a(G706), .b(G742), .O(G763) );
nand2 gate251( .a(G257), .b(G745), .O(G764) );

  xor2  gate2633(.a(G745), .b(G709), .O(gate252inter0));
  nand2 gate2634(.a(gate252inter0), .b(s_298), .O(gate252inter1));
  and2  gate2635(.a(G745), .b(G709), .O(gate252inter2));
  inv1  gate2636(.a(s_298), .O(gate252inter3));
  inv1  gate2637(.a(s_299), .O(gate252inter4));
  nand2 gate2638(.a(gate252inter4), .b(gate252inter3), .O(gate252inter5));
  nor2  gate2639(.a(gate252inter5), .b(gate252inter2), .O(gate252inter6));
  inv1  gate2640(.a(G709), .O(gate252inter7));
  inv1  gate2641(.a(G745), .O(gate252inter8));
  nand2 gate2642(.a(gate252inter8), .b(gate252inter7), .O(gate252inter9));
  nand2 gate2643(.a(s_299), .b(gate252inter3), .O(gate252inter10));
  nor2  gate2644(.a(gate252inter10), .b(gate252inter9), .O(gate252inter11));
  nor2  gate2645(.a(gate252inter11), .b(gate252inter6), .O(gate252inter12));
  nand2 gate2646(.a(gate252inter12), .b(gate252inter1), .O(G765));

  xor2  gate729(.a(G748), .b(G260), .O(gate253inter0));
  nand2 gate730(.a(gate253inter0), .b(s_26), .O(gate253inter1));
  and2  gate731(.a(G748), .b(G260), .O(gate253inter2));
  inv1  gate732(.a(s_26), .O(gate253inter3));
  inv1  gate733(.a(s_27), .O(gate253inter4));
  nand2 gate734(.a(gate253inter4), .b(gate253inter3), .O(gate253inter5));
  nor2  gate735(.a(gate253inter5), .b(gate253inter2), .O(gate253inter6));
  inv1  gate736(.a(G260), .O(gate253inter7));
  inv1  gate737(.a(G748), .O(gate253inter8));
  nand2 gate738(.a(gate253inter8), .b(gate253inter7), .O(gate253inter9));
  nand2 gate739(.a(s_27), .b(gate253inter3), .O(gate253inter10));
  nor2  gate740(.a(gate253inter10), .b(gate253inter9), .O(gate253inter11));
  nor2  gate741(.a(gate253inter11), .b(gate253inter6), .O(gate253inter12));
  nand2 gate742(.a(gate253inter12), .b(gate253inter1), .O(G766));

  xor2  gate1737(.a(G748), .b(G712), .O(gate254inter0));
  nand2 gate1738(.a(gate254inter0), .b(s_170), .O(gate254inter1));
  and2  gate1739(.a(G748), .b(G712), .O(gate254inter2));
  inv1  gate1740(.a(s_170), .O(gate254inter3));
  inv1  gate1741(.a(s_171), .O(gate254inter4));
  nand2 gate1742(.a(gate254inter4), .b(gate254inter3), .O(gate254inter5));
  nor2  gate1743(.a(gate254inter5), .b(gate254inter2), .O(gate254inter6));
  inv1  gate1744(.a(G712), .O(gate254inter7));
  inv1  gate1745(.a(G748), .O(gate254inter8));
  nand2 gate1746(.a(gate254inter8), .b(gate254inter7), .O(gate254inter9));
  nand2 gate1747(.a(s_171), .b(gate254inter3), .O(gate254inter10));
  nor2  gate1748(.a(gate254inter10), .b(gate254inter9), .O(gate254inter11));
  nor2  gate1749(.a(gate254inter11), .b(gate254inter6), .O(gate254inter12));
  nand2 gate1750(.a(gate254inter12), .b(gate254inter1), .O(G767));

  xor2  gate1639(.a(G751), .b(G263), .O(gate255inter0));
  nand2 gate1640(.a(gate255inter0), .b(s_156), .O(gate255inter1));
  and2  gate1641(.a(G751), .b(G263), .O(gate255inter2));
  inv1  gate1642(.a(s_156), .O(gate255inter3));
  inv1  gate1643(.a(s_157), .O(gate255inter4));
  nand2 gate1644(.a(gate255inter4), .b(gate255inter3), .O(gate255inter5));
  nor2  gate1645(.a(gate255inter5), .b(gate255inter2), .O(gate255inter6));
  inv1  gate1646(.a(G263), .O(gate255inter7));
  inv1  gate1647(.a(G751), .O(gate255inter8));
  nand2 gate1648(.a(gate255inter8), .b(gate255inter7), .O(gate255inter9));
  nand2 gate1649(.a(s_157), .b(gate255inter3), .O(gate255inter10));
  nor2  gate1650(.a(gate255inter10), .b(gate255inter9), .O(gate255inter11));
  nor2  gate1651(.a(gate255inter11), .b(gate255inter6), .O(gate255inter12));
  nand2 gate1652(.a(gate255inter12), .b(gate255inter1), .O(G768));
nand2 gate256( .a(G715), .b(G751), .O(G769) );

  xor2  gate2465(.a(G755), .b(G754), .O(gate257inter0));
  nand2 gate2466(.a(gate257inter0), .b(s_274), .O(gate257inter1));
  and2  gate2467(.a(G755), .b(G754), .O(gate257inter2));
  inv1  gate2468(.a(s_274), .O(gate257inter3));
  inv1  gate2469(.a(s_275), .O(gate257inter4));
  nand2 gate2470(.a(gate257inter4), .b(gate257inter3), .O(gate257inter5));
  nor2  gate2471(.a(gate257inter5), .b(gate257inter2), .O(gate257inter6));
  inv1  gate2472(.a(G754), .O(gate257inter7));
  inv1  gate2473(.a(G755), .O(gate257inter8));
  nand2 gate2474(.a(gate257inter8), .b(gate257inter7), .O(gate257inter9));
  nand2 gate2475(.a(s_275), .b(gate257inter3), .O(gate257inter10));
  nor2  gate2476(.a(gate257inter10), .b(gate257inter9), .O(gate257inter11));
  nor2  gate2477(.a(gate257inter11), .b(gate257inter6), .O(gate257inter12));
  nand2 gate2478(.a(gate257inter12), .b(gate257inter1), .O(G770));

  xor2  gate1709(.a(G757), .b(G756), .O(gate258inter0));
  nand2 gate1710(.a(gate258inter0), .b(s_166), .O(gate258inter1));
  and2  gate1711(.a(G757), .b(G756), .O(gate258inter2));
  inv1  gate1712(.a(s_166), .O(gate258inter3));
  inv1  gate1713(.a(s_167), .O(gate258inter4));
  nand2 gate1714(.a(gate258inter4), .b(gate258inter3), .O(gate258inter5));
  nor2  gate1715(.a(gate258inter5), .b(gate258inter2), .O(gate258inter6));
  inv1  gate1716(.a(G756), .O(gate258inter7));
  inv1  gate1717(.a(G757), .O(gate258inter8));
  nand2 gate1718(.a(gate258inter8), .b(gate258inter7), .O(gate258inter9));
  nand2 gate1719(.a(s_167), .b(gate258inter3), .O(gate258inter10));
  nor2  gate1720(.a(gate258inter10), .b(gate258inter9), .O(gate258inter11));
  nor2  gate1721(.a(gate258inter11), .b(gate258inter6), .O(gate258inter12));
  nand2 gate1722(.a(gate258inter12), .b(gate258inter1), .O(G773));

  xor2  gate1457(.a(G759), .b(G758), .O(gate259inter0));
  nand2 gate1458(.a(gate259inter0), .b(s_130), .O(gate259inter1));
  and2  gate1459(.a(G759), .b(G758), .O(gate259inter2));
  inv1  gate1460(.a(s_130), .O(gate259inter3));
  inv1  gate1461(.a(s_131), .O(gate259inter4));
  nand2 gate1462(.a(gate259inter4), .b(gate259inter3), .O(gate259inter5));
  nor2  gate1463(.a(gate259inter5), .b(gate259inter2), .O(gate259inter6));
  inv1  gate1464(.a(G758), .O(gate259inter7));
  inv1  gate1465(.a(G759), .O(gate259inter8));
  nand2 gate1466(.a(gate259inter8), .b(gate259inter7), .O(gate259inter9));
  nand2 gate1467(.a(s_131), .b(gate259inter3), .O(gate259inter10));
  nor2  gate1468(.a(gate259inter10), .b(gate259inter9), .O(gate259inter11));
  nor2  gate1469(.a(gate259inter11), .b(gate259inter6), .O(gate259inter12));
  nand2 gate1470(.a(gate259inter12), .b(gate259inter1), .O(G776));
nand2 gate260( .a(G760), .b(G761), .O(G779) );

  xor2  gate1653(.a(G763), .b(G762), .O(gate261inter0));
  nand2 gate1654(.a(gate261inter0), .b(s_158), .O(gate261inter1));
  and2  gate1655(.a(G763), .b(G762), .O(gate261inter2));
  inv1  gate1656(.a(s_158), .O(gate261inter3));
  inv1  gate1657(.a(s_159), .O(gate261inter4));
  nand2 gate1658(.a(gate261inter4), .b(gate261inter3), .O(gate261inter5));
  nor2  gate1659(.a(gate261inter5), .b(gate261inter2), .O(gate261inter6));
  inv1  gate1660(.a(G762), .O(gate261inter7));
  inv1  gate1661(.a(G763), .O(gate261inter8));
  nand2 gate1662(.a(gate261inter8), .b(gate261inter7), .O(gate261inter9));
  nand2 gate1663(.a(s_159), .b(gate261inter3), .O(gate261inter10));
  nor2  gate1664(.a(gate261inter10), .b(gate261inter9), .O(gate261inter11));
  nor2  gate1665(.a(gate261inter11), .b(gate261inter6), .O(gate261inter12));
  nand2 gate1666(.a(gate261inter12), .b(gate261inter1), .O(G782));
nand2 gate262( .a(G764), .b(G765), .O(G785) );

  xor2  gate659(.a(G767), .b(G766), .O(gate263inter0));
  nand2 gate660(.a(gate263inter0), .b(s_16), .O(gate263inter1));
  and2  gate661(.a(G767), .b(G766), .O(gate263inter2));
  inv1  gate662(.a(s_16), .O(gate263inter3));
  inv1  gate663(.a(s_17), .O(gate263inter4));
  nand2 gate664(.a(gate263inter4), .b(gate263inter3), .O(gate263inter5));
  nor2  gate665(.a(gate263inter5), .b(gate263inter2), .O(gate263inter6));
  inv1  gate666(.a(G766), .O(gate263inter7));
  inv1  gate667(.a(G767), .O(gate263inter8));
  nand2 gate668(.a(gate263inter8), .b(gate263inter7), .O(gate263inter9));
  nand2 gate669(.a(s_17), .b(gate263inter3), .O(gate263inter10));
  nor2  gate670(.a(gate263inter10), .b(gate263inter9), .O(gate263inter11));
  nor2  gate671(.a(gate263inter11), .b(gate263inter6), .O(gate263inter12));
  nand2 gate672(.a(gate263inter12), .b(gate263inter1), .O(G788));

  xor2  gate1443(.a(G769), .b(G768), .O(gate264inter0));
  nand2 gate1444(.a(gate264inter0), .b(s_128), .O(gate264inter1));
  and2  gate1445(.a(G769), .b(G768), .O(gate264inter2));
  inv1  gate1446(.a(s_128), .O(gate264inter3));
  inv1  gate1447(.a(s_129), .O(gate264inter4));
  nand2 gate1448(.a(gate264inter4), .b(gate264inter3), .O(gate264inter5));
  nor2  gate1449(.a(gate264inter5), .b(gate264inter2), .O(gate264inter6));
  inv1  gate1450(.a(G768), .O(gate264inter7));
  inv1  gate1451(.a(G769), .O(gate264inter8));
  nand2 gate1452(.a(gate264inter8), .b(gate264inter7), .O(gate264inter9));
  nand2 gate1453(.a(s_129), .b(gate264inter3), .O(gate264inter10));
  nor2  gate1454(.a(gate264inter10), .b(gate264inter9), .O(gate264inter11));
  nor2  gate1455(.a(gate264inter11), .b(gate264inter6), .O(gate264inter12));
  nand2 gate1456(.a(gate264inter12), .b(gate264inter1), .O(G791));

  xor2  gate2073(.a(G770), .b(G642), .O(gate265inter0));
  nand2 gate2074(.a(gate265inter0), .b(s_218), .O(gate265inter1));
  and2  gate2075(.a(G770), .b(G642), .O(gate265inter2));
  inv1  gate2076(.a(s_218), .O(gate265inter3));
  inv1  gate2077(.a(s_219), .O(gate265inter4));
  nand2 gate2078(.a(gate265inter4), .b(gate265inter3), .O(gate265inter5));
  nor2  gate2079(.a(gate265inter5), .b(gate265inter2), .O(gate265inter6));
  inv1  gate2080(.a(G642), .O(gate265inter7));
  inv1  gate2081(.a(G770), .O(gate265inter8));
  nand2 gate2082(.a(gate265inter8), .b(gate265inter7), .O(gate265inter9));
  nand2 gate2083(.a(s_219), .b(gate265inter3), .O(gate265inter10));
  nor2  gate2084(.a(gate265inter10), .b(gate265inter9), .O(gate265inter11));
  nor2  gate2085(.a(gate265inter11), .b(gate265inter6), .O(gate265inter12));
  nand2 gate2086(.a(gate265inter12), .b(gate265inter1), .O(G794));
nand2 gate266( .a(G645), .b(G773), .O(G797) );
nand2 gate267( .a(G648), .b(G776), .O(G800) );

  xor2  gate1163(.a(G779), .b(G651), .O(gate268inter0));
  nand2 gate1164(.a(gate268inter0), .b(s_88), .O(gate268inter1));
  and2  gate1165(.a(G779), .b(G651), .O(gate268inter2));
  inv1  gate1166(.a(s_88), .O(gate268inter3));
  inv1  gate1167(.a(s_89), .O(gate268inter4));
  nand2 gate1168(.a(gate268inter4), .b(gate268inter3), .O(gate268inter5));
  nor2  gate1169(.a(gate268inter5), .b(gate268inter2), .O(gate268inter6));
  inv1  gate1170(.a(G651), .O(gate268inter7));
  inv1  gate1171(.a(G779), .O(gate268inter8));
  nand2 gate1172(.a(gate268inter8), .b(gate268inter7), .O(gate268inter9));
  nand2 gate1173(.a(s_89), .b(gate268inter3), .O(gate268inter10));
  nor2  gate1174(.a(gate268inter10), .b(gate268inter9), .O(gate268inter11));
  nor2  gate1175(.a(gate268inter11), .b(gate268inter6), .O(gate268inter12));
  nand2 gate1176(.a(gate268inter12), .b(gate268inter1), .O(G803));
nand2 gate269( .a(G654), .b(G782), .O(G806) );

  xor2  gate589(.a(G785), .b(G657), .O(gate270inter0));
  nand2 gate590(.a(gate270inter0), .b(s_6), .O(gate270inter1));
  and2  gate591(.a(G785), .b(G657), .O(gate270inter2));
  inv1  gate592(.a(s_6), .O(gate270inter3));
  inv1  gate593(.a(s_7), .O(gate270inter4));
  nand2 gate594(.a(gate270inter4), .b(gate270inter3), .O(gate270inter5));
  nor2  gate595(.a(gate270inter5), .b(gate270inter2), .O(gate270inter6));
  inv1  gate596(.a(G657), .O(gate270inter7));
  inv1  gate597(.a(G785), .O(gate270inter8));
  nand2 gate598(.a(gate270inter8), .b(gate270inter7), .O(gate270inter9));
  nand2 gate599(.a(s_7), .b(gate270inter3), .O(gate270inter10));
  nor2  gate600(.a(gate270inter10), .b(gate270inter9), .O(gate270inter11));
  nor2  gate601(.a(gate270inter11), .b(gate270inter6), .O(gate270inter12));
  nand2 gate602(.a(gate270inter12), .b(gate270inter1), .O(G809));
nand2 gate271( .a(G660), .b(G788), .O(G812) );
nand2 gate272( .a(G663), .b(G791), .O(G815) );

  xor2  gate2437(.a(G794), .b(G642), .O(gate273inter0));
  nand2 gate2438(.a(gate273inter0), .b(s_270), .O(gate273inter1));
  and2  gate2439(.a(G794), .b(G642), .O(gate273inter2));
  inv1  gate2440(.a(s_270), .O(gate273inter3));
  inv1  gate2441(.a(s_271), .O(gate273inter4));
  nand2 gate2442(.a(gate273inter4), .b(gate273inter3), .O(gate273inter5));
  nor2  gate2443(.a(gate273inter5), .b(gate273inter2), .O(gate273inter6));
  inv1  gate2444(.a(G642), .O(gate273inter7));
  inv1  gate2445(.a(G794), .O(gate273inter8));
  nand2 gate2446(.a(gate273inter8), .b(gate273inter7), .O(gate273inter9));
  nand2 gate2447(.a(s_271), .b(gate273inter3), .O(gate273inter10));
  nor2  gate2448(.a(gate273inter10), .b(gate273inter9), .O(gate273inter11));
  nor2  gate2449(.a(gate273inter11), .b(gate273inter6), .O(gate273inter12));
  nand2 gate2450(.a(gate273inter12), .b(gate273inter1), .O(G818));

  xor2  gate855(.a(G794), .b(G770), .O(gate274inter0));
  nand2 gate856(.a(gate274inter0), .b(s_44), .O(gate274inter1));
  and2  gate857(.a(G794), .b(G770), .O(gate274inter2));
  inv1  gate858(.a(s_44), .O(gate274inter3));
  inv1  gate859(.a(s_45), .O(gate274inter4));
  nand2 gate860(.a(gate274inter4), .b(gate274inter3), .O(gate274inter5));
  nor2  gate861(.a(gate274inter5), .b(gate274inter2), .O(gate274inter6));
  inv1  gate862(.a(G770), .O(gate274inter7));
  inv1  gate863(.a(G794), .O(gate274inter8));
  nand2 gate864(.a(gate274inter8), .b(gate274inter7), .O(gate274inter9));
  nand2 gate865(.a(s_45), .b(gate274inter3), .O(gate274inter10));
  nor2  gate866(.a(gate274inter10), .b(gate274inter9), .O(gate274inter11));
  nor2  gate867(.a(gate274inter11), .b(gate274inter6), .O(gate274inter12));
  nand2 gate868(.a(gate274inter12), .b(gate274inter1), .O(G819));

  xor2  gate1695(.a(G797), .b(G645), .O(gate275inter0));
  nand2 gate1696(.a(gate275inter0), .b(s_164), .O(gate275inter1));
  and2  gate1697(.a(G797), .b(G645), .O(gate275inter2));
  inv1  gate1698(.a(s_164), .O(gate275inter3));
  inv1  gate1699(.a(s_165), .O(gate275inter4));
  nand2 gate1700(.a(gate275inter4), .b(gate275inter3), .O(gate275inter5));
  nor2  gate1701(.a(gate275inter5), .b(gate275inter2), .O(gate275inter6));
  inv1  gate1702(.a(G645), .O(gate275inter7));
  inv1  gate1703(.a(G797), .O(gate275inter8));
  nand2 gate1704(.a(gate275inter8), .b(gate275inter7), .O(gate275inter9));
  nand2 gate1705(.a(s_165), .b(gate275inter3), .O(gate275inter10));
  nor2  gate1706(.a(gate275inter10), .b(gate275inter9), .O(gate275inter11));
  nor2  gate1707(.a(gate275inter11), .b(gate275inter6), .O(gate275inter12));
  nand2 gate1708(.a(gate275inter12), .b(gate275inter1), .O(G820));
nand2 gate276( .a(G773), .b(G797), .O(G821) );
nand2 gate277( .a(G648), .b(G800), .O(G822) );
nand2 gate278( .a(G776), .b(G800), .O(G823) );

  xor2  gate2143(.a(G803), .b(G651), .O(gate279inter0));
  nand2 gate2144(.a(gate279inter0), .b(s_228), .O(gate279inter1));
  and2  gate2145(.a(G803), .b(G651), .O(gate279inter2));
  inv1  gate2146(.a(s_228), .O(gate279inter3));
  inv1  gate2147(.a(s_229), .O(gate279inter4));
  nand2 gate2148(.a(gate279inter4), .b(gate279inter3), .O(gate279inter5));
  nor2  gate2149(.a(gate279inter5), .b(gate279inter2), .O(gate279inter6));
  inv1  gate2150(.a(G651), .O(gate279inter7));
  inv1  gate2151(.a(G803), .O(gate279inter8));
  nand2 gate2152(.a(gate279inter8), .b(gate279inter7), .O(gate279inter9));
  nand2 gate2153(.a(s_229), .b(gate279inter3), .O(gate279inter10));
  nor2  gate2154(.a(gate279inter10), .b(gate279inter9), .O(gate279inter11));
  nor2  gate2155(.a(gate279inter11), .b(gate279inter6), .O(gate279inter12));
  nand2 gate2156(.a(gate279inter12), .b(gate279inter1), .O(G824));
nand2 gate280( .a(G779), .b(G803), .O(G825) );
nand2 gate281( .a(G654), .b(G806), .O(G826) );

  xor2  gate771(.a(G806), .b(G782), .O(gate282inter0));
  nand2 gate772(.a(gate282inter0), .b(s_32), .O(gate282inter1));
  and2  gate773(.a(G806), .b(G782), .O(gate282inter2));
  inv1  gate774(.a(s_32), .O(gate282inter3));
  inv1  gate775(.a(s_33), .O(gate282inter4));
  nand2 gate776(.a(gate282inter4), .b(gate282inter3), .O(gate282inter5));
  nor2  gate777(.a(gate282inter5), .b(gate282inter2), .O(gate282inter6));
  inv1  gate778(.a(G782), .O(gate282inter7));
  inv1  gate779(.a(G806), .O(gate282inter8));
  nand2 gate780(.a(gate282inter8), .b(gate282inter7), .O(gate282inter9));
  nand2 gate781(.a(s_33), .b(gate282inter3), .O(gate282inter10));
  nor2  gate782(.a(gate282inter10), .b(gate282inter9), .O(gate282inter11));
  nor2  gate783(.a(gate282inter11), .b(gate282inter6), .O(gate282inter12));
  nand2 gate784(.a(gate282inter12), .b(gate282inter1), .O(G827));

  xor2  gate1555(.a(G809), .b(G657), .O(gate283inter0));
  nand2 gate1556(.a(gate283inter0), .b(s_144), .O(gate283inter1));
  and2  gate1557(.a(G809), .b(G657), .O(gate283inter2));
  inv1  gate1558(.a(s_144), .O(gate283inter3));
  inv1  gate1559(.a(s_145), .O(gate283inter4));
  nand2 gate1560(.a(gate283inter4), .b(gate283inter3), .O(gate283inter5));
  nor2  gate1561(.a(gate283inter5), .b(gate283inter2), .O(gate283inter6));
  inv1  gate1562(.a(G657), .O(gate283inter7));
  inv1  gate1563(.a(G809), .O(gate283inter8));
  nand2 gate1564(.a(gate283inter8), .b(gate283inter7), .O(gate283inter9));
  nand2 gate1565(.a(s_145), .b(gate283inter3), .O(gate283inter10));
  nor2  gate1566(.a(gate283inter10), .b(gate283inter9), .O(gate283inter11));
  nor2  gate1567(.a(gate283inter11), .b(gate283inter6), .O(gate283inter12));
  nand2 gate1568(.a(gate283inter12), .b(gate283inter1), .O(G828));

  xor2  gate2255(.a(G809), .b(G785), .O(gate284inter0));
  nand2 gate2256(.a(gate284inter0), .b(s_244), .O(gate284inter1));
  and2  gate2257(.a(G809), .b(G785), .O(gate284inter2));
  inv1  gate2258(.a(s_244), .O(gate284inter3));
  inv1  gate2259(.a(s_245), .O(gate284inter4));
  nand2 gate2260(.a(gate284inter4), .b(gate284inter3), .O(gate284inter5));
  nor2  gate2261(.a(gate284inter5), .b(gate284inter2), .O(gate284inter6));
  inv1  gate2262(.a(G785), .O(gate284inter7));
  inv1  gate2263(.a(G809), .O(gate284inter8));
  nand2 gate2264(.a(gate284inter8), .b(gate284inter7), .O(gate284inter9));
  nand2 gate2265(.a(s_245), .b(gate284inter3), .O(gate284inter10));
  nor2  gate2266(.a(gate284inter10), .b(gate284inter9), .O(gate284inter11));
  nor2  gate2267(.a(gate284inter11), .b(gate284inter6), .O(gate284inter12));
  nand2 gate2268(.a(gate284inter12), .b(gate284inter1), .O(G829));

  xor2  gate1961(.a(G812), .b(G660), .O(gate285inter0));
  nand2 gate1962(.a(gate285inter0), .b(s_202), .O(gate285inter1));
  and2  gate1963(.a(G812), .b(G660), .O(gate285inter2));
  inv1  gate1964(.a(s_202), .O(gate285inter3));
  inv1  gate1965(.a(s_203), .O(gate285inter4));
  nand2 gate1966(.a(gate285inter4), .b(gate285inter3), .O(gate285inter5));
  nor2  gate1967(.a(gate285inter5), .b(gate285inter2), .O(gate285inter6));
  inv1  gate1968(.a(G660), .O(gate285inter7));
  inv1  gate1969(.a(G812), .O(gate285inter8));
  nand2 gate1970(.a(gate285inter8), .b(gate285inter7), .O(gate285inter9));
  nand2 gate1971(.a(s_203), .b(gate285inter3), .O(gate285inter10));
  nor2  gate1972(.a(gate285inter10), .b(gate285inter9), .O(gate285inter11));
  nor2  gate1973(.a(gate285inter11), .b(gate285inter6), .O(gate285inter12));
  nand2 gate1974(.a(gate285inter12), .b(gate285inter1), .O(G830));
nand2 gate286( .a(G788), .b(G812), .O(G831) );

  xor2  gate1807(.a(G815), .b(G663), .O(gate287inter0));
  nand2 gate1808(.a(gate287inter0), .b(s_180), .O(gate287inter1));
  and2  gate1809(.a(G815), .b(G663), .O(gate287inter2));
  inv1  gate1810(.a(s_180), .O(gate287inter3));
  inv1  gate1811(.a(s_181), .O(gate287inter4));
  nand2 gate1812(.a(gate287inter4), .b(gate287inter3), .O(gate287inter5));
  nor2  gate1813(.a(gate287inter5), .b(gate287inter2), .O(gate287inter6));
  inv1  gate1814(.a(G663), .O(gate287inter7));
  inv1  gate1815(.a(G815), .O(gate287inter8));
  nand2 gate1816(.a(gate287inter8), .b(gate287inter7), .O(gate287inter9));
  nand2 gate1817(.a(s_181), .b(gate287inter3), .O(gate287inter10));
  nor2  gate1818(.a(gate287inter10), .b(gate287inter9), .O(gate287inter11));
  nor2  gate1819(.a(gate287inter11), .b(gate287inter6), .O(gate287inter12));
  nand2 gate1820(.a(gate287inter12), .b(gate287inter1), .O(G832));
nand2 gate288( .a(G791), .b(G815), .O(G833) );
nand2 gate289( .a(G818), .b(G819), .O(G834) );
nand2 gate290( .a(G820), .b(G821), .O(G847) );
nand2 gate291( .a(G822), .b(G823), .O(G860) );

  xor2  gate2381(.a(G825), .b(G824), .O(gate292inter0));
  nand2 gate2382(.a(gate292inter0), .b(s_262), .O(gate292inter1));
  and2  gate2383(.a(G825), .b(G824), .O(gate292inter2));
  inv1  gate2384(.a(s_262), .O(gate292inter3));
  inv1  gate2385(.a(s_263), .O(gate292inter4));
  nand2 gate2386(.a(gate292inter4), .b(gate292inter3), .O(gate292inter5));
  nor2  gate2387(.a(gate292inter5), .b(gate292inter2), .O(gate292inter6));
  inv1  gate2388(.a(G824), .O(gate292inter7));
  inv1  gate2389(.a(G825), .O(gate292inter8));
  nand2 gate2390(.a(gate292inter8), .b(gate292inter7), .O(gate292inter9));
  nand2 gate2391(.a(s_263), .b(gate292inter3), .O(gate292inter10));
  nor2  gate2392(.a(gate292inter10), .b(gate292inter9), .O(gate292inter11));
  nor2  gate2393(.a(gate292inter11), .b(gate292inter6), .O(gate292inter12));
  nand2 gate2394(.a(gate292inter12), .b(gate292inter1), .O(G873));
nand2 gate293( .a(G828), .b(G829), .O(G886) );

  xor2  gate2185(.a(G833), .b(G832), .O(gate294inter0));
  nand2 gate2186(.a(gate294inter0), .b(s_234), .O(gate294inter1));
  and2  gate2187(.a(G833), .b(G832), .O(gate294inter2));
  inv1  gate2188(.a(s_234), .O(gate294inter3));
  inv1  gate2189(.a(s_235), .O(gate294inter4));
  nand2 gate2190(.a(gate294inter4), .b(gate294inter3), .O(gate294inter5));
  nor2  gate2191(.a(gate294inter5), .b(gate294inter2), .O(gate294inter6));
  inv1  gate2192(.a(G832), .O(gate294inter7));
  inv1  gate2193(.a(G833), .O(gate294inter8));
  nand2 gate2194(.a(gate294inter8), .b(gate294inter7), .O(gate294inter9));
  nand2 gate2195(.a(s_235), .b(gate294inter3), .O(gate294inter10));
  nor2  gate2196(.a(gate294inter10), .b(gate294inter9), .O(gate294inter11));
  nor2  gate2197(.a(gate294inter11), .b(gate294inter6), .O(gate294inter12));
  nand2 gate2198(.a(gate294inter12), .b(gate294inter1), .O(G899));

  xor2  gate827(.a(G831), .b(G830), .O(gate295inter0));
  nand2 gate828(.a(gate295inter0), .b(s_40), .O(gate295inter1));
  and2  gate829(.a(G831), .b(G830), .O(gate295inter2));
  inv1  gate830(.a(s_40), .O(gate295inter3));
  inv1  gate831(.a(s_41), .O(gate295inter4));
  nand2 gate832(.a(gate295inter4), .b(gate295inter3), .O(gate295inter5));
  nor2  gate833(.a(gate295inter5), .b(gate295inter2), .O(gate295inter6));
  inv1  gate834(.a(G830), .O(gate295inter7));
  inv1  gate835(.a(G831), .O(gate295inter8));
  nand2 gate836(.a(gate295inter8), .b(gate295inter7), .O(gate295inter9));
  nand2 gate837(.a(s_41), .b(gate295inter3), .O(gate295inter10));
  nor2  gate838(.a(gate295inter10), .b(gate295inter9), .O(gate295inter11));
  nor2  gate839(.a(gate295inter11), .b(gate295inter6), .O(gate295inter12));
  nand2 gate840(.a(gate295inter12), .b(gate295inter1), .O(G912));
nand2 gate296( .a(G826), .b(G827), .O(G925) );
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );
nand2 gate387( .a(G1), .b(G1036), .O(G1132) );

  xor2  gate1597(.a(G1039), .b(G2), .O(gate388inter0));
  nand2 gate1598(.a(gate388inter0), .b(s_150), .O(gate388inter1));
  and2  gate1599(.a(G1039), .b(G2), .O(gate388inter2));
  inv1  gate1600(.a(s_150), .O(gate388inter3));
  inv1  gate1601(.a(s_151), .O(gate388inter4));
  nand2 gate1602(.a(gate388inter4), .b(gate388inter3), .O(gate388inter5));
  nor2  gate1603(.a(gate388inter5), .b(gate388inter2), .O(gate388inter6));
  inv1  gate1604(.a(G2), .O(gate388inter7));
  inv1  gate1605(.a(G1039), .O(gate388inter8));
  nand2 gate1606(.a(gate388inter8), .b(gate388inter7), .O(gate388inter9));
  nand2 gate1607(.a(s_151), .b(gate388inter3), .O(gate388inter10));
  nor2  gate1608(.a(gate388inter10), .b(gate388inter9), .O(gate388inter11));
  nor2  gate1609(.a(gate388inter11), .b(gate388inter6), .O(gate388inter12));
  nand2 gate1610(.a(gate388inter12), .b(gate388inter1), .O(G1135));

  xor2  gate2003(.a(G1042), .b(G3), .O(gate389inter0));
  nand2 gate2004(.a(gate389inter0), .b(s_208), .O(gate389inter1));
  and2  gate2005(.a(G1042), .b(G3), .O(gate389inter2));
  inv1  gate2006(.a(s_208), .O(gate389inter3));
  inv1  gate2007(.a(s_209), .O(gate389inter4));
  nand2 gate2008(.a(gate389inter4), .b(gate389inter3), .O(gate389inter5));
  nor2  gate2009(.a(gate389inter5), .b(gate389inter2), .O(gate389inter6));
  inv1  gate2010(.a(G3), .O(gate389inter7));
  inv1  gate2011(.a(G1042), .O(gate389inter8));
  nand2 gate2012(.a(gate389inter8), .b(gate389inter7), .O(gate389inter9));
  nand2 gate2013(.a(s_209), .b(gate389inter3), .O(gate389inter10));
  nor2  gate2014(.a(gate389inter10), .b(gate389inter9), .O(gate389inter11));
  nor2  gate2015(.a(gate389inter11), .b(gate389inter6), .O(gate389inter12));
  nand2 gate2016(.a(gate389inter12), .b(gate389inter1), .O(G1138));
nand2 gate390( .a(G4), .b(G1045), .O(G1141) );

  xor2  gate2171(.a(G1048), .b(G5), .O(gate391inter0));
  nand2 gate2172(.a(gate391inter0), .b(s_232), .O(gate391inter1));
  and2  gate2173(.a(G1048), .b(G5), .O(gate391inter2));
  inv1  gate2174(.a(s_232), .O(gate391inter3));
  inv1  gate2175(.a(s_233), .O(gate391inter4));
  nand2 gate2176(.a(gate391inter4), .b(gate391inter3), .O(gate391inter5));
  nor2  gate2177(.a(gate391inter5), .b(gate391inter2), .O(gate391inter6));
  inv1  gate2178(.a(G5), .O(gate391inter7));
  inv1  gate2179(.a(G1048), .O(gate391inter8));
  nand2 gate2180(.a(gate391inter8), .b(gate391inter7), .O(gate391inter9));
  nand2 gate2181(.a(s_233), .b(gate391inter3), .O(gate391inter10));
  nor2  gate2182(.a(gate391inter10), .b(gate391inter9), .O(gate391inter11));
  nor2  gate2183(.a(gate391inter11), .b(gate391inter6), .O(gate391inter12));
  nand2 gate2184(.a(gate391inter12), .b(gate391inter1), .O(G1144));

  xor2  gate1177(.a(G1051), .b(G6), .O(gate392inter0));
  nand2 gate1178(.a(gate392inter0), .b(s_90), .O(gate392inter1));
  and2  gate1179(.a(G1051), .b(G6), .O(gate392inter2));
  inv1  gate1180(.a(s_90), .O(gate392inter3));
  inv1  gate1181(.a(s_91), .O(gate392inter4));
  nand2 gate1182(.a(gate392inter4), .b(gate392inter3), .O(gate392inter5));
  nor2  gate1183(.a(gate392inter5), .b(gate392inter2), .O(gate392inter6));
  inv1  gate1184(.a(G6), .O(gate392inter7));
  inv1  gate1185(.a(G1051), .O(gate392inter8));
  nand2 gate1186(.a(gate392inter8), .b(gate392inter7), .O(gate392inter9));
  nand2 gate1187(.a(s_91), .b(gate392inter3), .O(gate392inter10));
  nor2  gate1188(.a(gate392inter10), .b(gate392inter9), .O(gate392inter11));
  nor2  gate1189(.a(gate392inter11), .b(gate392inter6), .O(gate392inter12));
  nand2 gate1190(.a(gate392inter12), .b(gate392inter1), .O(G1147));
nand2 gate393( .a(G7), .b(G1054), .O(G1150) );
nand2 gate394( .a(G8), .b(G1057), .O(G1153) );
nand2 gate395( .a(G9), .b(G1060), .O(G1156) );

  xor2  gate743(.a(G1063), .b(G10), .O(gate396inter0));
  nand2 gate744(.a(gate396inter0), .b(s_28), .O(gate396inter1));
  and2  gate745(.a(G1063), .b(G10), .O(gate396inter2));
  inv1  gate746(.a(s_28), .O(gate396inter3));
  inv1  gate747(.a(s_29), .O(gate396inter4));
  nand2 gate748(.a(gate396inter4), .b(gate396inter3), .O(gate396inter5));
  nor2  gate749(.a(gate396inter5), .b(gate396inter2), .O(gate396inter6));
  inv1  gate750(.a(G10), .O(gate396inter7));
  inv1  gate751(.a(G1063), .O(gate396inter8));
  nand2 gate752(.a(gate396inter8), .b(gate396inter7), .O(gate396inter9));
  nand2 gate753(.a(s_29), .b(gate396inter3), .O(gate396inter10));
  nor2  gate754(.a(gate396inter10), .b(gate396inter9), .O(gate396inter11));
  nor2  gate755(.a(gate396inter11), .b(gate396inter6), .O(gate396inter12));
  nand2 gate756(.a(gate396inter12), .b(gate396inter1), .O(G1159));
nand2 gate397( .a(G11), .b(G1066), .O(G1162) );
nand2 gate398( .a(G12), .b(G1069), .O(G1165) );
nand2 gate399( .a(G13), .b(G1072), .O(G1168) );
nand2 gate400( .a(G14), .b(G1075), .O(G1171) );

  xor2  gate2367(.a(G1078), .b(G15), .O(gate401inter0));
  nand2 gate2368(.a(gate401inter0), .b(s_260), .O(gate401inter1));
  and2  gate2369(.a(G1078), .b(G15), .O(gate401inter2));
  inv1  gate2370(.a(s_260), .O(gate401inter3));
  inv1  gate2371(.a(s_261), .O(gate401inter4));
  nand2 gate2372(.a(gate401inter4), .b(gate401inter3), .O(gate401inter5));
  nor2  gate2373(.a(gate401inter5), .b(gate401inter2), .O(gate401inter6));
  inv1  gate2374(.a(G15), .O(gate401inter7));
  inv1  gate2375(.a(G1078), .O(gate401inter8));
  nand2 gate2376(.a(gate401inter8), .b(gate401inter7), .O(gate401inter9));
  nand2 gate2377(.a(s_261), .b(gate401inter3), .O(gate401inter10));
  nor2  gate2378(.a(gate401inter10), .b(gate401inter9), .O(gate401inter11));
  nor2  gate2379(.a(gate401inter11), .b(gate401inter6), .O(gate401inter12));
  nand2 gate2380(.a(gate401inter12), .b(gate401inter1), .O(G1174));

  xor2  gate1135(.a(G1081), .b(G16), .O(gate402inter0));
  nand2 gate1136(.a(gate402inter0), .b(s_84), .O(gate402inter1));
  and2  gate1137(.a(G1081), .b(G16), .O(gate402inter2));
  inv1  gate1138(.a(s_84), .O(gate402inter3));
  inv1  gate1139(.a(s_85), .O(gate402inter4));
  nand2 gate1140(.a(gate402inter4), .b(gate402inter3), .O(gate402inter5));
  nor2  gate1141(.a(gate402inter5), .b(gate402inter2), .O(gate402inter6));
  inv1  gate1142(.a(G16), .O(gate402inter7));
  inv1  gate1143(.a(G1081), .O(gate402inter8));
  nand2 gate1144(.a(gate402inter8), .b(gate402inter7), .O(gate402inter9));
  nand2 gate1145(.a(s_85), .b(gate402inter3), .O(gate402inter10));
  nor2  gate1146(.a(gate402inter10), .b(gate402inter9), .O(gate402inter11));
  nor2  gate1147(.a(gate402inter11), .b(gate402inter6), .O(gate402inter12));
  nand2 gate1148(.a(gate402inter12), .b(gate402inter1), .O(G1177));

  xor2  gate561(.a(G1084), .b(G17), .O(gate403inter0));
  nand2 gate562(.a(gate403inter0), .b(s_2), .O(gate403inter1));
  and2  gate563(.a(G1084), .b(G17), .O(gate403inter2));
  inv1  gate564(.a(s_2), .O(gate403inter3));
  inv1  gate565(.a(s_3), .O(gate403inter4));
  nand2 gate566(.a(gate403inter4), .b(gate403inter3), .O(gate403inter5));
  nor2  gate567(.a(gate403inter5), .b(gate403inter2), .O(gate403inter6));
  inv1  gate568(.a(G17), .O(gate403inter7));
  inv1  gate569(.a(G1084), .O(gate403inter8));
  nand2 gate570(.a(gate403inter8), .b(gate403inter7), .O(gate403inter9));
  nand2 gate571(.a(s_3), .b(gate403inter3), .O(gate403inter10));
  nor2  gate572(.a(gate403inter10), .b(gate403inter9), .O(gate403inter11));
  nor2  gate573(.a(gate403inter11), .b(gate403inter6), .O(gate403inter12));
  nand2 gate574(.a(gate403inter12), .b(gate403inter1), .O(G1180));

  xor2  gate2619(.a(G1087), .b(G18), .O(gate404inter0));
  nand2 gate2620(.a(gate404inter0), .b(s_296), .O(gate404inter1));
  and2  gate2621(.a(G1087), .b(G18), .O(gate404inter2));
  inv1  gate2622(.a(s_296), .O(gate404inter3));
  inv1  gate2623(.a(s_297), .O(gate404inter4));
  nand2 gate2624(.a(gate404inter4), .b(gate404inter3), .O(gate404inter5));
  nor2  gate2625(.a(gate404inter5), .b(gate404inter2), .O(gate404inter6));
  inv1  gate2626(.a(G18), .O(gate404inter7));
  inv1  gate2627(.a(G1087), .O(gate404inter8));
  nand2 gate2628(.a(gate404inter8), .b(gate404inter7), .O(gate404inter9));
  nand2 gate2629(.a(s_297), .b(gate404inter3), .O(gate404inter10));
  nor2  gate2630(.a(gate404inter10), .b(gate404inter9), .O(gate404inter11));
  nor2  gate2631(.a(gate404inter11), .b(gate404inter6), .O(gate404inter12));
  nand2 gate2632(.a(gate404inter12), .b(gate404inter1), .O(G1183));

  xor2  gate547(.a(G1090), .b(G19), .O(gate405inter0));
  nand2 gate548(.a(gate405inter0), .b(s_0), .O(gate405inter1));
  and2  gate549(.a(G1090), .b(G19), .O(gate405inter2));
  inv1  gate550(.a(s_0), .O(gate405inter3));
  inv1  gate551(.a(s_1), .O(gate405inter4));
  nand2 gate552(.a(gate405inter4), .b(gate405inter3), .O(gate405inter5));
  nor2  gate553(.a(gate405inter5), .b(gate405inter2), .O(gate405inter6));
  inv1  gate554(.a(G19), .O(gate405inter7));
  inv1  gate555(.a(G1090), .O(gate405inter8));
  nand2 gate556(.a(gate405inter8), .b(gate405inter7), .O(gate405inter9));
  nand2 gate557(.a(s_1), .b(gate405inter3), .O(gate405inter10));
  nor2  gate558(.a(gate405inter10), .b(gate405inter9), .O(gate405inter11));
  nor2  gate559(.a(gate405inter11), .b(gate405inter6), .O(gate405inter12));
  nand2 gate560(.a(gate405inter12), .b(gate405inter1), .O(G1186));
nand2 gate406( .a(G20), .b(G1093), .O(G1189) );
nand2 gate407( .a(G21), .b(G1096), .O(G1192) );
nand2 gate408( .a(G22), .b(G1099), .O(G1195) );

  xor2  gate2311(.a(G1102), .b(G23), .O(gate409inter0));
  nand2 gate2312(.a(gate409inter0), .b(s_252), .O(gate409inter1));
  and2  gate2313(.a(G1102), .b(G23), .O(gate409inter2));
  inv1  gate2314(.a(s_252), .O(gate409inter3));
  inv1  gate2315(.a(s_253), .O(gate409inter4));
  nand2 gate2316(.a(gate409inter4), .b(gate409inter3), .O(gate409inter5));
  nor2  gate2317(.a(gate409inter5), .b(gate409inter2), .O(gate409inter6));
  inv1  gate2318(.a(G23), .O(gate409inter7));
  inv1  gate2319(.a(G1102), .O(gate409inter8));
  nand2 gate2320(.a(gate409inter8), .b(gate409inter7), .O(gate409inter9));
  nand2 gate2321(.a(s_253), .b(gate409inter3), .O(gate409inter10));
  nor2  gate2322(.a(gate409inter10), .b(gate409inter9), .O(gate409inter11));
  nor2  gate2323(.a(gate409inter11), .b(gate409inter6), .O(gate409inter12));
  nand2 gate2324(.a(gate409inter12), .b(gate409inter1), .O(G1198));

  xor2  gate1793(.a(G1105), .b(G24), .O(gate410inter0));
  nand2 gate1794(.a(gate410inter0), .b(s_178), .O(gate410inter1));
  and2  gate1795(.a(G1105), .b(G24), .O(gate410inter2));
  inv1  gate1796(.a(s_178), .O(gate410inter3));
  inv1  gate1797(.a(s_179), .O(gate410inter4));
  nand2 gate1798(.a(gate410inter4), .b(gate410inter3), .O(gate410inter5));
  nor2  gate1799(.a(gate410inter5), .b(gate410inter2), .O(gate410inter6));
  inv1  gate1800(.a(G24), .O(gate410inter7));
  inv1  gate1801(.a(G1105), .O(gate410inter8));
  nand2 gate1802(.a(gate410inter8), .b(gate410inter7), .O(gate410inter9));
  nand2 gate1803(.a(s_179), .b(gate410inter3), .O(gate410inter10));
  nor2  gate1804(.a(gate410inter10), .b(gate410inter9), .O(gate410inter11));
  nor2  gate1805(.a(gate410inter11), .b(gate410inter6), .O(gate410inter12));
  nand2 gate1806(.a(gate410inter12), .b(gate410inter1), .O(G1201));
nand2 gate411( .a(G25), .b(G1108), .O(G1204) );
nand2 gate412( .a(G26), .b(G1111), .O(G1207) );
nand2 gate413( .a(G27), .b(G1114), .O(G1210) );
nand2 gate414( .a(G28), .b(G1117), .O(G1213) );

  xor2  gate2227(.a(G1120), .b(G29), .O(gate415inter0));
  nand2 gate2228(.a(gate415inter0), .b(s_240), .O(gate415inter1));
  and2  gate2229(.a(G1120), .b(G29), .O(gate415inter2));
  inv1  gate2230(.a(s_240), .O(gate415inter3));
  inv1  gate2231(.a(s_241), .O(gate415inter4));
  nand2 gate2232(.a(gate415inter4), .b(gate415inter3), .O(gate415inter5));
  nor2  gate2233(.a(gate415inter5), .b(gate415inter2), .O(gate415inter6));
  inv1  gate2234(.a(G29), .O(gate415inter7));
  inv1  gate2235(.a(G1120), .O(gate415inter8));
  nand2 gate2236(.a(gate415inter8), .b(gate415inter7), .O(gate415inter9));
  nand2 gate2237(.a(s_241), .b(gate415inter3), .O(gate415inter10));
  nor2  gate2238(.a(gate415inter10), .b(gate415inter9), .O(gate415inter11));
  nor2  gate2239(.a(gate415inter11), .b(gate415inter6), .O(gate415inter12));
  nand2 gate2240(.a(gate415inter12), .b(gate415inter1), .O(G1216));
nand2 gate416( .a(G30), .b(G1123), .O(G1219) );
nand2 gate417( .a(G31), .b(G1126), .O(G1222) );

  xor2  gate1275(.a(G1129), .b(G32), .O(gate418inter0));
  nand2 gate1276(.a(gate418inter0), .b(s_104), .O(gate418inter1));
  and2  gate1277(.a(G1129), .b(G32), .O(gate418inter2));
  inv1  gate1278(.a(s_104), .O(gate418inter3));
  inv1  gate1279(.a(s_105), .O(gate418inter4));
  nand2 gate1280(.a(gate418inter4), .b(gate418inter3), .O(gate418inter5));
  nor2  gate1281(.a(gate418inter5), .b(gate418inter2), .O(gate418inter6));
  inv1  gate1282(.a(G32), .O(gate418inter7));
  inv1  gate1283(.a(G1129), .O(gate418inter8));
  nand2 gate1284(.a(gate418inter8), .b(gate418inter7), .O(gate418inter9));
  nand2 gate1285(.a(s_105), .b(gate418inter3), .O(gate418inter10));
  nor2  gate1286(.a(gate418inter10), .b(gate418inter9), .O(gate418inter11));
  nor2  gate1287(.a(gate418inter11), .b(gate418inter6), .O(gate418inter12));
  nand2 gate1288(.a(gate418inter12), .b(gate418inter1), .O(G1225));
nand2 gate419( .a(G1), .b(G1132), .O(G1228) );

  xor2  gate2017(.a(G1132), .b(G1036), .O(gate420inter0));
  nand2 gate2018(.a(gate420inter0), .b(s_210), .O(gate420inter1));
  and2  gate2019(.a(G1132), .b(G1036), .O(gate420inter2));
  inv1  gate2020(.a(s_210), .O(gate420inter3));
  inv1  gate2021(.a(s_211), .O(gate420inter4));
  nand2 gate2022(.a(gate420inter4), .b(gate420inter3), .O(gate420inter5));
  nor2  gate2023(.a(gate420inter5), .b(gate420inter2), .O(gate420inter6));
  inv1  gate2024(.a(G1036), .O(gate420inter7));
  inv1  gate2025(.a(G1132), .O(gate420inter8));
  nand2 gate2026(.a(gate420inter8), .b(gate420inter7), .O(gate420inter9));
  nand2 gate2027(.a(s_211), .b(gate420inter3), .O(gate420inter10));
  nor2  gate2028(.a(gate420inter10), .b(gate420inter9), .O(gate420inter11));
  nor2  gate2029(.a(gate420inter11), .b(gate420inter6), .O(gate420inter12));
  nand2 gate2030(.a(gate420inter12), .b(gate420inter1), .O(G1229));
nand2 gate421( .a(G2), .b(G1135), .O(G1230) );
nand2 gate422( .a(G1039), .b(G1135), .O(G1231) );
nand2 gate423( .a(G3), .b(G1138), .O(G1232) );

  xor2  gate2689(.a(G1138), .b(G1042), .O(gate424inter0));
  nand2 gate2690(.a(gate424inter0), .b(s_306), .O(gate424inter1));
  and2  gate2691(.a(G1138), .b(G1042), .O(gate424inter2));
  inv1  gate2692(.a(s_306), .O(gate424inter3));
  inv1  gate2693(.a(s_307), .O(gate424inter4));
  nand2 gate2694(.a(gate424inter4), .b(gate424inter3), .O(gate424inter5));
  nor2  gate2695(.a(gate424inter5), .b(gate424inter2), .O(gate424inter6));
  inv1  gate2696(.a(G1042), .O(gate424inter7));
  inv1  gate2697(.a(G1138), .O(gate424inter8));
  nand2 gate2698(.a(gate424inter8), .b(gate424inter7), .O(gate424inter9));
  nand2 gate2699(.a(s_307), .b(gate424inter3), .O(gate424inter10));
  nor2  gate2700(.a(gate424inter10), .b(gate424inter9), .O(gate424inter11));
  nor2  gate2701(.a(gate424inter11), .b(gate424inter6), .O(gate424inter12));
  nand2 gate2702(.a(gate424inter12), .b(gate424inter1), .O(G1233));
nand2 gate425( .a(G4), .b(G1141), .O(G1234) );

  xor2  gate953(.a(G1141), .b(G1045), .O(gate426inter0));
  nand2 gate954(.a(gate426inter0), .b(s_58), .O(gate426inter1));
  and2  gate955(.a(G1141), .b(G1045), .O(gate426inter2));
  inv1  gate956(.a(s_58), .O(gate426inter3));
  inv1  gate957(.a(s_59), .O(gate426inter4));
  nand2 gate958(.a(gate426inter4), .b(gate426inter3), .O(gate426inter5));
  nor2  gate959(.a(gate426inter5), .b(gate426inter2), .O(gate426inter6));
  inv1  gate960(.a(G1045), .O(gate426inter7));
  inv1  gate961(.a(G1141), .O(gate426inter8));
  nand2 gate962(.a(gate426inter8), .b(gate426inter7), .O(gate426inter9));
  nand2 gate963(.a(s_59), .b(gate426inter3), .O(gate426inter10));
  nor2  gate964(.a(gate426inter10), .b(gate426inter9), .O(gate426inter11));
  nor2  gate965(.a(gate426inter11), .b(gate426inter6), .O(gate426inter12));
  nand2 gate966(.a(gate426inter12), .b(gate426inter1), .O(G1235));
nand2 gate427( .a(G5), .b(G1144), .O(G1236) );
nand2 gate428( .a(G1048), .b(G1144), .O(G1237) );
nand2 gate429( .a(G6), .b(G1147), .O(G1238) );

  xor2  gate1065(.a(G1147), .b(G1051), .O(gate430inter0));
  nand2 gate1066(.a(gate430inter0), .b(s_74), .O(gate430inter1));
  and2  gate1067(.a(G1147), .b(G1051), .O(gate430inter2));
  inv1  gate1068(.a(s_74), .O(gate430inter3));
  inv1  gate1069(.a(s_75), .O(gate430inter4));
  nand2 gate1070(.a(gate430inter4), .b(gate430inter3), .O(gate430inter5));
  nor2  gate1071(.a(gate430inter5), .b(gate430inter2), .O(gate430inter6));
  inv1  gate1072(.a(G1051), .O(gate430inter7));
  inv1  gate1073(.a(G1147), .O(gate430inter8));
  nand2 gate1074(.a(gate430inter8), .b(gate430inter7), .O(gate430inter9));
  nand2 gate1075(.a(s_75), .b(gate430inter3), .O(gate430inter10));
  nor2  gate1076(.a(gate430inter10), .b(gate430inter9), .O(gate430inter11));
  nor2  gate1077(.a(gate430inter11), .b(gate430inter6), .O(gate430inter12));
  nand2 gate1078(.a(gate430inter12), .b(gate430inter1), .O(G1239));
nand2 gate431( .a(G7), .b(G1150), .O(G1240) );
nand2 gate432( .a(G1054), .b(G1150), .O(G1241) );
nand2 gate433( .a(G8), .b(G1153), .O(G1242) );
nand2 gate434( .a(G1057), .b(G1153), .O(G1243) );
nand2 gate435( .a(G9), .b(G1156), .O(G1244) );

  xor2  gate1611(.a(G1156), .b(G1060), .O(gate436inter0));
  nand2 gate1612(.a(gate436inter0), .b(s_152), .O(gate436inter1));
  and2  gate1613(.a(G1156), .b(G1060), .O(gate436inter2));
  inv1  gate1614(.a(s_152), .O(gate436inter3));
  inv1  gate1615(.a(s_153), .O(gate436inter4));
  nand2 gate1616(.a(gate436inter4), .b(gate436inter3), .O(gate436inter5));
  nor2  gate1617(.a(gate436inter5), .b(gate436inter2), .O(gate436inter6));
  inv1  gate1618(.a(G1060), .O(gate436inter7));
  inv1  gate1619(.a(G1156), .O(gate436inter8));
  nand2 gate1620(.a(gate436inter8), .b(gate436inter7), .O(gate436inter9));
  nand2 gate1621(.a(s_153), .b(gate436inter3), .O(gate436inter10));
  nor2  gate1622(.a(gate436inter10), .b(gate436inter9), .O(gate436inter11));
  nor2  gate1623(.a(gate436inter11), .b(gate436inter6), .O(gate436inter12));
  nand2 gate1624(.a(gate436inter12), .b(gate436inter1), .O(G1245));
nand2 gate437( .a(G10), .b(G1159), .O(G1246) );

  xor2  gate813(.a(G1159), .b(G1063), .O(gate438inter0));
  nand2 gate814(.a(gate438inter0), .b(s_38), .O(gate438inter1));
  and2  gate815(.a(G1159), .b(G1063), .O(gate438inter2));
  inv1  gate816(.a(s_38), .O(gate438inter3));
  inv1  gate817(.a(s_39), .O(gate438inter4));
  nand2 gate818(.a(gate438inter4), .b(gate438inter3), .O(gate438inter5));
  nor2  gate819(.a(gate438inter5), .b(gate438inter2), .O(gate438inter6));
  inv1  gate820(.a(G1063), .O(gate438inter7));
  inv1  gate821(.a(G1159), .O(gate438inter8));
  nand2 gate822(.a(gate438inter8), .b(gate438inter7), .O(gate438inter9));
  nand2 gate823(.a(s_39), .b(gate438inter3), .O(gate438inter10));
  nor2  gate824(.a(gate438inter10), .b(gate438inter9), .O(gate438inter11));
  nor2  gate825(.a(gate438inter11), .b(gate438inter6), .O(gate438inter12));
  nand2 gate826(.a(gate438inter12), .b(gate438inter1), .O(G1247));

  xor2  gate575(.a(G1162), .b(G11), .O(gate439inter0));
  nand2 gate576(.a(gate439inter0), .b(s_4), .O(gate439inter1));
  and2  gate577(.a(G1162), .b(G11), .O(gate439inter2));
  inv1  gate578(.a(s_4), .O(gate439inter3));
  inv1  gate579(.a(s_5), .O(gate439inter4));
  nand2 gate580(.a(gate439inter4), .b(gate439inter3), .O(gate439inter5));
  nor2  gate581(.a(gate439inter5), .b(gate439inter2), .O(gate439inter6));
  inv1  gate582(.a(G11), .O(gate439inter7));
  inv1  gate583(.a(G1162), .O(gate439inter8));
  nand2 gate584(.a(gate439inter8), .b(gate439inter7), .O(gate439inter9));
  nand2 gate585(.a(s_5), .b(gate439inter3), .O(gate439inter10));
  nor2  gate586(.a(gate439inter10), .b(gate439inter9), .O(gate439inter11));
  nor2  gate587(.a(gate439inter11), .b(gate439inter6), .O(gate439inter12));
  nand2 gate588(.a(gate439inter12), .b(gate439inter1), .O(G1248));
nand2 gate440( .a(G1066), .b(G1162), .O(G1249) );

  xor2  gate1569(.a(G1165), .b(G12), .O(gate441inter0));
  nand2 gate1570(.a(gate441inter0), .b(s_146), .O(gate441inter1));
  and2  gate1571(.a(G1165), .b(G12), .O(gate441inter2));
  inv1  gate1572(.a(s_146), .O(gate441inter3));
  inv1  gate1573(.a(s_147), .O(gate441inter4));
  nand2 gate1574(.a(gate441inter4), .b(gate441inter3), .O(gate441inter5));
  nor2  gate1575(.a(gate441inter5), .b(gate441inter2), .O(gate441inter6));
  inv1  gate1576(.a(G12), .O(gate441inter7));
  inv1  gate1577(.a(G1165), .O(gate441inter8));
  nand2 gate1578(.a(gate441inter8), .b(gate441inter7), .O(gate441inter9));
  nand2 gate1579(.a(s_147), .b(gate441inter3), .O(gate441inter10));
  nor2  gate1580(.a(gate441inter10), .b(gate441inter9), .O(gate441inter11));
  nor2  gate1581(.a(gate441inter11), .b(gate441inter6), .O(gate441inter12));
  nand2 gate1582(.a(gate441inter12), .b(gate441inter1), .O(G1250));
nand2 gate442( .a(G1069), .b(G1165), .O(G1251) );
nand2 gate443( .a(G13), .b(G1168), .O(G1252) );

  xor2  gate785(.a(G1168), .b(G1072), .O(gate444inter0));
  nand2 gate786(.a(gate444inter0), .b(s_34), .O(gate444inter1));
  and2  gate787(.a(G1168), .b(G1072), .O(gate444inter2));
  inv1  gate788(.a(s_34), .O(gate444inter3));
  inv1  gate789(.a(s_35), .O(gate444inter4));
  nand2 gate790(.a(gate444inter4), .b(gate444inter3), .O(gate444inter5));
  nor2  gate791(.a(gate444inter5), .b(gate444inter2), .O(gate444inter6));
  inv1  gate792(.a(G1072), .O(gate444inter7));
  inv1  gate793(.a(G1168), .O(gate444inter8));
  nand2 gate794(.a(gate444inter8), .b(gate444inter7), .O(gate444inter9));
  nand2 gate795(.a(s_35), .b(gate444inter3), .O(gate444inter10));
  nor2  gate796(.a(gate444inter10), .b(gate444inter9), .O(gate444inter11));
  nor2  gate797(.a(gate444inter11), .b(gate444inter6), .O(gate444inter12));
  nand2 gate798(.a(gate444inter12), .b(gate444inter1), .O(G1253));
nand2 gate445( .a(G14), .b(G1171), .O(G1254) );

  xor2  gate1303(.a(G1171), .b(G1075), .O(gate446inter0));
  nand2 gate1304(.a(gate446inter0), .b(s_108), .O(gate446inter1));
  and2  gate1305(.a(G1171), .b(G1075), .O(gate446inter2));
  inv1  gate1306(.a(s_108), .O(gate446inter3));
  inv1  gate1307(.a(s_109), .O(gate446inter4));
  nand2 gate1308(.a(gate446inter4), .b(gate446inter3), .O(gate446inter5));
  nor2  gate1309(.a(gate446inter5), .b(gate446inter2), .O(gate446inter6));
  inv1  gate1310(.a(G1075), .O(gate446inter7));
  inv1  gate1311(.a(G1171), .O(gate446inter8));
  nand2 gate1312(.a(gate446inter8), .b(gate446inter7), .O(gate446inter9));
  nand2 gate1313(.a(s_109), .b(gate446inter3), .O(gate446inter10));
  nor2  gate1314(.a(gate446inter10), .b(gate446inter9), .O(gate446inter11));
  nor2  gate1315(.a(gate446inter11), .b(gate446inter6), .O(gate446inter12));
  nand2 gate1316(.a(gate446inter12), .b(gate446inter1), .O(G1255));
nand2 gate447( .a(G15), .b(G1174), .O(G1256) );
nand2 gate448( .a(G1078), .b(G1174), .O(G1257) );
nand2 gate449( .a(G16), .b(G1177), .O(G1258) );

  xor2  gate2507(.a(G1177), .b(G1081), .O(gate450inter0));
  nand2 gate2508(.a(gate450inter0), .b(s_280), .O(gate450inter1));
  and2  gate2509(.a(G1177), .b(G1081), .O(gate450inter2));
  inv1  gate2510(.a(s_280), .O(gate450inter3));
  inv1  gate2511(.a(s_281), .O(gate450inter4));
  nand2 gate2512(.a(gate450inter4), .b(gate450inter3), .O(gate450inter5));
  nor2  gate2513(.a(gate450inter5), .b(gate450inter2), .O(gate450inter6));
  inv1  gate2514(.a(G1081), .O(gate450inter7));
  inv1  gate2515(.a(G1177), .O(gate450inter8));
  nand2 gate2516(.a(gate450inter8), .b(gate450inter7), .O(gate450inter9));
  nand2 gate2517(.a(s_281), .b(gate450inter3), .O(gate450inter10));
  nor2  gate2518(.a(gate450inter10), .b(gate450inter9), .O(gate450inter11));
  nor2  gate2519(.a(gate450inter11), .b(gate450inter6), .O(gate450inter12));
  nand2 gate2520(.a(gate450inter12), .b(gate450inter1), .O(G1259));

  xor2  gate2647(.a(G1180), .b(G17), .O(gate451inter0));
  nand2 gate2648(.a(gate451inter0), .b(s_300), .O(gate451inter1));
  and2  gate2649(.a(G1180), .b(G17), .O(gate451inter2));
  inv1  gate2650(.a(s_300), .O(gate451inter3));
  inv1  gate2651(.a(s_301), .O(gate451inter4));
  nand2 gate2652(.a(gate451inter4), .b(gate451inter3), .O(gate451inter5));
  nor2  gate2653(.a(gate451inter5), .b(gate451inter2), .O(gate451inter6));
  inv1  gate2654(.a(G17), .O(gate451inter7));
  inv1  gate2655(.a(G1180), .O(gate451inter8));
  nand2 gate2656(.a(gate451inter8), .b(gate451inter7), .O(gate451inter9));
  nand2 gate2657(.a(s_301), .b(gate451inter3), .O(gate451inter10));
  nor2  gate2658(.a(gate451inter10), .b(gate451inter9), .O(gate451inter11));
  nor2  gate2659(.a(gate451inter11), .b(gate451inter6), .O(gate451inter12));
  nand2 gate2660(.a(gate451inter12), .b(gate451inter1), .O(G1260));
nand2 gate452( .a(G1084), .b(G1180), .O(G1261) );

  xor2  gate2451(.a(G1183), .b(G18), .O(gate453inter0));
  nand2 gate2452(.a(gate453inter0), .b(s_272), .O(gate453inter1));
  and2  gate2453(.a(G1183), .b(G18), .O(gate453inter2));
  inv1  gate2454(.a(s_272), .O(gate453inter3));
  inv1  gate2455(.a(s_273), .O(gate453inter4));
  nand2 gate2456(.a(gate453inter4), .b(gate453inter3), .O(gate453inter5));
  nor2  gate2457(.a(gate453inter5), .b(gate453inter2), .O(gate453inter6));
  inv1  gate2458(.a(G18), .O(gate453inter7));
  inv1  gate2459(.a(G1183), .O(gate453inter8));
  nand2 gate2460(.a(gate453inter8), .b(gate453inter7), .O(gate453inter9));
  nand2 gate2461(.a(s_273), .b(gate453inter3), .O(gate453inter10));
  nor2  gate2462(.a(gate453inter10), .b(gate453inter9), .O(gate453inter11));
  nor2  gate2463(.a(gate453inter11), .b(gate453inter6), .O(gate453inter12));
  nand2 gate2464(.a(gate453inter12), .b(gate453inter1), .O(G1262));

  xor2  gate1191(.a(G1183), .b(G1087), .O(gate454inter0));
  nand2 gate1192(.a(gate454inter0), .b(s_92), .O(gate454inter1));
  and2  gate1193(.a(G1183), .b(G1087), .O(gate454inter2));
  inv1  gate1194(.a(s_92), .O(gate454inter3));
  inv1  gate1195(.a(s_93), .O(gate454inter4));
  nand2 gate1196(.a(gate454inter4), .b(gate454inter3), .O(gate454inter5));
  nor2  gate1197(.a(gate454inter5), .b(gate454inter2), .O(gate454inter6));
  inv1  gate1198(.a(G1087), .O(gate454inter7));
  inv1  gate1199(.a(G1183), .O(gate454inter8));
  nand2 gate1200(.a(gate454inter8), .b(gate454inter7), .O(gate454inter9));
  nand2 gate1201(.a(s_93), .b(gate454inter3), .O(gate454inter10));
  nor2  gate1202(.a(gate454inter10), .b(gate454inter9), .O(gate454inter11));
  nor2  gate1203(.a(gate454inter11), .b(gate454inter6), .O(gate454inter12));
  nand2 gate1204(.a(gate454inter12), .b(gate454inter1), .O(G1263));
nand2 gate455( .a(G19), .b(G1186), .O(G1264) );
nand2 gate456( .a(G1090), .b(G1186), .O(G1265) );

  xor2  gate2059(.a(G1189), .b(G20), .O(gate457inter0));
  nand2 gate2060(.a(gate457inter0), .b(s_216), .O(gate457inter1));
  and2  gate2061(.a(G1189), .b(G20), .O(gate457inter2));
  inv1  gate2062(.a(s_216), .O(gate457inter3));
  inv1  gate2063(.a(s_217), .O(gate457inter4));
  nand2 gate2064(.a(gate457inter4), .b(gate457inter3), .O(gate457inter5));
  nor2  gate2065(.a(gate457inter5), .b(gate457inter2), .O(gate457inter6));
  inv1  gate2066(.a(G20), .O(gate457inter7));
  inv1  gate2067(.a(G1189), .O(gate457inter8));
  nand2 gate2068(.a(gate457inter8), .b(gate457inter7), .O(gate457inter9));
  nand2 gate2069(.a(s_217), .b(gate457inter3), .O(gate457inter10));
  nor2  gate2070(.a(gate457inter10), .b(gate457inter9), .O(gate457inter11));
  nor2  gate2071(.a(gate457inter11), .b(gate457inter6), .O(gate457inter12));
  nand2 gate2072(.a(gate457inter12), .b(gate457inter1), .O(G1266));
nand2 gate458( .a(G1093), .b(G1189), .O(G1267) );
nand2 gate459( .a(G21), .b(G1192), .O(G1268) );

  xor2  gate1751(.a(G1192), .b(G1096), .O(gate460inter0));
  nand2 gate1752(.a(gate460inter0), .b(s_172), .O(gate460inter1));
  and2  gate1753(.a(G1192), .b(G1096), .O(gate460inter2));
  inv1  gate1754(.a(s_172), .O(gate460inter3));
  inv1  gate1755(.a(s_173), .O(gate460inter4));
  nand2 gate1756(.a(gate460inter4), .b(gate460inter3), .O(gate460inter5));
  nor2  gate1757(.a(gate460inter5), .b(gate460inter2), .O(gate460inter6));
  inv1  gate1758(.a(G1096), .O(gate460inter7));
  inv1  gate1759(.a(G1192), .O(gate460inter8));
  nand2 gate1760(.a(gate460inter8), .b(gate460inter7), .O(gate460inter9));
  nand2 gate1761(.a(s_173), .b(gate460inter3), .O(gate460inter10));
  nor2  gate1762(.a(gate460inter10), .b(gate460inter9), .O(gate460inter11));
  nor2  gate1763(.a(gate460inter11), .b(gate460inter6), .O(gate460inter12));
  nand2 gate1764(.a(gate460inter12), .b(gate460inter1), .O(G1269));

  xor2  gate841(.a(G1195), .b(G22), .O(gate461inter0));
  nand2 gate842(.a(gate461inter0), .b(s_42), .O(gate461inter1));
  and2  gate843(.a(G1195), .b(G22), .O(gate461inter2));
  inv1  gate844(.a(s_42), .O(gate461inter3));
  inv1  gate845(.a(s_43), .O(gate461inter4));
  nand2 gate846(.a(gate461inter4), .b(gate461inter3), .O(gate461inter5));
  nor2  gate847(.a(gate461inter5), .b(gate461inter2), .O(gate461inter6));
  inv1  gate848(.a(G22), .O(gate461inter7));
  inv1  gate849(.a(G1195), .O(gate461inter8));
  nand2 gate850(.a(gate461inter8), .b(gate461inter7), .O(gate461inter9));
  nand2 gate851(.a(s_43), .b(gate461inter3), .O(gate461inter10));
  nor2  gate852(.a(gate461inter10), .b(gate461inter9), .O(gate461inter11));
  nor2  gate853(.a(gate461inter11), .b(gate461inter6), .O(gate461inter12));
  nand2 gate854(.a(gate461inter12), .b(gate461inter1), .O(G1270));
nand2 gate462( .a(G1099), .b(G1195), .O(G1271) );
nand2 gate463( .a(G23), .b(G1198), .O(G1272) );
nand2 gate464( .a(G1102), .b(G1198), .O(G1273) );
nand2 gate465( .a(G24), .b(G1201), .O(G1274) );
nand2 gate466( .a(G1105), .b(G1201), .O(G1275) );
nand2 gate467( .a(G25), .b(G1204), .O(G1276) );

  xor2  gate1037(.a(G1204), .b(G1108), .O(gate468inter0));
  nand2 gate1038(.a(gate468inter0), .b(s_70), .O(gate468inter1));
  and2  gate1039(.a(G1204), .b(G1108), .O(gate468inter2));
  inv1  gate1040(.a(s_70), .O(gate468inter3));
  inv1  gate1041(.a(s_71), .O(gate468inter4));
  nand2 gate1042(.a(gate468inter4), .b(gate468inter3), .O(gate468inter5));
  nor2  gate1043(.a(gate468inter5), .b(gate468inter2), .O(gate468inter6));
  inv1  gate1044(.a(G1108), .O(gate468inter7));
  inv1  gate1045(.a(G1204), .O(gate468inter8));
  nand2 gate1046(.a(gate468inter8), .b(gate468inter7), .O(gate468inter9));
  nand2 gate1047(.a(s_71), .b(gate468inter3), .O(gate468inter10));
  nor2  gate1048(.a(gate468inter10), .b(gate468inter9), .O(gate468inter11));
  nor2  gate1049(.a(gate468inter11), .b(gate468inter6), .O(gate468inter12));
  nand2 gate1050(.a(gate468inter12), .b(gate468inter1), .O(G1277));

  xor2  gate1541(.a(G1207), .b(G26), .O(gate469inter0));
  nand2 gate1542(.a(gate469inter0), .b(s_142), .O(gate469inter1));
  and2  gate1543(.a(G1207), .b(G26), .O(gate469inter2));
  inv1  gate1544(.a(s_142), .O(gate469inter3));
  inv1  gate1545(.a(s_143), .O(gate469inter4));
  nand2 gate1546(.a(gate469inter4), .b(gate469inter3), .O(gate469inter5));
  nor2  gate1547(.a(gate469inter5), .b(gate469inter2), .O(gate469inter6));
  inv1  gate1548(.a(G26), .O(gate469inter7));
  inv1  gate1549(.a(G1207), .O(gate469inter8));
  nand2 gate1550(.a(gate469inter8), .b(gate469inter7), .O(gate469inter9));
  nand2 gate1551(.a(s_143), .b(gate469inter3), .O(gate469inter10));
  nor2  gate1552(.a(gate469inter10), .b(gate469inter9), .O(gate469inter11));
  nor2  gate1553(.a(gate469inter11), .b(gate469inter6), .O(gate469inter12));
  nand2 gate1554(.a(gate469inter12), .b(gate469inter1), .O(G1278));
nand2 gate470( .a(G1111), .b(G1207), .O(G1279) );

  xor2  gate2605(.a(G1210), .b(G27), .O(gate471inter0));
  nand2 gate2606(.a(gate471inter0), .b(s_294), .O(gate471inter1));
  and2  gate2607(.a(G1210), .b(G27), .O(gate471inter2));
  inv1  gate2608(.a(s_294), .O(gate471inter3));
  inv1  gate2609(.a(s_295), .O(gate471inter4));
  nand2 gate2610(.a(gate471inter4), .b(gate471inter3), .O(gate471inter5));
  nor2  gate2611(.a(gate471inter5), .b(gate471inter2), .O(gate471inter6));
  inv1  gate2612(.a(G27), .O(gate471inter7));
  inv1  gate2613(.a(G1210), .O(gate471inter8));
  nand2 gate2614(.a(gate471inter8), .b(gate471inter7), .O(gate471inter9));
  nand2 gate2615(.a(s_295), .b(gate471inter3), .O(gate471inter10));
  nor2  gate2616(.a(gate471inter10), .b(gate471inter9), .O(gate471inter11));
  nor2  gate2617(.a(gate471inter11), .b(gate471inter6), .O(gate471inter12));
  nand2 gate2618(.a(gate471inter12), .b(gate471inter1), .O(G1280));

  xor2  gate1009(.a(G1210), .b(G1114), .O(gate472inter0));
  nand2 gate1010(.a(gate472inter0), .b(s_66), .O(gate472inter1));
  and2  gate1011(.a(G1210), .b(G1114), .O(gate472inter2));
  inv1  gate1012(.a(s_66), .O(gate472inter3));
  inv1  gate1013(.a(s_67), .O(gate472inter4));
  nand2 gate1014(.a(gate472inter4), .b(gate472inter3), .O(gate472inter5));
  nor2  gate1015(.a(gate472inter5), .b(gate472inter2), .O(gate472inter6));
  inv1  gate1016(.a(G1114), .O(gate472inter7));
  inv1  gate1017(.a(G1210), .O(gate472inter8));
  nand2 gate1018(.a(gate472inter8), .b(gate472inter7), .O(gate472inter9));
  nand2 gate1019(.a(s_67), .b(gate472inter3), .O(gate472inter10));
  nor2  gate1020(.a(gate472inter10), .b(gate472inter9), .O(gate472inter11));
  nor2  gate1021(.a(gate472inter11), .b(gate472inter6), .O(gate472inter12));
  nand2 gate1022(.a(gate472inter12), .b(gate472inter1), .O(G1281));
nand2 gate473( .a(G28), .b(G1213), .O(G1282) );
nand2 gate474( .a(G1117), .b(G1213), .O(G1283) );
nand2 gate475( .a(G29), .b(G1216), .O(G1284) );

  xor2  gate2241(.a(G1216), .b(G1120), .O(gate476inter0));
  nand2 gate2242(.a(gate476inter0), .b(s_242), .O(gate476inter1));
  and2  gate2243(.a(G1216), .b(G1120), .O(gate476inter2));
  inv1  gate2244(.a(s_242), .O(gate476inter3));
  inv1  gate2245(.a(s_243), .O(gate476inter4));
  nand2 gate2246(.a(gate476inter4), .b(gate476inter3), .O(gate476inter5));
  nor2  gate2247(.a(gate476inter5), .b(gate476inter2), .O(gate476inter6));
  inv1  gate2248(.a(G1120), .O(gate476inter7));
  inv1  gate2249(.a(G1216), .O(gate476inter8));
  nand2 gate2250(.a(gate476inter8), .b(gate476inter7), .O(gate476inter9));
  nand2 gate2251(.a(s_243), .b(gate476inter3), .O(gate476inter10));
  nor2  gate2252(.a(gate476inter10), .b(gate476inter9), .O(gate476inter11));
  nor2  gate2253(.a(gate476inter11), .b(gate476inter6), .O(gate476inter12));
  nand2 gate2254(.a(gate476inter12), .b(gate476inter1), .O(G1285));
nand2 gate477( .a(G30), .b(G1219), .O(G1286) );
nand2 gate478( .a(G1123), .b(G1219), .O(G1287) );
nand2 gate479( .a(G31), .b(G1222), .O(G1288) );

  xor2  gate1415(.a(G1222), .b(G1126), .O(gate480inter0));
  nand2 gate1416(.a(gate480inter0), .b(s_124), .O(gate480inter1));
  and2  gate1417(.a(G1222), .b(G1126), .O(gate480inter2));
  inv1  gate1418(.a(s_124), .O(gate480inter3));
  inv1  gate1419(.a(s_125), .O(gate480inter4));
  nand2 gate1420(.a(gate480inter4), .b(gate480inter3), .O(gate480inter5));
  nor2  gate1421(.a(gate480inter5), .b(gate480inter2), .O(gate480inter6));
  inv1  gate1422(.a(G1126), .O(gate480inter7));
  inv1  gate1423(.a(G1222), .O(gate480inter8));
  nand2 gate1424(.a(gate480inter8), .b(gate480inter7), .O(gate480inter9));
  nand2 gate1425(.a(s_125), .b(gate480inter3), .O(gate480inter10));
  nor2  gate1426(.a(gate480inter10), .b(gate480inter9), .O(gate480inter11));
  nor2  gate1427(.a(gate480inter11), .b(gate480inter6), .O(gate480inter12));
  nand2 gate1428(.a(gate480inter12), .b(gate480inter1), .O(G1289));

  xor2  gate1723(.a(G1225), .b(G32), .O(gate481inter0));
  nand2 gate1724(.a(gate481inter0), .b(s_168), .O(gate481inter1));
  and2  gate1725(.a(G1225), .b(G32), .O(gate481inter2));
  inv1  gate1726(.a(s_168), .O(gate481inter3));
  inv1  gate1727(.a(s_169), .O(gate481inter4));
  nand2 gate1728(.a(gate481inter4), .b(gate481inter3), .O(gate481inter5));
  nor2  gate1729(.a(gate481inter5), .b(gate481inter2), .O(gate481inter6));
  inv1  gate1730(.a(G32), .O(gate481inter7));
  inv1  gate1731(.a(G1225), .O(gate481inter8));
  nand2 gate1732(.a(gate481inter8), .b(gate481inter7), .O(gate481inter9));
  nand2 gate1733(.a(s_169), .b(gate481inter3), .O(gate481inter10));
  nor2  gate1734(.a(gate481inter10), .b(gate481inter9), .O(gate481inter11));
  nor2  gate1735(.a(gate481inter11), .b(gate481inter6), .O(gate481inter12));
  nand2 gate1736(.a(gate481inter12), .b(gate481inter1), .O(G1290));
nand2 gate482( .a(G1129), .b(G1225), .O(G1291) );
nand2 gate483( .a(G1228), .b(G1229), .O(G1292) );
nand2 gate484( .a(G1230), .b(G1231), .O(G1293) );

  xor2  gate1905(.a(G1233), .b(G1232), .O(gate485inter0));
  nand2 gate1906(.a(gate485inter0), .b(s_194), .O(gate485inter1));
  and2  gate1907(.a(G1233), .b(G1232), .O(gate485inter2));
  inv1  gate1908(.a(s_194), .O(gate485inter3));
  inv1  gate1909(.a(s_195), .O(gate485inter4));
  nand2 gate1910(.a(gate485inter4), .b(gate485inter3), .O(gate485inter5));
  nor2  gate1911(.a(gate485inter5), .b(gate485inter2), .O(gate485inter6));
  inv1  gate1912(.a(G1232), .O(gate485inter7));
  inv1  gate1913(.a(G1233), .O(gate485inter8));
  nand2 gate1914(.a(gate485inter8), .b(gate485inter7), .O(gate485inter9));
  nand2 gate1915(.a(s_195), .b(gate485inter3), .O(gate485inter10));
  nor2  gate1916(.a(gate485inter10), .b(gate485inter9), .O(gate485inter11));
  nor2  gate1917(.a(gate485inter11), .b(gate485inter6), .O(gate485inter12));
  nand2 gate1918(.a(gate485inter12), .b(gate485inter1), .O(G1294));
nand2 gate486( .a(G1234), .b(G1235), .O(G1295) );
nand2 gate487( .a(G1236), .b(G1237), .O(G1296) );

  xor2  gate1373(.a(G1239), .b(G1238), .O(gate488inter0));
  nand2 gate1374(.a(gate488inter0), .b(s_118), .O(gate488inter1));
  and2  gate1375(.a(G1239), .b(G1238), .O(gate488inter2));
  inv1  gate1376(.a(s_118), .O(gate488inter3));
  inv1  gate1377(.a(s_119), .O(gate488inter4));
  nand2 gate1378(.a(gate488inter4), .b(gate488inter3), .O(gate488inter5));
  nor2  gate1379(.a(gate488inter5), .b(gate488inter2), .O(gate488inter6));
  inv1  gate1380(.a(G1238), .O(gate488inter7));
  inv1  gate1381(.a(G1239), .O(gate488inter8));
  nand2 gate1382(.a(gate488inter8), .b(gate488inter7), .O(gate488inter9));
  nand2 gate1383(.a(s_119), .b(gate488inter3), .O(gate488inter10));
  nor2  gate1384(.a(gate488inter10), .b(gate488inter9), .O(gate488inter11));
  nor2  gate1385(.a(gate488inter11), .b(gate488inter6), .O(gate488inter12));
  nand2 gate1386(.a(gate488inter12), .b(gate488inter1), .O(G1297));
nand2 gate489( .a(G1240), .b(G1241), .O(G1298) );

  xor2  gate631(.a(G1243), .b(G1242), .O(gate490inter0));
  nand2 gate632(.a(gate490inter0), .b(s_12), .O(gate490inter1));
  and2  gate633(.a(G1243), .b(G1242), .O(gate490inter2));
  inv1  gate634(.a(s_12), .O(gate490inter3));
  inv1  gate635(.a(s_13), .O(gate490inter4));
  nand2 gate636(.a(gate490inter4), .b(gate490inter3), .O(gate490inter5));
  nor2  gate637(.a(gate490inter5), .b(gate490inter2), .O(gate490inter6));
  inv1  gate638(.a(G1242), .O(gate490inter7));
  inv1  gate639(.a(G1243), .O(gate490inter8));
  nand2 gate640(.a(gate490inter8), .b(gate490inter7), .O(gate490inter9));
  nand2 gate641(.a(s_13), .b(gate490inter3), .O(gate490inter10));
  nor2  gate642(.a(gate490inter10), .b(gate490inter9), .O(gate490inter11));
  nor2  gate643(.a(gate490inter11), .b(gate490inter6), .O(gate490inter12));
  nand2 gate644(.a(gate490inter12), .b(gate490inter1), .O(G1299));
nand2 gate491( .a(G1244), .b(G1245), .O(G1300) );

  xor2  gate2675(.a(G1247), .b(G1246), .O(gate492inter0));
  nand2 gate2676(.a(gate492inter0), .b(s_304), .O(gate492inter1));
  and2  gate2677(.a(G1247), .b(G1246), .O(gate492inter2));
  inv1  gate2678(.a(s_304), .O(gate492inter3));
  inv1  gate2679(.a(s_305), .O(gate492inter4));
  nand2 gate2680(.a(gate492inter4), .b(gate492inter3), .O(gate492inter5));
  nor2  gate2681(.a(gate492inter5), .b(gate492inter2), .O(gate492inter6));
  inv1  gate2682(.a(G1246), .O(gate492inter7));
  inv1  gate2683(.a(G1247), .O(gate492inter8));
  nand2 gate2684(.a(gate492inter8), .b(gate492inter7), .O(gate492inter9));
  nand2 gate2685(.a(s_305), .b(gate492inter3), .O(gate492inter10));
  nor2  gate2686(.a(gate492inter10), .b(gate492inter9), .O(gate492inter11));
  nor2  gate2687(.a(gate492inter11), .b(gate492inter6), .O(gate492inter12));
  nand2 gate2688(.a(gate492inter12), .b(gate492inter1), .O(G1301));
nand2 gate493( .a(G1248), .b(G1249), .O(G1302) );
nand2 gate494( .a(G1250), .b(G1251), .O(G1303) );
nand2 gate495( .a(G1252), .b(G1253), .O(G1304) );
nand2 gate496( .a(G1254), .b(G1255), .O(G1305) );

  xor2  gate1891(.a(G1257), .b(G1256), .O(gate497inter0));
  nand2 gate1892(.a(gate497inter0), .b(s_192), .O(gate497inter1));
  and2  gate1893(.a(G1257), .b(G1256), .O(gate497inter2));
  inv1  gate1894(.a(s_192), .O(gate497inter3));
  inv1  gate1895(.a(s_193), .O(gate497inter4));
  nand2 gate1896(.a(gate497inter4), .b(gate497inter3), .O(gate497inter5));
  nor2  gate1897(.a(gate497inter5), .b(gate497inter2), .O(gate497inter6));
  inv1  gate1898(.a(G1256), .O(gate497inter7));
  inv1  gate1899(.a(G1257), .O(gate497inter8));
  nand2 gate1900(.a(gate497inter8), .b(gate497inter7), .O(gate497inter9));
  nand2 gate1901(.a(s_193), .b(gate497inter3), .O(gate497inter10));
  nor2  gate1902(.a(gate497inter10), .b(gate497inter9), .O(gate497inter11));
  nor2  gate1903(.a(gate497inter11), .b(gate497inter6), .O(gate497inter12));
  nand2 gate1904(.a(gate497inter12), .b(gate497inter1), .O(G1306));
nand2 gate498( .a(G1258), .b(G1259), .O(G1307) );
nand2 gate499( .a(G1260), .b(G1261), .O(G1308) );

  xor2  gate1667(.a(G1263), .b(G1262), .O(gate500inter0));
  nand2 gate1668(.a(gate500inter0), .b(s_160), .O(gate500inter1));
  and2  gate1669(.a(G1263), .b(G1262), .O(gate500inter2));
  inv1  gate1670(.a(s_160), .O(gate500inter3));
  inv1  gate1671(.a(s_161), .O(gate500inter4));
  nand2 gate1672(.a(gate500inter4), .b(gate500inter3), .O(gate500inter5));
  nor2  gate1673(.a(gate500inter5), .b(gate500inter2), .O(gate500inter6));
  inv1  gate1674(.a(G1262), .O(gate500inter7));
  inv1  gate1675(.a(G1263), .O(gate500inter8));
  nand2 gate1676(.a(gate500inter8), .b(gate500inter7), .O(gate500inter9));
  nand2 gate1677(.a(s_161), .b(gate500inter3), .O(gate500inter10));
  nor2  gate1678(.a(gate500inter10), .b(gate500inter9), .O(gate500inter11));
  nor2  gate1679(.a(gate500inter11), .b(gate500inter6), .O(gate500inter12));
  nand2 gate1680(.a(gate500inter12), .b(gate500inter1), .O(G1309));
nand2 gate501( .a(G1264), .b(G1265), .O(G1310) );

  xor2  gate2535(.a(G1267), .b(G1266), .O(gate502inter0));
  nand2 gate2536(.a(gate502inter0), .b(s_284), .O(gate502inter1));
  and2  gate2537(.a(G1267), .b(G1266), .O(gate502inter2));
  inv1  gate2538(.a(s_284), .O(gate502inter3));
  inv1  gate2539(.a(s_285), .O(gate502inter4));
  nand2 gate2540(.a(gate502inter4), .b(gate502inter3), .O(gate502inter5));
  nor2  gate2541(.a(gate502inter5), .b(gate502inter2), .O(gate502inter6));
  inv1  gate2542(.a(G1266), .O(gate502inter7));
  inv1  gate2543(.a(G1267), .O(gate502inter8));
  nand2 gate2544(.a(gate502inter8), .b(gate502inter7), .O(gate502inter9));
  nand2 gate2545(.a(s_285), .b(gate502inter3), .O(gate502inter10));
  nor2  gate2546(.a(gate502inter10), .b(gate502inter9), .O(gate502inter11));
  nor2  gate2547(.a(gate502inter11), .b(gate502inter6), .O(gate502inter12));
  nand2 gate2548(.a(gate502inter12), .b(gate502inter1), .O(G1311));
nand2 gate503( .a(G1268), .b(G1269), .O(G1312) );
nand2 gate504( .a(G1270), .b(G1271), .O(G1313) );
nand2 gate505( .a(G1272), .b(G1273), .O(G1314) );
nand2 gate506( .a(G1274), .b(G1275), .O(G1315) );

  xor2  gate1625(.a(G1277), .b(G1276), .O(gate507inter0));
  nand2 gate1626(.a(gate507inter0), .b(s_154), .O(gate507inter1));
  and2  gate1627(.a(G1277), .b(G1276), .O(gate507inter2));
  inv1  gate1628(.a(s_154), .O(gate507inter3));
  inv1  gate1629(.a(s_155), .O(gate507inter4));
  nand2 gate1630(.a(gate507inter4), .b(gate507inter3), .O(gate507inter5));
  nor2  gate1631(.a(gate507inter5), .b(gate507inter2), .O(gate507inter6));
  inv1  gate1632(.a(G1276), .O(gate507inter7));
  inv1  gate1633(.a(G1277), .O(gate507inter8));
  nand2 gate1634(.a(gate507inter8), .b(gate507inter7), .O(gate507inter9));
  nand2 gate1635(.a(s_155), .b(gate507inter3), .O(gate507inter10));
  nor2  gate1636(.a(gate507inter10), .b(gate507inter9), .O(gate507inter11));
  nor2  gate1637(.a(gate507inter11), .b(gate507inter6), .O(gate507inter12));
  nand2 gate1638(.a(gate507inter12), .b(gate507inter1), .O(G1316));

  xor2  gate2031(.a(G1279), .b(G1278), .O(gate508inter0));
  nand2 gate2032(.a(gate508inter0), .b(s_212), .O(gate508inter1));
  and2  gate2033(.a(G1279), .b(G1278), .O(gate508inter2));
  inv1  gate2034(.a(s_212), .O(gate508inter3));
  inv1  gate2035(.a(s_213), .O(gate508inter4));
  nand2 gate2036(.a(gate508inter4), .b(gate508inter3), .O(gate508inter5));
  nor2  gate2037(.a(gate508inter5), .b(gate508inter2), .O(gate508inter6));
  inv1  gate2038(.a(G1278), .O(gate508inter7));
  inv1  gate2039(.a(G1279), .O(gate508inter8));
  nand2 gate2040(.a(gate508inter8), .b(gate508inter7), .O(gate508inter9));
  nand2 gate2041(.a(s_213), .b(gate508inter3), .O(gate508inter10));
  nor2  gate2042(.a(gate508inter10), .b(gate508inter9), .O(gate508inter11));
  nor2  gate2043(.a(gate508inter11), .b(gate508inter6), .O(gate508inter12));
  nand2 gate2044(.a(gate508inter12), .b(gate508inter1), .O(G1317));
nand2 gate509( .a(G1280), .b(G1281), .O(G1318) );
nand2 gate510( .a(G1282), .b(G1283), .O(G1319) );
nand2 gate511( .a(G1284), .b(G1285), .O(G1320) );

  xor2  gate1345(.a(G1287), .b(G1286), .O(gate512inter0));
  nand2 gate1346(.a(gate512inter0), .b(s_114), .O(gate512inter1));
  and2  gate1347(.a(G1287), .b(G1286), .O(gate512inter2));
  inv1  gate1348(.a(s_114), .O(gate512inter3));
  inv1  gate1349(.a(s_115), .O(gate512inter4));
  nand2 gate1350(.a(gate512inter4), .b(gate512inter3), .O(gate512inter5));
  nor2  gate1351(.a(gate512inter5), .b(gate512inter2), .O(gate512inter6));
  inv1  gate1352(.a(G1286), .O(gate512inter7));
  inv1  gate1353(.a(G1287), .O(gate512inter8));
  nand2 gate1354(.a(gate512inter8), .b(gate512inter7), .O(gate512inter9));
  nand2 gate1355(.a(s_115), .b(gate512inter3), .O(gate512inter10));
  nor2  gate1356(.a(gate512inter10), .b(gate512inter9), .O(gate512inter11));
  nor2  gate1357(.a(gate512inter11), .b(gate512inter6), .O(gate512inter12));
  nand2 gate1358(.a(gate512inter12), .b(gate512inter1), .O(G1321));
nand2 gate513( .a(G1288), .b(G1289), .O(G1322) );
nand2 gate514( .a(G1290), .b(G1291), .O(G1323) );
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule