module c499 (N1,N5,N9,N13,N17,N21,N25,N29,N33,N37,
             N41,N45,N49,N53,N57,N61,N65,N69,N73,N77,
             N81,N85,N89,N93,N97,N101,N105,N109,N113,N117,
             N121,N125,N129,N130,N131,N132,N133,N134,N135,N136,
             N137,N724,N725,N726,N727,N728,N729,N730,N731,N732,
             N733,N734,N735,N736,N737,N738,N739,N740,N741,N742,
             N743,N744,N745,N746,N747,N748,N749,N750,N751,N752,
             N753,N754,N755);

input N1,N5,N9,N13,N17,N21,N25,N29,N33,N37,
      N41,N45,N49,N53,N57,N61,N65,N69,N73,N77,
      N81,N85,N89,N93,N97,N101,N105,N109,N113,N117,
      N121,N125,N129,N130,N131,N132,N133,N134,N135,N136,
      N137;//RE__PI;

input s_0,s_1;//RE__ALLOW(00,01,10,11);
input s_2,s_3;//RE__ALLOW(00,01,10,11);
input s_4,s_5;//RE__ALLOW(00,01,10,11);
input s_6,s_7;//RE__ALLOW(00,01,10,11);
input s_8,s_9;//RE__ALLOW(00,01,10,11);
input s_10,s_11;//RE__ALLOW(00,01,10,11);
input s_12,s_13;//RE__ALLOW(00,01,10,11);
input s_14,s_15;//RE__ALLOW(00,01,10,11);
input s_16,s_17;//RE__ALLOW(00,01,10,11);
input s_18,s_19;//RE__ALLOW(00,01,10,11);
input s_20,s_21;//RE__ALLOW(00,01,10,11);
input s_22,s_23;//RE__ALLOW(00,01,10,11);
input s_24,s_25;//RE__ALLOW(00,01,10,11);
input s_26,s_27;//RE__ALLOW(00,01,10,11);
input s_28,s_29;//RE__ALLOW(00,01,10,11);
input s_30,s_31;//RE__ALLOW(00,01,10,11);
input s_32,s_33;//RE__ALLOW(00,01,10,11);
input s_34,s_35;//RE__ALLOW(00,01,10,11);
input s_36,s_37;//RE__ALLOW(00,01,10,11);
input s_38,s_39;//RE__ALLOW(00,01,10,11);
input s_40,s_41;//RE__ALLOW(00,01,10,11);
output N724,N725,N726,N727,N728,N729,N730,N731,N732,N733,
       N734,N735,N736,N737,N738,N739,N740,N741,N742,N743,
       N744,N745,N746,N747,N748,N749,N750,N751,N752,N753,
       N754,N755;

wire N250,N251,N252,N253,N254,N255,N256,N257,N258,N259,
     N260,N261,N262,N263,N264,N265,N266,N267,N268,N269,
     N270,N271,N272,N273,N274,N275,N276,N277,N278,N279,
     N280,N281,N282,N283,N284,N285,N286,N287,N288,N289,
     N290,N293,N296,N299,N302,N305,N308,N311,N314,N315,
     N316,N317,N318,N319,N320,N321,N338,N339,N340,N341,
     N342,N343,N344,N345,N346,N347,N348,N349,N350,N351,
     N352,N353,N354,N367,N380,N393,N406,N419,N432,N445,
     N554,N555,N556,N557,N558,N559,N560,N561,N562,N563,
     N564,N565,N566,N567,N568,N569,N570,N571,N572,N573,
     N574,N575,N576,N577,N578,N579,N580,N581,N582,N583,
     N584,N585,N586,N587,N588,N589,N590,N591,N592,N593,
     N594,N595,N596,N597,N598,N599,N600,N601,N602,N607,
     N620,N625,N630,N635,N640,N645,N650,N655,N692,N693,
     N694,N695,N696,N697,N698,N699,N700,N701,N702,N703,
     N704,N705,N706,N707,N708,N709,N710,N711,N712,N713,
     N714,N715,N716,N717,N718,N719,N720,N721,N722,N723, gate181inter0, gate181inter1, gate181inter2, gate181inter3, gate181inter4, gate181inter5, gate181inter6, gate181inter7, gate181inter8, gate181inter9, gate181inter10, gate181inter11, gate181inter12, gate192inter0, gate192inter1, gate192inter2, gate192inter3, gate192inter4, gate192inter5, gate192inter6, gate192inter7, gate192inter8, gate192inter9, gate192inter10, gate192inter11, gate192inter12, gate47inter0, gate47inter1, gate47inter2, gate47inter3, gate47inter4, gate47inter5, gate47inter6, gate47inter7, gate47inter8, gate47inter9, gate47inter10, gate47inter11, gate47inter12, gate180inter0, gate180inter1, gate180inter2, gate180inter3, gate180inter4, gate180inter5, gate180inter6, gate180inter7, gate180inter8, gate180inter9, gate180inter10, gate180inter11, gate180inter12, gate33inter0, gate33inter1, gate33inter2, gate33inter3, gate33inter4, gate33inter5, gate33inter6, gate33inter7, gate33inter8, gate33inter9, gate33inter10, gate33inter11, gate33inter12, gate174inter0, gate174inter1, gate174inter2, gate174inter3, gate174inter4, gate174inter5, gate174inter6, gate174inter7, gate174inter8, gate174inter9, gate174inter10, gate174inter11, gate174inter12, gate41inter0, gate41inter1, gate41inter2, gate41inter3, gate41inter4, gate41inter5, gate41inter6, gate41inter7, gate41inter8, gate41inter9, gate41inter10, gate41inter11, gate41inter12, gate26inter0, gate26inter1, gate26inter2, gate26inter3, gate26inter4, gate26inter5, gate26inter6, gate26inter7, gate26inter8, gate26inter9, gate26inter10, gate26inter11, gate26inter12, gate50inter0, gate50inter1, gate50inter2, gate50inter3, gate50inter4, gate50inter5, gate50inter6, gate50inter7, gate50inter8, gate50inter9, gate50inter10, gate50inter11, gate50inter12, gate15inter0, gate15inter1, gate15inter2, gate15inter3, gate15inter4, gate15inter5, gate15inter6, gate15inter7, gate15inter8, gate15inter9, gate15inter10, gate15inter11, gate15inter12, gate51inter0, gate51inter1, gate51inter2, gate51inter3, gate51inter4, gate51inter5, gate51inter6, gate51inter7, gate51inter8, gate51inter9, gate51inter10, gate51inter11, gate51inter12, gate188inter0, gate188inter1, gate188inter2, gate188inter3, gate188inter4, gate188inter5, gate188inter6, gate188inter7, gate188inter8, gate188inter9, gate188inter10, gate188inter11, gate188inter12, gate172inter0, gate172inter1, gate172inter2, gate172inter3, gate172inter4, gate172inter5, gate172inter6, gate172inter7, gate172inter8, gate172inter9, gate172inter10, gate172inter11, gate172inter12, gate13inter0, gate13inter1, gate13inter2, gate13inter3, gate13inter4, gate13inter5, gate13inter6, gate13inter7, gate13inter8, gate13inter9, gate13inter10, gate13inter11, gate13inter12, gate56inter0, gate56inter1, gate56inter2, gate56inter3, gate56inter4, gate56inter5, gate56inter6, gate56inter7, gate56inter8, gate56inter9, gate56inter10, gate56inter11, gate56inter12, gate185inter0, gate185inter1, gate185inter2, gate185inter3, gate185inter4, gate185inter5, gate185inter6, gate185inter7, gate185inter8, gate185inter9, gate185inter10, gate185inter11, gate185inter12, gate78inter0, gate78inter1, gate78inter2, gate78inter3, gate78inter4, gate78inter5, gate78inter6, gate78inter7, gate78inter8, gate78inter9, gate78inter10, gate78inter11, gate78inter12, gate48inter0, gate48inter1, gate48inter2, gate48inter3, gate48inter4, gate48inter5, gate48inter6, gate48inter7, gate48inter8, gate48inter9, gate48inter10, gate48inter11, gate48inter12, gate52inter0, gate52inter1, gate52inter2, gate52inter3, gate52inter4, gate52inter5, gate52inter6, gate52inter7, gate52inter8, gate52inter9, gate52inter10, gate52inter11, gate52inter12, gate49inter0, gate49inter1, gate49inter2, gate49inter3, gate49inter4, gate49inter5, gate49inter6, gate49inter7, gate49inter8, gate49inter9, gate49inter10, gate49inter11, gate49inter12, gate75inter0, gate75inter1, gate75inter2, gate75inter3, gate75inter4, gate75inter5, gate75inter6, gate75inter7, gate75inter8, gate75inter9, gate75inter10, gate75inter11, gate75inter12;



xor2 gate1( .a(N1), .b(N5), .O(N250) );
xor2 gate2( .a(N9), .b(N13), .O(N251) );
xor2 gate3( .a(N17), .b(N21), .O(N252) );
xor2 gate4( .a(N25), .b(N29), .O(N253) );
xor2 gate5( .a(N33), .b(N37), .O(N254) );
xor2 gate6( .a(N41), .b(N45), .O(N255) );
xor2 gate7( .a(N49), .b(N53), .O(N256) );
xor2 gate8( .a(N57), .b(N61), .O(N257) );
xor2 gate9( .a(N65), .b(N69), .O(N258) );
xor2 gate10( .a(N73), .b(N77), .O(N259) );
xor2 gate11( .a(N81), .b(N85), .O(N260) );
xor2 gate12( .a(N89), .b(N93), .O(N261) );

  xor2  gate385(.a(N101), .b(N97), .O(gate13inter0));
  nand2 gate386(.a(gate13inter0), .b(s_26), .O(gate13inter1));
  and2  gate387(.a(N101), .b(N97), .O(gate13inter2));
  inv1  gate388(.a(s_26), .O(gate13inter3));
  inv1  gate389(.a(s_27), .O(gate13inter4));
  nand2 gate390(.a(gate13inter4), .b(gate13inter3), .O(gate13inter5));
  nor2  gate391(.a(gate13inter5), .b(gate13inter2), .O(gate13inter6));
  inv1  gate392(.a(N97), .O(gate13inter7));
  inv1  gate393(.a(N101), .O(gate13inter8));
  nand2 gate394(.a(gate13inter8), .b(gate13inter7), .O(gate13inter9));
  nand2 gate395(.a(s_27), .b(gate13inter3), .O(gate13inter10));
  nor2  gate396(.a(gate13inter10), .b(gate13inter9), .O(gate13inter11));
  nor2  gate397(.a(gate13inter11), .b(gate13inter6), .O(gate13inter12));
  nand2 gate398(.a(gate13inter12), .b(gate13inter1), .O(N262));
xor2 gate14( .a(N105), .b(N109), .O(N263) );

  xor2  gate329(.a(N117), .b(N113), .O(gate15inter0));
  nand2 gate330(.a(gate15inter0), .b(s_18), .O(gate15inter1));
  and2  gate331(.a(N117), .b(N113), .O(gate15inter2));
  inv1  gate332(.a(s_18), .O(gate15inter3));
  inv1  gate333(.a(s_19), .O(gate15inter4));
  nand2 gate334(.a(gate15inter4), .b(gate15inter3), .O(gate15inter5));
  nor2  gate335(.a(gate15inter5), .b(gate15inter2), .O(gate15inter6));
  inv1  gate336(.a(N113), .O(gate15inter7));
  inv1  gate337(.a(N117), .O(gate15inter8));
  nand2 gate338(.a(gate15inter8), .b(gate15inter7), .O(gate15inter9));
  nand2 gate339(.a(s_19), .b(gate15inter3), .O(gate15inter10));
  nor2  gate340(.a(gate15inter10), .b(gate15inter9), .O(gate15inter11));
  nor2  gate341(.a(gate15inter11), .b(gate15inter6), .O(gate15inter12));
  nand2 gate342(.a(gate15inter12), .b(gate15inter1), .O(N264));
xor2 gate16( .a(N121), .b(N125), .O(N265) );
and2 gate17( .a(N129), .b(N137), .O(N266) );
and2 gate18( .a(N130), .b(N137), .O(N267) );
and2 gate19( .a(N131), .b(N137), .O(N268) );
and2 gate20( .a(N132), .b(N137), .O(N269) );
and2 gate21( .a(N133), .b(N137), .O(N270) );
and2 gate22( .a(N134), .b(N137), .O(N271) );
and2 gate23( .a(N135), .b(N137), .O(N272) );
and2 gate24( .a(N136), .b(N137), .O(N273) );
xor2 gate25( .a(N1), .b(N17), .O(N274) );

  xor2  gate301(.a(N49), .b(N33), .O(gate26inter0));
  nand2 gate302(.a(gate26inter0), .b(s_14), .O(gate26inter1));
  and2  gate303(.a(N49), .b(N33), .O(gate26inter2));
  inv1  gate304(.a(s_14), .O(gate26inter3));
  inv1  gate305(.a(s_15), .O(gate26inter4));
  nand2 gate306(.a(gate26inter4), .b(gate26inter3), .O(gate26inter5));
  nor2  gate307(.a(gate26inter5), .b(gate26inter2), .O(gate26inter6));
  inv1  gate308(.a(N33), .O(gate26inter7));
  inv1  gate309(.a(N49), .O(gate26inter8));
  nand2 gate310(.a(gate26inter8), .b(gate26inter7), .O(gate26inter9));
  nand2 gate311(.a(s_15), .b(gate26inter3), .O(gate26inter10));
  nor2  gate312(.a(gate26inter10), .b(gate26inter9), .O(gate26inter11));
  nor2  gate313(.a(gate26inter11), .b(gate26inter6), .O(gate26inter12));
  nand2 gate314(.a(gate26inter12), .b(gate26inter1), .O(N275));
xor2 gate27( .a(N5), .b(N21), .O(N276) );
xor2 gate28( .a(N37), .b(N53), .O(N277) );
xor2 gate29( .a(N9), .b(N25), .O(N278) );
xor2 gate30( .a(N41), .b(N57), .O(N279) );
xor2 gate31( .a(N13), .b(N29), .O(N280) );
xor2 gate32( .a(N45), .b(N61), .O(N281) );

  xor2  gate259(.a(N81), .b(N65), .O(gate33inter0));
  nand2 gate260(.a(gate33inter0), .b(s_8), .O(gate33inter1));
  and2  gate261(.a(N81), .b(N65), .O(gate33inter2));
  inv1  gate262(.a(s_8), .O(gate33inter3));
  inv1  gate263(.a(s_9), .O(gate33inter4));
  nand2 gate264(.a(gate33inter4), .b(gate33inter3), .O(gate33inter5));
  nor2  gate265(.a(gate33inter5), .b(gate33inter2), .O(gate33inter6));
  inv1  gate266(.a(N65), .O(gate33inter7));
  inv1  gate267(.a(N81), .O(gate33inter8));
  nand2 gate268(.a(gate33inter8), .b(gate33inter7), .O(gate33inter9));
  nand2 gate269(.a(s_9), .b(gate33inter3), .O(gate33inter10));
  nor2  gate270(.a(gate33inter10), .b(gate33inter9), .O(gate33inter11));
  nor2  gate271(.a(gate33inter11), .b(gate33inter6), .O(gate33inter12));
  nand2 gate272(.a(gate33inter12), .b(gate33inter1), .O(N282));
xor2 gate34( .a(N97), .b(N113), .O(N283) );
xor2 gate35( .a(N69), .b(N85), .O(N284) );
xor2 gate36( .a(N101), .b(N117), .O(N285) );
xor2 gate37( .a(N73), .b(N89), .O(N286) );
xor2 gate38( .a(N105), .b(N121), .O(N287) );
xor2 gate39( .a(N77), .b(N93), .O(N288) );
xor2 gate40( .a(N109), .b(N125), .O(N289) );

  xor2  gate287(.a(N251), .b(N250), .O(gate41inter0));
  nand2 gate288(.a(gate41inter0), .b(s_12), .O(gate41inter1));
  and2  gate289(.a(N251), .b(N250), .O(gate41inter2));
  inv1  gate290(.a(s_12), .O(gate41inter3));
  inv1  gate291(.a(s_13), .O(gate41inter4));
  nand2 gate292(.a(gate41inter4), .b(gate41inter3), .O(gate41inter5));
  nor2  gate293(.a(gate41inter5), .b(gate41inter2), .O(gate41inter6));
  inv1  gate294(.a(N250), .O(gate41inter7));
  inv1  gate295(.a(N251), .O(gate41inter8));
  nand2 gate296(.a(gate41inter8), .b(gate41inter7), .O(gate41inter9));
  nand2 gate297(.a(s_13), .b(gate41inter3), .O(gate41inter10));
  nor2  gate298(.a(gate41inter10), .b(gate41inter9), .O(gate41inter11));
  nor2  gate299(.a(gate41inter11), .b(gate41inter6), .O(gate41inter12));
  nand2 gate300(.a(gate41inter12), .b(gate41inter1), .O(N290));
xor2 gate42( .a(N252), .b(N253), .O(N293) );
xor2 gate43( .a(N254), .b(N255), .O(N296) );
xor2 gate44( .a(N256), .b(N257), .O(N299) );
xor2 gate45( .a(N258), .b(N259), .O(N302) );
xor2 gate46( .a(N260), .b(N261), .O(N305) );

  xor2  gate231(.a(N263), .b(N262), .O(gate47inter0));
  nand2 gate232(.a(gate47inter0), .b(s_4), .O(gate47inter1));
  and2  gate233(.a(N263), .b(N262), .O(gate47inter2));
  inv1  gate234(.a(s_4), .O(gate47inter3));
  inv1  gate235(.a(s_5), .O(gate47inter4));
  nand2 gate236(.a(gate47inter4), .b(gate47inter3), .O(gate47inter5));
  nor2  gate237(.a(gate47inter5), .b(gate47inter2), .O(gate47inter6));
  inv1  gate238(.a(N262), .O(gate47inter7));
  inv1  gate239(.a(N263), .O(gate47inter8));
  nand2 gate240(.a(gate47inter8), .b(gate47inter7), .O(gate47inter9));
  nand2 gate241(.a(s_5), .b(gate47inter3), .O(gate47inter10));
  nor2  gate242(.a(gate47inter10), .b(gate47inter9), .O(gate47inter11));
  nor2  gate243(.a(gate47inter11), .b(gate47inter6), .O(gate47inter12));
  nand2 gate244(.a(gate47inter12), .b(gate47inter1), .O(N308));

  xor2  gate441(.a(N265), .b(N264), .O(gate48inter0));
  nand2 gate442(.a(gate48inter0), .b(s_34), .O(gate48inter1));
  and2  gate443(.a(N265), .b(N264), .O(gate48inter2));
  inv1  gate444(.a(s_34), .O(gate48inter3));
  inv1  gate445(.a(s_35), .O(gate48inter4));
  nand2 gate446(.a(gate48inter4), .b(gate48inter3), .O(gate48inter5));
  nor2  gate447(.a(gate48inter5), .b(gate48inter2), .O(gate48inter6));
  inv1  gate448(.a(N264), .O(gate48inter7));
  inv1  gate449(.a(N265), .O(gate48inter8));
  nand2 gate450(.a(gate48inter8), .b(gate48inter7), .O(gate48inter9));
  nand2 gate451(.a(s_35), .b(gate48inter3), .O(gate48inter10));
  nor2  gate452(.a(gate48inter10), .b(gate48inter9), .O(gate48inter11));
  nor2  gate453(.a(gate48inter11), .b(gate48inter6), .O(gate48inter12));
  nand2 gate454(.a(gate48inter12), .b(gate48inter1), .O(N311));

  xor2  gate469(.a(N275), .b(N274), .O(gate49inter0));
  nand2 gate470(.a(gate49inter0), .b(s_38), .O(gate49inter1));
  and2  gate471(.a(N275), .b(N274), .O(gate49inter2));
  inv1  gate472(.a(s_38), .O(gate49inter3));
  inv1  gate473(.a(s_39), .O(gate49inter4));
  nand2 gate474(.a(gate49inter4), .b(gate49inter3), .O(gate49inter5));
  nor2  gate475(.a(gate49inter5), .b(gate49inter2), .O(gate49inter6));
  inv1  gate476(.a(N274), .O(gate49inter7));
  inv1  gate477(.a(N275), .O(gate49inter8));
  nand2 gate478(.a(gate49inter8), .b(gate49inter7), .O(gate49inter9));
  nand2 gate479(.a(s_39), .b(gate49inter3), .O(gate49inter10));
  nor2  gate480(.a(gate49inter10), .b(gate49inter9), .O(gate49inter11));
  nor2  gate481(.a(gate49inter11), .b(gate49inter6), .O(gate49inter12));
  nand2 gate482(.a(gate49inter12), .b(gate49inter1), .O(N314));

  xor2  gate315(.a(N277), .b(N276), .O(gate50inter0));
  nand2 gate316(.a(gate50inter0), .b(s_16), .O(gate50inter1));
  and2  gate317(.a(N277), .b(N276), .O(gate50inter2));
  inv1  gate318(.a(s_16), .O(gate50inter3));
  inv1  gate319(.a(s_17), .O(gate50inter4));
  nand2 gate320(.a(gate50inter4), .b(gate50inter3), .O(gate50inter5));
  nor2  gate321(.a(gate50inter5), .b(gate50inter2), .O(gate50inter6));
  inv1  gate322(.a(N276), .O(gate50inter7));
  inv1  gate323(.a(N277), .O(gate50inter8));
  nand2 gate324(.a(gate50inter8), .b(gate50inter7), .O(gate50inter9));
  nand2 gate325(.a(s_17), .b(gate50inter3), .O(gate50inter10));
  nor2  gate326(.a(gate50inter10), .b(gate50inter9), .O(gate50inter11));
  nor2  gate327(.a(gate50inter11), .b(gate50inter6), .O(gate50inter12));
  nand2 gate328(.a(gate50inter12), .b(gate50inter1), .O(N315));

  xor2  gate343(.a(N279), .b(N278), .O(gate51inter0));
  nand2 gate344(.a(gate51inter0), .b(s_20), .O(gate51inter1));
  and2  gate345(.a(N279), .b(N278), .O(gate51inter2));
  inv1  gate346(.a(s_20), .O(gate51inter3));
  inv1  gate347(.a(s_21), .O(gate51inter4));
  nand2 gate348(.a(gate51inter4), .b(gate51inter3), .O(gate51inter5));
  nor2  gate349(.a(gate51inter5), .b(gate51inter2), .O(gate51inter6));
  inv1  gate350(.a(N278), .O(gate51inter7));
  inv1  gate351(.a(N279), .O(gate51inter8));
  nand2 gate352(.a(gate51inter8), .b(gate51inter7), .O(gate51inter9));
  nand2 gate353(.a(s_21), .b(gate51inter3), .O(gate51inter10));
  nor2  gate354(.a(gate51inter10), .b(gate51inter9), .O(gate51inter11));
  nor2  gate355(.a(gate51inter11), .b(gate51inter6), .O(gate51inter12));
  nand2 gate356(.a(gate51inter12), .b(gate51inter1), .O(N316));

  xor2  gate455(.a(N281), .b(N280), .O(gate52inter0));
  nand2 gate456(.a(gate52inter0), .b(s_36), .O(gate52inter1));
  and2  gate457(.a(N281), .b(N280), .O(gate52inter2));
  inv1  gate458(.a(s_36), .O(gate52inter3));
  inv1  gate459(.a(s_37), .O(gate52inter4));
  nand2 gate460(.a(gate52inter4), .b(gate52inter3), .O(gate52inter5));
  nor2  gate461(.a(gate52inter5), .b(gate52inter2), .O(gate52inter6));
  inv1  gate462(.a(N280), .O(gate52inter7));
  inv1  gate463(.a(N281), .O(gate52inter8));
  nand2 gate464(.a(gate52inter8), .b(gate52inter7), .O(gate52inter9));
  nand2 gate465(.a(s_37), .b(gate52inter3), .O(gate52inter10));
  nor2  gate466(.a(gate52inter10), .b(gate52inter9), .O(gate52inter11));
  nor2  gate467(.a(gate52inter11), .b(gate52inter6), .O(gate52inter12));
  nand2 gate468(.a(gate52inter12), .b(gate52inter1), .O(N317));
xor2 gate53( .a(N282), .b(N283), .O(N318) );
xor2 gate54( .a(N284), .b(N285), .O(N319) );
xor2 gate55( .a(N286), .b(N287), .O(N320) );

  xor2  gate399(.a(N289), .b(N288), .O(gate56inter0));
  nand2 gate400(.a(gate56inter0), .b(s_28), .O(gate56inter1));
  and2  gate401(.a(N289), .b(N288), .O(gate56inter2));
  inv1  gate402(.a(s_28), .O(gate56inter3));
  inv1  gate403(.a(s_29), .O(gate56inter4));
  nand2 gate404(.a(gate56inter4), .b(gate56inter3), .O(gate56inter5));
  nor2  gate405(.a(gate56inter5), .b(gate56inter2), .O(gate56inter6));
  inv1  gate406(.a(N288), .O(gate56inter7));
  inv1  gate407(.a(N289), .O(gate56inter8));
  nand2 gate408(.a(gate56inter8), .b(gate56inter7), .O(gate56inter9));
  nand2 gate409(.a(s_29), .b(gate56inter3), .O(gate56inter10));
  nor2  gate410(.a(gate56inter10), .b(gate56inter9), .O(gate56inter11));
  nor2  gate411(.a(gate56inter11), .b(gate56inter6), .O(gate56inter12));
  nand2 gate412(.a(gate56inter12), .b(gate56inter1), .O(N321));
xor2 gate57( .a(N290), .b(N293), .O(N338) );
xor2 gate58( .a(N296), .b(N299), .O(N339) );
xor2 gate59( .a(N290), .b(N296), .O(N340) );
xor2 gate60( .a(N293), .b(N299), .O(N341) );
xor2 gate61( .a(N302), .b(N305), .O(N342) );
xor2 gate62( .a(N308), .b(N311), .O(N343) );
xor2 gate63( .a(N302), .b(N308), .O(N344) );
xor2 gate64( .a(N305), .b(N311), .O(N345) );
xor2 gate65( .a(N266), .b(N342), .O(N346) );
xor2 gate66( .a(N267), .b(N343), .O(N347) );
xor2 gate67( .a(N268), .b(N344), .O(N348) );
xor2 gate68( .a(N269), .b(N345), .O(N349) );
xor2 gate69( .a(N270), .b(N338), .O(N350) );
xor2 gate70( .a(N271), .b(N339), .O(N351) );
xor2 gate71( .a(N272), .b(N340), .O(N352) );
xor2 gate72( .a(N273), .b(N341), .O(N353) );
xor2 gate73( .a(N314), .b(N346), .O(N354) );
xor2 gate74( .a(N315), .b(N347), .O(N367) );

  xor2  gate483(.a(N348), .b(N316), .O(gate75inter0));
  nand2 gate484(.a(gate75inter0), .b(s_40), .O(gate75inter1));
  and2  gate485(.a(N348), .b(N316), .O(gate75inter2));
  inv1  gate486(.a(s_40), .O(gate75inter3));
  inv1  gate487(.a(s_41), .O(gate75inter4));
  nand2 gate488(.a(gate75inter4), .b(gate75inter3), .O(gate75inter5));
  nor2  gate489(.a(gate75inter5), .b(gate75inter2), .O(gate75inter6));
  inv1  gate490(.a(N316), .O(gate75inter7));
  inv1  gate491(.a(N348), .O(gate75inter8));
  nand2 gate492(.a(gate75inter8), .b(gate75inter7), .O(gate75inter9));
  nand2 gate493(.a(s_41), .b(gate75inter3), .O(gate75inter10));
  nor2  gate494(.a(gate75inter10), .b(gate75inter9), .O(gate75inter11));
  nor2  gate495(.a(gate75inter11), .b(gate75inter6), .O(gate75inter12));
  nand2 gate496(.a(gate75inter12), .b(gate75inter1), .O(N380));
xor2 gate76( .a(N317), .b(N349), .O(N393) );
xor2 gate77( .a(N318), .b(N350), .O(N406) );

  xor2  gate427(.a(N351), .b(N319), .O(gate78inter0));
  nand2 gate428(.a(gate78inter0), .b(s_32), .O(gate78inter1));
  and2  gate429(.a(N351), .b(N319), .O(gate78inter2));
  inv1  gate430(.a(s_32), .O(gate78inter3));
  inv1  gate431(.a(s_33), .O(gate78inter4));
  nand2 gate432(.a(gate78inter4), .b(gate78inter3), .O(gate78inter5));
  nor2  gate433(.a(gate78inter5), .b(gate78inter2), .O(gate78inter6));
  inv1  gate434(.a(N319), .O(gate78inter7));
  inv1  gate435(.a(N351), .O(gate78inter8));
  nand2 gate436(.a(gate78inter8), .b(gate78inter7), .O(gate78inter9));
  nand2 gate437(.a(s_33), .b(gate78inter3), .O(gate78inter10));
  nor2  gate438(.a(gate78inter10), .b(gate78inter9), .O(gate78inter11));
  nor2  gate439(.a(gate78inter11), .b(gate78inter6), .O(gate78inter12));
  nand2 gate440(.a(gate78inter12), .b(gate78inter1), .O(N419));
xor2 gate79( .a(N320), .b(N352), .O(N432) );
xor2 gate80( .a(N321), .b(N353), .O(N445) );
inv1 gate81( .a(N354), .O(N554) );
inv1 gate82( .a(N367), .O(N555) );
inv1 gate83( .a(N380), .O(N556) );
inv1 gate84( .a(N354), .O(N557) );
inv1 gate85( .a(N367), .O(N558) );
inv1 gate86( .a(N393), .O(N559) );
inv1 gate87( .a(N354), .O(N560) );
inv1 gate88( .a(N380), .O(N561) );
inv1 gate89( .a(N393), .O(N562) );
inv1 gate90( .a(N367), .O(N563) );
inv1 gate91( .a(N380), .O(N564) );
inv1 gate92( .a(N393), .O(N565) );
inv1 gate93( .a(N419), .O(N566) );
inv1 gate94( .a(N445), .O(N567) );
inv1 gate95( .a(N419), .O(N568) );
inv1 gate96( .a(N432), .O(N569) );
inv1 gate97( .a(N406), .O(N570) );
inv1 gate98( .a(N445), .O(N571) );
inv1 gate99( .a(N406), .O(N572) );
inv1 gate100( .a(N432), .O(N573) );
inv1 gate101( .a(N406), .O(N574) );
inv1 gate102( .a(N419), .O(N575) );
inv1 gate103( .a(N432), .O(N576) );
inv1 gate104( .a(N406), .O(N577) );
inv1 gate105( .a(N419), .O(N578) );
inv1 gate106( .a(N445), .O(N579) );
inv1 gate107( .a(N406), .O(N580) );
inv1 gate108( .a(N432), .O(N581) );
inv1 gate109( .a(N445), .O(N582) );
inv1 gate110( .a(N419), .O(N583) );
inv1 gate111( .a(N432), .O(N584) );
inv1 gate112( .a(N445), .O(N585) );
inv1 gate113( .a(N367), .O(N586) );
inv1 gate114( .a(N393), .O(N587) );
inv1 gate115( .a(N367), .O(N588) );
inv1 gate116( .a(N380), .O(N589) );
inv1 gate117( .a(N354), .O(N590) );
inv1 gate118( .a(N393), .O(N591) );
inv1 gate119( .a(N354), .O(N592) );
inv1 gate120( .a(N380), .O(N593) );
and4 gate121( .a(N554), .b(N555), .c(N556), .d(N393), .O(N594) );
and4 gate122( .a(N557), .b(N558), .c(N380), .d(N559), .O(N595) );
and4 gate123( .a(N560), .b(N367), .c(N561), .d(N562), .O(N596) );
and4 gate124( .a(N354), .b(N563), .c(N564), .d(N565), .O(N597) );
and4 gate125( .a(N574), .b(N575), .c(N576), .d(N445), .O(N598) );
and4 gate126( .a(N577), .b(N578), .c(N432), .d(N579), .O(N599) );
and4 gate127( .a(N580), .b(N419), .c(N581), .d(N582), .O(N600) );
and4 gate128( .a(N406), .b(N583), .c(N584), .d(N585), .O(N601) );
or4 gate129( .a(N594), .b(N595), .c(N596), .d(N597), .O(N602) );
or4 gate130( .a(N598), .b(N599), .c(N600), .d(N601), .O(N607) );
and5 gate131( .a(N406), .b(N566), .c(N432), .d(N567), .e(N602), .O(N620) );
and5 gate132( .a(N406), .b(N568), .c(N569), .d(N445), .e(N602), .O(N625) );
and5 gate133( .a(N570), .b(N419), .c(N432), .d(N571), .e(N602), .O(N630) );
and5 gate134( .a(N572), .b(N419), .c(N573), .d(N445), .e(N602), .O(N635) );
and5 gate135( .a(N354), .b(N586), .c(N380), .d(N587), .e(N607), .O(N640) );
and5 gate136( .a(N354), .b(N588), .c(N589), .d(N393), .e(N607), .O(N645) );
and5 gate137( .a(N590), .b(N367), .c(N380), .d(N591), .e(N607), .O(N650) );
and5 gate138( .a(N592), .b(N367), .c(N593), .d(N393), .e(N607), .O(N655) );
and2 gate139( .a(N354), .b(N620), .O(N692) );
and2 gate140( .a(N367), .b(N620), .O(N693) );
and2 gate141( .a(N380), .b(N620), .O(N694) );
and2 gate142( .a(N393), .b(N620), .O(N695) );
and2 gate143( .a(N354), .b(N625), .O(N696) );
and2 gate144( .a(N367), .b(N625), .O(N697) );
and2 gate145( .a(N380), .b(N625), .O(N698) );
and2 gate146( .a(N393), .b(N625), .O(N699) );
and2 gate147( .a(N354), .b(N630), .O(N700) );
and2 gate148( .a(N367), .b(N630), .O(N701) );
and2 gate149( .a(N380), .b(N630), .O(N702) );
and2 gate150( .a(N393), .b(N630), .O(N703) );
and2 gate151( .a(N354), .b(N635), .O(N704) );
and2 gate152( .a(N367), .b(N635), .O(N705) );
and2 gate153( .a(N380), .b(N635), .O(N706) );
and2 gate154( .a(N393), .b(N635), .O(N707) );
and2 gate155( .a(N406), .b(N640), .O(N708) );
and2 gate156( .a(N419), .b(N640), .O(N709) );
and2 gate157( .a(N432), .b(N640), .O(N710) );
and2 gate158( .a(N445), .b(N640), .O(N711) );
and2 gate159( .a(N406), .b(N645), .O(N712) );
and2 gate160( .a(N419), .b(N645), .O(N713) );
and2 gate161( .a(N432), .b(N645), .O(N714) );
and2 gate162( .a(N445), .b(N645), .O(N715) );
and2 gate163( .a(N406), .b(N650), .O(N716) );
and2 gate164( .a(N419), .b(N650), .O(N717) );
and2 gate165( .a(N432), .b(N650), .O(N718) );
and2 gate166( .a(N445), .b(N650), .O(N719) );
and2 gate167( .a(N406), .b(N655), .O(N720) );
and2 gate168( .a(N419), .b(N655), .O(N721) );
and2 gate169( .a(N432), .b(N655), .O(N722) );
and2 gate170( .a(N445), .b(N655), .O(N723) );
xor2 gate171( .a(N1), .b(N692), .O(N724) );

  xor2  gate371(.a(N693), .b(N5), .O(gate172inter0));
  nand2 gate372(.a(gate172inter0), .b(s_24), .O(gate172inter1));
  and2  gate373(.a(N693), .b(N5), .O(gate172inter2));
  inv1  gate374(.a(s_24), .O(gate172inter3));
  inv1  gate375(.a(s_25), .O(gate172inter4));
  nand2 gate376(.a(gate172inter4), .b(gate172inter3), .O(gate172inter5));
  nor2  gate377(.a(gate172inter5), .b(gate172inter2), .O(gate172inter6));
  inv1  gate378(.a(N5), .O(gate172inter7));
  inv1  gate379(.a(N693), .O(gate172inter8));
  nand2 gate380(.a(gate172inter8), .b(gate172inter7), .O(gate172inter9));
  nand2 gate381(.a(s_25), .b(gate172inter3), .O(gate172inter10));
  nor2  gate382(.a(gate172inter10), .b(gate172inter9), .O(gate172inter11));
  nor2  gate383(.a(gate172inter11), .b(gate172inter6), .O(gate172inter12));
  nand2 gate384(.a(gate172inter12), .b(gate172inter1), .O(N725));
xor2 gate173( .a(N9), .b(N694), .O(N726) );

  xor2  gate273(.a(N695), .b(N13), .O(gate174inter0));
  nand2 gate274(.a(gate174inter0), .b(s_10), .O(gate174inter1));
  and2  gate275(.a(N695), .b(N13), .O(gate174inter2));
  inv1  gate276(.a(s_10), .O(gate174inter3));
  inv1  gate277(.a(s_11), .O(gate174inter4));
  nand2 gate278(.a(gate174inter4), .b(gate174inter3), .O(gate174inter5));
  nor2  gate279(.a(gate174inter5), .b(gate174inter2), .O(gate174inter6));
  inv1  gate280(.a(N13), .O(gate174inter7));
  inv1  gate281(.a(N695), .O(gate174inter8));
  nand2 gate282(.a(gate174inter8), .b(gate174inter7), .O(gate174inter9));
  nand2 gate283(.a(s_11), .b(gate174inter3), .O(gate174inter10));
  nor2  gate284(.a(gate174inter10), .b(gate174inter9), .O(gate174inter11));
  nor2  gate285(.a(gate174inter11), .b(gate174inter6), .O(gate174inter12));
  nand2 gate286(.a(gate174inter12), .b(gate174inter1), .O(N727));
xor2 gate175( .a(N17), .b(N696), .O(N728) );
xor2 gate176( .a(N21), .b(N697), .O(N729) );
xor2 gate177( .a(N25), .b(N698), .O(N730) );
xor2 gate178( .a(N29), .b(N699), .O(N731) );
xor2 gate179( .a(N33), .b(N700), .O(N732) );

  xor2  gate245(.a(N701), .b(N37), .O(gate180inter0));
  nand2 gate246(.a(gate180inter0), .b(s_6), .O(gate180inter1));
  and2  gate247(.a(N701), .b(N37), .O(gate180inter2));
  inv1  gate248(.a(s_6), .O(gate180inter3));
  inv1  gate249(.a(s_7), .O(gate180inter4));
  nand2 gate250(.a(gate180inter4), .b(gate180inter3), .O(gate180inter5));
  nor2  gate251(.a(gate180inter5), .b(gate180inter2), .O(gate180inter6));
  inv1  gate252(.a(N37), .O(gate180inter7));
  inv1  gate253(.a(N701), .O(gate180inter8));
  nand2 gate254(.a(gate180inter8), .b(gate180inter7), .O(gate180inter9));
  nand2 gate255(.a(s_7), .b(gate180inter3), .O(gate180inter10));
  nor2  gate256(.a(gate180inter10), .b(gate180inter9), .O(gate180inter11));
  nor2  gate257(.a(gate180inter11), .b(gate180inter6), .O(gate180inter12));
  nand2 gate258(.a(gate180inter12), .b(gate180inter1), .O(N733));

  xor2  gate203(.a(N702), .b(N41), .O(gate181inter0));
  nand2 gate204(.a(gate181inter0), .b(s_0), .O(gate181inter1));
  and2  gate205(.a(N702), .b(N41), .O(gate181inter2));
  inv1  gate206(.a(s_0), .O(gate181inter3));
  inv1  gate207(.a(s_1), .O(gate181inter4));
  nand2 gate208(.a(gate181inter4), .b(gate181inter3), .O(gate181inter5));
  nor2  gate209(.a(gate181inter5), .b(gate181inter2), .O(gate181inter6));
  inv1  gate210(.a(N41), .O(gate181inter7));
  inv1  gate211(.a(N702), .O(gate181inter8));
  nand2 gate212(.a(gate181inter8), .b(gate181inter7), .O(gate181inter9));
  nand2 gate213(.a(s_1), .b(gate181inter3), .O(gate181inter10));
  nor2  gate214(.a(gate181inter10), .b(gate181inter9), .O(gate181inter11));
  nor2  gate215(.a(gate181inter11), .b(gate181inter6), .O(gate181inter12));
  nand2 gate216(.a(gate181inter12), .b(gate181inter1), .O(N734));
xor2 gate182( .a(N45), .b(N703), .O(N735) );
xor2 gate183( .a(N49), .b(N704), .O(N736) );
xor2 gate184( .a(N53), .b(N705), .O(N737) );

  xor2  gate413(.a(N706), .b(N57), .O(gate185inter0));
  nand2 gate414(.a(gate185inter0), .b(s_30), .O(gate185inter1));
  and2  gate415(.a(N706), .b(N57), .O(gate185inter2));
  inv1  gate416(.a(s_30), .O(gate185inter3));
  inv1  gate417(.a(s_31), .O(gate185inter4));
  nand2 gate418(.a(gate185inter4), .b(gate185inter3), .O(gate185inter5));
  nor2  gate419(.a(gate185inter5), .b(gate185inter2), .O(gate185inter6));
  inv1  gate420(.a(N57), .O(gate185inter7));
  inv1  gate421(.a(N706), .O(gate185inter8));
  nand2 gate422(.a(gate185inter8), .b(gate185inter7), .O(gate185inter9));
  nand2 gate423(.a(s_31), .b(gate185inter3), .O(gate185inter10));
  nor2  gate424(.a(gate185inter10), .b(gate185inter9), .O(gate185inter11));
  nor2  gate425(.a(gate185inter11), .b(gate185inter6), .O(gate185inter12));
  nand2 gate426(.a(gate185inter12), .b(gate185inter1), .O(N738));
xor2 gate186( .a(N61), .b(N707), .O(N739) );
xor2 gate187( .a(N65), .b(N708), .O(N740) );

  xor2  gate357(.a(N709), .b(N69), .O(gate188inter0));
  nand2 gate358(.a(gate188inter0), .b(s_22), .O(gate188inter1));
  and2  gate359(.a(N709), .b(N69), .O(gate188inter2));
  inv1  gate360(.a(s_22), .O(gate188inter3));
  inv1  gate361(.a(s_23), .O(gate188inter4));
  nand2 gate362(.a(gate188inter4), .b(gate188inter3), .O(gate188inter5));
  nor2  gate363(.a(gate188inter5), .b(gate188inter2), .O(gate188inter6));
  inv1  gate364(.a(N69), .O(gate188inter7));
  inv1  gate365(.a(N709), .O(gate188inter8));
  nand2 gate366(.a(gate188inter8), .b(gate188inter7), .O(gate188inter9));
  nand2 gate367(.a(s_23), .b(gate188inter3), .O(gate188inter10));
  nor2  gate368(.a(gate188inter10), .b(gate188inter9), .O(gate188inter11));
  nor2  gate369(.a(gate188inter11), .b(gate188inter6), .O(gate188inter12));
  nand2 gate370(.a(gate188inter12), .b(gate188inter1), .O(N741));
xor2 gate189( .a(N73), .b(N710), .O(N742) );
xor2 gate190( .a(N77), .b(N711), .O(N743) );
xor2 gate191( .a(N81), .b(N712), .O(N744) );

  xor2  gate217(.a(N713), .b(N85), .O(gate192inter0));
  nand2 gate218(.a(gate192inter0), .b(s_2), .O(gate192inter1));
  and2  gate219(.a(N713), .b(N85), .O(gate192inter2));
  inv1  gate220(.a(s_2), .O(gate192inter3));
  inv1  gate221(.a(s_3), .O(gate192inter4));
  nand2 gate222(.a(gate192inter4), .b(gate192inter3), .O(gate192inter5));
  nor2  gate223(.a(gate192inter5), .b(gate192inter2), .O(gate192inter6));
  inv1  gate224(.a(N85), .O(gate192inter7));
  inv1  gate225(.a(N713), .O(gate192inter8));
  nand2 gate226(.a(gate192inter8), .b(gate192inter7), .O(gate192inter9));
  nand2 gate227(.a(s_3), .b(gate192inter3), .O(gate192inter10));
  nor2  gate228(.a(gate192inter10), .b(gate192inter9), .O(gate192inter11));
  nor2  gate229(.a(gate192inter11), .b(gate192inter6), .O(gate192inter12));
  nand2 gate230(.a(gate192inter12), .b(gate192inter1), .O(N745));
xor2 gate193( .a(N89), .b(N714), .O(N746) );
xor2 gate194( .a(N93), .b(N715), .O(N747) );
xor2 gate195( .a(N97), .b(N716), .O(N748) );
xor2 gate196( .a(N101), .b(N717), .O(N749) );
xor2 gate197( .a(N105), .b(N718), .O(N750) );
xor2 gate198( .a(N109), .b(N719), .O(N751) );
xor2 gate199( .a(N113), .b(N720), .O(N752) );
xor2 gate200( .a(N117), .b(N721), .O(N753) );
xor2 gate201( .a(N121), .b(N722), .O(N754) );
xor2 gate202( .a(N125), .b(N723), .O(N755) );

endmodule