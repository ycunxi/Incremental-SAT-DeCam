module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);

input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;//RE__PI;

input s_0,s_1;//RE__ALLOW(00,01,10,11);
input s_2,s_3;//RE__ALLOW(00,01,10,11);
input s_4,s_5;//RE__ALLOW(00,01,10,11);
input s_6,s_7;//RE__ALLOW(00,01,10,11);
input s_8,s_9;//RE__ALLOW(00,01,10,11);
input s_10,s_11;//RE__ALLOW(00,01,10,11);
input s_12,s_13;//RE__ALLOW(00,01,10,11);
input s_14,s_15;//RE__ALLOW(00,01,10,11);
input s_16,s_17;//RE__ALLOW(00,01,10,11);
input s_18,s_19;//RE__ALLOW(00,01,10,11);
input s_20,s_21;//RE__ALLOW(00,01,10,11);
input s_22,s_23;//RE__ALLOW(00,01,10,11);
input s_24,s_25;//RE__ALLOW(00,01,10,11);
input s_26,s_27;//RE__ALLOW(00,01,10,11);
input s_28,s_29;//RE__ALLOW(00,01,10,11);
input s_30,s_31;//RE__ALLOW(00,01,10,11);
input s_32,s_33;//RE__ALLOW(00,01,10,11);
input s_34,s_35;//RE__ALLOW(00,01,10,11);
input s_36,s_37;//RE__ALLOW(00,01,10,11);
input s_38,s_39;//RE__ALLOW(00,01,10,11);
input s_40,s_41;//RE__ALLOW(00,01,10,11);
input s_42,s_43;//RE__ALLOW(00,01,10,11);
input s_44,s_45;//RE__ALLOW(00,01,10,11);
input s_46,s_47;//RE__ALLOW(00,01,10,11);
input s_48,s_49;//RE__ALLOW(00,01,10,11);
input s_50,s_51;//RE__ALLOW(00,01,10,11);
input s_52,s_53;//RE__ALLOW(00,01,10,11);
input s_54,s_55;//RE__ALLOW(00,01,10,11);
input s_56,s_57;//RE__ALLOW(00,01,10,11);
input s_58,s_59;//RE__ALLOW(00,01,10,11);
input s_60,s_61;//RE__ALLOW(00,01,10,11);
input s_62,s_63;//RE__ALLOW(00,01,10,11);
input s_64,s_65;//RE__ALLOW(00,01,10,11);
input s_66,s_67;//RE__ALLOW(00,01,10,11);
input s_68,s_69;//RE__ALLOW(00,01,10,11);
input s_70,s_71;//RE__ALLOW(00,01,10,11);
input s_72,s_73;//RE__ALLOW(00,01,10,11);
input s_74,s_75;//RE__ALLOW(00,01,10,11);
input s_76,s_77;//RE__ALLOW(00,01,10,11);
input s_78,s_79;//RE__ALLOW(00,01,10,11);
input s_80,s_81;//RE__ALLOW(00,01,10,11);
input s_82,s_83;//RE__ALLOW(00,01,10,11);
input s_84,s_85;//RE__ALLOW(00,01,10,11);
input s_86,s_87;//RE__ALLOW(00,01,10,11);
input s_88,s_89;//RE__ALLOW(00,01,10,11);
input s_90,s_91;//RE__ALLOW(00,01,10,11);
input s_92,s_93;//RE__ALLOW(00,01,10,11);
input s_94,s_95;//RE__ALLOW(00,01,10,11);
input s_96,s_97;//RE__ALLOW(00,01,10,11);
input s_98,s_99;//RE__ALLOW(00,01,10,11);
input s_100,s_101;//RE__ALLOW(00,01,10,11);
input s_102,s_103;//RE__ALLOW(00,01,10,11);
input s_104,s_105;//RE__ALLOW(00,01,10,11);
input s_106,s_107;//RE__ALLOW(00,01,10,11);
input s_108,s_109;//RE__ALLOW(00,01,10,11);
input s_110,s_111;//RE__ALLOW(00,01,10,11);
input s_112,s_113;//RE__ALLOW(00,01,10,11);
input s_114,s_115;//RE__ALLOW(00,01,10,11);
input s_116,s_117;//RE__ALLOW(00,01,10,11);
input s_118,s_119;//RE__ALLOW(00,01,10,11);
input s_120,s_121;//RE__ALLOW(00,01,10,11);
input s_122,s_123;//RE__ALLOW(00,01,10,11);
input s_124,s_125;//RE__ALLOW(00,01,10,11);
input s_126,s_127;//RE__ALLOW(00,01,10,11);
input s_128,s_129;//RE__ALLOW(00,01,10,11);
input s_130,s_131;//RE__ALLOW(00,01,10,11);
input s_132,s_133;//RE__ALLOW(00,01,10,11);
input s_134,s_135;//RE__ALLOW(00,01,10,11);
input s_136,s_137;//RE__ALLOW(00,01,10,11);
input s_138,s_139;//RE__ALLOW(00,01,10,11);
input s_140,s_141;//RE__ALLOW(00,01,10,11);
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;

  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate165inter0, gate165inter1, gate165inter2, gate165inter3, gate165inter4, gate165inter5, gate165inter6, gate165inter7, gate165inter8, gate165inter9, gate165inter10, gate165inter11, gate165inter12, gate92inter0, gate92inter1, gate92inter2, gate92inter3, gate92inter4, gate92inter5, gate92inter6, gate92inter7, gate92inter8, gate92inter9, gate92inter10, gate92inter11, gate92inter12, gate455inter0, gate455inter1, gate455inter2, gate455inter3, gate455inter4, gate455inter5, gate455inter6, gate455inter7, gate455inter8, gate455inter9, gate455inter10, gate455inter11, gate455inter12, gate251inter0, gate251inter1, gate251inter2, gate251inter3, gate251inter4, gate251inter5, gate251inter6, gate251inter7, gate251inter8, gate251inter9, gate251inter10, gate251inter11, gate251inter12, gate53inter0, gate53inter1, gate53inter2, gate53inter3, gate53inter4, gate53inter5, gate53inter6, gate53inter7, gate53inter8, gate53inter9, gate53inter10, gate53inter11, gate53inter12, gate124inter0, gate124inter1, gate124inter2, gate124inter3, gate124inter4, gate124inter5, gate124inter6, gate124inter7, gate124inter8, gate124inter9, gate124inter10, gate124inter11, gate124inter12, gate248inter0, gate248inter1, gate248inter2, gate248inter3, gate248inter4, gate248inter5, gate248inter6, gate248inter7, gate248inter8, gate248inter9, gate248inter10, gate248inter11, gate248inter12, gate148inter0, gate148inter1, gate148inter2, gate148inter3, gate148inter4, gate148inter5, gate148inter6, gate148inter7, gate148inter8, gate148inter9, gate148inter10, gate148inter11, gate148inter12, gate151inter0, gate151inter1, gate151inter2, gate151inter3, gate151inter4, gate151inter5, gate151inter6, gate151inter7, gate151inter8, gate151inter9, gate151inter10, gate151inter11, gate151inter12, gate210inter0, gate210inter1, gate210inter2, gate210inter3, gate210inter4, gate210inter5, gate210inter6, gate210inter7, gate210inter8, gate210inter9, gate210inter10, gate210inter11, gate210inter12, gate97inter0, gate97inter1, gate97inter2, gate97inter3, gate97inter4, gate97inter5, gate97inter6, gate97inter7, gate97inter8, gate97inter9, gate97inter10, gate97inter11, gate97inter12, gate206inter0, gate206inter1, gate206inter2, gate206inter3, gate206inter4, gate206inter5, gate206inter6, gate206inter7, gate206inter8, gate206inter9, gate206inter10, gate206inter11, gate206inter12, gate272inter0, gate272inter1, gate272inter2, gate272inter3, gate272inter4, gate272inter5, gate272inter6, gate272inter7, gate272inter8, gate272inter9, gate272inter10, gate272inter11, gate272inter12, gate217inter0, gate217inter1, gate217inter2, gate217inter3, gate217inter4, gate217inter5, gate217inter6, gate217inter7, gate217inter8, gate217inter9, gate217inter10, gate217inter11, gate217inter12, gate243inter0, gate243inter1, gate243inter2, gate243inter3, gate243inter4, gate243inter5, gate243inter6, gate243inter7, gate243inter8, gate243inter9, gate243inter10, gate243inter11, gate243inter12, gate130inter0, gate130inter1, gate130inter2, gate130inter3, gate130inter4, gate130inter5, gate130inter6, gate130inter7, gate130inter8, gate130inter9, gate130inter10, gate130inter11, gate130inter12, gate25inter0, gate25inter1, gate25inter2, gate25inter3, gate25inter4, gate25inter5, gate25inter6, gate25inter7, gate25inter8, gate25inter9, gate25inter10, gate25inter11, gate25inter12, gate250inter0, gate250inter1, gate250inter2, gate250inter3, gate250inter4, gate250inter5, gate250inter6, gate250inter7, gate250inter8, gate250inter9, gate250inter10, gate250inter11, gate250inter12, gate21inter0, gate21inter1, gate21inter2, gate21inter3, gate21inter4, gate21inter5, gate21inter6, gate21inter7, gate21inter8, gate21inter9, gate21inter10, gate21inter11, gate21inter12, gate214inter0, gate214inter1, gate214inter2, gate214inter3, gate214inter4, gate214inter5, gate214inter6, gate214inter7, gate214inter8, gate214inter9, gate214inter10, gate214inter11, gate214inter12, gate438inter0, gate438inter1, gate438inter2, gate438inter3, gate438inter4, gate438inter5, gate438inter6, gate438inter7, gate438inter8, gate438inter9, gate438inter10, gate438inter11, gate438inter12, gate17inter0, gate17inter1, gate17inter2, gate17inter3, gate17inter4, gate17inter5, gate17inter6, gate17inter7, gate17inter8, gate17inter9, gate17inter10, gate17inter11, gate17inter12, gate93inter0, gate93inter1, gate93inter2, gate93inter3, gate93inter4, gate93inter5, gate93inter6, gate93inter7, gate93inter8, gate93inter9, gate93inter10, gate93inter11, gate93inter12, gate427inter0, gate427inter1, gate427inter2, gate427inter3, gate427inter4, gate427inter5, gate427inter6, gate427inter7, gate427inter8, gate427inter9, gate427inter10, gate427inter11, gate427inter12, gate36inter0, gate36inter1, gate36inter2, gate36inter3, gate36inter4, gate36inter5, gate36inter6, gate36inter7, gate36inter8, gate36inter9, gate36inter10, gate36inter11, gate36inter12, gate12inter0, gate12inter1, gate12inter2, gate12inter3, gate12inter4, gate12inter5, gate12inter6, gate12inter7, gate12inter8, gate12inter9, gate12inter10, gate12inter11, gate12inter12, gate187inter0, gate187inter1, gate187inter2, gate187inter3, gate187inter4, gate187inter5, gate187inter6, gate187inter7, gate187inter8, gate187inter9, gate187inter10, gate187inter11, gate187inter12, gate41inter0, gate41inter1, gate41inter2, gate41inter3, gate41inter4, gate41inter5, gate41inter6, gate41inter7, gate41inter8, gate41inter9, gate41inter10, gate41inter11, gate41inter12, gate512inter0, gate512inter1, gate512inter2, gate512inter3, gate512inter4, gate512inter5, gate512inter6, gate512inter7, gate512inter8, gate512inter9, gate512inter10, gate512inter11, gate512inter12, gate78inter0, gate78inter1, gate78inter2, gate78inter3, gate78inter4, gate78inter5, gate78inter6, gate78inter7, gate78inter8, gate78inter9, gate78inter10, gate78inter11, gate78inter12, gate452inter0, gate452inter1, gate452inter2, gate452inter3, gate452inter4, gate452inter5, gate452inter6, gate452inter7, gate452inter8, gate452inter9, gate452inter10, gate452inter11, gate452inter12, gate129inter0, gate129inter1, gate129inter2, gate129inter3, gate129inter4, gate129inter5, gate129inter6, gate129inter7, gate129inter8, gate129inter9, gate129inter10, gate129inter11, gate129inter12, gate501inter0, gate501inter1, gate501inter2, gate501inter3, gate501inter4, gate501inter5, gate501inter6, gate501inter7, gate501inter8, gate501inter9, gate501inter10, gate501inter11, gate501inter12, gate184inter0, gate184inter1, gate184inter2, gate184inter3, gate184inter4, gate184inter5, gate184inter6, gate184inter7, gate184inter8, gate184inter9, gate184inter10, gate184inter11, gate184inter12, gate446inter0, gate446inter1, gate446inter2, gate446inter3, gate446inter4, gate446inter5, gate446inter6, gate446inter7, gate446inter8, gate446inter9, gate446inter10, gate446inter11, gate446inter12, gate267inter0, gate267inter1, gate267inter2, gate267inter3, gate267inter4, gate267inter5, gate267inter6, gate267inter7, gate267inter8, gate267inter9, gate267inter10, gate267inter11, gate267inter12, gate459inter0, gate459inter1, gate459inter2, gate459inter3, gate459inter4, gate459inter5, gate459inter6, gate459inter7, gate459inter8, gate459inter9, gate459inter10, gate459inter11, gate459inter12, gate145inter0, gate145inter1, gate145inter2, gate145inter3, gate145inter4, gate145inter5, gate145inter6, gate145inter7, gate145inter8, gate145inter9, gate145inter10, gate145inter11, gate145inter12, gate141inter0, gate141inter1, gate141inter2, gate141inter3, gate141inter4, gate141inter5, gate141inter6, gate141inter7, gate141inter8, gate141inter9, gate141inter10, gate141inter11, gate141inter12, gate134inter0, gate134inter1, gate134inter2, gate134inter3, gate134inter4, gate134inter5, gate134inter6, gate134inter7, gate134inter8, gate134inter9, gate134inter10, gate134inter11, gate134inter12, gate176inter0, gate176inter1, gate176inter2, gate176inter3, gate176inter4, gate176inter5, gate176inter6, gate176inter7, gate176inter8, gate176inter9, gate176inter10, gate176inter11, gate176inter12, gate185inter0, gate185inter1, gate185inter2, gate185inter3, gate185inter4, gate185inter5, gate185inter6, gate185inter7, gate185inter8, gate185inter9, gate185inter10, gate185inter11, gate185inter12, gate125inter0, gate125inter1, gate125inter2, gate125inter3, gate125inter4, gate125inter5, gate125inter6, gate125inter7, gate125inter8, gate125inter9, gate125inter10, gate125inter11, gate125inter12, gate288inter0, gate288inter1, gate288inter2, gate288inter3, gate288inter4, gate288inter5, gate288inter6, gate288inter7, gate288inter8, gate288inter9, gate288inter10, gate288inter11, gate288inter12, gate278inter0, gate278inter1, gate278inter2, gate278inter3, gate278inter4, gate278inter5, gate278inter6, gate278inter7, gate278inter8, gate278inter9, gate278inter10, gate278inter11, gate278inter12, gate434inter0, gate434inter1, gate434inter2, gate434inter3, gate434inter4, gate434inter5, gate434inter6, gate434inter7, gate434inter8, gate434inter9, gate434inter10, gate434inter11, gate434inter12, gate491inter0, gate491inter1, gate491inter2, gate491inter3, gate491inter4, gate491inter5, gate491inter6, gate491inter7, gate491inter8, gate491inter9, gate491inter10, gate491inter11, gate491inter12, gate69inter0, gate69inter1, gate69inter2, gate69inter3, gate69inter4, gate69inter5, gate69inter6, gate69inter7, gate69inter8, gate69inter9, gate69inter10, gate69inter11, gate69inter12, gate295inter0, gate295inter1, gate295inter2, gate295inter3, gate295inter4, gate295inter5, gate295inter6, gate295inter7, gate295inter8, gate295inter9, gate295inter10, gate295inter11, gate295inter12, gate292inter0, gate292inter1, gate292inter2, gate292inter3, gate292inter4, gate292inter5, gate292inter6, gate292inter7, gate292inter8, gate292inter9, gate292inter10, gate292inter11, gate292inter12, gate126inter0, gate126inter1, gate126inter2, gate126inter3, gate126inter4, gate126inter5, gate126inter6, gate126inter7, gate126inter8, gate126inter9, gate126inter10, gate126inter11, gate126inter12, gate264inter0, gate264inter1, gate264inter2, gate264inter3, gate264inter4, gate264inter5, gate264inter6, gate264inter7, gate264inter8, gate264inter9, gate264inter10, gate264inter11, gate264inter12, gate10inter0, gate10inter1, gate10inter2, gate10inter3, gate10inter4, gate10inter5, gate10inter6, gate10inter7, gate10inter8, gate10inter9, gate10inter10, gate10inter11, gate10inter12, gate139inter0, gate139inter1, gate139inter2, gate139inter3, gate139inter4, gate139inter5, gate139inter6, gate139inter7, gate139inter8, gate139inter9, gate139inter10, gate139inter11, gate139inter12, gate508inter0, gate508inter1, gate508inter2, gate508inter3, gate508inter4, gate508inter5, gate508inter6, gate508inter7, gate508inter8, gate508inter9, gate508inter10, gate508inter11, gate508inter12, gate390inter0, gate390inter1, gate390inter2, gate390inter3, gate390inter4, gate390inter5, gate390inter6, gate390inter7, gate390inter8, gate390inter9, gate390inter10, gate390inter11, gate390inter12, gate137inter0, gate137inter1, gate137inter2, gate137inter3, gate137inter4, gate137inter5, gate137inter6, gate137inter7, gate137inter8, gate137inter9, gate137inter10, gate137inter11, gate137inter12, gate259inter0, gate259inter1, gate259inter2, gate259inter3, gate259inter4, gate259inter5, gate259inter6, gate259inter7, gate259inter8, gate259inter9, gate259inter10, gate259inter11, gate259inter12, gate44inter0, gate44inter1, gate44inter2, gate44inter3, gate44inter4, gate44inter5, gate44inter6, gate44inter7, gate44inter8, gate44inter9, gate44inter10, gate44inter11, gate44inter12, gate233inter0, gate233inter1, gate233inter2, gate233inter3, gate233inter4, gate233inter5, gate233inter6, gate233inter7, gate233inter8, gate233inter9, gate233inter10, gate233inter11, gate233inter12, gate503inter0, gate503inter1, gate503inter2, gate503inter3, gate503inter4, gate503inter5, gate503inter6, gate503inter7, gate503inter8, gate503inter9, gate503inter10, gate503inter11, gate503inter12, gate425inter0, gate425inter1, gate425inter2, gate425inter3, gate425inter4, gate425inter5, gate425inter6, gate425inter7, gate425inter8, gate425inter9, gate425inter10, gate425inter11, gate425inter12, gate26inter0, gate26inter1, gate26inter2, gate26inter3, gate26inter4, gate26inter5, gate26inter6, gate26inter7, gate26inter8, gate26inter9, gate26inter10, gate26inter11, gate26inter12, gate231inter0, gate231inter1, gate231inter2, gate231inter3, gate231inter4, gate231inter5, gate231inter6, gate231inter7, gate231inter8, gate231inter9, gate231inter10, gate231inter11, gate231inter12, gate192inter0, gate192inter1, gate192inter2, gate192inter3, gate192inter4, gate192inter5, gate192inter6, gate192inter7, gate192inter8, gate192inter9, gate192inter10, gate192inter11, gate192inter12, gate46inter0, gate46inter1, gate46inter2, gate46inter3, gate46inter4, gate46inter5, gate46inter6, gate46inter7, gate46inter8, gate46inter9, gate46inter10, gate46inter11, gate46inter12, gate204inter0, gate204inter1, gate204inter2, gate204inter3, gate204inter4, gate204inter5, gate204inter6, gate204inter7, gate204inter8, gate204inter9, gate204inter10, gate204inter11, gate204inter12, gate191inter0, gate191inter1, gate191inter2, gate191inter3, gate191inter4, gate191inter5, gate191inter6, gate191inter7, gate191inter8, gate191inter9, gate191inter10, gate191inter11, gate191inter12, gate87inter0, gate87inter1, gate87inter2, gate87inter3, gate87inter4, gate87inter5, gate87inter6, gate87inter7, gate87inter8, gate87inter9, gate87inter10, gate87inter11, gate87inter12, gate441inter0, gate441inter1, gate441inter2, gate441inter3, gate441inter4, gate441inter5, gate441inter6, gate441inter7, gate441inter8, gate441inter9, gate441inter10, gate441inter11, gate441inter12, gate22inter0, gate22inter1, gate22inter2, gate22inter3, gate22inter4, gate22inter5, gate22inter6, gate22inter7, gate22inter8, gate22inter9, gate22inter10, gate22inter11, gate22inter12;



and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );
nand2 gate9( .a(G1), .b(G2), .O(G266) );

  xor2  gate1275(.a(G4), .b(G3), .O(gate10inter0));
  nand2 gate1276(.a(gate10inter0), .b(s_104), .O(gate10inter1));
  and2  gate1277(.a(G4), .b(G3), .O(gate10inter2));
  inv1  gate1278(.a(s_104), .O(gate10inter3));
  inv1  gate1279(.a(s_105), .O(gate10inter4));
  nand2 gate1280(.a(gate10inter4), .b(gate10inter3), .O(gate10inter5));
  nor2  gate1281(.a(gate10inter5), .b(gate10inter2), .O(gate10inter6));
  inv1  gate1282(.a(G3), .O(gate10inter7));
  inv1  gate1283(.a(G4), .O(gate10inter8));
  nand2 gate1284(.a(gate10inter8), .b(gate10inter7), .O(gate10inter9));
  nand2 gate1285(.a(s_105), .b(gate10inter3), .O(gate10inter10));
  nor2  gate1286(.a(gate10inter10), .b(gate10inter9), .O(gate10inter11));
  nor2  gate1287(.a(gate10inter11), .b(gate10inter6), .O(gate10inter12));
  nand2 gate1288(.a(gate10inter12), .b(gate10inter1), .O(G269));
nand2 gate11( .a(G5), .b(G6), .O(G272) );

  xor2  gate897(.a(G8), .b(G7), .O(gate12inter0));
  nand2 gate898(.a(gate12inter0), .b(s_50), .O(gate12inter1));
  and2  gate899(.a(G8), .b(G7), .O(gate12inter2));
  inv1  gate900(.a(s_50), .O(gate12inter3));
  inv1  gate901(.a(s_51), .O(gate12inter4));
  nand2 gate902(.a(gate12inter4), .b(gate12inter3), .O(gate12inter5));
  nor2  gate903(.a(gate12inter5), .b(gate12inter2), .O(gate12inter6));
  inv1  gate904(.a(G7), .O(gate12inter7));
  inv1  gate905(.a(G8), .O(gate12inter8));
  nand2 gate906(.a(gate12inter8), .b(gate12inter7), .O(gate12inter9));
  nand2 gate907(.a(s_51), .b(gate12inter3), .O(gate12inter10));
  nor2  gate908(.a(gate12inter10), .b(gate12inter9), .O(gate12inter11));
  nor2  gate909(.a(gate12inter11), .b(gate12inter6), .O(gate12inter12));
  nand2 gate910(.a(gate12inter12), .b(gate12inter1), .O(G275));
nand2 gate13( .a(G9), .b(G10), .O(G278) );
nand2 gate14( .a(G11), .b(G12), .O(G281) );
nand2 gate15( .a(G13), .b(G14), .O(G284) );
nand2 gate16( .a(G15), .b(G16), .O(G287) );

  xor2  gate841(.a(G18), .b(G17), .O(gate17inter0));
  nand2 gate842(.a(gate17inter0), .b(s_42), .O(gate17inter1));
  and2  gate843(.a(G18), .b(G17), .O(gate17inter2));
  inv1  gate844(.a(s_42), .O(gate17inter3));
  inv1  gate845(.a(s_43), .O(gate17inter4));
  nand2 gate846(.a(gate17inter4), .b(gate17inter3), .O(gate17inter5));
  nor2  gate847(.a(gate17inter5), .b(gate17inter2), .O(gate17inter6));
  inv1  gate848(.a(G17), .O(gate17inter7));
  inv1  gate849(.a(G18), .O(gate17inter8));
  nand2 gate850(.a(gate17inter8), .b(gate17inter7), .O(gate17inter9));
  nand2 gate851(.a(s_43), .b(gate17inter3), .O(gate17inter10));
  nor2  gate852(.a(gate17inter10), .b(gate17inter9), .O(gate17inter11));
  nor2  gate853(.a(gate17inter11), .b(gate17inter6), .O(gate17inter12));
  nand2 gate854(.a(gate17inter12), .b(gate17inter1), .O(G290));
nand2 gate18( .a(G19), .b(G20), .O(G293) );
nand2 gate19( .a(G21), .b(G22), .O(G296) );
nand2 gate20( .a(G23), .b(G24), .O(G299) );

  xor2  gate799(.a(G26), .b(G25), .O(gate21inter0));
  nand2 gate800(.a(gate21inter0), .b(s_36), .O(gate21inter1));
  and2  gate801(.a(G26), .b(G25), .O(gate21inter2));
  inv1  gate802(.a(s_36), .O(gate21inter3));
  inv1  gate803(.a(s_37), .O(gate21inter4));
  nand2 gate804(.a(gate21inter4), .b(gate21inter3), .O(gate21inter5));
  nor2  gate805(.a(gate21inter5), .b(gate21inter2), .O(gate21inter6));
  inv1  gate806(.a(G25), .O(gate21inter7));
  inv1  gate807(.a(G26), .O(gate21inter8));
  nand2 gate808(.a(gate21inter8), .b(gate21inter7), .O(gate21inter9));
  nand2 gate809(.a(s_37), .b(gate21inter3), .O(gate21inter10));
  nor2  gate810(.a(gate21inter10), .b(gate21inter9), .O(gate21inter11));
  nor2  gate811(.a(gate21inter11), .b(gate21inter6), .O(gate21inter12));
  nand2 gate812(.a(gate21inter12), .b(gate21inter1), .O(G302));

  xor2  gate1527(.a(G28), .b(G27), .O(gate22inter0));
  nand2 gate1528(.a(gate22inter0), .b(s_140), .O(gate22inter1));
  and2  gate1529(.a(G28), .b(G27), .O(gate22inter2));
  inv1  gate1530(.a(s_140), .O(gate22inter3));
  inv1  gate1531(.a(s_141), .O(gate22inter4));
  nand2 gate1532(.a(gate22inter4), .b(gate22inter3), .O(gate22inter5));
  nor2  gate1533(.a(gate22inter5), .b(gate22inter2), .O(gate22inter6));
  inv1  gate1534(.a(G27), .O(gate22inter7));
  inv1  gate1535(.a(G28), .O(gate22inter8));
  nand2 gate1536(.a(gate22inter8), .b(gate22inter7), .O(gate22inter9));
  nand2 gate1537(.a(s_141), .b(gate22inter3), .O(gate22inter10));
  nor2  gate1538(.a(gate22inter10), .b(gate22inter9), .O(gate22inter11));
  nor2  gate1539(.a(gate22inter11), .b(gate22inter6), .O(gate22inter12));
  nand2 gate1540(.a(gate22inter12), .b(gate22inter1), .O(G305));
nand2 gate23( .a(G29), .b(G30), .O(G308) );
nand2 gate24( .a(G31), .b(G32), .O(G311) );

  xor2  gate771(.a(G5), .b(G1), .O(gate25inter0));
  nand2 gate772(.a(gate25inter0), .b(s_32), .O(gate25inter1));
  and2  gate773(.a(G5), .b(G1), .O(gate25inter2));
  inv1  gate774(.a(s_32), .O(gate25inter3));
  inv1  gate775(.a(s_33), .O(gate25inter4));
  nand2 gate776(.a(gate25inter4), .b(gate25inter3), .O(gate25inter5));
  nor2  gate777(.a(gate25inter5), .b(gate25inter2), .O(gate25inter6));
  inv1  gate778(.a(G1), .O(gate25inter7));
  inv1  gate779(.a(G5), .O(gate25inter8));
  nand2 gate780(.a(gate25inter8), .b(gate25inter7), .O(gate25inter9));
  nand2 gate781(.a(s_33), .b(gate25inter3), .O(gate25inter10));
  nor2  gate782(.a(gate25inter10), .b(gate25inter9), .O(gate25inter11));
  nor2  gate783(.a(gate25inter11), .b(gate25inter6), .O(gate25inter12));
  nand2 gate784(.a(gate25inter12), .b(gate25inter1), .O(G314));

  xor2  gate1415(.a(G13), .b(G9), .O(gate26inter0));
  nand2 gate1416(.a(gate26inter0), .b(s_124), .O(gate26inter1));
  and2  gate1417(.a(G13), .b(G9), .O(gate26inter2));
  inv1  gate1418(.a(s_124), .O(gate26inter3));
  inv1  gate1419(.a(s_125), .O(gate26inter4));
  nand2 gate1420(.a(gate26inter4), .b(gate26inter3), .O(gate26inter5));
  nor2  gate1421(.a(gate26inter5), .b(gate26inter2), .O(gate26inter6));
  inv1  gate1422(.a(G9), .O(gate26inter7));
  inv1  gate1423(.a(G13), .O(gate26inter8));
  nand2 gate1424(.a(gate26inter8), .b(gate26inter7), .O(gate26inter9));
  nand2 gate1425(.a(s_125), .b(gate26inter3), .O(gate26inter10));
  nor2  gate1426(.a(gate26inter10), .b(gate26inter9), .O(gate26inter11));
  nor2  gate1427(.a(gate26inter11), .b(gate26inter6), .O(gate26inter12));
  nand2 gate1428(.a(gate26inter12), .b(gate26inter1), .O(G317));
nand2 gate27( .a(G2), .b(G6), .O(G320) );
nand2 gate28( .a(G10), .b(G14), .O(G323) );
nand2 gate29( .a(G3), .b(G7), .O(G326) );
nand2 gate30( .a(G11), .b(G15), .O(G329) );
nand2 gate31( .a(G4), .b(G8), .O(G332) );
nand2 gate32( .a(G12), .b(G16), .O(G335) );
nand2 gate33( .a(G17), .b(G21), .O(G338) );
nand2 gate34( .a(G25), .b(G29), .O(G341) );
nand2 gate35( .a(G18), .b(G22), .O(G344) );

  xor2  gate883(.a(G30), .b(G26), .O(gate36inter0));
  nand2 gate884(.a(gate36inter0), .b(s_48), .O(gate36inter1));
  and2  gate885(.a(G30), .b(G26), .O(gate36inter2));
  inv1  gate886(.a(s_48), .O(gate36inter3));
  inv1  gate887(.a(s_49), .O(gate36inter4));
  nand2 gate888(.a(gate36inter4), .b(gate36inter3), .O(gate36inter5));
  nor2  gate889(.a(gate36inter5), .b(gate36inter2), .O(gate36inter6));
  inv1  gate890(.a(G26), .O(gate36inter7));
  inv1  gate891(.a(G30), .O(gate36inter8));
  nand2 gate892(.a(gate36inter8), .b(gate36inter7), .O(gate36inter9));
  nand2 gate893(.a(s_49), .b(gate36inter3), .O(gate36inter10));
  nor2  gate894(.a(gate36inter10), .b(gate36inter9), .O(gate36inter11));
  nor2  gate895(.a(gate36inter11), .b(gate36inter6), .O(gate36inter12));
  nand2 gate896(.a(gate36inter12), .b(gate36inter1), .O(G347));
nand2 gate37( .a(G19), .b(G23), .O(G350) );
nand2 gate38( .a(G27), .b(G31), .O(G353) );
nand2 gate39( .a(G20), .b(G24), .O(G356) );
nand2 gate40( .a(G28), .b(G32), .O(G359) );

  xor2  gate925(.a(G266), .b(G1), .O(gate41inter0));
  nand2 gate926(.a(gate41inter0), .b(s_54), .O(gate41inter1));
  and2  gate927(.a(G266), .b(G1), .O(gate41inter2));
  inv1  gate928(.a(s_54), .O(gate41inter3));
  inv1  gate929(.a(s_55), .O(gate41inter4));
  nand2 gate930(.a(gate41inter4), .b(gate41inter3), .O(gate41inter5));
  nor2  gate931(.a(gate41inter5), .b(gate41inter2), .O(gate41inter6));
  inv1  gate932(.a(G1), .O(gate41inter7));
  inv1  gate933(.a(G266), .O(gate41inter8));
  nand2 gate934(.a(gate41inter8), .b(gate41inter7), .O(gate41inter9));
  nand2 gate935(.a(s_55), .b(gate41inter3), .O(gate41inter10));
  nor2  gate936(.a(gate41inter10), .b(gate41inter9), .O(gate41inter11));
  nor2  gate937(.a(gate41inter11), .b(gate41inter6), .O(gate41inter12));
  nand2 gate938(.a(gate41inter12), .b(gate41inter1), .O(G362));
nand2 gate42( .a(G2), .b(G266), .O(G363) );
nand2 gate43( .a(G3), .b(G269), .O(G364) );

  xor2  gate1359(.a(G269), .b(G4), .O(gate44inter0));
  nand2 gate1360(.a(gate44inter0), .b(s_116), .O(gate44inter1));
  and2  gate1361(.a(G269), .b(G4), .O(gate44inter2));
  inv1  gate1362(.a(s_116), .O(gate44inter3));
  inv1  gate1363(.a(s_117), .O(gate44inter4));
  nand2 gate1364(.a(gate44inter4), .b(gate44inter3), .O(gate44inter5));
  nor2  gate1365(.a(gate44inter5), .b(gate44inter2), .O(gate44inter6));
  inv1  gate1366(.a(G4), .O(gate44inter7));
  inv1  gate1367(.a(G269), .O(gate44inter8));
  nand2 gate1368(.a(gate44inter8), .b(gate44inter7), .O(gate44inter9));
  nand2 gate1369(.a(s_117), .b(gate44inter3), .O(gate44inter10));
  nor2  gate1370(.a(gate44inter10), .b(gate44inter9), .O(gate44inter11));
  nor2  gate1371(.a(gate44inter11), .b(gate44inter6), .O(gate44inter12));
  nand2 gate1372(.a(gate44inter12), .b(gate44inter1), .O(G365));
nand2 gate45( .a(G5), .b(G272), .O(G366) );

  xor2  gate1457(.a(G272), .b(G6), .O(gate46inter0));
  nand2 gate1458(.a(gate46inter0), .b(s_130), .O(gate46inter1));
  and2  gate1459(.a(G272), .b(G6), .O(gate46inter2));
  inv1  gate1460(.a(s_130), .O(gate46inter3));
  inv1  gate1461(.a(s_131), .O(gate46inter4));
  nand2 gate1462(.a(gate46inter4), .b(gate46inter3), .O(gate46inter5));
  nor2  gate1463(.a(gate46inter5), .b(gate46inter2), .O(gate46inter6));
  inv1  gate1464(.a(G6), .O(gate46inter7));
  inv1  gate1465(.a(G272), .O(gate46inter8));
  nand2 gate1466(.a(gate46inter8), .b(gate46inter7), .O(gate46inter9));
  nand2 gate1467(.a(s_131), .b(gate46inter3), .O(gate46inter10));
  nor2  gate1468(.a(gate46inter10), .b(gate46inter9), .O(gate46inter11));
  nor2  gate1469(.a(gate46inter11), .b(gate46inter6), .O(gate46inter12));
  nand2 gate1470(.a(gate46inter12), .b(gate46inter1), .O(G367));
nand2 gate47( .a(G7), .b(G275), .O(G368) );
nand2 gate48( .a(G8), .b(G275), .O(G369) );
nand2 gate49( .a(G9), .b(G278), .O(G370) );
nand2 gate50( .a(G10), .b(G278), .O(G371) );
nand2 gate51( .a(G11), .b(G281), .O(G372) );
nand2 gate52( .a(G12), .b(G281), .O(G373) );

  xor2  gate603(.a(G284), .b(G13), .O(gate53inter0));
  nand2 gate604(.a(gate53inter0), .b(s_8), .O(gate53inter1));
  and2  gate605(.a(G284), .b(G13), .O(gate53inter2));
  inv1  gate606(.a(s_8), .O(gate53inter3));
  inv1  gate607(.a(s_9), .O(gate53inter4));
  nand2 gate608(.a(gate53inter4), .b(gate53inter3), .O(gate53inter5));
  nor2  gate609(.a(gate53inter5), .b(gate53inter2), .O(gate53inter6));
  inv1  gate610(.a(G13), .O(gate53inter7));
  inv1  gate611(.a(G284), .O(gate53inter8));
  nand2 gate612(.a(gate53inter8), .b(gate53inter7), .O(gate53inter9));
  nand2 gate613(.a(s_9), .b(gate53inter3), .O(gate53inter10));
  nor2  gate614(.a(gate53inter10), .b(gate53inter9), .O(gate53inter11));
  nor2  gate615(.a(gate53inter11), .b(gate53inter6), .O(gate53inter12));
  nand2 gate616(.a(gate53inter12), .b(gate53inter1), .O(G374));
nand2 gate54( .a(G14), .b(G284), .O(G375) );
nand2 gate55( .a(G15), .b(G287), .O(G376) );
nand2 gate56( .a(G16), .b(G287), .O(G377) );
nand2 gate57( .a(G17), .b(G290), .O(G378) );
nand2 gate58( .a(G18), .b(G290), .O(G379) );
nand2 gate59( .a(G19), .b(G293), .O(G380) );
nand2 gate60( .a(G20), .b(G293), .O(G381) );
nand2 gate61( .a(G21), .b(G296), .O(G382) );
nand2 gate62( .a(G22), .b(G296), .O(G383) );
nand2 gate63( .a(G23), .b(G299), .O(G384) );
nand2 gate64( .a(G24), .b(G299), .O(G385) );
nand2 gate65( .a(G25), .b(G302), .O(G386) );
nand2 gate66( .a(G26), .b(G302), .O(G387) );
nand2 gate67( .a(G27), .b(G305), .O(G388) );
nand2 gate68( .a(G28), .b(G305), .O(G389) );

  xor2  gate1205(.a(G308), .b(G29), .O(gate69inter0));
  nand2 gate1206(.a(gate69inter0), .b(s_94), .O(gate69inter1));
  and2  gate1207(.a(G308), .b(G29), .O(gate69inter2));
  inv1  gate1208(.a(s_94), .O(gate69inter3));
  inv1  gate1209(.a(s_95), .O(gate69inter4));
  nand2 gate1210(.a(gate69inter4), .b(gate69inter3), .O(gate69inter5));
  nor2  gate1211(.a(gate69inter5), .b(gate69inter2), .O(gate69inter6));
  inv1  gate1212(.a(G29), .O(gate69inter7));
  inv1  gate1213(.a(G308), .O(gate69inter8));
  nand2 gate1214(.a(gate69inter8), .b(gate69inter7), .O(gate69inter9));
  nand2 gate1215(.a(s_95), .b(gate69inter3), .O(gate69inter10));
  nor2  gate1216(.a(gate69inter10), .b(gate69inter9), .O(gate69inter11));
  nor2  gate1217(.a(gate69inter11), .b(gate69inter6), .O(gate69inter12));
  nand2 gate1218(.a(gate69inter12), .b(gate69inter1), .O(G390));
nand2 gate70( .a(G30), .b(G308), .O(G391) );
nand2 gate71( .a(G31), .b(G311), .O(G392) );
nand2 gate72( .a(G32), .b(G311), .O(G393) );
nand2 gate73( .a(G1), .b(G314), .O(G394) );
nand2 gate74( .a(G5), .b(G314), .O(G395) );
nand2 gate75( .a(G9), .b(G317), .O(G396) );
nand2 gate76( .a(G13), .b(G317), .O(G397) );
nand2 gate77( .a(G2), .b(G320), .O(G398) );

  xor2  gate953(.a(G320), .b(G6), .O(gate78inter0));
  nand2 gate954(.a(gate78inter0), .b(s_58), .O(gate78inter1));
  and2  gate955(.a(G320), .b(G6), .O(gate78inter2));
  inv1  gate956(.a(s_58), .O(gate78inter3));
  inv1  gate957(.a(s_59), .O(gate78inter4));
  nand2 gate958(.a(gate78inter4), .b(gate78inter3), .O(gate78inter5));
  nor2  gate959(.a(gate78inter5), .b(gate78inter2), .O(gate78inter6));
  inv1  gate960(.a(G6), .O(gate78inter7));
  inv1  gate961(.a(G320), .O(gate78inter8));
  nand2 gate962(.a(gate78inter8), .b(gate78inter7), .O(gate78inter9));
  nand2 gate963(.a(s_59), .b(gate78inter3), .O(gate78inter10));
  nor2  gate964(.a(gate78inter10), .b(gate78inter9), .O(gate78inter11));
  nor2  gate965(.a(gate78inter11), .b(gate78inter6), .O(gate78inter12));
  nand2 gate966(.a(gate78inter12), .b(gate78inter1), .O(G399));
nand2 gate79( .a(G10), .b(G323), .O(G400) );
nand2 gate80( .a(G14), .b(G323), .O(G401) );
nand2 gate81( .a(G3), .b(G326), .O(G402) );
nand2 gate82( .a(G7), .b(G326), .O(G403) );
nand2 gate83( .a(G11), .b(G329), .O(G404) );
nand2 gate84( .a(G15), .b(G329), .O(G405) );
nand2 gate85( .a(G4), .b(G332), .O(G406) );
nand2 gate86( .a(G8), .b(G332), .O(G407) );

  xor2  gate1499(.a(G335), .b(G12), .O(gate87inter0));
  nand2 gate1500(.a(gate87inter0), .b(s_136), .O(gate87inter1));
  and2  gate1501(.a(G335), .b(G12), .O(gate87inter2));
  inv1  gate1502(.a(s_136), .O(gate87inter3));
  inv1  gate1503(.a(s_137), .O(gate87inter4));
  nand2 gate1504(.a(gate87inter4), .b(gate87inter3), .O(gate87inter5));
  nor2  gate1505(.a(gate87inter5), .b(gate87inter2), .O(gate87inter6));
  inv1  gate1506(.a(G12), .O(gate87inter7));
  inv1  gate1507(.a(G335), .O(gate87inter8));
  nand2 gate1508(.a(gate87inter8), .b(gate87inter7), .O(gate87inter9));
  nand2 gate1509(.a(s_137), .b(gate87inter3), .O(gate87inter10));
  nor2  gate1510(.a(gate87inter10), .b(gate87inter9), .O(gate87inter11));
  nor2  gate1511(.a(gate87inter11), .b(gate87inter6), .O(gate87inter12));
  nand2 gate1512(.a(gate87inter12), .b(gate87inter1), .O(G408));
nand2 gate88( .a(G16), .b(G335), .O(G409) );
nand2 gate89( .a(G17), .b(G338), .O(G410) );
nand2 gate90( .a(G21), .b(G338), .O(G411) );
nand2 gate91( .a(G25), .b(G341), .O(G412) );

  xor2  gate561(.a(G341), .b(G29), .O(gate92inter0));
  nand2 gate562(.a(gate92inter0), .b(s_2), .O(gate92inter1));
  and2  gate563(.a(G341), .b(G29), .O(gate92inter2));
  inv1  gate564(.a(s_2), .O(gate92inter3));
  inv1  gate565(.a(s_3), .O(gate92inter4));
  nand2 gate566(.a(gate92inter4), .b(gate92inter3), .O(gate92inter5));
  nor2  gate567(.a(gate92inter5), .b(gate92inter2), .O(gate92inter6));
  inv1  gate568(.a(G29), .O(gate92inter7));
  inv1  gate569(.a(G341), .O(gate92inter8));
  nand2 gate570(.a(gate92inter8), .b(gate92inter7), .O(gate92inter9));
  nand2 gate571(.a(s_3), .b(gate92inter3), .O(gate92inter10));
  nor2  gate572(.a(gate92inter10), .b(gate92inter9), .O(gate92inter11));
  nor2  gate573(.a(gate92inter11), .b(gate92inter6), .O(gate92inter12));
  nand2 gate574(.a(gate92inter12), .b(gate92inter1), .O(G413));

  xor2  gate855(.a(G344), .b(G18), .O(gate93inter0));
  nand2 gate856(.a(gate93inter0), .b(s_44), .O(gate93inter1));
  and2  gate857(.a(G344), .b(G18), .O(gate93inter2));
  inv1  gate858(.a(s_44), .O(gate93inter3));
  inv1  gate859(.a(s_45), .O(gate93inter4));
  nand2 gate860(.a(gate93inter4), .b(gate93inter3), .O(gate93inter5));
  nor2  gate861(.a(gate93inter5), .b(gate93inter2), .O(gate93inter6));
  inv1  gate862(.a(G18), .O(gate93inter7));
  inv1  gate863(.a(G344), .O(gate93inter8));
  nand2 gate864(.a(gate93inter8), .b(gate93inter7), .O(gate93inter9));
  nand2 gate865(.a(s_45), .b(gate93inter3), .O(gate93inter10));
  nor2  gate866(.a(gate93inter10), .b(gate93inter9), .O(gate93inter11));
  nor2  gate867(.a(gate93inter11), .b(gate93inter6), .O(gate93inter12));
  nand2 gate868(.a(gate93inter12), .b(gate93inter1), .O(G414));
nand2 gate94( .a(G22), .b(G344), .O(G415) );
nand2 gate95( .a(G26), .b(G347), .O(G416) );
nand2 gate96( .a(G30), .b(G347), .O(G417) );

  xor2  gate687(.a(G350), .b(G19), .O(gate97inter0));
  nand2 gate688(.a(gate97inter0), .b(s_20), .O(gate97inter1));
  and2  gate689(.a(G350), .b(G19), .O(gate97inter2));
  inv1  gate690(.a(s_20), .O(gate97inter3));
  inv1  gate691(.a(s_21), .O(gate97inter4));
  nand2 gate692(.a(gate97inter4), .b(gate97inter3), .O(gate97inter5));
  nor2  gate693(.a(gate97inter5), .b(gate97inter2), .O(gate97inter6));
  inv1  gate694(.a(G19), .O(gate97inter7));
  inv1  gate695(.a(G350), .O(gate97inter8));
  nand2 gate696(.a(gate97inter8), .b(gate97inter7), .O(gate97inter9));
  nand2 gate697(.a(s_21), .b(gate97inter3), .O(gate97inter10));
  nor2  gate698(.a(gate97inter10), .b(gate97inter9), .O(gate97inter11));
  nor2  gate699(.a(gate97inter11), .b(gate97inter6), .O(gate97inter12));
  nand2 gate700(.a(gate97inter12), .b(gate97inter1), .O(G418));
nand2 gate98( .a(G23), .b(G350), .O(G419) );
nand2 gate99( .a(G27), .b(G353), .O(G420) );
nand2 gate100( .a(G31), .b(G353), .O(G421) );
nand2 gate101( .a(G20), .b(G356), .O(G422) );
nand2 gate102( .a(G24), .b(G356), .O(G423) );
nand2 gate103( .a(G28), .b(G359), .O(G424) );
nand2 gate104( .a(G32), .b(G359), .O(G425) );
nand2 gate105( .a(G362), .b(G363), .O(G426) );
nand2 gate106( .a(G364), .b(G365), .O(G429) );
nand2 gate107( .a(G366), .b(G367), .O(G432) );
nand2 gate108( .a(G368), .b(G369), .O(G435) );
nand2 gate109( .a(G370), .b(G371), .O(G438) );
nand2 gate110( .a(G372), .b(G373), .O(G441) );
nand2 gate111( .a(G374), .b(G375), .O(G444) );
nand2 gate112( .a(G376), .b(G377), .O(G447) );
nand2 gate113( .a(G378), .b(G379), .O(G450) );
nand2 gate114( .a(G380), .b(G381), .O(G453) );
nand2 gate115( .a(G382), .b(G383), .O(G456) );
nand2 gate116( .a(G384), .b(G385), .O(G459) );
nand2 gate117( .a(G386), .b(G387), .O(G462) );
nand2 gate118( .a(G388), .b(G389), .O(G465) );
nand2 gate119( .a(G390), .b(G391), .O(G468) );
nand2 gate120( .a(G392), .b(G393), .O(G471) );
nand2 gate121( .a(G394), .b(G395), .O(G474) );
nand2 gate122( .a(G396), .b(G397), .O(G477) );
nand2 gate123( .a(G398), .b(G399), .O(G480) );

  xor2  gate617(.a(G401), .b(G400), .O(gate124inter0));
  nand2 gate618(.a(gate124inter0), .b(s_10), .O(gate124inter1));
  and2  gate619(.a(G401), .b(G400), .O(gate124inter2));
  inv1  gate620(.a(s_10), .O(gate124inter3));
  inv1  gate621(.a(s_11), .O(gate124inter4));
  nand2 gate622(.a(gate124inter4), .b(gate124inter3), .O(gate124inter5));
  nor2  gate623(.a(gate124inter5), .b(gate124inter2), .O(gate124inter6));
  inv1  gate624(.a(G400), .O(gate124inter7));
  inv1  gate625(.a(G401), .O(gate124inter8));
  nand2 gate626(.a(gate124inter8), .b(gate124inter7), .O(gate124inter9));
  nand2 gate627(.a(s_11), .b(gate124inter3), .O(gate124inter10));
  nor2  gate628(.a(gate124inter10), .b(gate124inter9), .O(gate124inter11));
  nor2  gate629(.a(gate124inter11), .b(gate124inter6), .O(gate124inter12));
  nand2 gate630(.a(gate124inter12), .b(gate124inter1), .O(G483));

  xor2  gate1135(.a(G403), .b(G402), .O(gate125inter0));
  nand2 gate1136(.a(gate125inter0), .b(s_84), .O(gate125inter1));
  and2  gate1137(.a(G403), .b(G402), .O(gate125inter2));
  inv1  gate1138(.a(s_84), .O(gate125inter3));
  inv1  gate1139(.a(s_85), .O(gate125inter4));
  nand2 gate1140(.a(gate125inter4), .b(gate125inter3), .O(gate125inter5));
  nor2  gate1141(.a(gate125inter5), .b(gate125inter2), .O(gate125inter6));
  inv1  gate1142(.a(G402), .O(gate125inter7));
  inv1  gate1143(.a(G403), .O(gate125inter8));
  nand2 gate1144(.a(gate125inter8), .b(gate125inter7), .O(gate125inter9));
  nand2 gate1145(.a(s_85), .b(gate125inter3), .O(gate125inter10));
  nor2  gate1146(.a(gate125inter10), .b(gate125inter9), .O(gate125inter11));
  nor2  gate1147(.a(gate125inter11), .b(gate125inter6), .O(gate125inter12));
  nand2 gate1148(.a(gate125inter12), .b(gate125inter1), .O(G486));

  xor2  gate1247(.a(G405), .b(G404), .O(gate126inter0));
  nand2 gate1248(.a(gate126inter0), .b(s_100), .O(gate126inter1));
  and2  gate1249(.a(G405), .b(G404), .O(gate126inter2));
  inv1  gate1250(.a(s_100), .O(gate126inter3));
  inv1  gate1251(.a(s_101), .O(gate126inter4));
  nand2 gate1252(.a(gate126inter4), .b(gate126inter3), .O(gate126inter5));
  nor2  gate1253(.a(gate126inter5), .b(gate126inter2), .O(gate126inter6));
  inv1  gate1254(.a(G404), .O(gate126inter7));
  inv1  gate1255(.a(G405), .O(gate126inter8));
  nand2 gate1256(.a(gate126inter8), .b(gate126inter7), .O(gate126inter9));
  nand2 gate1257(.a(s_101), .b(gate126inter3), .O(gate126inter10));
  nor2  gate1258(.a(gate126inter10), .b(gate126inter9), .O(gate126inter11));
  nor2  gate1259(.a(gate126inter11), .b(gate126inter6), .O(gate126inter12));
  nand2 gate1260(.a(gate126inter12), .b(gate126inter1), .O(G489));
nand2 gate127( .a(G406), .b(G407), .O(G492) );
nand2 gate128( .a(G408), .b(G409), .O(G495) );

  xor2  gate981(.a(G411), .b(G410), .O(gate129inter0));
  nand2 gate982(.a(gate129inter0), .b(s_62), .O(gate129inter1));
  and2  gate983(.a(G411), .b(G410), .O(gate129inter2));
  inv1  gate984(.a(s_62), .O(gate129inter3));
  inv1  gate985(.a(s_63), .O(gate129inter4));
  nand2 gate986(.a(gate129inter4), .b(gate129inter3), .O(gate129inter5));
  nor2  gate987(.a(gate129inter5), .b(gate129inter2), .O(gate129inter6));
  inv1  gate988(.a(G410), .O(gate129inter7));
  inv1  gate989(.a(G411), .O(gate129inter8));
  nand2 gate990(.a(gate129inter8), .b(gate129inter7), .O(gate129inter9));
  nand2 gate991(.a(s_63), .b(gate129inter3), .O(gate129inter10));
  nor2  gate992(.a(gate129inter10), .b(gate129inter9), .O(gate129inter11));
  nor2  gate993(.a(gate129inter11), .b(gate129inter6), .O(gate129inter12));
  nand2 gate994(.a(gate129inter12), .b(gate129inter1), .O(G498));

  xor2  gate757(.a(G413), .b(G412), .O(gate130inter0));
  nand2 gate758(.a(gate130inter0), .b(s_30), .O(gate130inter1));
  and2  gate759(.a(G413), .b(G412), .O(gate130inter2));
  inv1  gate760(.a(s_30), .O(gate130inter3));
  inv1  gate761(.a(s_31), .O(gate130inter4));
  nand2 gate762(.a(gate130inter4), .b(gate130inter3), .O(gate130inter5));
  nor2  gate763(.a(gate130inter5), .b(gate130inter2), .O(gate130inter6));
  inv1  gate764(.a(G412), .O(gate130inter7));
  inv1  gate765(.a(G413), .O(gate130inter8));
  nand2 gate766(.a(gate130inter8), .b(gate130inter7), .O(gate130inter9));
  nand2 gate767(.a(s_31), .b(gate130inter3), .O(gate130inter10));
  nor2  gate768(.a(gate130inter10), .b(gate130inter9), .O(gate130inter11));
  nor2  gate769(.a(gate130inter11), .b(gate130inter6), .O(gate130inter12));
  nand2 gate770(.a(gate130inter12), .b(gate130inter1), .O(G501));
nand2 gate131( .a(G414), .b(G415), .O(G504) );
nand2 gate132( .a(G416), .b(G417), .O(G507) );
nand2 gate133( .a(G418), .b(G419), .O(G510) );

  xor2  gate1093(.a(G421), .b(G420), .O(gate134inter0));
  nand2 gate1094(.a(gate134inter0), .b(s_78), .O(gate134inter1));
  and2  gate1095(.a(G421), .b(G420), .O(gate134inter2));
  inv1  gate1096(.a(s_78), .O(gate134inter3));
  inv1  gate1097(.a(s_79), .O(gate134inter4));
  nand2 gate1098(.a(gate134inter4), .b(gate134inter3), .O(gate134inter5));
  nor2  gate1099(.a(gate134inter5), .b(gate134inter2), .O(gate134inter6));
  inv1  gate1100(.a(G420), .O(gate134inter7));
  inv1  gate1101(.a(G421), .O(gate134inter8));
  nand2 gate1102(.a(gate134inter8), .b(gate134inter7), .O(gate134inter9));
  nand2 gate1103(.a(s_79), .b(gate134inter3), .O(gate134inter10));
  nor2  gate1104(.a(gate134inter10), .b(gate134inter9), .O(gate134inter11));
  nor2  gate1105(.a(gate134inter11), .b(gate134inter6), .O(gate134inter12));
  nand2 gate1106(.a(gate134inter12), .b(gate134inter1), .O(G513));
nand2 gate135( .a(G422), .b(G423), .O(G516) );
nand2 gate136( .a(G424), .b(G425), .O(G519) );

  xor2  gate1331(.a(G429), .b(G426), .O(gate137inter0));
  nand2 gate1332(.a(gate137inter0), .b(s_112), .O(gate137inter1));
  and2  gate1333(.a(G429), .b(G426), .O(gate137inter2));
  inv1  gate1334(.a(s_112), .O(gate137inter3));
  inv1  gate1335(.a(s_113), .O(gate137inter4));
  nand2 gate1336(.a(gate137inter4), .b(gate137inter3), .O(gate137inter5));
  nor2  gate1337(.a(gate137inter5), .b(gate137inter2), .O(gate137inter6));
  inv1  gate1338(.a(G426), .O(gate137inter7));
  inv1  gate1339(.a(G429), .O(gate137inter8));
  nand2 gate1340(.a(gate137inter8), .b(gate137inter7), .O(gate137inter9));
  nand2 gate1341(.a(s_113), .b(gate137inter3), .O(gate137inter10));
  nor2  gate1342(.a(gate137inter10), .b(gate137inter9), .O(gate137inter11));
  nor2  gate1343(.a(gate137inter11), .b(gate137inter6), .O(gate137inter12));
  nand2 gate1344(.a(gate137inter12), .b(gate137inter1), .O(G522));
nand2 gate138( .a(G432), .b(G435), .O(G525) );

  xor2  gate1289(.a(G441), .b(G438), .O(gate139inter0));
  nand2 gate1290(.a(gate139inter0), .b(s_106), .O(gate139inter1));
  and2  gate1291(.a(G441), .b(G438), .O(gate139inter2));
  inv1  gate1292(.a(s_106), .O(gate139inter3));
  inv1  gate1293(.a(s_107), .O(gate139inter4));
  nand2 gate1294(.a(gate139inter4), .b(gate139inter3), .O(gate139inter5));
  nor2  gate1295(.a(gate139inter5), .b(gate139inter2), .O(gate139inter6));
  inv1  gate1296(.a(G438), .O(gate139inter7));
  inv1  gate1297(.a(G441), .O(gate139inter8));
  nand2 gate1298(.a(gate139inter8), .b(gate139inter7), .O(gate139inter9));
  nand2 gate1299(.a(s_107), .b(gate139inter3), .O(gate139inter10));
  nor2  gate1300(.a(gate139inter10), .b(gate139inter9), .O(gate139inter11));
  nor2  gate1301(.a(gate139inter11), .b(gate139inter6), .O(gate139inter12));
  nand2 gate1302(.a(gate139inter12), .b(gate139inter1), .O(G528));
nand2 gate140( .a(G444), .b(G447), .O(G531) );

  xor2  gate1079(.a(G453), .b(G450), .O(gate141inter0));
  nand2 gate1080(.a(gate141inter0), .b(s_76), .O(gate141inter1));
  and2  gate1081(.a(G453), .b(G450), .O(gate141inter2));
  inv1  gate1082(.a(s_76), .O(gate141inter3));
  inv1  gate1083(.a(s_77), .O(gate141inter4));
  nand2 gate1084(.a(gate141inter4), .b(gate141inter3), .O(gate141inter5));
  nor2  gate1085(.a(gate141inter5), .b(gate141inter2), .O(gate141inter6));
  inv1  gate1086(.a(G450), .O(gate141inter7));
  inv1  gate1087(.a(G453), .O(gate141inter8));
  nand2 gate1088(.a(gate141inter8), .b(gate141inter7), .O(gate141inter9));
  nand2 gate1089(.a(s_77), .b(gate141inter3), .O(gate141inter10));
  nor2  gate1090(.a(gate141inter10), .b(gate141inter9), .O(gate141inter11));
  nor2  gate1091(.a(gate141inter11), .b(gate141inter6), .O(gate141inter12));
  nand2 gate1092(.a(gate141inter12), .b(gate141inter1), .O(G534));
nand2 gate142( .a(G456), .b(G459), .O(G537) );
nand2 gate143( .a(G462), .b(G465), .O(G540) );
nand2 gate144( .a(G468), .b(G471), .O(G543) );

  xor2  gate1065(.a(G477), .b(G474), .O(gate145inter0));
  nand2 gate1066(.a(gate145inter0), .b(s_74), .O(gate145inter1));
  and2  gate1067(.a(G477), .b(G474), .O(gate145inter2));
  inv1  gate1068(.a(s_74), .O(gate145inter3));
  inv1  gate1069(.a(s_75), .O(gate145inter4));
  nand2 gate1070(.a(gate145inter4), .b(gate145inter3), .O(gate145inter5));
  nor2  gate1071(.a(gate145inter5), .b(gate145inter2), .O(gate145inter6));
  inv1  gate1072(.a(G474), .O(gate145inter7));
  inv1  gate1073(.a(G477), .O(gate145inter8));
  nand2 gate1074(.a(gate145inter8), .b(gate145inter7), .O(gate145inter9));
  nand2 gate1075(.a(s_75), .b(gate145inter3), .O(gate145inter10));
  nor2  gate1076(.a(gate145inter10), .b(gate145inter9), .O(gate145inter11));
  nor2  gate1077(.a(gate145inter11), .b(gate145inter6), .O(gate145inter12));
  nand2 gate1078(.a(gate145inter12), .b(gate145inter1), .O(G546));
nand2 gate146( .a(G480), .b(G483), .O(G549) );
nand2 gate147( .a(G486), .b(G489), .O(G552) );

  xor2  gate645(.a(G495), .b(G492), .O(gate148inter0));
  nand2 gate646(.a(gate148inter0), .b(s_14), .O(gate148inter1));
  and2  gate647(.a(G495), .b(G492), .O(gate148inter2));
  inv1  gate648(.a(s_14), .O(gate148inter3));
  inv1  gate649(.a(s_15), .O(gate148inter4));
  nand2 gate650(.a(gate148inter4), .b(gate148inter3), .O(gate148inter5));
  nor2  gate651(.a(gate148inter5), .b(gate148inter2), .O(gate148inter6));
  inv1  gate652(.a(G492), .O(gate148inter7));
  inv1  gate653(.a(G495), .O(gate148inter8));
  nand2 gate654(.a(gate148inter8), .b(gate148inter7), .O(gate148inter9));
  nand2 gate655(.a(s_15), .b(gate148inter3), .O(gate148inter10));
  nor2  gate656(.a(gate148inter10), .b(gate148inter9), .O(gate148inter11));
  nor2  gate657(.a(gate148inter11), .b(gate148inter6), .O(gate148inter12));
  nand2 gate658(.a(gate148inter12), .b(gate148inter1), .O(G555));
nand2 gate149( .a(G498), .b(G501), .O(G558) );
nand2 gate150( .a(G504), .b(G507), .O(G561) );

  xor2  gate659(.a(G513), .b(G510), .O(gate151inter0));
  nand2 gate660(.a(gate151inter0), .b(s_16), .O(gate151inter1));
  and2  gate661(.a(G513), .b(G510), .O(gate151inter2));
  inv1  gate662(.a(s_16), .O(gate151inter3));
  inv1  gate663(.a(s_17), .O(gate151inter4));
  nand2 gate664(.a(gate151inter4), .b(gate151inter3), .O(gate151inter5));
  nor2  gate665(.a(gate151inter5), .b(gate151inter2), .O(gate151inter6));
  inv1  gate666(.a(G510), .O(gate151inter7));
  inv1  gate667(.a(G513), .O(gate151inter8));
  nand2 gate668(.a(gate151inter8), .b(gate151inter7), .O(gate151inter9));
  nand2 gate669(.a(s_17), .b(gate151inter3), .O(gate151inter10));
  nor2  gate670(.a(gate151inter10), .b(gate151inter9), .O(gate151inter11));
  nor2  gate671(.a(gate151inter11), .b(gate151inter6), .O(gate151inter12));
  nand2 gate672(.a(gate151inter12), .b(gate151inter1), .O(G564));
nand2 gate152( .a(G516), .b(G519), .O(G567) );
nand2 gate153( .a(G426), .b(G522), .O(G570) );
nand2 gate154( .a(G429), .b(G522), .O(G571) );
nand2 gate155( .a(G432), .b(G525), .O(G572) );
nand2 gate156( .a(G435), .b(G525), .O(G573) );
nand2 gate157( .a(G438), .b(G528), .O(G574) );
nand2 gate158( .a(G441), .b(G528), .O(G575) );
nand2 gate159( .a(G444), .b(G531), .O(G576) );
nand2 gate160( .a(G447), .b(G531), .O(G577) );
nand2 gate161( .a(G450), .b(G534), .O(G578) );
nand2 gate162( .a(G453), .b(G534), .O(G579) );
nand2 gate163( .a(G456), .b(G537), .O(G580) );
nand2 gate164( .a(G459), .b(G537), .O(G581) );

  xor2  gate547(.a(G540), .b(G462), .O(gate165inter0));
  nand2 gate548(.a(gate165inter0), .b(s_0), .O(gate165inter1));
  and2  gate549(.a(G540), .b(G462), .O(gate165inter2));
  inv1  gate550(.a(s_0), .O(gate165inter3));
  inv1  gate551(.a(s_1), .O(gate165inter4));
  nand2 gate552(.a(gate165inter4), .b(gate165inter3), .O(gate165inter5));
  nor2  gate553(.a(gate165inter5), .b(gate165inter2), .O(gate165inter6));
  inv1  gate554(.a(G462), .O(gate165inter7));
  inv1  gate555(.a(G540), .O(gate165inter8));
  nand2 gate556(.a(gate165inter8), .b(gate165inter7), .O(gate165inter9));
  nand2 gate557(.a(s_1), .b(gate165inter3), .O(gate165inter10));
  nor2  gate558(.a(gate165inter10), .b(gate165inter9), .O(gate165inter11));
  nor2  gate559(.a(gate165inter11), .b(gate165inter6), .O(gate165inter12));
  nand2 gate560(.a(gate165inter12), .b(gate165inter1), .O(G582));
nand2 gate166( .a(G465), .b(G540), .O(G583) );
nand2 gate167( .a(G468), .b(G543), .O(G584) );
nand2 gate168( .a(G471), .b(G543), .O(G585) );
nand2 gate169( .a(G474), .b(G546), .O(G586) );
nand2 gate170( .a(G477), .b(G546), .O(G587) );
nand2 gate171( .a(G480), .b(G549), .O(G588) );
nand2 gate172( .a(G483), .b(G549), .O(G589) );
nand2 gate173( .a(G486), .b(G552), .O(G590) );
nand2 gate174( .a(G489), .b(G552), .O(G591) );
nand2 gate175( .a(G492), .b(G555), .O(G592) );

  xor2  gate1107(.a(G555), .b(G495), .O(gate176inter0));
  nand2 gate1108(.a(gate176inter0), .b(s_80), .O(gate176inter1));
  and2  gate1109(.a(G555), .b(G495), .O(gate176inter2));
  inv1  gate1110(.a(s_80), .O(gate176inter3));
  inv1  gate1111(.a(s_81), .O(gate176inter4));
  nand2 gate1112(.a(gate176inter4), .b(gate176inter3), .O(gate176inter5));
  nor2  gate1113(.a(gate176inter5), .b(gate176inter2), .O(gate176inter6));
  inv1  gate1114(.a(G495), .O(gate176inter7));
  inv1  gate1115(.a(G555), .O(gate176inter8));
  nand2 gate1116(.a(gate176inter8), .b(gate176inter7), .O(gate176inter9));
  nand2 gate1117(.a(s_81), .b(gate176inter3), .O(gate176inter10));
  nor2  gate1118(.a(gate176inter10), .b(gate176inter9), .O(gate176inter11));
  nor2  gate1119(.a(gate176inter11), .b(gate176inter6), .O(gate176inter12));
  nand2 gate1120(.a(gate176inter12), .b(gate176inter1), .O(G593));
nand2 gate177( .a(G498), .b(G558), .O(G594) );
nand2 gate178( .a(G501), .b(G558), .O(G595) );
nand2 gate179( .a(G504), .b(G561), .O(G596) );
nand2 gate180( .a(G507), .b(G561), .O(G597) );
nand2 gate181( .a(G510), .b(G564), .O(G598) );
nand2 gate182( .a(G513), .b(G564), .O(G599) );
nand2 gate183( .a(G516), .b(G567), .O(G600) );

  xor2  gate1009(.a(G567), .b(G519), .O(gate184inter0));
  nand2 gate1010(.a(gate184inter0), .b(s_66), .O(gate184inter1));
  and2  gate1011(.a(G567), .b(G519), .O(gate184inter2));
  inv1  gate1012(.a(s_66), .O(gate184inter3));
  inv1  gate1013(.a(s_67), .O(gate184inter4));
  nand2 gate1014(.a(gate184inter4), .b(gate184inter3), .O(gate184inter5));
  nor2  gate1015(.a(gate184inter5), .b(gate184inter2), .O(gate184inter6));
  inv1  gate1016(.a(G519), .O(gate184inter7));
  inv1  gate1017(.a(G567), .O(gate184inter8));
  nand2 gate1018(.a(gate184inter8), .b(gate184inter7), .O(gate184inter9));
  nand2 gate1019(.a(s_67), .b(gate184inter3), .O(gate184inter10));
  nor2  gate1020(.a(gate184inter10), .b(gate184inter9), .O(gate184inter11));
  nor2  gate1021(.a(gate184inter11), .b(gate184inter6), .O(gate184inter12));
  nand2 gate1022(.a(gate184inter12), .b(gate184inter1), .O(G601));

  xor2  gate1121(.a(G571), .b(G570), .O(gate185inter0));
  nand2 gate1122(.a(gate185inter0), .b(s_82), .O(gate185inter1));
  and2  gate1123(.a(G571), .b(G570), .O(gate185inter2));
  inv1  gate1124(.a(s_82), .O(gate185inter3));
  inv1  gate1125(.a(s_83), .O(gate185inter4));
  nand2 gate1126(.a(gate185inter4), .b(gate185inter3), .O(gate185inter5));
  nor2  gate1127(.a(gate185inter5), .b(gate185inter2), .O(gate185inter6));
  inv1  gate1128(.a(G570), .O(gate185inter7));
  inv1  gate1129(.a(G571), .O(gate185inter8));
  nand2 gate1130(.a(gate185inter8), .b(gate185inter7), .O(gate185inter9));
  nand2 gate1131(.a(s_83), .b(gate185inter3), .O(gate185inter10));
  nor2  gate1132(.a(gate185inter10), .b(gate185inter9), .O(gate185inter11));
  nor2  gate1133(.a(gate185inter11), .b(gate185inter6), .O(gate185inter12));
  nand2 gate1134(.a(gate185inter12), .b(gate185inter1), .O(G602));
nand2 gate186( .a(G572), .b(G573), .O(G607) );

  xor2  gate911(.a(G575), .b(G574), .O(gate187inter0));
  nand2 gate912(.a(gate187inter0), .b(s_52), .O(gate187inter1));
  and2  gate913(.a(G575), .b(G574), .O(gate187inter2));
  inv1  gate914(.a(s_52), .O(gate187inter3));
  inv1  gate915(.a(s_53), .O(gate187inter4));
  nand2 gate916(.a(gate187inter4), .b(gate187inter3), .O(gate187inter5));
  nor2  gate917(.a(gate187inter5), .b(gate187inter2), .O(gate187inter6));
  inv1  gate918(.a(G574), .O(gate187inter7));
  inv1  gate919(.a(G575), .O(gate187inter8));
  nand2 gate920(.a(gate187inter8), .b(gate187inter7), .O(gate187inter9));
  nand2 gate921(.a(s_53), .b(gate187inter3), .O(gate187inter10));
  nor2  gate922(.a(gate187inter10), .b(gate187inter9), .O(gate187inter11));
  nor2  gate923(.a(gate187inter11), .b(gate187inter6), .O(gate187inter12));
  nand2 gate924(.a(gate187inter12), .b(gate187inter1), .O(G612));
nand2 gate188( .a(G576), .b(G577), .O(G617) );
nand2 gate189( .a(G578), .b(G579), .O(G622) );
nand2 gate190( .a(G580), .b(G581), .O(G627) );

  xor2  gate1485(.a(G583), .b(G582), .O(gate191inter0));
  nand2 gate1486(.a(gate191inter0), .b(s_134), .O(gate191inter1));
  and2  gate1487(.a(G583), .b(G582), .O(gate191inter2));
  inv1  gate1488(.a(s_134), .O(gate191inter3));
  inv1  gate1489(.a(s_135), .O(gate191inter4));
  nand2 gate1490(.a(gate191inter4), .b(gate191inter3), .O(gate191inter5));
  nor2  gate1491(.a(gate191inter5), .b(gate191inter2), .O(gate191inter6));
  inv1  gate1492(.a(G582), .O(gate191inter7));
  inv1  gate1493(.a(G583), .O(gate191inter8));
  nand2 gate1494(.a(gate191inter8), .b(gate191inter7), .O(gate191inter9));
  nand2 gate1495(.a(s_135), .b(gate191inter3), .O(gate191inter10));
  nor2  gate1496(.a(gate191inter10), .b(gate191inter9), .O(gate191inter11));
  nor2  gate1497(.a(gate191inter11), .b(gate191inter6), .O(gate191inter12));
  nand2 gate1498(.a(gate191inter12), .b(gate191inter1), .O(G632));

  xor2  gate1443(.a(G585), .b(G584), .O(gate192inter0));
  nand2 gate1444(.a(gate192inter0), .b(s_128), .O(gate192inter1));
  and2  gate1445(.a(G585), .b(G584), .O(gate192inter2));
  inv1  gate1446(.a(s_128), .O(gate192inter3));
  inv1  gate1447(.a(s_129), .O(gate192inter4));
  nand2 gate1448(.a(gate192inter4), .b(gate192inter3), .O(gate192inter5));
  nor2  gate1449(.a(gate192inter5), .b(gate192inter2), .O(gate192inter6));
  inv1  gate1450(.a(G584), .O(gate192inter7));
  inv1  gate1451(.a(G585), .O(gate192inter8));
  nand2 gate1452(.a(gate192inter8), .b(gate192inter7), .O(gate192inter9));
  nand2 gate1453(.a(s_129), .b(gate192inter3), .O(gate192inter10));
  nor2  gate1454(.a(gate192inter10), .b(gate192inter9), .O(gate192inter11));
  nor2  gate1455(.a(gate192inter11), .b(gate192inter6), .O(gate192inter12));
  nand2 gate1456(.a(gate192inter12), .b(gate192inter1), .O(G637));
nand2 gate193( .a(G586), .b(G587), .O(G642) );
nand2 gate194( .a(G588), .b(G589), .O(G645) );
nand2 gate195( .a(G590), .b(G591), .O(G648) );
nand2 gate196( .a(G592), .b(G593), .O(G651) );
nand2 gate197( .a(G594), .b(G595), .O(G654) );
nand2 gate198( .a(G596), .b(G597), .O(G657) );
nand2 gate199( .a(G598), .b(G599), .O(G660) );
nand2 gate200( .a(G600), .b(G601), .O(G663) );
nand2 gate201( .a(G602), .b(G607), .O(G666) );
nand2 gate202( .a(G612), .b(G617), .O(G669) );
nand2 gate203( .a(G602), .b(G612), .O(G672) );

  xor2  gate1471(.a(G617), .b(G607), .O(gate204inter0));
  nand2 gate1472(.a(gate204inter0), .b(s_132), .O(gate204inter1));
  and2  gate1473(.a(G617), .b(G607), .O(gate204inter2));
  inv1  gate1474(.a(s_132), .O(gate204inter3));
  inv1  gate1475(.a(s_133), .O(gate204inter4));
  nand2 gate1476(.a(gate204inter4), .b(gate204inter3), .O(gate204inter5));
  nor2  gate1477(.a(gate204inter5), .b(gate204inter2), .O(gate204inter6));
  inv1  gate1478(.a(G607), .O(gate204inter7));
  inv1  gate1479(.a(G617), .O(gate204inter8));
  nand2 gate1480(.a(gate204inter8), .b(gate204inter7), .O(gate204inter9));
  nand2 gate1481(.a(s_133), .b(gate204inter3), .O(gate204inter10));
  nor2  gate1482(.a(gate204inter10), .b(gate204inter9), .O(gate204inter11));
  nor2  gate1483(.a(gate204inter11), .b(gate204inter6), .O(gate204inter12));
  nand2 gate1484(.a(gate204inter12), .b(gate204inter1), .O(G675));
nand2 gate205( .a(G622), .b(G627), .O(G678) );

  xor2  gate701(.a(G637), .b(G632), .O(gate206inter0));
  nand2 gate702(.a(gate206inter0), .b(s_22), .O(gate206inter1));
  and2  gate703(.a(G637), .b(G632), .O(gate206inter2));
  inv1  gate704(.a(s_22), .O(gate206inter3));
  inv1  gate705(.a(s_23), .O(gate206inter4));
  nand2 gate706(.a(gate206inter4), .b(gate206inter3), .O(gate206inter5));
  nor2  gate707(.a(gate206inter5), .b(gate206inter2), .O(gate206inter6));
  inv1  gate708(.a(G632), .O(gate206inter7));
  inv1  gate709(.a(G637), .O(gate206inter8));
  nand2 gate710(.a(gate206inter8), .b(gate206inter7), .O(gate206inter9));
  nand2 gate711(.a(s_23), .b(gate206inter3), .O(gate206inter10));
  nor2  gate712(.a(gate206inter10), .b(gate206inter9), .O(gate206inter11));
  nor2  gate713(.a(gate206inter11), .b(gate206inter6), .O(gate206inter12));
  nand2 gate714(.a(gate206inter12), .b(gate206inter1), .O(G681));
nand2 gate207( .a(G622), .b(G632), .O(G684) );
nand2 gate208( .a(G627), .b(G637), .O(G687) );
nand2 gate209( .a(G602), .b(G666), .O(G690) );

  xor2  gate673(.a(G666), .b(G607), .O(gate210inter0));
  nand2 gate674(.a(gate210inter0), .b(s_18), .O(gate210inter1));
  and2  gate675(.a(G666), .b(G607), .O(gate210inter2));
  inv1  gate676(.a(s_18), .O(gate210inter3));
  inv1  gate677(.a(s_19), .O(gate210inter4));
  nand2 gate678(.a(gate210inter4), .b(gate210inter3), .O(gate210inter5));
  nor2  gate679(.a(gate210inter5), .b(gate210inter2), .O(gate210inter6));
  inv1  gate680(.a(G607), .O(gate210inter7));
  inv1  gate681(.a(G666), .O(gate210inter8));
  nand2 gate682(.a(gate210inter8), .b(gate210inter7), .O(gate210inter9));
  nand2 gate683(.a(s_19), .b(gate210inter3), .O(gate210inter10));
  nor2  gate684(.a(gate210inter10), .b(gate210inter9), .O(gate210inter11));
  nor2  gate685(.a(gate210inter11), .b(gate210inter6), .O(gate210inter12));
  nand2 gate686(.a(gate210inter12), .b(gate210inter1), .O(G691));
nand2 gate211( .a(G612), .b(G669), .O(G692) );
nand2 gate212( .a(G617), .b(G669), .O(G693) );
nand2 gate213( .a(G602), .b(G672), .O(G694) );

  xor2  gate813(.a(G672), .b(G612), .O(gate214inter0));
  nand2 gate814(.a(gate214inter0), .b(s_38), .O(gate214inter1));
  and2  gate815(.a(G672), .b(G612), .O(gate214inter2));
  inv1  gate816(.a(s_38), .O(gate214inter3));
  inv1  gate817(.a(s_39), .O(gate214inter4));
  nand2 gate818(.a(gate214inter4), .b(gate214inter3), .O(gate214inter5));
  nor2  gate819(.a(gate214inter5), .b(gate214inter2), .O(gate214inter6));
  inv1  gate820(.a(G612), .O(gate214inter7));
  inv1  gate821(.a(G672), .O(gate214inter8));
  nand2 gate822(.a(gate214inter8), .b(gate214inter7), .O(gate214inter9));
  nand2 gate823(.a(s_39), .b(gate214inter3), .O(gate214inter10));
  nor2  gate824(.a(gate214inter10), .b(gate214inter9), .O(gate214inter11));
  nor2  gate825(.a(gate214inter11), .b(gate214inter6), .O(gate214inter12));
  nand2 gate826(.a(gate214inter12), .b(gate214inter1), .O(G695));
nand2 gate215( .a(G607), .b(G675), .O(G696) );
nand2 gate216( .a(G617), .b(G675), .O(G697) );

  xor2  gate729(.a(G678), .b(G622), .O(gate217inter0));
  nand2 gate730(.a(gate217inter0), .b(s_26), .O(gate217inter1));
  and2  gate731(.a(G678), .b(G622), .O(gate217inter2));
  inv1  gate732(.a(s_26), .O(gate217inter3));
  inv1  gate733(.a(s_27), .O(gate217inter4));
  nand2 gate734(.a(gate217inter4), .b(gate217inter3), .O(gate217inter5));
  nor2  gate735(.a(gate217inter5), .b(gate217inter2), .O(gate217inter6));
  inv1  gate736(.a(G622), .O(gate217inter7));
  inv1  gate737(.a(G678), .O(gate217inter8));
  nand2 gate738(.a(gate217inter8), .b(gate217inter7), .O(gate217inter9));
  nand2 gate739(.a(s_27), .b(gate217inter3), .O(gate217inter10));
  nor2  gate740(.a(gate217inter10), .b(gate217inter9), .O(gate217inter11));
  nor2  gate741(.a(gate217inter11), .b(gate217inter6), .O(gate217inter12));
  nand2 gate742(.a(gate217inter12), .b(gate217inter1), .O(G698));
nand2 gate218( .a(G627), .b(G678), .O(G699) );
nand2 gate219( .a(G632), .b(G681), .O(G700) );
nand2 gate220( .a(G637), .b(G681), .O(G701) );
nand2 gate221( .a(G622), .b(G684), .O(G702) );
nand2 gate222( .a(G632), .b(G684), .O(G703) );
nand2 gate223( .a(G627), .b(G687), .O(G704) );
nand2 gate224( .a(G637), .b(G687), .O(G705) );
nand2 gate225( .a(G690), .b(G691), .O(G706) );
nand2 gate226( .a(G692), .b(G693), .O(G709) );
nand2 gate227( .a(G694), .b(G695), .O(G712) );
nand2 gate228( .a(G696), .b(G697), .O(G715) );
nand2 gate229( .a(G698), .b(G699), .O(G718) );
nand2 gate230( .a(G700), .b(G701), .O(G721) );

  xor2  gate1429(.a(G703), .b(G702), .O(gate231inter0));
  nand2 gate1430(.a(gate231inter0), .b(s_126), .O(gate231inter1));
  and2  gate1431(.a(G703), .b(G702), .O(gate231inter2));
  inv1  gate1432(.a(s_126), .O(gate231inter3));
  inv1  gate1433(.a(s_127), .O(gate231inter4));
  nand2 gate1434(.a(gate231inter4), .b(gate231inter3), .O(gate231inter5));
  nor2  gate1435(.a(gate231inter5), .b(gate231inter2), .O(gate231inter6));
  inv1  gate1436(.a(G702), .O(gate231inter7));
  inv1  gate1437(.a(G703), .O(gate231inter8));
  nand2 gate1438(.a(gate231inter8), .b(gate231inter7), .O(gate231inter9));
  nand2 gate1439(.a(s_127), .b(gate231inter3), .O(gate231inter10));
  nor2  gate1440(.a(gate231inter10), .b(gate231inter9), .O(gate231inter11));
  nor2  gate1441(.a(gate231inter11), .b(gate231inter6), .O(gate231inter12));
  nand2 gate1442(.a(gate231inter12), .b(gate231inter1), .O(G724));
nand2 gate232( .a(G704), .b(G705), .O(G727) );

  xor2  gate1373(.a(G718), .b(G242), .O(gate233inter0));
  nand2 gate1374(.a(gate233inter0), .b(s_118), .O(gate233inter1));
  and2  gate1375(.a(G718), .b(G242), .O(gate233inter2));
  inv1  gate1376(.a(s_118), .O(gate233inter3));
  inv1  gate1377(.a(s_119), .O(gate233inter4));
  nand2 gate1378(.a(gate233inter4), .b(gate233inter3), .O(gate233inter5));
  nor2  gate1379(.a(gate233inter5), .b(gate233inter2), .O(gate233inter6));
  inv1  gate1380(.a(G242), .O(gate233inter7));
  inv1  gate1381(.a(G718), .O(gate233inter8));
  nand2 gate1382(.a(gate233inter8), .b(gate233inter7), .O(gate233inter9));
  nand2 gate1383(.a(s_119), .b(gate233inter3), .O(gate233inter10));
  nor2  gate1384(.a(gate233inter10), .b(gate233inter9), .O(gate233inter11));
  nor2  gate1385(.a(gate233inter11), .b(gate233inter6), .O(gate233inter12));
  nand2 gate1386(.a(gate233inter12), .b(gate233inter1), .O(G730));
nand2 gate234( .a(G245), .b(G721), .O(G733) );
nand2 gate235( .a(G248), .b(G724), .O(G736) );
nand2 gate236( .a(G251), .b(G727), .O(G739) );
nand2 gate237( .a(G254), .b(G706), .O(G742) );
nand2 gate238( .a(G257), .b(G709), .O(G745) );
nand2 gate239( .a(G260), .b(G712), .O(G748) );
nand2 gate240( .a(G263), .b(G715), .O(G751) );
nand2 gate241( .a(G242), .b(G730), .O(G754) );
nand2 gate242( .a(G718), .b(G730), .O(G755) );

  xor2  gate743(.a(G733), .b(G245), .O(gate243inter0));
  nand2 gate744(.a(gate243inter0), .b(s_28), .O(gate243inter1));
  and2  gate745(.a(G733), .b(G245), .O(gate243inter2));
  inv1  gate746(.a(s_28), .O(gate243inter3));
  inv1  gate747(.a(s_29), .O(gate243inter4));
  nand2 gate748(.a(gate243inter4), .b(gate243inter3), .O(gate243inter5));
  nor2  gate749(.a(gate243inter5), .b(gate243inter2), .O(gate243inter6));
  inv1  gate750(.a(G245), .O(gate243inter7));
  inv1  gate751(.a(G733), .O(gate243inter8));
  nand2 gate752(.a(gate243inter8), .b(gate243inter7), .O(gate243inter9));
  nand2 gate753(.a(s_29), .b(gate243inter3), .O(gate243inter10));
  nor2  gate754(.a(gate243inter10), .b(gate243inter9), .O(gate243inter11));
  nor2  gate755(.a(gate243inter11), .b(gate243inter6), .O(gate243inter12));
  nand2 gate756(.a(gate243inter12), .b(gate243inter1), .O(G756));
nand2 gate244( .a(G721), .b(G733), .O(G757) );
nand2 gate245( .a(G248), .b(G736), .O(G758) );
nand2 gate246( .a(G724), .b(G736), .O(G759) );
nand2 gate247( .a(G251), .b(G739), .O(G760) );

  xor2  gate631(.a(G739), .b(G727), .O(gate248inter0));
  nand2 gate632(.a(gate248inter0), .b(s_12), .O(gate248inter1));
  and2  gate633(.a(G739), .b(G727), .O(gate248inter2));
  inv1  gate634(.a(s_12), .O(gate248inter3));
  inv1  gate635(.a(s_13), .O(gate248inter4));
  nand2 gate636(.a(gate248inter4), .b(gate248inter3), .O(gate248inter5));
  nor2  gate637(.a(gate248inter5), .b(gate248inter2), .O(gate248inter6));
  inv1  gate638(.a(G727), .O(gate248inter7));
  inv1  gate639(.a(G739), .O(gate248inter8));
  nand2 gate640(.a(gate248inter8), .b(gate248inter7), .O(gate248inter9));
  nand2 gate641(.a(s_13), .b(gate248inter3), .O(gate248inter10));
  nor2  gate642(.a(gate248inter10), .b(gate248inter9), .O(gate248inter11));
  nor2  gate643(.a(gate248inter11), .b(gate248inter6), .O(gate248inter12));
  nand2 gate644(.a(gate248inter12), .b(gate248inter1), .O(G761));
nand2 gate249( .a(G254), .b(G742), .O(G762) );

  xor2  gate785(.a(G742), .b(G706), .O(gate250inter0));
  nand2 gate786(.a(gate250inter0), .b(s_34), .O(gate250inter1));
  and2  gate787(.a(G742), .b(G706), .O(gate250inter2));
  inv1  gate788(.a(s_34), .O(gate250inter3));
  inv1  gate789(.a(s_35), .O(gate250inter4));
  nand2 gate790(.a(gate250inter4), .b(gate250inter3), .O(gate250inter5));
  nor2  gate791(.a(gate250inter5), .b(gate250inter2), .O(gate250inter6));
  inv1  gate792(.a(G706), .O(gate250inter7));
  inv1  gate793(.a(G742), .O(gate250inter8));
  nand2 gate794(.a(gate250inter8), .b(gate250inter7), .O(gate250inter9));
  nand2 gate795(.a(s_35), .b(gate250inter3), .O(gate250inter10));
  nor2  gate796(.a(gate250inter10), .b(gate250inter9), .O(gate250inter11));
  nor2  gate797(.a(gate250inter11), .b(gate250inter6), .O(gate250inter12));
  nand2 gate798(.a(gate250inter12), .b(gate250inter1), .O(G763));

  xor2  gate589(.a(G745), .b(G257), .O(gate251inter0));
  nand2 gate590(.a(gate251inter0), .b(s_6), .O(gate251inter1));
  and2  gate591(.a(G745), .b(G257), .O(gate251inter2));
  inv1  gate592(.a(s_6), .O(gate251inter3));
  inv1  gate593(.a(s_7), .O(gate251inter4));
  nand2 gate594(.a(gate251inter4), .b(gate251inter3), .O(gate251inter5));
  nor2  gate595(.a(gate251inter5), .b(gate251inter2), .O(gate251inter6));
  inv1  gate596(.a(G257), .O(gate251inter7));
  inv1  gate597(.a(G745), .O(gate251inter8));
  nand2 gate598(.a(gate251inter8), .b(gate251inter7), .O(gate251inter9));
  nand2 gate599(.a(s_7), .b(gate251inter3), .O(gate251inter10));
  nor2  gate600(.a(gate251inter10), .b(gate251inter9), .O(gate251inter11));
  nor2  gate601(.a(gate251inter11), .b(gate251inter6), .O(gate251inter12));
  nand2 gate602(.a(gate251inter12), .b(gate251inter1), .O(G764));
nand2 gate252( .a(G709), .b(G745), .O(G765) );
nand2 gate253( .a(G260), .b(G748), .O(G766) );
nand2 gate254( .a(G712), .b(G748), .O(G767) );
nand2 gate255( .a(G263), .b(G751), .O(G768) );
nand2 gate256( .a(G715), .b(G751), .O(G769) );
nand2 gate257( .a(G754), .b(G755), .O(G770) );
nand2 gate258( .a(G756), .b(G757), .O(G773) );

  xor2  gate1345(.a(G759), .b(G758), .O(gate259inter0));
  nand2 gate1346(.a(gate259inter0), .b(s_114), .O(gate259inter1));
  and2  gate1347(.a(G759), .b(G758), .O(gate259inter2));
  inv1  gate1348(.a(s_114), .O(gate259inter3));
  inv1  gate1349(.a(s_115), .O(gate259inter4));
  nand2 gate1350(.a(gate259inter4), .b(gate259inter3), .O(gate259inter5));
  nor2  gate1351(.a(gate259inter5), .b(gate259inter2), .O(gate259inter6));
  inv1  gate1352(.a(G758), .O(gate259inter7));
  inv1  gate1353(.a(G759), .O(gate259inter8));
  nand2 gate1354(.a(gate259inter8), .b(gate259inter7), .O(gate259inter9));
  nand2 gate1355(.a(s_115), .b(gate259inter3), .O(gate259inter10));
  nor2  gate1356(.a(gate259inter10), .b(gate259inter9), .O(gate259inter11));
  nor2  gate1357(.a(gate259inter11), .b(gate259inter6), .O(gate259inter12));
  nand2 gate1358(.a(gate259inter12), .b(gate259inter1), .O(G776));
nand2 gate260( .a(G760), .b(G761), .O(G779) );
nand2 gate261( .a(G762), .b(G763), .O(G782) );
nand2 gate262( .a(G764), .b(G765), .O(G785) );
nand2 gate263( .a(G766), .b(G767), .O(G788) );

  xor2  gate1261(.a(G769), .b(G768), .O(gate264inter0));
  nand2 gate1262(.a(gate264inter0), .b(s_102), .O(gate264inter1));
  and2  gate1263(.a(G769), .b(G768), .O(gate264inter2));
  inv1  gate1264(.a(s_102), .O(gate264inter3));
  inv1  gate1265(.a(s_103), .O(gate264inter4));
  nand2 gate1266(.a(gate264inter4), .b(gate264inter3), .O(gate264inter5));
  nor2  gate1267(.a(gate264inter5), .b(gate264inter2), .O(gate264inter6));
  inv1  gate1268(.a(G768), .O(gate264inter7));
  inv1  gate1269(.a(G769), .O(gate264inter8));
  nand2 gate1270(.a(gate264inter8), .b(gate264inter7), .O(gate264inter9));
  nand2 gate1271(.a(s_103), .b(gate264inter3), .O(gate264inter10));
  nor2  gate1272(.a(gate264inter10), .b(gate264inter9), .O(gate264inter11));
  nor2  gate1273(.a(gate264inter11), .b(gate264inter6), .O(gate264inter12));
  nand2 gate1274(.a(gate264inter12), .b(gate264inter1), .O(G791));
nand2 gate265( .a(G642), .b(G770), .O(G794) );
nand2 gate266( .a(G645), .b(G773), .O(G797) );

  xor2  gate1037(.a(G776), .b(G648), .O(gate267inter0));
  nand2 gate1038(.a(gate267inter0), .b(s_70), .O(gate267inter1));
  and2  gate1039(.a(G776), .b(G648), .O(gate267inter2));
  inv1  gate1040(.a(s_70), .O(gate267inter3));
  inv1  gate1041(.a(s_71), .O(gate267inter4));
  nand2 gate1042(.a(gate267inter4), .b(gate267inter3), .O(gate267inter5));
  nor2  gate1043(.a(gate267inter5), .b(gate267inter2), .O(gate267inter6));
  inv1  gate1044(.a(G648), .O(gate267inter7));
  inv1  gate1045(.a(G776), .O(gate267inter8));
  nand2 gate1046(.a(gate267inter8), .b(gate267inter7), .O(gate267inter9));
  nand2 gate1047(.a(s_71), .b(gate267inter3), .O(gate267inter10));
  nor2  gate1048(.a(gate267inter10), .b(gate267inter9), .O(gate267inter11));
  nor2  gate1049(.a(gate267inter11), .b(gate267inter6), .O(gate267inter12));
  nand2 gate1050(.a(gate267inter12), .b(gate267inter1), .O(G800));
nand2 gate268( .a(G651), .b(G779), .O(G803) );
nand2 gate269( .a(G654), .b(G782), .O(G806) );
nand2 gate270( .a(G657), .b(G785), .O(G809) );
nand2 gate271( .a(G660), .b(G788), .O(G812) );

  xor2  gate715(.a(G791), .b(G663), .O(gate272inter0));
  nand2 gate716(.a(gate272inter0), .b(s_24), .O(gate272inter1));
  and2  gate717(.a(G791), .b(G663), .O(gate272inter2));
  inv1  gate718(.a(s_24), .O(gate272inter3));
  inv1  gate719(.a(s_25), .O(gate272inter4));
  nand2 gate720(.a(gate272inter4), .b(gate272inter3), .O(gate272inter5));
  nor2  gate721(.a(gate272inter5), .b(gate272inter2), .O(gate272inter6));
  inv1  gate722(.a(G663), .O(gate272inter7));
  inv1  gate723(.a(G791), .O(gate272inter8));
  nand2 gate724(.a(gate272inter8), .b(gate272inter7), .O(gate272inter9));
  nand2 gate725(.a(s_25), .b(gate272inter3), .O(gate272inter10));
  nor2  gate726(.a(gate272inter10), .b(gate272inter9), .O(gate272inter11));
  nor2  gate727(.a(gate272inter11), .b(gate272inter6), .O(gate272inter12));
  nand2 gate728(.a(gate272inter12), .b(gate272inter1), .O(G815));
nand2 gate273( .a(G642), .b(G794), .O(G818) );
nand2 gate274( .a(G770), .b(G794), .O(G819) );
nand2 gate275( .a(G645), .b(G797), .O(G820) );
nand2 gate276( .a(G773), .b(G797), .O(G821) );
nand2 gate277( .a(G648), .b(G800), .O(G822) );

  xor2  gate1163(.a(G800), .b(G776), .O(gate278inter0));
  nand2 gate1164(.a(gate278inter0), .b(s_88), .O(gate278inter1));
  and2  gate1165(.a(G800), .b(G776), .O(gate278inter2));
  inv1  gate1166(.a(s_88), .O(gate278inter3));
  inv1  gate1167(.a(s_89), .O(gate278inter4));
  nand2 gate1168(.a(gate278inter4), .b(gate278inter3), .O(gate278inter5));
  nor2  gate1169(.a(gate278inter5), .b(gate278inter2), .O(gate278inter6));
  inv1  gate1170(.a(G776), .O(gate278inter7));
  inv1  gate1171(.a(G800), .O(gate278inter8));
  nand2 gate1172(.a(gate278inter8), .b(gate278inter7), .O(gate278inter9));
  nand2 gate1173(.a(s_89), .b(gate278inter3), .O(gate278inter10));
  nor2  gate1174(.a(gate278inter10), .b(gate278inter9), .O(gate278inter11));
  nor2  gate1175(.a(gate278inter11), .b(gate278inter6), .O(gate278inter12));
  nand2 gate1176(.a(gate278inter12), .b(gate278inter1), .O(G823));
nand2 gate279( .a(G651), .b(G803), .O(G824) );
nand2 gate280( .a(G779), .b(G803), .O(G825) );
nand2 gate281( .a(G654), .b(G806), .O(G826) );
nand2 gate282( .a(G782), .b(G806), .O(G827) );
nand2 gate283( .a(G657), .b(G809), .O(G828) );
nand2 gate284( .a(G785), .b(G809), .O(G829) );
nand2 gate285( .a(G660), .b(G812), .O(G830) );
nand2 gate286( .a(G788), .b(G812), .O(G831) );
nand2 gate287( .a(G663), .b(G815), .O(G832) );

  xor2  gate1149(.a(G815), .b(G791), .O(gate288inter0));
  nand2 gate1150(.a(gate288inter0), .b(s_86), .O(gate288inter1));
  and2  gate1151(.a(G815), .b(G791), .O(gate288inter2));
  inv1  gate1152(.a(s_86), .O(gate288inter3));
  inv1  gate1153(.a(s_87), .O(gate288inter4));
  nand2 gate1154(.a(gate288inter4), .b(gate288inter3), .O(gate288inter5));
  nor2  gate1155(.a(gate288inter5), .b(gate288inter2), .O(gate288inter6));
  inv1  gate1156(.a(G791), .O(gate288inter7));
  inv1  gate1157(.a(G815), .O(gate288inter8));
  nand2 gate1158(.a(gate288inter8), .b(gate288inter7), .O(gate288inter9));
  nand2 gate1159(.a(s_87), .b(gate288inter3), .O(gate288inter10));
  nor2  gate1160(.a(gate288inter10), .b(gate288inter9), .O(gate288inter11));
  nor2  gate1161(.a(gate288inter11), .b(gate288inter6), .O(gate288inter12));
  nand2 gate1162(.a(gate288inter12), .b(gate288inter1), .O(G833));
nand2 gate289( .a(G818), .b(G819), .O(G834) );
nand2 gate290( .a(G820), .b(G821), .O(G847) );
nand2 gate291( .a(G822), .b(G823), .O(G860) );

  xor2  gate1233(.a(G825), .b(G824), .O(gate292inter0));
  nand2 gate1234(.a(gate292inter0), .b(s_98), .O(gate292inter1));
  and2  gate1235(.a(G825), .b(G824), .O(gate292inter2));
  inv1  gate1236(.a(s_98), .O(gate292inter3));
  inv1  gate1237(.a(s_99), .O(gate292inter4));
  nand2 gate1238(.a(gate292inter4), .b(gate292inter3), .O(gate292inter5));
  nor2  gate1239(.a(gate292inter5), .b(gate292inter2), .O(gate292inter6));
  inv1  gate1240(.a(G824), .O(gate292inter7));
  inv1  gate1241(.a(G825), .O(gate292inter8));
  nand2 gate1242(.a(gate292inter8), .b(gate292inter7), .O(gate292inter9));
  nand2 gate1243(.a(s_99), .b(gate292inter3), .O(gate292inter10));
  nor2  gate1244(.a(gate292inter10), .b(gate292inter9), .O(gate292inter11));
  nor2  gate1245(.a(gate292inter11), .b(gate292inter6), .O(gate292inter12));
  nand2 gate1246(.a(gate292inter12), .b(gate292inter1), .O(G873));
nand2 gate293( .a(G828), .b(G829), .O(G886) );
nand2 gate294( .a(G832), .b(G833), .O(G899) );

  xor2  gate1219(.a(G831), .b(G830), .O(gate295inter0));
  nand2 gate1220(.a(gate295inter0), .b(s_96), .O(gate295inter1));
  and2  gate1221(.a(G831), .b(G830), .O(gate295inter2));
  inv1  gate1222(.a(s_96), .O(gate295inter3));
  inv1  gate1223(.a(s_97), .O(gate295inter4));
  nand2 gate1224(.a(gate295inter4), .b(gate295inter3), .O(gate295inter5));
  nor2  gate1225(.a(gate295inter5), .b(gate295inter2), .O(gate295inter6));
  inv1  gate1226(.a(G830), .O(gate295inter7));
  inv1  gate1227(.a(G831), .O(gate295inter8));
  nand2 gate1228(.a(gate295inter8), .b(gate295inter7), .O(gate295inter9));
  nand2 gate1229(.a(s_97), .b(gate295inter3), .O(gate295inter10));
  nor2  gate1230(.a(gate295inter10), .b(gate295inter9), .O(gate295inter11));
  nor2  gate1231(.a(gate295inter11), .b(gate295inter6), .O(gate295inter12));
  nand2 gate1232(.a(gate295inter12), .b(gate295inter1), .O(G912));
nand2 gate296( .a(G826), .b(G827), .O(G925) );
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );
nand2 gate387( .a(G1), .b(G1036), .O(G1132) );
nand2 gate388( .a(G2), .b(G1039), .O(G1135) );
nand2 gate389( .a(G3), .b(G1042), .O(G1138) );

  xor2  gate1317(.a(G1045), .b(G4), .O(gate390inter0));
  nand2 gate1318(.a(gate390inter0), .b(s_110), .O(gate390inter1));
  and2  gate1319(.a(G1045), .b(G4), .O(gate390inter2));
  inv1  gate1320(.a(s_110), .O(gate390inter3));
  inv1  gate1321(.a(s_111), .O(gate390inter4));
  nand2 gate1322(.a(gate390inter4), .b(gate390inter3), .O(gate390inter5));
  nor2  gate1323(.a(gate390inter5), .b(gate390inter2), .O(gate390inter6));
  inv1  gate1324(.a(G4), .O(gate390inter7));
  inv1  gate1325(.a(G1045), .O(gate390inter8));
  nand2 gate1326(.a(gate390inter8), .b(gate390inter7), .O(gate390inter9));
  nand2 gate1327(.a(s_111), .b(gate390inter3), .O(gate390inter10));
  nor2  gate1328(.a(gate390inter10), .b(gate390inter9), .O(gate390inter11));
  nor2  gate1329(.a(gate390inter11), .b(gate390inter6), .O(gate390inter12));
  nand2 gate1330(.a(gate390inter12), .b(gate390inter1), .O(G1141));
nand2 gate391( .a(G5), .b(G1048), .O(G1144) );
nand2 gate392( .a(G6), .b(G1051), .O(G1147) );
nand2 gate393( .a(G7), .b(G1054), .O(G1150) );
nand2 gate394( .a(G8), .b(G1057), .O(G1153) );
nand2 gate395( .a(G9), .b(G1060), .O(G1156) );
nand2 gate396( .a(G10), .b(G1063), .O(G1159) );
nand2 gate397( .a(G11), .b(G1066), .O(G1162) );
nand2 gate398( .a(G12), .b(G1069), .O(G1165) );
nand2 gate399( .a(G13), .b(G1072), .O(G1168) );
nand2 gate400( .a(G14), .b(G1075), .O(G1171) );
nand2 gate401( .a(G15), .b(G1078), .O(G1174) );
nand2 gate402( .a(G16), .b(G1081), .O(G1177) );
nand2 gate403( .a(G17), .b(G1084), .O(G1180) );
nand2 gate404( .a(G18), .b(G1087), .O(G1183) );
nand2 gate405( .a(G19), .b(G1090), .O(G1186) );
nand2 gate406( .a(G20), .b(G1093), .O(G1189) );
nand2 gate407( .a(G21), .b(G1096), .O(G1192) );
nand2 gate408( .a(G22), .b(G1099), .O(G1195) );
nand2 gate409( .a(G23), .b(G1102), .O(G1198) );
nand2 gate410( .a(G24), .b(G1105), .O(G1201) );
nand2 gate411( .a(G25), .b(G1108), .O(G1204) );
nand2 gate412( .a(G26), .b(G1111), .O(G1207) );
nand2 gate413( .a(G27), .b(G1114), .O(G1210) );
nand2 gate414( .a(G28), .b(G1117), .O(G1213) );
nand2 gate415( .a(G29), .b(G1120), .O(G1216) );
nand2 gate416( .a(G30), .b(G1123), .O(G1219) );
nand2 gate417( .a(G31), .b(G1126), .O(G1222) );
nand2 gate418( .a(G32), .b(G1129), .O(G1225) );
nand2 gate419( .a(G1), .b(G1132), .O(G1228) );
nand2 gate420( .a(G1036), .b(G1132), .O(G1229) );
nand2 gate421( .a(G2), .b(G1135), .O(G1230) );
nand2 gate422( .a(G1039), .b(G1135), .O(G1231) );
nand2 gate423( .a(G3), .b(G1138), .O(G1232) );
nand2 gate424( .a(G1042), .b(G1138), .O(G1233) );

  xor2  gate1401(.a(G1141), .b(G4), .O(gate425inter0));
  nand2 gate1402(.a(gate425inter0), .b(s_122), .O(gate425inter1));
  and2  gate1403(.a(G1141), .b(G4), .O(gate425inter2));
  inv1  gate1404(.a(s_122), .O(gate425inter3));
  inv1  gate1405(.a(s_123), .O(gate425inter4));
  nand2 gate1406(.a(gate425inter4), .b(gate425inter3), .O(gate425inter5));
  nor2  gate1407(.a(gate425inter5), .b(gate425inter2), .O(gate425inter6));
  inv1  gate1408(.a(G4), .O(gate425inter7));
  inv1  gate1409(.a(G1141), .O(gate425inter8));
  nand2 gate1410(.a(gate425inter8), .b(gate425inter7), .O(gate425inter9));
  nand2 gate1411(.a(s_123), .b(gate425inter3), .O(gate425inter10));
  nor2  gate1412(.a(gate425inter10), .b(gate425inter9), .O(gate425inter11));
  nor2  gate1413(.a(gate425inter11), .b(gate425inter6), .O(gate425inter12));
  nand2 gate1414(.a(gate425inter12), .b(gate425inter1), .O(G1234));
nand2 gate426( .a(G1045), .b(G1141), .O(G1235) );

  xor2  gate869(.a(G1144), .b(G5), .O(gate427inter0));
  nand2 gate870(.a(gate427inter0), .b(s_46), .O(gate427inter1));
  and2  gate871(.a(G1144), .b(G5), .O(gate427inter2));
  inv1  gate872(.a(s_46), .O(gate427inter3));
  inv1  gate873(.a(s_47), .O(gate427inter4));
  nand2 gate874(.a(gate427inter4), .b(gate427inter3), .O(gate427inter5));
  nor2  gate875(.a(gate427inter5), .b(gate427inter2), .O(gate427inter6));
  inv1  gate876(.a(G5), .O(gate427inter7));
  inv1  gate877(.a(G1144), .O(gate427inter8));
  nand2 gate878(.a(gate427inter8), .b(gate427inter7), .O(gate427inter9));
  nand2 gate879(.a(s_47), .b(gate427inter3), .O(gate427inter10));
  nor2  gate880(.a(gate427inter10), .b(gate427inter9), .O(gate427inter11));
  nor2  gate881(.a(gate427inter11), .b(gate427inter6), .O(gate427inter12));
  nand2 gate882(.a(gate427inter12), .b(gate427inter1), .O(G1236));
nand2 gate428( .a(G1048), .b(G1144), .O(G1237) );
nand2 gate429( .a(G6), .b(G1147), .O(G1238) );
nand2 gate430( .a(G1051), .b(G1147), .O(G1239) );
nand2 gate431( .a(G7), .b(G1150), .O(G1240) );
nand2 gate432( .a(G1054), .b(G1150), .O(G1241) );
nand2 gate433( .a(G8), .b(G1153), .O(G1242) );

  xor2  gate1177(.a(G1153), .b(G1057), .O(gate434inter0));
  nand2 gate1178(.a(gate434inter0), .b(s_90), .O(gate434inter1));
  and2  gate1179(.a(G1153), .b(G1057), .O(gate434inter2));
  inv1  gate1180(.a(s_90), .O(gate434inter3));
  inv1  gate1181(.a(s_91), .O(gate434inter4));
  nand2 gate1182(.a(gate434inter4), .b(gate434inter3), .O(gate434inter5));
  nor2  gate1183(.a(gate434inter5), .b(gate434inter2), .O(gate434inter6));
  inv1  gate1184(.a(G1057), .O(gate434inter7));
  inv1  gate1185(.a(G1153), .O(gate434inter8));
  nand2 gate1186(.a(gate434inter8), .b(gate434inter7), .O(gate434inter9));
  nand2 gate1187(.a(s_91), .b(gate434inter3), .O(gate434inter10));
  nor2  gate1188(.a(gate434inter10), .b(gate434inter9), .O(gate434inter11));
  nor2  gate1189(.a(gate434inter11), .b(gate434inter6), .O(gate434inter12));
  nand2 gate1190(.a(gate434inter12), .b(gate434inter1), .O(G1243));
nand2 gate435( .a(G9), .b(G1156), .O(G1244) );
nand2 gate436( .a(G1060), .b(G1156), .O(G1245) );
nand2 gate437( .a(G10), .b(G1159), .O(G1246) );

  xor2  gate827(.a(G1159), .b(G1063), .O(gate438inter0));
  nand2 gate828(.a(gate438inter0), .b(s_40), .O(gate438inter1));
  and2  gate829(.a(G1159), .b(G1063), .O(gate438inter2));
  inv1  gate830(.a(s_40), .O(gate438inter3));
  inv1  gate831(.a(s_41), .O(gate438inter4));
  nand2 gate832(.a(gate438inter4), .b(gate438inter3), .O(gate438inter5));
  nor2  gate833(.a(gate438inter5), .b(gate438inter2), .O(gate438inter6));
  inv1  gate834(.a(G1063), .O(gate438inter7));
  inv1  gate835(.a(G1159), .O(gate438inter8));
  nand2 gate836(.a(gate438inter8), .b(gate438inter7), .O(gate438inter9));
  nand2 gate837(.a(s_41), .b(gate438inter3), .O(gate438inter10));
  nor2  gate838(.a(gate438inter10), .b(gate438inter9), .O(gate438inter11));
  nor2  gate839(.a(gate438inter11), .b(gate438inter6), .O(gate438inter12));
  nand2 gate840(.a(gate438inter12), .b(gate438inter1), .O(G1247));
nand2 gate439( .a(G11), .b(G1162), .O(G1248) );
nand2 gate440( .a(G1066), .b(G1162), .O(G1249) );

  xor2  gate1513(.a(G1165), .b(G12), .O(gate441inter0));
  nand2 gate1514(.a(gate441inter0), .b(s_138), .O(gate441inter1));
  and2  gate1515(.a(G1165), .b(G12), .O(gate441inter2));
  inv1  gate1516(.a(s_138), .O(gate441inter3));
  inv1  gate1517(.a(s_139), .O(gate441inter4));
  nand2 gate1518(.a(gate441inter4), .b(gate441inter3), .O(gate441inter5));
  nor2  gate1519(.a(gate441inter5), .b(gate441inter2), .O(gate441inter6));
  inv1  gate1520(.a(G12), .O(gate441inter7));
  inv1  gate1521(.a(G1165), .O(gate441inter8));
  nand2 gate1522(.a(gate441inter8), .b(gate441inter7), .O(gate441inter9));
  nand2 gate1523(.a(s_139), .b(gate441inter3), .O(gate441inter10));
  nor2  gate1524(.a(gate441inter10), .b(gate441inter9), .O(gate441inter11));
  nor2  gate1525(.a(gate441inter11), .b(gate441inter6), .O(gate441inter12));
  nand2 gate1526(.a(gate441inter12), .b(gate441inter1), .O(G1250));
nand2 gate442( .a(G1069), .b(G1165), .O(G1251) );
nand2 gate443( .a(G13), .b(G1168), .O(G1252) );
nand2 gate444( .a(G1072), .b(G1168), .O(G1253) );
nand2 gate445( .a(G14), .b(G1171), .O(G1254) );

  xor2  gate1023(.a(G1171), .b(G1075), .O(gate446inter0));
  nand2 gate1024(.a(gate446inter0), .b(s_68), .O(gate446inter1));
  and2  gate1025(.a(G1171), .b(G1075), .O(gate446inter2));
  inv1  gate1026(.a(s_68), .O(gate446inter3));
  inv1  gate1027(.a(s_69), .O(gate446inter4));
  nand2 gate1028(.a(gate446inter4), .b(gate446inter3), .O(gate446inter5));
  nor2  gate1029(.a(gate446inter5), .b(gate446inter2), .O(gate446inter6));
  inv1  gate1030(.a(G1075), .O(gate446inter7));
  inv1  gate1031(.a(G1171), .O(gate446inter8));
  nand2 gate1032(.a(gate446inter8), .b(gate446inter7), .O(gate446inter9));
  nand2 gate1033(.a(s_69), .b(gate446inter3), .O(gate446inter10));
  nor2  gate1034(.a(gate446inter10), .b(gate446inter9), .O(gate446inter11));
  nor2  gate1035(.a(gate446inter11), .b(gate446inter6), .O(gate446inter12));
  nand2 gate1036(.a(gate446inter12), .b(gate446inter1), .O(G1255));
nand2 gate447( .a(G15), .b(G1174), .O(G1256) );
nand2 gate448( .a(G1078), .b(G1174), .O(G1257) );
nand2 gate449( .a(G16), .b(G1177), .O(G1258) );
nand2 gate450( .a(G1081), .b(G1177), .O(G1259) );
nand2 gate451( .a(G17), .b(G1180), .O(G1260) );

  xor2  gate967(.a(G1180), .b(G1084), .O(gate452inter0));
  nand2 gate968(.a(gate452inter0), .b(s_60), .O(gate452inter1));
  and2  gate969(.a(G1180), .b(G1084), .O(gate452inter2));
  inv1  gate970(.a(s_60), .O(gate452inter3));
  inv1  gate971(.a(s_61), .O(gate452inter4));
  nand2 gate972(.a(gate452inter4), .b(gate452inter3), .O(gate452inter5));
  nor2  gate973(.a(gate452inter5), .b(gate452inter2), .O(gate452inter6));
  inv1  gate974(.a(G1084), .O(gate452inter7));
  inv1  gate975(.a(G1180), .O(gate452inter8));
  nand2 gate976(.a(gate452inter8), .b(gate452inter7), .O(gate452inter9));
  nand2 gate977(.a(s_61), .b(gate452inter3), .O(gate452inter10));
  nor2  gate978(.a(gate452inter10), .b(gate452inter9), .O(gate452inter11));
  nor2  gate979(.a(gate452inter11), .b(gate452inter6), .O(gate452inter12));
  nand2 gate980(.a(gate452inter12), .b(gate452inter1), .O(G1261));
nand2 gate453( .a(G18), .b(G1183), .O(G1262) );
nand2 gate454( .a(G1087), .b(G1183), .O(G1263) );

  xor2  gate575(.a(G1186), .b(G19), .O(gate455inter0));
  nand2 gate576(.a(gate455inter0), .b(s_4), .O(gate455inter1));
  and2  gate577(.a(G1186), .b(G19), .O(gate455inter2));
  inv1  gate578(.a(s_4), .O(gate455inter3));
  inv1  gate579(.a(s_5), .O(gate455inter4));
  nand2 gate580(.a(gate455inter4), .b(gate455inter3), .O(gate455inter5));
  nor2  gate581(.a(gate455inter5), .b(gate455inter2), .O(gate455inter6));
  inv1  gate582(.a(G19), .O(gate455inter7));
  inv1  gate583(.a(G1186), .O(gate455inter8));
  nand2 gate584(.a(gate455inter8), .b(gate455inter7), .O(gate455inter9));
  nand2 gate585(.a(s_5), .b(gate455inter3), .O(gate455inter10));
  nor2  gate586(.a(gate455inter10), .b(gate455inter9), .O(gate455inter11));
  nor2  gate587(.a(gate455inter11), .b(gate455inter6), .O(gate455inter12));
  nand2 gate588(.a(gate455inter12), .b(gate455inter1), .O(G1264));
nand2 gate456( .a(G1090), .b(G1186), .O(G1265) );
nand2 gate457( .a(G20), .b(G1189), .O(G1266) );
nand2 gate458( .a(G1093), .b(G1189), .O(G1267) );

  xor2  gate1051(.a(G1192), .b(G21), .O(gate459inter0));
  nand2 gate1052(.a(gate459inter0), .b(s_72), .O(gate459inter1));
  and2  gate1053(.a(G1192), .b(G21), .O(gate459inter2));
  inv1  gate1054(.a(s_72), .O(gate459inter3));
  inv1  gate1055(.a(s_73), .O(gate459inter4));
  nand2 gate1056(.a(gate459inter4), .b(gate459inter3), .O(gate459inter5));
  nor2  gate1057(.a(gate459inter5), .b(gate459inter2), .O(gate459inter6));
  inv1  gate1058(.a(G21), .O(gate459inter7));
  inv1  gate1059(.a(G1192), .O(gate459inter8));
  nand2 gate1060(.a(gate459inter8), .b(gate459inter7), .O(gate459inter9));
  nand2 gate1061(.a(s_73), .b(gate459inter3), .O(gate459inter10));
  nor2  gate1062(.a(gate459inter10), .b(gate459inter9), .O(gate459inter11));
  nor2  gate1063(.a(gate459inter11), .b(gate459inter6), .O(gate459inter12));
  nand2 gate1064(.a(gate459inter12), .b(gate459inter1), .O(G1268));
nand2 gate460( .a(G1096), .b(G1192), .O(G1269) );
nand2 gate461( .a(G22), .b(G1195), .O(G1270) );
nand2 gate462( .a(G1099), .b(G1195), .O(G1271) );
nand2 gate463( .a(G23), .b(G1198), .O(G1272) );
nand2 gate464( .a(G1102), .b(G1198), .O(G1273) );
nand2 gate465( .a(G24), .b(G1201), .O(G1274) );
nand2 gate466( .a(G1105), .b(G1201), .O(G1275) );
nand2 gate467( .a(G25), .b(G1204), .O(G1276) );
nand2 gate468( .a(G1108), .b(G1204), .O(G1277) );
nand2 gate469( .a(G26), .b(G1207), .O(G1278) );
nand2 gate470( .a(G1111), .b(G1207), .O(G1279) );
nand2 gate471( .a(G27), .b(G1210), .O(G1280) );
nand2 gate472( .a(G1114), .b(G1210), .O(G1281) );
nand2 gate473( .a(G28), .b(G1213), .O(G1282) );
nand2 gate474( .a(G1117), .b(G1213), .O(G1283) );
nand2 gate475( .a(G29), .b(G1216), .O(G1284) );
nand2 gate476( .a(G1120), .b(G1216), .O(G1285) );
nand2 gate477( .a(G30), .b(G1219), .O(G1286) );
nand2 gate478( .a(G1123), .b(G1219), .O(G1287) );
nand2 gate479( .a(G31), .b(G1222), .O(G1288) );
nand2 gate480( .a(G1126), .b(G1222), .O(G1289) );
nand2 gate481( .a(G32), .b(G1225), .O(G1290) );
nand2 gate482( .a(G1129), .b(G1225), .O(G1291) );
nand2 gate483( .a(G1228), .b(G1229), .O(G1292) );
nand2 gate484( .a(G1230), .b(G1231), .O(G1293) );
nand2 gate485( .a(G1232), .b(G1233), .O(G1294) );
nand2 gate486( .a(G1234), .b(G1235), .O(G1295) );
nand2 gate487( .a(G1236), .b(G1237), .O(G1296) );
nand2 gate488( .a(G1238), .b(G1239), .O(G1297) );
nand2 gate489( .a(G1240), .b(G1241), .O(G1298) );
nand2 gate490( .a(G1242), .b(G1243), .O(G1299) );

  xor2  gate1191(.a(G1245), .b(G1244), .O(gate491inter0));
  nand2 gate1192(.a(gate491inter0), .b(s_92), .O(gate491inter1));
  and2  gate1193(.a(G1245), .b(G1244), .O(gate491inter2));
  inv1  gate1194(.a(s_92), .O(gate491inter3));
  inv1  gate1195(.a(s_93), .O(gate491inter4));
  nand2 gate1196(.a(gate491inter4), .b(gate491inter3), .O(gate491inter5));
  nor2  gate1197(.a(gate491inter5), .b(gate491inter2), .O(gate491inter6));
  inv1  gate1198(.a(G1244), .O(gate491inter7));
  inv1  gate1199(.a(G1245), .O(gate491inter8));
  nand2 gate1200(.a(gate491inter8), .b(gate491inter7), .O(gate491inter9));
  nand2 gate1201(.a(s_93), .b(gate491inter3), .O(gate491inter10));
  nor2  gate1202(.a(gate491inter10), .b(gate491inter9), .O(gate491inter11));
  nor2  gate1203(.a(gate491inter11), .b(gate491inter6), .O(gate491inter12));
  nand2 gate1204(.a(gate491inter12), .b(gate491inter1), .O(G1300));
nand2 gate492( .a(G1246), .b(G1247), .O(G1301) );
nand2 gate493( .a(G1248), .b(G1249), .O(G1302) );
nand2 gate494( .a(G1250), .b(G1251), .O(G1303) );
nand2 gate495( .a(G1252), .b(G1253), .O(G1304) );
nand2 gate496( .a(G1254), .b(G1255), .O(G1305) );
nand2 gate497( .a(G1256), .b(G1257), .O(G1306) );
nand2 gate498( .a(G1258), .b(G1259), .O(G1307) );
nand2 gate499( .a(G1260), .b(G1261), .O(G1308) );
nand2 gate500( .a(G1262), .b(G1263), .O(G1309) );

  xor2  gate995(.a(G1265), .b(G1264), .O(gate501inter0));
  nand2 gate996(.a(gate501inter0), .b(s_64), .O(gate501inter1));
  and2  gate997(.a(G1265), .b(G1264), .O(gate501inter2));
  inv1  gate998(.a(s_64), .O(gate501inter3));
  inv1  gate999(.a(s_65), .O(gate501inter4));
  nand2 gate1000(.a(gate501inter4), .b(gate501inter3), .O(gate501inter5));
  nor2  gate1001(.a(gate501inter5), .b(gate501inter2), .O(gate501inter6));
  inv1  gate1002(.a(G1264), .O(gate501inter7));
  inv1  gate1003(.a(G1265), .O(gate501inter8));
  nand2 gate1004(.a(gate501inter8), .b(gate501inter7), .O(gate501inter9));
  nand2 gate1005(.a(s_65), .b(gate501inter3), .O(gate501inter10));
  nor2  gate1006(.a(gate501inter10), .b(gate501inter9), .O(gate501inter11));
  nor2  gate1007(.a(gate501inter11), .b(gate501inter6), .O(gate501inter12));
  nand2 gate1008(.a(gate501inter12), .b(gate501inter1), .O(G1310));
nand2 gate502( .a(G1266), .b(G1267), .O(G1311) );

  xor2  gate1387(.a(G1269), .b(G1268), .O(gate503inter0));
  nand2 gate1388(.a(gate503inter0), .b(s_120), .O(gate503inter1));
  and2  gate1389(.a(G1269), .b(G1268), .O(gate503inter2));
  inv1  gate1390(.a(s_120), .O(gate503inter3));
  inv1  gate1391(.a(s_121), .O(gate503inter4));
  nand2 gate1392(.a(gate503inter4), .b(gate503inter3), .O(gate503inter5));
  nor2  gate1393(.a(gate503inter5), .b(gate503inter2), .O(gate503inter6));
  inv1  gate1394(.a(G1268), .O(gate503inter7));
  inv1  gate1395(.a(G1269), .O(gate503inter8));
  nand2 gate1396(.a(gate503inter8), .b(gate503inter7), .O(gate503inter9));
  nand2 gate1397(.a(s_121), .b(gate503inter3), .O(gate503inter10));
  nor2  gate1398(.a(gate503inter10), .b(gate503inter9), .O(gate503inter11));
  nor2  gate1399(.a(gate503inter11), .b(gate503inter6), .O(gate503inter12));
  nand2 gate1400(.a(gate503inter12), .b(gate503inter1), .O(G1312));
nand2 gate504( .a(G1270), .b(G1271), .O(G1313) );
nand2 gate505( .a(G1272), .b(G1273), .O(G1314) );
nand2 gate506( .a(G1274), .b(G1275), .O(G1315) );
nand2 gate507( .a(G1276), .b(G1277), .O(G1316) );

  xor2  gate1303(.a(G1279), .b(G1278), .O(gate508inter0));
  nand2 gate1304(.a(gate508inter0), .b(s_108), .O(gate508inter1));
  and2  gate1305(.a(G1279), .b(G1278), .O(gate508inter2));
  inv1  gate1306(.a(s_108), .O(gate508inter3));
  inv1  gate1307(.a(s_109), .O(gate508inter4));
  nand2 gate1308(.a(gate508inter4), .b(gate508inter3), .O(gate508inter5));
  nor2  gate1309(.a(gate508inter5), .b(gate508inter2), .O(gate508inter6));
  inv1  gate1310(.a(G1278), .O(gate508inter7));
  inv1  gate1311(.a(G1279), .O(gate508inter8));
  nand2 gate1312(.a(gate508inter8), .b(gate508inter7), .O(gate508inter9));
  nand2 gate1313(.a(s_109), .b(gate508inter3), .O(gate508inter10));
  nor2  gate1314(.a(gate508inter10), .b(gate508inter9), .O(gate508inter11));
  nor2  gate1315(.a(gate508inter11), .b(gate508inter6), .O(gate508inter12));
  nand2 gate1316(.a(gate508inter12), .b(gate508inter1), .O(G1317));
nand2 gate509( .a(G1280), .b(G1281), .O(G1318) );
nand2 gate510( .a(G1282), .b(G1283), .O(G1319) );
nand2 gate511( .a(G1284), .b(G1285), .O(G1320) );

  xor2  gate939(.a(G1287), .b(G1286), .O(gate512inter0));
  nand2 gate940(.a(gate512inter0), .b(s_56), .O(gate512inter1));
  and2  gate941(.a(G1287), .b(G1286), .O(gate512inter2));
  inv1  gate942(.a(s_56), .O(gate512inter3));
  inv1  gate943(.a(s_57), .O(gate512inter4));
  nand2 gate944(.a(gate512inter4), .b(gate512inter3), .O(gate512inter5));
  nor2  gate945(.a(gate512inter5), .b(gate512inter2), .O(gate512inter6));
  inv1  gate946(.a(G1286), .O(gate512inter7));
  inv1  gate947(.a(G1287), .O(gate512inter8));
  nand2 gate948(.a(gate512inter8), .b(gate512inter7), .O(gate512inter9));
  nand2 gate949(.a(s_57), .b(gate512inter3), .O(gate512inter10));
  nor2  gate950(.a(gate512inter10), .b(gate512inter9), .O(gate512inter11));
  nor2  gate951(.a(gate512inter11), .b(gate512inter6), .O(gate512inter12));
  nand2 gate952(.a(gate512inter12), .b(gate512inter1), .O(G1321));
nand2 gate513( .a(G1288), .b(G1289), .O(G1322) );
nand2 gate514( .a(G1290), .b(G1291), .O(G1323) );
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule