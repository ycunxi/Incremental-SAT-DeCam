module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);

input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;//RE__PI;

input s_0,s_1;//RE__ALLOW(00,01,10,11);
input s_2,s_3;//RE__ALLOW(00,01,10,11);
input s_4,s_5;//RE__ALLOW(00,01,10,11);
input s_6,s_7;//RE__ALLOW(00,01,10,11);
input s_8,s_9;//RE__ALLOW(00,01,10,11);
input s_10,s_11;//RE__ALLOW(00,01,10,11);
input s_12,s_13;//RE__ALLOW(00,01,10,11);
input s_14,s_15;//RE__ALLOW(00,01,10,11);
input s_16,s_17;//RE__ALLOW(00,01,10,11);
input s_18,s_19;//RE__ALLOW(00,01,10,11);
input s_20,s_21;//RE__ALLOW(00,01,10,11);
input s_22,s_23;//RE__ALLOW(00,01,10,11);
input s_24,s_25;//RE__ALLOW(00,01,10,11);
input s_26,s_27;//RE__ALLOW(00,01,10,11);
input s_28,s_29;//RE__ALLOW(00,01,10,11);
input s_30,s_31;//RE__ALLOW(00,01,10,11);
input s_32,s_33;//RE__ALLOW(00,01,10,11);
input s_34,s_35;//RE__ALLOW(00,01,10,11);
input s_36,s_37;//RE__ALLOW(00,01,10,11);
input s_38,s_39;//RE__ALLOW(00,01,10,11);
input s_40,s_41;//RE__ALLOW(00,01,10,11);
input s_42,s_43;//RE__ALLOW(00,01,10,11);
input s_44,s_45;//RE__ALLOW(00,01,10,11);
input s_46,s_47;//RE__ALLOW(00,01,10,11);
input s_48,s_49;//RE__ALLOW(00,01,10,11);
input s_50,s_51;//RE__ALLOW(00,01,10,11);
input s_52,s_53;//RE__ALLOW(00,01,10,11);
input s_54,s_55;//RE__ALLOW(00,01,10,11);
input s_56,s_57;//RE__ALLOW(00,01,10,11);
input s_58,s_59;//RE__ALLOW(00,01,10,11);
input s_60,s_61;//RE__ALLOW(00,01,10,11);
input s_62,s_63;//RE__ALLOW(00,01,10,11);
input s_64,s_65;//RE__ALLOW(00,01,10,11);
input s_66,s_67;//RE__ALLOW(00,01,10,11);
input s_68,s_69;//RE__ALLOW(00,01,10,11);
input s_70,s_71;//RE__ALLOW(00,01,10,11);
input s_72,s_73;//RE__ALLOW(00,01,10,11);
input s_74,s_75;//RE__ALLOW(00,01,10,11);
input s_76,s_77;//RE__ALLOW(00,01,10,11);
input s_78,s_79;//RE__ALLOW(00,01,10,11);
input s_80,s_81;//RE__ALLOW(00,01,10,11);
input s_82,s_83;//RE__ALLOW(00,01,10,11);
input s_84,s_85;//RE__ALLOW(00,01,10,11);
input s_86,s_87;//RE__ALLOW(00,01,10,11);
input s_88,s_89;//RE__ALLOW(00,01,10,11);
input s_90,s_91;//RE__ALLOW(00,01,10,11);
input s_92,s_93;//RE__ALLOW(00,01,10,11);
input s_94,s_95;//RE__ALLOW(00,01,10,11);
input s_96,s_97;//RE__ALLOW(00,01,10,11);
input s_98,s_99;//RE__ALLOW(00,01,10,11);
input s_100,s_101;//RE__ALLOW(00,01,10,11);
input s_102,s_103;//RE__ALLOW(00,01,10,11);
input s_104,s_105;//RE__ALLOW(00,01,10,11);
input s_106,s_107;//RE__ALLOW(00,01,10,11);
input s_108,s_109;//RE__ALLOW(00,01,10,11);
input s_110,s_111;//RE__ALLOW(00,01,10,11);
input s_112,s_113;//RE__ALLOW(00,01,10,11);
input s_114,s_115;//RE__ALLOW(00,01,10,11);
input s_116,s_117;//RE__ALLOW(00,01,10,11);
input s_118,s_119;//RE__ALLOW(00,01,10,11);
input s_120,s_121;//RE__ALLOW(00,01,10,11);
input s_122,s_123;//RE__ALLOW(00,01,10,11);
input s_124,s_125;//RE__ALLOW(00,01,10,11);
input s_126,s_127;//RE__ALLOW(00,01,10,11);
input s_128,s_129;//RE__ALLOW(00,01,10,11);
input s_130,s_131;//RE__ALLOW(00,01,10,11);
input s_132,s_133;//RE__ALLOW(00,01,10,11);
input s_134,s_135;//RE__ALLOW(00,01,10,11);
input s_136,s_137;//RE__ALLOW(00,01,10,11);
input s_138,s_139;//RE__ALLOW(00,01,10,11);
input s_140,s_141;//RE__ALLOW(00,01,10,11);
input s_142,s_143;//RE__ALLOW(00,01,10,11);
input s_144,s_145;//RE__ALLOW(00,01,10,11);
input s_146,s_147;//RE__ALLOW(00,01,10,11);
input s_148,s_149;//RE__ALLOW(00,01,10,11);
input s_150,s_151;//RE__ALLOW(00,01,10,11);
input s_152,s_153;//RE__ALLOW(00,01,10,11);
input s_154,s_155;//RE__ALLOW(00,01,10,11);
input s_156,s_157;//RE__ALLOW(00,01,10,11);
input s_158,s_159;//RE__ALLOW(00,01,10,11);
input s_160,s_161;//RE__ALLOW(00,01,10,11);
input s_162,s_163;//RE__ALLOW(00,01,10,11);
input s_164,s_165;//RE__ALLOW(00,01,10,11);
input s_166,s_167;//RE__ALLOW(00,01,10,11);
input s_168,s_169;//RE__ALLOW(00,01,10,11);
input s_170,s_171;//RE__ALLOW(00,01,10,11);
input s_172,s_173;//RE__ALLOW(00,01,10,11);
input s_174,s_175;//RE__ALLOW(00,01,10,11);
input s_176,s_177;//RE__ALLOW(00,01,10,11);
input s_178,s_179;//RE__ALLOW(00,01,10,11);
input s_180,s_181;//RE__ALLOW(00,01,10,11);
input s_182,s_183;//RE__ALLOW(00,01,10,11);
input s_184,s_185;//RE__ALLOW(00,01,10,11);
input s_186,s_187;//RE__ALLOW(00,01,10,11);
input s_188,s_189;//RE__ALLOW(00,01,10,11);
input s_190,s_191;//RE__ALLOW(00,01,10,11);
input s_192,s_193;//RE__ALLOW(00,01,10,11);
input s_194,s_195;//RE__ALLOW(00,01,10,11);
input s_196,s_197;//RE__ALLOW(00,01,10,11);
input s_198,s_199;//RE__ALLOW(00,01,10,11);
input s_200,s_201;//RE__ALLOW(00,01,10,11);
input s_202,s_203;//RE__ALLOW(00,01,10,11);
input s_204,s_205;//RE__ALLOW(00,01,10,11);
input s_206,s_207;//RE__ALLOW(00,01,10,11);
input s_208,s_209;//RE__ALLOW(00,01,10,11);
input s_210,s_211;//RE__ALLOW(00,01,10,11);
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;

  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate513inter0, gate513inter1, gate513inter2, gate513inter3, gate513inter4, gate513inter5, gate513inter6, gate513inter7, gate513inter8, gate513inter9, gate513inter10, gate513inter11, gate513inter12, gate204inter0, gate204inter1, gate204inter2, gate204inter3, gate204inter4, gate204inter5, gate204inter6, gate204inter7, gate204inter8, gate204inter9, gate204inter10, gate204inter11, gate204inter12, gate100inter0, gate100inter1, gate100inter2, gate100inter3, gate100inter4, gate100inter5, gate100inter6, gate100inter7, gate100inter8, gate100inter9, gate100inter10, gate100inter11, gate100inter12, gate82inter0, gate82inter1, gate82inter2, gate82inter3, gate82inter4, gate82inter5, gate82inter6, gate82inter7, gate82inter8, gate82inter9, gate82inter10, gate82inter11, gate82inter12, gate76inter0, gate76inter1, gate76inter2, gate76inter3, gate76inter4, gate76inter5, gate76inter6, gate76inter7, gate76inter8, gate76inter9, gate76inter10, gate76inter11, gate76inter12, gate289inter0, gate289inter1, gate289inter2, gate289inter3, gate289inter4, gate289inter5, gate289inter6, gate289inter7, gate289inter8, gate289inter9, gate289inter10, gate289inter11, gate289inter12, gate86inter0, gate86inter1, gate86inter2, gate86inter3, gate86inter4, gate86inter5, gate86inter6, gate86inter7, gate86inter8, gate86inter9, gate86inter10, gate86inter11, gate86inter12, gate290inter0, gate290inter1, gate290inter2, gate290inter3, gate290inter4, gate290inter5, gate290inter6, gate290inter7, gate290inter8, gate290inter9, gate290inter10, gate290inter11, gate290inter12, gate401inter0, gate401inter1, gate401inter2, gate401inter3, gate401inter4, gate401inter5, gate401inter6, gate401inter7, gate401inter8, gate401inter9, gate401inter10, gate401inter11, gate401inter12, gate55inter0, gate55inter1, gate55inter2, gate55inter3, gate55inter4, gate55inter5, gate55inter6, gate55inter7, gate55inter8, gate55inter9, gate55inter10, gate55inter11, gate55inter12, gate123inter0, gate123inter1, gate123inter2, gate123inter3, gate123inter4, gate123inter5, gate123inter6, gate123inter7, gate123inter8, gate123inter9, gate123inter10, gate123inter11, gate123inter12, gate33inter0, gate33inter1, gate33inter2, gate33inter3, gate33inter4, gate33inter5, gate33inter6, gate33inter7, gate33inter8, gate33inter9, gate33inter10, gate33inter11, gate33inter12, gate262inter0, gate262inter1, gate262inter2, gate262inter3, gate262inter4, gate262inter5, gate262inter6, gate262inter7, gate262inter8, gate262inter9, gate262inter10, gate262inter11, gate262inter12, gate281inter0, gate281inter1, gate281inter2, gate281inter3, gate281inter4, gate281inter5, gate281inter6, gate281inter7, gate281inter8, gate281inter9, gate281inter10, gate281inter11, gate281inter12, gate469inter0, gate469inter1, gate469inter2, gate469inter3, gate469inter4, gate469inter5, gate469inter6, gate469inter7, gate469inter8, gate469inter9, gate469inter10, gate469inter11, gate469inter12, gate398inter0, gate398inter1, gate398inter2, gate398inter3, gate398inter4, gate398inter5, gate398inter6, gate398inter7, gate398inter8, gate398inter9, gate398inter10, gate398inter11, gate398inter12, gate28inter0, gate28inter1, gate28inter2, gate28inter3, gate28inter4, gate28inter5, gate28inter6, gate28inter7, gate28inter8, gate28inter9, gate28inter10, gate28inter11, gate28inter12, gate287inter0, gate287inter1, gate287inter2, gate287inter3, gate287inter4, gate287inter5, gate287inter6, gate287inter7, gate287inter8, gate287inter9, gate287inter10, gate287inter11, gate287inter12, gate80inter0, gate80inter1, gate80inter2, gate80inter3, gate80inter4, gate80inter5, gate80inter6, gate80inter7, gate80inter8, gate80inter9, gate80inter10, gate80inter11, gate80inter12, gate68inter0, gate68inter1, gate68inter2, gate68inter3, gate68inter4, gate68inter5, gate68inter6, gate68inter7, gate68inter8, gate68inter9, gate68inter10, gate68inter11, gate68inter12, gate498inter0, gate498inter1, gate498inter2, gate498inter3, gate498inter4, gate498inter5, gate498inter6, gate498inter7, gate498inter8, gate498inter9, gate498inter10, gate498inter11, gate498inter12, gate505inter0, gate505inter1, gate505inter2, gate505inter3, gate505inter4, gate505inter5, gate505inter6, gate505inter7, gate505inter8, gate505inter9, gate505inter10, gate505inter11, gate505inter12, gate128inter0, gate128inter1, gate128inter2, gate128inter3, gate128inter4, gate128inter5, gate128inter6, gate128inter7, gate128inter8, gate128inter9, gate128inter10, gate128inter11, gate128inter12, gate152inter0, gate152inter1, gate152inter2, gate152inter3, gate152inter4, gate152inter5, gate152inter6, gate152inter7, gate152inter8, gate152inter9, gate152inter10, gate152inter11, gate152inter12, gate22inter0, gate22inter1, gate22inter2, gate22inter3, gate22inter4, gate22inter5, gate22inter6, gate22inter7, gate22inter8, gate22inter9, gate22inter10, gate22inter11, gate22inter12, gate488inter0, gate488inter1, gate488inter2, gate488inter3, gate488inter4, gate488inter5, gate488inter6, gate488inter7, gate488inter8, gate488inter9, gate488inter10, gate488inter11, gate488inter12, gate176inter0, gate176inter1, gate176inter2, gate176inter3, gate176inter4, gate176inter5, gate176inter6, gate176inter7, gate176inter8, gate176inter9, gate176inter10, gate176inter11, gate176inter12, gate37inter0, gate37inter1, gate37inter2, gate37inter3, gate37inter4, gate37inter5, gate37inter6, gate37inter7, gate37inter8, gate37inter9, gate37inter10, gate37inter11, gate37inter12, gate233inter0, gate233inter1, gate233inter2, gate233inter3, gate233inter4, gate233inter5, gate233inter6, gate233inter7, gate233inter8, gate233inter9, gate233inter10, gate233inter11, gate233inter12, gate444inter0, gate444inter1, gate444inter2, gate444inter3, gate444inter4, gate444inter5, gate444inter6, gate444inter7, gate444inter8, gate444inter9, gate444inter10, gate444inter11, gate444inter12, gate507inter0, gate507inter1, gate507inter2, gate507inter3, gate507inter4, gate507inter5, gate507inter6, gate507inter7, gate507inter8, gate507inter9, gate507inter10, gate507inter11, gate507inter12, gate158inter0, gate158inter1, gate158inter2, gate158inter3, gate158inter4, gate158inter5, gate158inter6, gate158inter7, gate158inter8, gate158inter9, gate158inter10, gate158inter11, gate158inter12, gate195inter0, gate195inter1, gate195inter2, gate195inter3, gate195inter4, gate195inter5, gate195inter6, gate195inter7, gate195inter8, gate195inter9, gate195inter10, gate195inter11, gate195inter12, gate451inter0, gate451inter1, gate451inter2, gate451inter3, gate451inter4, gate451inter5, gate451inter6, gate451inter7, gate451inter8, gate451inter9, gate451inter10, gate451inter11, gate451inter12, gate34inter0, gate34inter1, gate34inter2, gate34inter3, gate34inter4, gate34inter5, gate34inter6, gate34inter7, gate34inter8, gate34inter9, gate34inter10, gate34inter11, gate34inter12, gate166inter0, gate166inter1, gate166inter2, gate166inter3, gate166inter4, gate166inter5, gate166inter6, gate166inter7, gate166inter8, gate166inter9, gate166inter10, gate166inter11, gate166inter12, gate452inter0, gate452inter1, gate452inter2, gate452inter3, gate452inter4, gate452inter5, gate452inter6, gate452inter7, gate452inter8, gate452inter9, gate452inter10, gate452inter11, gate452inter12, gate118inter0, gate118inter1, gate118inter2, gate118inter3, gate118inter4, gate118inter5, gate118inter6, gate118inter7, gate118inter8, gate118inter9, gate118inter10, gate118inter11, gate118inter12, gate127inter0, gate127inter1, gate127inter2, gate127inter3, gate127inter4, gate127inter5, gate127inter6, gate127inter7, gate127inter8, gate127inter9, gate127inter10, gate127inter11, gate127inter12, gate391inter0, gate391inter1, gate391inter2, gate391inter3, gate391inter4, gate391inter5, gate391inter6, gate391inter7, gate391inter8, gate391inter9, gate391inter10, gate391inter11, gate391inter12, gate285inter0, gate285inter1, gate285inter2, gate285inter3, gate285inter4, gate285inter5, gate285inter6, gate285inter7, gate285inter8, gate285inter9, gate285inter10, gate285inter11, gate285inter12, gate436inter0, gate436inter1, gate436inter2, gate436inter3, gate436inter4, gate436inter5, gate436inter6, gate436inter7, gate436inter8, gate436inter9, gate436inter10, gate436inter11, gate436inter12, gate144inter0, gate144inter1, gate144inter2, gate144inter3, gate144inter4, gate144inter5, gate144inter6, gate144inter7, gate144inter8, gate144inter9, gate144inter10, gate144inter11, gate144inter12, gate23inter0, gate23inter1, gate23inter2, gate23inter3, gate23inter4, gate23inter5, gate23inter6, gate23inter7, gate23inter8, gate23inter9, gate23inter10, gate23inter11, gate23inter12, gate491inter0, gate491inter1, gate491inter2, gate491inter3, gate491inter4, gate491inter5, gate491inter6, gate491inter7, gate491inter8, gate491inter9, gate491inter10, gate491inter11, gate491inter12, gate225inter0, gate225inter1, gate225inter2, gate225inter3, gate225inter4, gate225inter5, gate225inter6, gate225inter7, gate225inter8, gate225inter9, gate225inter10, gate225inter11, gate225inter12, gate163inter0, gate163inter1, gate163inter2, gate163inter3, gate163inter4, gate163inter5, gate163inter6, gate163inter7, gate163inter8, gate163inter9, gate163inter10, gate163inter11, gate163inter12, gate410inter0, gate410inter1, gate410inter2, gate410inter3, gate410inter4, gate410inter5, gate410inter6, gate410inter7, gate410inter8, gate410inter9, gate410inter10, gate410inter11, gate410inter12, gate492inter0, gate492inter1, gate492inter2, gate492inter3, gate492inter4, gate492inter5, gate492inter6, gate492inter7, gate492inter8, gate492inter9, gate492inter10, gate492inter11, gate492inter12, gate227inter0, gate227inter1, gate227inter2, gate227inter3, gate227inter4, gate227inter5, gate227inter6, gate227inter7, gate227inter8, gate227inter9, gate227inter10, gate227inter11, gate227inter12, gate61inter0, gate61inter1, gate61inter2, gate61inter3, gate61inter4, gate61inter5, gate61inter6, gate61inter7, gate61inter8, gate61inter9, gate61inter10, gate61inter11, gate61inter12, gate63inter0, gate63inter1, gate63inter2, gate63inter3, gate63inter4, gate63inter5, gate63inter6, gate63inter7, gate63inter8, gate63inter9, gate63inter10, gate63inter11, gate63inter12, gate243inter0, gate243inter1, gate243inter2, gate243inter3, gate243inter4, gate243inter5, gate243inter6, gate243inter7, gate243inter8, gate243inter9, gate243inter10, gate243inter11, gate243inter12, gate266inter0, gate266inter1, gate266inter2, gate266inter3, gate266inter4, gate266inter5, gate266inter6, gate266inter7, gate266inter8, gate266inter9, gate266inter10, gate266inter11, gate266inter12, gate89inter0, gate89inter1, gate89inter2, gate89inter3, gate89inter4, gate89inter5, gate89inter6, gate89inter7, gate89inter8, gate89inter9, gate89inter10, gate89inter11, gate89inter12, gate280inter0, gate280inter1, gate280inter2, gate280inter3, gate280inter4, gate280inter5, gate280inter6, gate280inter7, gate280inter8, gate280inter9, gate280inter10, gate280inter11, gate280inter12, gate210inter0, gate210inter1, gate210inter2, gate210inter3, gate210inter4, gate210inter5, gate210inter6, gate210inter7, gate210inter8, gate210inter9, gate210inter10, gate210inter11, gate210inter12, gate60inter0, gate60inter1, gate60inter2, gate60inter3, gate60inter4, gate60inter5, gate60inter6, gate60inter7, gate60inter8, gate60inter9, gate60inter10, gate60inter11, gate60inter12, gate114inter0, gate114inter1, gate114inter2, gate114inter3, gate114inter4, gate114inter5, gate114inter6, gate114inter7, gate114inter8, gate114inter9, gate114inter10, gate114inter11, gate114inter12, gate194inter0, gate194inter1, gate194inter2, gate194inter3, gate194inter4, gate194inter5, gate194inter6, gate194inter7, gate194inter8, gate194inter9, gate194inter10, gate194inter11, gate194inter12, gate235inter0, gate235inter1, gate235inter2, gate235inter3, gate235inter4, gate235inter5, gate235inter6, gate235inter7, gate235inter8, gate235inter9, gate235inter10, gate235inter11, gate235inter12, gate18inter0, gate18inter1, gate18inter2, gate18inter3, gate18inter4, gate18inter5, gate18inter6, gate18inter7, gate18inter8, gate18inter9, gate18inter10, gate18inter11, gate18inter12, gate190inter0, gate190inter1, gate190inter2, gate190inter3, gate190inter4, gate190inter5, gate190inter6, gate190inter7, gate190inter8, gate190inter9, gate190inter10, gate190inter11, gate190inter12, gate71inter0, gate71inter1, gate71inter2, gate71inter3, gate71inter4, gate71inter5, gate71inter6, gate71inter7, gate71inter8, gate71inter9, gate71inter10, gate71inter11, gate71inter12, gate431inter0, gate431inter1, gate431inter2, gate431inter3, gate431inter4, gate431inter5, gate431inter6, gate431inter7, gate431inter8, gate431inter9, gate431inter10, gate431inter11, gate431inter12, gate508inter0, gate508inter1, gate508inter2, gate508inter3, gate508inter4, gate508inter5, gate508inter6, gate508inter7, gate508inter8, gate508inter9, gate508inter10, gate508inter11, gate508inter12, gate460inter0, gate460inter1, gate460inter2, gate460inter3, gate460inter4, gate460inter5, gate460inter6, gate460inter7, gate460inter8, gate460inter9, gate460inter10, gate460inter11, gate460inter12, gate222inter0, gate222inter1, gate222inter2, gate222inter3, gate222inter4, gate222inter5, gate222inter6, gate222inter7, gate222inter8, gate222inter9, gate222inter10, gate222inter11, gate222inter12, gate138inter0, gate138inter1, gate138inter2, gate138inter3, gate138inter4, gate138inter5, gate138inter6, gate138inter7, gate138inter8, gate138inter9, gate138inter10, gate138inter11, gate138inter12, gate145inter0, gate145inter1, gate145inter2, gate145inter3, gate145inter4, gate145inter5, gate145inter6, gate145inter7, gate145inter8, gate145inter9, gate145inter10, gate145inter11, gate145inter12, gate107inter0, gate107inter1, gate107inter2, gate107inter3, gate107inter4, gate107inter5, gate107inter6, gate107inter7, gate107inter8, gate107inter9, gate107inter10, gate107inter11, gate107inter12, gate171inter0, gate171inter1, gate171inter2, gate171inter3, gate171inter4, gate171inter5, gate171inter6, gate171inter7, gate171inter8, gate171inter9, gate171inter10, gate171inter11, gate171inter12, gate263inter0, gate263inter1, gate263inter2, gate263inter3, gate263inter4, gate263inter5, gate263inter6, gate263inter7, gate263inter8, gate263inter9, gate263inter10, gate263inter11, gate263inter12, gate155inter0, gate155inter1, gate155inter2, gate155inter3, gate155inter4, gate155inter5, gate155inter6, gate155inter7, gate155inter8, gate155inter9, gate155inter10, gate155inter11, gate155inter12, gate173inter0, gate173inter1, gate173inter2, gate173inter3, gate173inter4, gate173inter5, gate173inter6, gate173inter7, gate173inter8, gate173inter9, gate173inter10, gate173inter11, gate173inter12, gate474inter0, gate474inter1, gate474inter2, gate474inter3, gate474inter4, gate474inter5, gate474inter6, gate474inter7, gate474inter8, gate474inter9, gate474inter10, gate474inter11, gate474inter12, gate75inter0, gate75inter1, gate75inter2, gate75inter3, gate75inter4, gate75inter5, gate75inter6, gate75inter7, gate75inter8, gate75inter9, gate75inter10, gate75inter11, gate75inter12, gate84inter0, gate84inter1, gate84inter2, gate84inter3, gate84inter4, gate84inter5, gate84inter6, gate84inter7, gate84inter8, gate84inter9, gate84inter10, gate84inter11, gate84inter12, gate504inter0, gate504inter1, gate504inter2, gate504inter3, gate504inter4, gate504inter5, gate504inter6, gate504inter7, gate504inter8, gate504inter9, gate504inter10, gate504inter11, gate504inter12, gate25inter0, gate25inter1, gate25inter2, gate25inter3, gate25inter4, gate25inter5, gate25inter6, gate25inter7, gate25inter8, gate25inter9, gate25inter10, gate25inter11, gate25inter12, gate132inter0, gate132inter1, gate132inter2, gate132inter3, gate132inter4, gate132inter5, gate132inter6, gate132inter7, gate132inter8, gate132inter9, gate132inter10, gate132inter11, gate132inter12, gate267inter0, gate267inter1, gate267inter2, gate267inter3, gate267inter4, gate267inter5, gate267inter6, gate267inter7, gate267inter8, gate267inter9, gate267inter10, gate267inter11, gate267inter12, gate30inter0, gate30inter1, gate30inter2, gate30inter3, gate30inter4, gate30inter5, gate30inter6, gate30inter7, gate30inter8, gate30inter9, gate30inter10, gate30inter11, gate30inter12, gate98inter0, gate98inter1, gate98inter2, gate98inter3, gate98inter4, gate98inter5, gate98inter6, gate98inter7, gate98inter8, gate98inter9, gate98inter10, gate98inter11, gate98inter12, gate205inter0, gate205inter1, gate205inter2, gate205inter3, gate205inter4, gate205inter5, gate205inter6, gate205inter7, gate205inter8, gate205inter9, gate205inter10, gate205inter11, gate205inter12, gate493inter0, gate493inter1, gate493inter2, gate493inter3, gate493inter4, gate493inter5, gate493inter6, gate493inter7, gate493inter8, gate493inter9, gate493inter10, gate493inter11, gate493inter12, gate150inter0, gate150inter1, gate150inter2, gate150inter3, gate150inter4, gate150inter5, gate150inter6, gate150inter7, gate150inter8, gate150inter9, gate150inter10, gate150inter11, gate150inter12, gate119inter0, gate119inter1, gate119inter2, gate119inter3, gate119inter4, gate119inter5, gate119inter6, gate119inter7, gate119inter8, gate119inter9, gate119inter10, gate119inter11, gate119inter12, gate39inter0, gate39inter1, gate39inter2, gate39inter3, gate39inter4, gate39inter5, gate39inter6, gate39inter7, gate39inter8, gate39inter9, gate39inter10, gate39inter11, gate39inter12, gate224inter0, gate224inter1, gate224inter2, gate224inter3, gate224inter4, gate224inter5, gate224inter6, gate224inter7, gate224inter8, gate224inter9, gate224inter10, gate224inter11, gate224inter12, gate111inter0, gate111inter1, gate111inter2, gate111inter3, gate111inter4, gate111inter5, gate111inter6, gate111inter7, gate111inter8, gate111inter9, gate111inter10, gate111inter11, gate111inter12, gate247inter0, gate247inter1, gate247inter2, gate247inter3, gate247inter4, gate247inter5, gate247inter6, gate247inter7, gate247inter8, gate247inter9, gate247inter10, gate247inter11, gate247inter12, gate16inter0, gate16inter1, gate16inter2, gate16inter3, gate16inter4, gate16inter5, gate16inter6, gate16inter7, gate16inter8, gate16inter9, gate16inter10, gate16inter11, gate16inter12, gate295inter0, gate295inter1, gate295inter2, gate295inter3, gate295inter4, gate295inter5, gate295inter6, gate295inter7, gate295inter8, gate295inter9, gate295inter10, gate295inter11, gate295inter12, gate46inter0, gate46inter1, gate46inter2, gate46inter3, gate46inter4, gate46inter5, gate46inter6, gate46inter7, gate46inter8, gate46inter9, gate46inter10, gate46inter11, gate46inter12, gate237inter0, gate237inter1, gate237inter2, gate237inter3, gate237inter4, gate237inter5, gate237inter6, gate237inter7, gate237inter8, gate237inter9, gate237inter10, gate237inter11, gate237inter12, gate477inter0, gate477inter1, gate477inter2, gate477inter3, gate477inter4, gate477inter5, gate477inter6, gate477inter7, gate477inter8, gate477inter9, gate477inter10, gate477inter11, gate477inter12, gate261inter0, gate261inter1, gate261inter2, gate261inter3, gate261inter4, gate261inter5, gate261inter6, gate261inter7, gate261inter8, gate261inter9, gate261inter10, gate261inter11, gate261inter12, gate167inter0, gate167inter1, gate167inter2, gate167inter3, gate167inter4, gate167inter5, gate167inter6, gate167inter7, gate167inter8, gate167inter9, gate167inter10, gate167inter11, gate167inter12, gate213inter0, gate213inter1, gate213inter2, gate213inter3, gate213inter4, gate213inter5, gate213inter6, gate213inter7, gate213inter8, gate213inter9, gate213inter10, gate213inter11, gate213inter12, gate430inter0, gate430inter1, gate430inter2, gate430inter3, gate430inter4, gate430inter5, gate430inter6, gate430inter7, gate430inter8, gate430inter9, gate430inter10, gate430inter11, gate430inter12, gate105inter0, gate105inter1, gate105inter2, gate105inter3, gate105inter4, gate105inter5, gate105inter6, gate105inter7, gate105inter8, gate105inter9, gate105inter10, gate105inter11, gate105inter12, gate284inter0, gate284inter1, gate284inter2, gate284inter3, gate284inter4, gate284inter5, gate284inter6, gate284inter7, gate284inter8, gate284inter9, gate284inter10, gate284inter11, gate284inter12, gate482inter0, gate482inter1, gate482inter2, gate482inter3, gate482inter4, gate482inter5, gate482inter6, gate482inter7, gate482inter8, gate482inter9, gate482inter10, gate482inter11, gate482inter12, gate294inter0, gate294inter1, gate294inter2, gate294inter3, gate294inter4, gate294inter5, gate294inter6, gate294inter7, gate294inter8, gate294inter9, gate294inter10, gate294inter11, gate294inter12, gate229inter0, gate229inter1, gate229inter2, gate229inter3, gate229inter4, gate229inter5, gate229inter6, gate229inter7, gate229inter8, gate229inter9, gate229inter10, gate229inter11, gate229inter12;



and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );
nand2 gate9( .a(G1), .b(G2), .O(G266) );
nand2 gate10( .a(G3), .b(G4), .O(G269) );
nand2 gate11( .a(G5), .b(G6), .O(G272) );
nand2 gate12( .a(G7), .b(G8), .O(G275) );
nand2 gate13( .a(G9), .b(G10), .O(G278) );
nand2 gate14( .a(G11), .b(G12), .O(G281) );
nand2 gate15( .a(G13), .b(G14), .O(G284) );

  xor2  gate1835(.a(G16), .b(G15), .O(gate16inter0));
  nand2 gate1836(.a(gate16inter0), .b(s_184), .O(gate16inter1));
  and2  gate1837(.a(G16), .b(G15), .O(gate16inter2));
  inv1  gate1838(.a(s_184), .O(gate16inter3));
  inv1  gate1839(.a(s_185), .O(gate16inter4));
  nand2 gate1840(.a(gate16inter4), .b(gate16inter3), .O(gate16inter5));
  nor2  gate1841(.a(gate16inter5), .b(gate16inter2), .O(gate16inter6));
  inv1  gate1842(.a(G15), .O(gate16inter7));
  inv1  gate1843(.a(G16), .O(gate16inter8));
  nand2 gate1844(.a(gate16inter8), .b(gate16inter7), .O(gate16inter9));
  nand2 gate1845(.a(s_185), .b(gate16inter3), .O(gate16inter10));
  nor2  gate1846(.a(gate16inter10), .b(gate16inter9), .O(gate16inter11));
  nor2  gate1847(.a(gate16inter11), .b(gate16inter6), .O(gate16inter12));
  nand2 gate1848(.a(gate16inter12), .b(gate16inter1), .O(G287));
nand2 gate17( .a(G17), .b(G18), .O(G290) );

  xor2  gate1401(.a(G20), .b(G19), .O(gate18inter0));
  nand2 gate1402(.a(gate18inter0), .b(s_122), .O(gate18inter1));
  and2  gate1403(.a(G20), .b(G19), .O(gate18inter2));
  inv1  gate1404(.a(s_122), .O(gate18inter3));
  inv1  gate1405(.a(s_123), .O(gate18inter4));
  nand2 gate1406(.a(gate18inter4), .b(gate18inter3), .O(gate18inter5));
  nor2  gate1407(.a(gate18inter5), .b(gate18inter2), .O(gate18inter6));
  inv1  gate1408(.a(G19), .O(gate18inter7));
  inv1  gate1409(.a(G20), .O(gate18inter8));
  nand2 gate1410(.a(gate18inter8), .b(gate18inter7), .O(gate18inter9));
  nand2 gate1411(.a(s_123), .b(gate18inter3), .O(gate18inter10));
  nor2  gate1412(.a(gate18inter10), .b(gate18inter9), .O(gate18inter11));
  nor2  gate1413(.a(gate18inter11), .b(gate18inter6), .O(gate18inter12));
  nand2 gate1414(.a(gate18inter12), .b(gate18inter1), .O(G293));
nand2 gate19( .a(G21), .b(G22), .O(G296) );
nand2 gate20( .a(G23), .b(G24), .O(G299) );
nand2 gate21( .a(G25), .b(G26), .O(G302) );

  xor2  gate883(.a(G28), .b(G27), .O(gate22inter0));
  nand2 gate884(.a(gate22inter0), .b(s_48), .O(gate22inter1));
  and2  gate885(.a(G28), .b(G27), .O(gate22inter2));
  inv1  gate886(.a(s_48), .O(gate22inter3));
  inv1  gate887(.a(s_49), .O(gate22inter4));
  nand2 gate888(.a(gate22inter4), .b(gate22inter3), .O(gate22inter5));
  nor2  gate889(.a(gate22inter5), .b(gate22inter2), .O(gate22inter6));
  inv1  gate890(.a(G27), .O(gate22inter7));
  inv1  gate891(.a(G28), .O(gate22inter8));
  nand2 gate892(.a(gate22inter8), .b(gate22inter7), .O(gate22inter9));
  nand2 gate893(.a(s_49), .b(gate22inter3), .O(gate22inter10));
  nor2  gate894(.a(gate22inter10), .b(gate22inter9), .O(gate22inter11));
  nor2  gate895(.a(gate22inter11), .b(gate22inter6), .O(gate22inter12));
  nand2 gate896(.a(gate22inter12), .b(gate22inter1), .O(G305));

  xor2  gate1149(.a(G30), .b(G29), .O(gate23inter0));
  nand2 gate1150(.a(gate23inter0), .b(s_86), .O(gate23inter1));
  and2  gate1151(.a(G30), .b(G29), .O(gate23inter2));
  inv1  gate1152(.a(s_86), .O(gate23inter3));
  inv1  gate1153(.a(s_87), .O(gate23inter4));
  nand2 gate1154(.a(gate23inter4), .b(gate23inter3), .O(gate23inter5));
  nor2  gate1155(.a(gate23inter5), .b(gate23inter2), .O(gate23inter6));
  inv1  gate1156(.a(G29), .O(gate23inter7));
  inv1  gate1157(.a(G30), .O(gate23inter8));
  nand2 gate1158(.a(gate23inter8), .b(gate23inter7), .O(gate23inter9));
  nand2 gate1159(.a(s_87), .b(gate23inter3), .O(gate23inter10));
  nor2  gate1160(.a(gate23inter10), .b(gate23inter9), .O(gate23inter11));
  nor2  gate1161(.a(gate23inter11), .b(gate23inter6), .O(gate23inter12));
  nand2 gate1162(.a(gate23inter12), .b(gate23inter1), .O(G308));
nand2 gate24( .a(G31), .b(G32), .O(G311) );

  xor2  gate1653(.a(G5), .b(G1), .O(gate25inter0));
  nand2 gate1654(.a(gate25inter0), .b(s_158), .O(gate25inter1));
  and2  gate1655(.a(G5), .b(G1), .O(gate25inter2));
  inv1  gate1656(.a(s_158), .O(gate25inter3));
  inv1  gate1657(.a(s_159), .O(gate25inter4));
  nand2 gate1658(.a(gate25inter4), .b(gate25inter3), .O(gate25inter5));
  nor2  gate1659(.a(gate25inter5), .b(gate25inter2), .O(gate25inter6));
  inv1  gate1660(.a(G1), .O(gate25inter7));
  inv1  gate1661(.a(G5), .O(gate25inter8));
  nand2 gate1662(.a(gate25inter8), .b(gate25inter7), .O(gate25inter9));
  nand2 gate1663(.a(s_159), .b(gate25inter3), .O(gate25inter10));
  nor2  gate1664(.a(gate25inter10), .b(gate25inter9), .O(gate25inter11));
  nor2  gate1665(.a(gate25inter11), .b(gate25inter6), .O(gate25inter12));
  nand2 gate1666(.a(gate25inter12), .b(gate25inter1), .O(G314));
nand2 gate26( .a(G9), .b(G13), .O(G317) );
nand2 gate27( .a(G2), .b(G6), .O(G320) );

  xor2  gate771(.a(G14), .b(G10), .O(gate28inter0));
  nand2 gate772(.a(gate28inter0), .b(s_32), .O(gate28inter1));
  and2  gate773(.a(G14), .b(G10), .O(gate28inter2));
  inv1  gate774(.a(s_32), .O(gate28inter3));
  inv1  gate775(.a(s_33), .O(gate28inter4));
  nand2 gate776(.a(gate28inter4), .b(gate28inter3), .O(gate28inter5));
  nor2  gate777(.a(gate28inter5), .b(gate28inter2), .O(gate28inter6));
  inv1  gate778(.a(G10), .O(gate28inter7));
  inv1  gate779(.a(G14), .O(gate28inter8));
  nand2 gate780(.a(gate28inter8), .b(gate28inter7), .O(gate28inter9));
  nand2 gate781(.a(s_33), .b(gate28inter3), .O(gate28inter10));
  nor2  gate782(.a(gate28inter10), .b(gate28inter9), .O(gate28inter11));
  nor2  gate783(.a(gate28inter11), .b(gate28inter6), .O(gate28inter12));
  nand2 gate784(.a(gate28inter12), .b(gate28inter1), .O(G323));
nand2 gate29( .a(G3), .b(G7), .O(G326) );

  xor2  gate1695(.a(G15), .b(G11), .O(gate30inter0));
  nand2 gate1696(.a(gate30inter0), .b(s_164), .O(gate30inter1));
  and2  gate1697(.a(G15), .b(G11), .O(gate30inter2));
  inv1  gate1698(.a(s_164), .O(gate30inter3));
  inv1  gate1699(.a(s_165), .O(gate30inter4));
  nand2 gate1700(.a(gate30inter4), .b(gate30inter3), .O(gate30inter5));
  nor2  gate1701(.a(gate30inter5), .b(gate30inter2), .O(gate30inter6));
  inv1  gate1702(.a(G11), .O(gate30inter7));
  inv1  gate1703(.a(G15), .O(gate30inter8));
  nand2 gate1704(.a(gate30inter8), .b(gate30inter7), .O(gate30inter9));
  nand2 gate1705(.a(s_165), .b(gate30inter3), .O(gate30inter10));
  nor2  gate1706(.a(gate30inter10), .b(gate30inter9), .O(gate30inter11));
  nor2  gate1707(.a(gate30inter11), .b(gate30inter6), .O(gate30inter12));
  nand2 gate1708(.a(gate30inter12), .b(gate30inter1), .O(G329));
nand2 gate31( .a(G4), .b(G8), .O(G332) );
nand2 gate32( .a(G12), .b(G16), .O(G335) );

  xor2  gate701(.a(G21), .b(G17), .O(gate33inter0));
  nand2 gate702(.a(gate33inter0), .b(s_22), .O(gate33inter1));
  and2  gate703(.a(G21), .b(G17), .O(gate33inter2));
  inv1  gate704(.a(s_22), .O(gate33inter3));
  inv1  gate705(.a(s_23), .O(gate33inter4));
  nand2 gate706(.a(gate33inter4), .b(gate33inter3), .O(gate33inter5));
  nor2  gate707(.a(gate33inter5), .b(gate33inter2), .O(gate33inter6));
  inv1  gate708(.a(G17), .O(gate33inter7));
  inv1  gate709(.a(G21), .O(gate33inter8));
  nand2 gate710(.a(gate33inter8), .b(gate33inter7), .O(gate33inter9));
  nand2 gate711(.a(s_23), .b(gate33inter3), .O(gate33inter10));
  nor2  gate712(.a(gate33inter10), .b(gate33inter9), .O(gate33inter11));
  nor2  gate713(.a(gate33inter11), .b(gate33inter6), .O(gate33inter12));
  nand2 gate714(.a(gate33inter12), .b(gate33inter1), .O(G338));

  xor2  gate1023(.a(G29), .b(G25), .O(gate34inter0));
  nand2 gate1024(.a(gate34inter0), .b(s_68), .O(gate34inter1));
  and2  gate1025(.a(G29), .b(G25), .O(gate34inter2));
  inv1  gate1026(.a(s_68), .O(gate34inter3));
  inv1  gate1027(.a(s_69), .O(gate34inter4));
  nand2 gate1028(.a(gate34inter4), .b(gate34inter3), .O(gate34inter5));
  nor2  gate1029(.a(gate34inter5), .b(gate34inter2), .O(gate34inter6));
  inv1  gate1030(.a(G25), .O(gate34inter7));
  inv1  gate1031(.a(G29), .O(gate34inter8));
  nand2 gate1032(.a(gate34inter8), .b(gate34inter7), .O(gate34inter9));
  nand2 gate1033(.a(s_69), .b(gate34inter3), .O(gate34inter10));
  nor2  gate1034(.a(gate34inter10), .b(gate34inter9), .O(gate34inter11));
  nor2  gate1035(.a(gate34inter11), .b(gate34inter6), .O(gate34inter12));
  nand2 gate1036(.a(gate34inter12), .b(gate34inter1), .O(G341));
nand2 gate35( .a(G18), .b(G22), .O(G344) );
nand2 gate36( .a(G26), .b(G30), .O(G347) );

  xor2  gate925(.a(G23), .b(G19), .O(gate37inter0));
  nand2 gate926(.a(gate37inter0), .b(s_54), .O(gate37inter1));
  and2  gate927(.a(G23), .b(G19), .O(gate37inter2));
  inv1  gate928(.a(s_54), .O(gate37inter3));
  inv1  gate929(.a(s_55), .O(gate37inter4));
  nand2 gate930(.a(gate37inter4), .b(gate37inter3), .O(gate37inter5));
  nor2  gate931(.a(gate37inter5), .b(gate37inter2), .O(gate37inter6));
  inv1  gate932(.a(G19), .O(gate37inter7));
  inv1  gate933(.a(G23), .O(gate37inter8));
  nand2 gate934(.a(gate37inter8), .b(gate37inter7), .O(gate37inter9));
  nand2 gate935(.a(s_55), .b(gate37inter3), .O(gate37inter10));
  nor2  gate936(.a(gate37inter10), .b(gate37inter9), .O(gate37inter11));
  nor2  gate937(.a(gate37inter11), .b(gate37inter6), .O(gate37inter12));
  nand2 gate938(.a(gate37inter12), .b(gate37inter1), .O(G350));
nand2 gate38( .a(G27), .b(G31), .O(G353) );

  xor2  gate1779(.a(G24), .b(G20), .O(gate39inter0));
  nand2 gate1780(.a(gate39inter0), .b(s_176), .O(gate39inter1));
  and2  gate1781(.a(G24), .b(G20), .O(gate39inter2));
  inv1  gate1782(.a(s_176), .O(gate39inter3));
  inv1  gate1783(.a(s_177), .O(gate39inter4));
  nand2 gate1784(.a(gate39inter4), .b(gate39inter3), .O(gate39inter5));
  nor2  gate1785(.a(gate39inter5), .b(gate39inter2), .O(gate39inter6));
  inv1  gate1786(.a(G20), .O(gate39inter7));
  inv1  gate1787(.a(G24), .O(gate39inter8));
  nand2 gate1788(.a(gate39inter8), .b(gate39inter7), .O(gate39inter9));
  nand2 gate1789(.a(s_177), .b(gate39inter3), .O(gate39inter10));
  nor2  gate1790(.a(gate39inter10), .b(gate39inter9), .O(gate39inter11));
  nor2  gate1791(.a(gate39inter11), .b(gate39inter6), .O(gate39inter12));
  nand2 gate1792(.a(gate39inter12), .b(gate39inter1), .O(G356));
nand2 gate40( .a(G28), .b(G32), .O(G359) );
nand2 gate41( .a(G1), .b(G266), .O(G362) );
nand2 gate42( .a(G2), .b(G266), .O(G363) );
nand2 gate43( .a(G3), .b(G269), .O(G364) );
nand2 gate44( .a(G4), .b(G269), .O(G365) );
nand2 gate45( .a(G5), .b(G272), .O(G366) );

  xor2  gate1863(.a(G272), .b(G6), .O(gate46inter0));
  nand2 gate1864(.a(gate46inter0), .b(s_188), .O(gate46inter1));
  and2  gate1865(.a(G272), .b(G6), .O(gate46inter2));
  inv1  gate1866(.a(s_188), .O(gate46inter3));
  inv1  gate1867(.a(s_189), .O(gate46inter4));
  nand2 gate1868(.a(gate46inter4), .b(gate46inter3), .O(gate46inter5));
  nor2  gate1869(.a(gate46inter5), .b(gate46inter2), .O(gate46inter6));
  inv1  gate1870(.a(G6), .O(gate46inter7));
  inv1  gate1871(.a(G272), .O(gate46inter8));
  nand2 gate1872(.a(gate46inter8), .b(gate46inter7), .O(gate46inter9));
  nand2 gate1873(.a(s_189), .b(gate46inter3), .O(gate46inter10));
  nor2  gate1874(.a(gate46inter10), .b(gate46inter9), .O(gate46inter11));
  nor2  gate1875(.a(gate46inter11), .b(gate46inter6), .O(gate46inter12));
  nand2 gate1876(.a(gate46inter12), .b(gate46inter1), .O(G367));
nand2 gate47( .a(G7), .b(G275), .O(G368) );
nand2 gate48( .a(G8), .b(G275), .O(G369) );
nand2 gate49( .a(G9), .b(G278), .O(G370) );
nand2 gate50( .a(G10), .b(G278), .O(G371) );
nand2 gate51( .a(G11), .b(G281), .O(G372) );
nand2 gate52( .a(G12), .b(G281), .O(G373) );
nand2 gate53( .a(G13), .b(G284), .O(G374) );
nand2 gate54( .a(G14), .b(G284), .O(G375) );

  xor2  gate673(.a(G287), .b(G15), .O(gate55inter0));
  nand2 gate674(.a(gate55inter0), .b(s_18), .O(gate55inter1));
  and2  gate675(.a(G287), .b(G15), .O(gate55inter2));
  inv1  gate676(.a(s_18), .O(gate55inter3));
  inv1  gate677(.a(s_19), .O(gate55inter4));
  nand2 gate678(.a(gate55inter4), .b(gate55inter3), .O(gate55inter5));
  nor2  gate679(.a(gate55inter5), .b(gate55inter2), .O(gate55inter6));
  inv1  gate680(.a(G15), .O(gate55inter7));
  inv1  gate681(.a(G287), .O(gate55inter8));
  nand2 gate682(.a(gate55inter8), .b(gate55inter7), .O(gate55inter9));
  nand2 gate683(.a(s_19), .b(gate55inter3), .O(gate55inter10));
  nor2  gate684(.a(gate55inter10), .b(gate55inter9), .O(gate55inter11));
  nor2  gate685(.a(gate55inter11), .b(gate55inter6), .O(gate55inter12));
  nand2 gate686(.a(gate55inter12), .b(gate55inter1), .O(G376));
nand2 gate56( .a(G16), .b(G287), .O(G377) );
nand2 gate57( .a(G17), .b(G290), .O(G378) );
nand2 gate58( .a(G18), .b(G290), .O(G379) );
nand2 gate59( .a(G19), .b(G293), .O(G380) );

  xor2  gate1345(.a(G293), .b(G20), .O(gate60inter0));
  nand2 gate1346(.a(gate60inter0), .b(s_114), .O(gate60inter1));
  and2  gate1347(.a(G293), .b(G20), .O(gate60inter2));
  inv1  gate1348(.a(s_114), .O(gate60inter3));
  inv1  gate1349(.a(s_115), .O(gate60inter4));
  nand2 gate1350(.a(gate60inter4), .b(gate60inter3), .O(gate60inter5));
  nor2  gate1351(.a(gate60inter5), .b(gate60inter2), .O(gate60inter6));
  inv1  gate1352(.a(G20), .O(gate60inter7));
  inv1  gate1353(.a(G293), .O(gate60inter8));
  nand2 gate1354(.a(gate60inter8), .b(gate60inter7), .O(gate60inter9));
  nand2 gate1355(.a(s_115), .b(gate60inter3), .O(gate60inter10));
  nor2  gate1356(.a(gate60inter10), .b(gate60inter9), .O(gate60inter11));
  nor2  gate1357(.a(gate60inter11), .b(gate60inter6), .O(gate60inter12));
  nand2 gate1358(.a(gate60inter12), .b(gate60inter1), .O(G381));

  xor2  gate1247(.a(G296), .b(G21), .O(gate61inter0));
  nand2 gate1248(.a(gate61inter0), .b(s_100), .O(gate61inter1));
  and2  gate1249(.a(G296), .b(G21), .O(gate61inter2));
  inv1  gate1250(.a(s_100), .O(gate61inter3));
  inv1  gate1251(.a(s_101), .O(gate61inter4));
  nand2 gate1252(.a(gate61inter4), .b(gate61inter3), .O(gate61inter5));
  nor2  gate1253(.a(gate61inter5), .b(gate61inter2), .O(gate61inter6));
  inv1  gate1254(.a(G21), .O(gate61inter7));
  inv1  gate1255(.a(G296), .O(gate61inter8));
  nand2 gate1256(.a(gate61inter8), .b(gate61inter7), .O(gate61inter9));
  nand2 gate1257(.a(s_101), .b(gate61inter3), .O(gate61inter10));
  nor2  gate1258(.a(gate61inter10), .b(gate61inter9), .O(gate61inter11));
  nor2  gate1259(.a(gate61inter11), .b(gate61inter6), .O(gate61inter12));
  nand2 gate1260(.a(gate61inter12), .b(gate61inter1), .O(G382));
nand2 gate62( .a(G22), .b(G296), .O(G383) );

  xor2  gate1261(.a(G299), .b(G23), .O(gate63inter0));
  nand2 gate1262(.a(gate63inter0), .b(s_102), .O(gate63inter1));
  and2  gate1263(.a(G299), .b(G23), .O(gate63inter2));
  inv1  gate1264(.a(s_102), .O(gate63inter3));
  inv1  gate1265(.a(s_103), .O(gate63inter4));
  nand2 gate1266(.a(gate63inter4), .b(gate63inter3), .O(gate63inter5));
  nor2  gate1267(.a(gate63inter5), .b(gate63inter2), .O(gate63inter6));
  inv1  gate1268(.a(G23), .O(gate63inter7));
  inv1  gate1269(.a(G299), .O(gate63inter8));
  nand2 gate1270(.a(gate63inter8), .b(gate63inter7), .O(gate63inter9));
  nand2 gate1271(.a(s_103), .b(gate63inter3), .O(gate63inter10));
  nor2  gate1272(.a(gate63inter10), .b(gate63inter9), .O(gate63inter11));
  nor2  gate1273(.a(gate63inter11), .b(gate63inter6), .O(gate63inter12));
  nand2 gate1274(.a(gate63inter12), .b(gate63inter1), .O(G384));
nand2 gate64( .a(G24), .b(G299), .O(G385) );
nand2 gate65( .a(G25), .b(G302), .O(G386) );
nand2 gate66( .a(G26), .b(G302), .O(G387) );
nand2 gate67( .a(G27), .b(G305), .O(G388) );

  xor2  gate813(.a(G305), .b(G28), .O(gate68inter0));
  nand2 gate814(.a(gate68inter0), .b(s_38), .O(gate68inter1));
  and2  gate815(.a(G305), .b(G28), .O(gate68inter2));
  inv1  gate816(.a(s_38), .O(gate68inter3));
  inv1  gate817(.a(s_39), .O(gate68inter4));
  nand2 gate818(.a(gate68inter4), .b(gate68inter3), .O(gate68inter5));
  nor2  gate819(.a(gate68inter5), .b(gate68inter2), .O(gate68inter6));
  inv1  gate820(.a(G28), .O(gate68inter7));
  inv1  gate821(.a(G305), .O(gate68inter8));
  nand2 gate822(.a(gate68inter8), .b(gate68inter7), .O(gate68inter9));
  nand2 gate823(.a(s_39), .b(gate68inter3), .O(gate68inter10));
  nor2  gate824(.a(gate68inter10), .b(gate68inter9), .O(gate68inter11));
  nor2  gate825(.a(gate68inter11), .b(gate68inter6), .O(gate68inter12));
  nand2 gate826(.a(gate68inter12), .b(gate68inter1), .O(G389));
nand2 gate69( .a(G29), .b(G308), .O(G390) );
nand2 gate70( .a(G30), .b(G308), .O(G391) );

  xor2  gate1429(.a(G311), .b(G31), .O(gate71inter0));
  nand2 gate1430(.a(gate71inter0), .b(s_126), .O(gate71inter1));
  and2  gate1431(.a(G311), .b(G31), .O(gate71inter2));
  inv1  gate1432(.a(s_126), .O(gate71inter3));
  inv1  gate1433(.a(s_127), .O(gate71inter4));
  nand2 gate1434(.a(gate71inter4), .b(gate71inter3), .O(gate71inter5));
  nor2  gate1435(.a(gate71inter5), .b(gate71inter2), .O(gate71inter6));
  inv1  gate1436(.a(G31), .O(gate71inter7));
  inv1  gate1437(.a(G311), .O(gate71inter8));
  nand2 gate1438(.a(gate71inter8), .b(gate71inter7), .O(gate71inter9));
  nand2 gate1439(.a(s_127), .b(gate71inter3), .O(gate71inter10));
  nor2  gate1440(.a(gate71inter10), .b(gate71inter9), .O(gate71inter11));
  nor2  gate1441(.a(gate71inter11), .b(gate71inter6), .O(gate71inter12));
  nand2 gate1442(.a(gate71inter12), .b(gate71inter1), .O(G392));
nand2 gate72( .a(G32), .b(G311), .O(G393) );
nand2 gate73( .a(G1), .b(G314), .O(G394) );
nand2 gate74( .a(G5), .b(G314), .O(G395) );

  xor2  gate1611(.a(G317), .b(G9), .O(gate75inter0));
  nand2 gate1612(.a(gate75inter0), .b(s_152), .O(gate75inter1));
  and2  gate1613(.a(G317), .b(G9), .O(gate75inter2));
  inv1  gate1614(.a(s_152), .O(gate75inter3));
  inv1  gate1615(.a(s_153), .O(gate75inter4));
  nand2 gate1616(.a(gate75inter4), .b(gate75inter3), .O(gate75inter5));
  nor2  gate1617(.a(gate75inter5), .b(gate75inter2), .O(gate75inter6));
  inv1  gate1618(.a(G9), .O(gate75inter7));
  inv1  gate1619(.a(G317), .O(gate75inter8));
  nand2 gate1620(.a(gate75inter8), .b(gate75inter7), .O(gate75inter9));
  nand2 gate1621(.a(s_153), .b(gate75inter3), .O(gate75inter10));
  nor2  gate1622(.a(gate75inter10), .b(gate75inter9), .O(gate75inter11));
  nor2  gate1623(.a(gate75inter11), .b(gate75inter6), .O(gate75inter12));
  nand2 gate1624(.a(gate75inter12), .b(gate75inter1), .O(G396));

  xor2  gate603(.a(G317), .b(G13), .O(gate76inter0));
  nand2 gate604(.a(gate76inter0), .b(s_8), .O(gate76inter1));
  and2  gate605(.a(G317), .b(G13), .O(gate76inter2));
  inv1  gate606(.a(s_8), .O(gate76inter3));
  inv1  gate607(.a(s_9), .O(gate76inter4));
  nand2 gate608(.a(gate76inter4), .b(gate76inter3), .O(gate76inter5));
  nor2  gate609(.a(gate76inter5), .b(gate76inter2), .O(gate76inter6));
  inv1  gate610(.a(G13), .O(gate76inter7));
  inv1  gate611(.a(G317), .O(gate76inter8));
  nand2 gate612(.a(gate76inter8), .b(gate76inter7), .O(gate76inter9));
  nand2 gate613(.a(s_9), .b(gate76inter3), .O(gate76inter10));
  nor2  gate614(.a(gate76inter10), .b(gate76inter9), .O(gate76inter11));
  nor2  gate615(.a(gate76inter11), .b(gate76inter6), .O(gate76inter12));
  nand2 gate616(.a(gate76inter12), .b(gate76inter1), .O(G397));
nand2 gate77( .a(G2), .b(G320), .O(G398) );
nand2 gate78( .a(G6), .b(G320), .O(G399) );
nand2 gate79( .a(G10), .b(G323), .O(G400) );

  xor2  gate799(.a(G323), .b(G14), .O(gate80inter0));
  nand2 gate800(.a(gate80inter0), .b(s_36), .O(gate80inter1));
  and2  gate801(.a(G323), .b(G14), .O(gate80inter2));
  inv1  gate802(.a(s_36), .O(gate80inter3));
  inv1  gate803(.a(s_37), .O(gate80inter4));
  nand2 gate804(.a(gate80inter4), .b(gate80inter3), .O(gate80inter5));
  nor2  gate805(.a(gate80inter5), .b(gate80inter2), .O(gate80inter6));
  inv1  gate806(.a(G14), .O(gate80inter7));
  inv1  gate807(.a(G323), .O(gate80inter8));
  nand2 gate808(.a(gate80inter8), .b(gate80inter7), .O(gate80inter9));
  nand2 gate809(.a(s_37), .b(gate80inter3), .O(gate80inter10));
  nor2  gate810(.a(gate80inter10), .b(gate80inter9), .O(gate80inter11));
  nor2  gate811(.a(gate80inter11), .b(gate80inter6), .O(gate80inter12));
  nand2 gate812(.a(gate80inter12), .b(gate80inter1), .O(G401));
nand2 gate81( .a(G3), .b(G326), .O(G402) );

  xor2  gate589(.a(G326), .b(G7), .O(gate82inter0));
  nand2 gate590(.a(gate82inter0), .b(s_6), .O(gate82inter1));
  and2  gate591(.a(G326), .b(G7), .O(gate82inter2));
  inv1  gate592(.a(s_6), .O(gate82inter3));
  inv1  gate593(.a(s_7), .O(gate82inter4));
  nand2 gate594(.a(gate82inter4), .b(gate82inter3), .O(gate82inter5));
  nor2  gate595(.a(gate82inter5), .b(gate82inter2), .O(gate82inter6));
  inv1  gate596(.a(G7), .O(gate82inter7));
  inv1  gate597(.a(G326), .O(gate82inter8));
  nand2 gate598(.a(gate82inter8), .b(gate82inter7), .O(gate82inter9));
  nand2 gate599(.a(s_7), .b(gate82inter3), .O(gate82inter10));
  nor2  gate600(.a(gate82inter10), .b(gate82inter9), .O(gate82inter11));
  nor2  gate601(.a(gate82inter11), .b(gate82inter6), .O(gate82inter12));
  nand2 gate602(.a(gate82inter12), .b(gate82inter1), .O(G403));
nand2 gate83( .a(G11), .b(G329), .O(G404) );

  xor2  gate1625(.a(G329), .b(G15), .O(gate84inter0));
  nand2 gate1626(.a(gate84inter0), .b(s_154), .O(gate84inter1));
  and2  gate1627(.a(G329), .b(G15), .O(gate84inter2));
  inv1  gate1628(.a(s_154), .O(gate84inter3));
  inv1  gate1629(.a(s_155), .O(gate84inter4));
  nand2 gate1630(.a(gate84inter4), .b(gate84inter3), .O(gate84inter5));
  nor2  gate1631(.a(gate84inter5), .b(gate84inter2), .O(gate84inter6));
  inv1  gate1632(.a(G15), .O(gate84inter7));
  inv1  gate1633(.a(G329), .O(gate84inter8));
  nand2 gate1634(.a(gate84inter8), .b(gate84inter7), .O(gate84inter9));
  nand2 gate1635(.a(s_155), .b(gate84inter3), .O(gate84inter10));
  nor2  gate1636(.a(gate84inter10), .b(gate84inter9), .O(gate84inter11));
  nor2  gate1637(.a(gate84inter11), .b(gate84inter6), .O(gate84inter12));
  nand2 gate1638(.a(gate84inter12), .b(gate84inter1), .O(G405));
nand2 gate85( .a(G4), .b(G332), .O(G406) );

  xor2  gate631(.a(G332), .b(G8), .O(gate86inter0));
  nand2 gate632(.a(gate86inter0), .b(s_12), .O(gate86inter1));
  and2  gate633(.a(G332), .b(G8), .O(gate86inter2));
  inv1  gate634(.a(s_12), .O(gate86inter3));
  inv1  gate635(.a(s_13), .O(gate86inter4));
  nand2 gate636(.a(gate86inter4), .b(gate86inter3), .O(gate86inter5));
  nor2  gate637(.a(gate86inter5), .b(gate86inter2), .O(gate86inter6));
  inv1  gate638(.a(G8), .O(gate86inter7));
  inv1  gate639(.a(G332), .O(gate86inter8));
  nand2 gate640(.a(gate86inter8), .b(gate86inter7), .O(gate86inter9));
  nand2 gate641(.a(s_13), .b(gate86inter3), .O(gate86inter10));
  nor2  gate642(.a(gate86inter10), .b(gate86inter9), .O(gate86inter11));
  nor2  gate643(.a(gate86inter11), .b(gate86inter6), .O(gate86inter12));
  nand2 gate644(.a(gate86inter12), .b(gate86inter1), .O(G407));
nand2 gate87( .a(G12), .b(G335), .O(G408) );
nand2 gate88( .a(G16), .b(G335), .O(G409) );

  xor2  gate1303(.a(G338), .b(G17), .O(gate89inter0));
  nand2 gate1304(.a(gate89inter0), .b(s_108), .O(gate89inter1));
  and2  gate1305(.a(G338), .b(G17), .O(gate89inter2));
  inv1  gate1306(.a(s_108), .O(gate89inter3));
  inv1  gate1307(.a(s_109), .O(gate89inter4));
  nand2 gate1308(.a(gate89inter4), .b(gate89inter3), .O(gate89inter5));
  nor2  gate1309(.a(gate89inter5), .b(gate89inter2), .O(gate89inter6));
  inv1  gate1310(.a(G17), .O(gate89inter7));
  inv1  gate1311(.a(G338), .O(gate89inter8));
  nand2 gate1312(.a(gate89inter8), .b(gate89inter7), .O(gate89inter9));
  nand2 gate1313(.a(s_109), .b(gate89inter3), .O(gate89inter10));
  nor2  gate1314(.a(gate89inter10), .b(gate89inter9), .O(gate89inter11));
  nor2  gate1315(.a(gate89inter11), .b(gate89inter6), .O(gate89inter12));
  nand2 gate1316(.a(gate89inter12), .b(gate89inter1), .O(G410));
nand2 gate90( .a(G21), .b(G338), .O(G411) );
nand2 gate91( .a(G25), .b(G341), .O(G412) );
nand2 gate92( .a(G29), .b(G341), .O(G413) );
nand2 gate93( .a(G18), .b(G344), .O(G414) );
nand2 gate94( .a(G22), .b(G344), .O(G415) );
nand2 gate95( .a(G26), .b(G347), .O(G416) );
nand2 gate96( .a(G30), .b(G347), .O(G417) );
nand2 gate97( .a(G19), .b(G350), .O(G418) );

  xor2  gate1709(.a(G350), .b(G23), .O(gate98inter0));
  nand2 gate1710(.a(gate98inter0), .b(s_166), .O(gate98inter1));
  and2  gate1711(.a(G350), .b(G23), .O(gate98inter2));
  inv1  gate1712(.a(s_166), .O(gate98inter3));
  inv1  gate1713(.a(s_167), .O(gate98inter4));
  nand2 gate1714(.a(gate98inter4), .b(gate98inter3), .O(gate98inter5));
  nor2  gate1715(.a(gate98inter5), .b(gate98inter2), .O(gate98inter6));
  inv1  gate1716(.a(G23), .O(gate98inter7));
  inv1  gate1717(.a(G350), .O(gate98inter8));
  nand2 gate1718(.a(gate98inter8), .b(gate98inter7), .O(gate98inter9));
  nand2 gate1719(.a(s_167), .b(gate98inter3), .O(gate98inter10));
  nor2  gate1720(.a(gate98inter10), .b(gate98inter9), .O(gate98inter11));
  nor2  gate1721(.a(gate98inter11), .b(gate98inter6), .O(gate98inter12));
  nand2 gate1722(.a(gate98inter12), .b(gate98inter1), .O(G419));
nand2 gate99( .a(G27), .b(G353), .O(G420) );

  xor2  gate575(.a(G353), .b(G31), .O(gate100inter0));
  nand2 gate576(.a(gate100inter0), .b(s_4), .O(gate100inter1));
  and2  gate577(.a(G353), .b(G31), .O(gate100inter2));
  inv1  gate578(.a(s_4), .O(gate100inter3));
  inv1  gate579(.a(s_5), .O(gate100inter4));
  nand2 gate580(.a(gate100inter4), .b(gate100inter3), .O(gate100inter5));
  nor2  gate581(.a(gate100inter5), .b(gate100inter2), .O(gate100inter6));
  inv1  gate582(.a(G31), .O(gate100inter7));
  inv1  gate583(.a(G353), .O(gate100inter8));
  nand2 gate584(.a(gate100inter8), .b(gate100inter7), .O(gate100inter9));
  nand2 gate585(.a(s_5), .b(gate100inter3), .O(gate100inter10));
  nor2  gate586(.a(gate100inter10), .b(gate100inter9), .O(gate100inter11));
  nor2  gate587(.a(gate100inter11), .b(gate100inter6), .O(gate100inter12));
  nand2 gate588(.a(gate100inter12), .b(gate100inter1), .O(G421));
nand2 gate101( .a(G20), .b(G356), .O(G422) );
nand2 gate102( .a(G24), .b(G356), .O(G423) );
nand2 gate103( .a(G28), .b(G359), .O(G424) );
nand2 gate104( .a(G32), .b(G359), .O(G425) );

  xor2  gate1961(.a(G363), .b(G362), .O(gate105inter0));
  nand2 gate1962(.a(gate105inter0), .b(s_202), .O(gate105inter1));
  and2  gate1963(.a(G363), .b(G362), .O(gate105inter2));
  inv1  gate1964(.a(s_202), .O(gate105inter3));
  inv1  gate1965(.a(s_203), .O(gate105inter4));
  nand2 gate1966(.a(gate105inter4), .b(gate105inter3), .O(gate105inter5));
  nor2  gate1967(.a(gate105inter5), .b(gate105inter2), .O(gate105inter6));
  inv1  gate1968(.a(G362), .O(gate105inter7));
  inv1  gate1969(.a(G363), .O(gate105inter8));
  nand2 gate1970(.a(gate105inter8), .b(gate105inter7), .O(gate105inter9));
  nand2 gate1971(.a(s_203), .b(gate105inter3), .O(gate105inter10));
  nor2  gate1972(.a(gate105inter10), .b(gate105inter9), .O(gate105inter11));
  nor2  gate1973(.a(gate105inter11), .b(gate105inter6), .O(gate105inter12));
  nand2 gate1974(.a(gate105inter12), .b(gate105inter1), .O(G426));
nand2 gate106( .a(G364), .b(G365), .O(G429) );

  xor2  gate1527(.a(G367), .b(G366), .O(gate107inter0));
  nand2 gate1528(.a(gate107inter0), .b(s_140), .O(gate107inter1));
  and2  gate1529(.a(G367), .b(G366), .O(gate107inter2));
  inv1  gate1530(.a(s_140), .O(gate107inter3));
  inv1  gate1531(.a(s_141), .O(gate107inter4));
  nand2 gate1532(.a(gate107inter4), .b(gate107inter3), .O(gate107inter5));
  nor2  gate1533(.a(gate107inter5), .b(gate107inter2), .O(gate107inter6));
  inv1  gate1534(.a(G366), .O(gate107inter7));
  inv1  gate1535(.a(G367), .O(gate107inter8));
  nand2 gate1536(.a(gate107inter8), .b(gate107inter7), .O(gate107inter9));
  nand2 gate1537(.a(s_141), .b(gate107inter3), .O(gate107inter10));
  nor2  gate1538(.a(gate107inter10), .b(gate107inter9), .O(gate107inter11));
  nor2  gate1539(.a(gate107inter11), .b(gate107inter6), .O(gate107inter12));
  nand2 gate1540(.a(gate107inter12), .b(gate107inter1), .O(G432));
nand2 gate108( .a(G368), .b(G369), .O(G435) );
nand2 gate109( .a(G370), .b(G371), .O(G438) );
nand2 gate110( .a(G372), .b(G373), .O(G441) );

  xor2  gate1807(.a(G375), .b(G374), .O(gate111inter0));
  nand2 gate1808(.a(gate111inter0), .b(s_180), .O(gate111inter1));
  and2  gate1809(.a(G375), .b(G374), .O(gate111inter2));
  inv1  gate1810(.a(s_180), .O(gate111inter3));
  inv1  gate1811(.a(s_181), .O(gate111inter4));
  nand2 gate1812(.a(gate111inter4), .b(gate111inter3), .O(gate111inter5));
  nor2  gate1813(.a(gate111inter5), .b(gate111inter2), .O(gate111inter6));
  inv1  gate1814(.a(G374), .O(gate111inter7));
  inv1  gate1815(.a(G375), .O(gate111inter8));
  nand2 gate1816(.a(gate111inter8), .b(gate111inter7), .O(gate111inter9));
  nand2 gate1817(.a(s_181), .b(gate111inter3), .O(gate111inter10));
  nor2  gate1818(.a(gate111inter10), .b(gate111inter9), .O(gate111inter11));
  nor2  gate1819(.a(gate111inter11), .b(gate111inter6), .O(gate111inter12));
  nand2 gate1820(.a(gate111inter12), .b(gate111inter1), .O(G444));
nand2 gate112( .a(G376), .b(G377), .O(G447) );
nand2 gate113( .a(G378), .b(G379), .O(G450) );

  xor2  gate1359(.a(G381), .b(G380), .O(gate114inter0));
  nand2 gate1360(.a(gate114inter0), .b(s_116), .O(gate114inter1));
  and2  gate1361(.a(G381), .b(G380), .O(gate114inter2));
  inv1  gate1362(.a(s_116), .O(gate114inter3));
  inv1  gate1363(.a(s_117), .O(gate114inter4));
  nand2 gate1364(.a(gate114inter4), .b(gate114inter3), .O(gate114inter5));
  nor2  gate1365(.a(gate114inter5), .b(gate114inter2), .O(gate114inter6));
  inv1  gate1366(.a(G380), .O(gate114inter7));
  inv1  gate1367(.a(G381), .O(gate114inter8));
  nand2 gate1368(.a(gate114inter8), .b(gate114inter7), .O(gate114inter9));
  nand2 gate1369(.a(s_117), .b(gate114inter3), .O(gate114inter10));
  nor2  gate1370(.a(gate114inter10), .b(gate114inter9), .O(gate114inter11));
  nor2  gate1371(.a(gate114inter11), .b(gate114inter6), .O(gate114inter12));
  nand2 gate1372(.a(gate114inter12), .b(gate114inter1), .O(G453));
nand2 gate115( .a(G382), .b(G383), .O(G456) );
nand2 gate116( .a(G384), .b(G385), .O(G459) );
nand2 gate117( .a(G386), .b(G387), .O(G462) );

  xor2  gate1065(.a(G389), .b(G388), .O(gate118inter0));
  nand2 gate1066(.a(gate118inter0), .b(s_74), .O(gate118inter1));
  and2  gate1067(.a(G389), .b(G388), .O(gate118inter2));
  inv1  gate1068(.a(s_74), .O(gate118inter3));
  inv1  gate1069(.a(s_75), .O(gate118inter4));
  nand2 gate1070(.a(gate118inter4), .b(gate118inter3), .O(gate118inter5));
  nor2  gate1071(.a(gate118inter5), .b(gate118inter2), .O(gate118inter6));
  inv1  gate1072(.a(G388), .O(gate118inter7));
  inv1  gate1073(.a(G389), .O(gate118inter8));
  nand2 gate1074(.a(gate118inter8), .b(gate118inter7), .O(gate118inter9));
  nand2 gate1075(.a(s_75), .b(gate118inter3), .O(gate118inter10));
  nor2  gate1076(.a(gate118inter10), .b(gate118inter9), .O(gate118inter11));
  nor2  gate1077(.a(gate118inter11), .b(gate118inter6), .O(gate118inter12));
  nand2 gate1078(.a(gate118inter12), .b(gate118inter1), .O(G465));

  xor2  gate1765(.a(G391), .b(G390), .O(gate119inter0));
  nand2 gate1766(.a(gate119inter0), .b(s_174), .O(gate119inter1));
  and2  gate1767(.a(G391), .b(G390), .O(gate119inter2));
  inv1  gate1768(.a(s_174), .O(gate119inter3));
  inv1  gate1769(.a(s_175), .O(gate119inter4));
  nand2 gate1770(.a(gate119inter4), .b(gate119inter3), .O(gate119inter5));
  nor2  gate1771(.a(gate119inter5), .b(gate119inter2), .O(gate119inter6));
  inv1  gate1772(.a(G390), .O(gate119inter7));
  inv1  gate1773(.a(G391), .O(gate119inter8));
  nand2 gate1774(.a(gate119inter8), .b(gate119inter7), .O(gate119inter9));
  nand2 gate1775(.a(s_175), .b(gate119inter3), .O(gate119inter10));
  nor2  gate1776(.a(gate119inter10), .b(gate119inter9), .O(gate119inter11));
  nor2  gate1777(.a(gate119inter11), .b(gate119inter6), .O(gate119inter12));
  nand2 gate1778(.a(gate119inter12), .b(gate119inter1), .O(G468));
nand2 gate120( .a(G392), .b(G393), .O(G471) );
nand2 gate121( .a(G394), .b(G395), .O(G474) );
nand2 gate122( .a(G396), .b(G397), .O(G477) );

  xor2  gate687(.a(G399), .b(G398), .O(gate123inter0));
  nand2 gate688(.a(gate123inter0), .b(s_20), .O(gate123inter1));
  and2  gate689(.a(G399), .b(G398), .O(gate123inter2));
  inv1  gate690(.a(s_20), .O(gate123inter3));
  inv1  gate691(.a(s_21), .O(gate123inter4));
  nand2 gate692(.a(gate123inter4), .b(gate123inter3), .O(gate123inter5));
  nor2  gate693(.a(gate123inter5), .b(gate123inter2), .O(gate123inter6));
  inv1  gate694(.a(G398), .O(gate123inter7));
  inv1  gate695(.a(G399), .O(gate123inter8));
  nand2 gate696(.a(gate123inter8), .b(gate123inter7), .O(gate123inter9));
  nand2 gate697(.a(s_21), .b(gate123inter3), .O(gate123inter10));
  nor2  gate698(.a(gate123inter10), .b(gate123inter9), .O(gate123inter11));
  nor2  gate699(.a(gate123inter11), .b(gate123inter6), .O(gate123inter12));
  nand2 gate700(.a(gate123inter12), .b(gate123inter1), .O(G480));
nand2 gate124( .a(G400), .b(G401), .O(G483) );
nand2 gate125( .a(G402), .b(G403), .O(G486) );
nand2 gate126( .a(G404), .b(G405), .O(G489) );

  xor2  gate1079(.a(G407), .b(G406), .O(gate127inter0));
  nand2 gate1080(.a(gate127inter0), .b(s_76), .O(gate127inter1));
  and2  gate1081(.a(G407), .b(G406), .O(gate127inter2));
  inv1  gate1082(.a(s_76), .O(gate127inter3));
  inv1  gate1083(.a(s_77), .O(gate127inter4));
  nand2 gate1084(.a(gate127inter4), .b(gate127inter3), .O(gate127inter5));
  nor2  gate1085(.a(gate127inter5), .b(gate127inter2), .O(gate127inter6));
  inv1  gate1086(.a(G406), .O(gate127inter7));
  inv1  gate1087(.a(G407), .O(gate127inter8));
  nand2 gate1088(.a(gate127inter8), .b(gate127inter7), .O(gate127inter9));
  nand2 gate1089(.a(s_77), .b(gate127inter3), .O(gate127inter10));
  nor2  gate1090(.a(gate127inter10), .b(gate127inter9), .O(gate127inter11));
  nor2  gate1091(.a(gate127inter11), .b(gate127inter6), .O(gate127inter12));
  nand2 gate1092(.a(gate127inter12), .b(gate127inter1), .O(G492));

  xor2  gate855(.a(G409), .b(G408), .O(gate128inter0));
  nand2 gate856(.a(gate128inter0), .b(s_44), .O(gate128inter1));
  and2  gate857(.a(G409), .b(G408), .O(gate128inter2));
  inv1  gate858(.a(s_44), .O(gate128inter3));
  inv1  gate859(.a(s_45), .O(gate128inter4));
  nand2 gate860(.a(gate128inter4), .b(gate128inter3), .O(gate128inter5));
  nor2  gate861(.a(gate128inter5), .b(gate128inter2), .O(gate128inter6));
  inv1  gate862(.a(G408), .O(gate128inter7));
  inv1  gate863(.a(G409), .O(gate128inter8));
  nand2 gate864(.a(gate128inter8), .b(gate128inter7), .O(gate128inter9));
  nand2 gate865(.a(s_45), .b(gate128inter3), .O(gate128inter10));
  nor2  gate866(.a(gate128inter10), .b(gate128inter9), .O(gate128inter11));
  nor2  gate867(.a(gate128inter11), .b(gate128inter6), .O(gate128inter12));
  nand2 gate868(.a(gate128inter12), .b(gate128inter1), .O(G495));
nand2 gate129( .a(G410), .b(G411), .O(G498) );
nand2 gate130( .a(G412), .b(G413), .O(G501) );
nand2 gate131( .a(G414), .b(G415), .O(G504) );

  xor2  gate1667(.a(G417), .b(G416), .O(gate132inter0));
  nand2 gate1668(.a(gate132inter0), .b(s_160), .O(gate132inter1));
  and2  gate1669(.a(G417), .b(G416), .O(gate132inter2));
  inv1  gate1670(.a(s_160), .O(gate132inter3));
  inv1  gate1671(.a(s_161), .O(gate132inter4));
  nand2 gate1672(.a(gate132inter4), .b(gate132inter3), .O(gate132inter5));
  nor2  gate1673(.a(gate132inter5), .b(gate132inter2), .O(gate132inter6));
  inv1  gate1674(.a(G416), .O(gate132inter7));
  inv1  gate1675(.a(G417), .O(gate132inter8));
  nand2 gate1676(.a(gate132inter8), .b(gate132inter7), .O(gate132inter9));
  nand2 gate1677(.a(s_161), .b(gate132inter3), .O(gate132inter10));
  nor2  gate1678(.a(gate132inter10), .b(gate132inter9), .O(gate132inter11));
  nor2  gate1679(.a(gate132inter11), .b(gate132inter6), .O(gate132inter12));
  nand2 gate1680(.a(gate132inter12), .b(gate132inter1), .O(G507));
nand2 gate133( .a(G418), .b(G419), .O(G510) );
nand2 gate134( .a(G420), .b(G421), .O(G513) );
nand2 gate135( .a(G422), .b(G423), .O(G516) );
nand2 gate136( .a(G424), .b(G425), .O(G519) );
nand2 gate137( .a(G426), .b(G429), .O(G522) );

  xor2  gate1499(.a(G435), .b(G432), .O(gate138inter0));
  nand2 gate1500(.a(gate138inter0), .b(s_136), .O(gate138inter1));
  and2  gate1501(.a(G435), .b(G432), .O(gate138inter2));
  inv1  gate1502(.a(s_136), .O(gate138inter3));
  inv1  gate1503(.a(s_137), .O(gate138inter4));
  nand2 gate1504(.a(gate138inter4), .b(gate138inter3), .O(gate138inter5));
  nor2  gate1505(.a(gate138inter5), .b(gate138inter2), .O(gate138inter6));
  inv1  gate1506(.a(G432), .O(gate138inter7));
  inv1  gate1507(.a(G435), .O(gate138inter8));
  nand2 gate1508(.a(gate138inter8), .b(gate138inter7), .O(gate138inter9));
  nand2 gate1509(.a(s_137), .b(gate138inter3), .O(gate138inter10));
  nor2  gate1510(.a(gate138inter10), .b(gate138inter9), .O(gate138inter11));
  nor2  gate1511(.a(gate138inter11), .b(gate138inter6), .O(gate138inter12));
  nand2 gate1512(.a(gate138inter12), .b(gate138inter1), .O(G525));
nand2 gate139( .a(G438), .b(G441), .O(G528) );
nand2 gate140( .a(G444), .b(G447), .O(G531) );
nand2 gate141( .a(G450), .b(G453), .O(G534) );
nand2 gate142( .a(G456), .b(G459), .O(G537) );
nand2 gate143( .a(G462), .b(G465), .O(G540) );

  xor2  gate1135(.a(G471), .b(G468), .O(gate144inter0));
  nand2 gate1136(.a(gate144inter0), .b(s_84), .O(gate144inter1));
  and2  gate1137(.a(G471), .b(G468), .O(gate144inter2));
  inv1  gate1138(.a(s_84), .O(gate144inter3));
  inv1  gate1139(.a(s_85), .O(gate144inter4));
  nand2 gate1140(.a(gate144inter4), .b(gate144inter3), .O(gate144inter5));
  nor2  gate1141(.a(gate144inter5), .b(gate144inter2), .O(gate144inter6));
  inv1  gate1142(.a(G468), .O(gate144inter7));
  inv1  gate1143(.a(G471), .O(gate144inter8));
  nand2 gate1144(.a(gate144inter8), .b(gate144inter7), .O(gate144inter9));
  nand2 gate1145(.a(s_85), .b(gate144inter3), .O(gate144inter10));
  nor2  gate1146(.a(gate144inter10), .b(gate144inter9), .O(gate144inter11));
  nor2  gate1147(.a(gate144inter11), .b(gate144inter6), .O(gate144inter12));
  nand2 gate1148(.a(gate144inter12), .b(gate144inter1), .O(G543));

  xor2  gate1513(.a(G477), .b(G474), .O(gate145inter0));
  nand2 gate1514(.a(gate145inter0), .b(s_138), .O(gate145inter1));
  and2  gate1515(.a(G477), .b(G474), .O(gate145inter2));
  inv1  gate1516(.a(s_138), .O(gate145inter3));
  inv1  gate1517(.a(s_139), .O(gate145inter4));
  nand2 gate1518(.a(gate145inter4), .b(gate145inter3), .O(gate145inter5));
  nor2  gate1519(.a(gate145inter5), .b(gate145inter2), .O(gate145inter6));
  inv1  gate1520(.a(G474), .O(gate145inter7));
  inv1  gate1521(.a(G477), .O(gate145inter8));
  nand2 gate1522(.a(gate145inter8), .b(gate145inter7), .O(gate145inter9));
  nand2 gate1523(.a(s_139), .b(gate145inter3), .O(gate145inter10));
  nor2  gate1524(.a(gate145inter10), .b(gate145inter9), .O(gate145inter11));
  nor2  gate1525(.a(gate145inter11), .b(gate145inter6), .O(gate145inter12));
  nand2 gate1526(.a(gate145inter12), .b(gate145inter1), .O(G546));
nand2 gate146( .a(G480), .b(G483), .O(G549) );
nand2 gate147( .a(G486), .b(G489), .O(G552) );
nand2 gate148( .a(G492), .b(G495), .O(G555) );
nand2 gate149( .a(G498), .b(G501), .O(G558) );

  xor2  gate1751(.a(G507), .b(G504), .O(gate150inter0));
  nand2 gate1752(.a(gate150inter0), .b(s_172), .O(gate150inter1));
  and2  gate1753(.a(G507), .b(G504), .O(gate150inter2));
  inv1  gate1754(.a(s_172), .O(gate150inter3));
  inv1  gate1755(.a(s_173), .O(gate150inter4));
  nand2 gate1756(.a(gate150inter4), .b(gate150inter3), .O(gate150inter5));
  nor2  gate1757(.a(gate150inter5), .b(gate150inter2), .O(gate150inter6));
  inv1  gate1758(.a(G504), .O(gate150inter7));
  inv1  gate1759(.a(G507), .O(gate150inter8));
  nand2 gate1760(.a(gate150inter8), .b(gate150inter7), .O(gate150inter9));
  nand2 gate1761(.a(s_173), .b(gate150inter3), .O(gate150inter10));
  nor2  gate1762(.a(gate150inter10), .b(gate150inter9), .O(gate150inter11));
  nor2  gate1763(.a(gate150inter11), .b(gate150inter6), .O(gate150inter12));
  nand2 gate1764(.a(gate150inter12), .b(gate150inter1), .O(G561));
nand2 gate151( .a(G510), .b(G513), .O(G564) );

  xor2  gate869(.a(G519), .b(G516), .O(gate152inter0));
  nand2 gate870(.a(gate152inter0), .b(s_46), .O(gate152inter1));
  and2  gate871(.a(G519), .b(G516), .O(gate152inter2));
  inv1  gate872(.a(s_46), .O(gate152inter3));
  inv1  gate873(.a(s_47), .O(gate152inter4));
  nand2 gate874(.a(gate152inter4), .b(gate152inter3), .O(gate152inter5));
  nor2  gate875(.a(gate152inter5), .b(gate152inter2), .O(gate152inter6));
  inv1  gate876(.a(G516), .O(gate152inter7));
  inv1  gate877(.a(G519), .O(gate152inter8));
  nand2 gate878(.a(gate152inter8), .b(gate152inter7), .O(gate152inter9));
  nand2 gate879(.a(s_47), .b(gate152inter3), .O(gate152inter10));
  nor2  gate880(.a(gate152inter10), .b(gate152inter9), .O(gate152inter11));
  nor2  gate881(.a(gate152inter11), .b(gate152inter6), .O(gate152inter12));
  nand2 gate882(.a(gate152inter12), .b(gate152inter1), .O(G567));
nand2 gate153( .a(G426), .b(G522), .O(G570) );
nand2 gate154( .a(G429), .b(G522), .O(G571) );

  xor2  gate1569(.a(G525), .b(G432), .O(gate155inter0));
  nand2 gate1570(.a(gate155inter0), .b(s_146), .O(gate155inter1));
  and2  gate1571(.a(G525), .b(G432), .O(gate155inter2));
  inv1  gate1572(.a(s_146), .O(gate155inter3));
  inv1  gate1573(.a(s_147), .O(gate155inter4));
  nand2 gate1574(.a(gate155inter4), .b(gate155inter3), .O(gate155inter5));
  nor2  gate1575(.a(gate155inter5), .b(gate155inter2), .O(gate155inter6));
  inv1  gate1576(.a(G432), .O(gate155inter7));
  inv1  gate1577(.a(G525), .O(gate155inter8));
  nand2 gate1578(.a(gate155inter8), .b(gate155inter7), .O(gate155inter9));
  nand2 gate1579(.a(s_147), .b(gate155inter3), .O(gate155inter10));
  nor2  gate1580(.a(gate155inter10), .b(gate155inter9), .O(gate155inter11));
  nor2  gate1581(.a(gate155inter11), .b(gate155inter6), .O(gate155inter12));
  nand2 gate1582(.a(gate155inter12), .b(gate155inter1), .O(G572));
nand2 gate156( .a(G435), .b(G525), .O(G573) );
nand2 gate157( .a(G438), .b(G528), .O(G574) );

  xor2  gate981(.a(G528), .b(G441), .O(gate158inter0));
  nand2 gate982(.a(gate158inter0), .b(s_62), .O(gate158inter1));
  and2  gate983(.a(G528), .b(G441), .O(gate158inter2));
  inv1  gate984(.a(s_62), .O(gate158inter3));
  inv1  gate985(.a(s_63), .O(gate158inter4));
  nand2 gate986(.a(gate158inter4), .b(gate158inter3), .O(gate158inter5));
  nor2  gate987(.a(gate158inter5), .b(gate158inter2), .O(gate158inter6));
  inv1  gate988(.a(G441), .O(gate158inter7));
  inv1  gate989(.a(G528), .O(gate158inter8));
  nand2 gate990(.a(gate158inter8), .b(gate158inter7), .O(gate158inter9));
  nand2 gate991(.a(s_63), .b(gate158inter3), .O(gate158inter10));
  nor2  gate992(.a(gate158inter10), .b(gate158inter9), .O(gate158inter11));
  nor2  gate993(.a(gate158inter11), .b(gate158inter6), .O(gate158inter12));
  nand2 gate994(.a(gate158inter12), .b(gate158inter1), .O(G575));
nand2 gate159( .a(G444), .b(G531), .O(G576) );
nand2 gate160( .a(G447), .b(G531), .O(G577) );
nand2 gate161( .a(G450), .b(G534), .O(G578) );
nand2 gate162( .a(G453), .b(G534), .O(G579) );

  xor2  gate1191(.a(G537), .b(G456), .O(gate163inter0));
  nand2 gate1192(.a(gate163inter0), .b(s_92), .O(gate163inter1));
  and2  gate1193(.a(G537), .b(G456), .O(gate163inter2));
  inv1  gate1194(.a(s_92), .O(gate163inter3));
  inv1  gate1195(.a(s_93), .O(gate163inter4));
  nand2 gate1196(.a(gate163inter4), .b(gate163inter3), .O(gate163inter5));
  nor2  gate1197(.a(gate163inter5), .b(gate163inter2), .O(gate163inter6));
  inv1  gate1198(.a(G456), .O(gate163inter7));
  inv1  gate1199(.a(G537), .O(gate163inter8));
  nand2 gate1200(.a(gate163inter8), .b(gate163inter7), .O(gate163inter9));
  nand2 gate1201(.a(s_93), .b(gate163inter3), .O(gate163inter10));
  nor2  gate1202(.a(gate163inter10), .b(gate163inter9), .O(gate163inter11));
  nor2  gate1203(.a(gate163inter11), .b(gate163inter6), .O(gate163inter12));
  nand2 gate1204(.a(gate163inter12), .b(gate163inter1), .O(G580));
nand2 gate164( .a(G459), .b(G537), .O(G581) );
nand2 gate165( .a(G462), .b(G540), .O(G582) );

  xor2  gate1037(.a(G540), .b(G465), .O(gate166inter0));
  nand2 gate1038(.a(gate166inter0), .b(s_70), .O(gate166inter1));
  and2  gate1039(.a(G540), .b(G465), .O(gate166inter2));
  inv1  gate1040(.a(s_70), .O(gate166inter3));
  inv1  gate1041(.a(s_71), .O(gate166inter4));
  nand2 gate1042(.a(gate166inter4), .b(gate166inter3), .O(gate166inter5));
  nor2  gate1043(.a(gate166inter5), .b(gate166inter2), .O(gate166inter6));
  inv1  gate1044(.a(G465), .O(gate166inter7));
  inv1  gate1045(.a(G540), .O(gate166inter8));
  nand2 gate1046(.a(gate166inter8), .b(gate166inter7), .O(gate166inter9));
  nand2 gate1047(.a(s_71), .b(gate166inter3), .O(gate166inter10));
  nor2  gate1048(.a(gate166inter10), .b(gate166inter9), .O(gate166inter11));
  nor2  gate1049(.a(gate166inter11), .b(gate166inter6), .O(gate166inter12));
  nand2 gate1050(.a(gate166inter12), .b(gate166inter1), .O(G583));

  xor2  gate1919(.a(G543), .b(G468), .O(gate167inter0));
  nand2 gate1920(.a(gate167inter0), .b(s_196), .O(gate167inter1));
  and2  gate1921(.a(G543), .b(G468), .O(gate167inter2));
  inv1  gate1922(.a(s_196), .O(gate167inter3));
  inv1  gate1923(.a(s_197), .O(gate167inter4));
  nand2 gate1924(.a(gate167inter4), .b(gate167inter3), .O(gate167inter5));
  nor2  gate1925(.a(gate167inter5), .b(gate167inter2), .O(gate167inter6));
  inv1  gate1926(.a(G468), .O(gate167inter7));
  inv1  gate1927(.a(G543), .O(gate167inter8));
  nand2 gate1928(.a(gate167inter8), .b(gate167inter7), .O(gate167inter9));
  nand2 gate1929(.a(s_197), .b(gate167inter3), .O(gate167inter10));
  nor2  gate1930(.a(gate167inter10), .b(gate167inter9), .O(gate167inter11));
  nor2  gate1931(.a(gate167inter11), .b(gate167inter6), .O(gate167inter12));
  nand2 gate1932(.a(gate167inter12), .b(gate167inter1), .O(G584));
nand2 gate168( .a(G471), .b(G543), .O(G585) );
nand2 gate169( .a(G474), .b(G546), .O(G586) );
nand2 gate170( .a(G477), .b(G546), .O(G587) );

  xor2  gate1541(.a(G549), .b(G480), .O(gate171inter0));
  nand2 gate1542(.a(gate171inter0), .b(s_142), .O(gate171inter1));
  and2  gate1543(.a(G549), .b(G480), .O(gate171inter2));
  inv1  gate1544(.a(s_142), .O(gate171inter3));
  inv1  gate1545(.a(s_143), .O(gate171inter4));
  nand2 gate1546(.a(gate171inter4), .b(gate171inter3), .O(gate171inter5));
  nor2  gate1547(.a(gate171inter5), .b(gate171inter2), .O(gate171inter6));
  inv1  gate1548(.a(G480), .O(gate171inter7));
  inv1  gate1549(.a(G549), .O(gate171inter8));
  nand2 gate1550(.a(gate171inter8), .b(gate171inter7), .O(gate171inter9));
  nand2 gate1551(.a(s_143), .b(gate171inter3), .O(gate171inter10));
  nor2  gate1552(.a(gate171inter10), .b(gate171inter9), .O(gate171inter11));
  nor2  gate1553(.a(gate171inter11), .b(gate171inter6), .O(gate171inter12));
  nand2 gate1554(.a(gate171inter12), .b(gate171inter1), .O(G588));
nand2 gate172( .a(G483), .b(G549), .O(G589) );

  xor2  gate1583(.a(G552), .b(G486), .O(gate173inter0));
  nand2 gate1584(.a(gate173inter0), .b(s_148), .O(gate173inter1));
  and2  gate1585(.a(G552), .b(G486), .O(gate173inter2));
  inv1  gate1586(.a(s_148), .O(gate173inter3));
  inv1  gate1587(.a(s_149), .O(gate173inter4));
  nand2 gate1588(.a(gate173inter4), .b(gate173inter3), .O(gate173inter5));
  nor2  gate1589(.a(gate173inter5), .b(gate173inter2), .O(gate173inter6));
  inv1  gate1590(.a(G486), .O(gate173inter7));
  inv1  gate1591(.a(G552), .O(gate173inter8));
  nand2 gate1592(.a(gate173inter8), .b(gate173inter7), .O(gate173inter9));
  nand2 gate1593(.a(s_149), .b(gate173inter3), .O(gate173inter10));
  nor2  gate1594(.a(gate173inter10), .b(gate173inter9), .O(gate173inter11));
  nor2  gate1595(.a(gate173inter11), .b(gate173inter6), .O(gate173inter12));
  nand2 gate1596(.a(gate173inter12), .b(gate173inter1), .O(G590));
nand2 gate174( .a(G489), .b(G552), .O(G591) );
nand2 gate175( .a(G492), .b(G555), .O(G592) );

  xor2  gate911(.a(G555), .b(G495), .O(gate176inter0));
  nand2 gate912(.a(gate176inter0), .b(s_52), .O(gate176inter1));
  and2  gate913(.a(G555), .b(G495), .O(gate176inter2));
  inv1  gate914(.a(s_52), .O(gate176inter3));
  inv1  gate915(.a(s_53), .O(gate176inter4));
  nand2 gate916(.a(gate176inter4), .b(gate176inter3), .O(gate176inter5));
  nor2  gate917(.a(gate176inter5), .b(gate176inter2), .O(gate176inter6));
  inv1  gate918(.a(G495), .O(gate176inter7));
  inv1  gate919(.a(G555), .O(gate176inter8));
  nand2 gate920(.a(gate176inter8), .b(gate176inter7), .O(gate176inter9));
  nand2 gate921(.a(s_53), .b(gate176inter3), .O(gate176inter10));
  nor2  gate922(.a(gate176inter10), .b(gate176inter9), .O(gate176inter11));
  nor2  gate923(.a(gate176inter11), .b(gate176inter6), .O(gate176inter12));
  nand2 gate924(.a(gate176inter12), .b(gate176inter1), .O(G593));
nand2 gate177( .a(G498), .b(G558), .O(G594) );
nand2 gate178( .a(G501), .b(G558), .O(G595) );
nand2 gate179( .a(G504), .b(G561), .O(G596) );
nand2 gate180( .a(G507), .b(G561), .O(G597) );
nand2 gate181( .a(G510), .b(G564), .O(G598) );
nand2 gate182( .a(G513), .b(G564), .O(G599) );
nand2 gate183( .a(G516), .b(G567), .O(G600) );
nand2 gate184( .a(G519), .b(G567), .O(G601) );
nand2 gate185( .a(G570), .b(G571), .O(G602) );
nand2 gate186( .a(G572), .b(G573), .O(G607) );
nand2 gate187( .a(G574), .b(G575), .O(G612) );
nand2 gate188( .a(G576), .b(G577), .O(G617) );
nand2 gate189( .a(G578), .b(G579), .O(G622) );

  xor2  gate1415(.a(G581), .b(G580), .O(gate190inter0));
  nand2 gate1416(.a(gate190inter0), .b(s_124), .O(gate190inter1));
  and2  gate1417(.a(G581), .b(G580), .O(gate190inter2));
  inv1  gate1418(.a(s_124), .O(gate190inter3));
  inv1  gate1419(.a(s_125), .O(gate190inter4));
  nand2 gate1420(.a(gate190inter4), .b(gate190inter3), .O(gate190inter5));
  nor2  gate1421(.a(gate190inter5), .b(gate190inter2), .O(gate190inter6));
  inv1  gate1422(.a(G580), .O(gate190inter7));
  inv1  gate1423(.a(G581), .O(gate190inter8));
  nand2 gate1424(.a(gate190inter8), .b(gate190inter7), .O(gate190inter9));
  nand2 gate1425(.a(s_125), .b(gate190inter3), .O(gate190inter10));
  nor2  gate1426(.a(gate190inter10), .b(gate190inter9), .O(gate190inter11));
  nor2  gate1427(.a(gate190inter11), .b(gate190inter6), .O(gate190inter12));
  nand2 gate1428(.a(gate190inter12), .b(gate190inter1), .O(G627));
nand2 gate191( .a(G582), .b(G583), .O(G632) );
nand2 gate192( .a(G584), .b(G585), .O(G637) );
nand2 gate193( .a(G586), .b(G587), .O(G642) );

  xor2  gate1373(.a(G589), .b(G588), .O(gate194inter0));
  nand2 gate1374(.a(gate194inter0), .b(s_118), .O(gate194inter1));
  and2  gate1375(.a(G589), .b(G588), .O(gate194inter2));
  inv1  gate1376(.a(s_118), .O(gate194inter3));
  inv1  gate1377(.a(s_119), .O(gate194inter4));
  nand2 gate1378(.a(gate194inter4), .b(gate194inter3), .O(gate194inter5));
  nor2  gate1379(.a(gate194inter5), .b(gate194inter2), .O(gate194inter6));
  inv1  gate1380(.a(G588), .O(gate194inter7));
  inv1  gate1381(.a(G589), .O(gate194inter8));
  nand2 gate1382(.a(gate194inter8), .b(gate194inter7), .O(gate194inter9));
  nand2 gate1383(.a(s_119), .b(gate194inter3), .O(gate194inter10));
  nor2  gate1384(.a(gate194inter10), .b(gate194inter9), .O(gate194inter11));
  nor2  gate1385(.a(gate194inter11), .b(gate194inter6), .O(gate194inter12));
  nand2 gate1386(.a(gate194inter12), .b(gate194inter1), .O(G645));

  xor2  gate995(.a(G591), .b(G590), .O(gate195inter0));
  nand2 gate996(.a(gate195inter0), .b(s_64), .O(gate195inter1));
  and2  gate997(.a(G591), .b(G590), .O(gate195inter2));
  inv1  gate998(.a(s_64), .O(gate195inter3));
  inv1  gate999(.a(s_65), .O(gate195inter4));
  nand2 gate1000(.a(gate195inter4), .b(gate195inter3), .O(gate195inter5));
  nor2  gate1001(.a(gate195inter5), .b(gate195inter2), .O(gate195inter6));
  inv1  gate1002(.a(G590), .O(gate195inter7));
  inv1  gate1003(.a(G591), .O(gate195inter8));
  nand2 gate1004(.a(gate195inter8), .b(gate195inter7), .O(gate195inter9));
  nand2 gate1005(.a(s_65), .b(gate195inter3), .O(gate195inter10));
  nor2  gate1006(.a(gate195inter10), .b(gate195inter9), .O(gate195inter11));
  nor2  gate1007(.a(gate195inter11), .b(gate195inter6), .O(gate195inter12));
  nand2 gate1008(.a(gate195inter12), .b(gate195inter1), .O(G648));
nand2 gate196( .a(G592), .b(G593), .O(G651) );
nand2 gate197( .a(G594), .b(G595), .O(G654) );
nand2 gate198( .a(G596), .b(G597), .O(G657) );
nand2 gate199( .a(G598), .b(G599), .O(G660) );
nand2 gate200( .a(G600), .b(G601), .O(G663) );
nand2 gate201( .a(G602), .b(G607), .O(G666) );
nand2 gate202( .a(G612), .b(G617), .O(G669) );
nand2 gate203( .a(G602), .b(G612), .O(G672) );

  xor2  gate561(.a(G617), .b(G607), .O(gate204inter0));
  nand2 gate562(.a(gate204inter0), .b(s_2), .O(gate204inter1));
  and2  gate563(.a(G617), .b(G607), .O(gate204inter2));
  inv1  gate564(.a(s_2), .O(gate204inter3));
  inv1  gate565(.a(s_3), .O(gate204inter4));
  nand2 gate566(.a(gate204inter4), .b(gate204inter3), .O(gate204inter5));
  nor2  gate567(.a(gate204inter5), .b(gate204inter2), .O(gate204inter6));
  inv1  gate568(.a(G607), .O(gate204inter7));
  inv1  gate569(.a(G617), .O(gate204inter8));
  nand2 gate570(.a(gate204inter8), .b(gate204inter7), .O(gate204inter9));
  nand2 gate571(.a(s_3), .b(gate204inter3), .O(gate204inter10));
  nor2  gate572(.a(gate204inter10), .b(gate204inter9), .O(gate204inter11));
  nor2  gate573(.a(gate204inter11), .b(gate204inter6), .O(gate204inter12));
  nand2 gate574(.a(gate204inter12), .b(gate204inter1), .O(G675));

  xor2  gate1723(.a(G627), .b(G622), .O(gate205inter0));
  nand2 gate1724(.a(gate205inter0), .b(s_168), .O(gate205inter1));
  and2  gate1725(.a(G627), .b(G622), .O(gate205inter2));
  inv1  gate1726(.a(s_168), .O(gate205inter3));
  inv1  gate1727(.a(s_169), .O(gate205inter4));
  nand2 gate1728(.a(gate205inter4), .b(gate205inter3), .O(gate205inter5));
  nor2  gate1729(.a(gate205inter5), .b(gate205inter2), .O(gate205inter6));
  inv1  gate1730(.a(G622), .O(gate205inter7));
  inv1  gate1731(.a(G627), .O(gate205inter8));
  nand2 gate1732(.a(gate205inter8), .b(gate205inter7), .O(gate205inter9));
  nand2 gate1733(.a(s_169), .b(gate205inter3), .O(gate205inter10));
  nor2  gate1734(.a(gate205inter10), .b(gate205inter9), .O(gate205inter11));
  nor2  gate1735(.a(gate205inter11), .b(gate205inter6), .O(gate205inter12));
  nand2 gate1736(.a(gate205inter12), .b(gate205inter1), .O(G678));
nand2 gate206( .a(G632), .b(G637), .O(G681) );
nand2 gate207( .a(G622), .b(G632), .O(G684) );
nand2 gate208( .a(G627), .b(G637), .O(G687) );
nand2 gate209( .a(G602), .b(G666), .O(G690) );

  xor2  gate1331(.a(G666), .b(G607), .O(gate210inter0));
  nand2 gate1332(.a(gate210inter0), .b(s_112), .O(gate210inter1));
  and2  gate1333(.a(G666), .b(G607), .O(gate210inter2));
  inv1  gate1334(.a(s_112), .O(gate210inter3));
  inv1  gate1335(.a(s_113), .O(gate210inter4));
  nand2 gate1336(.a(gate210inter4), .b(gate210inter3), .O(gate210inter5));
  nor2  gate1337(.a(gate210inter5), .b(gate210inter2), .O(gate210inter6));
  inv1  gate1338(.a(G607), .O(gate210inter7));
  inv1  gate1339(.a(G666), .O(gate210inter8));
  nand2 gate1340(.a(gate210inter8), .b(gate210inter7), .O(gate210inter9));
  nand2 gate1341(.a(s_113), .b(gate210inter3), .O(gate210inter10));
  nor2  gate1342(.a(gate210inter10), .b(gate210inter9), .O(gate210inter11));
  nor2  gate1343(.a(gate210inter11), .b(gate210inter6), .O(gate210inter12));
  nand2 gate1344(.a(gate210inter12), .b(gate210inter1), .O(G691));
nand2 gate211( .a(G612), .b(G669), .O(G692) );
nand2 gate212( .a(G617), .b(G669), .O(G693) );

  xor2  gate1933(.a(G672), .b(G602), .O(gate213inter0));
  nand2 gate1934(.a(gate213inter0), .b(s_198), .O(gate213inter1));
  and2  gate1935(.a(G672), .b(G602), .O(gate213inter2));
  inv1  gate1936(.a(s_198), .O(gate213inter3));
  inv1  gate1937(.a(s_199), .O(gate213inter4));
  nand2 gate1938(.a(gate213inter4), .b(gate213inter3), .O(gate213inter5));
  nor2  gate1939(.a(gate213inter5), .b(gate213inter2), .O(gate213inter6));
  inv1  gate1940(.a(G602), .O(gate213inter7));
  inv1  gate1941(.a(G672), .O(gate213inter8));
  nand2 gate1942(.a(gate213inter8), .b(gate213inter7), .O(gate213inter9));
  nand2 gate1943(.a(s_199), .b(gate213inter3), .O(gate213inter10));
  nor2  gate1944(.a(gate213inter10), .b(gate213inter9), .O(gate213inter11));
  nor2  gate1945(.a(gate213inter11), .b(gate213inter6), .O(gate213inter12));
  nand2 gate1946(.a(gate213inter12), .b(gate213inter1), .O(G694));
nand2 gate214( .a(G612), .b(G672), .O(G695) );
nand2 gate215( .a(G607), .b(G675), .O(G696) );
nand2 gate216( .a(G617), .b(G675), .O(G697) );
nand2 gate217( .a(G622), .b(G678), .O(G698) );
nand2 gate218( .a(G627), .b(G678), .O(G699) );
nand2 gate219( .a(G632), .b(G681), .O(G700) );
nand2 gate220( .a(G637), .b(G681), .O(G701) );
nand2 gate221( .a(G622), .b(G684), .O(G702) );

  xor2  gate1485(.a(G684), .b(G632), .O(gate222inter0));
  nand2 gate1486(.a(gate222inter0), .b(s_134), .O(gate222inter1));
  and2  gate1487(.a(G684), .b(G632), .O(gate222inter2));
  inv1  gate1488(.a(s_134), .O(gate222inter3));
  inv1  gate1489(.a(s_135), .O(gate222inter4));
  nand2 gate1490(.a(gate222inter4), .b(gate222inter3), .O(gate222inter5));
  nor2  gate1491(.a(gate222inter5), .b(gate222inter2), .O(gate222inter6));
  inv1  gate1492(.a(G632), .O(gate222inter7));
  inv1  gate1493(.a(G684), .O(gate222inter8));
  nand2 gate1494(.a(gate222inter8), .b(gate222inter7), .O(gate222inter9));
  nand2 gate1495(.a(s_135), .b(gate222inter3), .O(gate222inter10));
  nor2  gate1496(.a(gate222inter10), .b(gate222inter9), .O(gate222inter11));
  nor2  gate1497(.a(gate222inter11), .b(gate222inter6), .O(gate222inter12));
  nand2 gate1498(.a(gate222inter12), .b(gate222inter1), .O(G703));
nand2 gate223( .a(G627), .b(G687), .O(G704) );

  xor2  gate1793(.a(G687), .b(G637), .O(gate224inter0));
  nand2 gate1794(.a(gate224inter0), .b(s_178), .O(gate224inter1));
  and2  gate1795(.a(G687), .b(G637), .O(gate224inter2));
  inv1  gate1796(.a(s_178), .O(gate224inter3));
  inv1  gate1797(.a(s_179), .O(gate224inter4));
  nand2 gate1798(.a(gate224inter4), .b(gate224inter3), .O(gate224inter5));
  nor2  gate1799(.a(gate224inter5), .b(gate224inter2), .O(gate224inter6));
  inv1  gate1800(.a(G637), .O(gate224inter7));
  inv1  gate1801(.a(G687), .O(gate224inter8));
  nand2 gate1802(.a(gate224inter8), .b(gate224inter7), .O(gate224inter9));
  nand2 gate1803(.a(s_179), .b(gate224inter3), .O(gate224inter10));
  nor2  gate1804(.a(gate224inter10), .b(gate224inter9), .O(gate224inter11));
  nor2  gate1805(.a(gate224inter11), .b(gate224inter6), .O(gate224inter12));
  nand2 gate1806(.a(gate224inter12), .b(gate224inter1), .O(G705));

  xor2  gate1177(.a(G691), .b(G690), .O(gate225inter0));
  nand2 gate1178(.a(gate225inter0), .b(s_90), .O(gate225inter1));
  and2  gate1179(.a(G691), .b(G690), .O(gate225inter2));
  inv1  gate1180(.a(s_90), .O(gate225inter3));
  inv1  gate1181(.a(s_91), .O(gate225inter4));
  nand2 gate1182(.a(gate225inter4), .b(gate225inter3), .O(gate225inter5));
  nor2  gate1183(.a(gate225inter5), .b(gate225inter2), .O(gate225inter6));
  inv1  gate1184(.a(G690), .O(gate225inter7));
  inv1  gate1185(.a(G691), .O(gate225inter8));
  nand2 gate1186(.a(gate225inter8), .b(gate225inter7), .O(gate225inter9));
  nand2 gate1187(.a(s_91), .b(gate225inter3), .O(gate225inter10));
  nor2  gate1188(.a(gate225inter10), .b(gate225inter9), .O(gate225inter11));
  nor2  gate1189(.a(gate225inter11), .b(gate225inter6), .O(gate225inter12));
  nand2 gate1190(.a(gate225inter12), .b(gate225inter1), .O(G706));
nand2 gate226( .a(G692), .b(G693), .O(G709) );

  xor2  gate1233(.a(G695), .b(G694), .O(gate227inter0));
  nand2 gate1234(.a(gate227inter0), .b(s_98), .O(gate227inter1));
  and2  gate1235(.a(G695), .b(G694), .O(gate227inter2));
  inv1  gate1236(.a(s_98), .O(gate227inter3));
  inv1  gate1237(.a(s_99), .O(gate227inter4));
  nand2 gate1238(.a(gate227inter4), .b(gate227inter3), .O(gate227inter5));
  nor2  gate1239(.a(gate227inter5), .b(gate227inter2), .O(gate227inter6));
  inv1  gate1240(.a(G694), .O(gate227inter7));
  inv1  gate1241(.a(G695), .O(gate227inter8));
  nand2 gate1242(.a(gate227inter8), .b(gate227inter7), .O(gate227inter9));
  nand2 gate1243(.a(s_99), .b(gate227inter3), .O(gate227inter10));
  nor2  gate1244(.a(gate227inter10), .b(gate227inter9), .O(gate227inter11));
  nor2  gate1245(.a(gate227inter11), .b(gate227inter6), .O(gate227inter12));
  nand2 gate1246(.a(gate227inter12), .b(gate227inter1), .O(G712));
nand2 gate228( .a(G696), .b(G697), .O(G715) );

  xor2  gate2017(.a(G699), .b(G698), .O(gate229inter0));
  nand2 gate2018(.a(gate229inter0), .b(s_210), .O(gate229inter1));
  and2  gate2019(.a(G699), .b(G698), .O(gate229inter2));
  inv1  gate2020(.a(s_210), .O(gate229inter3));
  inv1  gate2021(.a(s_211), .O(gate229inter4));
  nand2 gate2022(.a(gate229inter4), .b(gate229inter3), .O(gate229inter5));
  nor2  gate2023(.a(gate229inter5), .b(gate229inter2), .O(gate229inter6));
  inv1  gate2024(.a(G698), .O(gate229inter7));
  inv1  gate2025(.a(G699), .O(gate229inter8));
  nand2 gate2026(.a(gate229inter8), .b(gate229inter7), .O(gate229inter9));
  nand2 gate2027(.a(s_211), .b(gate229inter3), .O(gate229inter10));
  nor2  gate2028(.a(gate229inter10), .b(gate229inter9), .O(gate229inter11));
  nor2  gate2029(.a(gate229inter11), .b(gate229inter6), .O(gate229inter12));
  nand2 gate2030(.a(gate229inter12), .b(gate229inter1), .O(G718));
nand2 gate230( .a(G700), .b(G701), .O(G721) );
nand2 gate231( .a(G702), .b(G703), .O(G724) );
nand2 gate232( .a(G704), .b(G705), .O(G727) );

  xor2  gate939(.a(G718), .b(G242), .O(gate233inter0));
  nand2 gate940(.a(gate233inter0), .b(s_56), .O(gate233inter1));
  and2  gate941(.a(G718), .b(G242), .O(gate233inter2));
  inv1  gate942(.a(s_56), .O(gate233inter3));
  inv1  gate943(.a(s_57), .O(gate233inter4));
  nand2 gate944(.a(gate233inter4), .b(gate233inter3), .O(gate233inter5));
  nor2  gate945(.a(gate233inter5), .b(gate233inter2), .O(gate233inter6));
  inv1  gate946(.a(G242), .O(gate233inter7));
  inv1  gate947(.a(G718), .O(gate233inter8));
  nand2 gate948(.a(gate233inter8), .b(gate233inter7), .O(gate233inter9));
  nand2 gate949(.a(s_57), .b(gate233inter3), .O(gate233inter10));
  nor2  gate950(.a(gate233inter10), .b(gate233inter9), .O(gate233inter11));
  nor2  gate951(.a(gate233inter11), .b(gate233inter6), .O(gate233inter12));
  nand2 gate952(.a(gate233inter12), .b(gate233inter1), .O(G730));
nand2 gate234( .a(G245), .b(G721), .O(G733) );

  xor2  gate1387(.a(G724), .b(G248), .O(gate235inter0));
  nand2 gate1388(.a(gate235inter0), .b(s_120), .O(gate235inter1));
  and2  gate1389(.a(G724), .b(G248), .O(gate235inter2));
  inv1  gate1390(.a(s_120), .O(gate235inter3));
  inv1  gate1391(.a(s_121), .O(gate235inter4));
  nand2 gate1392(.a(gate235inter4), .b(gate235inter3), .O(gate235inter5));
  nor2  gate1393(.a(gate235inter5), .b(gate235inter2), .O(gate235inter6));
  inv1  gate1394(.a(G248), .O(gate235inter7));
  inv1  gate1395(.a(G724), .O(gate235inter8));
  nand2 gate1396(.a(gate235inter8), .b(gate235inter7), .O(gate235inter9));
  nand2 gate1397(.a(s_121), .b(gate235inter3), .O(gate235inter10));
  nor2  gate1398(.a(gate235inter10), .b(gate235inter9), .O(gate235inter11));
  nor2  gate1399(.a(gate235inter11), .b(gate235inter6), .O(gate235inter12));
  nand2 gate1400(.a(gate235inter12), .b(gate235inter1), .O(G736));
nand2 gate236( .a(G251), .b(G727), .O(G739) );

  xor2  gate1877(.a(G706), .b(G254), .O(gate237inter0));
  nand2 gate1878(.a(gate237inter0), .b(s_190), .O(gate237inter1));
  and2  gate1879(.a(G706), .b(G254), .O(gate237inter2));
  inv1  gate1880(.a(s_190), .O(gate237inter3));
  inv1  gate1881(.a(s_191), .O(gate237inter4));
  nand2 gate1882(.a(gate237inter4), .b(gate237inter3), .O(gate237inter5));
  nor2  gate1883(.a(gate237inter5), .b(gate237inter2), .O(gate237inter6));
  inv1  gate1884(.a(G254), .O(gate237inter7));
  inv1  gate1885(.a(G706), .O(gate237inter8));
  nand2 gate1886(.a(gate237inter8), .b(gate237inter7), .O(gate237inter9));
  nand2 gate1887(.a(s_191), .b(gate237inter3), .O(gate237inter10));
  nor2  gate1888(.a(gate237inter10), .b(gate237inter9), .O(gate237inter11));
  nor2  gate1889(.a(gate237inter11), .b(gate237inter6), .O(gate237inter12));
  nand2 gate1890(.a(gate237inter12), .b(gate237inter1), .O(G742));
nand2 gate238( .a(G257), .b(G709), .O(G745) );
nand2 gate239( .a(G260), .b(G712), .O(G748) );
nand2 gate240( .a(G263), .b(G715), .O(G751) );
nand2 gate241( .a(G242), .b(G730), .O(G754) );
nand2 gate242( .a(G718), .b(G730), .O(G755) );

  xor2  gate1275(.a(G733), .b(G245), .O(gate243inter0));
  nand2 gate1276(.a(gate243inter0), .b(s_104), .O(gate243inter1));
  and2  gate1277(.a(G733), .b(G245), .O(gate243inter2));
  inv1  gate1278(.a(s_104), .O(gate243inter3));
  inv1  gate1279(.a(s_105), .O(gate243inter4));
  nand2 gate1280(.a(gate243inter4), .b(gate243inter3), .O(gate243inter5));
  nor2  gate1281(.a(gate243inter5), .b(gate243inter2), .O(gate243inter6));
  inv1  gate1282(.a(G245), .O(gate243inter7));
  inv1  gate1283(.a(G733), .O(gate243inter8));
  nand2 gate1284(.a(gate243inter8), .b(gate243inter7), .O(gate243inter9));
  nand2 gate1285(.a(s_105), .b(gate243inter3), .O(gate243inter10));
  nor2  gate1286(.a(gate243inter10), .b(gate243inter9), .O(gate243inter11));
  nor2  gate1287(.a(gate243inter11), .b(gate243inter6), .O(gate243inter12));
  nand2 gate1288(.a(gate243inter12), .b(gate243inter1), .O(G756));
nand2 gate244( .a(G721), .b(G733), .O(G757) );
nand2 gate245( .a(G248), .b(G736), .O(G758) );
nand2 gate246( .a(G724), .b(G736), .O(G759) );

  xor2  gate1821(.a(G739), .b(G251), .O(gate247inter0));
  nand2 gate1822(.a(gate247inter0), .b(s_182), .O(gate247inter1));
  and2  gate1823(.a(G739), .b(G251), .O(gate247inter2));
  inv1  gate1824(.a(s_182), .O(gate247inter3));
  inv1  gate1825(.a(s_183), .O(gate247inter4));
  nand2 gate1826(.a(gate247inter4), .b(gate247inter3), .O(gate247inter5));
  nor2  gate1827(.a(gate247inter5), .b(gate247inter2), .O(gate247inter6));
  inv1  gate1828(.a(G251), .O(gate247inter7));
  inv1  gate1829(.a(G739), .O(gate247inter8));
  nand2 gate1830(.a(gate247inter8), .b(gate247inter7), .O(gate247inter9));
  nand2 gate1831(.a(s_183), .b(gate247inter3), .O(gate247inter10));
  nor2  gate1832(.a(gate247inter10), .b(gate247inter9), .O(gate247inter11));
  nor2  gate1833(.a(gate247inter11), .b(gate247inter6), .O(gate247inter12));
  nand2 gate1834(.a(gate247inter12), .b(gate247inter1), .O(G760));
nand2 gate248( .a(G727), .b(G739), .O(G761) );
nand2 gate249( .a(G254), .b(G742), .O(G762) );
nand2 gate250( .a(G706), .b(G742), .O(G763) );
nand2 gate251( .a(G257), .b(G745), .O(G764) );
nand2 gate252( .a(G709), .b(G745), .O(G765) );
nand2 gate253( .a(G260), .b(G748), .O(G766) );
nand2 gate254( .a(G712), .b(G748), .O(G767) );
nand2 gate255( .a(G263), .b(G751), .O(G768) );
nand2 gate256( .a(G715), .b(G751), .O(G769) );
nand2 gate257( .a(G754), .b(G755), .O(G770) );
nand2 gate258( .a(G756), .b(G757), .O(G773) );
nand2 gate259( .a(G758), .b(G759), .O(G776) );
nand2 gate260( .a(G760), .b(G761), .O(G779) );

  xor2  gate1905(.a(G763), .b(G762), .O(gate261inter0));
  nand2 gate1906(.a(gate261inter0), .b(s_194), .O(gate261inter1));
  and2  gate1907(.a(G763), .b(G762), .O(gate261inter2));
  inv1  gate1908(.a(s_194), .O(gate261inter3));
  inv1  gate1909(.a(s_195), .O(gate261inter4));
  nand2 gate1910(.a(gate261inter4), .b(gate261inter3), .O(gate261inter5));
  nor2  gate1911(.a(gate261inter5), .b(gate261inter2), .O(gate261inter6));
  inv1  gate1912(.a(G762), .O(gate261inter7));
  inv1  gate1913(.a(G763), .O(gate261inter8));
  nand2 gate1914(.a(gate261inter8), .b(gate261inter7), .O(gate261inter9));
  nand2 gate1915(.a(s_195), .b(gate261inter3), .O(gate261inter10));
  nor2  gate1916(.a(gate261inter10), .b(gate261inter9), .O(gate261inter11));
  nor2  gate1917(.a(gate261inter11), .b(gate261inter6), .O(gate261inter12));
  nand2 gate1918(.a(gate261inter12), .b(gate261inter1), .O(G782));

  xor2  gate715(.a(G765), .b(G764), .O(gate262inter0));
  nand2 gate716(.a(gate262inter0), .b(s_24), .O(gate262inter1));
  and2  gate717(.a(G765), .b(G764), .O(gate262inter2));
  inv1  gate718(.a(s_24), .O(gate262inter3));
  inv1  gate719(.a(s_25), .O(gate262inter4));
  nand2 gate720(.a(gate262inter4), .b(gate262inter3), .O(gate262inter5));
  nor2  gate721(.a(gate262inter5), .b(gate262inter2), .O(gate262inter6));
  inv1  gate722(.a(G764), .O(gate262inter7));
  inv1  gate723(.a(G765), .O(gate262inter8));
  nand2 gate724(.a(gate262inter8), .b(gate262inter7), .O(gate262inter9));
  nand2 gate725(.a(s_25), .b(gate262inter3), .O(gate262inter10));
  nor2  gate726(.a(gate262inter10), .b(gate262inter9), .O(gate262inter11));
  nor2  gate727(.a(gate262inter11), .b(gate262inter6), .O(gate262inter12));
  nand2 gate728(.a(gate262inter12), .b(gate262inter1), .O(G785));

  xor2  gate1555(.a(G767), .b(G766), .O(gate263inter0));
  nand2 gate1556(.a(gate263inter0), .b(s_144), .O(gate263inter1));
  and2  gate1557(.a(G767), .b(G766), .O(gate263inter2));
  inv1  gate1558(.a(s_144), .O(gate263inter3));
  inv1  gate1559(.a(s_145), .O(gate263inter4));
  nand2 gate1560(.a(gate263inter4), .b(gate263inter3), .O(gate263inter5));
  nor2  gate1561(.a(gate263inter5), .b(gate263inter2), .O(gate263inter6));
  inv1  gate1562(.a(G766), .O(gate263inter7));
  inv1  gate1563(.a(G767), .O(gate263inter8));
  nand2 gate1564(.a(gate263inter8), .b(gate263inter7), .O(gate263inter9));
  nand2 gate1565(.a(s_145), .b(gate263inter3), .O(gate263inter10));
  nor2  gate1566(.a(gate263inter10), .b(gate263inter9), .O(gate263inter11));
  nor2  gate1567(.a(gate263inter11), .b(gate263inter6), .O(gate263inter12));
  nand2 gate1568(.a(gate263inter12), .b(gate263inter1), .O(G788));
nand2 gate264( .a(G768), .b(G769), .O(G791) );
nand2 gate265( .a(G642), .b(G770), .O(G794) );

  xor2  gate1289(.a(G773), .b(G645), .O(gate266inter0));
  nand2 gate1290(.a(gate266inter0), .b(s_106), .O(gate266inter1));
  and2  gate1291(.a(G773), .b(G645), .O(gate266inter2));
  inv1  gate1292(.a(s_106), .O(gate266inter3));
  inv1  gate1293(.a(s_107), .O(gate266inter4));
  nand2 gate1294(.a(gate266inter4), .b(gate266inter3), .O(gate266inter5));
  nor2  gate1295(.a(gate266inter5), .b(gate266inter2), .O(gate266inter6));
  inv1  gate1296(.a(G645), .O(gate266inter7));
  inv1  gate1297(.a(G773), .O(gate266inter8));
  nand2 gate1298(.a(gate266inter8), .b(gate266inter7), .O(gate266inter9));
  nand2 gate1299(.a(s_107), .b(gate266inter3), .O(gate266inter10));
  nor2  gate1300(.a(gate266inter10), .b(gate266inter9), .O(gate266inter11));
  nor2  gate1301(.a(gate266inter11), .b(gate266inter6), .O(gate266inter12));
  nand2 gate1302(.a(gate266inter12), .b(gate266inter1), .O(G797));

  xor2  gate1681(.a(G776), .b(G648), .O(gate267inter0));
  nand2 gate1682(.a(gate267inter0), .b(s_162), .O(gate267inter1));
  and2  gate1683(.a(G776), .b(G648), .O(gate267inter2));
  inv1  gate1684(.a(s_162), .O(gate267inter3));
  inv1  gate1685(.a(s_163), .O(gate267inter4));
  nand2 gate1686(.a(gate267inter4), .b(gate267inter3), .O(gate267inter5));
  nor2  gate1687(.a(gate267inter5), .b(gate267inter2), .O(gate267inter6));
  inv1  gate1688(.a(G648), .O(gate267inter7));
  inv1  gate1689(.a(G776), .O(gate267inter8));
  nand2 gate1690(.a(gate267inter8), .b(gate267inter7), .O(gate267inter9));
  nand2 gate1691(.a(s_163), .b(gate267inter3), .O(gate267inter10));
  nor2  gate1692(.a(gate267inter10), .b(gate267inter9), .O(gate267inter11));
  nor2  gate1693(.a(gate267inter11), .b(gate267inter6), .O(gate267inter12));
  nand2 gate1694(.a(gate267inter12), .b(gate267inter1), .O(G800));
nand2 gate268( .a(G651), .b(G779), .O(G803) );
nand2 gate269( .a(G654), .b(G782), .O(G806) );
nand2 gate270( .a(G657), .b(G785), .O(G809) );
nand2 gate271( .a(G660), .b(G788), .O(G812) );
nand2 gate272( .a(G663), .b(G791), .O(G815) );
nand2 gate273( .a(G642), .b(G794), .O(G818) );
nand2 gate274( .a(G770), .b(G794), .O(G819) );
nand2 gate275( .a(G645), .b(G797), .O(G820) );
nand2 gate276( .a(G773), .b(G797), .O(G821) );
nand2 gate277( .a(G648), .b(G800), .O(G822) );
nand2 gate278( .a(G776), .b(G800), .O(G823) );
nand2 gate279( .a(G651), .b(G803), .O(G824) );

  xor2  gate1317(.a(G803), .b(G779), .O(gate280inter0));
  nand2 gate1318(.a(gate280inter0), .b(s_110), .O(gate280inter1));
  and2  gate1319(.a(G803), .b(G779), .O(gate280inter2));
  inv1  gate1320(.a(s_110), .O(gate280inter3));
  inv1  gate1321(.a(s_111), .O(gate280inter4));
  nand2 gate1322(.a(gate280inter4), .b(gate280inter3), .O(gate280inter5));
  nor2  gate1323(.a(gate280inter5), .b(gate280inter2), .O(gate280inter6));
  inv1  gate1324(.a(G779), .O(gate280inter7));
  inv1  gate1325(.a(G803), .O(gate280inter8));
  nand2 gate1326(.a(gate280inter8), .b(gate280inter7), .O(gate280inter9));
  nand2 gate1327(.a(s_111), .b(gate280inter3), .O(gate280inter10));
  nor2  gate1328(.a(gate280inter10), .b(gate280inter9), .O(gate280inter11));
  nor2  gate1329(.a(gate280inter11), .b(gate280inter6), .O(gate280inter12));
  nand2 gate1330(.a(gate280inter12), .b(gate280inter1), .O(G825));

  xor2  gate729(.a(G806), .b(G654), .O(gate281inter0));
  nand2 gate730(.a(gate281inter0), .b(s_26), .O(gate281inter1));
  and2  gate731(.a(G806), .b(G654), .O(gate281inter2));
  inv1  gate732(.a(s_26), .O(gate281inter3));
  inv1  gate733(.a(s_27), .O(gate281inter4));
  nand2 gate734(.a(gate281inter4), .b(gate281inter3), .O(gate281inter5));
  nor2  gate735(.a(gate281inter5), .b(gate281inter2), .O(gate281inter6));
  inv1  gate736(.a(G654), .O(gate281inter7));
  inv1  gate737(.a(G806), .O(gate281inter8));
  nand2 gate738(.a(gate281inter8), .b(gate281inter7), .O(gate281inter9));
  nand2 gate739(.a(s_27), .b(gate281inter3), .O(gate281inter10));
  nor2  gate740(.a(gate281inter10), .b(gate281inter9), .O(gate281inter11));
  nor2  gate741(.a(gate281inter11), .b(gate281inter6), .O(gate281inter12));
  nand2 gate742(.a(gate281inter12), .b(gate281inter1), .O(G826));
nand2 gate282( .a(G782), .b(G806), .O(G827) );
nand2 gate283( .a(G657), .b(G809), .O(G828) );

  xor2  gate1975(.a(G809), .b(G785), .O(gate284inter0));
  nand2 gate1976(.a(gate284inter0), .b(s_204), .O(gate284inter1));
  and2  gate1977(.a(G809), .b(G785), .O(gate284inter2));
  inv1  gate1978(.a(s_204), .O(gate284inter3));
  inv1  gate1979(.a(s_205), .O(gate284inter4));
  nand2 gate1980(.a(gate284inter4), .b(gate284inter3), .O(gate284inter5));
  nor2  gate1981(.a(gate284inter5), .b(gate284inter2), .O(gate284inter6));
  inv1  gate1982(.a(G785), .O(gate284inter7));
  inv1  gate1983(.a(G809), .O(gate284inter8));
  nand2 gate1984(.a(gate284inter8), .b(gate284inter7), .O(gate284inter9));
  nand2 gate1985(.a(s_205), .b(gate284inter3), .O(gate284inter10));
  nor2  gate1986(.a(gate284inter10), .b(gate284inter9), .O(gate284inter11));
  nor2  gate1987(.a(gate284inter11), .b(gate284inter6), .O(gate284inter12));
  nand2 gate1988(.a(gate284inter12), .b(gate284inter1), .O(G829));

  xor2  gate1107(.a(G812), .b(G660), .O(gate285inter0));
  nand2 gate1108(.a(gate285inter0), .b(s_80), .O(gate285inter1));
  and2  gate1109(.a(G812), .b(G660), .O(gate285inter2));
  inv1  gate1110(.a(s_80), .O(gate285inter3));
  inv1  gate1111(.a(s_81), .O(gate285inter4));
  nand2 gate1112(.a(gate285inter4), .b(gate285inter3), .O(gate285inter5));
  nor2  gate1113(.a(gate285inter5), .b(gate285inter2), .O(gate285inter6));
  inv1  gate1114(.a(G660), .O(gate285inter7));
  inv1  gate1115(.a(G812), .O(gate285inter8));
  nand2 gate1116(.a(gate285inter8), .b(gate285inter7), .O(gate285inter9));
  nand2 gate1117(.a(s_81), .b(gate285inter3), .O(gate285inter10));
  nor2  gate1118(.a(gate285inter10), .b(gate285inter9), .O(gate285inter11));
  nor2  gate1119(.a(gate285inter11), .b(gate285inter6), .O(gate285inter12));
  nand2 gate1120(.a(gate285inter12), .b(gate285inter1), .O(G830));
nand2 gate286( .a(G788), .b(G812), .O(G831) );

  xor2  gate785(.a(G815), .b(G663), .O(gate287inter0));
  nand2 gate786(.a(gate287inter0), .b(s_34), .O(gate287inter1));
  and2  gate787(.a(G815), .b(G663), .O(gate287inter2));
  inv1  gate788(.a(s_34), .O(gate287inter3));
  inv1  gate789(.a(s_35), .O(gate287inter4));
  nand2 gate790(.a(gate287inter4), .b(gate287inter3), .O(gate287inter5));
  nor2  gate791(.a(gate287inter5), .b(gate287inter2), .O(gate287inter6));
  inv1  gate792(.a(G663), .O(gate287inter7));
  inv1  gate793(.a(G815), .O(gate287inter8));
  nand2 gate794(.a(gate287inter8), .b(gate287inter7), .O(gate287inter9));
  nand2 gate795(.a(s_35), .b(gate287inter3), .O(gate287inter10));
  nor2  gate796(.a(gate287inter10), .b(gate287inter9), .O(gate287inter11));
  nor2  gate797(.a(gate287inter11), .b(gate287inter6), .O(gate287inter12));
  nand2 gate798(.a(gate287inter12), .b(gate287inter1), .O(G832));
nand2 gate288( .a(G791), .b(G815), .O(G833) );

  xor2  gate617(.a(G819), .b(G818), .O(gate289inter0));
  nand2 gate618(.a(gate289inter0), .b(s_10), .O(gate289inter1));
  and2  gate619(.a(G819), .b(G818), .O(gate289inter2));
  inv1  gate620(.a(s_10), .O(gate289inter3));
  inv1  gate621(.a(s_11), .O(gate289inter4));
  nand2 gate622(.a(gate289inter4), .b(gate289inter3), .O(gate289inter5));
  nor2  gate623(.a(gate289inter5), .b(gate289inter2), .O(gate289inter6));
  inv1  gate624(.a(G818), .O(gate289inter7));
  inv1  gate625(.a(G819), .O(gate289inter8));
  nand2 gate626(.a(gate289inter8), .b(gate289inter7), .O(gate289inter9));
  nand2 gate627(.a(s_11), .b(gate289inter3), .O(gate289inter10));
  nor2  gate628(.a(gate289inter10), .b(gate289inter9), .O(gate289inter11));
  nor2  gate629(.a(gate289inter11), .b(gate289inter6), .O(gate289inter12));
  nand2 gate630(.a(gate289inter12), .b(gate289inter1), .O(G834));

  xor2  gate645(.a(G821), .b(G820), .O(gate290inter0));
  nand2 gate646(.a(gate290inter0), .b(s_14), .O(gate290inter1));
  and2  gate647(.a(G821), .b(G820), .O(gate290inter2));
  inv1  gate648(.a(s_14), .O(gate290inter3));
  inv1  gate649(.a(s_15), .O(gate290inter4));
  nand2 gate650(.a(gate290inter4), .b(gate290inter3), .O(gate290inter5));
  nor2  gate651(.a(gate290inter5), .b(gate290inter2), .O(gate290inter6));
  inv1  gate652(.a(G820), .O(gate290inter7));
  inv1  gate653(.a(G821), .O(gate290inter8));
  nand2 gate654(.a(gate290inter8), .b(gate290inter7), .O(gate290inter9));
  nand2 gate655(.a(s_15), .b(gate290inter3), .O(gate290inter10));
  nor2  gate656(.a(gate290inter10), .b(gate290inter9), .O(gate290inter11));
  nor2  gate657(.a(gate290inter11), .b(gate290inter6), .O(gate290inter12));
  nand2 gate658(.a(gate290inter12), .b(gate290inter1), .O(G847));
nand2 gate291( .a(G822), .b(G823), .O(G860) );
nand2 gate292( .a(G824), .b(G825), .O(G873) );
nand2 gate293( .a(G828), .b(G829), .O(G886) );

  xor2  gate2003(.a(G833), .b(G832), .O(gate294inter0));
  nand2 gate2004(.a(gate294inter0), .b(s_208), .O(gate294inter1));
  and2  gate2005(.a(G833), .b(G832), .O(gate294inter2));
  inv1  gate2006(.a(s_208), .O(gate294inter3));
  inv1  gate2007(.a(s_209), .O(gate294inter4));
  nand2 gate2008(.a(gate294inter4), .b(gate294inter3), .O(gate294inter5));
  nor2  gate2009(.a(gate294inter5), .b(gate294inter2), .O(gate294inter6));
  inv1  gate2010(.a(G832), .O(gate294inter7));
  inv1  gate2011(.a(G833), .O(gate294inter8));
  nand2 gate2012(.a(gate294inter8), .b(gate294inter7), .O(gate294inter9));
  nand2 gate2013(.a(s_209), .b(gate294inter3), .O(gate294inter10));
  nor2  gate2014(.a(gate294inter10), .b(gate294inter9), .O(gate294inter11));
  nor2  gate2015(.a(gate294inter11), .b(gate294inter6), .O(gate294inter12));
  nand2 gate2016(.a(gate294inter12), .b(gate294inter1), .O(G899));

  xor2  gate1849(.a(G831), .b(G830), .O(gate295inter0));
  nand2 gate1850(.a(gate295inter0), .b(s_186), .O(gate295inter1));
  and2  gate1851(.a(G831), .b(G830), .O(gate295inter2));
  inv1  gate1852(.a(s_186), .O(gate295inter3));
  inv1  gate1853(.a(s_187), .O(gate295inter4));
  nand2 gate1854(.a(gate295inter4), .b(gate295inter3), .O(gate295inter5));
  nor2  gate1855(.a(gate295inter5), .b(gate295inter2), .O(gate295inter6));
  inv1  gate1856(.a(G830), .O(gate295inter7));
  inv1  gate1857(.a(G831), .O(gate295inter8));
  nand2 gate1858(.a(gate295inter8), .b(gate295inter7), .O(gate295inter9));
  nand2 gate1859(.a(s_187), .b(gate295inter3), .O(gate295inter10));
  nor2  gate1860(.a(gate295inter10), .b(gate295inter9), .O(gate295inter11));
  nor2  gate1861(.a(gate295inter11), .b(gate295inter6), .O(gate295inter12));
  nand2 gate1862(.a(gate295inter12), .b(gate295inter1), .O(G912));
nand2 gate296( .a(G826), .b(G827), .O(G925) );
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );
nand2 gate387( .a(G1), .b(G1036), .O(G1132) );
nand2 gate388( .a(G2), .b(G1039), .O(G1135) );
nand2 gate389( .a(G3), .b(G1042), .O(G1138) );
nand2 gate390( .a(G4), .b(G1045), .O(G1141) );

  xor2  gate1093(.a(G1048), .b(G5), .O(gate391inter0));
  nand2 gate1094(.a(gate391inter0), .b(s_78), .O(gate391inter1));
  and2  gate1095(.a(G1048), .b(G5), .O(gate391inter2));
  inv1  gate1096(.a(s_78), .O(gate391inter3));
  inv1  gate1097(.a(s_79), .O(gate391inter4));
  nand2 gate1098(.a(gate391inter4), .b(gate391inter3), .O(gate391inter5));
  nor2  gate1099(.a(gate391inter5), .b(gate391inter2), .O(gate391inter6));
  inv1  gate1100(.a(G5), .O(gate391inter7));
  inv1  gate1101(.a(G1048), .O(gate391inter8));
  nand2 gate1102(.a(gate391inter8), .b(gate391inter7), .O(gate391inter9));
  nand2 gate1103(.a(s_79), .b(gate391inter3), .O(gate391inter10));
  nor2  gate1104(.a(gate391inter10), .b(gate391inter9), .O(gate391inter11));
  nor2  gate1105(.a(gate391inter11), .b(gate391inter6), .O(gate391inter12));
  nand2 gate1106(.a(gate391inter12), .b(gate391inter1), .O(G1144));
nand2 gate392( .a(G6), .b(G1051), .O(G1147) );
nand2 gate393( .a(G7), .b(G1054), .O(G1150) );
nand2 gate394( .a(G8), .b(G1057), .O(G1153) );
nand2 gate395( .a(G9), .b(G1060), .O(G1156) );
nand2 gate396( .a(G10), .b(G1063), .O(G1159) );
nand2 gate397( .a(G11), .b(G1066), .O(G1162) );

  xor2  gate757(.a(G1069), .b(G12), .O(gate398inter0));
  nand2 gate758(.a(gate398inter0), .b(s_30), .O(gate398inter1));
  and2  gate759(.a(G1069), .b(G12), .O(gate398inter2));
  inv1  gate760(.a(s_30), .O(gate398inter3));
  inv1  gate761(.a(s_31), .O(gate398inter4));
  nand2 gate762(.a(gate398inter4), .b(gate398inter3), .O(gate398inter5));
  nor2  gate763(.a(gate398inter5), .b(gate398inter2), .O(gate398inter6));
  inv1  gate764(.a(G12), .O(gate398inter7));
  inv1  gate765(.a(G1069), .O(gate398inter8));
  nand2 gate766(.a(gate398inter8), .b(gate398inter7), .O(gate398inter9));
  nand2 gate767(.a(s_31), .b(gate398inter3), .O(gate398inter10));
  nor2  gate768(.a(gate398inter10), .b(gate398inter9), .O(gate398inter11));
  nor2  gate769(.a(gate398inter11), .b(gate398inter6), .O(gate398inter12));
  nand2 gate770(.a(gate398inter12), .b(gate398inter1), .O(G1165));
nand2 gate399( .a(G13), .b(G1072), .O(G1168) );
nand2 gate400( .a(G14), .b(G1075), .O(G1171) );

  xor2  gate659(.a(G1078), .b(G15), .O(gate401inter0));
  nand2 gate660(.a(gate401inter0), .b(s_16), .O(gate401inter1));
  and2  gate661(.a(G1078), .b(G15), .O(gate401inter2));
  inv1  gate662(.a(s_16), .O(gate401inter3));
  inv1  gate663(.a(s_17), .O(gate401inter4));
  nand2 gate664(.a(gate401inter4), .b(gate401inter3), .O(gate401inter5));
  nor2  gate665(.a(gate401inter5), .b(gate401inter2), .O(gate401inter6));
  inv1  gate666(.a(G15), .O(gate401inter7));
  inv1  gate667(.a(G1078), .O(gate401inter8));
  nand2 gate668(.a(gate401inter8), .b(gate401inter7), .O(gate401inter9));
  nand2 gate669(.a(s_17), .b(gate401inter3), .O(gate401inter10));
  nor2  gate670(.a(gate401inter10), .b(gate401inter9), .O(gate401inter11));
  nor2  gate671(.a(gate401inter11), .b(gate401inter6), .O(gate401inter12));
  nand2 gate672(.a(gate401inter12), .b(gate401inter1), .O(G1174));
nand2 gate402( .a(G16), .b(G1081), .O(G1177) );
nand2 gate403( .a(G17), .b(G1084), .O(G1180) );
nand2 gate404( .a(G18), .b(G1087), .O(G1183) );
nand2 gate405( .a(G19), .b(G1090), .O(G1186) );
nand2 gate406( .a(G20), .b(G1093), .O(G1189) );
nand2 gate407( .a(G21), .b(G1096), .O(G1192) );
nand2 gate408( .a(G22), .b(G1099), .O(G1195) );
nand2 gate409( .a(G23), .b(G1102), .O(G1198) );

  xor2  gate1205(.a(G1105), .b(G24), .O(gate410inter0));
  nand2 gate1206(.a(gate410inter0), .b(s_94), .O(gate410inter1));
  and2  gate1207(.a(G1105), .b(G24), .O(gate410inter2));
  inv1  gate1208(.a(s_94), .O(gate410inter3));
  inv1  gate1209(.a(s_95), .O(gate410inter4));
  nand2 gate1210(.a(gate410inter4), .b(gate410inter3), .O(gate410inter5));
  nor2  gate1211(.a(gate410inter5), .b(gate410inter2), .O(gate410inter6));
  inv1  gate1212(.a(G24), .O(gate410inter7));
  inv1  gate1213(.a(G1105), .O(gate410inter8));
  nand2 gate1214(.a(gate410inter8), .b(gate410inter7), .O(gate410inter9));
  nand2 gate1215(.a(s_95), .b(gate410inter3), .O(gate410inter10));
  nor2  gate1216(.a(gate410inter10), .b(gate410inter9), .O(gate410inter11));
  nor2  gate1217(.a(gate410inter11), .b(gate410inter6), .O(gate410inter12));
  nand2 gate1218(.a(gate410inter12), .b(gate410inter1), .O(G1201));
nand2 gate411( .a(G25), .b(G1108), .O(G1204) );
nand2 gate412( .a(G26), .b(G1111), .O(G1207) );
nand2 gate413( .a(G27), .b(G1114), .O(G1210) );
nand2 gate414( .a(G28), .b(G1117), .O(G1213) );
nand2 gate415( .a(G29), .b(G1120), .O(G1216) );
nand2 gate416( .a(G30), .b(G1123), .O(G1219) );
nand2 gate417( .a(G31), .b(G1126), .O(G1222) );
nand2 gate418( .a(G32), .b(G1129), .O(G1225) );
nand2 gate419( .a(G1), .b(G1132), .O(G1228) );
nand2 gate420( .a(G1036), .b(G1132), .O(G1229) );
nand2 gate421( .a(G2), .b(G1135), .O(G1230) );
nand2 gate422( .a(G1039), .b(G1135), .O(G1231) );
nand2 gate423( .a(G3), .b(G1138), .O(G1232) );
nand2 gate424( .a(G1042), .b(G1138), .O(G1233) );
nand2 gate425( .a(G4), .b(G1141), .O(G1234) );
nand2 gate426( .a(G1045), .b(G1141), .O(G1235) );
nand2 gate427( .a(G5), .b(G1144), .O(G1236) );
nand2 gate428( .a(G1048), .b(G1144), .O(G1237) );
nand2 gate429( .a(G6), .b(G1147), .O(G1238) );

  xor2  gate1947(.a(G1147), .b(G1051), .O(gate430inter0));
  nand2 gate1948(.a(gate430inter0), .b(s_200), .O(gate430inter1));
  and2  gate1949(.a(G1147), .b(G1051), .O(gate430inter2));
  inv1  gate1950(.a(s_200), .O(gate430inter3));
  inv1  gate1951(.a(s_201), .O(gate430inter4));
  nand2 gate1952(.a(gate430inter4), .b(gate430inter3), .O(gate430inter5));
  nor2  gate1953(.a(gate430inter5), .b(gate430inter2), .O(gate430inter6));
  inv1  gate1954(.a(G1051), .O(gate430inter7));
  inv1  gate1955(.a(G1147), .O(gate430inter8));
  nand2 gate1956(.a(gate430inter8), .b(gate430inter7), .O(gate430inter9));
  nand2 gate1957(.a(s_201), .b(gate430inter3), .O(gate430inter10));
  nor2  gate1958(.a(gate430inter10), .b(gate430inter9), .O(gate430inter11));
  nor2  gate1959(.a(gate430inter11), .b(gate430inter6), .O(gate430inter12));
  nand2 gate1960(.a(gate430inter12), .b(gate430inter1), .O(G1239));

  xor2  gate1443(.a(G1150), .b(G7), .O(gate431inter0));
  nand2 gate1444(.a(gate431inter0), .b(s_128), .O(gate431inter1));
  and2  gate1445(.a(G1150), .b(G7), .O(gate431inter2));
  inv1  gate1446(.a(s_128), .O(gate431inter3));
  inv1  gate1447(.a(s_129), .O(gate431inter4));
  nand2 gate1448(.a(gate431inter4), .b(gate431inter3), .O(gate431inter5));
  nor2  gate1449(.a(gate431inter5), .b(gate431inter2), .O(gate431inter6));
  inv1  gate1450(.a(G7), .O(gate431inter7));
  inv1  gate1451(.a(G1150), .O(gate431inter8));
  nand2 gate1452(.a(gate431inter8), .b(gate431inter7), .O(gate431inter9));
  nand2 gate1453(.a(s_129), .b(gate431inter3), .O(gate431inter10));
  nor2  gate1454(.a(gate431inter10), .b(gate431inter9), .O(gate431inter11));
  nor2  gate1455(.a(gate431inter11), .b(gate431inter6), .O(gate431inter12));
  nand2 gate1456(.a(gate431inter12), .b(gate431inter1), .O(G1240));
nand2 gate432( .a(G1054), .b(G1150), .O(G1241) );
nand2 gate433( .a(G8), .b(G1153), .O(G1242) );
nand2 gate434( .a(G1057), .b(G1153), .O(G1243) );
nand2 gate435( .a(G9), .b(G1156), .O(G1244) );

  xor2  gate1121(.a(G1156), .b(G1060), .O(gate436inter0));
  nand2 gate1122(.a(gate436inter0), .b(s_82), .O(gate436inter1));
  and2  gate1123(.a(G1156), .b(G1060), .O(gate436inter2));
  inv1  gate1124(.a(s_82), .O(gate436inter3));
  inv1  gate1125(.a(s_83), .O(gate436inter4));
  nand2 gate1126(.a(gate436inter4), .b(gate436inter3), .O(gate436inter5));
  nor2  gate1127(.a(gate436inter5), .b(gate436inter2), .O(gate436inter6));
  inv1  gate1128(.a(G1060), .O(gate436inter7));
  inv1  gate1129(.a(G1156), .O(gate436inter8));
  nand2 gate1130(.a(gate436inter8), .b(gate436inter7), .O(gate436inter9));
  nand2 gate1131(.a(s_83), .b(gate436inter3), .O(gate436inter10));
  nor2  gate1132(.a(gate436inter10), .b(gate436inter9), .O(gate436inter11));
  nor2  gate1133(.a(gate436inter11), .b(gate436inter6), .O(gate436inter12));
  nand2 gate1134(.a(gate436inter12), .b(gate436inter1), .O(G1245));
nand2 gate437( .a(G10), .b(G1159), .O(G1246) );
nand2 gate438( .a(G1063), .b(G1159), .O(G1247) );
nand2 gate439( .a(G11), .b(G1162), .O(G1248) );
nand2 gate440( .a(G1066), .b(G1162), .O(G1249) );
nand2 gate441( .a(G12), .b(G1165), .O(G1250) );
nand2 gate442( .a(G1069), .b(G1165), .O(G1251) );
nand2 gate443( .a(G13), .b(G1168), .O(G1252) );

  xor2  gate953(.a(G1168), .b(G1072), .O(gate444inter0));
  nand2 gate954(.a(gate444inter0), .b(s_58), .O(gate444inter1));
  and2  gate955(.a(G1168), .b(G1072), .O(gate444inter2));
  inv1  gate956(.a(s_58), .O(gate444inter3));
  inv1  gate957(.a(s_59), .O(gate444inter4));
  nand2 gate958(.a(gate444inter4), .b(gate444inter3), .O(gate444inter5));
  nor2  gate959(.a(gate444inter5), .b(gate444inter2), .O(gate444inter6));
  inv1  gate960(.a(G1072), .O(gate444inter7));
  inv1  gate961(.a(G1168), .O(gate444inter8));
  nand2 gate962(.a(gate444inter8), .b(gate444inter7), .O(gate444inter9));
  nand2 gate963(.a(s_59), .b(gate444inter3), .O(gate444inter10));
  nor2  gate964(.a(gate444inter10), .b(gate444inter9), .O(gate444inter11));
  nor2  gate965(.a(gate444inter11), .b(gate444inter6), .O(gate444inter12));
  nand2 gate966(.a(gate444inter12), .b(gate444inter1), .O(G1253));
nand2 gate445( .a(G14), .b(G1171), .O(G1254) );
nand2 gate446( .a(G1075), .b(G1171), .O(G1255) );
nand2 gate447( .a(G15), .b(G1174), .O(G1256) );
nand2 gate448( .a(G1078), .b(G1174), .O(G1257) );
nand2 gate449( .a(G16), .b(G1177), .O(G1258) );
nand2 gate450( .a(G1081), .b(G1177), .O(G1259) );

  xor2  gate1009(.a(G1180), .b(G17), .O(gate451inter0));
  nand2 gate1010(.a(gate451inter0), .b(s_66), .O(gate451inter1));
  and2  gate1011(.a(G1180), .b(G17), .O(gate451inter2));
  inv1  gate1012(.a(s_66), .O(gate451inter3));
  inv1  gate1013(.a(s_67), .O(gate451inter4));
  nand2 gate1014(.a(gate451inter4), .b(gate451inter3), .O(gate451inter5));
  nor2  gate1015(.a(gate451inter5), .b(gate451inter2), .O(gate451inter6));
  inv1  gate1016(.a(G17), .O(gate451inter7));
  inv1  gate1017(.a(G1180), .O(gate451inter8));
  nand2 gate1018(.a(gate451inter8), .b(gate451inter7), .O(gate451inter9));
  nand2 gate1019(.a(s_67), .b(gate451inter3), .O(gate451inter10));
  nor2  gate1020(.a(gate451inter10), .b(gate451inter9), .O(gate451inter11));
  nor2  gate1021(.a(gate451inter11), .b(gate451inter6), .O(gate451inter12));
  nand2 gate1022(.a(gate451inter12), .b(gate451inter1), .O(G1260));

  xor2  gate1051(.a(G1180), .b(G1084), .O(gate452inter0));
  nand2 gate1052(.a(gate452inter0), .b(s_72), .O(gate452inter1));
  and2  gate1053(.a(G1180), .b(G1084), .O(gate452inter2));
  inv1  gate1054(.a(s_72), .O(gate452inter3));
  inv1  gate1055(.a(s_73), .O(gate452inter4));
  nand2 gate1056(.a(gate452inter4), .b(gate452inter3), .O(gate452inter5));
  nor2  gate1057(.a(gate452inter5), .b(gate452inter2), .O(gate452inter6));
  inv1  gate1058(.a(G1084), .O(gate452inter7));
  inv1  gate1059(.a(G1180), .O(gate452inter8));
  nand2 gate1060(.a(gate452inter8), .b(gate452inter7), .O(gate452inter9));
  nand2 gate1061(.a(s_73), .b(gate452inter3), .O(gate452inter10));
  nor2  gate1062(.a(gate452inter10), .b(gate452inter9), .O(gate452inter11));
  nor2  gate1063(.a(gate452inter11), .b(gate452inter6), .O(gate452inter12));
  nand2 gate1064(.a(gate452inter12), .b(gate452inter1), .O(G1261));
nand2 gate453( .a(G18), .b(G1183), .O(G1262) );
nand2 gate454( .a(G1087), .b(G1183), .O(G1263) );
nand2 gate455( .a(G19), .b(G1186), .O(G1264) );
nand2 gate456( .a(G1090), .b(G1186), .O(G1265) );
nand2 gate457( .a(G20), .b(G1189), .O(G1266) );
nand2 gate458( .a(G1093), .b(G1189), .O(G1267) );
nand2 gate459( .a(G21), .b(G1192), .O(G1268) );

  xor2  gate1471(.a(G1192), .b(G1096), .O(gate460inter0));
  nand2 gate1472(.a(gate460inter0), .b(s_132), .O(gate460inter1));
  and2  gate1473(.a(G1192), .b(G1096), .O(gate460inter2));
  inv1  gate1474(.a(s_132), .O(gate460inter3));
  inv1  gate1475(.a(s_133), .O(gate460inter4));
  nand2 gate1476(.a(gate460inter4), .b(gate460inter3), .O(gate460inter5));
  nor2  gate1477(.a(gate460inter5), .b(gate460inter2), .O(gate460inter6));
  inv1  gate1478(.a(G1096), .O(gate460inter7));
  inv1  gate1479(.a(G1192), .O(gate460inter8));
  nand2 gate1480(.a(gate460inter8), .b(gate460inter7), .O(gate460inter9));
  nand2 gate1481(.a(s_133), .b(gate460inter3), .O(gate460inter10));
  nor2  gate1482(.a(gate460inter10), .b(gate460inter9), .O(gate460inter11));
  nor2  gate1483(.a(gate460inter11), .b(gate460inter6), .O(gate460inter12));
  nand2 gate1484(.a(gate460inter12), .b(gate460inter1), .O(G1269));
nand2 gate461( .a(G22), .b(G1195), .O(G1270) );
nand2 gate462( .a(G1099), .b(G1195), .O(G1271) );
nand2 gate463( .a(G23), .b(G1198), .O(G1272) );
nand2 gate464( .a(G1102), .b(G1198), .O(G1273) );
nand2 gate465( .a(G24), .b(G1201), .O(G1274) );
nand2 gate466( .a(G1105), .b(G1201), .O(G1275) );
nand2 gate467( .a(G25), .b(G1204), .O(G1276) );
nand2 gate468( .a(G1108), .b(G1204), .O(G1277) );

  xor2  gate743(.a(G1207), .b(G26), .O(gate469inter0));
  nand2 gate744(.a(gate469inter0), .b(s_28), .O(gate469inter1));
  and2  gate745(.a(G1207), .b(G26), .O(gate469inter2));
  inv1  gate746(.a(s_28), .O(gate469inter3));
  inv1  gate747(.a(s_29), .O(gate469inter4));
  nand2 gate748(.a(gate469inter4), .b(gate469inter3), .O(gate469inter5));
  nor2  gate749(.a(gate469inter5), .b(gate469inter2), .O(gate469inter6));
  inv1  gate750(.a(G26), .O(gate469inter7));
  inv1  gate751(.a(G1207), .O(gate469inter8));
  nand2 gate752(.a(gate469inter8), .b(gate469inter7), .O(gate469inter9));
  nand2 gate753(.a(s_29), .b(gate469inter3), .O(gate469inter10));
  nor2  gate754(.a(gate469inter10), .b(gate469inter9), .O(gate469inter11));
  nor2  gate755(.a(gate469inter11), .b(gate469inter6), .O(gate469inter12));
  nand2 gate756(.a(gate469inter12), .b(gate469inter1), .O(G1278));
nand2 gate470( .a(G1111), .b(G1207), .O(G1279) );
nand2 gate471( .a(G27), .b(G1210), .O(G1280) );
nand2 gate472( .a(G1114), .b(G1210), .O(G1281) );
nand2 gate473( .a(G28), .b(G1213), .O(G1282) );

  xor2  gate1597(.a(G1213), .b(G1117), .O(gate474inter0));
  nand2 gate1598(.a(gate474inter0), .b(s_150), .O(gate474inter1));
  and2  gate1599(.a(G1213), .b(G1117), .O(gate474inter2));
  inv1  gate1600(.a(s_150), .O(gate474inter3));
  inv1  gate1601(.a(s_151), .O(gate474inter4));
  nand2 gate1602(.a(gate474inter4), .b(gate474inter3), .O(gate474inter5));
  nor2  gate1603(.a(gate474inter5), .b(gate474inter2), .O(gate474inter6));
  inv1  gate1604(.a(G1117), .O(gate474inter7));
  inv1  gate1605(.a(G1213), .O(gate474inter8));
  nand2 gate1606(.a(gate474inter8), .b(gate474inter7), .O(gate474inter9));
  nand2 gate1607(.a(s_151), .b(gate474inter3), .O(gate474inter10));
  nor2  gate1608(.a(gate474inter10), .b(gate474inter9), .O(gate474inter11));
  nor2  gate1609(.a(gate474inter11), .b(gate474inter6), .O(gate474inter12));
  nand2 gate1610(.a(gate474inter12), .b(gate474inter1), .O(G1283));
nand2 gate475( .a(G29), .b(G1216), .O(G1284) );
nand2 gate476( .a(G1120), .b(G1216), .O(G1285) );

  xor2  gate1891(.a(G1219), .b(G30), .O(gate477inter0));
  nand2 gate1892(.a(gate477inter0), .b(s_192), .O(gate477inter1));
  and2  gate1893(.a(G1219), .b(G30), .O(gate477inter2));
  inv1  gate1894(.a(s_192), .O(gate477inter3));
  inv1  gate1895(.a(s_193), .O(gate477inter4));
  nand2 gate1896(.a(gate477inter4), .b(gate477inter3), .O(gate477inter5));
  nor2  gate1897(.a(gate477inter5), .b(gate477inter2), .O(gate477inter6));
  inv1  gate1898(.a(G30), .O(gate477inter7));
  inv1  gate1899(.a(G1219), .O(gate477inter8));
  nand2 gate1900(.a(gate477inter8), .b(gate477inter7), .O(gate477inter9));
  nand2 gate1901(.a(s_193), .b(gate477inter3), .O(gate477inter10));
  nor2  gate1902(.a(gate477inter10), .b(gate477inter9), .O(gate477inter11));
  nor2  gate1903(.a(gate477inter11), .b(gate477inter6), .O(gate477inter12));
  nand2 gate1904(.a(gate477inter12), .b(gate477inter1), .O(G1286));
nand2 gate478( .a(G1123), .b(G1219), .O(G1287) );
nand2 gate479( .a(G31), .b(G1222), .O(G1288) );
nand2 gate480( .a(G1126), .b(G1222), .O(G1289) );
nand2 gate481( .a(G32), .b(G1225), .O(G1290) );

  xor2  gate1989(.a(G1225), .b(G1129), .O(gate482inter0));
  nand2 gate1990(.a(gate482inter0), .b(s_206), .O(gate482inter1));
  and2  gate1991(.a(G1225), .b(G1129), .O(gate482inter2));
  inv1  gate1992(.a(s_206), .O(gate482inter3));
  inv1  gate1993(.a(s_207), .O(gate482inter4));
  nand2 gate1994(.a(gate482inter4), .b(gate482inter3), .O(gate482inter5));
  nor2  gate1995(.a(gate482inter5), .b(gate482inter2), .O(gate482inter6));
  inv1  gate1996(.a(G1129), .O(gate482inter7));
  inv1  gate1997(.a(G1225), .O(gate482inter8));
  nand2 gate1998(.a(gate482inter8), .b(gate482inter7), .O(gate482inter9));
  nand2 gate1999(.a(s_207), .b(gate482inter3), .O(gate482inter10));
  nor2  gate2000(.a(gate482inter10), .b(gate482inter9), .O(gate482inter11));
  nor2  gate2001(.a(gate482inter11), .b(gate482inter6), .O(gate482inter12));
  nand2 gate2002(.a(gate482inter12), .b(gate482inter1), .O(G1291));
nand2 gate483( .a(G1228), .b(G1229), .O(G1292) );
nand2 gate484( .a(G1230), .b(G1231), .O(G1293) );
nand2 gate485( .a(G1232), .b(G1233), .O(G1294) );
nand2 gate486( .a(G1234), .b(G1235), .O(G1295) );
nand2 gate487( .a(G1236), .b(G1237), .O(G1296) );

  xor2  gate897(.a(G1239), .b(G1238), .O(gate488inter0));
  nand2 gate898(.a(gate488inter0), .b(s_50), .O(gate488inter1));
  and2  gate899(.a(G1239), .b(G1238), .O(gate488inter2));
  inv1  gate900(.a(s_50), .O(gate488inter3));
  inv1  gate901(.a(s_51), .O(gate488inter4));
  nand2 gate902(.a(gate488inter4), .b(gate488inter3), .O(gate488inter5));
  nor2  gate903(.a(gate488inter5), .b(gate488inter2), .O(gate488inter6));
  inv1  gate904(.a(G1238), .O(gate488inter7));
  inv1  gate905(.a(G1239), .O(gate488inter8));
  nand2 gate906(.a(gate488inter8), .b(gate488inter7), .O(gate488inter9));
  nand2 gate907(.a(s_51), .b(gate488inter3), .O(gate488inter10));
  nor2  gate908(.a(gate488inter10), .b(gate488inter9), .O(gate488inter11));
  nor2  gate909(.a(gate488inter11), .b(gate488inter6), .O(gate488inter12));
  nand2 gate910(.a(gate488inter12), .b(gate488inter1), .O(G1297));
nand2 gate489( .a(G1240), .b(G1241), .O(G1298) );
nand2 gate490( .a(G1242), .b(G1243), .O(G1299) );

  xor2  gate1163(.a(G1245), .b(G1244), .O(gate491inter0));
  nand2 gate1164(.a(gate491inter0), .b(s_88), .O(gate491inter1));
  and2  gate1165(.a(G1245), .b(G1244), .O(gate491inter2));
  inv1  gate1166(.a(s_88), .O(gate491inter3));
  inv1  gate1167(.a(s_89), .O(gate491inter4));
  nand2 gate1168(.a(gate491inter4), .b(gate491inter3), .O(gate491inter5));
  nor2  gate1169(.a(gate491inter5), .b(gate491inter2), .O(gate491inter6));
  inv1  gate1170(.a(G1244), .O(gate491inter7));
  inv1  gate1171(.a(G1245), .O(gate491inter8));
  nand2 gate1172(.a(gate491inter8), .b(gate491inter7), .O(gate491inter9));
  nand2 gate1173(.a(s_89), .b(gate491inter3), .O(gate491inter10));
  nor2  gate1174(.a(gate491inter10), .b(gate491inter9), .O(gate491inter11));
  nor2  gate1175(.a(gate491inter11), .b(gate491inter6), .O(gate491inter12));
  nand2 gate1176(.a(gate491inter12), .b(gate491inter1), .O(G1300));

  xor2  gate1219(.a(G1247), .b(G1246), .O(gate492inter0));
  nand2 gate1220(.a(gate492inter0), .b(s_96), .O(gate492inter1));
  and2  gate1221(.a(G1247), .b(G1246), .O(gate492inter2));
  inv1  gate1222(.a(s_96), .O(gate492inter3));
  inv1  gate1223(.a(s_97), .O(gate492inter4));
  nand2 gate1224(.a(gate492inter4), .b(gate492inter3), .O(gate492inter5));
  nor2  gate1225(.a(gate492inter5), .b(gate492inter2), .O(gate492inter6));
  inv1  gate1226(.a(G1246), .O(gate492inter7));
  inv1  gate1227(.a(G1247), .O(gate492inter8));
  nand2 gate1228(.a(gate492inter8), .b(gate492inter7), .O(gate492inter9));
  nand2 gate1229(.a(s_97), .b(gate492inter3), .O(gate492inter10));
  nor2  gate1230(.a(gate492inter10), .b(gate492inter9), .O(gate492inter11));
  nor2  gate1231(.a(gate492inter11), .b(gate492inter6), .O(gate492inter12));
  nand2 gate1232(.a(gate492inter12), .b(gate492inter1), .O(G1301));

  xor2  gate1737(.a(G1249), .b(G1248), .O(gate493inter0));
  nand2 gate1738(.a(gate493inter0), .b(s_170), .O(gate493inter1));
  and2  gate1739(.a(G1249), .b(G1248), .O(gate493inter2));
  inv1  gate1740(.a(s_170), .O(gate493inter3));
  inv1  gate1741(.a(s_171), .O(gate493inter4));
  nand2 gate1742(.a(gate493inter4), .b(gate493inter3), .O(gate493inter5));
  nor2  gate1743(.a(gate493inter5), .b(gate493inter2), .O(gate493inter6));
  inv1  gate1744(.a(G1248), .O(gate493inter7));
  inv1  gate1745(.a(G1249), .O(gate493inter8));
  nand2 gate1746(.a(gate493inter8), .b(gate493inter7), .O(gate493inter9));
  nand2 gate1747(.a(s_171), .b(gate493inter3), .O(gate493inter10));
  nor2  gate1748(.a(gate493inter10), .b(gate493inter9), .O(gate493inter11));
  nor2  gate1749(.a(gate493inter11), .b(gate493inter6), .O(gate493inter12));
  nand2 gate1750(.a(gate493inter12), .b(gate493inter1), .O(G1302));
nand2 gate494( .a(G1250), .b(G1251), .O(G1303) );
nand2 gate495( .a(G1252), .b(G1253), .O(G1304) );
nand2 gate496( .a(G1254), .b(G1255), .O(G1305) );
nand2 gate497( .a(G1256), .b(G1257), .O(G1306) );

  xor2  gate827(.a(G1259), .b(G1258), .O(gate498inter0));
  nand2 gate828(.a(gate498inter0), .b(s_40), .O(gate498inter1));
  and2  gate829(.a(G1259), .b(G1258), .O(gate498inter2));
  inv1  gate830(.a(s_40), .O(gate498inter3));
  inv1  gate831(.a(s_41), .O(gate498inter4));
  nand2 gate832(.a(gate498inter4), .b(gate498inter3), .O(gate498inter5));
  nor2  gate833(.a(gate498inter5), .b(gate498inter2), .O(gate498inter6));
  inv1  gate834(.a(G1258), .O(gate498inter7));
  inv1  gate835(.a(G1259), .O(gate498inter8));
  nand2 gate836(.a(gate498inter8), .b(gate498inter7), .O(gate498inter9));
  nand2 gate837(.a(s_41), .b(gate498inter3), .O(gate498inter10));
  nor2  gate838(.a(gate498inter10), .b(gate498inter9), .O(gate498inter11));
  nor2  gate839(.a(gate498inter11), .b(gate498inter6), .O(gate498inter12));
  nand2 gate840(.a(gate498inter12), .b(gate498inter1), .O(G1307));
nand2 gate499( .a(G1260), .b(G1261), .O(G1308) );
nand2 gate500( .a(G1262), .b(G1263), .O(G1309) );
nand2 gate501( .a(G1264), .b(G1265), .O(G1310) );
nand2 gate502( .a(G1266), .b(G1267), .O(G1311) );
nand2 gate503( .a(G1268), .b(G1269), .O(G1312) );

  xor2  gate1639(.a(G1271), .b(G1270), .O(gate504inter0));
  nand2 gate1640(.a(gate504inter0), .b(s_156), .O(gate504inter1));
  and2  gate1641(.a(G1271), .b(G1270), .O(gate504inter2));
  inv1  gate1642(.a(s_156), .O(gate504inter3));
  inv1  gate1643(.a(s_157), .O(gate504inter4));
  nand2 gate1644(.a(gate504inter4), .b(gate504inter3), .O(gate504inter5));
  nor2  gate1645(.a(gate504inter5), .b(gate504inter2), .O(gate504inter6));
  inv1  gate1646(.a(G1270), .O(gate504inter7));
  inv1  gate1647(.a(G1271), .O(gate504inter8));
  nand2 gate1648(.a(gate504inter8), .b(gate504inter7), .O(gate504inter9));
  nand2 gate1649(.a(s_157), .b(gate504inter3), .O(gate504inter10));
  nor2  gate1650(.a(gate504inter10), .b(gate504inter9), .O(gate504inter11));
  nor2  gate1651(.a(gate504inter11), .b(gate504inter6), .O(gate504inter12));
  nand2 gate1652(.a(gate504inter12), .b(gate504inter1), .O(G1313));

  xor2  gate841(.a(G1273), .b(G1272), .O(gate505inter0));
  nand2 gate842(.a(gate505inter0), .b(s_42), .O(gate505inter1));
  and2  gate843(.a(G1273), .b(G1272), .O(gate505inter2));
  inv1  gate844(.a(s_42), .O(gate505inter3));
  inv1  gate845(.a(s_43), .O(gate505inter4));
  nand2 gate846(.a(gate505inter4), .b(gate505inter3), .O(gate505inter5));
  nor2  gate847(.a(gate505inter5), .b(gate505inter2), .O(gate505inter6));
  inv1  gate848(.a(G1272), .O(gate505inter7));
  inv1  gate849(.a(G1273), .O(gate505inter8));
  nand2 gate850(.a(gate505inter8), .b(gate505inter7), .O(gate505inter9));
  nand2 gate851(.a(s_43), .b(gate505inter3), .O(gate505inter10));
  nor2  gate852(.a(gate505inter10), .b(gate505inter9), .O(gate505inter11));
  nor2  gate853(.a(gate505inter11), .b(gate505inter6), .O(gate505inter12));
  nand2 gate854(.a(gate505inter12), .b(gate505inter1), .O(G1314));
nand2 gate506( .a(G1274), .b(G1275), .O(G1315) );

  xor2  gate967(.a(G1277), .b(G1276), .O(gate507inter0));
  nand2 gate968(.a(gate507inter0), .b(s_60), .O(gate507inter1));
  and2  gate969(.a(G1277), .b(G1276), .O(gate507inter2));
  inv1  gate970(.a(s_60), .O(gate507inter3));
  inv1  gate971(.a(s_61), .O(gate507inter4));
  nand2 gate972(.a(gate507inter4), .b(gate507inter3), .O(gate507inter5));
  nor2  gate973(.a(gate507inter5), .b(gate507inter2), .O(gate507inter6));
  inv1  gate974(.a(G1276), .O(gate507inter7));
  inv1  gate975(.a(G1277), .O(gate507inter8));
  nand2 gate976(.a(gate507inter8), .b(gate507inter7), .O(gate507inter9));
  nand2 gate977(.a(s_61), .b(gate507inter3), .O(gate507inter10));
  nor2  gate978(.a(gate507inter10), .b(gate507inter9), .O(gate507inter11));
  nor2  gate979(.a(gate507inter11), .b(gate507inter6), .O(gate507inter12));
  nand2 gate980(.a(gate507inter12), .b(gate507inter1), .O(G1316));

  xor2  gate1457(.a(G1279), .b(G1278), .O(gate508inter0));
  nand2 gate1458(.a(gate508inter0), .b(s_130), .O(gate508inter1));
  and2  gate1459(.a(G1279), .b(G1278), .O(gate508inter2));
  inv1  gate1460(.a(s_130), .O(gate508inter3));
  inv1  gate1461(.a(s_131), .O(gate508inter4));
  nand2 gate1462(.a(gate508inter4), .b(gate508inter3), .O(gate508inter5));
  nor2  gate1463(.a(gate508inter5), .b(gate508inter2), .O(gate508inter6));
  inv1  gate1464(.a(G1278), .O(gate508inter7));
  inv1  gate1465(.a(G1279), .O(gate508inter8));
  nand2 gate1466(.a(gate508inter8), .b(gate508inter7), .O(gate508inter9));
  nand2 gate1467(.a(s_131), .b(gate508inter3), .O(gate508inter10));
  nor2  gate1468(.a(gate508inter10), .b(gate508inter9), .O(gate508inter11));
  nor2  gate1469(.a(gate508inter11), .b(gate508inter6), .O(gate508inter12));
  nand2 gate1470(.a(gate508inter12), .b(gate508inter1), .O(G1317));
nand2 gate509( .a(G1280), .b(G1281), .O(G1318) );
nand2 gate510( .a(G1282), .b(G1283), .O(G1319) );
nand2 gate511( .a(G1284), .b(G1285), .O(G1320) );
nand2 gate512( .a(G1286), .b(G1287), .O(G1321) );

  xor2  gate547(.a(G1289), .b(G1288), .O(gate513inter0));
  nand2 gate548(.a(gate513inter0), .b(s_0), .O(gate513inter1));
  and2  gate549(.a(G1289), .b(G1288), .O(gate513inter2));
  inv1  gate550(.a(s_0), .O(gate513inter3));
  inv1  gate551(.a(s_1), .O(gate513inter4));
  nand2 gate552(.a(gate513inter4), .b(gate513inter3), .O(gate513inter5));
  nor2  gate553(.a(gate513inter5), .b(gate513inter2), .O(gate513inter6));
  inv1  gate554(.a(G1288), .O(gate513inter7));
  inv1  gate555(.a(G1289), .O(gate513inter8));
  nand2 gate556(.a(gate513inter8), .b(gate513inter7), .O(gate513inter9));
  nand2 gate557(.a(s_1), .b(gate513inter3), .O(gate513inter10));
  nor2  gate558(.a(gate513inter10), .b(gate513inter9), .O(gate513inter11));
  nor2  gate559(.a(gate513inter11), .b(gate513inter6), .O(gate513inter12));
  nand2 gate560(.a(gate513inter12), .b(gate513inter1), .O(G1322));
nand2 gate514( .a(G1290), .b(G1291), .O(G1323) );
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule