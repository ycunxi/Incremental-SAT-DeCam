module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);

input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;//RE__PI;

input s_0,s_1;//RE__ALLOW(00,01,10,11);
input s_2,s_3;//RE__ALLOW(00,01,10,11);
input s_4,s_5;//RE__ALLOW(00,01,10,11);
input s_6,s_7;//RE__ALLOW(00,01,10,11);
input s_8,s_9;//RE__ALLOW(00,01,10,11);
input s_10,s_11;//RE__ALLOW(00,01,10,11);
input s_12,s_13;//RE__ALLOW(00,01,10,11);
input s_14,s_15;//RE__ALLOW(00,01,10,11);
input s_16,s_17;//RE__ALLOW(00,01,10,11);
input s_18,s_19;//RE__ALLOW(00,01,10,11);
input s_20,s_21;//RE__ALLOW(00,01,10,11);
input s_22,s_23;//RE__ALLOW(00,01,10,11);
input s_24,s_25;//RE__ALLOW(00,01,10,11);
input s_26,s_27;//RE__ALLOW(00,01,10,11);
input s_28,s_29;//RE__ALLOW(00,01,10,11);
input s_30,s_31;//RE__ALLOW(00,01,10,11);
input s_32,s_33;//RE__ALLOW(00,01,10,11);
input s_34,s_35;//RE__ALLOW(00,01,10,11);
input s_36,s_37;//RE__ALLOW(00,01,10,11);
input s_38,s_39;//RE__ALLOW(00,01,10,11);
input s_40,s_41;//RE__ALLOW(00,01,10,11);
input s_42,s_43;//RE__ALLOW(00,01,10,11);
input s_44,s_45;//RE__ALLOW(00,01,10,11);
input s_46,s_47;//RE__ALLOW(00,01,10,11);
input s_48,s_49;//RE__ALLOW(00,01,10,11);
input s_50,s_51;//RE__ALLOW(00,01,10,11);
input s_52,s_53;//RE__ALLOW(00,01,10,11);
input s_54,s_55;//RE__ALLOW(00,01,10,11);
input s_56,s_57;//RE__ALLOW(00,01,10,11);
input s_58,s_59;//RE__ALLOW(00,01,10,11);
input s_60,s_61;//RE__ALLOW(00,01,10,11);
input s_62,s_63;//RE__ALLOW(00,01,10,11);
input s_64,s_65;//RE__ALLOW(00,01,10,11);
input s_66,s_67;//RE__ALLOW(00,01,10,11);
input s_68,s_69;//RE__ALLOW(00,01,10,11);
input s_70,s_71;//RE__ALLOW(00,01,10,11);
input s_72,s_73;//RE__ALLOW(00,01,10,11);
input s_74,s_75;//RE__ALLOW(00,01,10,11);
input s_76,s_77;//RE__ALLOW(00,01,10,11);
input s_78,s_79;//RE__ALLOW(00,01,10,11);
input s_80,s_81;//RE__ALLOW(00,01,10,11);
input s_82,s_83;//RE__ALLOW(00,01,10,11);
input s_84,s_85;//RE__ALLOW(00,01,10,11);
input s_86,s_87;//RE__ALLOW(00,01,10,11);
input s_88,s_89;//RE__ALLOW(00,01,10,11);
input s_90,s_91;//RE__ALLOW(00,01,10,11);
input s_92,s_93;//RE__ALLOW(00,01,10,11);
input s_94,s_95;//RE__ALLOW(00,01,10,11);
input s_96,s_97;//RE__ALLOW(00,01,10,11);
input s_98,s_99;//RE__ALLOW(00,01,10,11);
input s_100,s_101;//RE__ALLOW(00,01,10,11);
input s_102,s_103;//RE__ALLOW(00,01,10,11);
input s_104,s_105;//RE__ALLOW(00,01,10,11);
input s_106,s_107;//RE__ALLOW(00,01,10,11);
input s_108,s_109;//RE__ALLOW(00,01,10,11);
input s_110,s_111;//RE__ALLOW(00,01,10,11);
input s_112,s_113;//RE__ALLOW(00,01,10,11);
input s_114,s_115;//RE__ALLOW(00,01,10,11);
input s_116,s_117;//RE__ALLOW(00,01,10,11);
input s_118,s_119;//RE__ALLOW(00,01,10,11);
input s_120,s_121;//RE__ALLOW(00,01,10,11);
input s_122,s_123;//RE__ALLOW(00,01,10,11);
input s_124,s_125;//RE__ALLOW(00,01,10,11);
input s_126,s_127;//RE__ALLOW(00,01,10,11);
input s_128,s_129;//RE__ALLOW(00,01,10,11);
input s_130,s_131;//RE__ALLOW(00,01,10,11);
input s_132,s_133;//RE__ALLOW(00,01,10,11);
input s_134,s_135;//RE__ALLOW(00,01,10,11);
input s_136,s_137;//RE__ALLOW(00,01,10,11);
input s_138,s_139;//RE__ALLOW(00,01,10,11);
input s_140,s_141;//RE__ALLOW(00,01,10,11);
input s_142,s_143;//RE__ALLOW(00,01,10,11);
input s_144,s_145;//RE__ALLOW(00,01,10,11);
input s_146,s_147;//RE__ALLOW(00,01,10,11);
input s_148,s_149;//RE__ALLOW(00,01,10,11);
input s_150,s_151;//RE__ALLOW(00,01,10,11);
input s_152,s_153;//RE__ALLOW(00,01,10,11);
input s_154,s_155;//RE__ALLOW(00,01,10,11);
input s_156,s_157;//RE__ALLOW(00,01,10,11);
input s_158,s_159;//RE__ALLOW(00,01,10,11);
input s_160,s_161;//RE__ALLOW(00,01,10,11);
input s_162,s_163;//RE__ALLOW(00,01,10,11);
input s_164,s_165;//RE__ALLOW(00,01,10,11);
input s_166,s_167;//RE__ALLOW(00,01,10,11);
input s_168,s_169;//RE__ALLOW(00,01,10,11);
input s_170,s_171;//RE__ALLOW(00,01,10,11);
input s_172,s_173;//RE__ALLOW(00,01,10,11);
input s_174,s_175;//RE__ALLOW(00,01,10,11);
input s_176,s_177;//RE__ALLOW(00,01,10,11);
input s_178,s_179;//RE__ALLOW(00,01,10,11);
input s_180,s_181;//RE__ALLOW(00,01,10,11);
input s_182,s_183;//RE__ALLOW(00,01,10,11);
input s_184,s_185;//RE__ALLOW(00,01,10,11);
input s_186,s_187;//RE__ALLOW(00,01,10,11);
input s_188,s_189;//RE__ALLOW(00,01,10,11);
input s_190,s_191;//RE__ALLOW(00,01,10,11);
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;

  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate271inter0, gate271inter1, gate271inter2, gate271inter3, gate271inter4, gate271inter5, gate271inter6, gate271inter7, gate271inter8, gate271inter9, gate271inter10, gate271inter11, gate271inter12, gate177inter0, gate177inter1, gate177inter2, gate177inter3, gate177inter4, gate177inter5, gate177inter6, gate177inter7, gate177inter8, gate177inter9, gate177inter10, gate177inter11, gate177inter12, gate160inter0, gate160inter1, gate160inter2, gate160inter3, gate160inter4, gate160inter5, gate160inter6, gate160inter7, gate160inter8, gate160inter9, gate160inter10, gate160inter11, gate160inter12, gate147inter0, gate147inter1, gate147inter2, gate147inter3, gate147inter4, gate147inter5, gate147inter6, gate147inter7, gate147inter8, gate147inter9, gate147inter10, gate147inter11, gate147inter12, gate482inter0, gate482inter1, gate482inter2, gate482inter3, gate482inter4, gate482inter5, gate482inter6, gate482inter7, gate482inter8, gate482inter9, gate482inter10, gate482inter11, gate482inter12, gate200inter0, gate200inter1, gate200inter2, gate200inter3, gate200inter4, gate200inter5, gate200inter6, gate200inter7, gate200inter8, gate200inter9, gate200inter10, gate200inter11, gate200inter12, gate259inter0, gate259inter1, gate259inter2, gate259inter3, gate259inter4, gate259inter5, gate259inter6, gate259inter7, gate259inter8, gate259inter9, gate259inter10, gate259inter11, gate259inter12, gate23inter0, gate23inter1, gate23inter2, gate23inter3, gate23inter4, gate23inter5, gate23inter6, gate23inter7, gate23inter8, gate23inter9, gate23inter10, gate23inter11, gate23inter12, gate463inter0, gate463inter1, gate463inter2, gate463inter3, gate463inter4, gate463inter5, gate463inter6, gate463inter7, gate463inter8, gate463inter9, gate463inter10, gate463inter11, gate463inter12, gate154inter0, gate154inter1, gate154inter2, gate154inter3, gate154inter4, gate154inter5, gate154inter6, gate154inter7, gate154inter8, gate154inter9, gate154inter10, gate154inter11, gate154inter12, gate494inter0, gate494inter1, gate494inter2, gate494inter3, gate494inter4, gate494inter5, gate494inter6, gate494inter7, gate494inter8, gate494inter9, gate494inter10, gate494inter11, gate494inter12, gate285inter0, gate285inter1, gate285inter2, gate285inter3, gate285inter4, gate285inter5, gate285inter6, gate285inter7, gate285inter8, gate285inter9, gate285inter10, gate285inter11, gate285inter12, gate410inter0, gate410inter1, gate410inter2, gate410inter3, gate410inter4, gate410inter5, gate410inter6, gate410inter7, gate410inter8, gate410inter9, gate410inter10, gate410inter11, gate410inter12, gate124inter0, gate124inter1, gate124inter2, gate124inter3, gate124inter4, gate124inter5, gate124inter6, gate124inter7, gate124inter8, gate124inter9, gate124inter10, gate124inter11, gate124inter12, gate220inter0, gate220inter1, gate220inter2, gate220inter3, gate220inter4, gate220inter5, gate220inter6, gate220inter7, gate220inter8, gate220inter9, gate220inter10, gate220inter11, gate220inter12, gate393inter0, gate393inter1, gate393inter2, gate393inter3, gate393inter4, gate393inter5, gate393inter6, gate393inter7, gate393inter8, gate393inter9, gate393inter10, gate393inter11, gate393inter12, gate508inter0, gate508inter1, gate508inter2, gate508inter3, gate508inter4, gate508inter5, gate508inter6, gate508inter7, gate508inter8, gate508inter9, gate508inter10, gate508inter11, gate508inter12, gate237inter0, gate237inter1, gate237inter2, gate237inter3, gate237inter4, gate237inter5, gate237inter6, gate237inter7, gate237inter8, gate237inter9, gate237inter10, gate237inter11, gate237inter12, gate246inter0, gate246inter1, gate246inter2, gate246inter3, gate246inter4, gate246inter5, gate246inter6, gate246inter7, gate246inter8, gate246inter9, gate246inter10, gate246inter11, gate246inter12, gate198inter0, gate198inter1, gate198inter2, gate198inter3, gate198inter4, gate198inter5, gate198inter6, gate198inter7, gate198inter8, gate198inter9, gate198inter10, gate198inter11, gate198inter12, gate12inter0, gate12inter1, gate12inter2, gate12inter3, gate12inter4, gate12inter5, gate12inter6, gate12inter7, gate12inter8, gate12inter9, gate12inter10, gate12inter11, gate12inter12, gate245inter0, gate245inter1, gate245inter2, gate245inter3, gate245inter4, gate245inter5, gate245inter6, gate245inter7, gate245inter8, gate245inter9, gate245inter10, gate245inter11, gate245inter12, gate507inter0, gate507inter1, gate507inter2, gate507inter3, gate507inter4, gate507inter5, gate507inter6, gate507inter7, gate507inter8, gate507inter9, gate507inter10, gate507inter11, gate507inter12, gate239inter0, gate239inter1, gate239inter2, gate239inter3, gate239inter4, gate239inter5, gate239inter6, gate239inter7, gate239inter8, gate239inter9, gate239inter10, gate239inter11, gate239inter12, gate458inter0, gate458inter1, gate458inter2, gate458inter3, gate458inter4, gate458inter5, gate458inter6, gate458inter7, gate458inter8, gate458inter9, gate458inter10, gate458inter11, gate458inter12, gate35inter0, gate35inter1, gate35inter2, gate35inter3, gate35inter4, gate35inter5, gate35inter6, gate35inter7, gate35inter8, gate35inter9, gate35inter10, gate35inter11, gate35inter12, gate243inter0, gate243inter1, gate243inter2, gate243inter3, gate243inter4, gate243inter5, gate243inter6, gate243inter7, gate243inter8, gate243inter9, gate243inter10, gate243inter11, gate243inter12, gate223inter0, gate223inter1, gate223inter2, gate223inter3, gate223inter4, gate223inter5, gate223inter6, gate223inter7, gate223inter8, gate223inter9, gate223inter10, gate223inter11, gate223inter12, gate483inter0, gate483inter1, gate483inter2, gate483inter3, gate483inter4, gate483inter5, gate483inter6, gate483inter7, gate483inter8, gate483inter9, gate483inter10, gate483inter11, gate483inter12, gate240inter0, gate240inter1, gate240inter2, gate240inter3, gate240inter4, gate240inter5, gate240inter6, gate240inter7, gate240inter8, gate240inter9, gate240inter10, gate240inter11, gate240inter12, gate446inter0, gate446inter1, gate446inter2, gate446inter3, gate446inter4, gate446inter5, gate446inter6, gate446inter7, gate446inter8, gate446inter9, gate446inter10, gate446inter11, gate446inter12, gate162inter0, gate162inter1, gate162inter2, gate162inter3, gate162inter4, gate162inter5, gate162inter6, gate162inter7, gate162inter8, gate162inter9, gate162inter10, gate162inter11, gate162inter12, gate19inter0, gate19inter1, gate19inter2, gate19inter3, gate19inter4, gate19inter5, gate19inter6, gate19inter7, gate19inter8, gate19inter9, gate19inter10, gate19inter11, gate19inter12, gate65inter0, gate65inter1, gate65inter2, gate65inter3, gate65inter4, gate65inter5, gate65inter6, gate65inter7, gate65inter8, gate65inter9, gate65inter10, gate65inter11, gate65inter12, gate195inter0, gate195inter1, gate195inter2, gate195inter3, gate195inter4, gate195inter5, gate195inter6, gate195inter7, gate195inter8, gate195inter9, gate195inter10, gate195inter11, gate195inter12, gate203inter0, gate203inter1, gate203inter2, gate203inter3, gate203inter4, gate203inter5, gate203inter6, gate203inter7, gate203inter8, gate203inter9, gate203inter10, gate203inter11, gate203inter12, gate452inter0, gate452inter1, gate452inter2, gate452inter3, gate452inter4, gate452inter5, gate452inter6, gate452inter7, gate452inter8, gate452inter9, gate452inter10, gate452inter11, gate452inter12, gate205inter0, gate205inter1, gate205inter2, gate205inter3, gate205inter4, gate205inter5, gate205inter6, gate205inter7, gate205inter8, gate205inter9, gate205inter10, gate205inter11, gate205inter12, gate112inter0, gate112inter1, gate112inter2, gate112inter3, gate112inter4, gate112inter5, gate112inter6, gate112inter7, gate112inter8, gate112inter9, gate112inter10, gate112inter11, gate112inter12, gate171inter0, gate171inter1, gate171inter2, gate171inter3, gate171inter4, gate171inter5, gate171inter6, gate171inter7, gate171inter8, gate171inter9, gate171inter10, gate171inter11, gate171inter12, gate164inter0, gate164inter1, gate164inter2, gate164inter3, gate164inter4, gate164inter5, gate164inter6, gate164inter7, gate164inter8, gate164inter9, gate164inter10, gate164inter11, gate164inter12, gate58inter0, gate58inter1, gate58inter2, gate58inter3, gate58inter4, gate58inter5, gate58inter6, gate58inter7, gate58inter8, gate58inter9, gate58inter10, gate58inter11, gate58inter12, gate481inter0, gate481inter1, gate481inter2, gate481inter3, gate481inter4, gate481inter5, gate481inter6, gate481inter7, gate481inter8, gate481inter9, gate481inter10, gate481inter11, gate481inter12, gate73inter0, gate73inter1, gate73inter2, gate73inter3, gate73inter4, gate73inter5, gate73inter6, gate73inter7, gate73inter8, gate73inter9, gate73inter10, gate73inter11, gate73inter12, gate136inter0, gate136inter1, gate136inter2, gate136inter3, gate136inter4, gate136inter5, gate136inter6, gate136inter7, gate136inter8, gate136inter9, gate136inter10, gate136inter11, gate136inter12, gate181inter0, gate181inter1, gate181inter2, gate181inter3, gate181inter4, gate181inter5, gate181inter6, gate181inter7, gate181inter8, gate181inter9, gate181inter10, gate181inter11, gate181inter12, gate395inter0, gate395inter1, gate395inter2, gate395inter3, gate395inter4, gate395inter5, gate395inter6, gate395inter7, gate395inter8, gate395inter9, gate395inter10, gate395inter11, gate395inter12, gate443inter0, gate443inter1, gate443inter2, gate443inter3, gate443inter4, gate443inter5, gate443inter6, gate443inter7, gate443inter8, gate443inter9, gate443inter10, gate443inter11, gate443inter12, gate447inter0, gate447inter1, gate447inter2, gate447inter3, gate447inter4, gate447inter5, gate447inter6, gate447inter7, gate447inter8, gate447inter9, gate447inter10, gate447inter11, gate447inter12, gate79inter0, gate79inter1, gate79inter2, gate79inter3, gate79inter4, gate79inter5, gate79inter6, gate79inter7, gate79inter8, gate79inter9, gate79inter10, gate79inter11, gate79inter12, gate216inter0, gate216inter1, gate216inter2, gate216inter3, gate216inter4, gate216inter5, gate216inter6, gate216inter7, gate216inter8, gate216inter9, gate216inter10, gate216inter11, gate216inter12, gate502inter0, gate502inter1, gate502inter2, gate502inter3, gate502inter4, gate502inter5, gate502inter6, gate502inter7, gate502inter8, gate502inter9, gate502inter10, gate502inter11, gate502inter12, gate262inter0, gate262inter1, gate262inter2, gate262inter3, gate262inter4, gate262inter5, gate262inter6, gate262inter7, gate262inter8, gate262inter9, gate262inter10, gate262inter11, gate262inter12, gate453inter0, gate453inter1, gate453inter2, gate453inter3, gate453inter4, gate453inter5, gate453inter6, gate453inter7, gate453inter8, gate453inter9, gate453inter10, gate453inter11, gate453inter12, gate102inter0, gate102inter1, gate102inter2, gate102inter3, gate102inter4, gate102inter5, gate102inter6, gate102inter7, gate102inter8, gate102inter9, gate102inter10, gate102inter11, gate102inter12, gate293inter0, gate293inter1, gate293inter2, gate293inter3, gate293inter4, gate293inter5, gate293inter6, gate293inter7, gate293inter8, gate293inter9, gate293inter10, gate293inter11, gate293inter12, gate94inter0, gate94inter1, gate94inter2, gate94inter3, gate94inter4, gate94inter5, gate94inter6, gate94inter7, gate94inter8, gate94inter9, gate94inter10, gate94inter11, gate94inter12, gate232inter0, gate232inter1, gate232inter2, gate232inter3, gate232inter4, gate232inter5, gate232inter6, gate232inter7, gate232inter8, gate232inter9, gate232inter10, gate232inter11, gate232inter12, gate430inter0, gate430inter1, gate430inter2, gate430inter3, gate430inter4, gate430inter5, gate430inter6, gate430inter7, gate430inter8, gate430inter9, gate430inter10, gate430inter11, gate430inter12, gate34inter0, gate34inter1, gate34inter2, gate34inter3, gate34inter4, gate34inter5, gate34inter6, gate34inter7, gate34inter8, gate34inter9, gate34inter10, gate34inter11, gate34inter12, gate97inter0, gate97inter1, gate97inter2, gate97inter3, gate97inter4, gate97inter5, gate97inter6, gate97inter7, gate97inter8, gate97inter9, gate97inter10, gate97inter11, gate97inter12, gate49inter0, gate49inter1, gate49inter2, gate49inter3, gate49inter4, gate49inter5, gate49inter6, gate49inter7, gate49inter8, gate49inter9, gate49inter10, gate49inter11, gate49inter12, gate399inter0, gate399inter1, gate399inter2, gate399inter3, gate399inter4, gate399inter5, gate399inter6, gate399inter7, gate399inter8, gate399inter9, gate399inter10, gate399inter11, gate399inter12, gate148inter0, gate148inter1, gate148inter2, gate148inter3, gate148inter4, gate148inter5, gate148inter6, gate148inter7, gate148inter8, gate148inter9, gate148inter10, gate148inter11, gate148inter12, gate41inter0, gate41inter1, gate41inter2, gate41inter3, gate41inter4, gate41inter5, gate41inter6, gate41inter7, gate41inter8, gate41inter9, gate41inter10, gate41inter11, gate41inter12, gate474inter0, gate474inter1, gate474inter2, gate474inter3, gate474inter4, gate474inter5, gate474inter6, gate474inter7, gate474inter8, gate474inter9, gate474inter10, gate474inter11, gate474inter12, gate224inter0, gate224inter1, gate224inter2, gate224inter3, gate224inter4, gate224inter5, gate224inter6, gate224inter7, gate224inter8, gate224inter9, gate224inter10, gate224inter11, gate224inter12, gate123inter0, gate123inter1, gate123inter2, gate123inter3, gate123inter4, gate123inter5, gate123inter6, gate123inter7, gate123inter8, gate123inter9, gate123inter10, gate123inter11, gate123inter12, gate449inter0, gate449inter1, gate449inter2, gate449inter3, gate449inter4, gate449inter5, gate449inter6, gate449inter7, gate449inter8, gate449inter9, gate449inter10, gate449inter11, gate449inter12, gate33inter0, gate33inter1, gate33inter2, gate33inter3, gate33inter4, gate33inter5, gate33inter6, gate33inter7, gate33inter8, gate33inter9, gate33inter10, gate33inter11, gate33inter12, gate120inter0, gate120inter1, gate120inter2, gate120inter3, gate120inter4, gate120inter5, gate120inter6, gate120inter7, gate120inter8, gate120inter9, gate120inter10, gate120inter11, gate120inter12, gate392inter0, gate392inter1, gate392inter2, gate392inter3, gate392inter4, gate392inter5, gate392inter6, gate392inter7, gate392inter8, gate392inter9, gate392inter10, gate392inter11, gate392inter12, gate153inter0, gate153inter1, gate153inter2, gate153inter3, gate153inter4, gate153inter5, gate153inter6, gate153inter7, gate153inter8, gate153inter9, gate153inter10, gate153inter11, gate153inter12, gate131inter0, gate131inter1, gate131inter2, gate131inter3, gate131inter4, gate131inter5, gate131inter6, gate131inter7, gate131inter8, gate131inter9, gate131inter10, gate131inter11, gate131inter12, gate501inter0, gate501inter1, gate501inter2, gate501inter3, gate501inter4, gate501inter5, gate501inter6, gate501inter7, gate501inter8, gate501inter9, gate501inter10, gate501inter11, gate501inter12, gate21inter0, gate21inter1, gate21inter2, gate21inter3, gate21inter4, gate21inter5, gate21inter6, gate21inter7, gate21inter8, gate21inter9, gate21inter10, gate21inter11, gate21inter12, gate255inter0, gate255inter1, gate255inter2, gate255inter3, gate255inter4, gate255inter5, gate255inter6, gate255inter7, gate255inter8, gate255inter9, gate255inter10, gate255inter11, gate255inter12, gate506inter0, gate506inter1, gate506inter2, gate506inter3, gate506inter4, gate506inter5, gate506inter6, gate506inter7, gate506inter8, gate506inter9, gate506inter10, gate506inter11, gate506inter12, gate283inter0, gate283inter1, gate283inter2, gate283inter3, gate283inter4, gate283inter5, gate283inter6, gate283inter7, gate283inter8, gate283inter9, gate283inter10, gate283inter11, gate283inter12, gate142inter0, gate142inter1, gate142inter2, gate142inter3, gate142inter4, gate142inter5, gate142inter6, gate142inter7, gate142inter8, gate142inter9, gate142inter10, gate142inter11, gate142inter12, gate37inter0, gate37inter1, gate37inter2, gate37inter3, gate37inter4, gate37inter5, gate37inter6, gate37inter7, gate37inter8, gate37inter9, gate37inter10, gate37inter11, gate37inter12, gate183inter0, gate183inter1, gate183inter2, gate183inter3, gate183inter4, gate183inter5, gate183inter6, gate183inter7, gate183inter8, gate183inter9, gate183inter10, gate183inter11, gate183inter12, gate74inter0, gate74inter1, gate74inter2, gate74inter3, gate74inter4, gate74inter5, gate74inter6, gate74inter7, gate74inter8, gate74inter9, gate74inter10, gate74inter11, gate74inter12, gate244inter0, gate244inter1, gate244inter2, gate244inter3, gate244inter4, gate244inter5, gate244inter6, gate244inter7, gate244inter8, gate244inter9, gate244inter10, gate244inter11, gate244inter12, gate57inter0, gate57inter1, gate57inter2, gate57inter3, gate57inter4, gate57inter5, gate57inter6, gate57inter7, gate57inter8, gate57inter9, gate57inter10, gate57inter11, gate57inter12, gate150inter0, gate150inter1, gate150inter2, gate150inter3, gate150inter4, gate150inter5, gate150inter6, gate150inter7, gate150inter8, gate150inter9, gate150inter10, gate150inter11, gate150inter12, gate420inter0, gate420inter1, gate420inter2, gate420inter3, gate420inter4, gate420inter5, gate420inter6, gate420inter7, gate420inter8, gate420inter9, gate420inter10, gate420inter11, gate420inter12, gate468inter0, gate468inter1, gate468inter2, gate468inter3, gate468inter4, gate468inter5, gate468inter6, gate468inter7, gate468inter8, gate468inter9, gate468inter10, gate468inter11, gate468inter12, gate432inter0, gate432inter1, gate432inter2, gate432inter3, gate432inter4, gate432inter5, gate432inter6, gate432inter7, gate432inter8, gate432inter9, gate432inter10, gate432inter11, gate432inter12, gate466inter0, gate466inter1, gate466inter2, gate466inter3, gate466inter4, gate466inter5, gate466inter6, gate466inter7, gate466inter8, gate466inter9, gate466inter10, gate466inter11, gate466inter12, gate173inter0, gate173inter1, gate173inter2, gate173inter3, gate173inter4, gate173inter5, gate173inter6, gate173inter7, gate173inter8, gate173inter9, gate173inter10, gate173inter11, gate173inter12, gate122inter0, gate122inter1, gate122inter2, gate122inter3, gate122inter4, gate122inter5, gate122inter6, gate122inter7, gate122inter8, gate122inter9, gate122inter10, gate122inter11, gate122inter12, gate107inter0, gate107inter1, gate107inter2, gate107inter3, gate107inter4, gate107inter5, gate107inter6, gate107inter7, gate107inter8, gate107inter9, gate107inter10, gate107inter11, gate107inter12, gate67inter0, gate67inter1, gate67inter2, gate67inter3, gate67inter4, gate67inter5, gate67inter6, gate67inter7, gate67inter8, gate67inter9, gate67inter10, gate67inter11, gate67inter12, gate419inter0, gate419inter1, gate419inter2, gate419inter3, gate419inter4, gate419inter5, gate419inter6, gate419inter7, gate419inter8, gate419inter9, gate419inter10, gate419inter11, gate419inter12, gate145inter0, gate145inter1, gate145inter2, gate145inter3, gate145inter4, gate145inter5, gate145inter6, gate145inter7, gate145inter8, gate145inter9, gate145inter10, gate145inter11, gate145inter12;



and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );
nand2 gate9( .a(G1), .b(G2), .O(G266) );
nand2 gate10( .a(G3), .b(G4), .O(G269) );
nand2 gate11( .a(G5), .b(G6), .O(G272) );

  xor2  gate827(.a(G8), .b(G7), .O(gate12inter0));
  nand2 gate828(.a(gate12inter0), .b(s_40), .O(gate12inter1));
  and2  gate829(.a(G8), .b(G7), .O(gate12inter2));
  inv1  gate830(.a(s_40), .O(gate12inter3));
  inv1  gate831(.a(s_41), .O(gate12inter4));
  nand2 gate832(.a(gate12inter4), .b(gate12inter3), .O(gate12inter5));
  nor2  gate833(.a(gate12inter5), .b(gate12inter2), .O(gate12inter6));
  inv1  gate834(.a(G7), .O(gate12inter7));
  inv1  gate835(.a(G8), .O(gate12inter8));
  nand2 gate836(.a(gate12inter8), .b(gate12inter7), .O(gate12inter9));
  nand2 gate837(.a(s_41), .b(gate12inter3), .O(gate12inter10));
  nor2  gate838(.a(gate12inter10), .b(gate12inter9), .O(gate12inter11));
  nor2  gate839(.a(gate12inter11), .b(gate12inter6), .O(gate12inter12));
  nand2 gate840(.a(gate12inter12), .b(gate12inter1), .O(G275));
nand2 gate13( .a(G9), .b(G10), .O(G278) );
nand2 gate14( .a(G11), .b(G12), .O(G281) );
nand2 gate15( .a(G13), .b(G14), .O(G284) );
nand2 gate16( .a(G15), .b(G16), .O(G287) );
nand2 gate17( .a(G17), .b(G18), .O(G290) );
nand2 gate18( .a(G19), .b(G20), .O(G293) );

  xor2  gate995(.a(G22), .b(G21), .O(gate19inter0));
  nand2 gate996(.a(gate19inter0), .b(s_64), .O(gate19inter1));
  and2  gate997(.a(G22), .b(G21), .O(gate19inter2));
  inv1  gate998(.a(s_64), .O(gate19inter3));
  inv1  gate999(.a(s_65), .O(gate19inter4));
  nand2 gate1000(.a(gate19inter4), .b(gate19inter3), .O(gate19inter5));
  nor2  gate1001(.a(gate19inter5), .b(gate19inter2), .O(gate19inter6));
  inv1  gate1002(.a(G21), .O(gate19inter7));
  inv1  gate1003(.a(G22), .O(gate19inter8));
  nand2 gate1004(.a(gate19inter8), .b(gate19inter7), .O(gate19inter9));
  nand2 gate1005(.a(s_65), .b(gate19inter3), .O(gate19inter10));
  nor2  gate1006(.a(gate19inter10), .b(gate19inter9), .O(gate19inter11));
  nor2  gate1007(.a(gate19inter11), .b(gate19inter6), .O(gate19inter12));
  nand2 gate1008(.a(gate19inter12), .b(gate19inter1), .O(G296));
nand2 gate20( .a(G23), .b(G24), .O(G299) );

  xor2  gate1597(.a(G26), .b(G25), .O(gate21inter0));
  nand2 gate1598(.a(gate21inter0), .b(s_150), .O(gate21inter1));
  and2  gate1599(.a(G26), .b(G25), .O(gate21inter2));
  inv1  gate1600(.a(s_150), .O(gate21inter3));
  inv1  gate1601(.a(s_151), .O(gate21inter4));
  nand2 gate1602(.a(gate21inter4), .b(gate21inter3), .O(gate21inter5));
  nor2  gate1603(.a(gate21inter5), .b(gate21inter2), .O(gate21inter6));
  inv1  gate1604(.a(G25), .O(gate21inter7));
  inv1  gate1605(.a(G26), .O(gate21inter8));
  nand2 gate1606(.a(gate21inter8), .b(gate21inter7), .O(gate21inter9));
  nand2 gate1607(.a(s_151), .b(gate21inter3), .O(gate21inter10));
  nor2  gate1608(.a(gate21inter10), .b(gate21inter9), .O(gate21inter11));
  nor2  gate1609(.a(gate21inter11), .b(gate21inter6), .O(gate21inter12));
  nand2 gate1610(.a(gate21inter12), .b(gate21inter1), .O(G302));
nand2 gate22( .a(G27), .b(G28), .O(G305) );

  xor2  gate645(.a(G30), .b(G29), .O(gate23inter0));
  nand2 gate646(.a(gate23inter0), .b(s_14), .O(gate23inter1));
  and2  gate647(.a(G30), .b(G29), .O(gate23inter2));
  inv1  gate648(.a(s_14), .O(gate23inter3));
  inv1  gate649(.a(s_15), .O(gate23inter4));
  nand2 gate650(.a(gate23inter4), .b(gate23inter3), .O(gate23inter5));
  nor2  gate651(.a(gate23inter5), .b(gate23inter2), .O(gate23inter6));
  inv1  gate652(.a(G29), .O(gate23inter7));
  inv1  gate653(.a(G30), .O(gate23inter8));
  nand2 gate654(.a(gate23inter8), .b(gate23inter7), .O(gate23inter9));
  nand2 gate655(.a(s_15), .b(gate23inter3), .O(gate23inter10));
  nor2  gate656(.a(gate23inter10), .b(gate23inter9), .O(gate23inter11));
  nor2  gate657(.a(gate23inter11), .b(gate23inter6), .O(gate23inter12));
  nand2 gate658(.a(gate23inter12), .b(gate23inter1), .O(G308));
nand2 gate24( .a(G31), .b(G32), .O(G311) );
nand2 gate25( .a(G1), .b(G5), .O(G314) );
nand2 gate26( .a(G9), .b(G13), .O(G317) );
nand2 gate27( .a(G2), .b(G6), .O(G320) );
nand2 gate28( .a(G10), .b(G14), .O(G323) );
nand2 gate29( .a(G3), .b(G7), .O(G326) );
nand2 gate30( .a(G11), .b(G15), .O(G329) );
nand2 gate31( .a(G4), .b(G8), .O(G332) );
nand2 gate32( .a(G12), .b(G16), .O(G335) );

  xor2  gate1513(.a(G21), .b(G17), .O(gate33inter0));
  nand2 gate1514(.a(gate33inter0), .b(s_138), .O(gate33inter1));
  and2  gate1515(.a(G21), .b(G17), .O(gate33inter2));
  inv1  gate1516(.a(s_138), .O(gate33inter3));
  inv1  gate1517(.a(s_139), .O(gate33inter4));
  nand2 gate1518(.a(gate33inter4), .b(gate33inter3), .O(gate33inter5));
  nor2  gate1519(.a(gate33inter5), .b(gate33inter2), .O(gate33inter6));
  inv1  gate1520(.a(G17), .O(gate33inter7));
  inv1  gate1521(.a(G21), .O(gate33inter8));
  nand2 gate1522(.a(gate33inter8), .b(gate33inter7), .O(gate33inter9));
  nand2 gate1523(.a(s_139), .b(gate33inter3), .O(gate33inter10));
  nor2  gate1524(.a(gate33inter10), .b(gate33inter9), .O(gate33inter11));
  nor2  gate1525(.a(gate33inter11), .b(gate33inter6), .O(gate33inter12));
  nand2 gate1526(.a(gate33inter12), .b(gate33inter1), .O(G338));

  xor2  gate1373(.a(G29), .b(G25), .O(gate34inter0));
  nand2 gate1374(.a(gate34inter0), .b(s_118), .O(gate34inter1));
  and2  gate1375(.a(G29), .b(G25), .O(gate34inter2));
  inv1  gate1376(.a(s_118), .O(gate34inter3));
  inv1  gate1377(.a(s_119), .O(gate34inter4));
  nand2 gate1378(.a(gate34inter4), .b(gate34inter3), .O(gate34inter5));
  nor2  gate1379(.a(gate34inter5), .b(gate34inter2), .O(gate34inter6));
  inv1  gate1380(.a(G25), .O(gate34inter7));
  inv1  gate1381(.a(G29), .O(gate34inter8));
  nand2 gate1382(.a(gate34inter8), .b(gate34inter7), .O(gate34inter9));
  nand2 gate1383(.a(s_119), .b(gate34inter3), .O(gate34inter10));
  nor2  gate1384(.a(gate34inter10), .b(gate34inter9), .O(gate34inter11));
  nor2  gate1385(.a(gate34inter11), .b(gate34inter6), .O(gate34inter12));
  nand2 gate1386(.a(gate34inter12), .b(gate34inter1), .O(G341));

  xor2  gate897(.a(G22), .b(G18), .O(gate35inter0));
  nand2 gate898(.a(gate35inter0), .b(s_50), .O(gate35inter1));
  and2  gate899(.a(G22), .b(G18), .O(gate35inter2));
  inv1  gate900(.a(s_50), .O(gate35inter3));
  inv1  gate901(.a(s_51), .O(gate35inter4));
  nand2 gate902(.a(gate35inter4), .b(gate35inter3), .O(gate35inter5));
  nor2  gate903(.a(gate35inter5), .b(gate35inter2), .O(gate35inter6));
  inv1  gate904(.a(G18), .O(gate35inter7));
  inv1  gate905(.a(G22), .O(gate35inter8));
  nand2 gate906(.a(gate35inter8), .b(gate35inter7), .O(gate35inter9));
  nand2 gate907(.a(s_51), .b(gate35inter3), .O(gate35inter10));
  nor2  gate908(.a(gate35inter10), .b(gate35inter9), .O(gate35inter11));
  nor2  gate909(.a(gate35inter11), .b(gate35inter6), .O(gate35inter12));
  nand2 gate910(.a(gate35inter12), .b(gate35inter1), .O(G344));
nand2 gate36( .a(G26), .b(G30), .O(G347) );

  xor2  gate1667(.a(G23), .b(G19), .O(gate37inter0));
  nand2 gate1668(.a(gate37inter0), .b(s_160), .O(gate37inter1));
  and2  gate1669(.a(G23), .b(G19), .O(gate37inter2));
  inv1  gate1670(.a(s_160), .O(gate37inter3));
  inv1  gate1671(.a(s_161), .O(gate37inter4));
  nand2 gate1672(.a(gate37inter4), .b(gate37inter3), .O(gate37inter5));
  nor2  gate1673(.a(gate37inter5), .b(gate37inter2), .O(gate37inter6));
  inv1  gate1674(.a(G19), .O(gate37inter7));
  inv1  gate1675(.a(G23), .O(gate37inter8));
  nand2 gate1676(.a(gate37inter8), .b(gate37inter7), .O(gate37inter9));
  nand2 gate1677(.a(s_161), .b(gate37inter3), .O(gate37inter10));
  nor2  gate1678(.a(gate37inter10), .b(gate37inter9), .O(gate37inter11));
  nor2  gate1679(.a(gate37inter11), .b(gate37inter6), .O(gate37inter12));
  nand2 gate1680(.a(gate37inter12), .b(gate37inter1), .O(G350));
nand2 gate38( .a(G27), .b(G31), .O(G353) );
nand2 gate39( .a(G20), .b(G24), .O(G356) );
nand2 gate40( .a(G28), .b(G32), .O(G359) );

  xor2  gate1443(.a(G266), .b(G1), .O(gate41inter0));
  nand2 gate1444(.a(gate41inter0), .b(s_128), .O(gate41inter1));
  and2  gate1445(.a(G266), .b(G1), .O(gate41inter2));
  inv1  gate1446(.a(s_128), .O(gate41inter3));
  inv1  gate1447(.a(s_129), .O(gate41inter4));
  nand2 gate1448(.a(gate41inter4), .b(gate41inter3), .O(gate41inter5));
  nor2  gate1449(.a(gate41inter5), .b(gate41inter2), .O(gate41inter6));
  inv1  gate1450(.a(G1), .O(gate41inter7));
  inv1  gate1451(.a(G266), .O(gate41inter8));
  nand2 gate1452(.a(gate41inter8), .b(gate41inter7), .O(gate41inter9));
  nand2 gate1453(.a(s_129), .b(gate41inter3), .O(gate41inter10));
  nor2  gate1454(.a(gate41inter10), .b(gate41inter9), .O(gate41inter11));
  nor2  gate1455(.a(gate41inter11), .b(gate41inter6), .O(gate41inter12));
  nand2 gate1456(.a(gate41inter12), .b(gate41inter1), .O(G362));
nand2 gate42( .a(G2), .b(G266), .O(G363) );
nand2 gate43( .a(G3), .b(G269), .O(G364) );
nand2 gate44( .a(G4), .b(G269), .O(G365) );
nand2 gate45( .a(G5), .b(G272), .O(G366) );
nand2 gate46( .a(G6), .b(G272), .O(G367) );
nand2 gate47( .a(G7), .b(G275), .O(G368) );
nand2 gate48( .a(G8), .b(G275), .O(G369) );

  xor2  gate1401(.a(G278), .b(G9), .O(gate49inter0));
  nand2 gate1402(.a(gate49inter0), .b(s_122), .O(gate49inter1));
  and2  gate1403(.a(G278), .b(G9), .O(gate49inter2));
  inv1  gate1404(.a(s_122), .O(gate49inter3));
  inv1  gate1405(.a(s_123), .O(gate49inter4));
  nand2 gate1406(.a(gate49inter4), .b(gate49inter3), .O(gate49inter5));
  nor2  gate1407(.a(gate49inter5), .b(gate49inter2), .O(gate49inter6));
  inv1  gate1408(.a(G9), .O(gate49inter7));
  inv1  gate1409(.a(G278), .O(gate49inter8));
  nand2 gate1410(.a(gate49inter8), .b(gate49inter7), .O(gate49inter9));
  nand2 gate1411(.a(s_123), .b(gate49inter3), .O(gate49inter10));
  nor2  gate1412(.a(gate49inter10), .b(gate49inter9), .O(gate49inter11));
  nor2  gate1413(.a(gate49inter11), .b(gate49inter6), .O(gate49inter12));
  nand2 gate1414(.a(gate49inter12), .b(gate49inter1), .O(G370));
nand2 gate50( .a(G10), .b(G278), .O(G371) );
nand2 gate51( .a(G11), .b(G281), .O(G372) );
nand2 gate52( .a(G12), .b(G281), .O(G373) );
nand2 gate53( .a(G13), .b(G284), .O(G374) );
nand2 gate54( .a(G14), .b(G284), .O(G375) );
nand2 gate55( .a(G15), .b(G287), .O(G376) );
nand2 gate56( .a(G16), .b(G287), .O(G377) );

  xor2  gate1723(.a(G290), .b(G17), .O(gate57inter0));
  nand2 gate1724(.a(gate57inter0), .b(s_168), .O(gate57inter1));
  and2  gate1725(.a(G290), .b(G17), .O(gate57inter2));
  inv1  gate1726(.a(s_168), .O(gate57inter3));
  inv1  gate1727(.a(s_169), .O(gate57inter4));
  nand2 gate1728(.a(gate57inter4), .b(gate57inter3), .O(gate57inter5));
  nor2  gate1729(.a(gate57inter5), .b(gate57inter2), .O(gate57inter6));
  inv1  gate1730(.a(G17), .O(gate57inter7));
  inv1  gate1731(.a(G290), .O(gate57inter8));
  nand2 gate1732(.a(gate57inter8), .b(gate57inter7), .O(gate57inter9));
  nand2 gate1733(.a(s_169), .b(gate57inter3), .O(gate57inter10));
  nor2  gate1734(.a(gate57inter10), .b(gate57inter9), .O(gate57inter11));
  nor2  gate1735(.a(gate57inter11), .b(gate57inter6), .O(gate57inter12));
  nand2 gate1736(.a(gate57inter12), .b(gate57inter1), .O(G378));

  xor2  gate1121(.a(G290), .b(G18), .O(gate58inter0));
  nand2 gate1122(.a(gate58inter0), .b(s_82), .O(gate58inter1));
  and2  gate1123(.a(G290), .b(G18), .O(gate58inter2));
  inv1  gate1124(.a(s_82), .O(gate58inter3));
  inv1  gate1125(.a(s_83), .O(gate58inter4));
  nand2 gate1126(.a(gate58inter4), .b(gate58inter3), .O(gate58inter5));
  nor2  gate1127(.a(gate58inter5), .b(gate58inter2), .O(gate58inter6));
  inv1  gate1128(.a(G18), .O(gate58inter7));
  inv1  gate1129(.a(G290), .O(gate58inter8));
  nand2 gate1130(.a(gate58inter8), .b(gate58inter7), .O(gate58inter9));
  nand2 gate1131(.a(s_83), .b(gate58inter3), .O(gate58inter10));
  nor2  gate1132(.a(gate58inter10), .b(gate58inter9), .O(gate58inter11));
  nor2  gate1133(.a(gate58inter11), .b(gate58inter6), .O(gate58inter12));
  nand2 gate1134(.a(gate58inter12), .b(gate58inter1), .O(G379));
nand2 gate59( .a(G19), .b(G293), .O(G380) );
nand2 gate60( .a(G20), .b(G293), .O(G381) );
nand2 gate61( .a(G21), .b(G296), .O(G382) );
nand2 gate62( .a(G22), .b(G296), .O(G383) );
nand2 gate63( .a(G23), .b(G299), .O(G384) );
nand2 gate64( .a(G24), .b(G299), .O(G385) );

  xor2  gate1009(.a(G302), .b(G25), .O(gate65inter0));
  nand2 gate1010(.a(gate65inter0), .b(s_66), .O(gate65inter1));
  and2  gate1011(.a(G302), .b(G25), .O(gate65inter2));
  inv1  gate1012(.a(s_66), .O(gate65inter3));
  inv1  gate1013(.a(s_67), .O(gate65inter4));
  nand2 gate1014(.a(gate65inter4), .b(gate65inter3), .O(gate65inter5));
  nor2  gate1015(.a(gate65inter5), .b(gate65inter2), .O(gate65inter6));
  inv1  gate1016(.a(G25), .O(gate65inter7));
  inv1  gate1017(.a(G302), .O(gate65inter8));
  nand2 gate1018(.a(gate65inter8), .b(gate65inter7), .O(gate65inter9));
  nand2 gate1019(.a(s_67), .b(gate65inter3), .O(gate65inter10));
  nor2  gate1020(.a(gate65inter10), .b(gate65inter9), .O(gate65inter11));
  nor2  gate1021(.a(gate65inter11), .b(gate65inter6), .O(gate65inter12));
  nand2 gate1022(.a(gate65inter12), .b(gate65inter1), .O(G386));
nand2 gate66( .a(G26), .b(G302), .O(G387) );

  xor2  gate1849(.a(G305), .b(G27), .O(gate67inter0));
  nand2 gate1850(.a(gate67inter0), .b(s_186), .O(gate67inter1));
  and2  gate1851(.a(G305), .b(G27), .O(gate67inter2));
  inv1  gate1852(.a(s_186), .O(gate67inter3));
  inv1  gate1853(.a(s_187), .O(gate67inter4));
  nand2 gate1854(.a(gate67inter4), .b(gate67inter3), .O(gate67inter5));
  nor2  gate1855(.a(gate67inter5), .b(gate67inter2), .O(gate67inter6));
  inv1  gate1856(.a(G27), .O(gate67inter7));
  inv1  gate1857(.a(G305), .O(gate67inter8));
  nand2 gate1858(.a(gate67inter8), .b(gate67inter7), .O(gate67inter9));
  nand2 gate1859(.a(s_187), .b(gate67inter3), .O(gate67inter10));
  nor2  gate1860(.a(gate67inter10), .b(gate67inter9), .O(gate67inter11));
  nor2  gate1861(.a(gate67inter11), .b(gate67inter6), .O(gate67inter12));
  nand2 gate1862(.a(gate67inter12), .b(gate67inter1), .O(G388));
nand2 gate68( .a(G28), .b(G305), .O(G389) );
nand2 gate69( .a(G29), .b(G308), .O(G390) );
nand2 gate70( .a(G30), .b(G308), .O(G391) );
nand2 gate71( .a(G31), .b(G311), .O(G392) );
nand2 gate72( .a(G32), .b(G311), .O(G393) );

  xor2  gate1149(.a(G314), .b(G1), .O(gate73inter0));
  nand2 gate1150(.a(gate73inter0), .b(s_86), .O(gate73inter1));
  and2  gate1151(.a(G314), .b(G1), .O(gate73inter2));
  inv1  gate1152(.a(s_86), .O(gate73inter3));
  inv1  gate1153(.a(s_87), .O(gate73inter4));
  nand2 gate1154(.a(gate73inter4), .b(gate73inter3), .O(gate73inter5));
  nor2  gate1155(.a(gate73inter5), .b(gate73inter2), .O(gate73inter6));
  inv1  gate1156(.a(G1), .O(gate73inter7));
  inv1  gate1157(.a(G314), .O(gate73inter8));
  nand2 gate1158(.a(gate73inter8), .b(gate73inter7), .O(gate73inter9));
  nand2 gate1159(.a(s_87), .b(gate73inter3), .O(gate73inter10));
  nor2  gate1160(.a(gate73inter10), .b(gate73inter9), .O(gate73inter11));
  nor2  gate1161(.a(gate73inter11), .b(gate73inter6), .O(gate73inter12));
  nand2 gate1162(.a(gate73inter12), .b(gate73inter1), .O(G394));

  xor2  gate1695(.a(G314), .b(G5), .O(gate74inter0));
  nand2 gate1696(.a(gate74inter0), .b(s_164), .O(gate74inter1));
  and2  gate1697(.a(G314), .b(G5), .O(gate74inter2));
  inv1  gate1698(.a(s_164), .O(gate74inter3));
  inv1  gate1699(.a(s_165), .O(gate74inter4));
  nand2 gate1700(.a(gate74inter4), .b(gate74inter3), .O(gate74inter5));
  nor2  gate1701(.a(gate74inter5), .b(gate74inter2), .O(gate74inter6));
  inv1  gate1702(.a(G5), .O(gate74inter7));
  inv1  gate1703(.a(G314), .O(gate74inter8));
  nand2 gate1704(.a(gate74inter8), .b(gate74inter7), .O(gate74inter9));
  nand2 gate1705(.a(s_165), .b(gate74inter3), .O(gate74inter10));
  nor2  gate1706(.a(gate74inter10), .b(gate74inter9), .O(gate74inter11));
  nor2  gate1707(.a(gate74inter11), .b(gate74inter6), .O(gate74inter12));
  nand2 gate1708(.a(gate74inter12), .b(gate74inter1), .O(G395));
nand2 gate75( .a(G9), .b(G317), .O(G396) );
nand2 gate76( .a(G13), .b(G317), .O(G397) );
nand2 gate77( .a(G2), .b(G320), .O(G398) );
nand2 gate78( .a(G6), .b(G320), .O(G399) );

  xor2  gate1233(.a(G323), .b(G10), .O(gate79inter0));
  nand2 gate1234(.a(gate79inter0), .b(s_98), .O(gate79inter1));
  and2  gate1235(.a(G323), .b(G10), .O(gate79inter2));
  inv1  gate1236(.a(s_98), .O(gate79inter3));
  inv1  gate1237(.a(s_99), .O(gate79inter4));
  nand2 gate1238(.a(gate79inter4), .b(gate79inter3), .O(gate79inter5));
  nor2  gate1239(.a(gate79inter5), .b(gate79inter2), .O(gate79inter6));
  inv1  gate1240(.a(G10), .O(gate79inter7));
  inv1  gate1241(.a(G323), .O(gate79inter8));
  nand2 gate1242(.a(gate79inter8), .b(gate79inter7), .O(gate79inter9));
  nand2 gate1243(.a(s_99), .b(gate79inter3), .O(gate79inter10));
  nor2  gate1244(.a(gate79inter10), .b(gate79inter9), .O(gate79inter11));
  nor2  gate1245(.a(gate79inter11), .b(gate79inter6), .O(gate79inter12));
  nand2 gate1246(.a(gate79inter12), .b(gate79inter1), .O(G400));
nand2 gate80( .a(G14), .b(G323), .O(G401) );
nand2 gate81( .a(G3), .b(G326), .O(G402) );
nand2 gate82( .a(G7), .b(G326), .O(G403) );
nand2 gate83( .a(G11), .b(G329), .O(G404) );
nand2 gate84( .a(G15), .b(G329), .O(G405) );
nand2 gate85( .a(G4), .b(G332), .O(G406) );
nand2 gate86( .a(G8), .b(G332), .O(G407) );
nand2 gate87( .a(G12), .b(G335), .O(G408) );
nand2 gate88( .a(G16), .b(G335), .O(G409) );
nand2 gate89( .a(G17), .b(G338), .O(G410) );
nand2 gate90( .a(G21), .b(G338), .O(G411) );
nand2 gate91( .a(G25), .b(G341), .O(G412) );
nand2 gate92( .a(G29), .b(G341), .O(G413) );
nand2 gate93( .a(G18), .b(G344), .O(G414) );

  xor2  gate1331(.a(G344), .b(G22), .O(gate94inter0));
  nand2 gate1332(.a(gate94inter0), .b(s_112), .O(gate94inter1));
  and2  gate1333(.a(G344), .b(G22), .O(gate94inter2));
  inv1  gate1334(.a(s_112), .O(gate94inter3));
  inv1  gate1335(.a(s_113), .O(gate94inter4));
  nand2 gate1336(.a(gate94inter4), .b(gate94inter3), .O(gate94inter5));
  nor2  gate1337(.a(gate94inter5), .b(gate94inter2), .O(gate94inter6));
  inv1  gate1338(.a(G22), .O(gate94inter7));
  inv1  gate1339(.a(G344), .O(gate94inter8));
  nand2 gate1340(.a(gate94inter8), .b(gate94inter7), .O(gate94inter9));
  nand2 gate1341(.a(s_113), .b(gate94inter3), .O(gate94inter10));
  nor2  gate1342(.a(gate94inter10), .b(gate94inter9), .O(gate94inter11));
  nor2  gate1343(.a(gate94inter11), .b(gate94inter6), .O(gate94inter12));
  nand2 gate1344(.a(gate94inter12), .b(gate94inter1), .O(G415));
nand2 gate95( .a(G26), .b(G347), .O(G416) );
nand2 gate96( .a(G30), .b(G347), .O(G417) );

  xor2  gate1387(.a(G350), .b(G19), .O(gate97inter0));
  nand2 gate1388(.a(gate97inter0), .b(s_120), .O(gate97inter1));
  and2  gate1389(.a(G350), .b(G19), .O(gate97inter2));
  inv1  gate1390(.a(s_120), .O(gate97inter3));
  inv1  gate1391(.a(s_121), .O(gate97inter4));
  nand2 gate1392(.a(gate97inter4), .b(gate97inter3), .O(gate97inter5));
  nor2  gate1393(.a(gate97inter5), .b(gate97inter2), .O(gate97inter6));
  inv1  gate1394(.a(G19), .O(gate97inter7));
  inv1  gate1395(.a(G350), .O(gate97inter8));
  nand2 gate1396(.a(gate97inter8), .b(gate97inter7), .O(gate97inter9));
  nand2 gate1397(.a(s_121), .b(gate97inter3), .O(gate97inter10));
  nor2  gate1398(.a(gate97inter10), .b(gate97inter9), .O(gate97inter11));
  nor2  gate1399(.a(gate97inter11), .b(gate97inter6), .O(gate97inter12));
  nand2 gate1400(.a(gate97inter12), .b(gate97inter1), .O(G418));
nand2 gate98( .a(G23), .b(G350), .O(G419) );
nand2 gate99( .a(G27), .b(G353), .O(G420) );
nand2 gate100( .a(G31), .b(G353), .O(G421) );
nand2 gate101( .a(G20), .b(G356), .O(G422) );

  xor2  gate1303(.a(G356), .b(G24), .O(gate102inter0));
  nand2 gate1304(.a(gate102inter0), .b(s_108), .O(gate102inter1));
  and2  gate1305(.a(G356), .b(G24), .O(gate102inter2));
  inv1  gate1306(.a(s_108), .O(gate102inter3));
  inv1  gate1307(.a(s_109), .O(gate102inter4));
  nand2 gate1308(.a(gate102inter4), .b(gate102inter3), .O(gate102inter5));
  nor2  gate1309(.a(gate102inter5), .b(gate102inter2), .O(gate102inter6));
  inv1  gate1310(.a(G24), .O(gate102inter7));
  inv1  gate1311(.a(G356), .O(gate102inter8));
  nand2 gate1312(.a(gate102inter8), .b(gate102inter7), .O(gate102inter9));
  nand2 gate1313(.a(s_109), .b(gate102inter3), .O(gate102inter10));
  nor2  gate1314(.a(gate102inter10), .b(gate102inter9), .O(gate102inter11));
  nor2  gate1315(.a(gate102inter11), .b(gate102inter6), .O(gate102inter12));
  nand2 gate1316(.a(gate102inter12), .b(gate102inter1), .O(G423));
nand2 gate103( .a(G28), .b(G359), .O(G424) );
nand2 gate104( .a(G32), .b(G359), .O(G425) );
nand2 gate105( .a(G362), .b(G363), .O(G426) );
nand2 gate106( .a(G364), .b(G365), .O(G429) );

  xor2  gate1835(.a(G367), .b(G366), .O(gate107inter0));
  nand2 gate1836(.a(gate107inter0), .b(s_184), .O(gate107inter1));
  and2  gate1837(.a(G367), .b(G366), .O(gate107inter2));
  inv1  gate1838(.a(s_184), .O(gate107inter3));
  inv1  gate1839(.a(s_185), .O(gate107inter4));
  nand2 gate1840(.a(gate107inter4), .b(gate107inter3), .O(gate107inter5));
  nor2  gate1841(.a(gate107inter5), .b(gate107inter2), .O(gate107inter6));
  inv1  gate1842(.a(G366), .O(gate107inter7));
  inv1  gate1843(.a(G367), .O(gate107inter8));
  nand2 gate1844(.a(gate107inter8), .b(gate107inter7), .O(gate107inter9));
  nand2 gate1845(.a(s_185), .b(gate107inter3), .O(gate107inter10));
  nor2  gate1846(.a(gate107inter10), .b(gate107inter9), .O(gate107inter11));
  nor2  gate1847(.a(gate107inter11), .b(gate107inter6), .O(gate107inter12));
  nand2 gate1848(.a(gate107inter12), .b(gate107inter1), .O(G432));
nand2 gate108( .a(G368), .b(G369), .O(G435) );
nand2 gate109( .a(G370), .b(G371), .O(G438) );
nand2 gate110( .a(G372), .b(G373), .O(G441) );
nand2 gate111( .a(G374), .b(G375), .O(G444) );

  xor2  gate1079(.a(G377), .b(G376), .O(gate112inter0));
  nand2 gate1080(.a(gate112inter0), .b(s_76), .O(gate112inter1));
  and2  gate1081(.a(G377), .b(G376), .O(gate112inter2));
  inv1  gate1082(.a(s_76), .O(gate112inter3));
  inv1  gate1083(.a(s_77), .O(gate112inter4));
  nand2 gate1084(.a(gate112inter4), .b(gate112inter3), .O(gate112inter5));
  nor2  gate1085(.a(gate112inter5), .b(gate112inter2), .O(gate112inter6));
  inv1  gate1086(.a(G376), .O(gate112inter7));
  inv1  gate1087(.a(G377), .O(gate112inter8));
  nand2 gate1088(.a(gate112inter8), .b(gate112inter7), .O(gate112inter9));
  nand2 gate1089(.a(s_77), .b(gate112inter3), .O(gate112inter10));
  nor2  gate1090(.a(gate112inter10), .b(gate112inter9), .O(gate112inter11));
  nor2  gate1091(.a(gate112inter11), .b(gate112inter6), .O(gate112inter12));
  nand2 gate1092(.a(gate112inter12), .b(gate112inter1), .O(G447));
nand2 gate113( .a(G378), .b(G379), .O(G450) );
nand2 gate114( .a(G380), .b(G381), .O(G453) );
nand2 gate115( .a(G382), .b(G383), .O(G456) );
nand2 gate116( .a(G384), .b(G385), .O(G459) );
nand2 gate117( .a(G386), .b(G387), .O(G462) );
nand2 gate118( .a(G388), .b(G389), .O(G465) );
nand2 gate119( .a(G390), .b(G391), .O(G468) );

  xor2  gate1527(.a(G393), .b(G392), .O(gate120inter0));
  nand2 gate1528(.a(gate120inter0), .b(s_140), .O(gate120inter1));
  and2  gate1529(.a(G393), .b(G392), .O(gate120inter2));
  inv1  gate1530(.a(s_140), .O(gate120inter3));
  inv1  gate1531(.a(s_141), .O(gate120inter4));
  nand2 gate1532(.a(gate120inter4), .b(gate120inter3), .O(gate120inter5));
  nor2  gate1533(.a(gate120inter5), .b(gate120inter2), .O(gate120inter6));
  inv1  gate1534(.a(G392), .O(gate120inter7));
  inv1  gate1535(.a(G393), .O(gate120inter8));
  nand2 gate1536(.a(gate120inter8), .b(gate120inter7), .O(gate120inter9));
  nand2 gate1537(.a(s_141), .b(gate120inter3), .O(gate120inter10));
  nor2  gate1538(.a(gate120inter10), .b(gate120inter9), .O(gate120inter11));
  nor2  gate1539(.a(gate120inter11), .b(gate120inter6), .O(gate120inter12));
  nand2 gate1540(.a(gate120inter12), .b(gate120inter1), .O(G471));
nand2 gate121( .a(G394), .b(G395), .O(G474) );

  xor2  gate1821(.a(G397), .b(G396), .O(gate122inter0));
  nand2 gate1822(.a(gate122inter0), .b(s_182), .O(gate122inter1));
  and2  gate1823(.a(G397), .b(G396), .O(gate122inter2));
  inv1  gate1824(.a(s_182), .O(gate122inter3));
  inv1  gate1825(.a(s_183), .O(gate122inter4));
  nand2 gate1826(.a(gate122inter4), .b(gate122inter3), .O(gate122inter5));
  nor2  gate1827(.a(gate122inter5), .b(gate122inter2), .O(gate122inter6));
  inv1  gate1828(.a(G396), .O(gate122inter7));
  inv1  gate1829(.a(G397), .O(gate122inter8));
  nand2 gate1830(.a(gate122inter8), .b(gate122inter7), .O(gate122inter9));
  nand2 gate1831(.a(s_183), .b(gate122inter3), .O(gate122inter10));
  nor2  gate1832(.a(gate122inter10), .b(gate122inter9), .O(gate122inter11));
  nor2  gate1833(.a(gate122inter11), .b(gate122inter6), .O(gate122inter12));
  nand2 gate1834(.a(gate122inter12), .b(gate122inter1), .O(G477));

  xor2  gate1485(.a(G399), .b(G398), .O(gate123inter0));
  nand2 gate1486(.a(gate123inter0), .b(s_134), .O(gate123inter1));
  and2  gate1487(.a(G399), .b(G398), .O(gate123inter2));
  inv1  gate1488(.a(s_134), .O(gate123inter3));
  inv1  gate1489(.a(s_135), .O(gate123inter4));
  nand2 gate1490(.a(gate123inter4), .b(gate123inter3), .O(gate123inter5));
  nor2  gate1491(.a(gate123inter5), .b(gate123inter2), .O(gate123inter6));
  inv1  gate1492(.a(G398), .O(gate123inter7));
  inv1  gate1493(.a(G399), .O(gate123inter8));
  nand2 gate1494(.a(gate123inter8), .b(gate123inter7), .O(gate123inter9));
  nand2 gate1495(.a(s_135), .b(gate123inter3), .O(gate123inter10));
  nor2  gate1496(.a(gate123inter10), .b(gate123inter9), .O(gate123inter11));
  nor2  gate1497(.a(gate123inter11), .b(gate123inter6), .O(gate123inter12));
  nand2 gate1498(.a(gate123inter12), .b(gate123inter1), .O(G480));

  xor2  gate729(.a(G401), .b(G400), .O(gate124inter0));
  nand2 gate730(.a(gate124inter0), .b(s_26), .O(gate124inter1));
  and2  gate731(.a(G401), .b(G400), .O(gate124inter2));
  inv1  gate732(.a(s_26), .O(gate124inter3));
  inv1  gate733(.a(s_27), .O(gate124inter4));
  nand2 gate734(.a(gate124inter4), .b(gate124inter3), .O(gate124inter5));
  nor2  gate735(.a(gate124inter5), .b(gate124inter2), .O(gate124inter6));
  inv1  gate736(.a(G400), .O(gate124inter7));
  inv1  gate737(.a(G401), .O(gate124inter8));
  nand2 gate738(.a(gate124inter8), .b(gate124inter7), .O(gate124inter9));
  nand2 gate739(.a(s_27), .b(gate124inter3), .O(gate124inter10));
  nor2  gate740(.a(gate124inter10), .b(gate124inter9), .O(gate124inter11));
  nor2  gate741(.a(gate124inter11), .b(gate124inter6), .O(gate124inter12));
  nand2 gate742(.a(gate124inter12), .b(gate124inter1), .O(G483));
nand2 gate125( .a(G402), .b(G403), .O(G486) );
nand2 gate126( .a(G404), .b(G405), .O(G489) );
nand2 gate127( .a(G406), .b(G407), .O(G492) );
nand2 gate128( .a(G408), .b(G409), .O(G495) );
nand2 gate129( .a(G410), .b(G411), .O(G498) );
nand2 gate130( .a(G412), .b(G413), .O(G501) );

  xor2  gate1569(.a(G415), .b(G414), .O(gate131inter0));
  nand2 gate1570(.a(gate131inter0), .b(s_146), .O(gate131inter1));
  and2  gate1571(.a(G415), .b(G414), .O(gate131inter2));
  inv1  gate1572(.a(s_146), .O(gate131inter3));
  inv1  gate1573(.a(s_147), .O(gate131inter4));
  nand2 gate1574(.a(gate131inter4), .b(gate131inter3), .O(gate131inter5));
  nor2  gate1575(.a(gate131inter5), .b(gate131inter2), .O(gate131inter6));
  inv1  gate1576(.a(G414), .O(gate131inter7));
  inv1  gate1577(.a(G415), .O(gate131inter8));
  nand2 gate1578(.a(gate131inter8), .b(gate131inter7), .O(gate131inter9));
  nand2 gate1579(.a(s_147), .b(gate131inter3), .O(gate131inter10));
  nor2  gate1580(.a(gate131inter10), .b(gate131inter9), .O(gate131inter11));
  nor2  gate1581(.a(gate131inter11), .b(gate131inter6), .O(gate131inter12));
  nand2 gate1582(.a(gate131inter12), .b(gate131inter1), .O(G504));
nand2 gate132( .a(G416), .b(G417), .O(G507) );
nand2 gate133( .a(G418), .b(G419), .O(G510) );
nand2 gate134( .a(G420), .b(G421), .O(G513) );
nand2 gate135( .a(G422), .b(G423), .O(G516) );

  xor2  gate1163(.a(G425), .b(G424), .O(gate136inter0));
  nand2 gate1164(.a(gate136inter0), .b(s_88), .O(gate136inter1));
  and2  gate1165(.a(G425), .b(G424), .O(gate136inter2));
  inv1  gate1166(.a(s_88), .O(gate136inter3));
  inv1  gate1167(.a(s_89), .O(gate136inter4));
  nand2 gate1168(.a(gate136inter4), .b(gate136inter3), .O(gate136inter5));
  nor2  gate1169(.a(gate136inter5), .b(gate136inter2), .O(gate136inter6));
  inv1  gate1170(.a(G424), .O(gate136inter7));
  inv1  gate1171(.a(G425), .O(gate136inter8));
  nand2 gate1172(.a(gate136inter8), .b(gate136inter7), .O(gate136inter9));
  nand2 gate1173(.a(s_89), .b(gate136inter3), .O(gate136inter10));
  nor2  gate1174(.a(gate136inter10), .b(gate136inter9), .O(gate136inter11));
  nor2  gate1175(.a(gate136inter11), .b(gate136inter6), .O(gate136inter12));
  nand2 gate1176(.a(gate136inter12), .b(gate136inter1), .O(G519));
nand2 gate137( .a(G426), .b(G429), .O(G522) );
nand2 gate138( .a(G432), .b(G435), .O(G525) );
nand2 gate139( .a(G438), .b(G441), .O(G528) );
nand2 gate140( .a(G444), .b(G447), .O(G531) );
nand2 gate141( .a(G450), .b(G453), .O(G534) );

  xor2  gate1653(.a(G459), .b(G456), .O(gate142inter0));
  nand2 gate1654(.a(gate142inter0), .b(s_158), .O(gate142inter1));
  and2  gate1655(.a(G459), .b(G456), .O(gate142inter2));
  inv1  gate1656(.a(s_158), .O(gate142inter3));
  inv1  gate1657(.a(s_159), .O(gate142inter4));
  nand2 gate1658(.a(gate142inter4), .b(gate142inter3), .O(gate142inter5));
  nor2  gate1659(.a(gate142inter5), .b(gate142inter2), .O(gate142inter6));
  inv1  gate1660(.a(G456), .O(gate142inter7));
  inv1  gate1661(.a(G459), .O(gate142inter8));
  nand2 gate1662(.a(gate142inter8), .b(gate142inter7), .O(gate142inter9));
  nand2 gate1663(.a(s_159), .b(gate142inter3), .O(gate142inter10));
  nor2  gate1664(.a(gate142inter10), .b(gate142inter9), .O(gate142inter11));
  nor2  gate1665(.a(gate142inter11), .b(gate142inter6), .O(gate142inter12));
  nand2 gate1666(.a(gate142inter12), .b(gate142inter1), .O(G537));
nand2 gate143( .a(G462), .b(G465), .O(G540) );
nand2 gate144( .a(G468), .b(G471), .O(G543) );

  xor2  gate1877(.a(G477), .b(G474), .O(gate145inter0));
  nand2 gate1878(.a(gate145inter0), .b(s_190), .O(gate145inter1));
  and2  gate1879(.a(G477), .b(G474), .O(gate145inter2));
  inv1  gate1880(.a(s_190), .O(gate145inter3));
  inv1  gate1881(.a(s_191), .O(gate145inter4));
  nand2 gate1882(.a(gate145inter4), .b(gate145inter3), .O(gate145inter5));
  nor2  gate1883(.a(gate145inter5), .b(gate145inter2), .O(gate145inter6));
  inv1  gate1884(.a(G474), .O(gate145inter7));
  inv1  gate1885(.a(G477), .O(gate145inter8));
  nand2 gate1886(.a(gate145inter8), .b(gate145inter7), .O(gate145inter9));
  nand2 gate1887(.a(s_191), .b(gate145inter3), .O(gate145inter10));
  nor2  gate1888(.a(gate145inter10), .b(gate145inter9), .O(gate145inter11));
  nor2  gate1889(.a(gate145inter11), .b(gate145inter6), .O(gate145inter12));
  nand2 gate1890(.a(gate145inter12), .b(gate145inter1), .O(G546));
nand2 gate146( .a(G480), .b(G483), .O(G549) );

  xor2  gate589(.a(G489), .b(G486), .O(gate147inter0));
  nand2 gate590(.a(gate147inter0), .b(s_6), .O(gate147inter1));
  and2  gate591(.a(G489), .b(G486), .O(gate147inter2));
  inv1  gate592(.a(s_6), .O(gate147inter3));
  inv1  gate593(.a(s_7), .O(gate147inter4));
  nand2 gate594(.a(gate147inter4), .b(gate147inter3), .O(gate147inter5));
  nor2  gate595(.a(gate147inter5), .b(gate147inter2), .O(gate147inter6));
  inv1  gate596(.a(G486), .O(gate147inter7));
  inv1  gate597(.a(G489), .O(gate147inter8));
  nand2 gate598(.a(gate147inter8), .b(gate147inter7), .O(gate147inter9));
  nand2 gate599(.a(s_7), .b(gate147inter3), .O(gate147inter10));
  nor2  gate600(.a(gate147inter10), .b(gate147inter9), .O(gate147inter11));
  nor2  gate601(.a(gate147inter11), .b(gate147inter6), .O(gate147inter12));
  nand2 gate602(.a(gate147inter12), .b(gate147inter1), .O(G552));

  xor2  gate1429(.a(G495), .b(G492), .O(gate148inter0));
  nand2 gate1430(.a(gate148inter0), .b(s_126), .O(gate148inter1));
  and2  gate1431(.a(G495), .b(G492), .O(gate148inter2));
  inv1  gate1432(.a(s_126), .O(gate148inter3));
  inv1  gate1433(.a(s_127), .O(gate148inter4));
  nand2 gate1434(.a(gate148inter4), .b(gate148inter3), .O(gate148inter5));
  nor2  gate1435(.a(gate148inter5), .b(gate148inter2), .O(gate148inter6));
  inv1  gate1436(.a(G492), .O(gate148inter7));
  inv1  gate1437(.a(G495), .O(gate148inter8));
  nand2 gate1438(.a(gate148inter8), .b(gate148inter7), .O(gate148inter9));
  nand2 gate1439(.a(s_127), .b(gate148inter3), .O(gate148inter10));
  nor2  gate1440(.a(gate148inter10), .b(gate148inter9), .O(gate148inter11));
  nor2  gate1441(.a(gate148inter11), .b(gate148inter6), .O(gate148inter12));
  nand2 gate1442(.a(gate148inter12), .b(gate148inter1), .O(G555));
nand2 gate149( .a(G498), .b(G501), .O(G558) );

  xor2  gate1737(.a(G507), .b(G504), .O(gate150inter0));
  nand2 gate1738(.a(gate150inter0), .b(s_170), .O(gate150inter1));
  and2  gate1739(.a(G507), .b(G504), .O(gate150inter2));
  inv1  gate1740(.a(s_170), .O(gate150inter3));
  inv1  gate1741(.a(s_171), .O(gate150inter4));
  nand2 gate1742(.a(gate150inter4), .b(gate150inter3), .O(gate150inter5));
  nor2  gate1743(.a(gate150inter5), .b(gate150inter2), .O(gate150inter6));
  inv1  gate1744(.a(G504), .O(gate150inter7));
  inv1  gate1745(.a(G507), .O(gate150inter8));
  nand2 gate1746(.a(gate150inter8), .b(gate150inter7), .O(gate150inter9));
  nand2 gate1747(.a(s_171), .b(gate150inter3), .O(gate150inter10));
  nor2  gate1748(.a(gate150inter10), .b(gate150inter9), .O(gate150inter11));
  nor2  gate1749(.a(gate150inter11), .b(gate150inter6), .O(gate150inter12));
  nand2 gate1750(.a(gate150inter12), .b(gate150inter1), .O(G561));
nand2 gate151( .a(G510), .b(G513), .O(G564) );
nand2 gate152( .a(G516), .b(G519), .O(G567) );

  xor2  gate1555(.a(G522), .b(G426), .O(gate153inter0));
  nand2 gate1556(.a(gate153inter0), .b(s_144), .O(gate153inter1));
  and2  gate1557(.a(G522), .b(G426), .O(gate153inter2));
  inv1  gate1558(.a(s_144), .O(gate153inter3));
  inv1  gate1559(.a(s_145), .O(gate153inter4));
  nand2 gate1560(.a(gate153inter4), .b(gate153inter3), .O(gate153inter5));
  nor2  gate1561(.a(gate153inter5), .b(gate153inter2), .O(gate153inter6));
  inv1  gate1562(.a(G426), .O(gate153inter7));
  inv1  gate1563(.a(G522), .O(gate153inter8));
  nand2 gate1564(.a(gate153inter8), .b(gate153inter7), .O(gate153inter9));
  nand2 gate1565(.a(s_145), .b(gate153inter3), .O(gate153inter10));
  nor2  gate1566(.a(gate153inter10), .b(gate153inter9), .O(gate153inter11));
  nor2  gate1567(.a(gate153inter11), .b(gate153inter6), .O(gate153inter12));
  nand2 gate1568(.a(gate153inter12), .b(gate153inter1), .O(G570));

  xor2  gate673(.a(G522), .b(G429), .O(gate154inter0));
  nand2 gate674(.a(gate154inter0), .b(s_18), .O(gate154inter1));
  and2  gate675(.a(G522), .b(G429), .O(gate154inter2));
  inv1  gate676(.a(s_18), .O(gate154inter3));
  inv1  gate677(.a(s_19), .O(gate154inter4));
  nand2 gate678(.a(gate154inter4), .b(gate154inter3), .O(gate154inter5));
  nor2  gate679(.a(gate154inter5), .b(gate154inter2), .O(gate154inter6));
  inv1  gate680(.a(G429), .O(gate154inter7));
  inv1  gate681(.a(G522), .O(gate154inter8));
  nand2 gate682(.a(gate154inter8), .b(gate154inter7), .O(gate154inter9));
  nand2 gate683(.a(s_19), .b(gate154inter3), .O(gate154inter10));
  nor2  gate684(.a(gate154inter10), .b(gate154inter9), .O(gate154inter11));
  nor2  gate685(.a(gate154inter11), .b(gate154inter6), .O(gate154inter12));
  nand2 gate686(.a(gate154inter12), .b(gate154inter1), .O(G571));
nand2 gate155( .a(G432), .b(G525), .O(G572) );
nand2 gate156( .a(G435), .b(G525), .O(G573) );
nand2 gate157( .a(G438), .b(G528), .O(G574) );
nand2 gate158( .a(G441), .b(G528), .O(G575) );
nand2 gate159( .a(G444), .b(G531), .O(G576) );

  xor2  gate575(.a(G531), .b(G447), .O(gate160inter0));
  nand2 gate576(.a(gate160inter0), .b(s_4), .O(gate160inter1));
  and2  gate577(.a(G531), .b(G447), .O(gate160inter2));
  inv1  gate578(.a(s_4), .O(gate160inter3));
  inv1  gate579(.a(s_5), .O(gate160inter4));
  nand2 gate580(.a(gate160inter4), .b(gate160inter3), .O(gate160inter5));
  nor2  gate581(.a(gate160inter5), .b(gate160inter2), .O(gate160inter6));
  inv1  gate582(.a(G447), .O(gate160inter7));
  inv1  gate583(.a(G531), .O(gate160inter8));
  nand2 gate584(.a(gate160inter8), .b(gate160inter7), .O(gate160inter9));
  nand2 gate585(.a(s_5), .b(gate160inter3), .O(gate160inter10));
  nor2  gate586(.a(gate160inter10), .b(gate160inter9), .O(gate160inter11));
  nor2  gate587(.a(gate160inter11), .b(gate160inter6), .O(gate160inter12));
  nand2 gate588(.a(gate160inter12), .b(gate160inter1), .O(G577));
nand2 gate161( .a(G450), .b(G534), .O(G578) );

  xor2  gate981(.a(G534), .b(G453), .O(gate162inter0));
  nand2 gate982(.a(gate162inter0), .b(s_62), .O(gate162inter1));
  and2  gate983(.a(G534), .b(G453), .O(gate162inter2));
  inv1  gate984(.a(s_62), .O(gate162inter3));
  inv1  gate985(.a(s_63), .O(gate162inter4));
  nand2 gate986(.a(gate162inter4), .b(gate162inter3), .O(gate162inter5));
  nor2  gate987(.a(gate162inter5), .b(gate162inter2), .O(gate162inter6));
  inv1  gate988(.a(G453), .O(gate162inter7));
  inv1  gate989(.a(G534), .O(gate162inter8));
  nand2 gate990(.a(gate162inter8), .b(gate162inter7), .O(gate162inter9));
  nand2 gate991(.a(s_63), .b(gate162inter3), .O(gate162inter10));
  nor2  gate992(.a(gate162inter10), .b(gate162inter9), .O(gate162inter11));
  nor2  gate993(.a(gate162inter11), .b(gate162inter6), .O(gate162inter12));
  nand2 gate994(.a(gate162inter12), .b(gate162inter1), .O(G579));
nand2 gate163( .a(G456), .b(G537), .O(G580) );

  xor2  gate1107(.a(G537), .b(G459), .O(gate164inter0));
  nand2 gate1108(.a(gate164inter0), .b(s_80), .O(gate164inter1));
  and2  gate1109(.a(G537), .b(G459), .O(gate164inter2));
  inv1  gate1110(.a(s_80), .O(gate164inter3));
  inv1  gate1111(.a(s_81), .O(gate164inter4));
  nand2 gate1112(.a(gate164inter4), .b(gate164inter3), .O(gate164inter5));
  nor2  gate1113(.a(gate164inter5), .b(gate164inter2), .O(gate164inter6));
  inv1  gate1114(.a(G459), .O(gate164inter7));
  inv1  gate1115(.a(G537), .O(gate164inter8));
  nand2 gate1116(.a(gate164inter8), .b(gate164inter7), .O(gate164inter9));
  nand2 gate1117(.a(s_81), .b(gate164inter3), .O(gate164inter10));
  nor2  gate1118(.a(gate164inter10), .b(gate164inter9), .O(gate164inter11));
  nor2  gate1119(.a(gate164inter11), .b(gate164inter6), .O(gate164inter12));
  nand2 gate1120(.a(gate164inter12), .b(gate164inter1), .O(G581));
nand2 gate165( .a(G462), .b(G540), .O(G582) );
nand2 gate166( .a(G465), .b(G540), .O(G583) );
nand2 gate167( .a(G468), .b(G543), .O(G584) );
nand2 gate168( .a(G471), .b(G543), .O(G585) );
nand2 gate169( .a(G474), .b(G546), .O(G586) );
nand2 gate170( .a(G477), .b(G546), .O(G587) );

  xor2  gate1093(.a(G549), .b(G480), .O(gate171inter0));
  nand2 gate1094(.a(gate171inter0), .b(s_78), .O(gate171inter1));
  and2  gate1095(.a(G549), .b(G480), .O(gate171inter2));
  inv1  gate1096(.a(s_78), .O(gate171inter3));
  inv1  gate1097(.a(s_79), .O(gate171inter4));
  nand2 gate1098(.a(gate171inter4), .b(gate171inter3), .O(gate171inter5));
  nor2  gate1099(.a(gate171inter5), .b(gate171inter2), .O(gate171inter6));
  inv1  gate1100(.a(G480), .O(gate171inter7));
  inv1  gate1101(.a(G549), .O(gate171inter8));
  nand2 gate1102(.a(gate171inter8), .b(gate171inter7), .O(gate171inter9));
  nand2 gate1103(.a(s_79), .b(gate171inter3), .O(gate171inter10));
  nor2  gate1104(.a(gate171inter10), .b(gate171inter9), .O(gate171inter11));
  nor2  gate1105(.a(gate171inter11), .b(gate171inter6), .O(gate171inter12));
  nand2 gate1106(.a(gate171inter12), .b(gate171inter1), .O(G588));
nand2 gate172( .a(G483), .b(G549), .O(G589) );

  xor2  gate1807(.a(G552), .b(G486), .O(gate173inter0));
  nand2 gate1808(.a(gate173inter0), .b(s_180), .O(gate173inter1));
  and2  gate1809(.a(G552), .b(G486), .O(gate173inter2));
  inv1  gate1810(.a(s_180), .O(gate173inter3));
  inv1  gate1811(.a(s_181), .O(gate173inter4));
  nand2 gate1812(.a(gate173inter4), .b(gate173inter3), .O(gate173inter5));
  nor2  gate1813(.a(gate173inter5), .b(gate173inter2), .O(gate173inter6));
  inv1  gate1814(.a(G486), .O(gate173inter7));
  inv1  gate1815(.a(G552), .O(gate173inter8));
  nand2 gate1816(.a(gate173inter8), .b(gate173inter7), .O(gate173inter9));
  nand2 gate1817(.a(s_181), .b(gate173inter3), .O(gate173inter10));
  nor2  gate1818(.a(gate173inter10), .b(gate173inter9), .O(gate173inter11));
  nor2  gate1819(.a(gate173inter11), .b(gate173inter6), .O(gate173inter12));
  nand2 gate1820(.a(gate173inter12), .b(gate173inter1), .O(G590));
nand2 gate174( .a(G489), .b(G552), .O(G591) );
nand2 gate175( .a(G492), .b(G555), .O(G592) );
nand2 gate176( .a(G495), .b(G555), .O(G593) );

  xor2  gate561(.a(G558), .b(G498), .O(gate177inter0));
  nand2 gate562(.a(gate177inter0), .b(s_2), .O(gate177inter1));
  and2  gate563(.a(G558), .b(G498), .O(gate177inter2));
  inv1  gate564(.a(s_2), .O(gate177inter3));
  inv1  gate565(.a(s_3), .O(gate177inter4));
  nand2 gate566(.a(gate177inter4), .b(gate177inter3), .O(gate177inter5));
  nor2  gate567(.a(gate177inter5), .b(gate177inter2), .O(gate177inter6));
  inv1  gate568(.a(G498), .O(gate177inter7));
  inv1  gate569(.a(G558), .O(gate177inter8));
  nand2 gate570(.a(gate177inter8), .b(gate177inter7), .O(gate177inter9));
  nand2 gate571(.a(s_3), .b(gate177inter3), .O(gate177inter10));
  nor2  gate572(.a(gate177inter10), .b(gate177inter9), .O(gate177inter11));
  nor2  gate573(.a(gate177inter11), .b(gate177inter6), .O(gate177inter12));
  nand2 gate574(.a(gate177inter12), .b(gate177inter1), .O(G594));
nand2 gate178( .a(G501), .b(G558), .O(G595) );
nand2 gate179( .a(G504), .b(G561), .O(G596) );
nand2 gate180( .a(G507), .b(G561), .O(G597) );

  xor2  gate1177(.a(G564), .b(G510), .O(gate181inter0));
  nand2 gate1178(.a(gate181inter0), .b(s_90), .O(gate181inter1));
  and2  gate1179(.a(G564), .b(G510), .O(gate181inter2));
  inv1  gate1180(.a(s_90), .O(gate181inter3));
  inv1  gate1181(.a(s_91), .O(gate181inter4));
  nand2 gate1182(.a(gate181inter4), .b(gate181inter3), .O(gate181inter5));
  nor2  gate1183(.a(gate181inter5), .b(gate181inter2), .O(gate181inter6));
  inv1  gate1184(.a(G510), .O(gate181inter7));
  inv1  gate1185(.a(G564), .O(gate181inter8));
  nand2 gate1186(.a(gate181inter8), .b(gate181inter7), .O(gate181inter9));
  nand2 gate1187(.a(s_91), .b(gate181inter3), .O(gate181inter10));
  nor2  gate1188(.a(gate181inter10), .b(gate181inter9), .O(gate181inter11));
  nor2  gate1189(.a(gate181inter11), .b(gate181inter6), .O(gate181inter12));
  nand2 gate1190(.a(gate181inter12), .b(gate181inter1), .O(G598));
nand2 gate182( .a(G513), .b(G564), .O(G599) );

  xor2  gate1681(.a(G567), .b(G516), .O(gate183inter0));
  nand2 gate1682(.a(gate183inter0), .b(s_162), .O(gate183inter1));
  and2  gate1683(.a(G567), .b(G516), .O(gate183inter2));
  inv1  gate1684(.a(s_162), .O(gate183inter3));
  inv1  gate1685(.a(s_163), .O(gate183inter4));
  nand2 gate1686(.a(gate183inter4), .b(gate183inter3), .O(gate183inter5));
  nor2  gate1687(.a(gate183inter5), .b(gate183inter2), .O(gate183inter6));
  inv1  gate1688(.a(G516), .O(gate183inter7));
  inv1  gate1689(.a(G567), .O(gate183inter8));
  nand2 gate1690(.a(gate183inter8), .b(gate183inter7), .O(gate183inter9));
  nand2 gate1691(.a(s_163), .b(gate183inter3), .O(gate183inter10));
  nor2  gate1692(.a(gate183inter10), .b(gate183inter9), .O(gate183inter11));
  nor2  gate1693(.a(gate183inter11), .b(gate183inter6), .O(gate183inter12));
  nand2 gate1694(.a(gate183inter12), .b(gate183inter1), .O(G600));
nand2 gate184( .a(G519), .b(G567), .O(G601) );
nand2 gate185( .a(G570), .b(G571), .O(G602) );
nand2 gate186( .a(G572), .b(G573), .O(G607) );
nand2 gate187( .a(G574), .b(G575), .O(G612) );
nand2 gate188( .a(G576), .b(G577), .O(G617) );
nand2 gate189( .a(G578), .b(G579), .O(G622) );
nand2 gate190( .a(G580), .b(G581), .O(G627) );
nand2 gate191( .a(G582), .b(G583), .O(G632) );
nand2 gate192( .a(G584), .b(G585), .O(G637) );
nand2 gate193( .a(G586), .b(G587), .O(G642) );
nand2 gate194( .a(G588), .b(G589), .O(G645) );

  xor2  gate1023(.a(G591), .b(G590), .O(gate195inter0));
  nand2 gate1024(.a(gate195inter0), .b(s_68), .O(gate195inter1));
  and2  gate1025(.a(G591), .b(G590), .O(gate195inter2));
  inv1  gate1026(.a(s_68), .O(gate195inter3));
  inv1  gate1027(.a(s_69), .O(gate195inter4));
  nand2 gate1028(.a(gate195inter4), .b(gate195inter3), .O(gate195inter5));
  nor2  gate1029(.a(gate195inter5), .b(gate195inter2), .O(gate195inter6));
  inv1  gate1030(.a(G590), .O(gate195inter7));
  inv1  gate1031(.a(G591), .O(gate195inter8));
  nand2 gate1032(.a(gate195inter8), .b(gate195inter7), .O(gate195inter9));
  nand2 gate1033(.a(s_69), .b(gate195inter3), .O(gate195inter10));
  nor2  gate1034(.a(gate195inter10), .b(gate195inter9), .O(gate195inter11));
  nor2  gate1035(.a(gate195inter11), .b(gate195inter6), .O(gate195inter12));
  nand2 gate1036(.a(gate195inter12), .b(gate195inter1), .O(G648));
nand2 gate196( .a(G592), .b(G593), .O(G651) );
nand2 gate197( .a(G594), .b(G595), .O(G654) );

  xor2  gate813(.a(G597), .b(G596), .O(gate198inter0));
  nand2 gate814(.a(gate198inter0), .b(s_38), .O(gate198inter1));
  and2  gate815(.a(G597), .b(G596), .O(gate198inter2));
  inv1  gate816(.a(s_38), .O(gate198inter3));
  inv1  gate817(.a(s_39), .O(gate198inter4));
  nand2 gate818(.a(gate198inter4), .b(gate198inter3), .O(gate198inter5));
  nor2  gate819(.a(gate198inter5), .b(gate198inter2), .O(gate198inter6));
  inv1  gate820(.a(G596), .O(gate198inter7));
  inv1  gate821(.a(G597), .O(gate198inter8));
  nand2 gate822(.a(gate198inter8), .b(gate198inter7), .O(gate198inter9));
  nand2 gate823(.a(s_39), .b(gate198inter3), .O(gate198inter10));
  nor2  gate824(.a(gate198inter10), .b(gate198inter9), .O(gate198inter11));
  nor2  gate825(.a(gate198inter11), .b(gate198inter6), .O(gate198inter12));
  nand2 gate826(.a(gate198inter12), .b(gate198inter1), .O(G657));
nand2 gate199( .a(G598), .b(G599), .O(G660) );

  xor2  gate617(.a(G601), .b(G600), .O(gate200inter0));
  nand2 gate618(.a(gate200inter0), .b(s_10), .O(gate200inter1));
  and2  gate619(.a(G601), .b(G600), .O(gate200inter2));
  inv1  gate620(.a(s_10), .O(gate200inter3));
  inv1  gate621(.a(s_11), .O(gate200inter4));
  nand2 gate622(.a(gate200inter4), .b(gate200inter3), .O(gate200inter5));
  nor2  gate623(.a(gate200inter5), .b(gate200inter2), .O(gate200inter6));
  inv1  gate624(.a(G600), .O(gate200inter7));
  inv1  gate625(.a(G601), .O(gate200inter8));
  nand2 gate626(.a(gate200inter8), .b(gate200inter7), .O(gate200inter9));
  nand2 gate627(.a(s_11), .b(gate200inter3), .O(gate200inter10));
  nor2  gate628(.a(gate200inter10), .b(gate200inter9), .O(gate200inter11));
  nor2  gate629(.a(gate200inter11), .b(gate200inter6), .O(gate200inter12));
  nand2 gate630(.a(gate200inter12), .b(gate200inter1), .O(G663));
nand2 gate201( .a(G602), .b(G607), .O(G666) );
nand2 gate202( .a(G612), .b(G617), .O(G669) );

  xor2  gate1037(.a(G612), .b(G602), .O(gate203inter0));
  nand2 gate1038(.a(gate203inter0), .b(s_70), .O(gate203inter1));
  and2  gate1039(.a(G612), .b(G602), .O(gate203inter2));
  inv1  gate1040(.a(s_70), .O(gate203inter3));
  inv1  gate1041(.a(s_71), .O(gate203inter4));
  nand2 gate1042(.a(gate203inter4), .b(gate203inter3), .O(gate203inter5));
  nor2  gate1043(.a(gate203inter5), .b(gate203inter2), .O(gate203inter6));
  inv1  gate1044(.a(G602), .O(gate203inter7));
  inv1  gate1045(.a(G612), .O(gate203inter8));
  nand2 gate1046(.a(gate203inter8), .b(gate203inter7), .O(gate203inter9));
  nand2 gate1047(.a(s_71), .b(gate203inter3), .O(gate203inter10));
  nor2  gate1048(.a(gate203inter10), .b(gate203inter9), .O(gate203inter11));
  nor2  gate1049(.a(gate203inter11), .b(gate203inter6), .O(gate203inter12));
  nand2 gate1050(.a(gate203inter12), .b(gate203inter1), .O(G672));
nand2 gate204( .a(G607), .b(G617), .O(G675) );

  xor2  gate1065(.a(G627), .b(G622), .O(gate205inter0));
  nand2 gate1066(.a(gate205inter0), .b(s_74), .O(gate205inter1));
  and2  gate1067(.a(G627), .b(G622), .O(gate205inter2));
  inv1  gate1068(.a(s_74), .O(gate205inter3));
  inv1  gate1069(.a(s_75), .O(gate205inter4));
  nand2 gate1070(.a(gate205inter4), .b(gate205inter3), .O(gate205inter5));
  nor2  gate1071(.a(gate205inter5), .b(gate205inter2), .O(gate205inter6));
  inv1  gate1072(.a(G622), .O(gate205inter7));
  inv1  gate1073(.a(G627), .O(gate205inter8));
  nand2 gate1074(.a(gate205inter8), .b(gate205inter7), .O(gate205inter9));
  nand2 gate1075(.a(s_75), .b(gate205inter3), .O(gate205inter10));
  nor2  gate1076(.a(gate205inter10), .b(gate205inter9), .O(gate205inter11));
  nor2  gate1077(.a(gate205inter11), .b(gate205inter6), .O(gate205inter12));
  nand2 gate1078(.a(gate205inter12), .b(gate205inter1), .O(G678));
nand2 gate206( .a(G632), .b(G637), .O(G681) );
nand2 gate207( .a(G622), .b(G632), .O(G684) );
nand2 gate208( .a(G627), .b(G637), .O(G687) );
nand2 gate209( .a(G602), .b(G666), .O(G690) );
nand2 gate210( .a(G607), .b(G666), .O(G691) );
nand2 gate211( .a(G612), .b(G669), .O(G692) );
nand2 gate212( .a(G617), .b(G669), .O(G693) );
nand2 gate213( .a(G602), .b(G672), .O(G694) );
nand2 gate214( .a(G612), .b(G672), .O(G695) );
nand2 gate215( .a(G607), .b(G675), .O(G696) );

  xor2  gate1247(.a(G675), .b(G617), .O(gate216inter0));
  nand2 gate1248(.a(gate216inter0), .b(s_100), .O(gate216inter1));
  and2  gate1249(.a(G675), .b(G617), .O(gate216inter2));
  inv1  gate1250(.a(s_100), .O(gate216inter3));
  inv1  gate1251(.a(s_101), .O(gate216inter4));
  nand2 gate1252(.a(gate216inter4), .b(gate216inter3), .O(gate216inter5));
  nor2  gate1253(.a(gate216inter5), .b(gate216inter2), .O(gate216inter6));
  inv1  gate1254(.a(G617), .O(gate216inter7));
  inv1  gate1255(.a(G675), .O(gate216inter8));
  nand2 gate1256(.a(gate216inter8), .b(gate216inter7), .O(gate216inter9));
  nand2 gate1257(.a(s_101), .b(gate216inter3), .O(gate216inter10));
  nor2  gate1258(.a(gate216inter10), .b(gate216inter9), .O(gate216inter11));
  nor2  gate1259(.a(gate216inter11), .b(gate216inter6), .O(gate216inter12));
  nand2 gate1260(.a(gate216inter12), .b(gate216inter1), .O(G697));
nand2 gate217( .a(G622), .b(G678), .O(G698) );
nand2 gate218( .a(G627), .b(G678), .O(G699) );
nand2 gate219( .a(G632), .b(G681), .O(G700) );

  xor2  gate743(.a(G681), .b(G637), .O(gate220inter0));
  nand2 gate744(.a(gate220inter0), .b(s_28), .O(gate220inter1));
  and2  gate745(.a(G681), .b(G637), .O(gate220inter2));
  inv1  gate746(.a(s_28), .O(gate220inter3));
  inv1  gate747(.a(s_29), .O(gate220inter4));
  nand2 gate748(.a(gate220inter4), .b(gate220inter3), .O(gate220inter5));
  nor2  gate749(.a(gate220inter5), .b(gate220inter2), .O(gate220inter6));
  inv1  gate750(.a(G637), .O(gate220inter7));
  inv1  gate751(.a(G681), .O(gate220inter8));
  nand2 gate752(.a(gate220inter8), .b(gate220inter7), .O(gate220inter9));
  nand2 gate753(.a(s_29), .b(gate220inter3), .O(gate220inter10));
  nor2  gate754(.a(gate220inter10), .b(gate220inter9), .O(gate220inter11));
  nor2  gate755(.a(gate220inter11), .b(gate220inter6), .O(gate220inter12));
  nand2 gate756(.a(gate220inter12), .b(gate220inter1), .O(G701));
nand2 gate221( .a(G622), .b(G684), .O(G702) );
nand2 gate222( .a(G632), .b(G684), .O(G703) );

  xor2  gate925(.a(G687), .b(G627), .O(gate223inter0));
  nand2 gate926(.a(gate223inter0), .b(s_54), .O(gate223inter1));
  and2  gate927(.a(G687), .b(G627), .O(gate223inter2));
  inv1  gate928(.a(s_54), .O(gate223inter3));
  inv1  gate929(.a(s_55), .O(gate223inter4));
  nand2 gate930(.a(gate223inter4), .b(gate223inter3), .O(gate223inter5));
  nor2  gate931(.a(gate223inter5), .b(gate223inter2), .O(gate223inter6));
  inv1  gate932(.a(G627), .O(gate223inter7));
  inv1  gate933(.a(G687), .O(gate223inter8));
  nand2 gate934(.a(gate223inter8), .b(gate223inter7), .O(gate223inter9));
  nand2 gate935(.a(s_55), .b(gate223inter3), .O(gate223inter10));
  nor2  gate936(.a(gate223inter10), .b(gate223inter9), .O(gate223inter11));
  nor2  gate937(.a(gate223inter11), .b(gate223inter6), .O(gate223inter12));
  nand2 gate938(.a(gate223inter12), .b(gate223inter1), .O(G704));

  xor2  gate1471(.a(G687), .b(G637), .O(gate224inter0));
  nand2 gate1472(.a(gate224inter0), .b(s_132), .O(gate224inter1));
  and2  gate1473(.a(G687), .b(G637), .O(gate224inter2));
  inv1  gate1474(.a(s_132), .O(gate224inter3));
  inv1  gate1475(.a(s_133), .O(gate224inter4));
  nand2 gate1476(.a(gate224inter4), .b(gate224inter3), .O(gate224inter5));
  nor2  gate1477(.a(gate224inter5), .b(gate224inter2), .O(gate224inter6));
  inv1  gate1478(.a(G637), .O(gate224inter7));
  inv1  gate1479(.a(G687), .O(gate224inter8));
  nand2 gate1480(.a(gate224inter8), .b(gate224inter7), .O(gate224inter9));
  nand2 gate1481(.a(s_133), .b(gate224inter3), .O(gate224inter10));
  nor2  gate1482(.a(gate224inter10), .b(gate224inter9), .O(gate224inter11));
  nor2  gate1483(.a(gate224inter11), .b(gate224inter6), .O(gate224inter12));
  nand2 gate1484(.a(gate224inter12), .b(gate224inter1), .O(G705));
nand2 gate225( .a(G690), .b(G691), .O(G706) );
nand2 gate226( .a(G692), .b(G693), .O(G709) );
nand2 gate227( .a(G694), .b(G695), .O(G712) );
nand2 gate228( .a(G696), .b(G697), .O(G715) );
nand2 gate229( .a(G698), .b(G699), .O(G718) );
nand2 gate230( .a(G700), .b(G701), .O(G721) );
nand2 gate231( .a(G702), .b(G703), .O(G724) );

  xor2  gate1345(.a(G705), .b(G704), .O(gate232inter0));
  nand2 gate1346(.a(gate232inter0), .b(s_114), .O(gate232inter1));
  and2  gate1347(.a(G705), .b(G704), .O(gate232inter2));
  inv1  gate1348(.a(s_114), .O(gate232inter3));
  inv1  gate1349(.a(s_115), .O(gate232inter4));
  nand2 gate1350(.a(gate232inter4), .b(gate232inter3), .O(gate232inter5));
  nor2  gate1351(.a(gate232inter5), .b(gate232inter2), .O(gate232inter6));
  inv1  gate1352(.a(G704), .O(gate232inter7));
  inv1  gate1353(.a(G705), .O(gate232inter8));
  nand2 gate1354(.a(gate232inter8), .b(gate232inter7), .O(gate232inter9));
  nand2 gate1355(.a(s_115), .b(gate232inter3), .O(gate232inter10));
  nor2  gate1356(.a(gate232inter10), .b(gate232inter9), .O(gate232inter11));
  nor2  gate1357(.a(gate232inter11), .b(gate232inter6), .O(gate232inter12));
  nand2 gate1358(.a(gate232inter12), .b(gate232inter1), .O(G727));
nand2 gate233( .a(G242), .b(G718), .O(G730) );
nand2 gate234( .a(G245), .b(G721), .O(G733) );
nand2 gate235( .a(G248), .b(G724), .O(G736) );
nand2 gate236( .a(G251), .b(G727), .O(G739) );

  xor2  gate785(.a(G706), .b(G254), .O(gate237inter0));
  nand2 gate786(.a(gate237inter0), .b(s_34), .O(gate237inter1));
  and2  gate787(.a(G706), .b(G254), .O(gate237inter2));
  inv1  gate788(.a(s_34), .O(gate237inter3));
  inv1  gate789(.a(s_35), .O(gate237inter4));
  nand2 gate790(.a(gate237inter4), .b(gate237inter3), .O(gate237inter5));
  nor2  gate791(.a(gate237inter5), .b(gate237inter2), .O(gate237inter6));
  inv1  gate792(.a(G254), .O(gate237inter7));
  inv1  gate793(.a(G706), .O(gate237inter8));
  nand2 gate794(.a(gate237inter8), .b(gate237inter7), .O(gate237inter9));
  nand2 gate795(.a(s_35), .b(gate237inter3), .O(gate237inter10));
  nor2  gate796(.a(gate237inter10), .b(gate237inter9), .O(gate237inter11));
  nor2  gate797(.a(gate237inter11), .b(gate237inter6), .O(gate237inter12));
  nand2 gate798(.a(gate237inter12), .b(gate237inter1), .O(G742));
nand2 gate238( .a(G257), .b(G709), .O(G745) );

  xor2  gate869(.a(G712), .b(G260), .O(gate239inter0));
  nand2 gate870(.a(gate239inter0), .b(s_46), .O(gate239inter1));
  and2  gate871(.a(G712), .b(G260), .O(gate239inter2));
  inv1  gate872(.a(s_46), .O(gate239inter3));
  inv1  gate873(.a(s_47), .O(gate239inter4));
  nand2 gate874(.a(gate239inter4), .b(gate239inter3), .O(gate239inter5));
  nor2  gate875(.a(gate239inter5), .b(gate239inter2), .O(gate239inter6));
  inv1  gate876(.a(G260), .O(gate239inter7));
  inv1  gate877(.a(G712), .O(gate239inter8));
  nand2 gate878(.a(gate239inter8), .b(gate239inter7), .O(gate239inter9));
  nand2 gate879(.a(s_47), .b(gate239inter3), .O(gate239inter10));
  nor2  gate880(.a(gate239inter10), .b(gate239inter9), .O(gate239inter11));
  nor2  gate881(.a(gate239inter11), .b(gate239inter6), .O(gate239inter12));
  nand2 gate882(.a(gate239inter12), .b(gate239inter1), .O(G748));

  xor2  gate953(.a(G715), .b(G263), .O(gate240inter0));
  nand2 gate954(.a(gate240inter0), .b(s_58), .O(gate240inter1));
  and2  gate955(.a(G715), .b(G263), .O(gate240inter2));
  inv1  gate956(.a(s_58), .O(gate240inter3));
  inv1  gate957(.a(s_59), .O(gate240inter4));
  nand2 gate958(.a(gate240inter4), .b(gate240inter3), .O(gate240inter5));
  nor2  gate959(.a(gate240inter5), .b(gate240inter2), .O(gate240inter6));
  inv1  gate960(.a(G263), .O(gate240inter7));
  inv1  gate961(.a(G715), .O(gate240inter8));
  nand2 gate962(.a(gate240inter8), .b(gate240inter7), .O(gate240inter9));
  nand2 gate963(.a(s_59), .b(gate240inter3), .O(gate240inter10));
  nor2  gate964(.a(gate240inter10), .b(gate240inter9), .O(gate240inter11));
  nor2  gate965(.a(gate240inter11), .b(gate240inter6), .O(gate240inter12));
  nand2 gate966(.a(gate240inter12), .b(gate240inter1), .O(G751));
nand2 gate241( .a(G242), .b(G730), .O(G754) );
nand2 gate242( .a(G718), .b(G730), .O(G755) );

  xor2  gate911(.a(G733), .b(G245), .O(gate243inter0));
  nand2 gate912(.a(gate243inter0), .b(s_52), .O(gate243inter1));
  and2  gate913(.a(G733), .b(G245), .O(gate243inter2));
  inv1  gate914(.a(s_52), .O(gate243inter3));
  inv1  gate915(.a(s_53), .O(gate243inter4));
  nand2 gate916(.a(gate243inter4), .b(gate243inter3), .O(gate243inter5));
  nor2  gate917(.a(gate243inter5), .b(gate243inter2), .O(gate243inter6));
  inv1  gate918(.a(G245), .O(gate243inter7));
  inv1  gate919(.a(G733), .O(gate243inter8));
  nand2 gate920(.a(gate243inter8), .b(gate243inter7), .O(gate243inter9));
  nand2 gate921(.a(s_53), .b(gate243inter3), .O(gate243inter10));
  nor2  gate922(.a(gate243inter10), .b(gate243inter9), .O(gate243inter11));
  nor2  gate923(.a(gate243inter11), .b(gate243inter6), .O(gate243inter12));
  nand2 gate924(.a(gate243inter12), .b(gate243inter1), .O(G756));

  xor2  gate1709(.a(G733), .b(G721), .O(gate244inter0));
  nand2 gate1710(.a(gate244inter0), .b(s_166), .O(gate244inter1));
  and2  gate1711(.a(G733), .b(G721), .O(gate244inter2));
  inv1  gate1712(.a(s_166), .O(gate244inter3));
  inv1  gate1713(.a(s_167), .O(gate244inter4));
  nand2 gate1714(.a(gate244inter4), .b(gate244inter3), .O(gate244inter5));
  nor2  gate1715(.a(gate244inter5), .b(gate244inter2), .O(gate244inter6));
  inv1  gate1716(.a(G721), .O(gate244inter7));
  inv1  gate1717(.a(G733), .O(gate244inter8));
  nand2 gate1718(.a(gate244inter8), .b(gate244inter7), .O(gate244inter9));
  nand2 gate1719(.a(s_167), .b(gate244inter3), .O(gate244inter10));
  nor2  gate1720(.a(gate244inter10), .b(gate244inter9), .O(gate244inter11));
  nor2  gate1721(.a(gate244inter11), .b(gate244inter6), .O(gate244inter12));
  nand2 gate1722(.a(gate244inter12), .b(gate244inter1), .O(G757));

  xor2  gate841(.a(G736), .b(G248), .O(gate245inter0));
  nand2 gate842(.a(gate245inter0), .b(s_42), .O(gate245inter1));
  and2  gate843(.a(G736), .b(G248), .O(gate245inter2));
  inv1  gate844(.a(s_42), .O(gate245inter3));
  inv1  gate845(.a(s_43), .O(gate245inter4));
  nand2 gate846(.a(gate245inter4), .b(gate245inter3), .O(gate245inter5));
  nor2  gate847(.a(gate245inter5), .b(gate245inter2), .O(gate245inter6));
  inv1  gate848(.a(G248), .O(gate245inter7));
  inv1  gate849(.a(G736), .O(gate245inter8));
  nand2 gate850(.a(gate245inter8), .b(gate245inter7), .O(gate245inter9));
  nand2 gate851(.a(s_43), .b(gate245inter3), .O(gate245inter10));
  nor2  gate852(.a(gate245inter10), .b(gate245inter9), .O(gate245inter11));
  nor2  gate853(.a(gate245inter11), .b(gate245inter6), .O(gate245inter12));
  nand2 gate854(.a(gate245inter12), .b(gate245inter1), .O(G758));

  xor2  gate799(.a(G736), .b(G724), .O(gate246inter0));
  nand2 gate800(.a(gate246inter0), .b(s_36), .O(gate246inter1));
  and2  gate801(.a(G736), .b(G724), .O(gate246inter2));
  inv1  gate802(.a(s_36), .O(gate246inter3));
  inv1  gate803(.a(s_37), .O(gate246inter4));
  nand2 gate804(.a(gate246inter4), .b(gate246inter3), .O(gate246inter5));
  nor2  gate805(.a(gate246inter5), .b(gate246inter2), .O(gate246inter6));
  inv1  gate806(.a(G724), .O(gate246inter7));
  inv1  gate807(.a(G736), .O(gate246inter8));
  nand2 gate808(.a(gate246inter8), .b(gate246inter7), .O(gate246inter9));
  nand2 gate809(.a(s_37), .b(gate246inter3), .O(gate246inter10));
  nor2  gate810(.a(gate246inter10), .b(gate246inter9), .O(gate246inter11));
  nor2  gate811(.a(gate246inter11), .b(gate246inter6), .O(gate246inter12));
  nand2 gate812(.a(gate246inter12), .b(gate246inter1), .O(G759));
nand2 gate247( .a(G251), .b(G739), .O(G760) );
nand2 gate248( .a(G727), .b(G739), .O(G761) );
nand2 gate249( .a(G254), .b(G742), .O(G762) );
nand2 gate250( .a(G706), .b(G742), .O(G763) );
nand2 gate251( .a(G257), .b(G745), .O(G764) );
nand2 gate252( .a(G709), .b(G745), .O(G765) );
nand2 gate253( .a(G260), .b(G748), .O(G766) );
nand2 gate254( .a(G712), .b(G748), .O(G767) );

  xor2  gate1611(.a(G751), .b(G263), .O(gate255inter0));
  nand2 gate1612(.a(gate255inter0), .b(s_152), .O(gate255inter1));
  and2  gate1613(.a(G751), .b(G263), .O(gate255inter2));
  inv1  gate1614(.a(s_152), .O(gate255inter3));
  inv1  gate1615(.a(s_153), .O(gate255inter4));
  nand2 gate1616(.a(gate255inter4), .b(gate255inter3), .O(gate255inter5));
  nor2  gate1617(.a(gate255inter5), .b(gate255inter2), .O(gate255inter6));
  inv1  gate1618(.a(G263), .O(gate255inter7));
  inv1  gate1619(.a(G751), .O(gate255inter8));
  nand2 gate1620(.a(gate255inter8), .b(gate255inter7), .O(gate255inter9));
  nand2 gate1621(.a(s_153), .b(gate255inter3), .O(gate255inter10));
  nor2  gate1622(.a(gate255inter10), .b(gate255inter9), .O(gate255inter11));
  nor2  gate1623(.a(gate255inter11), .b(gate255inter6), .O(gate255inter12));
  nand2 gate1624(.a(gate255inter12), .b(gate255inter1), .O(G768));
nand2 gate256( .a(G715), .b(G751), .O(G769) );
nand2 gate257( .a(G754), .b(G755), .O(G770) );
nand2 gate258( .a(G756), .b(G757), .O(G773) );

  xor2  gate631(.a(G759), .b(G758), .O(gate259inter0));
  nand2 gate632(.a(gate259inter0), .b(s_12), .O(gate259inter1));
  and2  gate633(.a(G759), .b(G758), .O(gate259inter2));
  inv1  gate634(.a(s_12), .O(gate259inter3));
  inv1  gate635(.a(s_13), .O(gate259inter4));
  nand2 gate636(.a(gate259inter4), .b(gate259inter3), .O(gate259inter5));
  nor2  gate637(.a(gate259inter5), .b(gate259inter2), .O(gate259inter6));
  inv1  gate638(.a(G758), .O(gate259inter7));
  inv1  gate639(.a(G759), .O(gate259inter8));
  nand2 gate640(.a(gate259inter8), .b(gate259inter7), .O(gate259inter9));
  nand2 gate641(.a(s_13), .b(gate259inter3), .O(gate259inter10));
  nor2  gate642(.a(gate259inter10), .b(gate259inter9), .O(gate259inter11));
  nor2  gate643(.a(gate259inter11), .b(gate259inter6), .O(gate259inter12));
  nand2 gate644(.a(gate259inter12), .b(gate259inter1), .O(G776));
nand2 gate260( .a(G760), .b(G761), .O(G779) );
nand2 gate261( .a(G762), .b(G763), .O(G782) );

  xor2  gate1275(.a(G765), .b(G764), .O(gate262inter0));
  nand2 gate1276(.a(gate262inter0), .b(s_104), .O(gate262inter1));
  and2  gate1277(.a(G765), .b(G764), .O(gate262inter2));
  inv1  gate1278(.a(s_104), .O(gate262inter3));
  inv1  gate1279(.a(s_105), .O(gate262inter4));
  nand2 gate1280(.a(gate262inter4), .b(gate262inter3), .O(gate262inter5));
  nor2  gate1281(.a(gate262inter5), .b(gate262inter2), .O(gate262inter6));
  inv1  gate1282(.a(G764), .O(gate262inter7));
  inv1  gate1283(.a(G765), .O(gate262inter8));
  nand2 gate1284(.a(gate262inter8), .b(gate262inter7), .O(gate262inter9));
  nand2 gate1285(.a(s_105), .b(gate262inter3), .O(gate262inter10));
  nor2  gate1286(.a(gate262inter10), .b(gate262inter9), .O(gate262inter11));
  nor2  gate1287(.a(gate262inter11), .b(gate262inter6), .O(gate262inter12));
  nand2 gate1288(.a(gate262inter12), .b(gate262inter1), .O(G785));
nand2 gate263( .a(G766), .b(G767), .O(G788) );
nand2 gate264( .a(G768), .b(G769), .O(G791) );
nand2 gate265( .a(G642), .b(G770), .O(G794) );
nand2 gate266( .a(G645), .b(G773), .O(G797) );
nand2 gate267( .a(G648), .b(G776), .O(G800) );
nand2 gate268( .a(G651), .b(G779), .O(G803) );
nand2 gate269( .a(G654), .b(G782), .O(G806) );
nand2 gate270( .a(G657), .b(G785), .O(G809) );

  xor2  gate547(.a(G788), .b(G660), .O(gate271inter0));
  nand2 gate548(.a(gate271inter0), .b(s_0), .O(gate271inter1));
  and2  gate549(.a(G788), .b(G660), .O(gate271inter2));
  inv1  gate550(.a(s_0), .O(gate271inter3));
  inv1  gate551(.a(s_1), .O(gate271inter4));
  nand2 gate552(.a(gate271inter4), .b(gate271inter3), .O(gate271inter5));
  nor2  gate553(.a(gate271inter5), .b(gate271inter2), .O(gate271inter6));
  inv1  gate554(.a(G660), .O(gate271inter7));
  inv1  gate555(.a(G788), .O(gate271inter8));
  nand2 gate556(.a(gate271inter8), .b(gate271inter7), .O(gate271inter9));
  nand2 gate557(.a(s_1), .b(gate271inter3), .O(gate271inter10));
  nor2  gate558(.a(gate271inter10), .b(gate271inter9), .O(gate271inter11));
  nor2  gate559(.a(gate271inter11), .b(gate271inter6), .O(gate271inter12));
  nand2 gate560(.a(gate271inter12), .b(gate271inter1), .O(G812));
nand2 gate272( .a(G663), .b(G791), .O(G815) );
nand2 gate273( .a(G642), .b(G794), .O(G818) );
nand2 gate274( .a(G770), .b(G794), .O(G819) );
nand2 gate275( .a(G645), .b(G797), .O(G820) );
nand2 gate276( .a(G773), .b(G797), .O(G821) );
nand2 gate277( .a(G648), .b(G800), .O(G822) );
nand2 gate278( .a(G776), .b(G800), .O(G823) );
nand2 gate279( .a(G651), .b(G803), .O(G824) );
nand2 gate280( .a(G779), .b(G803), .O(G825) );
nand2 gate281( .a(G654), .b(G806), .O(G826) );
nand2 gate282( .a(G782), .b(G806), .O(G827) );

  xor2  gate1639(.a(G809), .b(G657), .O(gate283inter0));
  nand2 gate1640(.a(gate283inter0), .b(s_156), .O(gate283inter1));
  and2  gate1641(.a(G809), .b(G657), .O(gate283inter2));
  inv1  gate1642(.a(s_156), .O(gate283inter3));
  inv1  gate1643(.a(s_157), .O(gate283inter4));
  nand2 gate1644(.a(gate283inter4), .b(gate283inter3), .O(gate283inter5));
  nor2  gate1645(.a(gate283inter5), .b(gate283inter2), .O(gate283inter6));
  inv1  gate1646(.a(G657), .O(gate283inter7));
  inv1  gate1647(.a(G809), .O(gate283inter8));
  nand2 gate1648(.a(gate283inter8), .b(gate283inter7), .O(gate283inter9));
  nand2 gate1649(.a(s_157), .b(gate283inter3), .O(gate283inter10));
  nor2  gate1650(.a(gate283inter10), .b(gate283inter9), .O(gate283inter11));
  nor2  gate1651(.a(gate283inter11), .b(gate283inter6), .O(gate283inter12));
  nand2 gate1652(.a(gate283inter12), .b(gate283inter1), .O(G828));
nand2 gate284( .a(G785), .b(G809), .O(G829) );

  xor2  gate701(.a(G812), .b(G660), .O(gate285inter0));
  nand2 gate702(.a(gate285inter0), .b(s_22), .O(gate285inter1));
  and2  gate703(.a(G812), .b(G660), .O(gate285inter2));
  inv1  gate704(.a(s_22), .O(gate285inter3));
  inv1  gate705(.a(s_23), .O(gate285inter4));
  nand2 gate706(.a(gate285inter4), .b(gate285inter3), .O(gate285inter5));
  nor2  gate707(.a(gate285inter5), .b(gate285inter2), .O(gate285inter6));
  inv1  gate708(.a(G660), .O(gate285inter7));
  inv1  gate709(.a(G812), .O(gate285inter8));
  nand2 gate710(.a(gate285inter8), .b(gate285inter7), .O(gate285inter9));
  nand2 gate711(.a(s_23), .b(gate285inter3), .O(gate285inter10));
  nor2  gate712(.a(gate285inter10), .b(gate285inter9), .O(gate285inter11));
  nor2  gate713(.a(gate285inter11), .b(gate285inter6), .O(gate285inter12));
  nand2 gate714(.a(gate285inter12), .b(gate285inter1), .O(G830));
nand2 gate286( .a(G788), .b(G812), .O(G831) );
nand2 gate287( .a(G663), .b(G815), .O(G832) );
nand2 gate288( .a(G791), .b(G815), .O(G833) );
nand2 gate289( .a(G818), .b(G819), .O(G834) );
nand2 gate290( .a(G820), .b(G821), .O(G847) );
nand2 gate291( .a(G822), .b(G823), .O(G860) );
nand2 gate292( .a(G824), .b(G825), .O(G873) );

  xor2  gate1317(.a(G829), .b(G828), .O(gate293inter0));
  nand2 gate1318(.a(gate293inter0), .b(s_110), .O(gate293inter1));
  and2  gate1319(.a(G829), .b(G828), .O(gate293inter2));
  inv1  gate1320(.a(s_110), .O(gate293inter3));
  inv1  gate1321(.a(s_111), .O(gate293inter4));
  nand2 gate1322(.a(gate293inter4), .b(gate293inter3), .O(gate293inter5));
  nor2  gate1323(.a(gate293inter5), .b(gate293inter2), .O(gate293inter6));
  inv1  gate1324(.a(G828), .O(gate293inter7));
  inv1  gate1325(.a(G829), .O(gate293inter8));
  nand2 gate1326(.a(gate293inter8), .b(gate293inter7), .O(gate293inter9));
  nand2 gate1327(.a(s_111), .b(gate293inter3), .O(gate293inter10));
  nor2  gate1328(.a(gate293inter10), .b(gate293inter9), .O(gate293inter11));
  nor2  gate1329(.a(gate293inter11), .b(gate293inter6), .O(gate293inter12));
  nand2 gate1330(.a(gate293inter12), .b(gate293inter1), .O(G886));
nand2 gate294( .a(G832), .b(G833), .O(G899) );
nand2 gate295( .a(G830), .b(G831), .O(G912) );
nand2 gate296( .a(G826), .b(G827), .O(G925) );
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );
nand2 gate387( .a(G1), .b(G1036), .O(G1132) );
nand2 gate388( .a(G2), .b(G1039), .O(G1135) );
nand2 gate389( .a(G3), .b(G1042), .O(G1138) );
nand2 gate390( .a(G4), .b(G1045), .O(G1141) );
nand2 gate391( .a(G5), .b(G1048), .O(G1144) );

  xor2  gate1541(.a(G1051), .b(G6), .O(gate392inter0));
  nand2 gate1542(.a(gate392inter0), .b(s_142), .O(gate392inter1));
  and2  gate1543(.a(G1051), .b(G6), .O(gate392inter2));
  inv1  gate1544(.a(s_142), .O(gate392inter3));
  inv1  gate1545(.a(s_143), .O(gate392inter4));
  nand2 gate1546(.a(gate392inter4), .b(gate392inter3), .O(gate392inter5));
  nor2  gate1547(.a(gate392inter5), .b(gate392inter2), .O(gate392inter6));
  inv1  gate1548(.a(G6), .O(gate392inter7));
  inv1  gate1549(.a(G1051), .O(gate392inter8));
  nand2 gate1550(.a(gate392inter8), .b(gate392inter7), .O(gate392inter9));
  nand2 gate1551(.a(s_143), .b(gate392inter3), .O(gate392inter10));
  nor2  gate1552(.a(gate392inter10), .b(gate392inter9), .O(gate392inter11));
  nor2  gate1553(.a(gate392inter11), .b(gate392inter6), .O(gate392inter12));
  nand2 gate1554(.a(gate392inter12), .b(gate392inter1), .O(G1147));

  xor2  gate757(.a(G1054), .b(G7), .O(gate393inter0));
  nand2 gate758(.a(gate393inter0), .b(s_30), .O(gate393inter1));
  and2  gate759(.a(G1054), .b(G7), .O(gate393inter2));
  inv1  gate760(.a(s_30), .O(gate393inter3));
  inv1  gate761(.a(s_31), .O(gate393inter4));
  nand2 gate762(.a(gate393inter4), .b(gate393inter3), .O(gate393inter5));
  nor2  gate763(.a(gate393inter5), .b(gate393inter2), .O(gate393inter6));
  inv1  gate764(.a(G7), .O(gate393inter7));
  inv1  gate765(.a(G1054), .O(gate393inter8));
  nand2 gate766(.a(gate393inter8), .b(gate393inter7), .O(gate393inter9));
  nand2 gate767(.a(s_31), .b(gate393inter3), .O(gate393inter10));
  nor2  gate768(.a(gate393inter10), .b(gate393inter9), .O(gate393inter11));
  nor2  gate769(.a(gate393inter11), .b(gate393inter6), .O(gate393inter12));
  nand2 gate770(.a(gate393inter12), .b(gate393inter1), .O(G1150));
nand2 gate394( .a(G8), .b(G1057), .O(G1153) );

  xor2  gate1191(.a(G1060), .b(G9), .O(gate395inter0));
  nand2 gate1192(.a(gate395inter0), .b(s_92), .O(gate395inter1));
  and2  gate1193(.a(G1060), .b(G9), .O(gate395inter2));
  inv1  gate1194(.a(s_92), .O(gate395inter3));
  inv1  gate1195(.a(s_93), .O(gate395inter4));
  nand2 gate1196(.a(gate395inter4), .b(gate395inter3), .O(gate395inter5));
  nor2  gate1197(.a(gate395inter5), .b(gate395inter2), .O(gate395inter6));
  inv1  gate1198(.a(G9), .O(gate395inter7));
  inv1  gate1199(.a(G1060), .O(gate395inter8));
  nand2 gate1200(.a(gate395inter8), .b(gate395inter7), .O(gate395inter9));
  nand2 gate1201(.a(s_93), .b(gate395inter3), .O(gate395inter10));
  nor2  gate1202(.a(gate395inter10), .b(gate395inter9), .O(gate395inter11));
  nor2  gate1203(.a(gate395inter11), .b(gate395inter6), .O(gate395inter12));
  nand2 gate1204(.a(gate395inter12), .b(gate395inter1), .O(G1156));
nand2 gate396( .a(G10), .b(G1063), .O(G1159) );
nand2 gate397( .a(G11), .b(G1066), .O(G1162) );
nand2 gate398( .a(G12), .b(G1069), .O(G1165) );

  xor2  gate1415(.a(G1072), .b(G13), .O(gate399inter0));
  nand2 gate1416(.a(gate399inter0), .b(s_124), .O(gate399inter1));
  and2  gate1417(.a(G1072), .b(G13), .O(gate399inter2));
  inv1  gate1418(.a(s_124), .O(gate399inter3));
  inv1  gate1419(.a(s_125), .O(gate399inter4));
  nand2 gate1420(.a(gate399inter4), .b(gate399inter3), .O(gate399inter5));
  nor2  gate1421(.a(gate399inter5), .b(gate399inter2), .O(gate399inter6));
  inv1  gate1422(.a(G13), .O(gate399inter7));
  inv1  gate1423(.a(G1072), .O(gate399inter8));
  nand2 gate1424(.a(gate399inter8), .b(gate399inter7), .O(gate399inter9));
  nand2 gate1425(.a(s_125), .b(gate399inter3), .O(gate399inter10));
  nor2  gate1426(.a(gate399inter10), .b(gate399inter9), .O(gate399inter11));
  nor2  gate1427(.a(gate399inter11), .b(gate399inter6), .O(gate399inter12));
  nand2 gate1428(.a(gate399inter12), .b(gate399inter1), .O(G1168));
nand2 gate400( .a(G14), .b(G1075), .O(G1171) );
nand2 gate401( .a(G15), .b(G1078), .O(G1174) );
nand2 gate402( .a(G16), .b(G1081), .O(G1177) );
nand2 gate403( .a(G17), .b(G1084), .O(G1180) );
nand2 gate404( .a(G18), .b(G1087), .O(G1183) );
nand2 gate405( .a(G19), .b(G1090), .O(G1186) );
nand2 gate406( .a(G20), .b(G1093), .O(G1189) );
nand2 gate407( .a(G21), .b(G1096), .O(G1192) );
nand2 gate408( .a(G22), .b(G1099), .O(G1195) );
nand2 gate409( .a(G23), .b(G1102), .O(G1198) );

  xor2  gate715(.a(G1105), .b(G24), .O(gate410inter0));
  nand2 gate716(.a(gate410inter0), .b(s_24), .O(gate410inter1));
  and2  gate717(.a(G1105), .b(G24), .O(gate410inter2));
  inv1  gate718(.a(s_24), .O(gate410inter3));
  inv1  gate719(.a(s_25), .O(gate410inter4));
  nand2 gate720(.a(gate410inter4), .b(gate410inter3), .O(gate410inter5));
  nor2  gate721(.a(gate410inter5), .b(gate410inter2), .O(gate410inter6));
  inv1  gate722(.a(G24), .O(gate410inter7));
  inv1  gate723(.a(G1105), .O(gate410inter8));
  nand2 gate724(.a(gate410inter8), .b(gate410inter7), .O(gate410inter9));
  nand2 gate725(.a(s_25), .b(gate410inter3), .O(gate410inter10));
  nor2  gate726(.a(gate410inter10), .b(gate410inter9), .O(gate410inter11));
  nor2  gate727(.a(gate410inter11), .b(gate410inter6), .O(gate410inter12));
  nand2 gate728(.a(gate410inter12), .b(gate410inter1), .O(G1201));
nand2 gate411( .a(G25), .b(G1108), .O(G1204) );
nand2 gate412( .a(G26), .b(G1111), .O(G1207) );
nand2 gate413( .a(G27), .b(G1114), .O(G1210) );
nand2 gate414( .a(G28), .b(G1117), .O(G1213) );
nand2 gate415( .a(G29), .b(G1120), .O(G1216) );
nand2 gate416( .a(G30), .b(G1123), .O(G1219) );
nand2 gate417( .a(G31), .b(G1126), .O(G1222) );
nand2 gate418( .a(G32), .b(G1129), .O(G1225) );

  xor2  gate1863(.a(G1132), .b(G1), .O(gate419inter0));
  nand2 gate1864(.a(gate419inter0), .b(s_188), .O(gate419inter1));
  and2  gate1865(.a(G1132), .b(G1), .O(gate419inter2));
  inv1  gate1866(.a(s_188), .O(gate419inter3));
  inv1  gate1867(.a(s_189), .O(gate419inter4));
  nand2 gate1868(.a(gate419inter4), .b(gate419inter3), .O(gate419inter5));
  nor2  gate1869(.a(gate419inter5), .b(gate419inter2), .O(gate419inter6));
  inv1  gate1870(.a(G1), .O(gate419inter7));
  inv1  gate1871(.a(G1132), .O(gate419inter8));
  nand2 gate1872(.a(gate419inter8), .b(gate419inter7), .O(gate419inter9));
  nand2 gate1873(.a(s_189), .b(gate419inter3), .O(gate419inter10));
  nor2  gate1874(.a(gate419inter10), .b(gate419inter9), .O(gate419inter11));
  nor2  gate1875(.a(gate419inter11), .b(gate419inter6), .O(gate419inter12));
  nand2 gate1876(.a(gate419inter12), .b(gate419inter1), .O(G1228));

  xor2  gate1751(.a(G1132), .b(G1036), .O(gate420inter0));
  nand2 gate1752(.a(gate420inter0), .b(s_172), .O(gate420inter1));
  and2  gate1753(.a(G1132), .b(G1036), .O(gate420inter2));
  inv1  gate1754(.a(s_172), .O(gate420inter3));
  inv1  gate1755(.a(s_173), .O(gate420inter4));
  nand2 gate1756(.a(gate420inter4), .b(gate420inter3), .O(gate420inter5));
  nor2  gate1757(.a(gate420inter5), .b(gate420inter2), .O(gate420inter6));
  inv1  gate1758(.a(G1036), .O(gate420inter7));
  inv1  gate1759(.a(G1132), .O(gate420inter8));
  nand2 gate1760(.a(gate420inter8), .b(gate420inter7), .O(gate420inter9));
  nand2 gate1761(.a(s_173), .b(gate420inter3), .O(gate420inter10));
  nor2  gate1762(.a(gate420inter10), .b(gate420inter9), .O(gate420inter11));
  nor2  gate1763(.a(gate420inter11), .b(gate420inter6), .O(gate420inter12));
  nand2 gate1764(.a(gate420inter12), .b(gate420inter1), .O(G1229));
nand2 gate421( .a(G2), .b(G1135), .O(G1230) );
nand2 gate422( .a(G1039), .b(G1135), .O(G1231) );
nand2 gate423( .a(G3), .b(G1138), .O(G1232) );
nand2 gate424( .a(G1042), .b(G1138), .O(G1233) );
nand2 gate425( .a(G4), .b(G1141), .O(G1234) );
nand2 gate426( .a(G1045), .b(G1141), .O(G1235) );
nand2 gate427( .a(G5), .b(G1144), .O(G1236) );
nand2 gate428( .a(G1048), .b(G1144), .O(G1237) );
nand2 gate429( .a(G6), .b(G1147), .O(G1238) );

  xor2  gate1359(.a(G1147), .b(G1051), .O(gate430inter0));
  nand2 gate1360(.a(gate430inter0), .b(s_116), .O(gate430inter1));
  and2  gate1361(.a(G1147), .b(G1051), .O(gate430inter2));
  inv1  gate1362(.a(s_116), .O(gate430inter3));
  inv1  gate1363(.a(s_117), .O(gate430inter4));
  nand2 gate1364(.a(gate430inter4), .b(gate430inter3), .O(gate430inter5));
  nor2  gate1365(.a(gate430inter5), .b(gate430inter2), .O(gate430inter6));
  inv1  gate1366(.a(G1051), .O(gate430inter7));
  inv1  gate1367(.a(G1147), .O(gate430inter8));
  nand2 gate1368(.a(gate430inter8), .b(gate430inter7), .O(gate430inter9));
  nand2 gate1369(.a(s_117), .b(gate430inter3), .O(gate430inter10));
  nor2  gate1370(.a(gate430inter10), .b(gate430inter9), .O(gate430inter11));
  nor2  gate1371(.a(gate430inter11), .b(gate430inter6), .O(gate430inter12));
  nand2 gate1372(.a(gate430inter12), .b(gate430inter1), .O(G1239));
nand2 gate431( .a(G7), .b(G1150), .O(G1240) );

  xor2  gate1779(.a(G1150), .b(G1054), .O(gate432inter0));
  nand2 gate1780(.a(gate432inter0), .b(s_176), .O(gate432inter1));
  and2  gate1781(.a(G1150), .b(G1054), .O(gate432inter2));
  inv1  gate1782(.a(s_176), .O(gate432inter3));
  inv1  gate1783(.a(s_177), .O(gate432inter4));
  nand2 gate1784(.a(gate432inter4), .b(gate432inter3), .O(gate432inter5));
  nor2  gate1785(.a(gate432inter5), .b(gate432inter2), .O(gate432inter6));
  inv1  gate1786(.a(G1054), .O(gate432inter7));
  inv1  gate1787(.a(G1150), .O(gate432inter8));
  nand2 gate1788(.a(gate432inter8), .b(gate432inter7), .O(gate432inter9));
  nand2 gate1789(.a(s_177), .b(gate432inter3), .O(gate432inter10));
  nor2  gate1790(.a(gate432inter10), .b(gate432inter9), .O(gate432inter11));
  nor2  gate1791(.a(gate432inter11), .b(gate432inter6), .O(gate432inter12));
  nand2 gate1792(.a(gate432inter12), .b(gate432inter1), .O(G1241));
nand2 gate433( .a(G8), .b(G1153), .O(G1242) );
nand2 gate434( .a(G1057), .b(G1153), .O(G1243) );
nand2 gate435( .a(G9), .b(G1156), .O(G1244) );
nand2 gate436( .a(G1060), .b(G1156), .O(G1245) );
nand2 gate437( .a(G10), .b(G1159), .O(G1246) );
nand2 gate438( .a(G1063), .b(G1159), .O(G1247) );
nand2 gate439( .a(G11), .b(G1162), .O(G1248) );
nand2 gate440( .a(G1066), .b(G1162), .O(G1249) );
nand2 gate441( .a(G12), .b(G1165), .O(G1250) );
nand2 gate442( .a(G1069), .b(G1165), .O(G1251) );

  xor2  gate1205(.a(G1168), .b(G13), .O(gate443inter0));
  nand2 gate1206(.a(gate443inter0), .b(s_94), .O(gate443inter1));
  and2  gate1207(.a(G1168), .b(G13), .O(gate443inter2));
  inv1  gate1208(.a(s_94), .O(gate443inter3));
  inv1  gate1209(.a(s_95), .O(gate443inter4));
  nand2 gate1210(.a(gate443inter4), .b(gate443inter3), .O(gate443inter5));
  nor2  gate1211(.a(gate443inter5), .b(gate443inter2), .O(gate443inter6));
  inv1  gate1212(.a(G13), .O(gate443inter7));
  inv1  gate1213(.a(G1168), .O(gate443inter8));
  nand2 gate1214(.a(gate443inter8), .b(gate443inter7), .O(gate443inter9));
  nand2 gate1215(.a(s_95), .b(gate443inter3), .O(gate443inter10));
  nor2  gate1216(.a(gate443inter10), .b(gate443inter9), .O(gate443inter11));
  nor2  gate1217(.a(gate443inter11), .b(gate443inter6), .O(gate443inter12));
  nand2 gate1218(.a(gate443inter12), .b(gate443inter1), .O(G1252));
nand2 gate444( .a(G1072), .b(G1168), .O(G1253) );
nand2 gate445( .a(G14), .b(G1171), .O(G1254) );

  xor2  gate967(.a(G1171), .b(G1075), .O(gate446inter0));
  nand2 gate968(.a(gate446inter0), .b(s_60), .O(gate446inter1));
  and2  gate969(.a(G1171), .b(G1075), .O(gate446inter2));
  inv1  gate970(.a(s_60), .O(gate446inter3));
  inv1  gate971(.a(s_61), .O(gate446inter4));
  nand2 gate972(.a(gate446inter4), .b(gate446inter3), .O(gate446inter5));
  nor2  gate973(.a(gate446inter5), .b(gate446inter2), .O(gate446inter6));
  inv1  gate974(.a(G1075), .O(gate446inter7));
  inv1  gate975(.a(G1171), .O(gate446inter8));
  nand2 gate976(.a(gate446inter8), .b(gate446inter7), .O(gate446inter9));
  nand2 gate977(.a(s_61), .b(gate446inter3), .O(gate446inter10));
  nor2  gate978(.a(gate446inter10), .b(gate446inter9), .O(gate446inter11));
  nor2  gate979(.a(gate446inter11), .b(gate446inter6), .O(gate446inter12));
  nand2 gate980(.a(gate446inter12), .b(gate446inter1), .O(G1255));

  xor2  gate1219(.a(G1174), .b(G15), .O(gate447inter0));
  nand2 gate1220(.a(gate447inter0), .b(s_96), .O(gate447inter1));
  and2  gate1221(.a(G1174), .b(G15), .O(gate447inter2));
  inv1  gate1222(.a(s_96), .O(gate447inter3));
  inv1  gate1223(.a(s_97), .O(gate447inter4));
  nand2 gate1224(.a(gate447inter4), .b(gate447inter3), .O(gate447inter5));
  nor2  gate1225(.a(gate447inter5), .b(gate447inter2), .O(gate447inter6));
  inv1  gate1226(.a(G15), .O(gate447inter7));
  inv1  gate1227(.a(G1174), .O(gate447inter8));
  nand2 gate1228(.a(gate447inter8), .b(gate447inter7), .O(gate447inter9));
  nand2 gate1229(.a(s_97), .b(gate447inter3), .O(gate447inter10));
  nor2  gate1230(.a(gate447inter10), .b(gate447inter9), .O(gate447inter11));
  nor2  gate1231(.a(gate447inter11), .b(gate447inter6), .O(gate447inter12));
  nand2 gate1232(.a(gate447inter12), .b(gate447inter1), .O(G1256));
nand2 gate448( .a(G1078), .b(G1174), .O(G1257) );

  xor2  gate1499(.a(G1177), .b(G16), .O(gate449inter0));
  nand2 gate1500(.a(gate449inter0), .b(s_136), .O(gate449inter1));
  and2  gate1501(.a(G1177), .b(G16), .O(gate449inter2));
  inv1  gate1502(.a(s_136), .O(gate449inter3));
  inv1  gate1503(.a(s_137), .O(gate449inter4));
  nand2 gate1504(.a(gate449inter4), .b(gate449inter3), .O(gate449inter5));
  nor2  gate1505(.a(gate449inter5), .b(gate449inter2), .O(gate449inter6));
  inv1  gate1506(.a(G16), .O(gate449inter7));
  inv1  gate1507(.a(G1177), .O(gate449inter8));
  nand2 gate1508(.a(gate449inter8), .b(gate449inter7), .O(gate449inter9));
  nand2 gate1509(.a(s_137), .b(gate449inter3), .O(gate449inter10));
  nor2  gate1510(.a(gate449inter10), .b(gate449inter9), .O(gate449inter11));
  nor2  gate1511(.a(gate449inter11), .b(gate449inter6), .O(gate449inter12));
  nand2 gate1512(.a(gate449inter12), .b(gate449inter1), .O(G1258));
nand2 gate450( .a(G1081), .b(G1177), .O(G1259) );
nand2 gate451( .a(G17), .b(G1180), .O(G1260) );

  xor2  gate1051(.a(G1180), .b(G1084), .O(gate452inter0));
  nand2 gate1052(.a(gate452inter0), .b(s_72), .O(gate452inter1));
  and2  gate1053(.a(G1180), .b(G1084), .O(gate452inter2));
  inv1  gate1054(.a(s_72), .O(gate452inter3));
  inv1  gate1055(.a(s_73), .O(gate452inter4));
  nand2 gate1056(.a(gate452inter4), .b(gate452inter3), .O(gate452inter5));
  nor2  gate1057(.a(gate452inter5), .b(gate452inter2), .O(gate452inter6));
  inv1  gate1058(.a(G1084), .O(gate452inter7));
  inv1  gate1059(.a(G1180), .O(gate452inter8));
  nand2 gate1060(.a(gate452inter8), .b(gate452inter7), .O(gate452inter9));
  nand2 gate1061(.a(s_73), .b(gate452inter3), .O(gate452inter10));
  nor2  gate1062(.a(gate452inter10), .b(gate452inter9), .O(gate452inter11));
  nor2  gate1063(.a(gate452inter11), .b(gate452inter6), .O(gate452inter12));
  nand2 gate1064(.a(gate452inter12), .b(gate452inter1), .O(G1261));

  xor2  gate1289(.a(G1183), .b(G18), .O(gate453inter0));
  nand2 gate1290(.a(gate453inter0), .b(s_106), .O(gate453inter1));
  and2  gate1291(.a(G1183), .b(G18), .O(gate453inter2));
  inv1  gate1292(.a(s_106), .O(gate453inter3));
  inv1  gate1293(.a(s_107), .O(gate453inter4));
  nand2 gate1294(.a(gate453inter4), .b(gate453inter3), .O(gate453inter5));
  nor2  gate1295(.a(gate453inter5), .b(gate453inter2), .O(gate453inter6));
  inv1  gate1296(.a(G18), .O(gate453inter7));
  inv1  gate1297(.a(G1183), .O(gate453inter8));
  nand2 gate1298(.a(gate453inter8), .b(gate453inter7), .O(gate453inter9));
  nand2 gate1299(.a(s_107), .b(gate453inter3), .O(gate453inter10));
  nor2  gate1300(.a(gate453inter10), .b(gate453inter9), .O(gate453inter11));
  nor2  gate1301(.a(gate453inter11), .b(gate453inter6), .O(gate453inter12));
  nand2 gate1302(.a(gate453inter12), .b(gate453inter1), .O(G1262));
nand2 gate454( .a(G1087), .b(G1183), .O(G1263) );
nand2 gate455( .a(G19), .b(G1186), .O(G1264) );
nand2 gate456( .a(G1090), .b(G1186), .O(G1265) );
nand2 gate457( .a(G20), .b(G1189), .O(G1266) );

  xor2  gate883(.a(G1189), .b(G1093), .O(gate458inter0));
  nand2 gate884(.a(gate458inter0), .b(s_48), .O(gate458inter1));
  and2  gate885(.a(G1189), .b(G1093), .O(gate458inter2));
  inv1  gate886(.a(s_48), .O(gate458inter3));
  inv1  gate887(.a(s_49), .O(gate458inter4));
  nand2 gate888(.a(gate458inter4), .b(gate458inter3), .O(gate458inter5));
  nor2  gate889(.a(gate458inter5), .b(gate458inter2), .O(gate458inter6));
  inv1  gate890(.a(G1093), .O(gate458inter7));
  inv1  gate891(.a(G1189), .O(gate458inter8));
  nand2 gate892(.a(gate458inter8), .b(gate458inter7), .O(gate458inter9));
  nand2 gate893(.a(s_49), .b(gate458inter3), .O(gate458inter10));
  nor2  gate894(.a(gate458inter10), .b(gate458inter9), .O(gate458inter11));
  nor2  gate895(.a(gate458inter11), .b(gate458inter6), .O(gate458inter12));
  nand2 gate896(.a(gate458inter12), .b(gate458inter1), .O(G1267));
nand2 gate459( .a(G21), .b(G1192), .O(G1268) );
nand2 gate460( .a(G1096), .b(G1192), .O(G1269) );
nand2 gate461( .a(G22), .b(G1195), .O(G1270) );
nand2 gate462( .a(G1099), .b(G1195), .O(G1271) );

  xor2  gate659(.a(G1198), .b(G23), .O(gate463inter0));
  nand2 gate660(.a(gate463inter0), .b(s_16), .O(gate463inter1));
  and2  gate661(.a(G1198), .b(G23), .O(gate463inter2));
  inv1  gate662(.a(s_16), .O(gate463inter3));
  inv1  gate663(.a(s_17), .O(gate463inter4));
  nand2 gate664(.a(gate463inter4), .b(gate463inter3), .O(gate463inter5));
  nor2  gate665(.a(gate463inter5), .b(gate463inter2), .O(gate463inter6));
  inv1  gate666(.a(G23), .O(gate463inter7));
  inv1  gate667(.a(G1198), .O(gate463inter8));
  nand2 gate668(.a(gate463inter8), .b(gate463inter7), .O(gate463inter9));
  nand2 gate669(.a(s_17), .b(gate463inter3), .O(gate463inter10));
  nor2  gate670(.a(gate463inter10), .b(gate463inter9), .O(gate463inter11));
  nor2  gate671(.a(gate463inter11), .b(gate463inter6), .O(gate463inter12));
  nand2 gate672(.a(gate463inter12), .b(gate463inter1), .O(G1272));
nand2 gate464( .a(G1102), .b(G1198), .O(G1273) );
nand2 gate465( .a(G24), .b(G1201), .O(G1274) );

  xor2  gate1793(.a(G1201), .b(G1105), .O(gate466inter0));
  nand2 gate1794(.a(gate466inter0), .b(s_178), .O(gate466inter1));
  and2  gate1795(.a(G1201), .b(G1105), .O(gate466inter2));
  inv1  gate1796(.a(s_178), .O(gate466inter3));
  inv1  gate1797(.a(s_179), .O(gate466inter4));
  nand2 gate1798(.a(gate466inter4), .b(gate466inter3), .O(gate466inter5));
  nor2  gate1799(.a(gate466inter5), .b(gate466inter2), .O(gate466inter6));
  inv1  gate1800(.a(G1105), .O(gate466inter7));
  inv1  gate1801(.a(G1201), .O(gate466inter8));
  nand2 gate1802(.a(gate466inter8), .b(gate466inter7), .O(gate466inter9));
  nand2 gate1803(.a(s_179), .b(gate466inter3), .O(gate466inter10));
  nor2  gate1804(.a(gate466inter10), .b(gate466inter9), .O(gate466inter11));
  nor2  gate1805(.a(gate466inter11), .b(gate466inter6), .O(gate466inter12));
  nand2 gate1806(.a(gate466inter12), .b(gate466inter1), .O(G1275));
nand2 gate467( .a(G25), .b(G1204), .O(G1276) );

  xor2  gate1765(.a(G1204), .b(G1108), .O(gate468inter0));
  nand2 gate1766(.a(gate468inter0), .b(s_174), .O(gate468inter1));
  and2  gate1767(.a(G1204), .b(G1108), .O(gate468inter2));
  inv1  gate1768(.a(s_174), .O(gate468inter3));
  inv1  gate1769(.a(s_175), .O(gate468inter4));
  nand2 gate1770(.a(gate468inter4), .b(gate468inter3), .O(gate468inter5));
  nor2  gate1771(.a(gate468inter5), .b(gate468inter2), .O(gate468inter6));
  inv1  gate1772(.a(G1108), .O(gate468inter7));
  inv1  gate1773(.a(G1204), .O(gate468inter8));
  nand2 gate1774(.a(gate468inter8), .b(gate468inter7), .O(gate468inter9));
  nand2 gate1775(.a(s_175), .b(gate468inter3), .O(gate468inter10));
  nor2  gate1776(.a(gate468inter10), .b(gate468inter9), .O(gate468inter11));
  nor2  gate1777(.a(gate468inter11), .b(gate468inter6), .O(gate468inter12));
  nand2 gate1778(.a(gate468inter12), .b(gate468inter1), .O(G1277));
nand2 gate469( .a(G26), .b(G1207), .O(G1278) );
nand2 gate470( .a(G1111), .b(G1207), .O(G1279) );
nand2 gate471( .a(G27), .b(G1210), .O(G1280) );
nand2 gate472( .a(G1114), .b(G1210), .O(G1281) );
nand2 gate473( .a(G28), .b(G1213), .O(G1282) );

  xor2  gate1457(.a(G1213), .b(G1117), .O(gate474inter0));
  nand2 gate1458(.a(gate474inter0), .b(s_130), .O(gate474inter1));
  and2  gate1459(.a(G1213), .b(G1117), .O(gate474inter2));
  inv1  gate1460(.a(s_130), .O(gate474inter3));
  inv1  gate1461(.a(s_131), .O(gate474inter4));
  nand2 gate1462(.a(gate474inter4), .b(gate474inter3), .O(gate474inter5));
  nor2  gate1463(.a(gate474inter5), .b(gate474inter2), .O(gate474inter6));
  inv1  gate1464(.a(G1117), .O(gate474inter7));
  inv1  gate1465(.a(G1213), .O(gate474inter8));
  nand2 gate1466(.a(gate474inter8), .b(gate474inter7), .O(gate474inter9));
  nand2 gate1467(.a(s_131), .b(gate474inter3), .O(gate474inter10));
  nor2  gate1468(.a(gate474inter10), .b(gate474inter9), .O(gate474inter11));
  nor2  gate1469(.a(gate474inter11), .b(gate474inter6), .O(gate474inter12));
  nand2 gate1470(.a(gate474inter12), .b(gate474inter1), .O(G1283));
nand2 gate475( .a(G29), .b(G1216), .O(G1284) );
nand2 gate476( .a(G1120), .b(G1216), .O(G1285) );
nand2 gate477( .a(G30), .b(G1219), .O(G1286) );
nand2 gate478( .a(G1123), .b(G1219), .O(G1287) );
nand2 gate479( .a(G31), .b(G1222), .O(G1288) );
nand2 gate480( .a(G1126), .b(G1222), .O(G1289) );

  xor2  gate1135(.a(G1225), .b(G32), .O(gate481inter0));
  nand2 gate1136(.a(gate481inter0), .b(s_84), .O(gate481inter1));
  and2  gate1137(.a(G1225), .b(G32), .O(gate481inter2));
  inv1  gate1138(.a(s_84), .O(gate481inter3));
  inv1  gate1139(.a(s_85), .O(gate481inter4));
  nand2 gate1140(.a(gate481inter4), .b(gate481inter3), .O(gate481inter5));
  nor2  gate1141(.a(gate481inter5), .b(gate481inter2), .O(gate481inter6));
  inv1  gate1142(.a(G32), .O(gate481inter7));
  inv1  gate1143(.a(G1225), .O(gate481inter8));
  nand2 gate1144(.a(gate481inter8), .b(gate481inter7), .O(gate481inter9));
  nand2 gate1145(.a(s_85), .b(gate481inter3), .O(gate481inter10));
  nor2  gate1146(.a(gate481inter10), .b(gate481inter9), .O(gate481inter11));
  nor2  gate1147(.a(gate481inter11), .b(gate481inter6), .O(gate481inter12));
  nand2 gate1148(.a(gate481inter12), .b(gate481inter1), .O(G1290));

  xor2  gate603(.a(G1225), .b(G1129), .O(gate482inter0));
  nand2 gate604(.a(gate482inter0), .b(s_8), .O(gate482inter1));
  and2  gate605(.a(G1225), .b(G1129), .O(gate482inter2));
  inv1  gate606(.a(s_8), .O(gate482inter3));
  inv1  gate607(.a(s_9), .O(gate482inter4));
  nand2 gate608(.a(gate482inter4), .b(gate482inter3), .O(gate482inter5));
  nor2  gate609(.a(gate482inter5), .b(gate482inter2), .O(gate482inter6));
  inv1  gate610(.a(G1129), .O(gate482inter7));
  inv1  gate611(.a(G1225), .O(gate482inter8));
  nand2 gate612(.a(gate482inter8), .b(gate482inter7), .O(gate482inter9));
  nand2 gate613(.a(s_9), .b(gate482inter3), .O(gate482inter10));
  nor2  gate614(.a(gate482inter10), .b(gate482inter9), .O(gate482inter11));
  nor2  gate615(.a(gate482inter11), .b(gate482inter6), .O(gate482inter12));
  nand2 gate616(.a(gate482inter12), .b(gate482inter1), .O(G1291));

  xor2  gate939(.a(G1229), .b(G1228), .O(gate483inter0));
  nand2 gate940(.a(gate483inter0), .b(s_56), .O(gate483inter1));
  and2  gate941(.a(G1229), .b(G1228), .O(gate483inter2));
  inv1  gate942(.a(s_56), .O(gate483inter3));
  inv1  gate943(.a(s_57), .O(gate483inter4));
  nand2 gate944(.a(gate483inter4), .b(gate483inter3), .O(gate483inter5));
  nor2  gate945(.a(gate483inter5), .b(gate483inter2), .O(gate483inter6));
  inv1  gate946(.a(G1228), .O(gate483inter7));
  inv1  gate947(.a(G1229), .O(gate483inter8));
  nand2 gate948(.a(gate483inter8), .b(gate483inter7), .O(gate483inter9));
  nand2 gate949(.a(s_57), .b(gate483inter3), .O(gate483inter10));
  nor2  gate950(.a(gate483inter10), .b(gate483inter9), .O(gate483inter11));
  nor2  gate951(.a(gate483inter11), .b(gate483inter6), .O(gate483inter12));
  nand2 gate952(.a(gate483inter12), .b(gate483inter1), .O(G1292));
nand2 gate484( .a(G1230), .b(G1231), .O(G1293) );
nand2 gate485( .a(G1232), .b(G1233), .O(G1294) );
nand2 gate486( .a(G1234), .b(G1235), .O(G1295) );
nand2 gate487( .a(G1236), .b(G1237), .O(G1296) );
nand2 gate488( .a(G1238), .b(G1239), .O(G1297) );
nand2 gate489( .a(G1240), .b(G1241), .O(G1298) );
nand2 gate490( .a(G1242), .b(G1243), .O(G1299) );
nand2 gate491( .a(G1244), .b(G1245), .O(G1300) );
nand2 gate492( .a(G1246), .b(G1247), .O(G1301) );
nand2 gate493( .a(G1248), .b(G1249), .O(G1302) );

  xor2  gate687(.a(G1251), .b(G1250), .O(gate494inter0));
  nand2 gate688(.a(gate494inter0), .b(s_20), .O(gate494inter1));
  and2  gate689(.a(G1251), .b(G1250), .O(gate494inter2));
  inv1  gate690(.a(s_20), .O(gate494inter3));
  inv1  gate691(.a(s_21), .O(gate494inter4));
  nand2 gate692(.a(gate494inter4), .b(gate494inter3), .O(gate494inter5));
  nor2  gate693(.a(gate494inter5), .b(gate494inter2), .O(gate494inter6));
  inv1  gate694(.a(G1250), .O(gate494inter7));
  inv1  gate695(.a(G1251), .O(gate494inter8));
  nand2 gate696(.a(gate494inter8), .b(gate494inter7), .O(gate494inter9));
  nand2 gate697(.a(s_21), .b(gate494inter3), .O(gate494inter10));
  nor2  gate698(.a(gate494inter10), .b(gate494inter9), .O(gate494inter11));
  nor2  gate699(.a(gate494inter11), .b(gate494inter6), .O(gate494inter12));
  nand2 gate700(.a(gate494inter12), .b(gate494inter1), .O(G1303));
nand2 gate495( .a(G1252), .b(G1253), .O(G1304) );
nand2 gate496( .a(G1254), .b(G1255), .O(G1305) );
nand2 gate497( .a(G1256), .b(G1257), .O(G1306) );
nand2 gate498( .a(G1258), .b(G1259), .O(G1307) );
nand2 gate499( .a(G1260), .b(G1261), .O(G1308) );
nand2 gate500( .a(G1262), .b(G1263), .O(G1309) );

  xor2  gate1583(.a(G1265), .b(G1264), .O(gate501inter0));
  nand2 gate1584(.a(gate501inter0), .b(s_148), .O(gate501inter1));
  and2  gate1585(.a(G1265), .b(G1264), .O(gate501inter2));
  inv1  gate1586(.a(s_148), .O(gate501inter3));
  inv1  gate1587(.a(s_149), .O(gate501inter4));
  nand2 gate1588(.a(gate501inter4), .b(gate501inter3), .O(gate501inter5));
  nor2  gate1589(.a(gate501inter5), .b(gate501inter2), .O(gate501inter6));
  inv1  gate1590(.a(G1264), .O(gate501inter7));
  inv1  gate1591(.a(G1265), .O(gate501inter8));
  nand2 gate1592(.a(gate501inter8), .b(gate501inter7), .O(gate501inter9));
  nand2 gate1593(.a(s_149), .b(gate501inter3), .O(gate501inter10));
  nor2  gate1594(.a(gate501inter10), .b(gate501inter9), .O(gate501inter11));
  nor2  gate1595(.a(gate501inter11), .b(gate501inter6), .O(gate501inter12));
  nand2 gate1596(.a(gate501inter12), .b(gate501inter1), .O(G1310));

  xor2  gate1261(.a(G1267), .b(G1266), .O(gate502inter0));
  nand2 gate1262(.a(gate502inter0), .b(s_102), .O(gate502inter1));
  and2  gate1263(.a(G1267), .b(G1266), .O(gate502inter2));
  inv1  gate1264(.a(s_102), .O(gate502inter3));
  inv1  gate1265(.a(s_103), .O(gate502inter4));
  nand2 gate1266(.a(gate502inter4), .b(gate502inter3), .O(gate502inter5));
  nor2  gate1267(.a(gate502inter5), .b(gate502inter2), .O(gate502inter6));
  inv1  gate1268(.a(G1266), .O(gate502inter7));
  inv1  gate1269(.a(G1267), .O(gate502inter8));
  nand2 gate1270(.a(gate502inter8), .b(gate502inter7), .O(gate502inter9));
  nand2 gate1271(.a(s_103), .b(gate502inter3), .O(gate502inter10));
  nor2  gate1272(.a(gate502inter10), .b(gate502inter9), .O(gate502inter11));
  nor2  gate1273(.a(gate502inter11), .b(gate502inter6), .O(gate502inter12));
  nand2 gate1274(.a(gate502inter12), .b(gate502inter1), .O(G1311));
nand2 gate503( .a(G1268), .b(G1269), .O(G1312) );
nand2 gate504( .a(G1270), .b(G1271), .O(G1313) );
nand2 gate505( .a(G1272), .b(G1273), .O(G1314) );

  xor2  gate1625(.a(G1275), .b(G1274), .O(gate506inter0));
  nand2 gate1626(.a(gate506inter0), .b(s_154), .O(gate506inter1));
  and2  gate1627(.a(G1275), .b(G1274), .O(gate506inter2));
  inv1  gate1628(.a(s_154), .O(gate506inter3));
  inv1  gate1629(.a(s_155), .O(gate506inter4));
  nand2 gate1630(.a(gate506inter4), .b(gate506inter3), .O(gate506inter5));
  nor2  gate1631(.a(gate506inter5), .b(gate506inter2), .O(gate506inter6));
  inv1  gate1632(.a(G1274), .O(gate506inter7));
  inv1  gate1633(.a(G1275), .O(gate506inter8));
  nand2 gate1634(.a(gate506inter8), .b(gate506inter7), .O(gate506inter9));
  nand2 gate1635(.a(s_155), .b(gate506inter3), .O(gate506inter10));
  nor2  gate1636(.a(gate506inter10), .b(gate506inter9), .O(gate506inter11));
  nor2  gate1637(.a(gate506inter11), .b(gate506inter6), .O(gate506inter12));
  nand2 gate1638(.a(gate506inter12), .b(gate506inter1), .O(G1315));

  xor2  gate855(.a(G1277), .b(G1276), .O(gate507inter0));
  nand2 gate856(.a(gate507inter0), .b(s_44), .O(gate507inter1));
  and2  gate857(.a(G1277), .b(G1276), .O(gate507inter2));
  inv1  gate858(.a(s_44), .O(gate507inter3));
  inv1  gate859(.a(s_45), .O(gate507inter4));
  nand2 gate860(.a(gate507inter4), .b(gate507inter3), .O(gate507inter5));
  nor2  gate861(.a(gate507inter5), .b(gate507inter2), .O(gate507inter6));
  inv1  gate862(.a(G1276), .O(gate507inter7));
  inv1  gate863(.a(G1277), .O(gate507inter8));
  nand2 gate864(.a(gate507inter8), .b(gate507inter7), .O(gate507inter9));
  nand2 gate865(.a(s_45), .b(gate507inter3), .O(gate507inter10));
  nor2  gate866(.a(gate507inter10), .b(gate507inter9), .O(gate507inter11));
  nor2  gate867(.a(gate507inter11), .b(gate507inter6), .O(gate507inter12));
  nand2 gate868(.a(gate507inter12), .b(gate507inter1), .O(G1316));

  xor2  gate771(.a(G1279), .b(G1278), .O(gate508inter0));
  nand2 gate772(.a(gate508inter0), .b(s_32), .O(gate508inter1));
  and2  gate773(.a(G1279), .b(G1278), .O(gate508inter2));
  inv1  gate774(.a(s_32), .O(gate508inter3));
  inv1  gate775(.a(s_33), .O(gate508inter4));
  nand2 gate776(.a(gate508inter4), .b(gate508inter3), .O(gate508inter5));
  nor2  gate777(.a(gate508inter5), .b(gate508inter2), .O(gate508inter6));
  inv1  gate778(.a(G1278), .O(gate508inter7));
  inv1  gate779(.a(G1279), .O(gate508inter8));
  nand2 gate780(.a(gate508inter8), .b(gate508inter7), .O(gate508inter9));
  nand2 gate781(.a(s_33), .b(gate508inter3), .O(gate508inter10));
  nor2  gate782(.a(gate508inter10), .b(gate508inter9), .O(gate508inter11));
  nor2  gate783(.a(gate508inter11), .b(gate508inter6), .O(gate508inter12));
  nand2 gate784(.a(gate508inter12), .b(gate508inter1), .O(G1317));
nand2 gate509( .a(G1280), .b(G1281), .O(G1318) );
nand2 gate510( .a(G1282), .b(G1283), .O(G1319) );
nand2 gate511( .a(G1284), .b(G1285), .O(G1320) );
nand2 gate512( .a(G1286), .b(G1287), .O(G1321) );
nand2 gate513( .a(G1288), .b(G1289), .O(G1322) );
nand2 gate514( .a(G1290), .b(G1291), .O(G1323) );
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule