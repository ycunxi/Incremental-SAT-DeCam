module c1908 (N1,N4,N7,N10,N13,N16,N19,N22,N25,N28,
              N31,N34,N37,N40,N43,N46,N49,N53,N56,N60,
              N63,N66,N69,N72,N76,N79,N82,N85,N88,N91,
              N94,N99,N104,N2753,N2754,N2755,N2756,N2762,N2767,N2768,
              N2779,N2780,N2781,N2782,N2783,N2784,N2785,N2786,N2787,N2811,
              N2886,N2887,N2888,N2889,N2890,N2891,N2892,N2899);
input N1,N4,N7,N10,N13,N16,N19,N22,N25,N28,
      N31,N34,N37,N40,N43,N46,N49,N53,N56,N60,
      N63,N66,N69,N72,N76,N79,N82,N85,N88,N91,
      N94,N99,N104;
  input s_0, s_1, s_2, s_3, s_4, s_5, s_6, s_7, s_8, s_9, s_10, s_11, s_12, s_13, s_14, s_15, s_16, s_17, s_18, s_19, s_20, s_21, s_22, s_23, s_24, s_25, s_26, s_27, s_28, s_29, s_30, s_31, s_32, s_33, s_34, s_35, s_36, s_37, s_38, s_39, s_40, s_41, s_42, s_43, s_44, s_45, s_46, s_47, s_48, s_49, s_50, s_51, s_52, s_53, s_54, s_55, s_56, s_57, s_58, s_59, s_60, s_61, s_62, s_63, s_64, s_65, s_66, s_67, s_68, s_69, s_70, s_71, s_72, s_73, s_74, s_75, s_76, s_77, s_78, s_79, s_80, s_81, s_82, s_83, s_84, s_85, s_86, s_87, s_88, s_89, s_90, s_91, s_92, s_93, s_94, s_95, s_96, s_97, s_98, s_99, s_100, s_101, s_102, s_103, s_104, s_105, s_106, s_107, s_108, s_109, s_110, s_111, s_112, s_113, s_114, s_115, s_116, s_117, s_118, s_119, s_120, s_121, s_122, s_123, s_124, s_125, s_126, s_127, s_128, s_129, s_130, s_131;
output N2753,N2754,N2755,N2756,N2762,N2767,N2768,N2779,N2780,N2781,
       N2782,N2783,N2784,N2785,N2786,N2787,N2811,N2886,N2887,N2888,
       N2889,N2890,N2891,N2892,N2899;
wire N190,N194,N197,N201,N206,N209,N212,N216,N220,N225,
     N229,N232,N235,N239,N243,N247,N251,N252,N253,N256,
     N257,N260,N263,N266,N269,N272,N275,N276,N277,N280,
     N283,N290,N297,N300,N303,N306,N313,N316,N319,N326,
     N331,N338,N343,N346,N349,N352,N355,N358,N361,N364,
     N367,N370,N373,N376,N379,N382,N385,N388,N534,N535,
     N536,N537,N538,N539,N540,N541,N542,N543,N544,N545,
     N546,N547,N548,N549,N550,N551,N552,N553,N554,N555,
     N556,N559,N562,N565,N568,N571,N574,N577,N580,N583,
     N586,N589,N592,N595,N598,N601,N602,N603,N608,N612,
     N616,N619,N622,N625,N628,N631,N634,N637,N640,N643,
     N646,N649,N652,N655,N658,N661,N664,N667,N670,N673,
     N676,N679,N682,N685,N688,N691,N694,N697,N700,N703,
     N706,N709,N712,N715,N718,N721,N724,N727,N730,N733,
     N736,N739,N742,N745,N748,N751,N886,N887,N888,N889,
     N890,N891,N892,N893,N894,N895,N896,N897,N898,N899,
     N903,N907,N910,N913,N914,N915,N916,N917,N918,N919,
     N920,N921,N922,N923,N926,N935,N938,N939,N942,N943,
     N946,N947,N950,N951,N954,N955,N958,N959,N962,N965,
     N968,N969,N972,N973,N976,N977,N980,N981,N984,N985,
     N988,N989,N990,N991,N992,N993,N994,N997,N998,N1001,
     N1002,N1003,N1004,N1005,N1006,N1007,N1008,N1009,N1010,N1013,
     N1016,N1019,N1022,N1025,N1028,N1031,N1034,N1037,N1040,N1043,
     N1046,N1049,N1054,N1055,N1063,N1064,N1067,N1068,N1119,N1120,
     N1121,N1122,N1128,N1129,N1130,N1131,N1132,N1133,N1148,N1149,
     N1150,N1151,N1152,N1153,N1154,N1155,N1156,N1157,N1158,N1159,
     N1160,N1161,N1162,N1163,N1164,N1167,N1168,N1171,N1188,N1205,
     N1206,N1207,N1208,N1209,N1210,N1211,N1212,N1213,N1214,N1215,
     N1216,N1217,N1218,N1219,N1220,N1221,N1222,N1223,N1224,N1225,
     N1226,N1227,N1228,N1229,N1230,N1231,N1232,N1235,N1238,N1239,
     N1240,N1241,N1242,N1243,N1246,N1249,N1252,N1255,N1258,N1261,
     N1264,N1267,N1309,N1310,N1311,N1312,N1313,N1314,N1315,N1316,
     N1317,N1318,N1319,N1322,N1327,N1328,N1334,N1344,N1345,N1346,
     N1348,N1349,N1350,N1351,N1352,N1355,N1358,N1361,N1364,N1367,
     N1370,N1373,N1376,N1379,N1383,N1386,N1387,N1388,N1389,N1390,
     N1393,N1396,N1397,N1398,N1399,N1409,N1412,N1413,N1416,N1419,
     N1433,N1434,N1438,N1439,N1440,N1443,N1444,N1445,N1446,N1447,
     N1448,N1451,N1452,N1453,N1454,N1455,N1456,N1457,N1458,N1459,
     N1460,N1461,N1462,N1463,N1464,N1468,N1469,N1470,N1471,N1472,
     N1475,N1476,N1478,N1481,N1484,N1487,N1488,N1489,N1490,N1491,
     N1492,N1493,N1494,N1495,N1496,N1498,N1499,N1500,N1501,N1504,
     N1510,N1513,N1514,N1517,N1520,N1521,N1522,N1526,N1527,N1528,
     N1529,N1530,N1531,N1532,N1534,N1537,N1540,N1546,N1554,N1557,
     N1561,N1567,N1568,N1569,N1571,N1576,N1588,N1591,N1593,N1594,
     N1595,N1596,N1600,N1603,N1606,N1609,N1612,N1615,N1620,N1623,
     N1635,N1636,N1638,N1639,N1640,N1643,N1647,N1651,N1658,N1661,
     N1664,N1671,N1672,N1675,N1677,N1678,N1679,N1680,N1681,N1682,
     N1683,N1685,N1688,N1697,N1701,N1706,N1707,N1708,N1709,N1710,
     N1711,N1712,N1713,N1714,N1717,N1720,N1721,N1723,N1727,N1728,
     N1730,N1731,N1734,N1740,N1741,N1742,N1746,N1747,N1748,N1751,
     N1759,N1761,N1762,N1763,N1764,N1768,N1769,N1772,N1773,N1774,
     N1777,N1783,N1784,N1785,N1786,N1787,N1788,N1791,N1792,N1795,
     N1796,N1798,N1801,N1802,N1807,N1808,N1809,N1810,N1812,N1815,
     N1818,N1821,N1822,N1823,N1824,N1825,N1826,N1827,N1830,N1837,
     N1838,N1841,N1848,N1849,N1850,N1852,N1855,N1856,N1857,N1858,
     N1864,N1865,N1866,N1869,N1872,N1875,N1878,N1879,N1882,N1883,
     N1884,N1885,N1889,N1895,N1896,N1897,N1898,N1902,N1910,N1911,
     N1912,N1913,N1915,N1919,N1920,N1921,N1922,N1923,N1924,N1927,
     N1930,N1933,N1936,N1937,N1938,N1941,N1942,N1944,N1947,N1950,
     N1953,N1958,N1961,N1965,N1968,N1975,N1976,N1977,N1978,N1979,
     N1980,N1985,N1987,N1999,N2000,N2002,N2003,N2004,N2005,N2006,
     N2007,N2008,N2009,N2012,N2013,N2014,N2015,N2016,N2018,N2019,
     N2020,N2021,N2022,N2023,N2024,N2025,N2026,N2027,N2030,N2033,
     N2036,N2037,N2038,N2039,N2040,N2041,N2042,N2047,N2052,N2055,
     N2060,N2061,N2062,N2067,N2068,N2071,N2076,N2077,N2078,N2081,
     N2086,N2089,N2104,N2119,N2129,N2143,N2148,N2151,N2196,N2199,
     N2202,N2205,N2214,N2215,N2216,N2217,N2222,N2223,N2224,N2225,
     N2226,N2227,N2228,N2229,N2230,N2231,N2232,N2233,N2234,N2235,
     N2236,N2237,N2240,N2241,N2244,N2245,N2250,N2253,N2256,N2257,
     N2260,N2263,N2266,N2269,N2272,N2279,N2286,N2297,N2315,N2326,
     N2340,N2353,N2361,N2375,N2384,N2385,N2386,N2426,N2427,N2537,
     N2540,N2543,N2546,N2549,N2552,N2555,N2558,N2561,N2564,N2567,
     N2570,N2573,N2576,N2594,N2597,N2600,N2603,N2606,N2611,N2614,
     N2617,N2620,N2627,N2628,N2629,N2630,N2631,N2632,N2633,N2634,
     N2639,N2642,N2645,N2648,N2651,N2655,N2658,N2661,N2664,N2669,
     N2670,N2671,N2672,N2673,N2674,N2675,N2676,N2682,N2683,N2688,
     N2689,N2690,N2691,N2710,N2720,N2721,N2722,N2723,N2724,N2725,
     N2726,N2727,N2728,N2729,N2730,N2731,N2732,N2733,N2734,N2735,
     N2736,N2737,N2738,N2739,N2740,N2741,N2742,N2743,N2744,N2745,
     N2746,N2747,N2750,N2757,N2758,N2759,N2760,N2761,N2763,N2764,
     N2765,N2766,N2773,N2776,N2788,N2789,N2800,N2807,N2808,N2809,
     N2810,N2812,N2815,N2818,N2821,N2824,N2827,N2828,N2829,N2843,
     N2846,N2850,N2851,N2852,N2853,N2854,N2857,N2858,N2859,N2860,
     N2861,N2862,N2863,N2866,N2867,N2868,N2869,N2870,N2871,N2872,
     N2873,N2874,N2875,N2876,N2877,N2878,N2879,N2880,N2881,N2882,
     N2883,N2895,N2896,N2897,N2898, gate750inter0, gate750inter1, gate750inter2, gate750inter3, gate750inter4, gate750inter5, gate750inter6, gate750inter7, gate750inter8, gate750inter9, gate750inter10, gate750inter11, gate750inter12, gate628inter0, gate628inter1, gate628inter2, gate628inter3, gate628inter4, gate628inter5, gate628inter6, gate628inter7, gate628inter8, gate628inter9, gate628inter10, gate628inter11, gate628inter12, gate414inter0, gate414inter1, gate414inter2, gate414inter3, gate414inter4, gate414inter5, gate414inter6, gate414inter7, gate414inter8, gate414inter9, gate414inter10, gate414inter11, gate414inter12, gate303inter0, gate303inter1, gate303inter2, gate303inter3, gate303inter4, gate303inter5, gate303inter6, gate303inter7, gate303inter8, gate303inter9, gate303inter10, gate303inter11, gate303inter12, gate547inter0, gate547inter1, gate547inter2, gate547inter3, gate547inter4, gate547inter5, gate547inter6, gate547inter7, gate547inter8, gate547inter9, gate547inter10, gate547inter11, gate547inter12, gate17inter0, gate17inter1, gate17inter2, gate17inter3, gate17inter4, gate17inter5, gate17inter6, gate17inter7, gate17inter8, gate17inter9, gate17inter10, gate17inter11, gate17inter12, gate677inter0, gate677inter1, gate677inter2, gate677inter3, gate677inter4, gate677inter5, gate677inter6, gate677inter7, gate677inter8, gate677inter9, gate677inter10, gate677inter11, gate677inter12, gate667inter0, gate667inter1, gate667inter2, gate667inter3, gate667inter4, gate667inter5, gate667inter6, gate667inter7, gate667inter8, gate667inter9, gate667inter10, gate667inter11, gate667inter12, gate259inter0, gate259inter1, gate259inter2, gate259inter3, gate259inter4, gate259inter5, gate259inter6, gate259inter7, gate259inter8, gate259inter9, gate259inter10, gate259inter11, gate259inter12, gate322inter0, gate322inter1, gate322inter2, gate322inter3, gate322inter4, gate322inter5, gate322inter6, gate322inter7, gate322inter8, gate322inter9, gate322inter10, gate322inter11, gate322inter12, gate498inter0, gate498inter1, gate498inter2, gate498inter3, gate498inter4, gate498inter5, gate498inter6, gate498inter7, gate498inter8, gate498inter9, gate498inter10, gate498inter11, gate498inter12, gate559inter0, gate559inter1, gate559inter2, gate559inter3, gate559inter4, gate559inter5, gate559inter6, gate559inter7, gate559inter8, gate559inter9, gate559inter10, gate559inter11, gate559inter12, gate556inter0, gate556inter1, gate556inter2, gate556inter3, gate556inter4, gate556inter5, gate556inter6, gate556inter7, gate556inter8, gate556inter9, gate556inter10, gate556inter11, gate556inter12, gate780inter0, gate780inter1, gate780inter2, gate780inter3, gate780inter4, gate780inter5, gate780inter6, gate780inter7, gate780inter8, gate780inter9, gate780inter10, gate780inter11, gate780inter12, gate237inter0, gate237inter1, gate237inter2, gate237inter3, gate237inter4, gate237inter5, gate237inter6, gate237inter7, gate237inter8, gate237inter9, gate237inter10, gate237inter11, gate237inter12, gate627inter0, gate627inter1, gate627inter2, gate627inter3, gate627inter4, gate627inter5, gate627inter6, gate627inter7, gate627inter8, gate627inter9, gate627inter10, gate627inter11, gate627inter12, gate767inter0, gate767inter1, gate767inter2, gate767inter3, gate767inter4, gate767inter5, gate767inter6, gate767inter7, gate767inter8, gate767inter9, gate767inter10, gate767inter11, gate767inter12, gate563inter0, gate563inter1, gate563inter2, gate563inter3, gate563inter4, gate563inter5, gate563inter6, gate563inter7, gate563inter8, gate563inter9, gate563inter10, gate563inter11, gate563inter12, gate421inter0, gate421inter1, gate421inter2, gate421inter3, gate421inter4, gate421inter5, gate421inter6, gate421inter7, gate421inter8, gate421inter9, gate421inter10, gate421inter11, gate421inter12, gate372inter0, gate372inter1, gate372inter2, gate372inter3, gate372inter4, gate372inter5, gate372inter6, gate372inter7, gate372inter8, gate372inter9, gate372inter10, gate372inter11, gate372inter12, gate404inter0, gate404inter1, gate404inter2, gate404inter3, gate404inter4, gate404inter5, gate404inter6, gate404inter7, gate404inter8, gate404inter9, gate404inter10, gate404inter11, gate404inter12, gate317inter0, gate317inter1, gate317inter2, gate317inter3, gate317inter4, gate317inter5, gate317inter6, gate317inter7, gate317inter8, gate317inter9, gate317inter10, gate317inter11, gate317inter12, gate345inter0, gate345inter1, gate345inter2, gate345inter3, gate345inter4, gate345inter5, gate345inter6, gate345inter7, gate345inter8, gate345inter9, gate345inter10, gate345inter11, gate345inter12, gate343inter0, gate343inter1, gate343inter2, gate343inter3, gate343inter4, gate343inter5, gate343inter6, gate343inter7, gate343inter8, gate343inter9, gate343inter10, gate343inter11, gate343inter12, gate362inter0, gate362inter1, gate362inter2, gate362inter3, gate362inter4, gate362inter5, gate362inter6, gate362inter7, gate362inter8, gate362inter9, gate362inter10, gate362inter11, gate362inter12, gate500inter0, gate500inter1, gate500inter2, gate500inter3, gate500inter4, gate500inter5, gate500inter6, gate500inter7, gate500inter8, gate500inter9, gate500inter10, gate500inter11, gate500inter12, gate298inter0, gate298inter1, gate298inter2, gate298inter3, gate298inter4, gate298inter5, gate298inter6, gate298inter7, gate298inter8, gate298inter9, gate298inter10, gate298inter11, gate298inter12, gate777inter0, gate777inter1, gate777inter2, gate777inter3, gate777inter4, gate777inter5, gate777inter6, gate777inter7, gate777inter8, gate777inter9, gate777inter10, gate777inter11, gate777inter12, gate336inter0, gate336inter1, gate336inter2, gate336inter3, gate336inter4, gate336inter5, gate336inter6, gate336inter7, gate336inter8, gate336inter9, gate336inter10, gate336inter11, gate336inter12, gate410inter0, gate410inter1, gate410inter2, gate410inter3, gate410inter4, gate410inter5, gate410inter6, gate410inter7, gate410inter8, gate410inter9, gate410inter10, gate410inter11, gate410inter12, gate488inter0, gate488inter1, gate488inter2, gate488inter3, gate488inter4, gate488inter5, gate488inter6, gate488inter7, gate488inter8, gate488inter9, gate488inter10, gate488inter11, gate488inter12, gate815inter0, gate815inter1, gate815inter2, gate815inter3, gate815inter4, gate815inter5, gate815inter6, gate815inter7, gate815inter8, gate815inter9, gate815inter10, gate815inter11, gate815inter12, gate601inter0, gate601inter1, gate601inter2, gate601inter3, gate601inter4, gate601inter5, gate601inter6, gate601inter7, gate601inter8, gate601inter9, gate601inter10, gate601inter11, gate601inter12, gate636inter0, gate636inter1, gate636inter2, gate636inter3, gate636inter4, gate636inter5, gate636inter6, gate636inter7, gate636inter8, gate636inter9, gate636inter10, gate636inter11, gate636inter12, gate640inter0, gate640inter1, gate640inter2, gate640inter3, gate640inter4, gate640inter5, gate640inter6, gate640inter7, gate640inter8, gate640inter9, gate640inter10, gate640inter11, gate640inter12, gate453inter0, gate453inter1, gate453inter2, gate453inter3, gate453inter4, gate453inter5, gate453inter6, gate453inter7, gate453inter8, gate453inter9, gate453inter10, gate453inter11, gate453inter12, gate860inter0, gate860inter1, gate860inter2, gate860inter3, gate860inter4, gate860inter5, gate860inter6, gate860inter7, gate860inter8, gate860inter9, gate860inter10, gate860inter11, gate860inter12, gate476inter0, gate476inter1, gate476inter2, gate476inter3, gate476inter4, gate476inter5, gate476inter6, gate476inter7, gate476inter8, gate476inter9, gate476inter10, gate476inter11, gate476inter12, gate161inter0, gate161inter1, gate161inter2, gate161inter3, gate161inter4, gate161inter5, gate161inter6, gate161inter7, gate161inter8, gate161inter9, gate161inter10, gate161inter11, gate161inter12, gate321inter0, gate321inter1, gate321inter2, gate321inter3, gate321inter4, gate321inter5, gate321inter6, gate321inter7, gate321inter8, gate321inter9, gate321inter10, gate321inter11, gate321inter12, gate558inter0, gate558inter1, gate558inter2, gate558inter3, gate558inter4, gate558inter5, gate558inter6, gate558inter7, gate558inter8, gate558inter9, gate558inter10, gate558inter11, gate558inter12, gate370inter0, gate370inter1, gate370inter2, gate370inter3, gate370inter4, gate370inter5, gate370inter6, gate370inter7, gate370inter8, gate370inter9, gate370inter10, gate370inter11, gate370inter12, gate513inter0, gate513inter1, gate513inter2, gate513inter3, gate513inter4, gate513inter5, gate513inter6, gate513inter7, gate513inter8, gate513inter9, gate513inter10, gate513inter11, gate513inter12, gate598inter0, gate598inter1, gate598inter2, gate598inter3, gate598inter4, gate598inter5, gate598inter6, gate598inter7, gate598inter8, gate598inter9, gate598inter10, gate598inter11, gate598inter12, gate574inter0, gate574inter1, gate574inter2, gate574inter3, gate574inter4, gate574inter5, gate574inter6, gate574inter7, gate574inter8, gate574inter9, gate574inter10, gate574inter11, gate574inter12, gate244inter0, gate244inter1, gate244inter2, gate244inter3, gate244inter4, gate244inter5, gate244inter6, gate244inter7, gate244inter8, gate244inter9, gate244inter10, gate244inter11, gate244inter12, gate363inter0, gate363inter1, gate363inter2, gate363inter3, gate363inter4, gate363inter5, gate363inter6, gate363inter7, gate363inter8, gate363inter9, gate363inter10, gate363inter11, gate363inter12, gate432inter0, gate432inter1, gate432inter2, gate432inter3, gate432inter4, gate432inter5, gate432inter6, gate432inter7, gate432inter8, gate432inter9, gate432inter10, gate432inter11, gate432inter12, gate600inter0, gate600inter1, gate600inter2, gate600inter3, gate600inter4, gate600inter5, gate600inter6, gate600inter7, gate600inter8, gate600inter9, gate600inter10, gate600inter11, gate600inter12, gate378inter0, gate378inter1, gate378inter2, gate378inter3, gate378inter4, gate378inter5, gate378inter6, gate378inter7, gate378inter8, gate378inter9, gate378inter10, gate378inter11, gate378inter12, gate626inter0, gate626inter1, gate626inter2, gate626inter3, gate626inter4, gate626inter5, gate626inter6, gate626inter7, gate626inter8, gate626inter9, gate626inter10, gate626inter11, gate626inter12, gate529inter0, gate529inter1, gate529inter2, gate529inter3, gate529inter4, gate529inter5, gate529inter6, gate529inter7, gate529inter8, gate529inter9, gate529inter10, gate529inter11, gate529inter12, gate775inter0, gate775inter1, gate775inter2, gate775inter3, gate775inter4, gate775inter5, gate775inter6, gate775inter7, gate775inter8, gate775inter9, gate775inter10, gate775inter11, gate775inter12, gate828inter0, gate828inter1, gate828inter2, gate828inter3, gate828inter4, gate828inter5, gate828inter6, gate828inter7, gate828inter8, gate828inter9, gate828inter10, gate828inter11, gate828inter12, gate682inter0, gate682inter1, gate682inter2, gate682inter3, gate682inter4, gate682inter5, gate682inter6, gate682inter7, gate682inter8, gate682inter9, gate682inter10, gate682inter11, gate682inter12, gate875inter0, gate875inter1, gate875inter2, gate875inter3, gate875inter4, gate875inter5, gate875inter6, gate875inter7, gate875inter8, gate875inter9, gate875inter10, gate875inter11, gate875inter12, gate684inter0, gate684inter1, gate684inter2, gate684inter3, gate684inter4, gate684inter5, gate684inter6, gate684inter7, gate684inter8, gate684inter9, gate684inter10, gate684inter11, gate684inter12, gate305inter0, gate305inter1, gate305inter2, gate305inter3, gate305inter4, gate305inter5, gate305inter6, gate305inter7, gate305inter8, gate305inter9, gate305inter10, gate305inter11, gate305inter12, gate561inter0, gate561inter1, gate561inter2, gate561inter3, gate561inter4, gate561inter5, gate561inter6, gate561inter7, gate561inter8, gate561inter9, gate561inter10, gate561inter11, gate561inter12, gate854inter0, gate854inter1, gate854inter2, gate854inter3, gate854inter4, gate854inter5, gate854inter6, gate854inter7, gate854inter8, gate854inter9, gate854inter10, gate854inter11, gate854inter12, gate516inter0, gate516inter1, gate516inter2, gate516inter3, gate516inter4, gate516inter5, gate516inter6, gate516inter7, gate516inter8, gate516inter9, gate516inter10, gate516inter11, gate516inter12, gate294inter0, gate294inter1, gate294inter2, gate294inter3, gate294inter4, gate294inter5, gate294inter6, gate294inter7, gate294inter8, gate294inter9, gate294inter10, gate294inter11, gate294inter12, gate822inter0, gate822inter1, gate822inter2, gate822inter3, gate822inter4, gate822inter5, gate822inter6, gate822inter7, gate822inter8, gate822inter9, gate822inter10, gate822inter11, gate822inter12, gate96inter0, gate96inter1, gate96inter2, gate96inter3, gate96inter4, gate96inter5, gate96inter6, gate96inter7, gate96inter8, gate96inter9, gate96inter10, gate96inter11, gate96inter12, gate236inter0, gate236inter1, gate236inter2, gate236inter3, gate236inter4, gate236inter5, gate236inter6, gate236inter7, gate236inter8, gate236inter9, gate236inter10, gate236inter11, gate236inter12, gate766inter0, gate766inter1, gate766inter2, gate766inter3, gate766inter4, gate766inter5, gate766inter6, gate766inter7, gate766inter8, gate766inter9, gate766inter10, gate766inter11, gate766inter12;


inv1 gate1( .a(N1), .O(N190) );
inv1 gate2( .a(N4), .O(N194) );
inv1 gate3( .a(N7), .O(N197) );
inv1 gate4( .a(N10), .O(N201) );
inv1 gate5( .a(N13), .O(N206) );
inv1 gate6( .a(N16), .O(N209) );
inv1 gate7( .a(N19), .O(N212) );
inv1 gate8( .a(N22), .O(N216) );
inv1 gate9( .a(N25), .O(N220) );
inv1 gate10( .a(N28), .O(N225) );
inv1 gate11( .a(N31), .O(N229) );
inv1 gate12( .a(N34), .O(N232) );
inv1 gate13( .a(N37), .O(N235) );
inv1 gate14( .a(N40), .O(N239) );
inv1 gate15( .a(N43), .O(N243) );
inv1 gate16( .a(N46), .O(N247) );

  xor2  gate951(.a(N88), .b(N63), .O(gate17inter0));
  nand2 gate952(.a(gate17inter0), .b(s_10), .O(gate17inter1));
  and2  gate953(.a(N88), .b(N63), .O(gate17inter2));
  inv1  gate954(.a(s_10), .O(gate17inter3));
  inv1  gate955(.a(s_11), .O(gate17inter4));
  nand2 gate956(.a(gate17inter4), .b(gate17inter3), .O(gate17inter5));
  nor2  gate957(.a(gate17inter5), .b(gate17inter2), .O(gate17inter6));
  inv1  gate958(.a(N63), .O(gate17inter7));
  inv1  gate959(.a(N88), .O(gate17inter8));
  nand2 gate960(.a(gate17inter8), .b(gate17inter7), .O(gate17inter9));
  nand2 gate961(.a(s_11), .b(gate17inter3), .O(gate17inter10));
  nor2  gate962(.a(gate17inter10), .b(gate17inter9), .O(gate17inter11));
  nor2  gate963(.a(gate17inter11), .b(gate17inter6), .O(gate17inter12));
  nand2 gate964(.a(gate17inter12), .b(gate17inter1), .O(N251));
nand2 gate18( .a(N66), .b(N91), .O(N252) );
inv1 gate19( .a(N72), .O(N253) );
inv1 gate20( .a(N72), .O(N256) );
buf1 gate21( .a(N69), .O(N257) );
buf1 gate22( .a(N69), .O(N260) );
inv1 gate23( .a(N76), .O(N263) );
inv1 gate24( .a(N79), .O(N266) );
inv1 gate25( .a(N82), .O(N269) );
inv1 gate26( .a(N85), .O(N272) );
inv1 gate27( .a(N104), .O(N275) );
inv1 gate28( .a(N104), .O(N276) );
inv1 gate29( .a(N88), .O(N277) );
inv1 gate30( .a(N91), .O(N280) );
buf1 gate31( .a(N94), .O(N283) );
inv1 gate32( .a(N94), .O(N290) );
buf1 gate33( .a(N94), .O(N297) );
inv1 gate34( .a(N94), .O(N300) );
buf1 gate35( .a(N99), .O(N303) );
inv1 gate36( .a(N99), .O(N306) );
inv1 gate37( .a(N99), .O(N313) );
buf1 gate38( .a(N104), .O(N316) );
inv1 gate39( .a(N104), .O(N319) );
buf1 gate40( .a(N104), .O(N326) );
buf1 gate41( .a(N104), .O(N331) );
inv1 gate42( .a(N104), .O(N338) );
buf1 gate43( .a(N1), .O(N343) );
buf1 gate44( .a(N4), .O(N346) );
buf1 gate45( .a(N7), .O(N349) );
buf1 gate46( .a(N10), .O(N352) );
buf1 gate47( .a(N13), .O(N355) );
buf1 gate48( .a(N16), .O(N358) );
buf1 gate49( .a(N19), .O(N361) );
buf1 gate50( .a(N22), .O(N364) );
buf1 gate51( .a(N25), .O(N367) );
buf1 gate52( .a(N28), .O(N370) );
buf1 gate53( .a(N31), .O(N373) );
buf1 gate54( .a(N34), .O(N376) );
buf1 gate55( .a(N37), .O(N379) );
buf1 gate56( .a(N40), .O(N382) );
buf1 gate57( .a(N43), .O(N385) );
buf1 gate58( .a(N46), .O(N388) );
inv1 gate59( .a(N343), .O(N534) );
inv1 gate60( .a(N346), .O(N535) );
inv1 gate61( .a(N349), .O(N536) );
inv1 gate62( .a(N352), .O(N537) );
inv1 gate63( .a(N355), .O(N538) );
inv1 gate64( .a(N358), .O(N539) );
inv1 gate65( .a(N361), .O(N540) );
inv1 gate66( .a(N364), .O(N541) );
inv1 gate67( .a(N367), .O(N542) );
inv1 gate68( .a(N370), .O(N543) );
inv1 gate69( .a(N373), .O(N544) );
inv1 gate70( .a(N376), .O(N545) );
inv1 gate71( .a(N379), .O(N546) );
inv1 gate72( .a(N382), .O(N547) );
inv1 gate73( .a(N385), .O(N548) );
inv1 gate74( .a(N388), .O(N549) );
nand2 gate75( .a(N306), .b(N331), .O(N550) );
nand2 gate76( .a(N306), .b(N331), .O(N551) );
nand2 gate77( .a(N306), .b(N331), .O(N552) );
nand2 gate78( .a(N306), .b(N331), .O(N553) );
nand2 gate79( .a(N306), .b(N331), .O(N554) );
nand2 gate80( .a(N306), .b(N331), .O(N555) );
buf1 gate81( .a(N190), .O(N556) );
buf1 gate82( .a(N194), .O(N559) );
buf1 gate83( .a(N206), .O(N562) );
buf1 gate84( .a(N209), .O(N565) );
buf1 gate85( .a(N225), .O(N568) );
buf1 gate86( .a(N243), .O(N571) );
and2 gate87( .a(N63), .b(N319), .O(N574) );
buf1 gate88( .a(N220), .O(N577) );
buf1 gate89( .a(N229), .O(N580) );
buf1 gate90( .a(N232), .O(N583) );
and2 gate91( .a(N66), .b(N319), .O(N586) );
buf1 gate92( .a(N239), .O(N589) );
and3 gate93( .a(N49), .b(N253), .c(N319), .O(N592) );
buf1 gate94( .a(N247), .O(N595) );
buf1 gate95( .a(N239), .O(N598) );

  xor2  gate1763(.a(N277), .b(N326), .O(gate96inter0));
  nand2 gate1764(.a(gate96inter0), .b(s_126), .O(gate96inter1));
  and2  gate1765(.a(N277), .b(N326), .O(gate96inter2));
  inv1  gate1766(.a(s_126), .O(gate96inter3));
  inv1  gate1767(.a(s_127), .O(gate96inter4));
  nand2 gate1768(.a(gate96inter4), .b(gate96inter3), .O(gate96inter5));
  nor2  gate1769(.a(gate96inter5), .b(gate96inter2), .O(gate96inter6));
  inv1  gate1770(.a(N326), .O(gate96inter7));
  inv1  gate1771(.a(N277), .O(gate96inter8));
  nand2 gate1772(.a(gate96inter8), .b(gate96inter7), .O(gate96inter9));
  nand2 gate1773(.a(s_127), .b(gate96inter3), .O(gate96inter10));
  nor2  gate1774(.a(gate96inter10), .b(gate96inter9), .O(gate96inter11));
  nor2  gate1775(.a(gate96inter11), .b(gate96inter6), .O(gate96inter12));
  nand2 gate1776(.a(gate96inter12), .b(gate96inter1), .O(N601));
nand2 gate97( .a(N326), .b(N280), .O(N602) );
nand2 gate98( .a(N260), .b(N72), .O(N603) );
nand2 gate99( .a(N260), .b(N300), .O(N608) );
nand2 gate100( .a(N256), .b(N300), .O(N612) );
buf1 gate101( .a(N201), .O(N616) );
buf1 gate102( .a(N216), .O(N619) );
buf1 gate103( .a(N220), .O(N622) );
buf1 gate104( .a(N239), .O(N625) );
buf1 gate105( .a(N190), .O(N628) );
buf1 gate106( .a(N190), .O(N631) );
buf1 gate107( .a(N194), .O(N634) );
buf1 gate108( .a(N229), .O(N637) );
buf1 gate109( .a(N197), .O(N640) );
and3 gate110( .a(N56), .b(N257), .c(N319), .O(N643) );
buf1 gate111( .a(N232), .O(N646) );
buf1 gate112( .a(N201), .O(N649) );
buf1 gate113( .a(N235), .O(N652) );
and3 gate114( .a(N60), .b(N257), .c(N319), .O(N655) );
buf1 gate115( .a(N263), .O(N658) );
buf1 gate116( .a(N263), .O(N661) );
buf1 gate117( .a(N266), .O(N664) );
buf1 gate118( .a(N266), .O(N667) );
buf1 gate119( .a(N269), .O(N670) );
buf1 gate120( .a(N269), .O(N673) );
buf1 gate121( .a(N272), .O(N676) );
buf1 gate122( .a(N272), .O(N679) );
and2 gate123( .a(N251), .b(N316), .O(N682) );
and2 gate124( .a(N252), .b(N316), .O(N685) );
buf1 gate125( .a(N197), .O(N688) );
buf1 gate126( .a(N197), .O(N691) );
buf1 gate127( .a(N212), .O(N694) );
buf1 gate128( .a(N212), .O(N697) );
buf1 gate129( .a(N247), .O(N700) );
buf1 gate130( .a(N247), .O(N703) );
buf1 gate131( .a(N235), .O(N706) );
buf1 gate132( .a(N235), .O(N709) );
buf1 gate133( .a(N201), .O(N712) );
buf1 gate134( .a(N201), .O(N715) );
buf1 gate135( .a(N206), .O(N718) );
buf1 gate136( .a(N216), .O(N721) );
and3 gate137( .a(N53), .b(N253), .c(N319), .O(N724) );
buf1 gate138( .a(N243), .O(N727) );
buf1 gate139( .a(N220), .O(N730) );
buf1 gate140( .a(N220), .O(N733) );
buf1 gate141( .a(N209), .O(N736) );
buf1 gate142( .a(N216), .O(N739) );
buf1 gate143( .a(N225), .O(N742) );
buf1 gate144( .a(N243), .O(N745) );
buf1 gate145( .a(N212), .O(N748) );
buf1 gate146( .a(N225), .O(N751) );
inv1 gate147( .a(N682), .O(N886) );
inv1 gate148( .a(N685), .O(N887) );
inv1 gate149( .a(N616), .O(N888) );
inv1 gate150( .a(N619), .O(N889) );
inv1 gate151( .a(N622), .O(N890) );
inv1 gate152( .a(N625), .O(N891) );
inv1 gate153( .a(N631), .O(N892) );
inv1 gate154( .a(N643), .O(N893) );
inv1 gate155( .a(N649), .O(N894) );
inv1 gate156( .a(N652), .O(N895) );
inv1 gate157( .a(N655), .O(N896) );
and2 gate158( .a(N49), .b(N612), .O(N897) );
and2 gate159( .a(N56), .b(N608), .O(N898) );
nand2 gate160( .a(N53), .b(N612), .O(N899) );

  xor2  gate1413(.a(N608), .b(N60), .O(gate161inter0));
  nand2 gate1414(.a(gate161inter0), .b(s_76), .O(gate161inter1));
  and2  gate1415(.a(N608), .b(N60), .O(gate161inter2));
  inv1  gate1416(.a(s_76), .O(gate161inter3));
  inv1  gate1417(.a(s_77), .O(gate161inter4));
  nand2 gate1418(.a(gate161inter4), .b(gate161inter3), .O(gate161inter5));
  nor2  gate1419(.a(gate161inter5), .b(gate161inter2), .O(gate161inter6));
  inv1  gate1420(.a(N60), .O(gate161inter7));
  inv1  gate1421(.a(N608), .O(gate161inter8));
  nand2 gate1422(.a(gate161inter8), .b(gate161inter7), .O(gate161inter9));
  nand2 gate1423(.a(s_77), .b(gate161inter3), .O(gate161inter10));
  nor2  gate1424(.a(gate161inter10), .b(gate161inter9), .O(gate161inter11));
  nor2  gate1425(.a(gate161inter11), .b(gate161inter6), .O(gate161inter12));
  nand2 gate1426(.a(gate161inter12), .b(gate161inter1), .O(N903));
nand2 gate162( .a(N49), .b(N612), .O(N907) );
nand2 gate163( .a(N56), .b(N608), .O(N910) );
inv1 gate164( .a(N661), .O(N913) );
inv1 gate165( .a(N658), .O(N914) );
inv1 gate166( .a(N667), .O(N915) );
inv1 gate167( .a(N664), .O(N916) );
inv1 gate168( .a(N673), .O(N917) );
inv1 gate169( .a(N670), .O(N918) );
inv1 gate170( .a(N679), .O(N919) );
inv1 gate171( .a(N676), .O(N920) );
nand4 gate172( .a(N277), .b(N297), .c(N326), .d(N603), .O(N921) );
nand4 gate173( .a(N280), .b(N297), .c(N326), .d(N603), .O(N922) );
nand3 gate174( .a(N303), .b(N338), .c(N603), .O(N923) );
and3 gate175( .a(N303), .b(N338), .c(N603), .O(N926) );
buf1 gate176( .a(N556), .O(N935) );
inv1 gate177( .a(N688), .O(N938) );
buf1 gate178( .a(N556), .O(N939) );
inv1 gate179( .a(N691), .O(N942) );
buf1 gate180( .a(N562), .O(N943) );
inv1 gate181( .a(N694), .O(N946) );
buf1 gate182( .a(N562), .O(N947) );
inv1 gate183( .a(N697), .O(N950) );
buf1 gate184( .a(N568), .O(N951) );
inv1 gate185( .a(N700), .O(N954) );
buf1 gate186( .a(N568), .O(N955) );
inv1 gate187( .a(N703), .O(N958) );
buf1 gate188( .a(N574), .O(N959) );
buf1 gate189( .a(N574), .O(N962) );
buf1 gate190( .a(N580), .O(N965) );
inv1 gate191( .a(N706), .O(N968) );
buf1 gate192( .a(N580), .O(N969) );
inv1 gate193( .a(N709), .O(N972) );
buf1 gate194( .a(N586), .O(N973) );
inv1 gate195( .a(N712), .O(N976) );
buf1 gate196( .a(N586), .O(N977) );
inv1 gate197( .a(N715), .O(N980) );
buf1 gate198( .a(N592), .O(N981) );
inv1 gate199( .a(N628), .O(N984) );
buf1 gate200( .a(N592), .O(N985) );
inv1 gate201( .a(N718), .O(N988) );
inv1 gate202( .a(N721), .O(N989) );
inv1 gate203( .a(N634), .O(N990) );
inv1 gate204( .a(N724), .O(N991) );
inv1 gate205( .a(N727), .O(N992) );
inv1 gate206( .a(N637), .O(N993) );
buf1 gate207( .a(N595), .O(N994) );
inv1 gate208( .a(N730), .O(N997) );
buf1 gate209( .a(N595), .O(N998) );
inv1 gate210( .a(N733), .O(N1001) );
inv1 gate211( .a(N736), .O(N1002) );
inv1 gate212( .a(N739), .O(N1003) );
inv1 gate213( .a(N640), .O(N1004) );
inv1 gate214( .a(N742), .O(N1005) );
inv1 gate215( .a(N745), .O(N1006) );
inv1 gate216( .a(N646), .O(N1007) );
inv1 gate217( .a(N748), .O(N1008) );
inv1 gate218( .a(N751), .O(N1009) );
buf1 gate219( .a(N559), .O(N1010) );
buf1 gate220( .a(N559), .O(N1013) );
buf1 gate221( .a(N565), .O(N1016) );
buf1 gate222( .a(N565), .O(N1019) );
buf1 gate223( .a(N571), .O(N1022) );
buf1 gate224( .a(N571), .O(N1025) );
buf1 gate225( .a(N577), .O(N1028) );
buf1 gate226( .a(N577), .O(N1031) );
buf1 gate227( .a(N583), .O(N1034) );
buf1 gate228( .a(N583), .O(N1037) );
buf1 gate229( .a(N589), .O(N1040) );
buf1 gate230( .a(N589), .O(N1043) );
buf1 gate231( .a(N598), .O(N1046) );
buf1 gate232( .a(N598), .O(N1049) );
nand2 gate233( .a(N619), .b(N888), .O(N1054) );
nand2 gate234( .a(N616), .b(N889), .O(N1055) );
nand2 gate235( .a(N625), .b(N890), .O(N1063) );

  xor2  gate1777(.a(N891), .b(N622), .O(gate236inter0));
  nand2 gate1778(.a(gate236inter0), .b(s_128), .O(gate236inter1));
  and2  gate1779(.a(N891), .b(N622), .O(gate236inter2));
  inv1  gate1780(.a(s_128), .O(gate236inter3));
  inv1  gate1781(.a(s_129), .O(gate236inter4));
  nand2 gate1782(.a(gate236inter4), .b(gate236inter3), .O(gate236inter5));
  nor2  gate1783(.a(gate236inter5), .b(gate236inter2), .O(gate236inter6));
  inv1  gate1784(.a(N622), .O(gate236inter7));
  inv1  gate1785(.a(N891), .O(gate236inter8));
  nand2 gate1786(.a(gate236inter8), .b(gate236inter7), .O(gate236inter9));
  nand2 gate1787(.a(s_129), .b(gate236inter3), .O(gate236inter10));
  nor2  gate1788(.a(gate236inter10), .b(gate236inter9), .O(gate236inter11));
  nor2  gate1789(.a(gate236inter11), .b(gate236inter6), .O(gate236inter12));
  nand2 gate1790(.a(gate236inter12), .b(gate236inter1), .O(N1064));

  xor2  gate1077(.a(N895), .b(N655), .O(gate237inter0));
  nand2 gate1078(.a(gate237inter0), .b(s_28), .O(gate237inter1));
  and2  gate1079(.a(N895), .b(N655), .O(gate237inter2));
  inv1  gate1080(.a(s_28), .O(gate237inter3));
  inv1  gate1081(.a(s_29), .O(gate237inter4));
  nand2 gate1082(.a(gate237inter4), .b(gate237inter3), .O(gate237inter5));
  nor2  gate1083(.a(gate237inter5), .b(gate237inter2), .O(gate237inter6));
  inv1  gate1084(.a(N655), .O(gate237inter7));
  inv1  gate1085(.a(N895), .O(gate237inter8));
  nand2 gate1086(.a(gate237inter8), .b(gate237inter7), .O(gate237inter9));
  nand2 gate1087(.a(s_29), .b(gate237inter3), .O(gate237inter10));
  nor2  gate1088(.a(gate237inter10), .b(gate237inter9), .O(gate237inter11));
  nor2  gate1089(.a(gate237inter11), .b(gate237inter6), .O(gate237inter12));
  nand2 gate1090(.a(gate237inter12), .b(gate237inter1), .O(N1067));
nand2 gate238( .a(N652), .b(N896), .O(N1068) );
nand2 gate239( .a(N721), .b(N988), .O(N1119) );
nand2 gate240( .a(N718), .b(N989), .O(N1120) );
nand2 gate241( .a(N727), .b(N991), .O(N1121) );
nand2 gate242( .a(N724), .b(N992), .O(N1122) );
nand2 gate243( .a(N739), .b(N1002), .O(N1128) );

  xor2  gate1511(.a(N1003), .b(N736), .O(gate244inter0));
  nand2 gate1512(.a(gate244inter0), .b(s_90), .O(gate244inter1));
  and2  gate1513(.a(N1003), .b(N736), .O(gate244inter2));
  inv1  gate1514(.a(s_90), .O(gate244inter3));
  inv1  gate1515(.a(s_91), .O(gate244inter4));
  nand2 gate1516(.a(gate244inter4), .b(gate244inter3), .O(gate244inter5));
  nor2  gate1517(.a(gate244inter5), .b(gate244inter2), .O(gate244inter6));
  inv1  gate1518(.a(N736), .O(gate244inter7));
  inv1  gate1519(.a(N1003), .O(gate244inter8));
  nand2 gate1520(.a(gate244inter8), .b(gate244inter7), .O(gate244inter9));
  nand2 gate1521(.a(s_91), .b(gate244inter3), .O(gate244inter10));
  nor2  gate1522(.a(gate244inter10), .b(gate244inter9), .O(gate244inter11));
  nor2  gate1523(.a(gate244inter11), .b(gate244inter6), .O(gate244inter12));
  nand2 gate1524(.a(gate244inter12), .b(gate244inter1), .O(N1129));
nand2 gate245( .a(N745), .b(N1005), .O(N1130) );
nand2 gate246( .a(N742), .b(N1006), .O(N1131) );
nand2 gate247( .a(N751), .b(N1008), .O(N1132) );
nand2 gate248( .a(N748), .b(N1009), .O(N1133) );
inv1 gate249( .a(N939), .O(N1148) );
inv1 gate250( .a(N935), .O(N1149) );
nand2 gate251( .a(N1054), .b(N1055), .O(N1150) );
inv1 gate252( .a(N943), .O(N1151) );
inv1 gate253( .a(N947), .O(N1152) );
inv1 gate254( .a(N955), .O(N1153) );
inv1 gate255( .a(N951), .O(N1154) );
inv1 gate256( .a(N962), .O(N1155) );
inv1 gate257( .a(N969), .O(N1156) );
inv1 gate258( .a(N977), .O(N1157) );

  xor2  gate993(.a(N1064), .b(N1063), .O(gate259inter0));
  nand2 gate994(.a(gate259inter0), .b(s_16), .O(gate259inter1));
  and2  gate995(.a(N1064), .b(N1063), .O(gate259inter2));
  inv1  gate996(.a(s_16), .O(gate259inter3));
  inv1  gate997(.a(s_17), .O(gate259inter4));
  nand2 gate998(.a(gate259inter4), .b(gate259inter3), .O(gate259inter5));
  nor2  gate999(.a(gate259inter5), .b(gate259inter2), .O(gate259inter6));
  inv1  gate1000(.a(N1063), .O(gate259inter7));
  inv1  gate1001(.a(N1064), .O(gate259inter8));
  nand2 gate1002(.a(gate259inter8), .b(gate259inter7), .O(gate259inter9));
  nand2 gate1003(.a(s_17), .b(gate259inter3), .O(gate259inter10));
  nor2  gate1004(.a(gate259inter10), .b(gate259inter9), .O(gate259inter11));
  nor2  gate1005(.a(gate259inter11), .b(gate259inter6), .O(gate259inter12));
  nand2 gate1006(.a(gate259inter12), .b(gate259inter1), .O(N1158));
inv1 gate260( .a(N985), .O(N1159) );
nand2 gate261( .a(N985), .b(N892), .O(N1160) );
inv1 gate262( .a(N998), .O(N1161) );
nand2 gate263( .a(N1067), .b(N1068), .O(N1162) );
inv1 gate264( .a(N899), .O(N1163) );
buf1 gate265( .a(N899), .O(N1164) );
inv1 gate266( .a(N903), .O(N1167) );
buf1 gate267( .a(N903), .O(N1168) );
nand2 gate268( .a(N921), .b(N923), .O(N1171) );
nand2 gate269( .a(N922), .b(N923), .O(N1188) );
inv1 gate270( .a(N1010), .O(N1205) );
nand2 gate271( .a(N1010), .b(N938), .O(N1206) );
inv1 gate272( .a(N1013), .O(N1207) );
nand2 gate273( .a(N1013), .b(N942), .O(N1208) );
inv1 gate274( .a(N1016), .O(N1209) );
nand2 gate275( .a(N1016), .b(N946), .O(N1210) );
inv1 gate276( .a(N1019), .O(N1211) );
nand2 gate277( .a(N1019), .b(N950), .O(N1212) );
inv1 gate278( .a(N1022), .O(N1213) );
nand2 gate279( .a(N1022), .b(N954), .O(N1214) );
inv1 gate280( .a(N1025), .O(N1215) );
nand2 gate281( .a(N1025), .b(N958), .O(N1216) );
inv1 gate282( .a(N1028), .O(N1217) );
inv1 gate283( .a(N959), .O(N1218) );
inv1 gate284( .a(N1031), .O(N1219) );
inv1 gate285( .a(N1034), .O(N1220) );
nand2 gate286( .a(N1034), .b(N968), .O(N1221) );
inv1 gate287( .a(N965), .O(N1222) );
inv1 gate288( .a(N1037), .O(N1223) );
nand2 gate289( .a(N1037), .b(N972), .O(N1224) );
inv1 gate290( .a(N1040), .O(N1225) );
nand2 gate291( .a(N1040), .b(N976), .O(N1226) );
inv1 gate292( .a(N973), .O(N1227) );
inv1 gate293( .a(N1043), .O(N1228) );

  xor2  gate1735(.a(N980), .b(N1043), .O(gate294inter0));
  nand2 gate1736(.a(gate294inter0), .b(s_122), .O(gate294inter1));
  and2  gate1737(.a(N980), .b(N1043), .O(gate294inter2));
  inv1  gate1738(.a(s_122), .O(gate294inter3));
  inv1  gate1739(.a(s_123), .O(gate294inter4));
  nand2 gate1740(.a(gate294inter4), .b(gate294inter3), .O(gate294inter5));
  nor2  gate1741(.a(gate294inter5), .b(gate294inter2), .O(gate294inter6));
  inv1  gate1742(.a(N1043), .O(gate294inter7));
  inv1  gate1743(.a(N980), .O(gate294inter8));
  nand2 gate1744(.a(gate294inter8), .b(gate294inter7), .O(gate294inter9));
  nand2 gate1745(.a(s_123), .b(gate294inter3), .O(gate294inter10));
  nor2  gate1746(.a(gate294inter10), .b(gate294inter9), .O(gate294inter11));
  nor2  gate1747(.a(gate294inter11), .b(gate294inter6), .O(gate294inter12));
  nand2 gate1748(.a(gate294inter12), .b(gate294inter1), .O(N1229));
inv1 gate295( .a(N981), .O(N1230) );
nand2 gate296( .a(N981), .b(N984), .O(N1231) );
nand2 gate297( .a(N1119), .b(N1120), .O(N1232) );

  xor2  gate1245(.a(N1122), .b(N1121), .O(gate298inter0));
  nand2 gate1246(.a(gate298inter0), .b(s_52), .O(gate298inter1));
  and2  gate1247(.a(N1122), .b(N1121), .O(gate298inter2));
  inv1  gate1248(.a(s_52), .O(gate298inter3));
  inv1  gate1249(.a(s_53), .O(gate298inter4));
  nand2 gate1250(.a(gate298inter4), .b(gate298inter3), .O(gate298inter5));
  nor2  gate1251(.a(gate298inter5), .b(gate298inter2), .O(gate298inter6));
  inv1  gate1252(.a(N1121), .O(gate298inter7));
  inv1  gate1253(.a(N1122), .O(gate298inter8));
  nand2 gate1254(.a(gate298inter8), .b(gate298inter7), .O(gate298inter9));
  nand2 gate1255(.a(s_53), .b(gate298inter3), .O(gate298inter10));
  nor2  gate1256(.a(gate298inter10), .b(gate298inter9), .O(gate298inter11));
  nor2  gate1257(.a(gate298inter11), .b(gate298inter6), .O(gate298inter12));
  nand2 gate1258(.a(gate298inter12), .b(gate298inter1), .O(N1235));
inv1 gate299( .a(N1046), .O(N1238) );
nand2 gate300( .a(N1046), .b(N997), .O(N1239) );
inv1 gate301( .a(N994), .O(N1240) );
inv1 gate302( .a(N1049), .O(N1241) );

  xor2  gate923(.a(N1001), .b(N1049), .O(gate303inter0));
  nand2 gate924(.a(gate303inter0), .b(s_6), .O(gate303inter1));
  and2  gate925(.a(N1001), .b(N1049), .O(gate303inter2));
  inv1  gate926(.a(s_6), .O(gate303inter3));
  inv1  gate927(.a(s_7), .O(gate303inter4));
  nand2 gate928(.a(gate303inter4), .b(gate303inter3), .O(gate303inter5));
  nor2  gate929(.a(gate303inter5), .b(gate303inter2), .O(gate303inter6));
  inv1  gate930(.a(N1049), .O(gate303inter7));
  inv1  gate931(.a(N1001), .O(gate303inter8));
  nand2 gate932(.a(gate303inter8), .b(gate303inter7), .O(gate303inter9));
  nand2 gate933(.a(s_7), .b(gate303inter3), .O(gate303inter10));
  nor2  gate934(.a(gate303inter10), .b(gate303inter9), .O(gate303inter11));
  nor2  gate935(.a(gate303inter11), .b(gate303inter6), .O(gate303inter12));
  nand2 gate936(.a(gate303inter12), .b(gate303inter1), .O(N1242));
nand2 gate304( .a(N1128), .b(N1129), .O(N1243) );

  xor2  gate1679(.a(N1131), .b(N1130), .O(gate305inter0));
  nand2 gate1680(.a(gate305inter0), .b(s_114), .O(gate305inter1));
  and2  gate1681(.a(N1131), .b(N1130), .O(gate305inter2));
  inv1  gate1682(.a(s_114), .O(gate305inter3));
  inv1  gate1683(.a(s_115), .O(gate305inter4));
  nand2 gate1684(.a(gate305inter4), .b(gate305inter3), .O(gate305inter5));
  nor2  gate1685(.a(gate305inter5), .b(gate305inter2), .O(gate305inter6));
  inv1  gate1686(.a(N1130), .O(gate305inter7));
  inv1  gate1687(.a(N1131), .O(gate305inter8));
  nand2 gate1688(.a(gate305inter8), .b(gate305inter7), .O(gate305inter9));
  nand2 gate1689(.a(s_115), .b(gate305inter3), .O(gate305inter10));
  nor2  gate1690(.a(gate305inter10), .b(gate305inter9), .O(gate305inter11));
  nor2  gate1691(.a(gate305inter11), .b(gate305inter6), .O(gate305inter12));
  nand2 gate1692(.a(gate305inter12), .b(gate305inter1), .O(N1246));
nand2 gate306( .a(N1132), .b(N1133), .O(N1249) );
buf1 gate307( .a(N907), .O(N1252) );
buf1 gate308( .a(N907), .O(N1255) );
buf1 gate309( .a(N910), .O(N1258) );
buf1 gate310( .a(N910), .O(N1261) );
inv1 gate311( .a(N1150), .O(N1264) );
nand2 gate312( .a(N631), .b(N1159), .O(N1267) );
nand2 gate313( .a(N688), .b(N1205), .O(N1309) );
nand2 gate314( .a(N691), .b(N1207), .O(N1310) );
nand2 gate315( .a(N694), .b(N1209), .O(N1311) );
nand2 gate316( .a(N697), .b(N1211), .O(N1312) );

  xor2  gate1175(.a(N1213), .b(N700), .O(gate317inter0));
  nand2 gate1176(.a(gate317inter0), .b(s_42), .O(gate317inter1));
  and2  gate1177(.a(N1213), .b(N700), .O(gate317inter2));
  inv1  gate1178(.a(s_42), .O(gate317inter3));
  inv1  gate1179(.a(s_43), .O(gate317inter4));
  nand2 gate1180(.a(gate317inter4), .b(gate317inter3), .O(gate317inter5));
  nor2  gate1181(.a(gate317inter5), .b(gate317inter2), .O(gate317inter6));
  inv1  gate1182(.a(N700), .O(gate317inter7));
  inv1  gate1183(.a(N1213), .O(gate317inter8));
  nand2 gate1184(.a(gate317inter8), .b(gate317inter7), .O(gate317inter9));
  nand2 gate1185(.a(s_43), .b(gate317inter3), .O(gate317inter10));
  nor2  gate1186(.a(gate317inter10), .b(gate317inter9), .O(gate317inter11));
  nor2  gate1187(.a(gate317inter11), .b(gate317inter6), .O(gate317inter12));
  nand2 gate1188(.a(gate317inter12), .b(gate317inter1), .O(N1313));
nand2 gate318( .a(N703), .b(N1215), .O(N1314) );
nand2 gate319( .a(N706), .b(N1220), .O(N1315) );
nand2 gate320( .a(N709), .b(N1223), .O(N1316) );

  xor2  gate1427(.a(N1225), .b(N712), .O(gate321inter0));
  nand2 gate1428(.a(gate321inter0), .b(s_78), .O(gate321inter1));
  and2  gate1429(.a(N1225), .b(N712), .O(gate321inter2));
  inv1  gate1430(.a(s_78), .O(gate321inter3));
  inv1  gate1431(.a(s_79), .O(gate321inter4));
  nand2 gate1432(.a(gate321inter4), .b(gate321inter3), .O(gate321inter5));
  nor2  gate1433(.a(gate321inter5), .b(gate321inter2), .O(gate321inter6));
  inv1  gate1434(.a(N712), .O(gate321inter7));
  inv1  gate1435(.a(N1225), .O(gate321inter8));
  nand2 gate1436(.a(gate321inter8), .b(gate321inter7), .O(gate321inter9));
  nand2 gate1437(.a(s_79), .b(gate321inter3), .O(gate321inter10));
  nor2  gate1438(.a(gate321inter10), .b(gate321inter9), .O(gate321inter11));
  nor2  gate1439(.a(gate321inter11), .b(gate321inter6), .O(gate321inter12));
  nand2 gate1440(.a(gate321inter12), .b(gate321inter1), .O(N1317));

  xor2  gate1007(.a(N1228), .b(N715), .O(gate322inter0));
  nand2 gate1008(.a(gate322inter0), .b(s_18), .O(gate322inter1));
  and2  gate1009(.a(N1228), .b(N715), .O(gate322inter2));
  inv1  gate1010(.a(s_18), .O(gate322inter3));
  inv1  gate1011(.a(s_19), .O(gate322inter4));
  nand2 gate1012(.a(gate322inter4), .b(gate322inter3), .O(gate322inter5));
  nor2  gate1013(.a(gate322inter5), .b(gate322inter2), .O(gate322inter6));
  inv1  gate1014(.a(N715), .O(gate322inter7));
  inv1  gate1015(.a(N1228), .O(gate322inter8));
  nand2 gate1016(.a(gate322inter8), .b(gate322inter7), .O(gate322inter9));
  nand2 gate1017(.a(s_19), .b(gate322inter3), .O(gate322inter10));
  nor2  gate1018(.a(gate322inter10), .b(gate322inter9), .O(gate322inter11));
  nor2  gate1019(.a(gate322inter11), .b(gate322inter6), .O(gate322inter12));
  nand2 gate1020(.a(gate322inter12), .b(gate322inter1), .O(N1318));
inv1 gate323( .a(N1158), .O(N1319) );
nand2 gate324( .a(N628), .b(N1230), .O(N1322) );
nand2 gate325( .a(N730), .b(N1238), .O(N1327) );
nand2 gate326( .a(N733), .b(N1241), .O(N1328) );
inv1 gate327( .a(N1162), .O(N1334) );
nand2 gate328( .a(N1267), .b(N1160), .O(N1344) );
nand2 gate329( .a(N1249), .b(N894), .O(N1345) );
inv1 gate330( .a(N1249), .O(N1346) );
inv1 gate331( .a(N1255), .O(N1348) );
inv1 gate332( .a(N1252), .O(N1349) );
inv1 gate333( .a(N1261), .O(N1350) );
inv1 gate334( .a(N1258), .O(N1351) );
nand2 gate335( .a(N1309), .b(N1206), .O(N1352) );

  xor2  gate1273(.a(N1208), .b(N1310), .O(gate336inter0));
  nand2 gate1274(.a(gate336inter0), .b(s_56), .O(gate336inter1));
  and2  gate1275(.a(N1208), .b(N1310), .O(gate336inter2));
  inv1  gate1276(.a(s_56), .O(gate336inter3));
  inv1  gate1277(.a(s_57), .O(gate336inter4));
  nand2 gate1278(.a(gate336inter4), .b(gate336inter3), .O(gate336inter5));
  nor2  gate1279(.a(gate336inter5), .b(gate336inter2), .O(gate336inter6));
  inv1  gate1280(.a(N1310), .O(gate336inter7));
  inv1  gate1281(.a(N1208), .O(gate336inter8));
  nand2 gate1282(.a(gate336inter8), .b(gate336inter7), .O(gate336inter9));
  nand2 gate1283(.a(s_57), .b(gate336inter3), .O(gate336inter10));
  nor2  gate1284(.a(gate336inter10), .b(gate336inter9), .O(gate336inter11));
  nor2  gate1285(.a(gate336inter11), .b(gate336inter6), .O(gate336inter12));
  nand2 gate1286(.a(gate336inter12), .b(gate336inter1), .O(N1355));
nand2 gate337( .a(N1311), .b(N1210), .O(N1358) );
nand2 gate338( .a(N1312), .b(N1212), .O(N1361) );
nand2 gate339( .a(N1313), .b(N1214), .O(N1364) );
nand2 gate340( .a(N1314), .b(N1216), .O(N1367) );
nand2 gate341( .a(N1315), .b(N1221), .O(N1370) );
nand2 gate342( .a(N1316), .b(N1224), .O(N1373) );

  xor2  gate1203(.a(N1226), .b(N1317), .O(gate343inter0));
  nand2 gate1204(.a(gate343inter0), .b(s_46), .O(gate343inter1));
  and2  gate1205(.a(N1226), .b(N1317), .O(gate343inter2));
  inv1  gate1206(.a(s_46), .O(gate343inter3));
  inv1  gate1207(.a(s_47), .O(gate343inter4));
  nand2 gate1208(.a(gate343inter4), .b(gate343inter3), .O(gate343inter5));
  nor2  gate1209(.a(gate343inter5), .b(gate343inter2), .O(gate343inter6));
  inv1  gate1210(.a(N1317), .O(gate343inter7));
  inv1  gate1211(.a(N1226), .O(gate343inter8));
  nand2 gate1212(.a(gate343inter8), .b(gate343inter7), .O(gate343inter9));
  nand2 gate1213(.a(s_47), .b(gate343inter3), .O(gate343inter10));
  nor2  gate1214(.a(gate343inter10), .b(gate343inter9), .O(gate343inter11));
  nor2  gate1215(.a(gate343inter11), .b(gate343inter6), .O(gate343inter12));
  nand2 gate1216(.a(gate343inter12), .b(gate343inter1), .O(N1376));
nand2 gate344( .a(N1318), .b(N1229), .O(N1379) );

  xor2  gate1189(.a(N1231), .b(N1322), .O(gate345inter0));
  nand2 gate1190(.a(gate345inter0), .b(s_44), .O(gate345inter1));
  and2  gate1191(.a(N1231), .b(N1322), .O(gate345inter2));
  inv1  gate1192(.a(s_44), .O(gate345inter3));
  inv1  gate1193(.a(s_45), .O(gate345inter4));
  nand2 gate1194(.a(gate345inter4), .b(gate345inter3), .O(gate345inter5));
  nor2  gate1195(.a(gate345inter5), .b(gate345inter2), .O(gate345inter6));
  inv1  gate1196(.a(N1322), .O(gate345inter7));
  inv1  gate1197(.a(N1231), .O(gate345inter8));
  nand2 gate1198(.a(gate345inter8), .b(gate345inter7), .O(gate345inter9));
  nand2 gate1199(.a(s_45), .b(gate345inter3), .O(gate345inter10));
  nor2  gate1200(.a(gate345inter10), .b(gate345inter9), .O(gate345inter11));
  nor2  gate1201(.a(gate345inter11), .b(gate345inter6), .O(gate345inter12));
  nand2 gate1202(.a(gate345inter12), .b(gate345inter1), .O(N1383));
inv1 gate346( .a(N1232), .O(N1386) );
nand2 gate347( .a(N1232), .b(N990), .O(N1387) );
inv1 gate348( .a(N1235), .O(N1388) );
nand2 gate349( .a(N1235), .b(N993), .O(N1389) );
nand2 gate350( .a(N1327), .b(N1239), .O(N1390) );
nand2 gate351( .a(N1328), .b(N1242), .O(N1393) );
inv1 gate352( .a(N1243), .O(N1396) );
nand2 gate353( .a(N1243), .b(N1004), .O(N1397) );
inv1 gate354( .a(N1246), .O(N1398) );
nand2 gate355( .a(N1246), .b(N1007), .O(N1399) );
inv1 gate356( .a(N1319), .O(N1409) );
nand2 gate357( .a(N649), .b(N1346), .O(N1412) );
inv1 gate358( .a(N1334), .O(N1413) );
buf1 gate359( .a(N1264), .O(N1416) );
buf1 gate360( .a(N1264), .O(N1419) );
nand2 gate361( .a(N634), .b(N1386), .O(N1433) );

  xor2  gate1217(.a(N1388), .b(N637), .O(gate362inter0));
  nand2 gate1218(.a(gate362inter0), .b(s_48), .O(gate362inter1));
  and2  gate1219(.a(N1388), .b(N637), .O(gate362inter2));
  inv1  gate1220(.a(s_48), .O(gate362inter3));
  inv1  gate1221(.a(s_49), .O(gate362inter4));
  nand2 gate1222(.a(gate362inter4), .b(gate362inter3), .O(gate362inter5));
  nor2  gate1223(.a(gate362inter5), .b(gate362inter2), .O(gate362inter6));
  inv1  gate1224(.a(N637), .O(gate362inter7));
  inv1  gate1225(.a(N1388), .O(gate362inter8));
  nand2 gate1226(.a(gate362inter8), .b(gate362inter7), .O(gate362inter9));
  nand2 gate1227(.a(s_49), .b(gate362inter3), .O(gate362inter10));
  nor2  gate1228(.a(gate362inter10), .b(gate362inter9), .O(gate362inter11));
  nor2  gate1229(.a(gate362inter11), .b(gate362inter6), .O(gate362inter12));
  nand2 gate1230(.a(gate362inter12), .b(gate362inter1), .O(N1434));

  xor2  gate1525(.a(N1396), .b(N640), .O(gate363inter0));
  nand2 gate1526(.a(gate363inter0), .b(s_92), .O(gate363inter1));
  and2  gate1527(.a(N1396), .b(N640), .O(gate363inter2));
  inv1  gate1528(.a(s_92), .O(gate363inter3));
  inv1  gate1529(.a(s_93), .O(gate363inter4));
  nand2 gate1530(.a(gate363inter4), .b(gate363inter3), .O(gate363inter5));
  nor2  gate1531(.a(gate363inter5), .b(gate363inter2), .O(gate363inter6));
  inv1  gate1532(.a(N640), .O(gate363inter7));
  inv1  gate1533(.a(N1396), .O(gate363inter8));
  nand2 gate1534(.a(gate363inter8), .b(gate363inter7), .O(gate363inter9));
  nand2 gate1535(.a(s_93), .b(gate363inter3), .O(gate363inter10));
  nor2  gate1536(.a(gate363inter10), .b(gate363inter9), .O(gate363inter11));
  nor2  gate1537(.a(gate363inter11), .b(gate363inter6), .O(gate363inter12));
  nand2 gate1538(.a(gate363inter12), .b(gate363inter1), .O(N1438));
nand2 gate364( .a(N646), .b(N1398), .O(N1439) );
inv1 gate365( .a(N1344), .O(N1440) );
nand2 gate366( .a(N1355), .b(N1148), .O(N1443) );
inv1 gate367( .a(N1355), .O(N1444) );
nand2 gate368( .a(N1352), .b(N1149), .O(N1445) );
inv1 gate369( .a(N1352), .O(N1446) );

  xor2  gate1455(.a(N1151), .b(N1358), .O(gate370inter0));
  nand2 gate1456(.a(gate370inter0), .b(s_82), .O(gate370inter1));
  and2  gate1457(.a(N1151), .b(N1358), .O(gate370inter2));
  inv1  gate1458(.a(s_82), .O(gate370inter3));
  inv1  gate1459(.a(s_83), .O(gate370inter4));
  nand2 gate1460(.a(gate370inter4), .b(gate370inter3), .O(gate370inter5));
  nor2  gate1461(.a(gate370inter5), .b(gate370inter2), .O(gate370inter6));
  inv1  gate1462(.a(N1358), .O(gate370inter7));
  inv1  gate1463(.a(N1151), .O(gate370inter8));
  nand2 gate1464(.a(gate370inter8), .b(gate370inter7), .O(gate370inter9));
  nand2 gate1465(.a(s_83), .b(gate370inter3), .O(gate370inter10));
  nor2  gate1466(.a(gate370inter10), .b(gate370inter9), .O(gate370inter11));
  nor2  gate1467(.a(gate370inter11), .b(gate370inter6), .O(gate370inter12));
  nand2 gate1468(.a(gate370inter12), .b(gate370inter1), .O(N1447));
inv1 gate371( .a(N1358), .O(N1448) );

  xor2  gate1147(.a(N1152), .b(N1361), .O(gate372inter0));
  nand2 gate1148(.a(gate372inter0), .b(s_38), .O(gate372inter1));
  and2  gate1149(.a(N1152), .b(N1361), .O(gate372inter2));
  inv1  gate1150(.a(s_38), .O(gate372inter3));
  inv1  gate1151(.a(s_39), .O(gate372inter4));
  nand2 gate1152(.a(gate372inter4), .b(gate372inter3), .O(gate372inter5));
  nor2  gate1153(.a(gate372inter5), .b(gate372inter2), .O(gate372inter6));
  inv1  gate1154(.a(N1361), .O(gate372inter7));
  inv1  gate1155(.a(N1152), .O(gate372inter8));
  nand2 gate1156(.a(gate372inter8), .b(gate372inter7), .O(gate372inter9));
  nand2 gate1157(.a(s_39), .b(gate372inter3), .O(gate372inter10));
  nor2  gate1158(.a(gate372inter10), .b(gate372inter9), .O(gate372inter11));
  nor2  gate1159(.a(gate372inter11), .b(gate372inter6), .O(gate372inter12));
  nand2 gate1160(.a(gate372inter12), .b(gate372inter1), .O(N1451));
inv1 gate373( .a(N1361), .O(N1452) );
nand2 gate374( .a(N1367), .b(N1153), .O(N1453) );
inv1 gate375( .a(N1367), .O(N1454) );
nand2 gate376( .a(N1364), .b(N1154), .O(N1455) );
inv1 gate377( .a(N1364), .O(N1456) );

  xor2  gate1567(.a(N1156), .b(N1373), .O(gate378inter0));
  nand2 gate1568(.a(gate378inter0), .b(s_98), .O(gate378inter1));
  and2  gate1569(.a(N1156), .b(N1373), .O(gate378inter2));
  inv1  gate1570(.a(s_98), .O(gate378inter3));
  inv1  gate1571(.a(s_99), .O(gate378inter4));
  nand2 gate1572(.a(gate378inter4), .b(gate378inter3), .O(gate378inter5));
  nor2  gate1573(.a(gate378inter5), .b(gate378inter2), .O(gate378inter6));
  inv1  gate1574(.a(N1373), .O(gate378inter7));
  inv1  gate1575(.a(N1156), .O(gate378inter8));
  nand2 gate1576(.a(gate378inter8), .b(gate378inter7), .O(gate378inter9));
  nand2 gate1577(.a(s_99), .b(gate378inter3), .O(gate378inter10));
  nor2  gate1578(.a(gate378inter10), .b(gate378inter9), .O(gate378inter11));
  nor2  gate1579(.a(gate378inter11), .b(gate378inter6), .O(gate378inter12));
  nand2 gate1580(.a(gate378inter12), .b(gate378inter1), .O(N1457));
inv1 gate379( .a(N1373), .O(N1458) );
nand2 gate380( .a(N1379), .b(N1157), .O(N1459) );
inv1 gate381( .a(N1379), .O(N1460) );
inv1 gate382( .a(N1383), .O(N1461) );
nand2 gate383( .a(N1393), .b(N1161), .O(N1462) );
inv1 gate384( .a(N1393), .O(N1463) );
nand2 gate385( .a(N1345), .b(N1412), .O(N1464) );
inv1 gate386( .a(N1370), .O(N1468) );
nand2 gate387( .a(N1370), .b(N1222), .O(N1469) );
inv1 gate388( .a(N1376), .O(N1470) );
nand2 gate389( .a(N1376), .b(N1227), .O(N1471) );
nand2 gate390( .a(N1387), .b(N1433), .O(N1472) );
inv1 gate391( .a(N1390), .O(N1475) );
nand2 gate392( .a(N1390), .b(N1240), .O(N1476) );
nand2 gate393( .a(N1389), .b(N1434), .O(N1478) );
nand2 gate394( .a(N1399), .b(N1439), .O(N1481) );
nand2 gate395( .a(N1397), .b(N1438), .O(N1484) );
nand2 gate396( .a(N939), .b(N1444), .O(N1487) );
nand2 gate397( .a(N935), .b(N1446), .O(N1488) );
nand2 gate398( .a(N943), .b(N1448), .O(N1489) );
inv1 gate399( .a(N1419), .O(N1490) );
inv1 gate400( .a(N1416), .O(N1491) );
nand2 gate401( .a(N947), .b(N1452), .O(N1492) );
nand2 gate402( .a(N955), .b(N1454), .O(N1493) );
nand2 gate403( .a(N951), .b(N1456), .O(N1494) );

  xor2  gate1161(.a(N1458), .b(N969), .O(gate404inter0));
  nand2 gate1162(.a(gate404inter0), .b(s_40), .O(gate404inter1));
  and2  gate1163(.a(N1458), .b(N969), .O(gate404inter2));
  inv1  gate1164(.a(s_40), .O(gate404inter3));
  inv1  gate1165(.a(s_41), .O(gate404inter4));
  nand2 gate1166(.a(gate404inter4), .b(gate404inter3), .O(gate404inter5));
  nor2  gate1167(.a(gate404inter5), .b(gate404inter2), .O(gate404inter6));
  inv1  gate1168(.a(N969), .O(gate404inter7));
  inv1  gate1169(.a(N1458), .O(gate404inter8));
  nand2 gate1170(.a(gate404inter8), .b(gate404inter7), .O(gate404inter9));
  nand2 gate1171(.a(s_41), .b(gate404inter3), .O(gate404inter10));
  nor2  gate1172(.a(gate404inter10), .b(gate404inter9), .O(gate404inter11));
  nor2  gate1173(.a(gate404inter11), .b(gate404inter6), .O(gate404inter12));
  nand2 gate1174(.a(gate404inter12), .b(gate404inter1), .O(N1495));
nand2 gate405( .a(N977), .b(N1460), .O(N1496) );
nand2 gate406( .a(N998), .b(N1463), .O(N1498) );
inv1 gate407( .a(N1440), .O(N1499) );
nand2 gate408( .a(N965), .b(N1468), .O(N1500) );
nand2 gate409( .a(N973), .b(N1470), .O(N1501) );

  xor2  gate1287(.a(N1475), .b(N994), .O(gate410inter0));
  nand2 gate1288(.a(gate410inter0), .b(s_58), .O(gate410inter1));
  and2  gate1289(.a(N1475), .b(N994), .O(gate410inter2));
  inv1  gate1290(.a(s_58), .O(gate410inter3));
  inv1  gate1291(.a(s_59), .O(gate410inter4));
  nand2 gate1292(.a(gate410inter4), .b(gate410inter3), .O(gate410inter5));
  nor2  gate1293(.a(gate410inter5), .b(gate410inter2), .O(gate410inter6));
  inv1  gate1294(.a(N994), .O(gate410inter7));
  inv1  gate1295(.a(N1475), .O(gate410inter8));
  nand2 gate1296(.a(gate410inter8), .b(gate410inter7), .O(gate410inter9));
  nand2 gate1297(.a(s_59), .b(gate410inter3), .O(gate410inter10));
  nor2  gate1298(.a(gate410inter10), .b(gate410inter9), .O(gate410inter11));
  nor2  gate1299(.a(gate410inter11), .b(gate410inter6), .O(gate410inter12));
  nand2 gate1300(.a(gate410inter12), .b(gate410inter1), .O(N1504));
inv1 gate411( .a(N1464), .O(N1510) );
nand2 gate412( .a(N1443), .b(N1487), .O(N1513) );
nand2 gate413( .a(N1445), .b(N1488), .O(N1514) );

  xor2  gate909(.a(N1489), .b(N1447), .O(gate414inter0));
  nand2 gate910(.a(gate414inter0), .b(s_4), .O(gate414inter1));
  and2  gate911(.a(N1489), .b(N1447), .O(gate414inter2));
  inv1  gate912(.a(s_4), .O(gate414inter3));
  inv1  gate913(.a(s_5), .O(gate414inter4));
  nand2 gate914(.a(gate414inter4), .b(gate414inter3), .O(gate414inter5));
  nor2  gate915(.a(gate414inter5), .b(gate414inter2), .O(gate414inter6));
  inv1  gate916(.a(N1447), .O(gate414inter7));
  inv1  gate917(.a(N1489), .O(gate414inter8));
  nand2 gate918(.a(gate414inter8), .b(gate414inter7), .O(gate414inter9));
  nand2 gate919(.a(s_5), .b(gate414inter3), .O(gate414inter10));
  nor2  gate920(.a(gate414inter10), .b(gate414inter9), .O(gate414inter11));
  nor2  gate921(.a(gate414inter11), .b(gate414inter6), .O(gate414inter12));
  nand2 gate922(.a(gate414inter12), .b(gate414inter1), .O(N1517));
nand2 gate415( .a(N1451), .b(N1492), .O(N1520) );
nand2 gate416( .a(N1453), .b(N1493), .O(N1521) );
nand2 gate417( .a(N1455), .b(N1494), .O(N1522) );
nand2 gate418( .a(N1457), .b(N1495), .O(N1526) );
nand2 gate419( .a(N1459), .b(N1496), .O(N1527) );
inv1 gate420( .a(N1472), .O(N1528) );

  xor2  gate1133(.a(N1498), .b(N1462), .O(gate421inter0));
  nand2 gate1134(.a(gate421inter0), .b(s_36), .O(gate421inter1));
  and2  gate1135(.a(N1498), .b(N1462), .O(gate421inter2));
  inv1  gate1136(.a(s_36), .O(gate421inter3));
  inv1  gate1137(.a(s_37), .O(gate421inter4));
  nand2 gate1138(.a(gate421inter4), .b(gate421inter3), .O(gate421inter5));
  nor2  gate1139(.a(gate421inter5), .b(gate421inter2), .O(gate421inter6));
  inv1  gate1140(.a(N1462), .O(gate421inter7));
  inv1  gate1141(.a(N1498), .O(gate421inter8));
  nand2 gate1142(.a(gate421inter8), .b(gate421inter7), .O(gate421inter9));
  nand2 gate1143(.a(s_37), .b(gate421inter3), .O(gate421inter10));
  nor2  gate1144(.a(gate421inter10), .b(gate421inter9), .O(gate421inter11));
  nor2  gate1145(.a(gate421inter11), .b(gate421inter6), .O(gate421inter12));
  nand2 gate1146(.a(gate421inter12), .b(gate421inter1), .O(N1529));
inv1 gate422( .a(N1478), .O(N1530) );
inv1 gate423( .a(N1481), .O(N1531) );
inv1 gate424( .a(N1484), .O(N1532) );
nand2 gate425( .a(N1471), .b(N1501), .O(N1534) );
nand2 gate426( .a(N1469), .b(N1500), .O(N1537) );
nand2 gate427( .a(N1476), .b(N1504), .O(N1540) );
inv1 gate428( .a(N1513), .O(N1546) );
inv1 gate429( .a(N1521), .O(N1554) );
inv1 gate430( .a(N1526), .O(N1557) );
inv1 gate431( .a(N1520), .O(N1561) );

  xor2  gate1539(.a(N1531), .b(N1484), .O(gate432inter0));
  nand2 gate1540(.a(gate432inter0), .b(s_94), .O(gate432inter1));
  and2  gate1541(.a(N1531), .b(N1484), .O(gate432inter2));
  inv1  gate1542(.a(s_94), .O(gate432inter3));
  inv1  gate1543(.a(s_95), .O(gate432inter4));
  nand2 gate1544(.a(gate432inter4), .b(gate432inter3), .O(gate432inter5));
  nor2  gate1545(.a(gate432inter5), .b(gate432inter2), .O(gate432inter6));
  inv1  gate1546(.a(N1484), .O(gate432inter7));
  inv1  gate1547(.a(N1531), .O(gate432inter8));
  nand2 gate1548(.a(gate432inter8), .b(gate432inter7), .O(gate432inter9));
  nand2 gate1549(.a(s_95), .b(gate432inter3), .O(gate432inter10));
  nor2  gate1550(.a(gate432inter10), .b(gate432inter9), .O(gate432inter11));
  nor2  gate1551(.a(gate432inter11), .b(gate432inter6), .O(gate432inter12));
  nand2 gate1552(.a(gate432inter12), .b(gate432inter1), .O(N1567));
nand2 gate433( .a(N1481), .b(N1532), .O(N1568) );
inv1 gate434( .a(N1510), .O(N1569) );
inv1 gate435( .a(N1527), .O(N1571) );
inv1 gate436( .a(N1529), .O(N1576) );
buf1 gate437( .a(N1522), .O(N1588) );
inv1 gate438( .a(N1534), .O(N1591) );
inv1 gate439( .a(N1537), .O(N1593) );
nand2 gate440( .a(N1540), .b(N1530), .O(N1594) );
inv1 gate441( .a(N1540), .O(N1595) );
nand2 gate442( .a(N1567), .b(N1568), .O(N1596) );
buf1 gate443( .a(N1517), .O(N1600) );
buf1 gate444( .a(N1517), .O(N1603) );
buf1 gate445( .a(N1522), .O(N1606) );
buf1 gate446( .a(N1522), .O(N1609) );
buf1 gate447( .a(N1514), .O(N1612) );
buf1 gate448( .a(N1514), .O(N1615) );
buf1 gate449( .a(N1557), .O(N1620) );
buf1 gate450( .a(N1554), .O(N1623) );
inv1 gate451( .a(N1571), .O(N1635) );
nand2 gate452( .a(N1478), .b(N1595), .O(N1636) );

  xor2  gate1371(.a(N1569), .b(N1576), .O(gate453inter0));
  nand2 gate1372(.a(gate453inter0), .b(s_70), .O(gate453inter1));
  and2  gate1373(.a(N1569), .b(N1576), .O(gate453inter2));
  inv1  gate1374(.a(s_70), .O(gate453inter3));
  inv1  gate1375(.a(s_71), .O(gate453inter4));
  nand2 gate1376(.a(gate453inter4), .b(gate453inter3), .O(gate453inter5));
  nor2  gate1377(.a(gate453inter5), .b(gate453inter2), .O(gate453inter6));
  inv1  gate1378(.a(N1576), .O(gate453inter7));
  inv1  gate1379(.a(N1569), .O(gate453inter8));
  nand2 gate1380(.a(gate453inter8), .b(gate453inter7), .O(gate453inter9));
  nand2 gate1381(.a(s_71), .b(gate453inter3), .O(gate453inter10));
  nor2  gate1382(.a(gate453inter10), .b(gate453inter9), .O(gate453inter11));
  nor2  gate1383(.a(gate453inter11), .b(gate453inter6), .O(gate453inter12));
  nand2 gate1384(.a(gate453inter12), .b(gate453inter1), .O(N1638));
inv1 gate454( .a(N1576), .O(N1639) );
buf1 gate455( .a(N1561), .O(N1640) );
buf1 gate456( .a(N1561), .O(N1643) );
buf1 gate457( .a(N1546), .O(N1647) );
buf1 gate458( .a(N1546), .O(N1651) );
buf1 gate459( .a(N1554), .O(N1658) );
buf1 gate460( .a(N1557), .O(N1661) );
buf1 gate461( .a(N1557), .O(N1664) );
nand2 gate462( .a(N1596), .b(N893), .O(N1671) );
inv1 gate463( .a(N1596), .O(N1672) );
inv1 gate464( .a(N1600), .O(N1675) );
inv1 gate465( .a(N1603), .O(N1677) );
nand2 gate466( .a(N1606), .b(N1217), .O(N1678) );
inv1 gate467( .a(N1606), .O(N1679) );
nand2 gate468( .a(N1609), .b(N1219), .O(N1680) );
inv1 gate469( .a(N1609), .O(N1681) );
inv1 gate470( .a(N1612), .O(N1682) );
inv1 gate471( .a(N1615), .O(N1683) );
nand2 gate472( .a(N1594), .b(N1636), .O(N1685) );
nand2 gate473( .a(N1510), .b(N1639), .O(N1688) );
buf1 gate474( .a(N1588), .O(N1697) );
buf1 gate475( .a(N1588), .O(N1701) );

  xor2  gate1399(.a(N1672), .b(N643), .O(gate476inter0));
  nand2 gate1400(.a(gate476inter0), .b(s_74), .O(gate476inter1));
  and2  gate1401(.a(N1672), .b(N643), .O(gate476inter2));
  inv1  gate1402(.a(s_74), .O(gate476inter3));
  inv1  gate1403(.a(s_75), .O(gate476inter4));
  nand2 gate1404(.a(gate476inter4), .b(gate476inter3), .O(gate476inter5));
  nor2  gate1405(.a(gate476inter5), .b(gate476inter2), .O(gate476inter6));
  inv1  gate1406(.a(N643), .O(gate476inter7));
  inv1  gate1407(.a(N1672), .O(gate476inter8));
  nand2 gate1408(.a(gate476inter8), .b(gate476inter7), .O(gate476inter9));
  nand2 gate1409(.a(s_75), .b(gate476inter3), .O(gate476inter10));
  nor2  gate1410(.a(gate476inter10), .b(gate476inter9), .O(gate476inter11));
  nor2  gate1411(.a(gate476inter11), .b(gate476inter6), .O(gate476inter12));
  nand2 gate1412(.a(gate476inter12), .b(gate476inter1), .O(N1706));
inv1 gate477( .a(N1643), .O(N1707) );
nand2 gate478( .a(N1647), .b(N1675), .O(N1708) );
inv1 gate479( .a(N1647), .O(N1709) );
nand2 gate480( .a(N1651), .b(N1677), .O(N1710) );
inv1 gate481( .a(N1651), .O(N1711) );
nand2 gate482( .a(N1028), .b(N1679), .O(N1712) );
nand2 gate483( .a(N1031), .b(N1681), .O(N1713) );
buf1 gate484( .a(N1620), .O(N1714) );
buf1 gate485( .a(N1620), .O(N1717) );
nand2 gate486( .a(N1658), .b(N1593), .O(N1720) );
inv1 gate487( .a(N1658), .O(N1721) );

  xor2  gate1301(.a(N1688), .b(N1638), .O(gate488inter0));
  nand2 gate1302(.a(gate488inter0), .b(s_60), .O(gate488inter1));
  and2  gate1303(.a(N1688), .b(N1638), .O(gate488inter2));
  inv1  gate1304(.a(s_60), .O(gate488inter3));
  inv1  gate1305(.a(s_61), .O(gate488inter4));
  nand2 gate1306(.a(gate488inter4), .b(gate488inter3), .O(gate488inter5));
  nor2  gate1307(.a(gate488inter5), .b(gate488inter2), .O(gate488inter6));
  inv1  gate1308(.a(N1638), .O(gate488inter7));
  inv1  gate1309(.a(N1688), .O(gate488inter8));
  nand2 gate1310(.a(gate488inter8), .b(gate488inter7), .O(gate488inter9));
  nand2 gate1311(.a(s_61), .b(gate488inter3), .O(gate488inter10));
  nor2  gate1312(.a(gate488inter10), .b(gate488inter9), .O(gate488inter11));
  nor2  gate1313(.a(gate488inter11), .b(gate488inter6), .O(gate488inter12));
  nand2 gate1314(.a(gate488inter12), .b(gate488inter1), .O(N1723));
inv1 gate489( .a(N1661), .O(N1727) );
inv1 gate490( .a(N1640), .O(N1728) );
inv1 gate491( .a(N1664), .O(N1730) );
buf1 gate492( .a(N1623), .O(N1731) );
buf1 gate493( .a(N1623), .O(N1734) );
nand2 gate494( .a(N1685), .b(N1528), .O(N1740) );
inv1 gate495( .a(N1685), .O(N1741) );
nand2 gate496( .a(N1671), .b(N1706), .O(N1742) );
nand2 gate497( .a(N1600), .b(N1709), .O(N1746) );

  xor2  gate1021(.a(N1711), .b(N1603), .O(gate498inter0));
  nand2 gate1022(.a(gate498inter0), .b(s_20), .O(gate498inter1));
  and2  gate1023(.a(N1711), .b(N1603), .O(gate498inter2));
  inv1  gate1024(.a(s_20), .O(gate498inter3));
  inv1  gate1025(.a(s_21), .O(gate498inter4));
  nand2 gate1026(.a(gate498inter4), .b(gate498inter3), .O(gate498inter5));
  nor2  gate1027(.a(gate498inter5), .b(gate498inter2), .O(gate498inter6));
  inv1  gate1028(.a(N1603), .O(gate498inter7));
  inv1  gate1029(.a(N1711), .O(gate498inter8));
  nand2 gate1030(.a(gate498inter8), .b(gate498inter7), .O(gate498inter9));
  nand2 gate1031(.a(s_21), .b(gate498inter3), .O(gate498inter10));
  nor2  gate1032(.a(gate498inter10), .b(gate498inter9), .O(gate498inter11));
  nor2  gate1033(.a(gate498inter11), .b(gate498inter6), .O(gate498inter12));
  nand2 gate1034(.a(gate498inter12), .b(gate498inter1), .O(N1747));
nand2 gate499( .a(N1678), .b(N1712), .O(N1748) );

  xor2  gate1231(.a(N1713), .b(N1680), .O(gate500inter0));
  nand2 gate1232(.a(gate500inter0), .b(s_50), .O(gate500inter1));
  and2  gate1233(.a(N1713), .b(N1680), .O(gate500inter2));
  inv1  gate1234(.a(s_50), .O(gate500inter3));
  inv1  gate1235(.a(s_51), .O(gate500inter4));
  nand2 gate1236(.a(gate500inter4), .b(gate500inter3), .O(gate500inter5));
  nor2  gate1237(.a(gate500inter5), .b(gate500inter2), .O(gate500inter6));
  inv1  gate1238(.a(N1680), .O(gate500inter7));
  inv1  gate1239(.a(N1713), .O(gate500inter8));
  nand2 gate1240(.a(gate500inter8), .b(gate500inter7), .O(gate500inter9));
  nand2 gate1241(.a(s_51), .b(gate500inter3), .O(gate500inter10));
  nor2  gate1242(.a(gate500inter10), .b(gate500inter9), .O(gate500inter11));
  nor2  gate1243(.a(gate500inter11), .b(gate500inter6), .O(gate500inter12));
  nand2 gate1244(.a(gate500inter12), .b(gate500inter1), .O(N1751));
nand2 gate501( .a(N1537), .b(N1721), .O(N1759) );
inv1 gate502( .a(N1697), .O(N1761) );
nand2 gate503( .a(N1697), .b(N1727), .O(N1762) );
inv1 gate504( .a(N1701), .O(N1763) );
nand2 gate505( .a(N1701), .b(N1730), .O(N1764) );
inv1 gate506( .a(N1717), .O(N1768) );
nand2 gate507( .a(N1472), .b(N1741), .O(N1769) );
nand2 gate508( .a(N1723), .b(N1413), .O(N1772) );
inv1 gate509( .a(N1723), .O(N1773) );
nand2 gate510( .a(N1708), .b(N1746), .O(N1774) );
nand2 gate511( .a(N1710), .b(N1747), .O(N1777) );
inv1 gate512( .a(N1731), .O(N1783) );

  xor2  gate1469(.a(N1682), .b(N1731), .O(gate513inter0));
  nand2 gate1470(.a(gate513inter0), .b(s_84), .O(gate513inter1));
  and2  gate1471(.a(N1682), .b(N1731), .O(gate513inter2));
  inv1  gate1472(.a(s_84), .O(gate513inter3));
  inv1  gate1473(.a(s_85), .O(gate513inter4));
  nand2 gate1474(.a(gate513inter4), .b(gate513inter3), .O(gate513inter5));
  nor2  gate1475(.a(gate513inter5), .b(gate513inter2), .O(gate513inter6));
  inv1  gate1476(.a(N1731), .O(gate513inter7));
  inv1  gate1477(.a(N1682), .O(gate513inter8));
  nand2 gate1478(.a(gate513inter8), .b(gate513inter7), .O(gate513inter9));
  nand2 gate1479(.a(s_85), .b(gate513inter3), .O(gate513inter10));
  nor2  gate1480(.a(gate513inter10), .b(gate513inter9), .O(gate513inter11));
  nor2  gate1481(.a(gate513inter11), .b(gate513inter6), .O(gate513inter12));
  nand2 gate1482(.a(gate513inter12), .b(gate513inter1), .O(N1784));
inv1 gate514( .a(N1714), .O(N1785) );
inv1 gate515( .a(N1734), .O(N1786) );

  xor2  gate1721(.a(N1683), .b(N1734), .O(gate516inter0));
  nand2 gate1722(.a(gate516inter0), .b(s_120), .O(gate516inter1));
  and2  gate1723(.a(N1683), .b(N1734), .O(gate516inter2));
  inv1  gate1724(.a(s_120), .O(gate516inter3));
  inv1  gate1725(.a(s_121), .O(gate516inter4));
  nand2 gate1726(.a(gate516inter4), .b(gate516inter3), .O(gate516inter5));
  nor2  gate1727(.a(gate516inter5), .b(gate516inter2), .O(gate516inter6));
  inv1  gate1728(.a(N1734), .O(gate516inter7));
  inv1  gate1729(.a(N1683), .O(gate516inter8));
  nand2 gate1730(.a(gate516inter8), .b(gate516inter7), .O(gate516inter9));
  nand2 gate1731(.a(s_121), .b(gate516inter3), .O(gate516inter10));
  nor2  gate1732(.a(gate516inter10), .b(gate516inter9), .O(gate516inter11));
  nor2  gate1733(.a(gate516inter11), .b(gate516inter6), .O(gate516inter12));
  nand2 gate1734(.a(gate516inter12), .b(gate516inter1), .O(N1787));
nand2 gate517( .a(N1720), .b(N1759), .O(N1788) );
nand2 gate518( .a(N1661), .b(N1761), .O(N1791) );
nand2 gate519( .a(N1664), .b(N1763), .O(N1792) );
nand2 gate520( .a(N1751), .b(N1155), .O(N1795) );
inv1 gate521( .a(N1751), .O(N1796) );
nand2 gate522( .a(N1740), .b(N1769), .O(N1798) );
nand2 gate523( .a(N1334), .b(N1773), .O(N1801) );
nand2 gate524( .a(N1742), .b(N290), .O(N1802) );
inv1 gate525( .a(N1748), .O(N1807) );
nand2 gate526( .a(N1748), .b(N1218), .O(N1808) );
nand2 gate527( .a(N1612), .b(N1783), .O(N1809) );
nand2 gate528( .a(N1615), .b(N1786), .O(N1810) );

  xor2  gate1595(.a(N1762), .b(N1791), .O(gate529inter0));
  nand2 gate1596(.a(gate529inter0), .b(s_102), .O(gate529inter1));
  and2  gate1597(.a(N1762), .b(N1791), .O(gate529inter2));
  inv1  gate1598(.a(s_102), .O(gate529inter3));
  inv1  gate1599(.a(s_103), .O(gate529inter4));
  nand2 gate1600(.a(gate529inter4), .b(gate529inter3), .O(gate529inter5));
  nor2  gate1601(.a(gate529inter5), .b(gate529inter2), .O(gate529inter6));
  inv1  gate1602(.a(N1791), .O(gate529inter7));
  inv1  gate1603(.a(N1762), .O(gate529inter8));
  nand2 gate1604(.a(gate529inter8), .b(gate529inter7), .O(gate529inter9));
  nand2 gate1605(.a(s_103), .b(gate529inter3), .O(gate529inter10));
  nor2  gate1606(.a(gate529inter10), .b(gate529inter9), .O(gate529inter11));
  nor2  gate1607(.a(gate529inter11), .b(gate529inter6), .O(gate529inter12));
  nand2 gate1608(.a(gate529inter12), .b(gate529inter1), .O(N1812));
nand2 gate530( .a(N1792), .b(N1764), .O(N1815) );
buf1 gate531( .a(N1742), .O(N1818) );
nand2 gate532( .a(N1777), .b(N1490), .O(N1821) );
inv1 gate533( .a(N1777), .O(N1822) );
nand2 gate534( .a(N1774), .b(N1491), .O(N1823) );
inv1 gate535( .a(N1774), .O(N1824) );
nand2 gate536( .a(N962), .b(N1796), .O(N1825) );
nand2 gate537( .a(N1788), .b(N1409), .O(N1826) );
inv1 gate538( .a(N1788), .O(N1827) );
nand2 gate539( .a(N1772), .b(N1801), .O(N1830) );
nand2 gate540( .a(N959), .b(N1807), .O(N1837) );
nand2 gate541( .a(N1809), .b(N1784), .O(N1838) );
nand2 gate542( .a(N1810), .b(N1787), .O(N1841) );
nand2 gate543( .a(N1419), .b(N1822), .O(N1848) );
nand2 gate544( .a(N1416), .b(N1824), .O(N1849) );
nand2 gate545( .a(N1795), .b(N1825), .O(N1850) );
nand2 gate546( .a(N1319), .b(N1827), .O(N1852) );

  xor2  gate937(.a(N1707), .b(N1815), .O(gate547inter0));
  nand2 gate938(.a(gate547inter0), .b(s_8), .O(gate547inter1));
  and2  gate939(.a(N1707), .b(N1815), .O(gate547inter2));
  inv1  gate940(.a(s_8), .O(gate547inter3));
  inv1  gate941(.a(s_9), .O(gate547inter4));
  nand2 gate942(.a(gate547inter4), .b(gate547inter3), .O(gate547inter5));
  nor2  gate943(.a(gate547inter5), .b(gate547inter2), .O(gate547inter6));
  inv1  gate944(.a(N1815), .O(gate547inter7));
  inv1  gate945(.a(N1707), .O(gate547inter8));
  nand2 gate946(.a(gate547inter8), .b(gate547inter7), .O(gate547inter9));
  nand2 gate947(.a(s_9), .b(gate547inter3), .O(gate547inter10));
  nor2  gate948(.a(gate547inter10), .b(gate547inter9), .O(gate547inter11));
  nor2  gate949(.a(gate547inter11), .b(gate547inter6), .O(gate547inter12));
  nand2 gate950(.a(gate547inter12), .b(gate547inter1), .O(N1855));
inv1 gate548( .a(N1815), .O(N1856) );
inv1 gate549( .a(N1818), .O(N1857) );
nand2 gate550( .a(N1798), .b(N290), .O(N1858) );
inv1 gate551( .a(N1812), .O(N1864) );
nand2 gate552( .a(N1812), .b(N1728), .O(N1865) );
buf1 gate553( .a(N1798), .O(N1866) );
buf1 gate554( .a(N1802), .O(N1869) );
buf1 gate555( .a(N1802), .O(N1872) );

  xor2  gate1049(.a(N1837), .b(N1808), .O(gate556inter0));
  nand2 gate1050(.a(gate556inter0), .b(s_24), .O(gate556inter1));
  and2  gate1051(.a(N1837), .b(N1808), .O(gate556inter2));
  inv1  gate1052(.a(s_24), .O(gate556inter3));
  inv1  gate1053(.a(s_25), .O(gate556inter4));
  nand2 gate1054(.a(gate556inter4), .b(gate556inter3), .O(gate556inter5));
  nor2  gate1055(.a(gate556inter5), .b(gate556inter2), .O(gate556inter6));
  inv1  gate1056(.a(N1808), .O(gate556inter7));
  inv1  gate1057(.a(N1837), .O(gate556inter8));
  nand2 gate1058(.a(gate556inter8), .b(gate556inter7), .O(gate556inter9));
  nand2 gate1059(.a(s_25), .b(gate556inter3), .O(gate556inter10));
  nor2  gate1060(.a(gate556inter10), .b(gate556inter9), .O(gate556inter11));
  nor2  gate1061(.a(gate556inter11), .b(gate556inter6), .O(gate556inter12));
  nand2 gate1062(.a(gate556inter12), .b(gate556inter1), .O(N1875));
nand2 gate557( .a(N1821), .b(N1848), .O(N1878) );

  xor2  gate1441(.a(N1849), .b(N1823), .O(gate558inter0));
  nand2 gate1442(.a(gate558inter0), .b(s_80), .O(gate558inter1));
  and2  gate1443(.a(N1849), .b(N1823), .O(gate558inter2));
  inv1  gate1444(.a(s_80), .O(gate558inter3));
  inv1  gate1445(.a(s_81), .O(gate558inter4));
  nand2 gate1446(.a(gate558inter4), .b(gate558inter3), .O(gate558inter5));
  nor2  gate1447(.a(gate558inter5), .b(gate558inter2), .O(gate558inter6));
  inv1  gate1448(.a(N1823), .O(gate558inter7));
  inv1  gate1449(.a(N1849), .O(gate558inter8));
  nand2 gate1450(.a(gate558inter8), .b(gate558inter7), .O(gate558inter9));
  nand2 gate1451(.a(s_81), .b(gate558inter3), .O(gate558inter10));
  nor2  gate1452(.a(gate558inter10), .b(gate558inter9), .O(gate558inter11));
  nor2  gate1453(.a(gate558inter11), .b(gate558inter6), .O(gate558inter12));
  nand2 gate1454(.a(gate558inter12), .b(gate558inter1), .O(N1879));

  xor2  gate1035(.a(N1768), .b(N1841), .O(gate559inter0));
  nand2 gate1036(.a(gate559inter0), .b(s_22), .O(gate559inter1));
  and2  gate1037(.a(N1768), .b(N1841), .O(gate559inter2));
  inv1  gate1038(.a(s_22), .O(gate559inter3));
  inv1  gate1039(.a(s_23), .O(gate559inter4));
  nand2 gate1040(.a(gate559inter4), .b(gate559inter3), .O(gate559inter5));
  nor2  gate1041(.a(gate559inter5), .b(gate559inter2), .O(gate559inter6));
  inv1  gate1042(.a(N1841), .O(gate559inter7));
  inv1  gate1043(.a(N1768), .O(gate559inter8));
  nand2 gate1044(.a(gate559inter8), .b(gate559inter7), .O(gate559inter9));
  nand2 gate1045(.a(s_23), .b(gate559inter3), .O(gate559inter10));
  nor2  gate1046(.a(gate559inter10), .b(gate559inter9), .O(gate559inter11));
  nor2  gate1047(.a(gate559inter11), .b(gate559inter6), .O(gate559inter12));
  nand2 gate1048(.a(gate559inter12), .b(gate559inter1), .O(N1882));
inv1 gate560( .a(N1841), .O(N1883) );

  xor2  gate1693(.a(N1852), .b(N1826), .O(gate561inter0));
  nand2 gate1694(.a(gate561inter0), .b(s_116), .O(gate561inter1));
  and2  gate1695(.a(N1852), .b(N1826), .O(gate561inter2));
  inv1  gate1696(.a(s_116), .O(gate561inter3));
  inv1  gate1697(.a(s_117), .O(gate561inter4));
  nand2 gate1698(.a(gate561inter4), .b(gate561inter3), .O(gate561inter5));
  nor2  gate1699(.a(gate561inter5), .b(gate561inter2), .O(gate561inter6));
  inv1  gate1700(.a(N1826), .O(gate561inter7));
  inv1  gate1701(.a(N1852), .O(gate561inter8));
  nand2 gate1702(.a(gate561inter8), .b(gate561inter7), .O(gate561inter9));
  nand2 gate1703(.a(s_117), .b(gate561inter3), .O(gate561inter10));
  nor2  gate1704(.a(gate561inter10), .b(gate561inter9), .O(gate561inter11));
  nor2  gate1705(.a(gate561inter11), .b(gate561inter6), .O(gate561inter12));
  nand2 gate1706(.a(gate561inter12), .b(gate561inter1), .O(N1884));
nand2 gate562( .a(N1643), .b(N1856), .O(N1885) );

  xor2  gate1119(.a(N290), .b(N1830), .O(gate563inter0));
  nand2 gate1120(.a(gate563inter0), .b(s_34), .O(gate563inter1));
  and2  gate1121(.a(N290), .b(N1830), .O(gate563inter2));
  inv1  gate1122(.a(s_34), .O(gate563inter3));
  inv1  gate1123(.a(s_35), .O(gate563inter4));
  nand2 gate1124(.a(gate563inter4), .b(gate563inter3), .O(gate563inter5));
  nor2  gate1125(.a(gate563inter5), .b(gate563inter2), .O(gate563inter6));
  inv1  gate1126(.a(N1830), .O(gate563inter7));
  inv1  gate1127(.a(N290), .O(gate563inter8));
  nand2 gate1128(.a(gate563inter8), .b(gate563inter7), .O(gate563inter9));
  nand2 gate1129(.a(s_35), .b(gate563inter3), .O(gate563inter10));
  nor2  gate1130(.a(gate563inter10), .b(gate563inter9), .O(gate563inter11));
  nor2  gate1131(.a(gate563inter11), .b(gate563inter6), .O(gate563inter12));
  nand2 gate1132(.a(gate563inter12), .b(gate563inter1), .O(N1889));
inv1 gate564( .a(N1838), .O(N1895) );
nand2 gate565( .a(N1838), .b(N1785), .O(N1896) );
nand2 gate566( .a(N1640), .b(N1864), .O(N1897) );
inv1 gate567( .a(N1850), .O(N1898) );
buf1 gate568( .a(N1830), .O(N1902) );
inv1 gate569( .a(N1878), .O(N1910) );
nand2 gate570( .a(N1717), .b(N1883), .O(N1911) );
inv1 gate571( .a(N1884), .O(N1912) );
nand2 gate572( .a(N1855), .b(N1885), .O(N1913) );
inv1 gate573( .a(N1866), .O(N1915) );

  xor2  gate1497(.a(N919), .b(N1872), .O(gate574inter0));
  nand2 gate1498(.a(gate574inter0), .b(s_88), .O(gate574inter1));
  and2  gate1499(.a(N919), .b(N1872), .O(gate574inter2));
  inv1  gate1500(.a(s_88), .O(gate574inter3));
  inv1  gate1501(.a(s_89), .O(gate574inter4));
  nand2 gate1502(.a(gate574inter4), .b(gate574inter3), .O(gate574inter5));
  nor2  gate1503(.a(gate574inter5), .b(gate574inter2), .O(gate574inter6));
  inv1  gate1504(.a(N1872), .O(gate574inter7));
  inv1  gate1505(.a(N919), .O(gate574inter8));
  nand2 gate1506(.a(gate574inter8), .b(gate574inter7), .O(gate574inter9));
  nand2 gate1507(.a(s_89), .b(gate574inter3), .O(gate574inter10));
  nor2  gate1508(.a(gate574inter10), .b(gate574inter9), .O(gate574inter11));
  nor2  gate1509(.a(gate574inter11), .b(gate574inter6), .O(gate574inter12));
  nand2 gate1510(.a(gate574inter12), .b(gate574inter1), .O(N1919));
inv1 gate575( .a(N1872), .O(N1920) );
nand2 gate576( .a(N1869), .b(N920), .O(N1921) );
inv1 gate577( .a(N1869), .O(N1922) );
inv1 gate578( .a(N1875), .O(N1923) );
nand2 gate579( .a(N1714), .b(N1895), .O(N1924) );
buf1 gate580( .a(N1858), .O(N1927) );
buf1 gate581( .a(N1858), .O(N1930) );
nand2 gate582( .a(N1865), .b(N1897), .O(N1933) );
nand2 gate583( .a(N1882), .b(N1911), .O(N1936) );
inv1 gate584( .a(N1898), .O(N1937) );
inv1 gate585( .a(N1902), .O(N1938) );
nand2 gate586( .a(N679), .b(N1920), .O(N1941) );
nand2 gate587( .a(N676), .b(N1922), .O(N1942) );
buf1 gate588( .a(N1879), .O(N1944) );
inv1 gate589( .a(N1913), .O(N1947) );
buf1 gate590( .a(N1889), .O(N1950) );
buf1 gate591( .a(N1889), .O(N1953) );
buf1 gate592( .a(N1879), .O(N1958) );
nand2 gate593( .a(N1896), .b(N1924), .O(N1961) );
and2 gate594( .a(N1910), .b(N601), .O(N1965) );
and2 gate595( .a(N602), .b(N1912), .O(N1968) );
nand2 gate596( .a(N1930), .b(N917), .O(N1975) );
inv1 gate597( .a(N1930), .O(N1976) );

  xor2  gate1483(.a(N918), .b(N1927), .O(gate598inter0));
  nand2 gate1484(.a(gate598inter0), .b(s_86), .O(gate598inter1));
  and2  gate1485(.a(N918), .b(N1927), .O(gate598inter2));
  inv1  gate1486(.a(s_86), .O(gate598inter3));
  inv1  gate1487(.a(s_87), .O(gate598inter4));
  nand2 gate1488(.a(gate598inter4), .b(gate598inter3), .O(gate598inter5));
  nor2  gate1489(.a(gate598inter5), .b(gate598inter2), .O(gate598inter6));
  inv1  gate1490(.a(N1927), .O(gate598inter7));
  inv1  gate1491(.a(N918), .O(gate598inter8));
  nand2 gate1492(.a(gate598inter8), .b(gate598inter7), .O(gate598inter9));
  nand2 gate1493(.a(s_87), .b(gate598inter3), .O(gate598inter10));
  nor2  gate1494(.a(gate598inter10), .b(gate598inter9), .O(gate598inter11));
  nor2  gate1495(.a(gate598inter11), .b(gate598inter6), .O(gate598inter12));
  nand2 gate1496(.a(gate598inter12), .b(gate598inter1), .O(N1977));
inv1 gate599( .a(N1927), .O(N1978) );

  xor2  gate1553(.a(N1941), .b(N1919), .O(gate600inter0));
  nand2 gate1554(.a(gate600inter0), .b(s_96), .O(gate600inter1));
  and2  gate1555(.a(N1941), .b(N1919), .O(gate600inter2));
  inv1  gate1556(.a(s_96), .O(gate600inter3));
  inv1  gate1557(.a(s_97), .O(gate600inter4));
  nand2 gate1558(.a(gate600inter4), .b(gate600inter3), .O(gate600inter5));
  nor2  gate1559(.a(gate600inter5), .b(gate600inter2), .O(gate600inter6));
  inv1  gate1560(.a(N1919), .O(gate600inter7));
  inv1  gate1561(.a(N1941), .O(gate600inter8));
  nand2 gate1562(.a(gate600inter8), .b(gate600inter7), .O(gate600inter9));
  nand2 gate1563(.a(s_97), .b(gate600inter3), .O(gate600inter10));
  nor2  gate1564(.a(gate600inter10), .b(gate600inter9), .O(gate600inter11));
  nor2  gate1565(.a(gate600inter11), .b(gate600inter6), .O(gate600inter12));
  nand2 gate1566(.a(gate600inter12), .b(gate600inter1), .O(N1979));

  xor2  gate1329(.a(N1942), .b(N1921), .O(gate601inter0));
  nand2 gate1330(.a(gate601inter0), .b(s_64), .O(gate601inter1));
  and2  gate1331(.a(N1942), .b(N1921), .O(gate601inter2));
  inv1  gate1332(.a(s_64), .O(gate601inter3));
  inv1  gate1333(.a(s_65), .O(gate601inter4));
  nand2 gate1334(.a(gate601inter4), .b(gate601inter3), .O(gate601inter5));
  nor2  gate1335(.a(gate601inter5), .b(gate601inter2), .O(gate601inter6));
  inv1  gate1336(.a(N1921), .O(gate601inter7));
  inv1  gate1337(.a(N1942), .O(gate601inter8));
  nand2 gate1338(.a(gate601inter8), .b(gate601inter7), .O(gate601inter9));
  nand2 gate1339(.a(s_65), .b(gate601inter3), .O(gate601inter10));
  nor2  gate1340(.a(gate601inter10), .b(gate601inter9), .O(gate601inter11));
  nor2  gate1341(.a(gate601inter11), .b(gate601inter6), .O(gate601inter12));
  nand2 gate1342(.a(gate601inter12), .b(gate601inter1), .O(N1980));
inv1 gate602( .a(N1933), .O(N1985) );
inv1 gate603( .a(N1936), .O(N1987) );
inv1 gate604( .a(N1944), .O(N1999) );
nand2 gate605( .a(N1944), .b(N1937), .O(N2000) );
inv1 gate606( .a(N1947), .O(N2002) );
nand2 gate607( .a(N1947), .b(N1499), .O(N2003) );
nand2 gate608( .a(N1953), .b(N1350), .O(N2004) );
inv1 gate609( .a(N1953), .O(N2005) );
nand2 gate610( .a(N1950), .b(N1351), .O(N2006) );
inv1 gate611( .a(N1950), .O(N2007) );
nand2 gate612( .a(N673), .b(N1976), .O(N2008) );
nand2 gate613( .a(N670), .b(N1978), .O(N2009) );
inv1 gate614( .a(N1979), .O(N2012) );
inv1 gate615( .a(N1958), .O(N2013) );
nand2 gate616( .a(N1958), .b(N1923), .O(N2014) );
inv1 gate617( .a(N1961), .O(N2015) );
nand2 gate618( .a(N1961), .b(N1635), .O(N2016) );
inv1 gate619( .a(N1965), .O(N2018) );
inv1 gate620( .a(N1968), .O(N2019) );
nand2 gate621( .a(N1898), .b(N1999), .O(N2020) );
inv1 gate622( .a(N1987), .O(N2021) );
nand2 gate623( .a(N1987), .b(N1591), .O(N2022) );
nand2 gate624( .a(N1440), .b(N2002), .O(N2023) );
nand2 gate625( .a(N1261), .b(N2005), .O(N2024) );

  xor2  gate1581(.a(N2007), .b(N1258), .O(gate626inter0));
  nand2 gate1582(.a(gate626inter0), .b(s_100), .O(gate626inter1));
  and2  gate1583(.a(N2007), .b(N1258), .O(gate626inter2));
  inv1  gate1584(.a(s_100), .O(gate626inter3));
  inv1  gate1585(.a(s_101), .O(gate626inter4));
  nand2 gate1586(.a(gate626inter4), .b(gate626inter3), .O(gate626inter5));
  nor2  gate1587(.a(gate626inter5), .b(gate626inter2), .O(gate626inter6));
  inv1  gate1588(.a(N1258), .O(gate626inter7));
  inv1  gate1589(.a(N2007), .O(gate626inter8));
  nand2 gate1590(.a(gate626inter8), .b(gate626inter7), .O(gate626inter9));
  nand2 gate1591(.a(s_101), .b(gate626inter3), .O(gate626inter10));
  nor2  gate1592(.a(gate626inter10), .b(gate626inter9), .O(gate626inter11));
  nor2  gate1593(.a(gate626inter11), .b(gate626inter6), .O(gate626inter12));
  nand2 gate1594(.a(gate626inter12), .b(gate626inter1), .O(N2025));

  xor2  gate1091(.a(N2008), .b(N1975), .O(gate627inter0));
  nand2 gate1092(.a(gate627inter0), .b(s_30), .O(gate627inter1));
  and2  gate1093(.a(N2008), .b(N1975), .O(gate627inter2));
  inv1  gate1094(.a(s_30), .O(gate627inter3));
  inv1  gate1095(.a(s_31), .O(gate627inter4));
  nand2 gate1096(.a(gate627inter4), .b(gate627inter3), .O(gate627inter5));
  nor2  gate1097(.a(gate627inter5), .b(gate627inter2), .O(gate627inter6));
  inv1  gate1098(.a(N1975), .O(gate627inter7));
  inv1  gate1099(.a(N2008), .O(gate627inter8));
  nand2 gate1100(.a(gate627inter8), .b(gate627inter7), .O(gate627inter9));
  nand2 gate1101(.a(s_31), .b(gate627inter3), .O(gate627inter10));
  nor2  gate1102(.a(gate627inter10), .b(gate627inter9), .O(gate627inter11));
  nor2  gate1103(.a(gate627inter11), .b(gate627inter6), .O(gate627inter12));
  nand2 gate1104(.a(gate627inter12), .b(gate627inter1), .O(N2026));

  xor2  gate895(.a(N2009), .b(N1977), .O(gate628inter0));
  nand2 gate896(.a(gate628inter0), .b(s_2), .O(gate628inter1));
  and2  gate897(.a(N2009), .b(N1977), .O(gate628inter2));
  inv1  gate898(.a(s_2), .O(gate628inter3));
  inv1  gate899(.a(s_3), .O(gate628inter4));
  nand2 gate900(.a(gate628inter4), .b(gate628inter3), .O(gate628inter5));
  nor2  gate901(.a(gate628inter5), .b(gate628inter2), .O(gate628inter6));
  inv1  gate902(.a(N1977), .O(gate628inter7));
  inv1  gate903(.a(N2009), .O(gate628inter8));
  nand2 gate904(.a(gate628inter8), .b(gate628inter7), .O(gate628inter9));
  nand2 gate905(.a(s_3), .b(gate628inter3), .O(gate628inter10));
  nor2  gate906(.a(gate628inter10), .b(gate628inter9), .O(gate628inter11));
  nor2  gate907(.a(gate628inter11), .b(gate628inter6), .O(gate628inter12));
  nand2 gate908(.a(gate628inter12), .b(gate628inter1), .O(N2027));
inv1 gate629( .a(N1980), .O(N2030) );
buf1 gate630( .a(N1980), .O(N2033) );
nand2 gate631( .a(N1875), .b(N2013), .O(N2036) );
nand2 gate632( .a(N1571), .b(N2015), .O(N2037) );
nand2 gate633( .a(N2020), .b(N2000), .O(N2038) );
nand2 gate634( .a(N1534), .b(N2021), .O(N2039) );
nand2 gate635( .a(N2023), .b(N2003), .O(N2040) );

  xor2  gate1343(.a(N2024), .b(N2004), .O(gate636inter0));
  nand2 gate1344(.a(gate636inter0), .b(s_66), .O(gate636inter1));
  and2  gate1345(.a(N2024), .b(N2004), .O(gate636inter2));
  inv1  gate1346(.a(s_66), .O(gate636inter3));
  inv1  gate1347(.a(s_67), .O(gate636inter4));
  nand2 gate1348(.a(gate636inter4), .b(gate636inter3), .O(gate636inter5));
  nor2  gate1349(.a(gate636inter5), .b(gate636inter2), .O(gate636inter6));
  inv1  gate1350(.a(N2004), .O(gate636inter7));
  inv1  gate1351(.a(N2024), .O(gate636inter8));
  nand2 gate1352(.a(gate636inter8), .b(gate636inter7), .O(gate636inter9));
  nand2 gate1353(.a(s_67), .b(gate636inter3), .O(gate636inter10));
  nor2  gate1354(.a(gate636inter10), .b(gate636inter9), .O(gate636inter11));
  nor2  gate1355(.a(gate636inter11), .b(gate636inter6), .O(gate636inter12));
  nand2 gate1356(.a(gate636inter12), .b(gate636inter1), .O(N2041));
nand2 gate637( .a(N2006), .b(N2025), .O(N2042) );
inv1 gate638( .a(N2026), .O(N2047) );
nand2 gate639( .a(N2036), .b(N2014), .O(N2052) );

  xor2  gate1357(.a(N2016), .b(N2037), .O(gate640inter0));
  nand2 gate1358(.a(gate640inter0), .b(s_68), .O(gate640inter1));
  and2  gate1359(.a(N2016), .b(N2037), .O(gate640inter2));
  inv1  gate1360(.a(s_68), .O(gate640inter3));
  inv1  gate1361(.a(s_69), .O(gate640inter4));
  nand2 gate1362(.a(gate640inter4), .b(gate640inter3), .O(gate640inter5));
  nor2  gate1363(.a(gate640inter5), .b(gate640inter2), .O(gate640inter6));
  inv1  gate1364(.a(N2037), .O(gate640inter7));
  inv1  gate1365(.a(N2016), .O(gate640inter8));
  nand2 gate1366(.a(gate640inter8), .b(gate640inter7), .O(gate640inter9));
  nand2 gate1367(.a(s_69), .b(gate640inter3), .O(gate640inter10));
  nor2  gate1368(.a(gate640inter10), .b(gate640inter9), .O(gate640inter11));
  nor2  gate1369(.a(gate640inter11), .b(gate640inter6), .O(gate640inter12));
  nand2 gate1370(.a(gate640inter12), .b(gate640inter1), .O(N2055));
inv1 gate641( .a(N2038), .O(N2060) );
nand2 gate642( .a(N2039), .b(N2022), .O(N2061) );
nand2 gate643( .a(N2040), .b(N290), .O(N2062) );
inv1 gate644( .a(N2041), .O(N2067) );
inv1 gate645( .a(N2027), .O(N2068) );
buf1 gate646( .a(N2027), .O(N2071) );
inv1 gate647( .a(N2052), .O(N2076) );
inv1 gate648( .a(N2055), .O(N2077) );
nand2 gate649( .a(N2060), .b(N290), .O(N2078) );
nand2 gate650( .a(N2061), .b(N290), .O(N2081) );
inv1 gate651( .a(N2042), .O(N2086) );
buf1 gate652( .a(N2042), .O(N2089) );
and2 gate653( .a(N2030), .b(N2068), .O(N2104) );
and2 gate654( .a(N2033), .b(N2068), .O(N2119) );
and2 gate655( .a(N2030), .b(N2071), .O(N2129) );
and2 gate656( .a(N2033), .b(N2071), .O(N2143) );
buf1 gate657( .a(N2062), .O(N2148) );
buf1 gate658( .a(N2062), .O(N2151) );
buf1 gate659( .a(N2078), .O(N2196) );
buf1 gate660( .a(N2078), .O(N2199) );
buf1 gate661( .a(N2081), .O(N2202) );
buf1 gate662( .a(N2081), .O(N2205) );
nand2 gate663( .a(N2151), .b(N915), .O(N2214) );
inv1 gate664( .a(N2151), .O(N2215) );
nand2 gate665( .a(N2148), .b(N916), .O(N2216) );
inv1 gate666( .a(N2148), .O(N2217) );

  xor2  gate979(.a(N1348), .b(N2199), .O(gate667inter0));
  nand2 gate980(.a(gate667inter0), .b(s_14), .O(gate667inter1));
  and2  gate981(.a(N1348), .b(N2199), .O(gate667inter2));
  inv1  gate982(.a(s_14), .O(gate667inter3));
  inv1  gate983(.a(s_15), .O(gate667inter4));
  nand2 gate984(.a(gate667inter4), .b(gate667inter3), .O(gate667inter5));
  nor2  gate985(.a(gate667inter5), .b(gate667inter2), .O(gate667inter6));
  inv1  gate986(.a(N2199), .O(gate667inter7));
  inv1  gate987(.a(N1348), .O(gate667inter8));
  nand2 gate988(.a(gate667inter8), .b(gate667inter7), .O(gate667inter9));
  nand2 gate989(.a(s_15), .b(gate667inter3), .O(gate667inter10));
  nor2  gate990(.a(gate667inter10), .b(gate667inter9), .O(gate667inter11));
  nor2  gate991(.a(gate667inter11), .b(gate667inter6), .O(gate667inter12));
  nand2 gate992(.a(gate667inter12), .b(gate667inter1), .O(N2222));
inv1 gate668( .a(N2199), .O(N2223) );
nand2 gate669( .a(N2196), .b(N1349), .O(N2224) );
inv1 gate670( .a(N2196), .O(N2225) );
nand2 gate671( .a(N2205), .b(N913), .O(N2226) );
inv1 gate672( .a(N2205), .O(N2227) );
nand2 gate673( .a(N2202), .b(N914), .O(N2228) );
inv1 gate674( .a(N2202), .O(N2229) );
nand2 gate675( .a(N667), .b(N2215), .O(N2230) );
nand2 gate676( .a(N664), .b(N2217), .O(N2231) );

  xor2  gate965(.a(N2223), .b(N1255), .O(gate677inter0));
  nand2 gate966(.a(gate677inter0), .b(s_12), .O(gate677inter1));
  and2  gate967(.a(N2223), .b(N1255), .O(gate677inter2));
  inv1  gate968(.a(s_12), .O(gate677inter3));
  inv1  gate969(.a(s_13), .O(gate677inter4));
  nand2 gate970(.a(gate677inter4), .b(gate677inter3), .O(gate677inter5));
  nor2  gate971(.a(gate677inter5), .b(gate677inter2), .O(gate677inter6));
  inv1  gate972(.a(N1255), .O(gate677inter7));
  inv1  gate973(.a(N2223), .O(gate677inter8));
  nand2 gate974(.a(gate677inter8), .b(gate677inter7), .O(gate677inter9));
  nand2 gate975(.a(s_13), .b(gate677inter3), .O(gate677inter10));
  nor2  gate976(.a(gate677inter10), .b(gate677inter9), .O(gate677inter11));
  nor2  gate977(.a(gate677inter11), .b(gate677inter6), .O(gate677inter12));
  nand2 gate978(.a(gate677inter12), .b(gate677inter1), .O(N2232));
nand2 gate678( .a(N1252), .b(N2225), .O(N2233) );
nand2 gate679( .a(N661), .b(N2227), .O(N2234) );
nand2 gate680( .a(N658), .b(N2229), .O(N2235) );
nand2 gate681( .a(N2214), .b(N2230), .O(N2236) );

  xor2  gate1637(.a(N2231), .b(N2216), .O(gate682inter0));
  nand2 gate1638(.a(gate682inter0), .b(s_108), .O(gate682inter1));
  and2  gate1639(.a(N2231), .b(N2216), .O(gate682inter2));
  inv1  gate1640(.a(s_108), .O(gate682inter3));
  inv1  gate1641(.a(s_109), .O(gate682inter4));
  nand2 gate1642(.a(gate682inter4), .b(gate682inter3), .O(gate682inter5));
  nor2  gate1643(.a(gate682inter5), .b(gate682inter2), .O(gate682inter6));
  inv1  gate1644(.a(N2216), .O(gate682inter7));
  inv1  gate1645(.a(N2231), .O(gate682inter8));
  nand2 gate1646(.a(gate682inter8), .b(gate682inter7), .O(gate682inter9));
  nand2 gate1647(.a(s_109), .b(gate682inter3), .O(gate682inter10));
  nor2  gate1648(.a(gate682inter10), .b(gate682inter9), .O(gate682inter11));
  nor2  gate1649(.a(gate682inter11), .b(gate682inter6), .O(gate682inter12));
  nand2 gate1650(.a(gate682inter12), .b(gate682inter1), .O(N2237));
nand2 gate683( .a(N2222), .b(N2232), .O(N2240) );

  xor2  gate1665(.a(N2233), .b(N2224), .O(gate684inter0));
  nand2 gate1666(.a(gate684inter0), .b(s_112), .O(gate684inter1));
  and2  gate1667(.a(N2233), .b(N2224), .O(gate684inter2));
  inv1  gate1668(.a(s_112), .O(gate684inter3));
  inv1  gate1669(.a(s_113), .O(gate684inter4));
  nand2 gate1670(.a(gate684inter4), .b(gate684inter3), .O(gate684inter5));
  nor2  gate1671(.a(gate684inter5), .b(gate684inter2), .O(gate684inter6));
  inv1  gate1672(.a(N2224), .O(gate684inter7));
  inv1  gate1673(.a(N2233), .O(gate684inter8));
  nand2 gate1674(.a(gate684inter8), .b(gate684inter7), .O(gate684inter9));
  nand2 gate1675(.a(s_113), .b(gate684inter3), .O(gate684inter10));
  nor2  gate1676(.a(gate684inter10), .b(gate684inter9), .O(gate684inter11));
  nor2  gate1677(.a(gate684inter11), .b(gate684inter6), .O(gate684inter12));
  nand2 gate1678(.a(gate684inter12), .b(gate684inter1), .O(N2241));
nand2 gate685( .a(N2226), .b(N2234), .O(N2244) );
nand2 gate686( .a(N2228), .b(N2235), .O(N2245) );
inv1 gate687( .a(N2236), .O(N2250) );
inv1 gate688( .a(N2240), .O(N2253) );
inv1 gate689( .a(N2244), .O(N2256) );
inv1 gate690( .a(N2237), .O(N2257) );
buf1 gate691( .a(N2237), .O(N2260) );
inv1 gate692( .a(N2241), .O(N2263) );
and2 gate693( .a(N1164), .b(N2241), .O(N2266) );
inv1 gate694( .a(N2245), .O(N2269) );
and2 gate695( .a(N1168), .b(N2245), .O(N2272) );
nand8 gate696( .a(N2067), .b(N2012), .c(N2047), .d(N2250), .e(N899), .f(N2256), .g(N2253), .h(N903), .O(N2279) );
buf1 gate697( .a(N2266), .O(N2286) );
buf1 gate698( .a(N2266), .O(N2297) );
buf1 gate699( .a(N2272), .O(N2315) );
buf1 gate700( .a(N2272), .O(N2326) );
and2 gate701( .a(N2086), .b(N2257), .O(N2340) );
and2 gate702( .a(N2089), .b(N2257), .O(N2353) );
and2 gate703( .a(N2086), .b(N2260), .O(N2361) );
and2 gate704( .a(N2089), .b(N2260), .O(N2375) );
and4 gate705( .a(N338), .b(N2279), .c(N313), .d(N313), .O(N2384) );
and2 gate706( .a(N1163), .b(N2263), .O(N2385) );
and2 gate707( .a(N1164), .b(N2263), .O(N2386) );
and2 gate708( .a(N1167), .b(N2269), .O(N2426) );
and2 gate709( .a(N1168), .b(N2269), .O(N2427) );
nand5 gate710( .a(N2286), .b(N2315), .c(N2361), .d(N2104), .e(N1171), .O(N2537) );
nand5 gate711( .a(N2286), .b(N2315), .c(N2340), .d(N2129), .e(N1171), .O(N2540) );
nand5 gate712( .a(N2286), .b(N2315), .c(N2340), .d(N2119), .e(N1171), .O(N2543) );
nand5 gate713( .a(N2286), .b(N2315), .c(N2353), .d(N2104), .e(N1171), .O(N2546) );
nand5 gate714( .a(N2297), .b(N2315), .c(N2375), .d(N2119), .e(N1188), .O(N2549) );
nand5 gate715( .a(N2297), .b(N2326), .c(N2361), .d(N2143), .e(N1188), .O(N2552) );
nand5 gate716( .a(N2297), .b(N2326), .c(N2375), .d(N2129), .e(N1188), .O(N2555) );
and5 gate717( .a(N2286), .b(N2315), .c(N2361), .d(N2104), .e(N1171), .O(N2558) );
and5 gate718( .a(N2286), .b(N2315), .c(N2340), .d(N2129), .e(N1171), .O(N2561) );
and5 gate719( .a(N2286), .b(N2315), .c(N2340), .d(N2119), .e(N1171), .O(N2564) );
and5 gate720( .a(N2286), .b(N2315), .c(N2353), .d(N2104), .e(N1171), .O(N2567) );
and5 gate721( .a(N2297), .b(N2315), .c(N2375), .d(N2119), .e(N1188), .O(N2570) );
and5 gate722( .a(N2297), .b(N2326), .c(N2361), .d(N2143), .e(N1188), .O(N2573) );
and5 gate723( .a(N2297), .b(N2326), .c(N2375), .d(N2129), .e(N1188), .O(N2576) );
nand5 gate724( .a(N2286), .b(N2427), .c(N2361), .d(N2129), .e(N1171), .O(N2594) );
nand5 gate725( .a(N2297), .b(N2427), .c(N2361), .d(N2119), .e(N1171), .O(N2597) );
nand5 gate726( .a(N2297), .b(N2427), .c(N2375), .d(N2104), .e(N1171), .O(N2600) );
nand5 gate727( .a(N2297), .b(N2427), .c(N2340), .d(N2143), .e(N1171), .O(N2603) );
nand5 gate728( .a(N2297), .b(N2427), .c(N2353), .d(N2129), .e(N1188), .O(N2606) );
nand5 gate729( .a(N2386), .b(N2326), .c(N2361), .d(N2129), .e(N1188), .O(N2611) );
nand5 gate730( .a(N2386), .b(N2326), .c(N2361), .d(N2119), .e(N1188), .O(N2614) );
nand5 gate731( .a(N2386), .b(N2326), .c(N2375), .d(N2104), .e(N1188), .O(N2617) );
nand5 gate732( .a(N2386), .b(N2326), .c(N2353), .d(N2129), .e(N1188), .O(N2620) );
nand5 gate733( .a(N2297), .b(N2427), .c(N2340), .d(N2104), .e(N926), .O(N2627) );
nand5 gate734( .a(N2386), .b(N2326), .c(N2340), .d(N2104), .e(N926), .O(N2628) );
nand5 gate735( .a(N2386), .b(N2427), .c(N2361), .d(N2104), .e(N926), .O(N2629) );
nand5 gate736( .a(N2386), .b(N2427), .c(N2340), .d(N2129), .e(N926), .O(N2630) );
nand5 gate737( .a(N2386), .b(N2427), .c(N2340), .d(N2119), .e(N926), .O(N2631) );
nand5 gate738( .a(N2386), .b(N2427), .c(N2353), .d(N2104), .e(N926), .O(N2632) );
nand5 gate739( .a(N2386), .b(N2426), .c(N2340), .d(N2104), .e(N926), .O(N2633) );
nand5 gate740( .a(N2385), .b(N2427), .c(N2340), .d(N2104), .e(N926), .O(N2634) );
and5 gate741( .a(N2286), .b(N2427), .c(N2361), .d(N2129), .e(N1171), .O(N2639) );
and5 gate742( .a(N2297), .b(N2427), .c(N2361), .d(N2119), .e(N1171), .O(N2642) );
and5 gate743( .a(N2297), .b(N2427), .c(N2375), .d(N2104), .e(N1171), .O(N2645) );
and5 gate744( .a(N2297), .b(N2427), .c(N2340), .d(N2143), .e(N1171), .O(N2648) );
and5 gate745( .a(N2297), .b(N2427), .c(N2353), .d(N2129), .e(N1188), .O(N2651) );
and5 gate746( .a(N2386), .b(N2326), .c(N2361), .d(N2129), .e(N1188), .O(N2655) );
and5 gate747( .a(N2386), .b(N2326), .c(N2361), .d(N2119), .e(N1188), .O(N2658) );
and5 gate748( .a(N2386), .b(N2326), .c(N2375), .d(N2104), .e(N1188), .O(N2661) );
and5 gate749( .a(N2386), .b(N2326), .c(N2353), .d(N2129), .e(N1188), .O(N2664) );

  xor2  gate881(.a(N534), .b(N2558), .O(gate750inter0));
  nand2 gate882(.a(gate750inter0), .b(s_0), .O(gate750inter1));
  and2  gate883(.a(N534), .b(N2558), .O(gate750inter2));
  inv1  gate884(.a(s_0), .O(gate750inter3));
  inv1  gate885(.a(s_1), .O(gate750inter4));
  nand2 gate886(.a(gate750inter4), .b(gate750inter3), .O(gate750inter5));
  nor2  gate887(.a(gate750inter5), .b(gate750inter2), .O(gate750inter6));
  inv1  gate888(.a(N2558), .O(gate750inter7));
  inv1  gate889(.a(N534), .O(gate750inter8));
  nand2 gate890(.a(gate750inter8), .b(gate750inter7), .O(gate750inter9));
  nand2 gate891(.a(s_1), .b(gate750inter3), .O(gate750inter10));
  nor2  gate892(.a(gate750inter10), .b(gate750inter9), .O(gate750inter11));
  nor2  gate893(.a(gate750inter11), .b(gate750inter6), .O(gate750inter12));
  nand2 gate894(.a(gate750inter12), .b(gate750inter1), .O(N2669));
inv1 gate751( .a(N2558), .O(N2670) );
nand2 gate752( .a(N2561), .b(N535), .O(N2671) );
inv1 gate753( .a(N2561), .O(N2672) );
nand2 gate754( .a(N2564), .b(N536), .O(N2673) );
inv1 gate755( .a(N2564), .O(N2674) );
nand2 gate756( .a(N2567), .b(N537), .O(N2675) );
inv1 gate757( .a(N2567), .O(N2676) );
nand2 gate758( .a(N2570), .b(N543), .O(N2682) );
inv1 gate759( .a(N2570), .O(N2683) );
nand2 gate760( .a(N2573), .b(N548), .O(N2688) );
inv1 gate761( .a(N2573), .O(N2689) );
nand2 gate762( .a(N2576), .b(N549), .O(N2690) );
inv1 gate763( .a(N2576), .O(N2691) );
and8 gate764( .a(N2627), .b(N2628), .c(N2629), .d(N2630), .e(N2631), .f(N2632), .g(N2633), .h(N2634), .O(N2710) );
nand2 gate765( .a(N343), .b(N2670), .O(N2720) );

  xor2  gate1791(.a(N2672), .b(N346), .O(gate766inter0));
  nand2 gate1792(.a(gate766inter0), .b(s_130), .O(gate766inter1));
  and2  gate1793(.a(N2672), .b(N346), .O(gate766inter2));
  inv1  gate1794(.a(s_130), .O(gate766inter3));
  inv1  gate1795(.a(s_131), .O(gate766inter4));
  nand2 gate1796(.a(gate766inter4), .b(gate766inter3), .O(gate766inter5));
  nor2  gate1797(.a(gate766inter5), .b(gate766inter2), .O(gate766inter6));
  inv1  gate1798(.a(N346), .O(gate766inter7));
  inv1  gate1799(.a(N2672), .O(gate766inter8));
  nand2 gate1800(.a(gate766inter8), .b(gate766inter7), .O(gate766inter9));
  nand2 gate1801(.a(s_131), .b(gate766inter3), .O(gate766inter10));
  nor2  gate1802(.a(gate766inter10), .b(gate766inter9), .O(gate766inter11));
  nor2  gate1803(.a(gate766inter11), .b(gate766inter6), .O(gate766inter12));
  nand2 gate1804(.a(gate766inter12), .b(gate766inter1), .O(N2721));

  xor2  gate1105(.a(N2674), .b(N349), .O(gate767inter0));
  nand2 gate1106(.a(gate767inter0), .b(s_32), .O(gate767inter1));
  and2  gate1107(.a(N2674), .b(N349), .O(gate767inter2));
  inv1  gate1108(.a(s_32), .O(gate767inter3));
  inv1  gate1109(.a(s_33), .O(gate767inter4));
  nand2 gate1110(.a(gate767inter4), .b(gate767inter3), .O(gate767inter5));
  nor2  gate1111(.a(gate767inter5), .b(gate767inter2), .O(gate767inter6));
  inv1  gate1112(.a(N349), .O(gate767inter7));
  inv1  gate1113(.a(N2674), .O(gate767inter8));
  nand2 gate1114(.a(gate767inter8), .b(gate767inter7), .O(gate767inter9));
  nand2 gate1115(.a(s_33), .b(gate767inter3), .O(gate767inter10));
  nor2  gate1116(.a(gate767inter10), .b(gate767inter9), .O(gate767inter11));
  nor2  gate1117(.a(gate767inter11), .b(gate767inter6), .O(gate767inter12));
  nand2 gate1118(.a(gate767inter12), .b(gate767inter1), .O(N2722));
nand2 gate768( .a(N352), .b(N2676), .O(N2723) );
nand2 gate769( .a(N2639), .b(N538), .O(N2724) );
inv1 gate770( .a(N2639), .O(N2725) );
nand2 gate771( .a(N2642), .b(N539), .O(N2726) );
inv1 gate772( .a(N2642), .O(N2727) );
nand2 gate773( .a(N2645), .b(N540), .O(N2728) );
inv1 gate774( .a(N2645), .O(N2729) );

  xor2  gate1609(.a(N541), .b(N2648), .O(gate775inter0));
  nand2 gate1610(.a(gate775inter0), .b(s_104), .O(gate775inter1));
  and2  gate1611(.a(N541), .b(N2648), .O(gate775inter2));
  inv1  gate1612(.a(s_104), .O(gate775inter3));
  inv1  gate1613(.a(s_105), .O(gate775inter4));
  nand2 gate1614(.a(gate775inter4), .b(gate775inter3), .O(gate775inter5));
  nor2  gate1615(.a(gate775inter5), .b(gate775inter2), .O(gate775inter6));
  inv1  gate1616(.a(N2648), .O(gate775inter7));
  inv1  gate1617(.a(N541), .O(gate775inter8));
  nand2 gate1618(.a(gate775inter8), .b(gate775inter7), .O(gate775inter9));
  nand2 gate1619(.a(s_105), .b(gate775inter3), .O(gate775inter10));
  nor2  gate1620(.a(gate775inter10), .b(gate775inter9), .O(gate775inter11));
  nor2  gate1621(.a(gate775inter11), .b(gate775inter6), .O(gate775inter12));
  nand2 gate1622(.a(gate775inter12), .b(gate775inter1), .O(N2730));
inv1 gate776( .a(N2648), .O(N2731) );

  xor2  gate1259(.a(N542), .b(N2651), .O(gate777inter0));
  nand2 gate1260(.a(gate777inter0), .b(s_54), .O(gate777inter1));
  and2  gate1261(.a(N542), .b(N2651), .O(gate777inter2));
  inv1  gate1262(.a(s_54), .O(gate777inter3));
  inv1  gate1263(.a(s_55), .O(gate777inter4));
  nand2 gate1264(.a(gate777inter4), .b(gate777inter3), .O(gate777inter5));
  nor2  gate1265(.a(gate777inter5), .b(gate777inter2), .O(gate777inter6));
  inv1  gate1266(.a(N2651), .O(gate777inter7));
  inv1  gate1267(.a(N542), .O(gate777inter8));
  nand2 gate1268(.a(gate777inter8), .b(gate777inter7), .O(gate777inter9));
  nand2 gate1269(.a(s_55), .b(gate777inter3), .O(gate777inter10));
  nor2  gate1270(.a(gate777inter10), .b(gate777inter9), .O(gate777inter11));
  nor2  gate1271(.a(gate777inter11), .b(gate777inter6), .O(gate777inter12));
  nand2 gate1272(.a(gate777inter12), .b(gate777inter1), .O(N2732));
inv1 gate778( .a(N2651), .O(N2733) );
nand2 gate779( .a(N370), .b(N2683), .O(N2734) );

  xor2  gate1063(.a(N544), .b(N2655), .O(gate780inter0));
  nand2 gate1064(.a(gate780inter0), .b(s_26), .O(gate780inter1));
  and2  gate1065(.a(N544), .b(N2655), .O(gate780inter2));
  inv1  gate1066(.a(s_26), .O(gate780inter3));
  inv1  gate1067(.a(s_27), .O(gate780inter4));
  nand2 gate1068(.a(gate780inter4), .b(gate780inter3), .O(gate780inter5));
  nor2  gate1069(.a(gate780inter5), .b(gate780inter2), .O(gate780inter6));
  inv1  gate1070(.a(N2655), .O(gate780inter7));
  inv1  gate1071(.a(N544), .O(gate780inter8));
  nand2 gate1072(.a(gate780inter8), .b(gate780inter7), .O(gate780inter9));
  nand2 gate1073(.a(s_27), .b(gate780inter3), .O(gate780inter10));
  nor2  gate1074(.a(gate780inter10), .b(gate780inter9), .O(gate780inter11));
  nor2  gate1075(.a(gate780inter11), .b(gate780inter6), .O(gate780inter12));
  nand2 gate1076(.a(gate780inter12), .b(gate780inter1), .O(N2735));
inv1 gate781( .a(N2655), .O(N2736) );
nand2 gate782( .a(N2658), .b(N545), .O(N2737) );
inv1 gate783( .a(N2658), .O(N2738) );
nand2 gate784( .a(N2661), .b(N546), .O(N2739) );
inv1 gate785( .a(N2661), .O(N2740) );
nand2 gate786( .a(N2664), .b(N547), .O(N2741) );
inv1 gate787( .a(N2664), .O(N2742) );
nand2 gate788( .a(N385), .b(N2689), .O(N2743) );
nand2 gate789( .a(N388), .b(N2691), .O(N2744) );
nand8 gate790( .a(N2537), .b(N2540), .c(N2543), .d(N2546), .e(N2594), .f(N2597), .g(N2600), .h(N2603), .O(N2745) );
nand8 gate791( .a(N2606), .b(N2549), .c(N2611), .d(N2614), .e(N2617), .f(N2620), .g(N2552), .h(N2555), .O(N2746) );
and8 gate792( .a(N2537), .b(N2540), .c(N2543), .d(N2546), .e(N2594), .f(N2597), .g(N2600), .h(N2603), .O(N2747) );
and8 gate793( .a(N2606), .b(N2549), .c(N2611), .d(N2614), .e(N2617), .f(N2620), .g(N2552), .h(N2555), .O(N2750) );
nand2 gate794( .a(N2669), .b(N2720), .O(N2753) );
nand2 gate795( .a(N2671), .b(N2721), .O(N2754) );
nand2 gate796( .a(N2673), .b(N2722), .O(N2755) );
nand2 gate797( .a(N2675), .b(N2723), .O(N2756) );
nand2 gate798( .a(N355), .b(N2725), .O(N2757) );
nand2 gate799( .a(N358), .b(N2727), .O(N2758) );
nand2 gate800( .a(N361), .b(N2729), .O(N2759) );
nand2 gate801( .a(N364), .b(N2731), .O(N2760) );
nand2 gate802( .a(N367), .b(N2733), .O(N2761) );
nand2 gate803( .a(N2682), .b(N2734), .O(N2762) );
nand2 gate804( .a(N373), .b(N2736), .O(N2763) );
nand2 gate805( .a(N376), .b(N2738), .O(N2764) );
nand2 gate806( .a(N379), .b(N2740), .O(N2765) );
nand2 gate807( .a(N382), .b(N2742), .O(N2766) );
nand2 gate808( .a(N2688), .b(N2743), .O(N2767) );
nand2 gate809( .a(N2690), .b(N2744), .O(N2768) );
and2 gate810( .a(N2745), .b(N275), .O(N2773) );
and2 gate811( .a(N2746), .b(N276), .O(N2776) );
nand2 gate812( .a(N2724), .b(N2757), .O(N2779) );
nand2 gate813( .a(N2726), .b(N2758), .O(N2780) );
nand2 gate814( .a(N2728), .b(N2759), .O(N2781) );

  xor2  gate1315(.a(N2760), .b(N2730), .O(gate815inter0));
  nand2 gate1316(.a(gate815inter0), .b(s_62), .O(gate815inter1));
  and2  gate1317(.a(N2760), .b(N2730), .O(gate815inter2));
  inv1  gate1318(.a(s_62), .O(gate815inter3));
  inv1  gate1319(.a(s_63), .O(gate815inter4));
  nand2 gate1320(.a(gate815inter4), .b(gate815inter3), .O(gate815inter5));
  nor2  gate1321(.a(gate815inter5), .b(gate815inter2), .O(gate815inter6));
  inv1  gate1322(.a(N2730), .O(gate815inter7));
  inv1  gate1323(.a(N2760), .O(gate815inter8));
  nand2 gate1324(.a(gate815inter8), .b(gate815inter7), .O(gate815inter9));
  nand2 gate1325(.a(s_63), .b(gate815inter3), .O(gate815inter10));
  nor2  gate1326(.a(gate815inter10), .b(gate815inter9), .O(gate815inter11));
  nor2  gate1327(.a(gate815inter11), .b(gate815inter6), .O(gate815inter12));
  nand2 gate1328(.a(gate815inter12), .b(gate815inter1), .O(N2782));
nand2 gate816( .a(N2732), .b(N2761), .O(N2783) );
nand2 gate817( .a(N2735), .b(N2763), .O(N2784) );
nand2 gate818( .a(N2737), .b(N2764), .O(N2785) );
nand2 gate819( .a(N2739), .b(N2765), .O(N2786) );
nand2 gate820( .a(N2741), .b(N2766), .O(N2787) );
and3 gate821( .a(N2747), .b(N2750), .c(N2710), .O(N2788) );

  xor2  gate1749(.a(N2750), .b(N2747), .O(gate822inter0));
  nand2 gate1750(.a(gate822inter0), .b(s_124), .O(gate822inter1));
  and2  gate1751(.a(N2750), .b(N2747), .O(gate822inter2));
  inv1  gate1752(.a(s_124), .O(gate822inter3));
  inv1  gate1753(.a(s_125), .O(gate822inter4));
  nand2 gate1754(.a(gate822inter4), .b(gate822inter3), .O(gate822inter5));
  nor2  gate1755(.a(gate822inter5), .b(gate822inter2), .O(gate822inter6));
  inv1  gate1756(.a(N2747), .O(gate822inter7));
  inv1  gate1757(.a(N2750), .O(gate822inter8));
  nand2 gate1758(.a(gate822inter8), .b(gate822inter7), .O(gate822inter9));
  nand2 gate1759(.a(s_125), .b(gate822inter3), .O(gate822inter10));
  nor2  gate1760(.a(gate822inter10), .b(gate822inter9), .O(gate822inter11));
  nor2  gate1761(.a(gate822inter11), .b(gate822inter6), .O(gate822inter12));
  nand2 gate1762(.a(gate822inter12), .b(gate822inter1), .O(N2789));
and4 gate823( .a(N338), .b(N2279), .c(N99), .d(N2788), .O(N2800) );
nand2 gate824( .a(N2773), .b(N2018), .O(N2807) );
inv1 gate825( .a(N2773), .O(N2808) );
nand2 gate826( .a(N2776), .b(N2019), .O(N2809) );
inv1 gate827( .a(N2776), .O(N2810) );

  xor2  gate1623(.a(N2800), .b(N2384), .O(gate828inter0));
  nand2 gate1624(.a(gate828inter0), .b(s_106), .O(gate828inter1));
  and2  gate1625(.a(N2800), .b(N2384), .O(gate828inter2));
  inv1  gate1626(.a(s_106), .O(gate828inter3));
  inv1  gate1627(.a(s_107), .O(gate828inter4));
  nand2 gate1628(.a(gate828inter4), .b(gate828inter3), .O(gate828inter5));
  nor2  gate1629(.a(gate828inter5), .b(gate828inter2), .O(gate828inter6));
  inv1  gate1630(.a(N2384), .O(gate828inter7));
  inv1  gate1631(.a(N2800), .O(gate828inter8));
  nand2 gate1632(.a(gate828inter8), .b(gate828inter7), .O(gate828inter9));
  nand2 gate1633(.a(s_107), .b(gate828inter3), .O(gate828inter10));
  nor2  gate1634(.a(gate828inter10), .b(gate828inter9), .O(gate828inter11));
  nor2  gate1635(.a(gate828inter11), .b(gate828inter6), .O(gate828inter12));
  nand2 gate1636(.a(gate828inter12), .b(gate828inter1), .O(N2811));
and3 gate829( .a(N897), .b(N283), .c(N2789), .O(N2812) );
and3 gate830( .a(N76), .b(N283), .c(N2789), .O(N2815) );
and3 gate831( .a(N82), .b(N283), .c(N2789), .O(N2818) );
and3 gate832( .a(N85), .b(N283), .c(N2789), .O(N2821) );
and3 gate833( .a(N898), .b(N283), .c(N2789), .O(N2824) );
nand2 gate834( .a(N1965), .b(N2808), .O(N2827) );
nand2 gate835( .a(N1968), .b(N2810), .O(N2828) );
and3 gate836( .a(N79), .b(N283), .c(N2789), .O(N2829) );
nand2 gate837( .a(N2807), .b(N2827), .O(N2843) );
nand2 gate838( .a(N2809), .b(N2828), .O(N2846) );
nand2 gate839( .a(N2812), .b(N2076), .O(N2850) );
nand2 gate840( .a(N2815), .b(N2077), .O(N2851) );
nand2 gate841( .a(N2818), .b(N1915), .O(N2852) );
nand2 gate842( .a(N2821), .b(N1857), .O(N2853) );
nand2 gate843( .a(N2824), .b(N1938), .O(N2854) );
inv1 gate844( .a(N2812), .O(N2857) );
inv1 gate845( .a(N2815), .O(N2858) );
inv1 gate846( .a(N2818), .O(N2859) );
inv1 gate847( .a(N2821), .O(N2860) );
inv1 gate848( .a(N2824), .O(N2861) );
inv1 gate849( .a(N2829), .O(N2862) );
nand2 gate850( .a(N2829), .b(N1985), .O(N2863) );
nand2 gate851( .a(N2052), .b(N2857), .O(N2866) );
nand2 gate852( .a(N2055), .b(N2858), .O(N2867) );
nand2 gate853( .a(N1866), .b(N2859), .O(N2868) );

  xor2  gate1707(.a(N2860), .b(N1818), .O(gate854inter0));
  nand2 gate1708(.a(gate854inter0), .b(s_118), .O(gate854inter1));
  and2  gate1709(.a(N2860), .b(N1818), .O(gate854inter2));
  inv1  gate1710(.a(s_118), .O(gate854inter3));
  inv1  gate1711(.a(s_119), .O(gate854inter4));
  nand2 gate1712(.a(gate854inter4), .b(gate854inter3), .O(gate854inter5));
  nor2  gate1713(.a(gate854inter5), .b(gate854inter2), .O(gate854inter6));
  inv1  gate1714(.a(N1818), .O(gate854inter7));
  inv1  gate1715(.a(N2860), .O(gate854inter8));
  nand2 gate1716(.a(gate854inter8), .b(gate854inter7), .O(gate854inter9));
  nand2 gate1717(.a(s_119), .b(gate854inter3), .O(gate854inter10));
  nor2  gate1718(.a(gate854inter10), .b(gate854inter9), .O(gate854inter11));
  nor2  gate1719(.a(gate854inter11), .b(gate854inter6), .O(gate854inter12));
  nand2 gate1720(.a(gate854inter12), .b(gate854inter1), .O(N2869));
nand2 gate855( .a(N1902), .b(N2861), .O(N2870) );
nand2 gate856( .a(N2843), .b(N886), .O(N2871) );
inv1 gate857( .a(N2843), .O(N2872) );
nand2 gate858( .a(N2846), .b(N887), .O(N2873) );
inv1 gate859( .a(N2846), .O(N2874) );

  xor2  gate1385(.a(N2862), .b(N1933), .O(gate860inter0));
  nand2 gate1386(.a(gate860inter0), .b(s_72), .O(gate860inter1));
  and2  gate1387(.a(N2862), .b(N1933), .O(gate860inter2));
  inv1  gate1388(.a(s_72), .O(gate860inter3));
  inv1  gate1389(.a(s_73), .O(gate860inter4));
  nand2 gate1390(.a(gate860inter4), .b(gate860inter3), .O(gate860inter5));
  nor2  gate1391(.a(gate860inter5), .b(gate860inter2), .O(gate860inter6));
  inv1  gate1392(.a(N1933), .O(gate860inter7));
  inv1  gate1393(.a(N2862), .O(gate860inter8));
  nand2 gate1394(.a(gate860inter8), .b(gate860inter7), .O(gate860inter9));
  nand2 gate1395(.a(s_73), .b(gate860inter3), .O(gate860inter10));
  nor2  gate1396(.a(gate860inter10), .b(gate860inter9), .O(gate860inter11));
  nor2  gate1397(.a(gate860inter11), .b(gate860inter6), .O(gate860inter12));
  nand2 gate1398(.a(gate860inter12), .b(gate860inter1), .O(N2875));
nand2 gate861( .a(N2866), .b(N2850), .O(N2876) );
nand2 gate862( .a(N2867), .b(N2851), .O(N2877) );
nand2 gate863( .a(N2868), .b(N2852), .O(N2878) );
nand2 gate864( .a(N2869), .b(N2853), .O(N2879) );
nand2 gate865( .a(N2870), .b(N2854), .O(N2880) );
nand2 gate866( .a(N682), .b(N2872), .O(N2881) );
nand2 gate867( .a(N685), .b(N2874), .O(N2882) );
nand2 gate868( .a(N2875), .b(N2863), .O(N2883) );
and2 gate869( .a(N2876), .b(N550), .O(N2886) );
and2 gate870( .a(N551), .b(N2877), .O(N2887) );
and2 gate871( .a(N553), .b(N2878), .O(N2888) );
and2 gate872( .a(N2879), .b(N554), .O(N2889) );
and2 gate873( .a(N555), .b(N2880), .O(N2890) );
nand2 gate874( .a(N2871), .b(N2881), .O(N2891) );

  xor2  gate1651(.a(N2882), .b(N2873), .O(gate875inter0));
  nand2 gate1652(.a(gate875inter0), .b(s_110), .O(gate875inter1));
  and2  gate1653(.a(N2882), .b(N2873), .O(gate875inter2));
  inv1  gate1654(.a(s_110), .O(gate875inter3));
  inv1  gate1655(.a(s_111), .O(gate875inter4));
  nand2 gate1656(.a(gate875inter4), .b(gate875inter3), .O(gate875inter5));
  nor2  gate1657(.a(gate875inter5), .b(gate875inter2), .O(gate875inter6));
  inv1  gate1658(.a(N2873), .O(gate875inter7));
  inv1  gate1659(.a(N2882), .O(gate875inter8));
  nand2 gate1660(.a(gate875inter8), .b(gate875inter7), .O(gate875inter9));
  nand2 gate1661(.a(s_111), .b(gate875inter3), .O(gate875inter10));
  nor2  gate1662(.a(gate875inter10), .b(gate875inter9), .O(gate875inter11));
  nor2  gate1663(.a(gate875inter11), .b(gate875inter6), .O(gate875inter12));
  nand2 gate1664(.a(gate875inter12), .b(gate875inter1), .O(N2892));
nand2 gate876( .a(N2883), .b(N1461), .O(N2895) );
inv1 gate877( .a(N2883), .O(N2896) );
nand2 gate878( .a(N1383), .b(N2896), .O(N2897) );
nand2 gate879( .a(N2895), .b(N2897), .O(N2898) );
and2 gate880( .a(N2898), .b(N552), .O(N2899) );

endmodule