module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);

input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;//RE__PI;

input s_0,s_1;//RE__ALLOW(00,01,10,11);
input s_2,s_3;//RE__ALLOW(00,01,10,11);
input s_4,s_5;//RE__ALLOW(00,01,10,11);
input s_6,s_7;//RE__ALLOW(00,01,10,11);
input s_8,s_9;//RE__ALLOW(00,01,10,11);
input s_10,s_11;//RE__ALLOW(00,01,10,11);
input s_12,s_13;//RE__ALLOW(00,01,10,11);
input s_14,s_15;//RE__ALLOW(00,01,10,11);
input s_16,s_17;//RE__ALLOW(00,01,10,11);
input s_18,s_19;//RE__ALLOW(00,01,10,11);
input s_20,s_21;//RE__ALLOW(00,01,10,11);
input s_22,s_23;//RE__ALLOW(00,01,10,11);
input s_24,s_25;//RE__ALLOW(00,01,10,11);
input s_26,s_27;//RE__ALLOW(00,01,10,11);
input s_28,s_29;//RE__ALLOW(00,01,10,11);
input s_30,s_31;//RE__ALLOW(00,01,10,11);
input s_32,s_33;//RE__ALLOW(00,01,10,11);
input s_34,s_35;//RE__ALLOW(00,01,10,11);
input s_36,s_37;//RE__ALLOW(00,01,10,11);
input s_38,s_39;//RE__ALLOW(00,01,10,11);
input s_40,s_41;//RE__ALLOW(00,01,10,11);
input s_42,s_43;//RE__ALLOW(00,01,10,11);
input s_44,s_45;//RE__ALLOW(00,01,10,11);
input s_46,s_47;//RE__ALLOW(00,01,10,11);
input s_48,s_49;//RE__ALLOW(00,01,10,11);
input s_50,s_51;//RE__ALLOW(00,01,10,11);
input s_52,s_53;//RE__ALLOW(00,01,10,11);
input s_54,s_55;//RE__ALLOW(00,01,10,11);
input s_56,s_57;//RE__ALLOW(00,01,10,11);
input s_58,s_59;//RE__ALLOW(00,01,10,11);
input s_60,s_61;//RE__ALLOW(00,01,10,11);
input s_62,s_63;//RE__ALLOW(00,01,10,11);
input s_64,s_65;//RE__ALLOW(00,01,10,11);
input s_66,s_67;//RE__ALLOW(00,01,10,11);
input s_68,s_69;//RE__ALLOW(00,01,10,11);
input s_70,s_71;//RE__ALLOW(00,01,10,11);
input s_72,s_73;//RE__ALLOW(00,01,10,11);
input s_74,s_75;//RE__ALLOW(00,01,10,11);
input s_76,s_77;//RE__ALLOW(00,01,10,11);
input s_78,s_79;//RE__ALLOW(00,01,10,11);
input s_80,s_81;//RE__ALLOW(00,01,10,11);
input s_82,s_83;//RE__ALLOW(00,01,10,11);
input s_84,s_85;//RE__ALLOW(00,01,10,11);
input s_86,s_87;//RE__ALLOW(00,01,10,11);
input s_88,s_89;//RE__ALLOW(00,01,10,11);
input s_90,s_91;//RE__ALLOW(00,01,10,11);
input s_92,s_93;//RE__ALLOW(00,01,10,11);
input s_94,s_95;//RE__ALLOW(00,01,10,11);
input s_96,s_97;//RE__ALLOW(00,01,10,11);
input s_98,s_99;//RE__ALLOW(00,01,10,11);
input s_100,s_101;//RE__ALLOW(00,01,10,11);
input s_102,s_103;//RE__ALLOW(00,01,10,11);
input s_104,s_105;//RE__ALLOW(00,01,10,11);
input s_106,s_107;//RE__ALLOW(00,01,10,11);
input s_108,s_109;//RE__ALLOW(00,01,10,11);
input s_110,s_111;//RE__ALLOW(00,01,10,11);
input s_112,s_113;//RE__ALLOW(00,01,10,11);
input s_114,s_115;//RE__ALLOW(00,01,10,11);
input s_116,s_117;//RE__ALLOW(00,01,10,11);
input s_118,s_119;//RE__ALLOW(00,01,10,11);
input s_120,s_121;//RE__ALLOW(00,01,10,11);
input s_122,s_123;//RE__ALLOW(00,01,10,11);
input s_124,s_125;//RE__ALLOW(00,01,10,11);
input s_126,s_127;//RE__ALLOW(00,01,10,11);
input s_128,s_129;//RE__ALLOW(00,01,10,11);
input s_130,s_131;//RE__ALLOW(00,01,10,11);
input s_132,s_133;//RE__ALLOW(00,01,10,11);
input s_134,s_135;//RE__ALLOW(00,01,10,11);
input s_136,s_137;//RE__ALLOW(00,01,10,11);
input s_138,s_139;//RE__ALLOW(00,01,10,11);
input s_140,s_141;//RE__ALLOW(00,01,10,11);
input s_142,s_143;//RE__ALLOW(00,01,10,11);
input s_144,s_145;//RE__ALLOW(00,01,10,11);
input s_146,s_147;//RE__ALLOW(00,01,10,11);
input s_148,s_149;//RE__ALLOW(00,01,10,11);
input s_150,s_151;//RE__ALLOW(00,01,10,11);
input s_152,s_153;//RE__ALLOW(00,01,10,11);
input s_154,s_155;//RE__ALLOW(00,01,10,11);
input s_156,s_157;//RE__ALLOW(00,01,10,11);
input s_158,s_159;//RE__ALLOW(00,01,10,11);
input s_160,s_161;//RE__ALLOW(00,01,10,11);
input s_162,s_163;//RE__ALLOW(00,01,10,11);
input s_164,s_165;//RE__ALLOW(00,01,10,11);
input s_166,s_167;//RE__ALLOW(00,01,10,11);
input s_168,s_169;//RE__ALLOW(00,01,10,11);
input s_170,s_171;//RE__ALLOW(00,01,10,11);
input s_172,s_173;//RE__ALLOW(00,01,10,11);
input s_174,s_175;//RE__ALLOW(00,01,10,11);
input s_176,s_177;//RE__ALLOW(00,01,10,11);
input s_178,s_179;//RE__ALLOW(00,01,10,11);
input s_180,s_181;//RE__ALLOW(00,01,10,11);
input s_182,s_183;//RE__ALLOW(00,01,10,11);
input s_184,s_185;//RE__ALLOW(00,01,10,11);
input s_186,s_187;//RE__ALLOW(00,01,10,11);
input s_188,s_189;//RE__ALLOW(00,01,10,11);
input s_190,s_191;//RE__ALLOW(00,01,10,11);
input s_192,s_193;//RE__ALLOW(00,01,10,11);
input s_194,s_195;//RE__ALLOW(00,01,10,11);
input s_196,s_197;//RE__ALLOW(00,01,10,11);
input s_198,s_199;//RE__ALLOW(00,01,10,11);
input s_200,s_201;//RE__ALLOW(00,01,10,11);
input s_202,s_203;//RE__ALLOW(00,01,10,11);
input s_204,s_205;//RE__ALLOW(00,01,10,11);
input s_206,s_207;//RE__ALLOW(00,01,10,11);
input s_208,s_209;//RE__ALLOW(00,01,10,11);
input s_210,s_211;//RE__ALLOW(00,01,10,11);
input s_212,s_213;//RE__ALLOW(00,01,10,11);
input s_214,s_215;//RE__ALLOW(00,01,10,11);
input s_216,s_217;//RE__ALLOW(00,01,10,11);
input s_218,s_219;//RE__ALLOW(00,01,10,11);
input s_220,s_221;//RE__ALLOW(00,01,10,11);
input s_222,s_223;//RE__ALLOW(00,01,10,11);
input s_224,s_225;//RE__ALLOW(00,01,10,11);
input s_226,s_227;//RE__ALLOW(00,01,10,11);
input s_228,s_229;//RE__ALLOW(00,01,10,11);
input s_230,s_231;//RE__ALLOW(00,01,10,11);
input s_232,s_233;//RE__ALLOW(00,01,10,11);
input s_234,s_235;//RE__ALLOW(00,01,10,11);
input s_236,s_237;//RE__ALLOW(00,01,10,11);
input s_238,s_239;//RE__ALLOW(00,01,10,11);
input s_240,s_241;//RE__ALLOW(00,01,10,11);
input s_242,s_243;//RE__ALLOW(00,01,10,11);
input s_244,s_245;//RE__ALLOW(00,01,10,11);
input s_246,s_247;//RE__ALLOW(00,01,10,11);
input s_248,s_249;//RE__ALLOW(00,01,10,11);
input s_250,s_251;//RE__ALLOW(00,01,10,11);
input s_252,s_253;//RE__ALLOW(00,01,10,11);
input s_254,s_255;//RE__ALLOW(00,01,10,11);
input s_256,s_257;//RE__ALLOW(00,01,10,11);
input s_258,s_259;//RE__ALLOW(00,01,10,11);
input s_260,s_261;//RE__ALLOW(00,01,10,11);
input s_262,s_263;//RE__ALLOW(00,01,10,11);
input s_264,s_265;//RE__ALLOW(00,01,10,11);
input s_266,s_267;//RE__ALLOW(00,01,10,11);
input s_268,s_269;//RE__ALLOW(00,01,10,11);
input s_270,s_271;//RE__ALLOW(00,01,10,11);
input s_272,s_273;//RE__ALLOW(00,01,10,11);
input s_274,s_275;//RE__ALLOW(00,01,10,11);
input s_276,s_277;//RE__ALLOW(00,01,10,11);
input s_278,s_279;//RE__ALLOW(00,01,10,11);
input s_280,s_281;//RE__ALLOW(00,01,10,11);
input s_282,s_283;//RE__ALLOW(00,01,10,11);
input s_284,s_285;//RE__ALLOW(00,01,10,11);
input s_286,s_287;//RE__ALLOW(00,01,10,11);
input s_288,s_289;//RE__ALLOW(00,01,10,11);
input s_290,s_291;//RE__ALLOW(00,01,10,11);
input s_292,s_293;//RE__ALLOW(00,01,10,11);
input s_294,s_295;//RE__ALLOW(00,01,10,11);
input s_296,s_297;//RE__ALLOW(00,01,10,11);
input s_298,s_299;//RE__ALLOW(00,01,10,11);
input s_300,s_301;//RE__ALLOW(00,01,10,11);
input s_302,s_303;//RE__ALLOW(00,01,10,11);
input s_304,s_305;//RE__ALLOW(00,01,10,11);
input s_306,s_307;//RE__ALLOW(00,01,10,11);
input s_308,s_309;//RE__ALLOW(00,01,10,11);
input s_310,s_311;//RE__ALLOW(00,01,10,11);
input s_312,s_313;//RE__ALLOW(00,01,10,11);
input s_314,s_315;//RE__ALLOW(00,01,10,11);
input s_316,s_317;//RE__ALLOW(00,01,10,11);
input s_318,s_319;//RE__ALLOW(00,01,10,11);
input s_320,s_321;//RE__ALLOW(00,01,10,11);
input s_322,s_323;//RE__ALLOW(00,01,10,11);
input s_324,s_325;//RE__ALLOW(00,01,10,11);
input s_326,s_327;//RE__ALLOW(00,01,10,11);
input s_328,s_329;//RE__ALLOW(00,01,10,11);
input s_330,s_331;//RE__ALLOW(00,01,10,11);
input s_332,s_333;//RE__ALLOW(00,01,10,11);
input s_334,s_335;//RE__ALLOW(00,01,10,11);
input s_336,s_337;//RE__ALLOW(00,01,10,11);
input s_338,s_339;//RE__ALLOW(00,01,10,11);
input s_340,s_341;//RE__ALLOW(00,01,10,11);
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;

  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate134inter0, gate134inter1, gate134inter2, gate134inter3, gate134inter4, gate134inter5, gate134inter6, gate134inter7, gate134inter8, gate134inter9, gate134inter10, gate134inter11, gate134inter12, gate453inter0, gate453inter1, gate453inter2, gate453inter3, gate453inter4, gate453inter5, gate453inter6, gate453inter7, gate453inter8, gate453inter9, gate453inter10, gate453inter11, gate453inter12, gate51inter0, gate51inter1, gate51inter2, gate51inter3, gate51inter4, gate51inter5, gate51inter6, gate51inter7, gate51inter8, gate51inter9, gate51inter10, gate51inter11, gate51inter12, gate66inter0, gate66inter1, gate66inter2, gate66inter3, gate66inter4, gate66inter5, gate66inter6, gate66inter7, gate66inter8, gate66inter9, gate66inter10, gate66inter11, gate66inter12, gate129inter0, gate129inter1, gate129inter2, gate129inter3, gate129inter4, gate129inter5, gate129inter6, gate129inter7, gate129inter8, gate129inter9, gate129inter10, gate129inter11, gate129inter12, gate491inter0, gate491inter1, gate491inter2, gate491inter3, gate491inter4, gate491inter5, gate491inter6, gate491inter7, gate491inter8, gate491inter9, gate491inter10, gate491inter11, gate491inter12, gate211inter0, gate211inter1, gate211inter2, gate211inter3, gate211inter4, gate211inter5, gate211inter6, gate211inter7, gate211inter8, gate211inter9, gate211inter10, gate211inter11, gate211inter12, gate175inter0, gate175inter1, gate175inter2, gate175inter3, gate175inter4, gate175inter5, gate175inter6, gate175inter7, gate175inter8, gate175inter9, gate175inter10, gate175inter11, gate175inter12, gate59inter0, gate59inter1, gate59inter2, gate59inter3, gate59inter4, gate59inter5, gate59inter6, gate59inter7, gate59inter8, gate59inter9, gate59inter10, gate59inter11, gate59inter12, gate502inter0, gate502inter1, gate502inter2, gate502inter3, gate502inter4, gate502inter5, gate502inter6, gate502inter7, gate502inter8, gate502inter9, gate502inter10, gate502inter11, gate502inter12, gate161inter0, gate161inter1, gate161inter2, gate161inter3, gate161inter4, gate161inter5, gate161inter6, gate161inter7, gate161inter8, gate161inter9, gate161inter10, gate161inter11, gate161inter12, gate275inter0, gate275inter1, gate275inter2, gate275inter3, gate275inter4, gate275inter5, gate275inter6, gate275inter7, gate275inter8, gate275inter9, gate275inter10, gate275inter11, gate275inter12, gate507inter0, gate507inter1, gate507inter2, gate507inter3, gate507inter4, gate507inter5, gate507inter6, gate507inter7, gate507inter8, gate507inter9, gate507inter10, gate507inter11, gate507inter12, gate168inter0, gate168inter1, gate168inter2, gate168inter3, gate168inter4, gate168inter5, gate168inter6, gate168inter7, gate168inter8, gate168inter9, gate168inter10, gate168inter11, gate168inter12, gate256inter0, gate256inter1, gate256inter2, gate256inter3, gate256inter4, gate256inter5, gate256inter6, gate256inter7, gate256inter8, gate256inter9, gate256inter10, gate256inter11, gate256inter12, gate396inter0, gate396inter1, gate396inter2, gate396inter3, gate396inter4, gate396inter5, gate396inter6, gate396inter7, gate396inter8, gate396inter9, gate396inter10, gate396inter11, gate396inter12, gate46inter0, gate46inter1, gate46inter2, gate46inter3, gate46inter4, gate46inter5, gate46inter6, gate46inter7, gate46inter8, gate46inter9, gate46inter10, gate46inter11, gate46inter12, gate292inter0, gate292inter1, gate292inter2, gate292inter3, gate292inter4, gate292inter5, gate292inter6, gate292inter7, gate292inter8, gate292inter9, gate292inter10, gate292inter11, gate292inter12, gate454inter0, gate454inter1, gate454inter2, gate454inter3, gate454inter4, gate454inter5, gate454inter6, gate454inter7, gate454inter8, gate454inter9, gate454inter10, gate454inter11, gate454inter12, gate249inter0, gate249inter1, gate249inter2, gate249inter3, gate249inter4, gate249inter5, gate249inter6, gate249inter7, gate249inter8, gate249inter9, gate249inter10, gate249inter11, gate249inter12, gate105inter0, gate105inter1, gate105inter2, gate105inter3, gate105inter4, gate105inter5, gate105inter6, gate105inter7, gate105inter8, gate105inter9, gate105inter10, gate105inter11, gate105inter12, gate447inter0, gate447inter1, gate447inter2, gate447inter3, gate447inter4, gate447inter5, gate447inter6, gate447inter7, gate447inter8, gate447inter9, gate447inter10, gate447inter11, gate447inter12, gate110inter0, gate110inter1, gate110inter2, gate110inter3, gate110inter4, gate110inter5, gate110inter6, gate110inter7, gate110inter8, gate110inter9, gate110inter10, gate110inter11, gate110inter12, gate235inter0, gate235inter1, gate235inter2, gate235inter3, gate235inter4, gate235inter5, gate235inter6, gate235inter7, gate235inter8, gate235inter9, gate235inter10, gate235inter11, gate235inter12, gate157inter0, gate157inter1, gate157inter2, gate157inter3, gate157inter4, gate157inter5, gate157inter6, gate157inter7, gate157inter8, gate157inter9, gate157inter10, gate157inter11, gate157inter12, gate180inter0, gate180inter1, gate180inter2, gate180inter3, gate180inter4, gate180inter5, gate180inter6, gate180inter7, gate180inter8, gate180inter9, gate180inter10, gate180inter11, gate180inter12, gate216inter0, gate216inter1, gate216inter2, gate216inter3, gate216inter4, gate216inter5, gate216inter6, gate216inter7, gate216inter8, gate216inter9, gate216inter10, gate216inter11, gate216inter12, gate483inter0, gate483inter1, gate483inter2, gate483inter3, gate483inter4, gate483inter5, gate483inter6, gate483inter7, gate483inter8, gate483inter9, gate483inter10, gate483inter11, gate483inter12, gate411inter0, gate411inter1, gate411inter2, gate411inter3, gate411inter4, gate411inter5, gate411inter6, gate411inter7, gate411inter8, gate411inter9, gate411inter10, gate411inter11, gate411inter12, gate248inter0, gate248inter1, gate248inter2, gate248inter3, gate248inter4, gate248inter5, gate248inter6, gate248inter7, gate248inter8, gate248inter9, gate248inter10, gate248inter11, gate248inter12, gate400inter0, gate400inter1, gate400inter2, gate400inter3, gate400inter4, gate400inter5, gate400inter6, gate400inter7, gate400inter8, gate400inter9, gate400inter10, gate400inter11, gate400inter12, gate63inter0, gate63inter1, gate63inter2, gate63inter3, gate63inter4, gate63inter5, gate63inter6, gate63inter7, gate63inter8, gate63inter9, gate63inter10, gate63inter11, gate63inter12, gate195inter0, gate195inter1, gate195inter2, gate195inter3, gate195inter4, gate195inter5, gate195inter6, gate195inter7, gate195inter8, gate195inter9, gate195inter10, gate195inter11, gate195inter12, gate153inter0, gate153inter1, gate153inter2, gate153inter3, gate153inter4, gate153inter5, gate153inter6, gate153inter7, gate153inter8, gate153inter9, gate153inter10, gate153inter11, gate153inter12, gate424inter0, gate424inter1, gate424inter2, gate424inter3, gate424inter4, gate424inter5, gate424inter6, gate424inter7, gate424inter8, gate424inter9, gate424inter10, gate424inter11, gate424inter12, gate77inter0, gate77inter1, gate77inter2, gate77inter3, gate77inter4, gate77inter5, gate77inter6, gate77inter7, gate77inter8, gate77inter9, gate77inter10, gate77inter11, gate77inter12, gate403inter0, gate403inter1, gate403inter2, gate403inter3, gate403inter4, gate403inter5, gate403inter6, gate403inter7, gate403inter8, gate403inter9, gate403inter10, gate403inter11, gate403inter12, gate250inter0, gate250inter1, gate250inter2, gate250inter3, gate250inter4, gate250inter5, gate250inter6, gate250inter7, gate250inter8, gate250inter9, gate250inter10, gate250inter11, gate250inter12, gate43inter0, gate43inter1, gate43inter2, gate43inter3, gate43inter4, gate43inter5, gate43inter6, gate43inter7, gate43inter8, gate43inter9, gate43inter10, gate43inter11, gate43inter12, gate271inter0, gate271inter1, gate271inter2, gate271inter3, gate271inter4, gate271inter5, gate271inter6, gate271inter7, gate271inter8, gate271inter9, gate271inter10, gate271inter11, gate271inter12, gate142inter0, gate142inter1, gate142inter2, gate142inter3, gate142inter4, gate142inter5, gate142inter6, gate142inter7, gate142inter8, gate142inter9, gate142inter10, gate142inter11, gate142inter12, gate64inter0, gate64inter1, gate64inter2, gate64inter3, gate64inter4, gate64inter5, gate64inter6, gate64inter7, gate64inter8, gate64inter9, gate64inter10, gate64inter11, gate64inter12, gate241inter0, gate241inter1, gate241inter2, gate241inter3, gate241inter4, gate241inter5, gate241inter6, gate241inter7, gate241inter8, gate241inter9, gate241inter10, gate241inter11, gate241inter12, gate442inter0, gate442inter1, gate442inter2, gate442inter3, gate442inter4, gate442inter5, gate442inter6, gate442inter7, gate442inter8, gate442inter9, gate442inter10, gate442inter11, gate442inter12, gate429inter0, gate429inter1, gate429inter2, gate429inter3, gate429inter4, gate429inter5, gate429inter6, gate429inter7, gate429inter8, gate429inter9, gate429inter10, gate429inter11, gate429inter12, gate408inter0, gate408inter1, gate408inter2, gate408inter3, gate408inter4, gate408inter5, gate408inter6, gate408inter7, gate408inter8, gate408inter9, gate408inter10, gate408inter11, gate408inter12, gate207inter0, gate207inter1, gate207inter2, gate207inter3, gate207inter4, gate207inter5, gate207inter6, gate207inter7, gate207inter8, gate207inter9, gate207inter10, gate207inter11, gate207inter12, gate407inter0, gate407inter1, gate407inter2, gate407inter3, gate407inter4, gate407inter5, gate407inter6, gate407inter7, gate407inter8, gate407inter9, gate407inter10, gate407inter11, gate407inter12, gate277inter0, gate277inter1, gate277inter2, gate277inter3, gate277inter4, gate277inter5, gate277inter6, gate277inter7, gate277inter8, gate277inter9, gate277inter10, gate277inter11, gate277inter12, gate81inter0, gate81inter1, gate81inter2, gate81inter3, gate81inter4, gate81inter5, gate81inter6, gate81inter7, gate81inter8, gate81inter9, gate81inter10, gate81inter11, gate81inter12, gate30inter0, gate30inter1, gate30inter2, gate30inter3, gate30inter4, gate30inter5, gate30inter6, gate30inter7, gate30inter8, gate30inter9, gate30inter10, gate30inter11, gate30inter12, gate481inter0, gate481inter1, gate481inter2, gate481inter3, gate481inter4, gate481inter5, gate481inter6, gate481inter7, gate481inter8, gate481inter9, gate481inter10, gate481inter11, gate481inter12, gate192inter0, gate192inter1, gate192inter2, gate192inter3, gate192inter4, gate192inter5, gate192inter6, gate192inter7, gate192inter8, gate192inter9, gate192inter10, gate192inter11, gate192inter12, gate280inter0, gate280inter1, gate280inter2, gate280inter3, gate280inter4, gate280inter5, gate280inter6, gate280inter7, gate280inter8, gate280inter9, gate280inter10, gate280inter11, gate280inter12, gate47inter0, gate47inter1, gate47inter2, gate47inter3, gate47inter4, gate47inter5, gate47inter6, gate47inter7, gate47inter8, gate47inter9, gate47inter10, gate47inter11, gate47inter12, gate84inter0, gate84inter1, gate84inter2, gate84inter3, gate84inter4, gate84inter5, gate84inter6, gate84inter7, gate84inter8, gate84inter9, gate84inter10, gate84inter11, gate84inter12, gate226inter0, gate226inter1, gate226inter2, gate226inter3, gate226inter4, gate226inter5, gate226inter6, gate226inter7, gate226inter8, gate226inter9, gate226inter10, gate226inter11, gate226inter12, gate261inter0, gate261inter1, gate261inter2, gate261inter3, gate261inter4, gate261inter5, gate261inter6, gate261inter7, gate261inter8, gate261inter9, gate261inter10, gate261inter11, gate261inter12, gate291inter0, gate291inter1, gate291inter2, gate291inter3, gate291inter4, gate291inter5, gate291inter6, gate291inter7, gate291inter8, gate291inter9, gate291inter10, gate291inter11, gate291inter12, gate49inter0, gate49inter1, gate49inter2, gate49inter3, gate49inter4, gate49inter5, gate49inter6, gate49inter7, gate49inter8, gate49inter9, gate49inter10, gate49inter11, gate49inter12, gate149inter0, gate149inter1, gate149inter2, gate149inter3, gate149inter4, gate149inter5, gate149inter6, gate149inter7, gate149inter8, gate149inter9, gate149inter10, gate149inter11, gate149inter12, gate20inter0, gate20inter1, gate20inter2, gate20inter3, gate20inter4, gate20inter5, gate20inter6, gate20inter7, gate20inter8, gate20inter9, gate20inter10, gate20inter11, gate20inter12, gate166inter0, gate166inter1, gate166inter2, gate166inter3, gate166inter4, gate166inter5, gate166inter6, gate166inter7, gate166inter8, gate166inter9, gate166inter10, gate166inter11, gate166inter12, gate270inter0, gate270inter1, gate270inter2, gate270inter3, gate270inter4, gate270inter5, gate270inter6, gate270inter7, gate270inter8, gate270inter9, gate270inter10, gate270inter11, gate270inter12, gate100inter0, gate100inter1, gate100inter2, gate100inter3, gate100inter4, gate100inter5, gate100inter6, gate100inter7, gate100inter8, gate100inter9, gate100inter10, gate100inter11, gate100inter12, gate266inter0, gate266inter1, gate266inter2, gate266inter3, gate266inter4, gate266inter5, gate266inter6, gate266inter7, gate266inter8, gate266inter9, gate266inter10, gate266inter11, gate266inter12, gate398inter0, gate398inter1, gate398inter2, gate398inter3, gate398inter4, gate398inter5, gate398inter6, gate398inter7, gate398inter8, gate398inter9, gate398inter10, gate398inter11, gate398inter12, gate120inter0, gate120inter1, gate120inter2, gate120inter3, gate120inter4, gate120inter5, gate120inter6, gate120inter7, gate120inter8, gate120inter9, gate120inter10, gate120inter11, gate120inter12, gate255inter0, gate255inter1, gate255inter2, gate255inter3, gate255inter4, gate255inter5, gate255inter6, gate255inter7, gate255inter8, gate255inter9, gate255inter10, gate255inter11, gate255inter12, gate487inter0, gate487inter1, gate487inter2, gate487inter3, gate487inter4, gate487inter5, gate487inter6, gate487inter7, gate487inter8, gate487inter9, gate487inter10, gate487inter11, gate487inter12, gate234inter0, gate234inter1, gate234inter2, gate234inter3, gate234inter4, gate234inter5, gate234inter6, gate234inter7, gate234inter8, gate234inter9, gate234inter10, gate234inter11, gate234inter12, gate111inter0, gate111inter1, gate111inter2, gate111inter3, gate111inter4, gate111inter5, gate111inter6, gate111inter7, gate111inter8, gate111inter9, gate111inter10, gate111inter11, gate111inter12, gate71inter0, gate71inter1, gate71inter2, gate71inter3, gate71inter4, gate71inter5, gate71inter6, gate71inter7, gate71inter8, gate71inter9, gate71inter10, gate71inter11, gate71inter12, gate267inter0, gate267inter1, gate267inter2, gate267inter3, gate267inter4, gate267inter5, gate267inter6, gate267inter7, gate267inter8, gate267inter9, gate267inter10, gate267inter11, gate267inter12, gate215inter0, gate215inter1, gate215inter2, gate215inter3, gate215inter4, gate215inter5, gate215inter6, gate215inter7, gate215inter8, gate215inter9, gate215inter10, gate215inter11, gate215inter12, gate511inter0, gate511inter1, gate511inter2, gate511inter3, gate511inter4, gate511inter5, gate511inter6, gate511inter7, gate511inter8, gate511inter9, gate511inter10, gate511inter11, gate511inter12, gate224inter0, gate224inter1, gate224inter2, gate224inter3, gate224inter4, gate224inter5, gate224inter6, gate224inter7, gate224inter8, gate224inter9, gate224inter10, gate224inter11, gate224inter12, gate184inter0, gate184inter1, gate184inter2, gate184inter3, gate184inter4, gate184inter5, gate184inter6, gate184inter7, gate184inter8, gate184inter9, gate184inter10, gate184inter11, gate184inter12, gate197inter0, gate197inter1, gate197inter2, gate197inter3, gate197inter4, gate197inter5, gate197inter6, gate197inter7, gate197inter8, gate197inter9, gate197inter10, gate197inter11, gate197inter12, gate148inter0, gate148inter1, gate148inter2, gate148inter3, gate148inter4, gate148inter5, gate148inter6, gate148inter7, gate148inter8, gate148inter9, gate148inter10, gate148inter11, gate148inter12, gate264inter0, gate264inter1, gate264inter2, gate264inter3, gate264inter4, gate264inter5, gate264inter6, gate264inter7, gate264inter8, gate264inter9, gate264inter10, gate264inter11, gate264inter12, gate274inter0, gate274inter1, gate274inter2, gate274inter3, gate274inter4, gate274inter5, gate274inter6, gate274inter7, gate274inter8, gate274inter9, gate274inter10, gate274inter11, gate274inter12, gate206inter0, gate206inter1, gate206inter2, gate206inter3, gate206inter4, gate206inter5, gate206inter6, gate206inter7, gate206inter8, gate206inter9, gate206inter10, gate206inter11, gate206inter12, gate21inter0, gate21inter1, gate21inter2, gate21inter3, gate21inter4, gate21inter5, gate21inter6, gate21inter7, gate21inter8, gate21inter9, gate21inter10, gate21inter11, gate21inter12, gate160inter0, gate160inter1, gate160inter2, gate160inter3, gate160inter4, gate160inter5, gate160inter6, gate160inter7, gate160inter8, gate160inter9, gate160inter10, gate160inter11, gate160inter12, gate397inter0, gate397inter1, gate397inter2, gate397inter3, gate397inter4, gate397inter5, gate397inter6, gate397inter7, gate397inter8, gate397inter9, gate397inter10, gate397inter11, gate397inter12, gate56inter0, gate56inter1, gate56inter2, gate56inter3, gate56inter4, gate56inter5, gate56inter6, gate56inter7, gate56inter8, gate56inter9, gate56inter10, gate56inter11, gate56inter12, gate477inter0, gate477inter1, gate477inter2, gate477inter3, gate477inter4, gate477inter5, gate477inter6, gate477inter7, gate477inter8, gate477inter9, gate477inter10, gate477inter11, gate477inter12, gate174inter0, gate174inter1, gate174inter2, gate174inter3, gate174inter4, gate174inter5, gate174inter6, gate174inter7, gate174inter8, gate174inter9, gate174inter10, gate174inter11, gate174inter12, gate75inter0, gate75inter1, gate75inter2, gate75inter3, gate75inter4, gate75inter5, gate75inter6, gate75inter7, gate75inter8, gate75inter9, gate75inter10, gate75inter11, gate75inter12, gate269inter0, gate269inter1, gate269inter2, gate269inter3, gate269inter4, gate269inter5, gate269inter6, gate269inter7, gate269inter8, gate269inter9, gate269inter10, gate269inter11, gate269inter12, gate413inter0, gate413inter1, gate413inter2, gate413inter3, gate413inter4, gate413inter5, gate413inter6, gate413inter7, gate413inter8, gate413inter9, gate413inter10, gate413inter11, gate413inter12, gate121inter0, gate121inter1, gate121inter2, gate121inter3, gate121inter4, gate121inter5, gate121inter6, gate121inter7, gate121inter8, gate121inter9, gate121inter10, gate121inter11, gate121inter12, gate479inter0, gate479inter1, gate479inter2, gate479inter3, gate479inter4, gate479inter5, gate479inter6, gate479inter7, gate479inter8, gate479inter9, gate479inter10, gate479inter11, gate479inter12, gate97inter0, gate97inter1, gate97inter2, gate97inter3, gate97inter4, gate97inter5, gate97inter6, gate97inter7, gate97inter8, gate97inter9, gate97inter10, gate97inter11, gate97inter12, gate452inter0, gate452inter1, gate452inter2, gate452inter3, gate452inter4, gate452inter5, gate452inter6, gate452inter7, gate452inter8, gate452inter9, gate452inter10, gate452inter11, gate452inter12, gate193inter0, gate193inter1, gate193inter2, gate193inter3, gate193inter4, gate193inter5, gate193inter6, gate193inter7, gate193inter8, gate193inter9, gate193inter10, gate193inter11, gate193inter12, gate132inter0, gate132inter1, gate132inter2, gate132inter3, gate132inter4, gate132inter5, gate132inter6, gate132inter7, gate132inter8, gate132inter9, gate132inter10, gate132inter11, gate132inter12, gate123inter0, gate123inter1, gate123inter2, gate123inter3, gate123inter4, gate123inter5, gate123inter6, gate123inter7, gate123inter8, gate123inter9, gate123inter10, gate123inter11, gate123inter12, gate495inter0, gate495inter1, gate495inter2, gate495inter3, gate495inter4, gate495inter5, gate495inter6, gate495inter7, gate495inter8, gate495inter9, gate495inter10, gate495inter11, gate495inter12, gate493inter0, gate493inter1, gate493inter2, gate493inter3, gate493inter4, gate493inter5, gate493inter6, gate493inter7, gate493inter8, gate493inter9, gate493inter10, gate493inter11, gate493inter12, gate69inter0, gate69inter1, gate69inter2, gate69inter3, gate69inter4, gate69inter5, gate69inter6, gate69inter7, gate69inter8, gate69inter9, gate69inter10, gate69inter11, gate69inter12, gate484inter0, gate484inter1, gate484inter2, gate484inter3, gate484inter4, gate484inter5, gate484inter6, gate484inter7, gate484inter8, gate484inter9, gate484inter10, gate484inter11, gate484inter12, gate422inter0, gate422inter1, gate422inter2, gate422inter3, gate422inter4, gate422inter5, gate422inter6, gate422inter7, gate422inter8, gate422inter9, gate422inter10, gate422inter11, gate422inter12, gate401inter0, gate401inter1, gate401inter2, gate401inter3, gate401inter4, gate401inter5, gate401inter6, gate401inter7, gate401inter8, gate401inter9, gate401inter10, gate401inter11, gate401inter12, gate44inter0, gate44inter1, gate44inter2, gate44inter3, gate44inter4, gate44inter5, gate44inter6, gate44inter7, gate44inter8, gate44inter9, gate44inter10, gate44inter11, gate44inter12, gate252inter0, gate252inter1, gate252inter2, gate252inter3, gate252inter4, gate252inter5, gate252inter6, gate252inter7, gate252inter8, gate252inter9, gate252inter10, gate252inter11, gate252inter12, gate428inter0, gate428inter1, gate428inter2, gate428inter3, gate428inter4, gate428inter5, gate428inter6, gate428inter7, gate428inter8, gate428inter9, gate428inter10, gate428inter11, gate428inter12, gate205inter0, gate205inter1, gate205inter2, gate205inter3, gate205inter4, gate205inter5, gate205inter6, gate205inter7, gate205inter8, gate205inter9, gate205inter10, gate205inter11, gate205inter12, gate164inter0, gate164inter1, gate164inter2, gate164inter3, gate164inter4, gate164inter5, gate164inter6, gate164inter7, gate164inter8, gate164inter9, gate164inter10, gate164inter11, gate164inter12, gate467inter0, gate467inter1, gate467inter2, gate467inter3, gate467inter4, gate467inter5, gate467inter6, gate467inter7, gate467inter8, gate467inter9, gate467inter10, gate467inter11, gate467inter12, gate217inter0, gate217inter1, gate217inter2, gate217inter3, gate217inter4, gate217inter5, gate217inter6, gate217inter7, gate217inter8, gate217inter9, gate217inter10, gate217inter11, gate217inter12, gate470inter0, gate470inter1, gate470inter2, gate470inter3, gate470inter4, gate470inter5, gate470inter6, gate470inter7, gate470inter8, gate470inter9, gate470inter10, gate470inter11, gate470inter12, gate202inter0, gate202inter1, gate202inter2, gate202inter3, gate202inter4, gate202inter5, gate202inter6, gate202inter7, gate202inter8, gate202inter9, gate202inter10, gate202inter11, gate202inter12, gate73inter0, gate73inter1, gate73inter2, gate73inter3, gate73inter4, gate73inter5, gate73inter6, gate73inter7, gate73inter8, gate73inter9, gate73inter10, gate73inter11, gate73inter12, gate116inter0, gate116inter1, gate116inter2, gate116inter3, gate116inter4, gate116inter5, gate116inter6, gate116inter7, gate116inter8, gate116inter9, gate116inter10, gate116inter11, gate116inter12, gate420inter0, gate420inter1, gate420inter2, gate420inter3, gate420inter4, gate420inter5, gate420inter6, gate420inter7, gate420inter8, gate420inter9, gate420inter10, gate420inter11, gate420inter12, gate170inter0, gate170inter1, gate170inter2, gate170inter3, gate170inter4, gate170inter5, gate170inter6, gate170inter7, gate170inter8, gate170inter9, gate170inter10, gate170inter11, gate170inter12, gate11inter0, gate11inter1, gate11inter2, gate11inter3, gate11inter4, gate11inter5, gate11inter6, gate11inter7, gate11inter8, gate11inter9, gate11inter10, gate11inter11, gate11inter12, gate40inter0, gate40inter1, gate40inter2, gate40inter3, gate40inter4, gate40inter5, gate40inter6, gate40inter7, gate40inter8, gate40inter9, gate40inter10, gate40inter11, gate40inter12, gate55inter0, gate55inter1, gate55inter2, gate55inter3, gate55inter4, gate55inter5, gate55inter6, gate55inter7, gate55inter8, gate55inter9, gate55inter10, gate55inter11, gate55inter12, gate93inter0, gate93inter1, gate93inter2, gate93inter3, gate93inter4, gate93inter5, gate93inter6, gate93inter7, gate93inter8, gate93inter9, gate93inter10, gate93inter11, gate93inter12, gate239inter0, gate239inter1, gate239inter2, gate239inter3, gate239inter4, gate239inter5, gate239inter6, gate239inter7, gate239inter8, gate239inter9, gate239inter10, gate239inter11, gate239inter12, gate212inter0, gate212inter1, gate212inter2, gate212inter3, gate212inter4, gate212inter5, gate212inter6, gate212inter7, gate212inter8, gate212inter9, gate212inter10, gate212inter11, gate212inter12, gate115inter0, gate115inter1, gate115inter2, gate115inter3, gate115inter4, gate115inter5, gate115inter6, gate115inter7, gate115inter8, gate115inter9, gate115inter10, gate115inter11, gate115inter12, gate141inter0, gate141inter1, gate141inter2, gate141inter3, gate141inter4, gate141inter5, gate141inter6, gate141inter7, gate141inter8, gate141inter9, gate141inter10, gate141inter11, gate141inter12, gate287inter0, gate287inter1, gate287inter2, gate287inter3, gate287inter4, gate287inter5, gate287inter6, gate287inter7, gate287inter8, gate287inter9, gate287inter10, gate287inter11, gate287inter12, gate86inter0, gate86inter1, gate86inter2, gate86inter3, gate86inter4, gate86inter5, gate86inter6, gate86inter7, gate86inter8, gate86inter9, gate86inter10, gate86inter11, gate86inter12, gate406inter0, gate406inter1, gate406inter2, gate406inter3, gate406inter4, gate406inter5, gate406inter6, gate406inter7, gate406inter8, gate406inter9, gate406inter10, gate406inter11, gate406inter12, gate434inter0, gate434inter1, gate434inter2, gate434inter3, gate434inter4, gate434inter5, gate434inter6, gate434inter7, gate434inter8, gate434inter9, gate434inter10, gate434inter11, gate434inter12, gate421inter0, gate421inter1, gate421inter2, gate421inter3, gate421inter4, gate421inter5, gate421inter6, gate421inter7, gate421inter8, gate421inter9, gate421inter10, gate421inter11, gate421inter12, gate19inter0, gate19inter1, gate19inter2, gate19inter3, gate19inter4, gate19inter5, gate19inter6, gate19inter7, gate19inter8, gate19inter9, gate19inter10, gate19inter11, gate19inter12, gate150inter0, gate150inter1, gate150inter2, gate150inter3, gate150inter4, gate150inter5, gate150inter6, gate150inter7, gate150inter8, gate150inter9, gate150inter10, gate150inter11, gate150inter12, gate191inter0, gate191inter1, gate191inter2, gate191inter3, gate191inter4, gate191inter5, gate191inter6, gate191inter7, gate191inter8, gate191inter9, gate191inter10, gate191inter11, gate191inter12, gate210inter0, gate210inter1, gate210inter2, gate210inter3, gate210inter4, gate210inter5, gate210inter6, gate210inter7, gate210inter8, gate210inter9, gate210inter10, gate210inter11, gate210inter12, gate485inter0, gate485inter1, gate485inter2, gate485inter3, gate485inter4, gate485inter5, gate485inter6, gate485inter7, gate485inter8, gate485inter9, gate485inter10, gate485inter11, gate485inter12, gate276inter0, gate276inter1, gate276inter2, gate276inter3, gate276inter4, gate276inter5, gate276inter6, gate276inter7, gate276inter8, gate276inter9, gate276inter10, gate276inter11, gate276inter12, gate506inter0, gate506inter1, gate506inter2, gate506inter3, gate506inter4, gate506inter5, gate506inter6, gate506inter7, gate506inter8, gate506inter9, gate506inter10, gate506inter11, gate506inter12, gate16inter0, gate16inter1, gate16inter2, gate16inter3, gate16inter4, gate16inter5, gate16inter6, gate16inter7, gate16inter8, gate16inter9, gate16inter10, gate16inter11, gate16inter12, gate448inter0, gate448inter1, gate448inter2, gate448inter3, gate448inter4, gate448inter5, gate448inter6, gate448inter7, gate448inter8, gate448inter9, gate448inter10, gate448inter11, gate448inter12, gate208inter0, gate208inter1, gate208inter2, gate208inter3, gate208inter4, gate208inter5, gate208inter6, gate208inter7, gate208inter8, gate208inter9, gate208inter10, gate208inter11, gate208inter12, gate113inter0, gate113inter1, gate113inter2, gate113inter3, gate113inter4, gate113inter5, gate113inter6, gate113inter7, gate113inter8, gate113inter9, gate113inter10, gate113inter11, gate113inter12, gate62inter0, gate62inter1, gate62inter2, gate62inter3, gate62inter4, gate62inter5, gate62inter6, gate62inter7, gate62inter8, gate62inter9, gate62inter10, gate62inter11, gate62inter12, gate72inter0, gate72inter1, gate72inter2, gate72inter3, gate72inter4, gate72inter5, gate72inter6, gate72inter7, gate72inter8, gate72inter9, gate72inter10, gate72inter11, gate72inter12, gate200inter0, gate200inter1, gate200inter2, gate200inter3, gate200inter4, gate200inter5, gate200inter6, gate200inter7, gate200inter8, gate200inter9, gate200inter10, gate200inter11, gate200inter12, gate469inter0, gate469inter1, gate469inter2, gate469inter3, gate469inter4, gate469inter5, gate469inter6, gate469inter7, gate469inter8, gate469inter9, gate469inter10, gate469inter11, gate469inter12, gate433inter0, gate433inter1, gate433inter2, gate433inter3, gate433inter4, gate433inter5, gate433inter6, gate433inter7, gate433inter8, gate433inter9, gate433inter10, gate433inter11, gate433inter12, gate92inter0, gate92inter1, gate92inter2, gate92inter3, gate92inter4, gate92inter5, gate92inter6, gate92inter7, gate92inter8, gate92inter9, gate92inter10, gate92inter11, gate92inter12, gate294inter0, gate294inter1, gate294inter2, gate294inter3, gate294inter4, gate294inter5, gate294inter6, gate294inter7, gate294inter8, gate294inter9, gate294inter10, gate294inter11, gate294inter12, gate50inter0, gate50inter1, gate50inter2, gate50inter3, gate50inter4, gate50inter5, gate50inter6, gate50inter7, gate50inter8, gate50inter9, gate50inter10, gate50inter11, gate50inter12, gate173inter0, gate173inter1, gate173inter2, gate173inter3, gate173inter4, gate173inter5, gate173inter6, gate173inter7, gate173inter8, gate173inter9, gate173inter10, gate173inter11, gate173inter12, gate169inter0, gate169inter1, gate169inter2, gate169inter3, gate169inter4, gate169inter5, gate169inter6, gate169inter7, gate169inter8, gate169inter9, gate169inter10, gate169inter11, gate169inter12, gate103inter0, gate103inter1, gate103inter2, gate103inter3, gate103inter4, gate103inter5, gate103inter6, gate103inter7, gate103inter8, gate103inter9, gate103inter10, gate103inter11, gate103inter12, gate133inter0, gate133inter1, gate133inter2, gate133inter3, gate133inter4, gate133inter5, gate133inter6, gate133inter7, gate133inter8, gate133inter9, gate133inter10, gate133inter11, gate133inter12, gate98inter0, gate98inter1, gate98inter2, gate98inter3, gate98inter4, gate98inter5, gate98inter6, gate98inter7, gate98inter8, gate98inter9, gate98inter10, gate98inter11, gate98inter12, gate293inter0, gate293inter1, gate293inter2, gate293inter3, gate293inter4, gate293inter5, gate293inter6, gate293inter7, gate293inter8, gate293inter9, gate293inter10, gate293inter11, gate293inter12, gate279inter0, gate279inter1, gate279inter2, gate279inter3, gate279inter4, gate279inter5, gate279inter6, gate279inter7, gate279inter8, gate279inter9, gate279inter10, gate279inter11, gate279inter12, gate23inter0, gate23inter1, gate23inter2, gate23inter3, gate23inter4, gate23inter5, gate23inter6, gate23inter7, gate23inter8, gate23inter9, gate23inter10, gate23inter11, gate23inter12, gate244inter0, gate244inter1, gate244inter2, gate244inter3, gate244inter4, gate244inter5, gate244inter6, gate244inter7, gate244inter8, gate244inter9, gate244inter10, gate244inter11, gate244inter12, gate171inter0, gate171inter1, gate171inter2, gate171inter3, gate171inter4, gate171inter5, gate171inter6, gate171inter7, gate171inter8, gate171inter9, gate171inter10, gate171inter11, gate171inter12, gate449inter0, gate449inter1, gate449inter2, gate449inter3, gate449inter4, gate449inter5, gate449inter6, gate449inter7, gate449inter8, gate449inter9, gate449inter10, gate449inter11, gate449inter12, gate38inter0, gate38inter1, gate38inter2, gate38inter3, gate38inter4, gate38inter5, gate38inter6, gate38inter7, gate38inter8, gate38inter9, gate38inter10, gate38inter11, gate38inter12, gate91inter0, gate91inter1, gate91inter2, gate91inter3, gate91inter4, gate91inter5, gate91inter6, gate91inter7, gate91inter8, gate91inter9, gate91inter10, gate91inter11, gate91inter12, gate96inter0, gate96inter1, gate96inter2, gate96inter3, gate96inter4, gate96inter5, gate96inter6, gate96inter7, gate96inter8, gate96inter9, gate96inter10, gate96inter11, gate96inter12, gate17inter0, gate17inter1, gate17inter2, gate17inter3, gate17inter4, gate17inter5, gate17inter6, gate17inter7, gate17inter8, gate17inter9, gate17inter10, gate17inter11, gate17inter12, gate482inter0, gate482inter1, gate482inter2, gate482inter3, gate482inter4, gate482inter5, gate482inter6, gate482inter7, gate482inter8, gate482inter9, gate482inter10, gate482inter11, gate482inter12, gate444inter0, gate444inter1, gate444inter2, gate444inter3, gate444inter4, gate444inter5, gate444inter6, gate444inter7, gate444inter8, gate444inter9, gate444inter10, gate444inter11, gate444inter12, gate106inter0, gate106inter1, gate106inter2, gate106inter3, gate106inter4, gate106inter5, gate106inter6, gate106inter7, gate106inter8, gate106inter9, gate106inter10, gate106inter11, gate106inter12, gate414inter0, gate414inter1, gate414inter2, gate414inter3, gate414inter4, gate414inter5, gate414inter6, gate414inter7, gate414inter8, gate414inter9, gate414inter10, gate414inter11, gate414inter12, gate296inter0, gate296inter1, gate296inter2, gate296inter3, gate296inter4, gate296inter5, gate296inter6, gate296inter7, gate296inter8, gate296inter9, gate296inter10, gate296inter11, gate296inter12, gate29inter0, gate29inter1, gate29inter2, gate29inter3, gate29inter4, gate29inter5, gate29inter6, gate29inter7, gate29inter8, gate29inter9, gate29inter10, gate29inter11, gate29inter12;



and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );
nand2 gate9( .a(G1), .b(G2), .O(G266) );
nand2 gate10( .a(G3), .b(G4), .O(G269) );

  xor2  gate2199(.a(G6), .b(G5), .O(gate11inter0));
  nand2 gate2200(.a(gate11inter0), .b(s_236), .O(gate11inter1));
  and2  gate2201(.a(G6), .b(G5), .O(gate11inter2));
  inv1  gate2202(.a(s_236), .O(gate11inter3));
  inv1  gate2203(.a(s_237), .O(gate11inter4));
  nand2 gate2204(.a(gate11inter4), .b(gate11inter3), .O(gate11inter5));
  nor2  gate2205(.a(gate11inter5), .b(gate11inter2), .O(gate11inter6));
  inv1  gate2206(.a(G5), .O(gate11inter7));
  inv1  gate2207(.a(G6), .O(gate11inter8));
  nand2 gate2208(.a(gate11inter8), .b(gate11inter7), .O(gate11inter9));
  nand2 gate2209(.a(s_237), .b(gate11inter3), .O(gate11inter10));
  nor2  gate2210(.a(gate11inter10), .b(gate11inter9), .O(gate11inter11));
  nor2  gate2211(.a(gate11inter11), .b(gate11inter6), .O(gate11inter12));
  nand2 gate2212(.a(gate11inter12), .b(gate11inter1), .O(G272));
nand2 gate12( .a(G7), .b(G8), .O(G275) );
nand2 gate13( .a(G9), .b(G10), .O(G278) );
nand2 gate14( .a(G11), .b(G12), .O(G281) );
nand2 gate15( .a(G13), .b(G14), .O(G284) );

  xor2  gate2479(.a(G16), .b(G15), .O(gate16inter0));
  nand2 gate2480(.a(gate16inter0), .b(s_276), .O(gate16inter1));
  and2  gate2481(.a(G16), .b(G15), .O(gate16inter2));
  inv1  gate2482(.a(s_276), .O(gate16inter3));
  inv1  gate2483(.a(s_277), .O(gate16inter4));
  nand2 gate2484(.a(gate16inter4), .b(gate16inter3), .O(gate16inter5));
  nor2  gate2485(.a(gate16inter5), .b(gate16inter2), .O(gate16inter6));
  inv1  gate2486(.a(G15), .O(gate16inter7));
  inv1  gate2487(.a(G16), .O(gate16inter8));
  nand2 gate2488(.a(gate16inter8), .b(gate16inter7), .O(gate16inter9));
  nand2 gate2489(.a(s_277), .b(gate16inter3), .O(gate16inter10));
  nor2  gate2490(.a(gate16inter10), .b(gate16inter9), .O(gate16inter11));
  nor2  gate2491(.a(gate16inter11), .b(gate16inter6), .O(gate16inter12));
  nand2 gate2492(.a(gate16inter12), .b(gate16inter1), .O(G287));

  xor2  gate2843(.a(G18), .b(G17), .O(gate17inter0));
  nand2 gate2844(.a(gate17inter0), .b(s_328), .O(gate17inter1));
  and2  gate2845(.a(G18), .b(G17), .O(gate17inter2));
  inv1  gate2846(.a(s_328), .O(gate17inter3));
  inv1  gate2847(.a(s_329), .O(gate17inter4));
  nand2 gate2848(.a(gate17inter4), .b(gate17inter3), .O(gate17inter5));
  nor2  gate2849(.a(gate17inter5), .b(gate17inter2), .O(gate17inter6));
  inv1  gate2850(.a(G17), .O(gate17inter7));
  inv1  gate2851(.a(G18), .O(gate17inter8));
  nand2 gate2852(.a(gate17inter8), .b(gate17inter7), .O(gate17inter9));
  nand2 gate2853(.a(s_329), .b(gate17inter3), .O(gate17inter10));
  nor2  gate2854(.a(gate17inter10), .b(gate17inter9), .O(gate17inter11));
  nor2  gate2855(.a(gate17inter11), .b(gate17inter6), .O(gate17inter12));
  nand2 gate2856(.a(gate17inter12), .b(gate17inter1), .O(G290));
nand2 gate18( .a(G19), .b(G20), .O(G293) );

  xor2  gate2381(.a(G22), .b(G21), .O(gate19inter0));
  nand2 gate2382(.a(gate19inter0), .b(s_262), .O(gate19inter1));
  and2  gate2383(.a(G22), .b(G21), .O(gate19inter2));
  inv1  gate2384(.a(s_262), .O(gate19inter3));
  inv1  gate2385(.a(s_263), .O(gate19inter4));
  nand2 gate2386(.a(gate19inter4), .b(gate19inter3), .O(gate19inter5));
  nor2  gate2387(.a(gate19inter5), .b(gate19inter2), .O(gate19inter6));
  inv1  gate2388(.a(G21), .O(gate19inter7));
  inv1  gate2389(.a(G22), .O(gate19inter8));
  nand2 gate2390(.a(gate19inter8), .b(gate19inter7), .O(gate19inter9));
  nand2 gate2391(.a(s_263), .b(gate19inter3), .O(gate19inter10));
  nor2  gate2392(.a(gate19inter10), .b(gate19inter9), .O(gate19inter11));
  nor2  gate2393(.a(gate19inter11), .b(gate19inter6), .O(gate19inter12));
  nand2 gate2394(.a(gate19inter12), .b(gate19inter1), .O(G296));

  xor2  gate1401(.a(G24), .b(G23), .O(gate20inter0));
  nand2 gate1402(.a(gate20inter0), .b(s_122), .O(gate20inter1));
  and2  gate1403(.a(G24), .b(G23), .O(gate20inter2));
  inv1  gate1404(.a(s_122), .O(gate20inter3));
  inv1  gate1405(.a(s_123), .O(gate20inter4));
  nand2 gate1406(.a(gate20inter4), .b(gate20inter3), .O(gate20inter5));
  nor2  gate1407(.a(gate20inter5), .b(gate20inter2), .O(gate20inter6));
  inv1  gate1408(.a(G23), .O(gate20inter7));
  inv1  gate1409(.a(G24), .O(gate20inter8));
  nand2 gate1410(.a(gate20inter8), .b(gate20inter7), .O(gate20inter9));
  nand2 gate1411(.a(s_123), .b(gate20inter3), .O(gate20inter10));
  nor2  gate1412(.a(gate20inter10), .b(gate20inter9), .O(gate20inter11));
  nor2  gate1413(.a(gate20inter11), .b(gate20inter6), .O(gate20inter12));
  nand2 gate1414(.a(gate20inter12), .b(gate20inter1), .O(G299));

  xor2  gate1709(.a(G26), .b(G25), .O(gate21inter0));
  nand2 gate1710(.a(gate21inter0), .b(s_166), .O(gate21inter1));
  and2  gate1711(.a(G26), .b(G25), .O(gate21inter2));
  inv1  gate1712(.a(s_166), .O(gate21inter3));
  inv1  gate1713(.a(s_167), .O(gate21inter4));
  nand2 gate1714(.a(gate21inter4), .b(gate21inter3), .O(gate21inter5));
  nor2  gate1715(.a(gate21inter5), .b(gate21inter2), .O(gate21inter6));
  inv1  gate1716(.a(G25), .O(gate21inter7));
  inv1  gate1717(.a(G26), .O(gate21inter8));
  nand2 gate1718(.a(gate21inter8), .b(gate21inter7), .O(gate21inter9));
  nand2 gate1719(.a(s_167), .b(gate21inter3), .O(gate21inter10));
  nor2  gate1720(.a(gate21inter10), .b(gate21inter9), .O(gate21inter11));
  nor2  gate1721(.a(gate21inter11), .b(gate21inter6), .O(gate21inter12));
  nand2 gate1722(.a(gate21inter12), .b(gate21inter1), .O(G302));
nand2 gate22( .a(G27), .b(G28), .O(G305) );

  xor2  gate2745(.a(G30), .b(G29), .O(gate23inter0));
  nand2 gate2746(.a(gate23inter0), .b(s_314), .O(gate23inter1));
  and2  gate2747(.a(G30), .b(G29), .O(gate23inter2));
  inv1  gate2748(.a(s_314), .O(gate23inter3));
  inv1  gate2749(.a(s_315), .O(gate23inter4));
  nand2 gate2750(.a(gate23inter4), .b(gate23inter3), .O(gate23inter5));
  nor2  gate2751(.a(gate23inter5), .b(gate23inter2), .O(gate23inter6));
  inv1  gate2752(.a(G29), .O(gate23inter7));
  inv1  gate2753(.a(G30), .O(gate23inter8));
  nand2 gate2754(.a(gate23inter8), .b(gate23inter7), .O(gate23inter9));
  nand2 gate2755(.a(s_315), .b(gate23inter3), .O(gate23inter10));
  nor2  gate2756(.a(gate23inter10), .b(gate23inter9), .O(gate23inter11));
  nor2  gate2757(.a(gate23inter11), .b(gate23inter6), .O(gate23inter12));
  nand2 gate2758(.a(gate23inter12), .b(gate23inter1), .O(G308));
nand2 gate24( .a(G31), .b(G32), .O(G311) );
nand2 gate25( .a(G1), .b(G5), .O(G314) );
nand2 gate26( .a(G9), .b(G13), .O(G317) );
nand2 gate27( .a(G2), .b(G6), .O(G320) );
nand2 gate28( .a(G10), .b(G14), .O(G323) );

  xor2  gate2927(.a(G7), .b(G3), .O(gate29inter0));
  nand2 gate2928(.a(gate29inter0), .b(s_340), .O(gate29inter1));
  and2  gate2929(.a(G7), .b(G3), .O(gate29inter2));
  inv1  gate2930(.a(s_340), .O(gate29inter3));
  inv1  gate2931(.a(s_341), .O(gate29inter4));
  nand2 gate2932(.a(gate29inter4), .b(gate29inter3), .O(gate29inter5));
  nor2  gate2933(.a(gate29inter5), .b(gate29inter2), .O(gate29inter6));
  inv1  gate2934(.a(G3), .O(gate29inter7));
  inv1  gate2935(.a(G7), .O(gate29inter8));
  nand2 gate2936(.a(gate29inter8), .b(gate29inter7), .O(gate29inter9));
  nand2 gate2937(.a(s_341), .b(gate29inter3), .O(gate29inter10));
  nor2  gate2938(.a(gate29inter10), .b(gate29inter9), .O(gate29inter11));
  nor2  gate2939(.a(gate29inter11), .b(gate29inter6), .O(gate29inter12));
  nand2 gate2940(.a(gate29inter12), .b(gate29inter1), .O(G326));

  xor2  gate1247(.a(G15), .b(G11), .O(gate30inter0));
  nand2 gate1248(.a(gate30inter0), .b(s_100), .O(gate30inter1));
  and2  gate1249(.a(G15), .b(G11), .O(gate30inter2));
  inv1  gate1250(.a(s_100), .O(gate30inter3));
  inv1  gate1251(.a(s_101), .O(gate30inter4));
  nand2 gate1252(.a(gate30inter4), .b(gate30inter3), .O(gate30inter5));
  nor2  gate1253(.a(gate30inter5), .b(gate30inter2), .O(gate30inter6));
  inv1  gate1254(.a(G11), .O(gate30inter7));
  inv1  gate1255(.a(G15), .O(gate30inter8));
  nand2 gate1256(.a(gate30inter8), .b(gate30inter7), .O(gate30inter9));
  nand2 gate1257(.a(s_101), .b(gate30inter3), .O(gate30inter10));
  nor2  gate1258(.a(gate30inter10), .b(gate30inter9), .O(gate30inter11));
  nor2  gate1259(.a(gate30inter11), .b(gate30inter6), .O(gate30inter12));
  nand2 gate1260(.a(gate30inter12), .b(gate30inter1), .O(G329));
nand2 gate31( .a(G4), .b(G8), .O(G332) );
nand2 gate32( .a(G12), .b(G16), .O(G335) );
nand2 gate33( .a(G17), .b(G21), .O(G338) );
nand2 gate34( .a(G25), .b(G29), .O(G341) );
nand2 gate35( .a(G18), .b(G22), .O(G344) );
nand2 gate36( .a(G26), .b(G30), .O(G347) );
nand2 gate37( .a(G19), .b(G23), .O(G350) );

  xor2  gate2801(.a(G31), .b(G27), .O(gate38inter0));
  nand2 gate2802(.a(gate38inter0), .b(s_322), .O(gate38inter1));
  and2  gate2803(.a(G31), .b(G27), .O(gate38inter2));
  inv1  gate2804(.a(s_322), .O(gate38inter3));
  inv1  gate2805(.a(s_323), .O(gate38inter4));
  nand2 gate2806(.a(gate38inter4), .b(gate38inter3), .O(gate38inter5));
  nor2  gate2807(.a(gate38inter5), .b(gate38inter2), .O(gate38inter6));
  inv1  gate2808(.a(G27), .O(gate38inter7));
  inv1  gate2809(.a(G31), .O(gate38inter8));
  nand2 gate2810(.a(gate38inter8), .b(gate38inter7), .O(gate38inter9));
  nand2 gate2811(.a(s_323), .b(gate38inter3), .O(gate38inter10));
  nor2  gate2812(.a(gate38inter10), .b(gate38inter9), .O(gate38inter11));
  nor2  gate2813(.a(gate38inter11), .b(gate38inter6), .O(gate38inter12));
  nand2 gate2814(.a(gate38inter12), .b(gate38inter1), .O(G353));
nand2 gate39( .a(G20), .b(G24), .O(G356) );

  xor2  gate2213(.a(G32), .b(G28), .O(gate40inter0));
  nand2 gate2214(.a(gate40inter0), .b(s_238), .O(gate40inter1));
  and2  gate2215(.a(G32), .b(G28), .O(gate40inter2));
  inv1  gate2216(.a(s_238), .O(gate40inter3));
  inv1  gate2217(.a(s_239), .O(gate40inter4));
  nand2 gate2218(.a(gate40inter4), .b(gate40inter3), .O(gate40inter5));
  nor2  gate2219(.a(gate40inter5), .b(gate40inter2), .O(gate40inter6));
  inv1  gate2220(.a(G28), .O(gate40inter7));
  inv1  gate2221(.a(G32), .O(gate40inter8));
  nand2 gate2222(.a(gate40inter8), .b(gate40inter7), .O(gate40inter9));
  nand2 gate2223(.a(s_239), .b(gate40inter3), .O(gate40inter10));
  nor2  gate2224(.a(gate40inter10), .b(gate40inter9), .O(gate40inter11));
  nor2  gate2225(.a(gate40inter11), .b(gate40inter6), .O(gate40inter12));
  nand2 gate2226(.a(gate40inter12), .b(gate40inter1), .O(G359));
nand2 gate41( .a(G1), .b(G266), .O(G362) );
nand2 gate42( .a(G2), .b(G266), .O(G363) );

  xor2  gate1079(.a(G269), .b(G3), .O(gate43inter0));
  nand2 gate1080(.a(gate43inter0), .b(s_76), .O(gate43inter1));
  and2  gate1081(.a(G269), .b(G3), .O(gate43inter2));
  inv1  gate1082(.a(s_76), .O(gate43inter3));
  inv1  gate1083(.a(s_77), .O(gate43inter4));
  nand2 gate1084(.a(gate43inter4), .b(gate43inter3), .O(gate43inter5));
  nor2  gate1085(.a(gate43inter5), .b(gate43inter2), .O(gate43inter6));
  inv1  gate1086(.a(G3), .O(gate43inter7));
  inv1  gate1087(.a(G269), .O(gate43inter8));
  nand2 gate1088(.a(gate43inter8), .b(gate43inter7), .O(gate43inter9));
  nand2 gate1089(.a(s_77), .b(gate43inter3), .O(gate43inter10));
  nor2  gate1090(.a(gate43inter10), .b(gate43inter9), .O(gate43inter11));
  nor2  gate1091(.a(gate43inter11), .b(gate43inter6), .O(gate43inter12));
  nand2 gate1092(.a(gate43inter12), .b(gate43inter1), .O(G364));

  xor2  gate2017(.a(G269), .b(G4), .O(gate44inter0));
  nand2 gate2018(.a(gate44inter0), .b(s_210), .O(gate44inter1));
  and2  gate2019(.a(G269), .b(G4), .O(gate44inter2));
  inv1  gate2020(.a(s_210), .O(gate44inter3));
  inv1  gate2021(.a(s_211), .O(gate44inter4));
  nand2 gate2022(.a(gate44inter4), .b(gate44inter3), .O(gate44inter5));
  nor2  gate2023(.a(gate44inter5), .b(gate44inter2), .O(gate44inter6));
  inv1  gate2024(.a(G4), .O(gate44inter7));
  inv1  gate2025(.a(G269), .O(gate44inter8));
  nand2 gate2026(.a(gate44inter8), .b(gate44inter7), .O(gate44inter9));
  nand2 gate2027(.a(s_211), .b(gate44inter3), .O(gate44inter10));
  nor2  gate2028(.a(gate44inter10), .b(gate44inter9), .O(gate44inter11));
  nor2  gate2029(.a(gate44inter11), .b(gate44inter6), .O(gate44inter12));
  nand2 gate2030(.a(gate44inter12), .b(gate44inter1), .O(G365));
nand2 gate45( .a(G5), .b(G272), .O(G366) );

  xor2  gate771(.a(G272), .b(G6), .O(gate46inter0));
  nand2 gate772(.a(gate46inter0), .b(s_32), .O(gate46inter1));
  and2  gate773(.a(G272), .b(G6), .O(gate46inter2));
  inv1  gate774(.a(s_32), .O(gate46inter3));
  inv1  gate775(.a(s_33), .O(gate46inter4));
  nand2 gate776(.a(gate46inter4), .b(gate46inter3), .O(gate46inter5));
  nor2  gate777(.a(gate46inter5), .b(gate46inter2), .O(gate46inter6));
  inv1  gate778(.a(G6), .O(gate46inter7));
  inv1  gate779(.a(G272), .O(gate46inter8));
  nand2 gate780(.a(gate46inter8), .b(gate46inter7), .O(gate46inter9));
  nand2 gate781(.a(s_33), .b(gate46inter3), .O(gate46inter10));
  nor2  gate782(.a(gate46inter10), .b(gate46inter9), .O(gate46inter11));
  nor2  gate783(.a(gate46inter11), .b(gate46inter6), .O(gate46inter12));
  nand2 gate784(.a(gate46inter12), .b(gate46inter1), .O(G367));

  xor2  gate1303(.a(G275), .b(G7), .O(gate47inter0));
  nand2 gate1304(.a(gate47inter0), .b(s_108), .O(gate47inter1));
  and2  gate1305(.a(G275), .b(G7), .O(gate47inter2));
  inv1  gate1306(.a(s_108), .O(gate47inter3));
  inv1  gate1307(.a(s_109), .O(gate47inter4));
  nand2 gate1308(.a(gate47inter4), .b(gate47inter3), .O(gate47inter5));
  nor2  gate1309(.a(gate47inter5), .b(gate47inter2), .O(gate47inter6));
  inv1  gate1310(.a(G7), .O(gate47inter7));
  inv1  gate1311(.a(G275), .O(gate47inter8));
  nand2 gate1312(.a(gate47inter8), .b(gate47inter7), .O(gate47inter9));
  nand2 gate1313(.a(s_109), .b(gate47inter3), .O(gate47inter10));
  nor2  gate1314(.a(gate47inter10), .b(gate47inter9), .O(gate47inter11));
  nor2  gate1315(.a(gate47inter11), .b(gate47inter6), .O(gate47inter12));
  nand2 gate1316(.a(gate47inter12), .b(gate47inter1), .O(G368));
nand2 gate48( .a(G8), .b(G275), .O(G369) );

  xor2  gate1373(.a(G278), .b(G9), .O(gate49inter0));
  nand2 gate1374(.a(gate49inter0), .b(s_118), .O(gate49inter1));
  and2  gate1375(.a(G278), .b(G9), .O(gate49inter2));
  inv1  gate1376(.a(s_118), .O(gate49inter3));
  inv1  gate1377(.a(s_119), .O(gate49inter4));
  nand2 gate1378(.a(gate49inter4), .b(gate49inter3), .O(gate49inter5));
  nor2  gate1379(.a(gate49inter5), .b(gate49inter2), .O(gate49inter6));
  inv1  gate1380(.a(G9), .O(gate49inter7));
  inv1  gate1381(.a(G278), .O(gate49inter8));
  nand2 gate1382(.a(gate49inter8), .b(gate49inter7), .O(gate49inter9));
  nand2 gate1383(.a(s_119), .b(gate49inter3), .O(gate49inter10));
  nor2  gate1384(.a(gate49inter10), .b(gate49inter9), .O(gate49inter11));
  nor2  gate1385(.a(gate49inter11), .b(gate49inter6), .O(gate49inter12));
  nand2 gate1386(.a(gate49inter12), .b(gate49inter1), .O(G370));

  xor2  gate2633(.a(G278), .b(G10), .O(gate50inter0));
  nand2 gate2634(.a(gate50inter0), .b(s_298), .O(gate50inter1));
  and2  gate2635(.a(G278), .b(G10), .O(gate50inter2));
  inv1  gate2636(.a(s_298), .O(gate50inter3));
  inv1  gate2637(.a(s_299), .O(gate50inter4));
  nand2 gate2638(.a(gate50inter4), .b(gate50inter3), .O(gate50inter5));
  nor2  gate2639(.a(gate50inter5), .b(gate50inter2), .O(gate50inter6));
  inv1  gate2640(.a(G10), .O(gate50inter7));
  inv1  gate2641(.a(G278), .O(gate50inter8));
  nand2 gate2642(.a(gate50inter8), .b(gate50inter7), .O(gate50inter9));
  nand2 gate2643(.a(s_299), .b(gate50inter3), .O(gate50inter10));
  nor2  gate2644(.a(gate50inter10), .b(gate50inter9), .O(gate50inter11));
  nor2  gate2645(.a(gate50inter11), .b(gate50inter6), .O(gate50inter12));
  nand2 gate2646(.a(gate50inter12), .b(gate50inter1), .O(G371));

  xor2  gate575(.a(G281), .b(G11), .O(gate51inter0));
  nand2 gate576(.a(gate51inter0), .b(s_4), .O(gate51inter1));
  and2  gate577(.a(G281), .b(G11), .O(gate51inter2));
  inv1  gate578(.a(s_4), .O(gate51inter3));
  inv1  gate579(.a(s_5), .O(gate51inter4));
  nand2 gate580(.a(gate51inter4), .b(gate51inter3), .O(gate51inter5));
  nor2  gate581(.a(gate51inter5), .b(gate51inter2), .O(gate51inter6));
  inv1  gate582(.a(G11), .O(gate51inter7));
  inv1  gate583(.a(G281), .O(gate51inter8));
  nand2 gate584(.a(gate51inter8), .b(gate51inter7), .O(gate51inter9));
  nand2 gate585(.a(s_5), .b(gate51inter3), .O(gate51inter10));
  nor2  gate586(.a(gate51inter10), .b(gate51inter9), .O(gate51inter11));
  nor2  gate587(.a(gate51inter11), .b(gate51inter6), .O(gate51inter12));
  nand2 gate588(.a(gate51inter12), .b(gate51inter1), .O(G372));
nand2 gate52( .a(G12), .b(G281), .O(G373) );
nand2 gate53( .a(G13), .b(G284), .O(G374) );
nand2 gate54( .a(G14), .b(G284), .O(G375) );

  xor2  gate2227(.a(G287), .b(G15), .O(gate55inter0));
  nand2 gate2228(.a(gate55inter0), .b(s_240), .O(gate55inter1));
  and2  gate2229(.a(G287), .b(G15), .O(gate55inter2));
  inv1  gate2230(.a(s_240), .O(gate55inter3));
  inv1  gate2231(.a(s_241), .O(gate55inter4));
  nand2 gate2232(.a(gate55inter4), .b(gate55inter3), .O(gate55inter5));
  nor2  gate2233(.a(gate55inter5), .b(gate55inter2), .O(gate55inter6));
  inv1  gate2234(.a(G15), .O(gate55inter7));
  inv1  gate2235(.a(G287), .O(gate55inter8));
  nand2 gate2236(.a(gate55inter8), .b(gate55inter7), .O(gate55inter9));
  nand2 gate2237(.a(s_241), .b(gate55inter3), .O(gate55inter10));
  nor2  gate2238(.a(gate55inter10), .b(gate55inter9), .O(gate55inter11));
  nor2  gate2239(.a(gate55inter11), .b(gate55inter6), .O(gate55inter12));
  nand2 gate2240(.a(gate55inter12), .b(gate55inter1), .O(G376));

  xor2  gate1751(.a(G287), .b(G16), .O(gate56inter0));
  nand2 gate1752(.a(gate56inter0), .b(s_172), .O(gate56inter1));
  and2  gate1753(.a(G287), .b(G16), .O(gate56inter2));
  inv1  gate1754(.a(s_172), .O(gate56inter3));
  inv1  gate1755(.a(s_173), .O(gate56inter4));
  nand2 gate1756(.a(gate56inter4), .b(gate56inter3), .O(gate56inter5));
  nor2  gate1757(.a(gate56inter5), .b(gate56inter2), .O(gate56inter6));
  inv1  gate1758(.a(G16), .O(gate56inter7));
  inv1  gate1759(.a(G287), .O(gate56inter8));
  nand2 gate1760(.a(gate56inter8), .b(gate56inter7), .O(gate56inter9));
  nand2 gate1761(.a(s_173), .b(gate56inter3), .O(gate56inter10));
  nor2  gate1762(.a(gate56inter10), .b(gate56inter9), .O(gate56inter11));
  nor2  gate1763(.a(gate56inter11), .b(gate56inter6), .O(gate56inter12));
  nand2 gate1764(.a(gate56inter12), .b(gate56inter1), .O(G377));
nand2 gate57( .a(G17), .b(G290), .O(G378) );
nand2 gate58( .a(G18), .b(G290), .O(G379) );

  xor2  gate659(.a(G293), .b(G19), .O(gate59inter0));
  nand2 gate660(.a(gate59inter0), .b(s_16), .O(gate59inter1));
  and2  gate661(.a(G293), .b(G19), .O(gate59inter2));
  inv1  gate662(.a(s_16), .O(gate59inter3));
  inv1  gate663(.a(s_17), .O(gate59inter4));
  nand2 gate664(.a(gate59inter4), .b(gate59inter3), .O(gate59inter5));
  nor2  gate665(.a(gate59inter5), .b(gate59inter2), .O(gate59inter6));
  inv1  gate666(.a(G19), .O(gate59inter7));
  inv1  gate667(.a(G293), .O(gate59inter8));
  nand2 gate668(.a(gate59inter8), .b(gate59inter7), .O(gate59inter9));
  nand2 gate669(.a(s_17), .b(gate59inter3), .O(gate59inter10));
  nor2  gate670(.a(gate59inter10), .b(gate59inter9), .O(gate59inter11));
  nor2  gate671(.a(gate59inter11), .b(gate59inter6), .O(gate59inter12));
  nand2 gate672(.a(gate59inter12), .b(gate59inter1), .O(G380));
nand2 gate60( .a(G20), .b(G293), .O(G381) );
nand2 gate61( .a(G21), .b(G296), .O(G382) );

  xor2  gate2535(.a(G296), .b(G22), .O(gate62inter0));
  nand2 gate2536(.a(gate62inter0), .b(s_284), .O(gate62inter1));
  and2  gate2537(.a(G296), .b(G22), .O(gate62inter2));
  inv1  gate2538(.a(s_284), .O(gate62inter3));
  inv1  gate2539(.a(s_285), .O(gate62inter4));
  nand2 gate2540(.a(gate62inter4), .b(gate62inter3), .O(gate62inter5));
  nor2  gate2541(.a(gate62inter5), .b(gate62inter2), .O(gate62inter6));
  inv1  gate2542(.a(G22), .O(gate62inter7));
  inv1  gate2543(.a(G296), .O(gate62inter8));
  nand2 gate2544(.a(gate62inter8), .b(gate62inter7), .O(gate62inter9));
  nand2 gate2545(.a(s_285), .b(gate62inter3), .O(gate62inter10));
  nor2  gate2546(.a(gate62inter10), .b(gate62inter9), .O(gate62inter11));
  nor2  gate2547(.a(gate62inter11), .b(gate62inter6), .O(gate62inter12));
  nand2 gate2548(.a(gate62inter12), .b(gate62inter1), .O(G383));

  xor2  gate981(.a(G299), .b(G23), .O(gate63inter0));
  nand2 gate982(.a(gate63inter0), .b(s_62), .O(gate63inter1));
  and2  gate983(.a(G299), .b(G23), .O(gate63inter2));
  inv1  gate984(.a(s_62), .O(gate63inter3));
  inv1  gate985(.a(s_63), .O(gate63inter4));
  nand2 gate986(.a(gate63inter4), .b(gate63inter3), .O(gate63inter5));
  nor2  gate987(.a(gate63inter5), .b(gate63inter2), .O(gate63inter6));
  inv1  gate988(.a(G23), .O(gate63inter7));
  inv1  gate989(.a(G299), .O(gate63inter8));
  nand2 gate990(.a(gate63inter8), .b(gate63inter7), .O(gate63inter9));
  nand2 gate991(.a(s_63), .b(gate63inter3), .O(gate63inter10));
  nor2  gate992(.a(gate63inter10), .b(gate63inter9), .O(gate63inter11));
  nor2  gate993(.a(gate63inter11), .b(gate63inter6), .O(gate63inter12));
  nand2 gate994(.a(gate63inter12), .b(gate63inter1), .O(G384));

  xor2  gate1121(.a(G299), .b(G24), .O(gate64inter0));
  nand2 gate1122(.a(gate64inter0), .b(s_82), .O(gate64inter1));
  and2  gate1123(.a(G299), .b(G24), .O(gate64inter2));
  inv1  gate1124(.a(s_82), .O(gate64inter3));
  inv1  gate1125(.a(s_83), .O(gate64inter4));
  nand2 gate1126(.a(gate64inter4), .b(gate64inter3), .O(gate64inter5));
  nor2  gate1127(.a(gate64inter5), .b(gate64inter2), .O(gate64inter6));
  inv1  gate1128(.a(G24), .O(gate64inter7));
  inv1  gate1129(.a(G299), .O(gate64inter8));
  nand2 gate1130(.a(gate64inter8), .b(gate64inter7), .O(gate64inter9));
  nand2 gate1131(.a(s_83), .b(gate64inter3), .O(gate64inter10));
  nor2  gate1132(.a(gate64inter10), .b(gate64inter9), .O(gate64inter11));
  nor2  gate1133(.a(gate64inter11), .b(gate64inter6), .O(gate64inter12));
  nand2 gate1134(.a(gate64inter12), .b(gate64inter1), .O(G385));
nand2 gate65( .a(G25), .b(G302), .O(G386) );

  xor2  gate589(.a(G302), .b(G26), .O(gate66inter0));
  nand2 gate590(.a(gate66inter0), .b(s_6), .O(gate66inter1));
  and2  gate591(.a(G302), .b(G26), .O(gate66inter2));
  inv1  gate592(.a(s_6), .O(gate66inter3));
  inv1  gate593(.a(s_7), .O(gate66inter4));
  nand2 gate594(.a(gate66inter4), .b(gate66inter3), .O(gate66inter5));
  nor2  gate595(.a(gate66inter5), .b(gate66inter2), .O(gate66inter6));
  inv1  gate596(.a(G26), .O(gate66inter7));
  inv1  gate597(.a(G302), .O(gate66inter8));
  nand2 gate598(.a(gate66inter8), .b(gate66inter7), .O(gate66inter9));
  nand2 gate599(.a(s_7), .b(gate66inter3), .O(gate66inter10));
  nor2  gate600(.a(gate66inter10), .b(gate66inter9), .O(gate66inter11));
  nor2  gate601(.a(gate66inter11), .b(gate66inter6), .O(gate66inter12));
  nand2 gate602(.a(gate66inter12), .b(gate66inter1), .O(G387));
nand2 gate67( .a(G27), .b(G305), .O(G388) );
nand2 gate68( .a(G28), .b(G305), .O(G389) );

  xor2  gate1961(.a(G308), .b(G29), .O(gate69inter0));
  nand2 gate1962(.a(gate69inter0), .b(s_202), .O(gate69inter1));
  and2  gate1963(.a(G308), .b(G29), .O(gate69inter2));
  inv1  gate1964(.a(s_202), .O(gate69inter3));
  inv1  gate1965(.a(s_203), .O(gate69inter4));
  nand2 gate1966(.a(gate69inter4), .b(gate69inter3), .O(gate69inter5));
  nor2  gate1967(.a(gate69inter5), .b(gate69inter2), .O(gate69inter6));
  inv1  gate1968(.a(G29), .O(gate69inter7));
  inv1  gate1969(.a(G308), .O(gate69inter8));
  nand2 gate1970(.a(gate69inter8), .b(gate69inter7), .O(gate69inter9));
  nand2 gate1971(.a(s_203), .b(gate69inter3), .O(gate69inter10));
  nor2  gate1972(.a(gate69inter10), .b(gate69inter9), .O(gate69inter11));
  nor2  gate1973(.a(gate69inter11), .b(gate69inter6), .O(gate69inter12));
  nand2 gate1974(.a(gate69inter12), .b(gate69inter1), .O(G390));
nand2 gate70( .a(G30), .b(G308), .O(G391) );

  xor2  gate1555(.a(G311), .b(G31), .O(gate71inter0));
  nand2 gate1556(.a(gate71inter0), .b(s_144), .O(gate71inter1));
  and2  gate1557(.a(G311), .b(G31), .O(gate71inter2));
  inv1  gate1558(.a(s_144), .O(gate71inter3));
  inv1  gate1559(.a(s_145), .O(gate71inter4));
  nand2 gate1560(.a(gate71inter4), .b(gate71inter3), .O(gate71inter5));
  nor2  gate1561(.a(gate71inter5), .b(gate71inter2), .O(gate71inter6));
  inv1  gate1562(.a(G31), .O(gate71inter7));
  inv1  gate1563(.a(G311), .O(gate71inter8));
  nand2 gate1564(.a(gate71inter8), .b(gate71inter7), .O(gate71inter9));
  nand2 gate1565(.a(s_145), .b(gate71inter3), .O(gate71inter10));
  nor2  gate1566(.a(gate71inter10), .b(gate71inter9), .O(gate71inter11));
  nor2  gate1567(.a(gate71inter11), .b(gate71inter6), .O(gate71inter12));
  nand2 gate1568(.a(gate71inter12), .b(gate71inter1), .O(G392));

  xor2  gate2549(.a(G311), .b(G32), .O(gate72inter0));
  nand2 gate2550(.a(gate72inter0), .b(s_286), .O(gate72inter1));
  and2  gate2551(.a(G311), .b(G32), .O(gate72inter2));
  inv1  gate2552(.a(s_286), .O(gate72inter3));
  inv1  gate2553(.a(s_287), .O(gate72inter4));
  nand2 gate2554(.a(gate72inter4), .b(gate72inter3), .O(gate72inter5));
  nor2  gate2555(.a(gate72inter5), .b(gate72inter2), .O(gate72inter6));
  inv1  gate2556(.a(G32), .O(gate72inter7));
  inv1  gate2557(.a(G311), .O(gate72inter8));
  nand2 gate2558(.a(gate72inter8), .b(gate72inter7), .O(gate72inter9));
  nand2 gate2559(.a(s_287), .b(gate72inter3), .O(gate72inter10));
  nor2  gate2560(.a(gate72inter10), .b(gate72inter9), .O(gate72inter11));
  nor2  gate2561(.a(gate72inter11), .b(gate72inter6), .O(gate72inter12));
  nand2 gate2562(.a(gate72inter12), .b(gate72inter1), .O(G393));

  xor2  gate2143(.a(G314), .b(G1), .O(gate73inter0));
  nand2 gate2144(.a(gate73inter0), .b(s_228), .O(gate73inter1));
  and2  gate2145(.a(G314), .b(G1), .O(gate73inter2));
  inv1  gate2146(.a(s_228), .O(gate73inter3));
  inv1  gate2147(.a(s_229), .O(gate73inter4));
  nand2 gate2148(.a(gate73inter4), .b(gate73inter3), .O(gate73inter5));
  nor2  gate2149(.a(gate73inter5), .b(gate73inter2), .O(gate73inter6));
  inv1  gate2150(.a(G1), .O(gate73inter7));
  inv1  gate2151(.a(G314), .O(gate73inter8));
  nand2 gate2152(.a(gate73inter8), .b(gate73inter7), .O(gate73inter9));
  nand2 gate2153(.a(s_229), .b(gate73inter3), .O(gate73inter10));
  nor2  gate2154(.a(gate73inter10), .b(gate73inter9), .O(gate73inter11));
  nor2  gate2155(.a(gate73inter11), .b(gate73inter6), .O(gate73inter12));
  nand2 gate2156(.a(gate73inter12), .b(gate73inter1), .O(G394));
nand2 gate74( .a(G5), .b(G314), .O(G395) );

  xor2  gate1793(.a(G317), .b(G9), .O(gate75inter0));
  nand2 gate1794(.a(gate75inter0), .b(s_178), .O(gate75inter1));
  and2  gate1795(.a(G317), .b(G9), .O(gate75inter2));
  inv1  gate1796(.a(s_178), .O(gate75inter3));
  inv1  gate1797(.a(s_179), .O(gate75inter4));
  nand2 gate1798(.a(gate75inter4), .b(gate75inter3), .O(gate75inter5));
  nor2  gate1799(.a(gate75inter5), .b(gate75inter2), .O(gate75inter6));
  inv1  gate1800(.a(G9), .O(gate75inter7));
  inv1  gate1801(.a(G317), .O(gate75inter8));
  nand2 gate1802(.a(gate75inter8), .b(gate75inter7), .O(gate75inter9));
  nand2 gate1803(.a(s_179), .b(gate75inter3), .O(gate75inter10));
  nor2  gate1804(.a(gate75inter10), .b(gate75inter9), .O(gate75inter11));
  nor2  gate1805(.a(gate75inter11), .b(gate75inter6), .O(gate75inter12));
  nand2 gate1806(.a(gate75inter12), .b(gate75inter1), .O(G396));
nand2 gate76( .a(G13), .b(G317), .O(G397) );

  xor2  gate1037(.a(G320), .b(G2), .O(gate77inter0));
  nand2 gate1038(.a(gate77inter0), .b(s_70), .O(gate77inter1));
  and2  gate1039(.a(G320), .b(G2), .O(gate77inter2));
  inv1  gate1040(.a(s_70), .O(gate77inter3));
  inv1  gate1041(.a(s_71), .O(gate77inter4));
  nand2 gate1042(.a(gate77inter4), .b(gate77inter3), .O(gate77inter5));
  nor2  gate1043(.a(gate77inter5), .b(gate77inter2), .O(gate77inter6));
  inv1  gate1044(.a(G2), .O(gate77inter7));
  inv1  gate1045(.a(G320), .O(gate77inter8));
  nand2 gate1046(.a(gate77inter8), .b(gate77inter7), .O(gate77inter9));
  nand2 gate1047(.a(s_71), .b(gate77inter3), .O(gate77inter10));
  nor2  gate1048(.a(gate77inter10), .b(gate77inter9), .O(gate77inter11));
  nor2  gate1049(.a(gate77inter11), .b(gate77inter6), .O(gate77inter12));
  nand2 gate1050(.a(gate77inter12), .b(gate77inter1), .O(G398));
nand2 gate78( .a(G6), .b(G320), .O(G399) );
nand2 gate79( .a(G10), .b(G323), .O(G400) );
nand2 gate80( .a(G14), .b(G323), .O(G401) );

  xor2  gate1233(.a(G326), .b(G3), .O(gate81inter0));
  nand2 gate1234(.a(gate81inter0), .b(s_98), .O(gate81inter1));
  and2  gate1235(.a(G326), .b(G3), .O(gate81inter2));
  inv1  gate1236(.a(s_98), .O(gate81inter3));
  inv1  gate1237(.a(s_99), .O(gate81inter4));
  nand2 gate1238(.a(gate81inter4), .b(gate81inter3), .O(gate81inter5));
  nor2  gate1239(.a(gate81inter5), .b(gate81inter2), .O(gate81inter6));
  inv1  gate1240(.a(G3), .O(gate81inter7));
  inv1  gate1241(.a(G326), .O(gate81inter8));
  nand2 gate1242(.a(gate81inter8), .b(gate81inter7), .O(gate81inter9));
  nand2 gate1243(.a(s_99), .b(gate81inter3), .O(gate81inter10));
  nor2  gate1244(.a(gate81inter10), .b(gate81inter9), .O(gate81inter11));
  nor2  gate1245(.a(gate81inter11), .b(gate81inter6), .O(gate81inter12));
  nand2 gate1246(.a(gate81inter12), .b(gate81inter1), .O(G402));
nand2 gate82( .a(G7), .b(G326), .O(G403) );
nand2 gate83( .a(G11), .b(G329), .O(G404) );

  xor2  gate1317(.a(G329), .b(G15), .O(gate84inter0));
  nand2 gate1318(.a(gate84inter0), .b(s_110), .O(gate84inter1));
  and2  gate1319(.a(G329), .b(G15), .O(gate84inter2));
  inv1  gate1320(.a(s_110), .O(gate84inter3));
  inv1  gate1321(.a(s_111), .O(gate84inter4));
  nand2 gate1322(.a(gate84inter4), .b(gate84inter3), .O(gate84inter5));
  nor2  gate1323(.a(gate84inter5), .b(gate84inter2), .O(gate84inter6));
  inv1  gate1324(.a(G15), .O(gate84inter7));
  inv1  gate1325(.a(G329), .O(gate84inter8));
  nand2 gate1326(.a(gate84inter8), .b(gate84inter7), .O(gate84inter9));
  nand2 gate1327(.a(s_111), .b(gate84inter3), .O(gate84inter10));
  nor2  gate1328(.a(gate84inter10), .b(gate84inter9), .O(gate84inter11));
  nor2  gate1329(.a(gate84inter11), .b(gate84inter6), .O(gate84inter12));
  nand2 gate1330(.a(gate84inter12), .b(gate84inter1), .O(G405));
nand2 gate85( .a(G4), .b(G332), .O(G406) );

  xor2  gate2325(.a(G332), .b(G8), .O(gate86inter0));
  nand2 gate2326(.a(gate86inter0), .b(s_254), .O(gate86inter1));
  and2  gate2327(.a(G332), .b(G8), .O(gate86inter2));
  inv1  gate2328(.a(s_254), .O(gate86inter3));
  inv1  gate2329(.a(s_255), .O(gate86inter4));
  nand2 gate2330(.a(gate86inter4), .b(gate86inter3), .O(gate86inter5));
  nor2  gate2331(.a(gate86inter5), .b(gate86inter2), .O(gate86inter6));
  inv1  gate2332(.a(G8), .O(gate86inter7));
  inv1  gate2333(.a(G332), .O(gate86inter8));
  nand2 gate2334(.a(gate86inter8), .b(gate86inter7), .O(gate86inter9));
  nand2 gate2335(.a(s_255), .b(gate86inter3), .O(gate86inter10));
  nor2  gate2336(.a(gate86inter10), .b(gate86inter9), .O(gate86inter11));
  nor2  gate2337(.a(gate86inter11), .b(gate86inter6), .O(gate86inter12));
  nand2 gate2338(.a(gate86inter12), .b(gate86inter1), .O(G407));
nand2 gate87( .a(G12), .b(G335), .O(G408) );
nand2 gate88( .a(G16), .b(G335), .O(G409) );
nand2 gate89( .a(G17), .b(G338), .O(G410) );
nand2 gate90( .a(G21), .b(G338), .O(G411) );

  xor2  gate2815(.a(G341), .b(G25), .O(gate91inter0));
  nand2 gate2816(.a(gate91inter0), .b(s_324), .O(gate91inter1));
  and2  gate2817(.a(G341), .b(G25), .O(gate91inter2));
  inv1  gate2818(.a(s_324), .O(gate91inter3));
  inv1  gate2819(.a(s_325), .O(gate91inter4));
  nand2 gate2820(.a(gate91inter4), .b(gate91inter3), .O(gate91inter5));
  nor2  gate2821(.a(gate91inter5), .b(gate91inter2), .O(gate91inter6));
  inv1  gate2822(.a(G25), .O(gate91inter7));
  inv1  gate2823(.a(G341), .O(gate91inter8));
  nand2 gate2824(.a(gate91inter8), .b(gate91inter7), .O(gate91inter9));
  nand2 gate2825(.a(s_325), .b(gate91inter3), .O(gate91inter10));
  nor2  gate2826(.a(gate91inter10), .b(gate91inter9), .O(gate91inter11));
  nor2  gate2827(.a(gate91inter11), .b(gate91inter6), .O(gate91inter12));
  nand2 gate2828(.a(gate91inter12), .b(gate91inter1), .O(G412));

  xor2  gate2605(.a(G341), .b(G29), .O(gate92inter0));
  nand2 gate2606(.a(gate92inter0), .b(s_294), .O(gate92inter1));
  and2  gate2607(.a(G341), .b(G29), .O(gate92inter2));
  inv1  gate2608(.a(s_294), .O(gate92inter3));
  inv1  gate2609(.a(s_295), .O(gate92inter4));
  nand2 gate2610(.a(gate92inter4), .b(gate92inter3), .O(gate92inter5));
  nor2  gate2611(.a(gate92inter5), .b(gate92inter2), .O(gate92inter6));
  inv1  gate2612(.a(G29), .O(gate92inter7));
  inv1  gate2613(.a(G341), .O(gate92inter8));
  nand2 gate2614(.a(gate92inter8), .b(gate92inter7), .O(gate92inter9));
  nand2 gate2615(.a(s_295), .b(gate92inter3), .O(gate92inter10));
  nor2  gate2616(.a(gate92inter10), .b(gate92inter9), .O(gate92inter11));
  nor2  gate2617(.a(gate92inter11), .b(gate92inter6), .O(gate92inter12));
  nand2 gate2618(.a(gate92inter12), .b(gate92inter1), .O(G413));

  xor2  gate2241(.a(G344), .b(G18), .O(gate93inter0));
  nand2 gate2242(.a(gate93inter0), .b(s_242), .O(gate93inter1));
  and2  gate2243(.a(G344), .b(G18), .O(gate93inter2));
  inv1  gate2244(.a(s_242), .O(gate93inter3));
  inv1  gate2245(.a(s_243), .O(gate93inter4));
  nand2 gate2246(.a(gate93inter4), .b(gate93inter3), .O(gate93inter5));
  nor2  gate2247(.a(gate93inter5), .b(gate93inter2), .O(gate93inter6));
  inv1  gate2248(.a(G18), .O(gate93inter7));
  inv1  gate2249(.a(G344), .O(gate93inter8));
  nand2 gate2250(.a(gate93inter8), .b(gate93inter7), .O(gate93inter9));
  nand2 gate2251(.a(s_243), .b(gate93inter3), .O(gate93inter10));
  nor2  gate2252(.a(gate93inter10), .b(gate93inter9), .O(gate93inter11));
  nor2  gate2253(.a(gate93inter11), .b(gate93inter6), .O(gate93inter12));
  nand2 gate2254(.a(gate93inter12), .b(gate93inter1), .O(G414));
nand2 gate94( .a(G22), .b(G344), .O(G415) );
nand2 gate95( .a(G26), .b(G347), .O(G416) );

  xor2  gate2829(.a(G347), .b(G30), .O(gate96inter0));
  nand2 gate2830(.a(gate96inter0), .b(s_326), .O(gate96inter1));
  and2  gate2831(.a(G347), .b(G30), .O(gate96inter2));
  inv1  gate2832(.a(s_326), .O(gate96inter3));
  inv1  gate2833(.a(s_327), .O(gate96inter4));
  nand2 gate2834(.a(gate96inter4), .b(gate96inter3), .O(gate96inter5));
  nor2  gate2835(.a(gate96inter5), .b(gate96inter2), .O(gate96inter6));
  inv1  gate2836(.a(G30), .O(gate96inter7));
  inv1  gate2837(.a(G347), .O(gate96inter8));
  nand2 gate2838(.a(gate96inter8), .b(gate96inter7), .O(gate96inter9));
  nand2 gate2839(.a(s_327), .b(gate96inter3), .O(gate96inter10));
  nor2  gate2840(.a(gate96inter10), .b(gate96inter9), .O(gate96inter11));
  nor2  gate2841(.a(gate96inter11), .b(gate96inter6), .O(gate96inter12));
  nand2 gate2842(.a(gate96inter12), .b(gate96inter1), .O(G417));

  xor2  gate1863(.a(G350), .b(G19), .O(gate97inter0));
  nand2 gate1864(.a(gate97inter0), .b(s_188), .O(gate97inter1));
  and2  gate1865(.a(G350), .b(G19), .O(gate97inter2));
  inv1  gate1866(.a(s_188), .O(gate97inter3));
  inv1  gate1867(.a(s_189), .O(gate97inter4));
  nand2 gate1868(.a(gate97inter4), .b(gate97inter3), .O(gate97inter5));
  nor2  gate1869(.a(gate97inter5), .b(gate97inter2), .O(gate97inter6));
  inv1  gate1870(.a(G19), .O(gate97inter7));
  inv1  gate1871(.a(G350), .O(gate97inter8));
  nand2 gate1872(.a(gate97inter8), .b(gate97inter7), .O(gate97inter9));
  nand2 gate1873(.a(s_189), .b(gate97inter3), .O(gate97inter10));
  nor2  gate1874(.a(gate97inter10), .b(gate97inter9), .O(gate97inter11));
  nor2  gate1875(.a(gate97inter11), .b(gate97inter6), .O(gate97inter12));
  nand2 gate1876(.a(gate97inter12), .b(gate97inter1), .O(G418));

  xor2  gate2703(.a(G350), .b(G23), .O(gate98inter0));
  nand2 gate2704(.a(gate98inter0), .b(s_308), .O(gate98inter1));
  and2  gate2705(.a(G350), .b(G23), .O(gate98inter2));
  inv1  gate2706(.a(s_308), .O(gate98inter3));
  inv1  gate2707(.a(s_309), .O(gate98inter4));
  nand2 gate2708(.a(gate98inter4), .b(gate98inter3), .O(gate98inter5));
  nor2  gate2709(.a(gate98inter5), .b(gate98inter2), .O(gate98inter6));
  inv1  gate2710(.a(G23), .O(gate98inter7));
  inv1  gate2711(.a(G350), .O(gate98inter8));
  nand2 gate2712(.a(gate98inter8), .b(gate98inter7), .O(gate98inter9));
  nand2 gate2713(.a(s_309), .b(gate98inter3), .O(gate98inter10));
  nor2  gate2714(.a(gate98inter10), .b(gate98inter9), .O(gate98inter11));
  nor2  gate2715(.a(gate98inter11), .b(gate98inter6), .O(gate98inter12));
  nand2 gate2716(.a(gate98inter12), .b(gate98inter1), .O(G419));
nand2 gate99( .a(G27), .b(G353), .O(G420) );

  xor2  gate1443(.a(G353), .b(G31), .O(gate100inter0));
  nand2 gate1444(.a(gate100inter0), .b(s_128), .O(gate100inter1));
  and2  gate1445(.a(G353), .b(G31), .O(gate100inter2));
  inv1  gate1446(.a(s_128), .O(gate100inter3));
  inv1  gate1447(.a(s_129), .O(gate100inter4));
  nand2 gate1448(.a(gate100inter4), .b(gate100inter3), .O(gate100inter5));
  nor2  gate1449(.a(gate100inter5), .b(gate100inter2), .O(gate100inter6));
  inv1  gate1450(.a(G31), .O(gate100inter7));
  inv1  gate1451(.a(G353), .O(gate100inter8));
  nand2 gate1452(.a(gate100inter8), .b(gate100inter7), .O(gate100inter9));
  nand2 gate1453(.a(s_129), .b(gate100inter3), .O(gate100inter10));
  nor2  gate1454(.a(gate100inter10), .b(gate100inter9), .O(gate100inter11));
  nor2  gate1455(.a(gate100inter11), .b(gate100inter6), .O(gate100inter12));
  nand2 gate1456(.a(gate100inter12), .b(gate100inter1), .O(G421));
nand2 gate101( .a(G20), .b(G356), .O(G422) );
nand2 gate102( .a(G24), .b(G356), .O(G423) );

  xor2  gate2675(.a(G359), .b(G28), .O(gate103inter0));
  nand2 gate2676(.a(gate103inter0), .b(s_304), .O(gate103inter1));
  and2  gate2677(.a(G359), .b(G28), .O(gate103inter2));
  inv1  gate2678(.a(s_304), .O(gate103inter3));
  inv1  gate2679(.a(s_305), .O(gate103inter4));
  nand2 gate2680(.a(gate103inter4), .b(gate103inter3), .O(gate103inter5));
  nor2  gate2681(.a(gate103inter5), .b(gate103inter2), .O(gate103inter6));
  inv1  gate2682(.a(G28), .O(gate103inter7));
  inv1  gate2683(.a(G359), .O(gate103inter8));
  nand2 gate2684(.a(gate103inter8), .b(gate103inter7), .O(gate103inter9));
  nand2 gate2685(.a(s_305), .b(gate103inter3), .O(gate103inter10));
  nor2  gate2686(.a(gate103inter10), .b(gate103inter9), .O(gate103inter11));
  nor2  gate2687(.a(gate103inter11), .b(gate103inter6), .O(gate103inter12));
  nand2 gate2688(.a(gate103inter12), .b(gate103inter1), .O(G424));
nand2 gate104( .a(G32), .b(G359), .O(G425) );

  xor2  gate827(.a(G363), .b(G362), .O(gate105inter0));
  nand2 gate828(.a(gate105inter0), .b(s_40), .O(gate105inter1));
  and2  gate829(.a(G363), .b(G362), .O(gate105inter2));
  inv1  gate830(.a(s_40), .O(gate105inter3));
  inv1  gate831(.a(s_41), .O(gate105inter4));
  nand2 gate832(.a(gate105inter4), .b(gate105inter3), .O(gate105inter5));
  nor2  gate833(.a(gate105inter5), .b(gate105inter2), .O(gate105inter6));
  inv1  gate834(.a(G362), .O(gate105inter7));
  inv1  gate835(.a(G363), .O(gate105inter8));
  nand2 gate836(.a(gate105inter8), .b(gate105inter7), .O(gate105inter9));
  nand2 gate837(.a(s_41), .b(gate105inter3), .O(gate105inter10));
  nor2  gate838(.a(gate105inter10), .b(gate105inter9), .O(gate105inter11));
  nor2  gate839(.a(gate105inter11), .b(gate105inter6), .O(gate105inter12));
  nand2 gate840(.a(gate105inter12), .b(gate105inter1), .O(G426));

  xor2  gate2885(.a(G365), .b(G364), .O(gate106inter0));
  nand2 gate2886(.a(gate106inter0), .b(s_334), .O(gate106inter1));
  and2  gate2887(.a(G365), .b(G364), .O(gate106inter2));
  inv1  gate2888(.a(s_334), .O(gate106inter3));
  inv1  gate2889(.a(s_335), .O(gate106inter4));
  nand2 gate2890(.a(gate106inter4), .b(gate106inter3), .O(gate106inter5));
  nor2  gate2891(.a(gate106inter5), .b(gate106inter2), .O(gate106inter6));
  inv1  gate2892(.a(G364), .O(gate106inter7));
  inv1  gate2893(.a(G365), .O(gate106inter8));
  nand2 gate2894(.a(gate106inter8), .b(gate106inter7), .O(gate106inter9));
  nand2 gate2895(.a(s_335), .b(gate106inter3), .O(gate106inter10));
  nor2  gate2896(.a(gate106inter10), .b(gate106inter9), .O(gate106inter11));
  nor2  gate2897(.a(gate106inter11), .b(gate106inter6), .O(gate106inter12));
  nand2 gate2898(.a(gate106inter12), .b(gate106inter1), .O(G429));
nand2 gate107( .a(G366), .b(G367), .O(G432) );
nand2 gate108( .a(G368), .b(G369), .O(G435) );
nand2 gate109( .a(G370), .b(G371), .O(G438) );

  xor2  gate855(.a(G373), .b(G372), .O(gate110inter0));
  nand2 gate856(.a(gate110inter0), .b(s_44), .O(gate110inter1));
  and2  gate857(.a(G373), .b(G372), .O(gate110inter2));
  inv1  gate858(.a(s_44), .O(gate110inter3));
  inv1  gate859(.a(s_45), .O(gate110inter4));
  nand2 gate860(.a(gate110inter4), .b(gate110inter3), .O(gate110inter5));
  nor2  gate861(.a(gate110inter5), .b(gate110inter2), .O(gate110inter6));
  inv1  gate862(.a(G372), .O(gate110inter7));
  inv1  gate863(.a(G373), .O(gate110inter8));
  nand2 gate864(.a(gate110inter8), .b(gate110inter7), .O(gate110inter9));
  nand2 gate865(.a(s_45), .b(gate110inter3), .O(gate110inter10));
  nor2  gate866(.a(gate110inter10), .b(gate110inter9), .O(gate110inter11));
  nor2  gate867(.a(gate110inter11), .b(gate110inter6), .O(gate110inter12));
  nand2 gate868(.a(gate110inter12), .b(gate110inter1), .O(G441));

  xor2  gate1541(.a(G375), .b(G374), .O(gate111inter0));
  nand2 gate1542(.a(gate111inter0), .b(s_142), .O(gate111inter1));
  and2  gate1543(.a(G375), .b(G374), .O(gate111inter2));
  inv1  gate1544(.a(s_142), .O(gate111inter3));
  inv1  gate1545(.a(s_143), .O(gate111inter4));
  nand2 gate1546(.a(gate111inter4), .b(gate111inter3), .O(gate111inter5));
  nor2  gate1547(.a(gate111inter5), .b(gate111inter2), .O(gate111inter6));
  inv1  gate1548(.a(G374), .O(gate111inter7));
  inv1  gate1549(.a(G375), .O(gate111inter8));
  nand2 gate1550(.a(gate111inter8), .b(gate111inter7), .O(gate111inter9));
  nand2 gate1551(.a(s_143), .b(gate111inter3), .O(gate111inter10));
  nor2  gate1552(.a(gate111inter10), .b(gate111inter9), .O(gate111inter11));
  nor2  gate1553(.a(gate111inter11), .b(gate111inter6), .O(gate111inter12));
  nand2 gate1554(.a(gate111inter12), .b(gate111inter1), .O(G444));
nand2 gate112( .a(G376), .b(G377), .O(G447) );

  xor2  gate2521(.a(G379), .b(G378), .O(gate113inter0));
  nand2 gate2522(.a(gate113inter0), .b(s_282), .O(gate113inter1));
  and2  gate2523(.a(G379), .b(G378), .O(gate113inter2));
  inv1  gate2524(.a(s_282), .O(gate113inter3));
  inv1  gate2525(.a(s_283), .O(gate113inter4));
  nand2 gate2526(.a(gate113inter4), .b(gate113inter3), .O(gate113inter5));
  nor2  gate2527(.a(gate113inter5), .b(gate113inter2), .O(gate113inter6));
  inv1  gate2528(.a(G378), .O(gate113inter7));
  inv1  gate2529(.a(G379), .O(gate113inter8));
  nand2 gate2530(.a(gate113inter8), .b(gate113inter7), .O(gate113inter9));
  nand2 gate2531(.a(s_283), .b(gate113inter3), .O(gate113inter10));
  nor2  gate2532(.a(gate113inter10), .b(gate113inter9), .O(gate113inter11));
  nor2  gate2533(.a(gate113inter11), .b(gate113inter6), .O(gate113inter12));
  nand2 gate2534(.a(gate113inter12), .b(gate113inter1), .O(G450));
nand2 gate114( .a(G380), .b(G381), .O(G453) );

  xor2  gate2283(.a(G383), .b(G382), .O(gate115inter0));
  nand2 gate2284(.a(gate115inter0), .b(s_248), .O(gate115inter1));
  and2  gate2285(.a(G383), .b(G382), .O(gate115inter2));
  inv1  gate2286(.a(s_248), .O(gate115inter3));
  inv1  gate2287(.a(s_249), .O(gate115inter4));
  nand2 gate2288(.a(gate115inter4), .b(gate115inter3), .O(gate115inter5));
  nor2  gate2289(.a(gate115inter5), .b(gate115inter2), .O(gate115inter6));
  inv1  gate2290(.a(G382), .O(gate115inter7));
  inv1  gate2291(.a(G383), .O(gate115inter8));
  nand2 gate2292(.a(gate115inter8), .b(gate115inter7), .O(gate115inter9));
  nand2 gate2293(.a(s_249), .b(gate115inter3), .O(gate115inter10));
  nor2  gate2294(.a(gate115inter10), .b(gate115inter9), .O(gate115inter11));
  nor2  gate2295(.a(gate115inter11), .b(gate115inter6), .O(gate115inter12));
  nand2 gate2296(.a(gate115inter12), .b(gate115inter1), .O(G456));

  xor2  gate2157(.a(G385), .b(G384), .O(gate116inter0));
  nand2 gate2158(.a(gate116inter0), .b(s_230), .O(gate116inter1));
  and2  gate2159(.a(G385), .b(G384), .O(gate116inter2));
  inv1  gate2160(.a(s_230), .O(gate116inter3));
  inv1  gate2161(.a(s_231), .O(gate116inter4));
  nand2 gate2162(.a(gate116inter4), .b(gate116inter3), .O(gate116inter5));
  nor2  gate2163(.a(gate116inter5), .b(gate116inter2), .O(gate116inter6));
  inv1  gate2164(.a(G384), .O(gate116inter7));
  inv1  gate2165(.a(G385), .O(gate116inter8));
  nand2 gate2166(.a(gate116inter8), .b(gate116inter7), .O(gate116inter9));
  nand2 gate2167(.a(s_231), .b(gate116inter3), .O(gate116inter10));
  nor2  gate2168(.a(gate116inter10), .b(gate116inter9), .O(gate116inter11));
  nor2  gate2169(.a(gate116inter11), .b(gate116inter6), .O(gate116inter12));
  nand2 gate2170(.a(gate116inter12), .b(gate116inter1), .O(G459));
nand2 gate117( .a(G386), .b(G387), .O(G462) );
nand2 gate118( .a(G388), .b(G389), .O(G465) );
nand2 gate119( .a(G390), .b(G391), .O(G468) );

  xor2  gate1485(.a(G393), .b(G392), .O(gate120inter0));
  nand2 gate1486(.a(gate120inter0), .b(s_134), .O(gate120inter1));
  and2  gate1487(.a(G393), .b(G392), .O(gate120inter2));
  inv1  gate1488(.a(s_134), .O(gate120inter3));
  inv1  gate1489(.a(s_135), .O(gate120inter4));
  nand2 gate1490(.a(gate120inter4), .b(gate120inter3), .O(gate120inter5));
  nor2  gate1491(.a(gate120inter5), .b(gate120inter2), .O(gate120inter6));
  inv1  gate1492(.a(G392), .O(gate120inter7));
  inv1  gate1493(.a(G393), .O(gate120inter8));
  nand2 gate1494(.a(gate120inter8), .b(gate120inter7), .O(gate120inter9));
  nand2 gate1495(.a(s_135), .b(gate120inter3), .O(gate120inter10));
  nor2  gate1496(.a(gate120inter10), .b(gate120inter9), .O(gate120inter11));
  nor2  gate1497(.a(gate120inter11), .b(gate120inter6), .O(gate120inter12));
  nand2 gate1498(.a(gate120inter12), .b(gate120inter1), .O(G471));

  xor2  gate1835(.a(G395), .b(G394), .O(gate121inter0));
  nand2 gate1836(.a(gate121inter0), .b(s_184), .O(gate121inter1));
  and2  gate1837(.a(G395), .b(G394), .O(gate121inter2));
  inv1  gate1838(.a(s_184), .O(gate121inter3));
  inv1  gate1839(.a(s_185), .O(gate121inter4));
  nand2 gate1840(.a(gate121inter4), .b(gate121inter3), .O(gate121inter5));
  nor2  gate1841(.a(gate121inter5), .b(gate121inter2), .O(gate121inter6));
  inv1  gate1842(.a(G394), .O(gate121inter7));
  inv1  gate1843(.a(G395), .O(gate121inter8));
  nand2 gate1844(.a(gate121inter8), .b(gate121inter7), .O(gate121inter9));
  nand2 gate1845(.a(s_185), .b(gate121inter3), .O(gate121inter10));
  nor2  gate1846(.a(gate121inter10), .b(gate121inter9), .O(gate121inter11));
  nor2  gate1847(.a(gate121inter11), .b(gate121inter6), .O(gate121inter12));
  nand2 gate1848(.a(gate121inter12), .b(gate121inter1), .O(G474));
nand2 gate122( .a(G396), .b(G397), .O(G477) );

  xor2  gate1919(.a(G399), .b(G398), .O(gate123inter0));
  nand2 gate1920(.a(gate123inter0), .b(s_196), .O(gate123inter1));
  and2  gate1921(.a(G399), .b(G398), .O(gate123inter2));
  inv1  gate1922(.a(s_196), .O(gate123inter3));
  inv1  gate1923(.a(s_197), .O(gate123inter4));
  nand2 gate1924(.a(gate123inter4), .b(gate123inter3), .O(gate123inter5));
  nor2  gate1925(.a(gate123inter5), .b(gate123inter2), .O(gate123inter6));
  inv1  gate1926(.a(G398), .O(gate123inter7));
  inv1  gate1927(.a(G399), .O(gate123inter8));
  nand2 gate1928(.a(gate123inter8), .b(gate123inter7), .O(gate123inter9));
  nand2 gate1929(.a(s_197), .b(gate123inter3), .O(gate123inter10));
  nor2  gate1930(.a(gate123inter10), .b(gate123inter9), .O(gate123inter11));
  nor2  gate1931(.a(gate123inter11), .b(gate123inter6), .O(gate123inter12));
  nand2 gate1932(.a(gate123inter12), .b(gate123inter1), .O(G480));
nand2 gate124( .a(G400), .b(G401), .O(G483) );
nand2 gate125( .a(G402), .b(G403), .O(G486) );
nand2 gate126( .a(G404), .b(G405), .O(G489) );
nand2 gate127( .a(G406), .b(G407), .O(G492) );
nand2 gate128( .a(G408), .b(G409), .O(G495) );

  xor2  gate603(.a(G411), .b(G410), .O(gate129inter0));
  nand2 gate604(.a(gate129inter0), .b(s_8), .O(gate129inter1));
  and2  gate605(.a(G411), .b(G410), .O(gate129inter2));
  inv1  gate606(.a(s_8), .O(gate129inter3));
  inv1  gate607(.a(s_9), .O(gate129inter4));
  nand2 gate608(.a(gate129inter4), .b(gate129inter3), .O(gate129inter5));
  nor2  gate609(.a(gate129inter5), .b(gate129inter2), .O(gate129inter6));
  inv1  gate610(.a(G410), .O(gate129inter7));
  inv1  gate611(.a(G411), .O(gate129inter8));
  nand2 gate612(.a(gate129inter8), .b(gate129inter7), .O(gate129inter9));
  nand2 gate613(.a(s_9), .b(gate129inter3), .O(gate129inter10));
  nor2  gate614(.a(gate129inter10), .b(gate129inter9), .O(gate129inter11));
  nor2  gate615(.a(gate129inter11), .b(gate129inter6), .O(gate129inter12));
  nand2 gate616(.a(gate129inter12), .b(gate129inter1), .O(G498));
nand2 gate130( .a(G412), .b(G413), .O(G501) );
nand2 gate131( .a(G414), .b(G415), .O(G504) );

  xor2  gate1905(.a(G417), .b(G416), .O(gate132inter0));
  nand2 gate1906(.a(gate132inter0), .b(s_194), .O(gate132inter1));
  and2  gate1907(.a(G417), .b(G416), .O(gate132inter2));
  inv1  gate1908(.a(s_194), .O(gate132inter3));
  inv1  gate1909(.a(s_195), .O(gate132inter4));
  nand2 gate1910(.a(gate132inter4), .b(gate132inter3), .O(gate132inter5));
  nor2  gate1911(.a(gate132inter5), .b(gate132inter2), .O(gate132inter6));
  inv1  gate1912(.a(G416), .O(gate132inter7));
  inv1  gate1913(.a(G417), .O(gate132inter8));
  nand2 gate1914(.a(gate132inter8), .b(gate132inter7), .O(gate132inter9));
  nand2 gate1915(.a(s_195), .b(gate132inter3), .O(gate132inter10));
  nor2  gate1916(.a(gate132inter10), .b(gate132inter9), .O(gate132inter11));
  nor2  gate1917(.a(gate132inter11), .b(gate132inter6), .O(gate132inter12));
  nand2 gate1918(.a(gate132inter12), .b(gate132inter1), .O(G507));

  xor2  gate2689(.a(G419), .b(G418), .O(gate133inter0));
  nand2 gate2690(.a(gate133inter0), .b(s_306), .O(gate133inter1));
  and2  gate2691(.a(G419), .b(G418), .O(gate133inter2));
  inv1  gate2692(.a(s_306), .O(gate133inter3));
  inv1  gate2693(.a(s_307), .O(gate133inter4));
  nand2 gate2694(.a(gate133inter4), .b(gate133inter3), .O(gate133inter5));
  nor2  gate2695(.a(gate133inter5), .b(gate133inter2), .O(gate133inter6));
  inv1  gate2696(.a(G418), .O(gate133inter7));
  inv1  gate2697(.a(G419), .O(gate133inter8));
  nand2 gate2698(.a(gate133inter8), .b(gate133inter7), .O(gate133inter9));
  nand2 gate2699(.a(s_307), .b(gate133inter3), .O(gate133inter10));
  nor2  gate2700(.a(gate133inter10), .b(gate133inter9), .O(gate133inter11));
  nor2  gate2701(.a(gate133inter11), .b(gate133inter6), .O(gate133inter12));
  nand2 gate2702(.a(gate133inter12), .b(gate133inter1), .O(G510));

  xor2  gate547(.a(G421), .b(G420), .O(gate134inter0));
  nand2 gate548(.a(gate134inter0), .b(s_0), .O(gate134inter1));
  and2  gate549(.a(G421), .b(G420), .O(gate134inter2));
  inv1  gate550(.a(s_0), .O(gate134inter3));
  inv1  gate551(.a(s_1), .O(gate134inter4));
  nand2 gate552(.a(gate134inter4), .b(gate134inter3), .O(gate134inter5));
  nor2  gate553(.a(gate134inter5), .b(gate134inter2), .O(gate134inter6));
  inv1  gate554(.a(G420), .O(gate134inter7));
  inv1  gate555(.a(G421), .O(gate134inter8));
  nand2 gate556(.a(gate134inter8), .b(gate134inter7), .O(gate134inter9));
  nand2 gate557(.a(s_1), .b(gate134inter3), .O(gate134inter10));
  nor2  gate558(.a(gate134inter10), .b(gate134inter9), .O(gate134inter11));
  nor2  gate559(.a(gate134inter11), .b(gate134inter6), .O(gate134inter12));
  nand2 gate560(.a(gate134inter12), .b(gate134inter1), .O(G513));
nand2 gate135( .a(G422), .b(G423), .O(G516) );
nand2 gate136( .a(G424), .b(G425), .O(G519) );
nand2 gate137( .a(G426), .b(G429), .O(G522) );
nand2 gate138( .a(G432), .b(G435), .O(G525) );
nand2 gate139( .a(G438), .b(G441), .O(G528) );
nand2 gate140( .a(G444), .b(G447), .O(G531) );

  xor2  gate2297(.a(G453), .b(G450), .O(gate141inter0));
  nand2 gate2298(.a(gate141inter0), .b(s_250), .O(gate141inter1));
  and2  gate2299(.a(G453), .b(G450), .O(gate141inter2));
  inv1  gate2300(.a(s_250), .O(gate141inter3));
  inv1  gate2301(.a(s_251), .O(gate141inter4));
  nand2 gate2302(.a(gate141inter4), .b(gate141inter3), .O(gate141inter5));
  nor2  gate2303(.a(gate141inter5), .b(gate141inter2), .O(gate141inter6));
  inv1  gate2304(.a(G450), .O(gate141inter7));
  inv1  gate2305(.a(G453), .O(gate141inter8));
  nand2 gate2306(.a(gate141inter8), .b(gate141inter7), .O(gate141inter9));
  nand2 gate2307(.a(s_251), .b(gate141inter3), .O(gate141inter10));
  nor2  gate2308(.a(gate141inter10), .b(gate141inter9), .O(gate141inter11));
  nor2  gate2309(.a(gate141inter11), .b(gate141inter6), .O(gate141inter12));
  nand2 gate2310(.a(gate141inter12), .b(gate141inter1), .O(G534));

  xor2  gate1107(.a(G459), .b(G456), .O(gate142inter0));
  nand2 gate1108(.a(gate142inter0), .b(s_80), .O(gate142inter1));
  and2  gate1109(.a(G459), .b(G456), .O(gate142inter2));
  inv1  gate1110(.a(s_80), .O(gate142inter3));
  inv1  gate1111(.a(s_81), .O(gate142inter4));
  nand2 gate1112(.a(gate142inter4), .b(gate142inter3), .O(gate142inter5));
  nor2  gate1113(.a(gate142inter5), .b(gate142inter2), .O(gate142inter6));
  inv1  gate1114(.a(G456), .O(gate142inter7));
  inv1  gate1115(.a(G459), .O(gate142inter8));
  nand2 gate1116(.a(gate142inter8), .b(gate142inter7), .O(gate142inter9));
  nand2 gate1117(.a(s_81), .b(gate142inter3), .O(gate142inter10));
  nor2  gate1118(.a(gate142inter10), .b(gate142inter9), .O(gate142inter11));
  nor2  gate1119(.a(gate142inter11), .b(gate142inter6), .O(gate142inter12));
  nand2 gate1120(.a(gate142inter12), .b(gate142inter1), .O(G537));
nand2 gate143( .a(G462), .b(G465), .O(G540) );
nand2 gate144( .a(G468), .b(G471), .O(G543) );
nand2 gate145( .a(G474), .b(G477), .O(G546) );
nand2 gate146( .a(G480), .b(G483), .O(G549) );
nand2 gate147( .a(G486), .b(G489), .O(G552) );

  xor2  gate1653(.a(G495), .b(G492), .O(gate148inter0));
  nand2 gate1654(.a(gate148inter0), .b(s_158), .O(gate148inter1));
  and2  gate1655(.a(G495), .b(G492), .O(gate148inter2));
  inv1  gate1656(.a(s_158), .O(gate148inter3));
  inv1  gate1657(.a(s_159), .O(gate148inter4));
  nand2 gate1658(.a(gate148inter4), .b(gate148inter3), .O(gate148inter5));
  nor2  gate1659(.a(gate148inter5), .b(gate148inter2), .O(gate148inter6));
  inv1  gate1660(.a(G492), .O(gate148inter7));
  inv1  gate1661(.a(G495), .O(gate148inter8));
  nand2 gate1662(.a(gate148inter8), .b(gate148inter7), .O(gate148inter9));
  nand2 gate1663(.a(s_159), .b(gate148inter3), .O(gate148inter10));
  nor2  gate1664(.a(gate148inter10), .b(gate148inter9), .O(gate148inter11));
  nor2  gate1665(.a(gate148inter11), .b(gate148inter6), .O(gate148inter12));
  nand2 gate1666(.a(gate148inter12), .b(gate148inter1), .O(G555));

  xor2  gate1387(.a(G501), .b(G498), .O(gate149inter0));
  nand2 gate1388(.a(gate149inter0), .b(s_120), .O(gate149inter1));
  and2  gate1389(.a(G501), .b(G498), .O(gate149inter2));
  inv1  gate1390(.a(s_120), .O(gate149inter3));
  inv1  gate1391(.a(s_121), .O(gate149inter4));
  nand2 gate1392(.a(gate149inter4), .b(gate149inter3), .O(gate149inter5));
  nor2  gate1393(.a(gate149inter5), .b(gate149inter2), .O(gate149inter6));
  inv1  gate1394(.a(G498), .O(gate149inter7));
  inv1  gate1395(.a(G501), .O(gate149inter8));
  nand2 gate1396(.a(gate149inter8), .b(gate149inter7), .O(gate149inter9));
  nand2 gate1397(.a(s_121), .b(gate149inter3), .O(gate149inter10));
  nor2  gate1398(.a(gate149inter10), .b(gate149inter9), .O(gate149inter11));
  nor2  gate1399(.a(gate149inter11), .b(gate149inter6), .O(gate149inter12));
  nand2 gate1400(.a(gate149inter12), .b(gate149inter1), .O(G558));

  xor2  gate2395(.a(G507), .b(G504), .O(gate150inter0));
  nand2 gate2396(.a(gate150inter0), .b(s_264), .O(gate150inter1));
  and2  gate2397(.a(G507), .b(G504), .O(gate150inter2));
  inv1  gate2398(.a(s_264), .O(gate150inter3));
  inv1  gate2399(.a(s_265), .O(gate150inter4));
  nand2 gate2400(.a(gate150inter4), .b(gate150inter3), .O(gate150inter5));
  nor2  gate2401(.a(gate150inter5), .b(gate150inter2), .O(gate150inter6));
  inv1  gate2402(.a(G504), .O(gate150inter7));
  inv1  gate2403(.a(G507), .O(gate150inter8));
  nand2 gate2404(.a(gate150inter8), .b(gate150inter7), .O(gate150inter9));
  nand2 gate2405(.a(s_265), .b(gate150inter3), .O(gate150inter10));
  nor2  gate2406(.a(gate150inter10), .b(gate150inter9), .O(gate150inter11));
  nor2  gate2407(.a(gate150inter11), .b(gate150inter6), .O(gate150inter12));
  nand2 gate2408(.a(gate150inter12), .b(gate150inter1), .O(G561));
nand2 gate151( .a(G510), .b(G513), .O(G564) );
nand2 gate152( .a(G516), .b(G519), .O(G567) );

  xor2  gate1009(.a(G522), .b(G426), .O(gate153inter0));
  nand2 gate1010(.a(gate153inter0), .b(s_66), .O(gate153inter1));
  and2  gate1011(.a(G522), .b(G426), .O(gate153inter2));
  inv1  gate1012(.a(s_66), .O(gate153inter3));
  inv1  gate1013(.a(s_67), .O(gate153inter4));
  nand2 gate1014(.a(gate153inter4), .b(gate153inter3), .O(gate153inter5));
  nor2  gate1015(.a(gate153inter5), .b(gate153inter2), .O(gate153inter6));
  inv1  gate1016(.a(G426), .O(gate153inter7));
  inv1  gate1017(.a(G522), .O(gate153inter8));
  nand2 gate1018(.a(gate153inter8), .b(gate153inter7), .O(gate153inter9));
  nand2 gate1019(.a(s_67), .b(gate153inter3), .O(gate153inter10));
  nor2  gate1020(.a(gate153inter10), .b(gate153inter9), .O(gate153inter11));
  nor2  gate1021(.a(gate153inter11), .b(gate153inter6), .O(gate153inter12));
  nand2 gate1022(.a(gate153inter12), .b(gate153inter1), .O(G570));
nand2 gate154( .a(G429), .b(G522), .O(G571) );
nand2 gate155( .a(G432), .b(G525), .O(G572) );
nand2 gate156( .a(G435), .b(G525), .O(G573) );

  xor2  gate883(.a(G528), .b(G438), .O(gate157inter0));
  nand2 gate884(.a(gate157inter0), .b(s_48), .O(gate157inter1));
  and2  gate885(.a(G528), .b(G438), .O(gate157inter2));
  inv1  gate886(.a(s_48), .O(gate157inter3));
  inv1  gate887(.a(s_49), .O(gate157inter4));
  nand2 gate888(.a(gate157inter4), .b(gate157inter3), .O(gate157inter5));
  nor2  gate889(.a(gate157inter5), .b(gate157inter2), .O(gate157inter6));
  inv1  gate890(.a(G438), .O(gate157inter7));
  inv1  gate891(.a(G528), .O(gate157inter8));
  nand2 gate892(.a(gate157inter8), .b(gate157inter7), .O(gate157inter9));
  nand2 gate893(.a(s_49), .b(gate157inter3), .O(gate157inter10));
  nor2  gate894(.a(gate157inter10), .b(gate157inter9), .O(gate157inter11));
  nor2  gate895(.a(gate157inter11), .b(gate157inter6), .O(gate157inter12));
  nand2 gate896(.a(gate157inter12), .b(gate157inter1), .O(G574));
nand2 gate158( .a(G441), .b(G528), .O(G575) );
nand2 gate159( .a(G444), .b(G531), .O(G576) );

  xor2  gate1723(.a(G531), .b(G447), .O(gate160inter0));
  nand2 gate1724(.a(gate160inter0), .b(s_168), .O(gate160inter1));
  and2  gate1725(.a(G531), .b(G447), .O(gate160inter2));
  inv1  gate1726(.a(s_168), .O(gate160inter3));
  inv1  gate1727(.a(s_169), .O(gate160inter4));
  nand2 gate1728(.a(gate160inter4), .b(gate160inter3), .O(gate160inter5));
  nor2  gate1729(.a(gate160inter5), .b(gate160inter2), .O(gate160inter6));
  inv1  gate1730(.a(G447), .O(gate160inter7));
  inv1  gate1731(.a(G531), .O(gate160inter8));
  nand2 gate1732(.a(gate160inter8), .b(gate160inter7), .O(gate160inter9));
  nand2 gate1733(.a(s_169), .b(gate160inter3), .O(gate160inter10));
  nor2  gate1734(.a(gate160inter10), .b(gate160inter9), .O(gate160inter11));
  nor2  gate1735(.a(gate160inter11), .b(gate160inter6), .O(gate160inter12));
  nand2 gate1736(.a(gate160inter12), .b(gate160inter1), .O(G577));

  xor2  gate687(.a(G534), .b(G450), .O(gate161inter0));
  nand2 gate688(.a(gate161inter0), .b(s_20), .O(gate161inter1));
  and2  gate689(.a(G534), .b(G450), .O(gate161inter2));
  inv1  gate690(.a(s_20), .O(gate161inter3));
  inv1  gate691(.a(s_21), .O(gate161inter4));
  nand2 gate692(.a(gate161inter4), .b(gate161inter3), .O(gate161inter5));
  nor2  gate693(.a(gate161inter5), .b(gate161inter2), .O(gate161inter6));
  inv1  gate694(.a(G450), .O(gate161inter7));
  inv1  gate695(.a(G534), .O(gate161inter8));
  nand2 gate696(.a(gate161inter8), .b(gate161inter7), .O(gate161inter9));
  nand2 gate697(.a(s_21), .b(gate161inter3), .O(gate161inter10));
  nor2  gate698(.a(gate161inter10), .b(gate161inter9), .O(gate161inter11));
  nor2  gate699(.a(gate161inter11), .b(gate161inter6), .O(gate161inter12));
  nand2 gate700(.a(gate161inter12), .b(gate161inter1), .O(G578));
nand2 gate162( .a(G453), .b(G534), .O(G579) );
nand2 gate163( .a(G456), .b(G537), .O(G580) );

  xor2  gate2073(.a(G537), .b(G459), .O(gate164inter0));
  nand2 gate2074(.a(gate164inter0), .b(s_218), .O(gate164inter1));
  and2  gate2075(.a(G537), .b(G459), .O(gate164inter2));
  inv1  gate2076(.a(s_218), .O(gate164inter3));
  inv1  gate2077(.a(s_219), .O(gate164inter4));
  nand2 gate2078(.a(gate164inter4), .b(gate164inter3), .O(gate164inter5));
  nor2  gate2079(.a(gate164inter5), .b(gate164inter2), .O(gate164inter6));
  inv1  gate2080(.a(G459), .O(gate164inter7));
  inv1  gate2081(.a(G537), .O(gate164inter8));
  nand2 gate2082(.a(gate164inter8), .b(gate164inter7), .O(gate164inter9));
  nand2 gate2083(.a(s_219), .b(gate164inter3), .O(gate164inter10));
  nor2  gate2084(.a(gate164inter10), .b(gate164inter9), .O(gate164inter11));
  nor2  gate2085(.a(gate164inter11), .b(gate164inter6), .O(gate164inter12));
  nand2 gate2086(.a(gate164inter12), .b(gate164inter1), .O(G581));
nand2 gate165( .a(G462), .b(G540), .O(G582) );

  xor2  gate1415(.a(G540), .b(G465), .O(gate166inter0));
  nand2 gate1416(.a(gate166inter0), .b(s_124), .O(gate166inter1));
  and2  gate1417(.a(G540), .b(G465), .O(gate166inter2));
  inv1  gate1418(.a(s_124), .O(gate166inter3));
  inv1  gate1419(.a(s_125), .O(gate166inter4));
  nand2 gate1420(.a(gate166inter4), .b(gate166inter3), .O(gate166inter5));
  nor2  gate1421(.a(gate166inter5), .b(gate166inter2), .O(gate166inter6));
  inv1  gate1422(.a(G465), .O(gate166inter7));
  inv1  gate1423(.a(G540), .O(gate166inter8));
  nand2 gate1424(.a(gate166inter8), .b(gate166inter7), .O(gate166inter9));
  nand2 gate1425(.a(s_125), .b(gate166inter3), .O(gate166inter10));
  nor2  gate1426(.a(gate166inter10), .b(gate166inter9), .O(gate166inter11));
  nor2  gate1427(.a(gate166inter11), .b(gate166inter6), .O(gate166inter12));
  nand2 gate1428(.a(gate166inter12), .b(gate166inter1), .O(G583));
nand2 gate167( .a(G468), .b(G543), .O(G584) );

  xor2  gate729(.a(G543), .b(G471), .O(gate168inter0));
  nand2 gate730(.a(gate168inter0), .b(s_26), .O(gate168inter1));
  and2  gate731(.a(G543), .b(G471), .O(gate168inter2));
  inv1  gate732(.a(s_26), .O(gate168inter3));
  inv1  gate733(.a(s_27), .O(gate168inter4));
  nand2 gate734(.a(gate168inter4), .b(gate168inter3), .O(gate168inter5));
  nor2  gate735(.a(gate168inter5), .b(gate168inter2), .O(gate168inter6));
  inv1  gate736(.a(G471), .O(gate168inter7));
  inv1  gate737(.a(G543), .O(gate168inter8));
  nand2 gate738(.a(gate168inter8), .b(gate168inter7), .O(gate168inter9));
  nand2 gate739(.a(s_27), .b(gate168inter3), .O(gate168inter10));
  nor2  gate740(.a(gate168inter10), .b(gate168inter9), .O(gate168inter11));
  nor2  gate741(.a(gate168inter11), .b(gate168inter6), .O(gate168inter12));
  nand2 gate742(.a(gate168inter12), .b(gate168inter1), .O(G585));

  xor2  gate2661(.a(G546), .b(G474), .O(gate169inter0));
  nand2 gate2662(.a(gate169inter0), .b(s_302), .O(gate169inter1));
  and2  gate2663(.a(G546), .b(G474), .O(gate169inter2));
  inv1  gate2664(.a(s_302), .O(gate169inter3));
  inv1  gate2665(.a(s_303), .O(gate169inter4));
  nand2 gate2666(.a(gate169inter4), .b(gate169inter3), .O(gate169inter5));
  nor2  gate2667(.a(gate169inter5), .b(gate169inter2), .O(gate169inter6));
  inv1  gate2668(.a(G474), .O(gate169inter7));
  inv1  gate2669(.a(G546), .O(gate169inter8));
  nand2 gate2670(.a(gate169inter8), .b(gate169inter7), .O(gate169inter9));
  nand2 gate2671(.a(s_303), .b(gate169inter3), .O(gate169inter10));
  nor2  gate2672(.a(gate169inter10), .b(gate169inter9), .O(gate169inter11));
  nor2  gate2673(.a(gate169inter11), .b(gate169inter6), .O(gate169inter12));
  nand2 gate2674(.a(gate169inter12), .b(gate169inter1), .O(G586));

  xor2  gate2185(.a(G546), .b(G477), .O(gate170inter0));
  nand2 gate2186(.a(gate170inter0), .b(s_234), .O(gate170inter1));
  and2  gate2187(.a(G546), .b(G477), .O(gate170inter2));
  inv1  gate2188(.a(s_234), .O(gate170inter3));
  inv1  gate2189(.a(s_235), .O(gate170inter4));
  nand2 gate2190(.a(gate170inter4), .b(gate170inter3), .O(gate170inter5));
  nor2  gate2191(.a(gate170inter5), .b(gate170inter2), .O(gate170inter6));
  inv1  gate2192(.a(G477), .O(gate170inter7));
  inv1  gate2193(.a(G546), .O(gate170inter8));
  nand2 gate2194(.a(gate170inter8), .b(gate170inter7), .O(gate170inter9));
  nand2 gate2195(.a(s_235), .b(gate170inter3), .O(gate170inter10));
  nor2  gate2196(.a(gate170inter10), .b(gate170inter9), .O(gate170inter11));
  nor2  gate2197(.a(gate170inter11), .b(gate170inter6), .O(gate170inter12));
  nand2 gate2198(.a(gate170inter12), .b(gate170inter1), .O(G587));

  xor2  gate2773(.a(G549), .b(G480), .O(gate171inter0));
  nand2 gate2774(.a(gate171inter0), .b(s_318), .O(gate171inter1));
  and2  gate2775(.a(G549), .b(G480), .O(gate171inter2));
  inv1  gate2776(.a(s_318), .O(gate171inter3));
  inv1  gate2777(.a(s_319), .O(gate171inter4));
  nand2 gate2778(.a(gate171inter4), .b(gate171inter3), .O(gate171inter5));
  nor2  gate2779(.a(gate171inter5), .b(gate171inter2), .O(gate171inter6));
  inv1  gate2780(.a(G480), .O(gate171inter7));
  inv1  gate2781(.a(G549), .O(gate171inter8));
  nand2 gate2782(.a(gate171inter8), .b(gate171inter7), .O(gate171inter9));
  nand2 gate2783(.a(s_319), .b(gate171inter3), .O(gate171inter10));
  nor2  gate2784(.a(gate171inter10), .b(gate171inter9), .O(gate171inter11));
  nor2  gate2785(.a(gate171inter11), .b(gate171inter6), .O(gate171inter12));
  nand2 gate2786(.a(gate171inter12), .b(gate171inter1), .O(G588));
nand2 gate172( .a(G483), .b(G549), .O(G589) );

  xor2  gate2647(.a(G552), .b(G486), .O(gate173inter0));
  nand2 gate2648(.a(gate173inter0), .b(s_300), .O(gate173inter1));
  and2  gate2649(.a(G552), .b(G486), .O(gate173inter2));
  inv1  gate2650(.a(s_300), .O(gate173inter3));
  inv1  gate2651(.a(s_301), .O(gate173inter4));
  nand2 gate2652(.a(gate173inter4), .b(gate173inter3), .O(gate173inter5));
  nor2  gate2653(.a(gate173inter5), .b(gate173inter2), .O(gate173inter6));
  inv1  gate2654(.a(G486), .O(gate173inter7));
  inv1  gate2655(.a(G552), .O(gate173inter8));
  nand2 gate2656(.a(gate173inter8), .b(gate173inter7), .O(gate173inter9));
  nand2 gate2657(.a(s_301), .b(gate173inter3), .O(gate173inter10));
  nor2  gate2658(.a(gate173inter10), .b(gate173inter9), .O(gate173inter11));
  nor2  gate2659(.a(gate173inter11), .b(gate173inter6), .O(gate173inter12));
  nand2 gate2660(.a(gate173inter12), .b(gate173inter1), .O(G590));

  xor2  gate1779(.a(G552), .b(G489), .O(gate174inter0));
  nand2 gate1780(.a(gate174inter0), .b(s_176), .O(gate174inter1));
  and2  gate1781(.a(G552), .b(G489), .O(gate174inter2));
  inv1  gate1782(.a(s_176), .O(gate174inter3));
  inv1  gate1783(.a(s_177), .O(gate174inter4));
  nand2 gate1784(.a(gate174inter4), .b(gate174inter3), .O(gate174inter5));
  nor2  gate1785(.a(gate174inter5), .b(gate174inter2), .O(gate174inter6));
  inv1  gate1786(.a(G489), .O(gate174inter7));
  inv1  gate1787(.a(G552), .O(gate174inter8));
  nand2 gate1788(.a(gate174inter8), .b(gate174inter7), .O(gate174inter9));
  nand2 gate1789(.a(s_177), .b(gate174inter3), .O(gate174inter10));
  nor2  gate1790(.a(gate174inter10), .b(gate174inter9), .O(gate174inter11));
  nor2  gate1791(.a(gate174inter11), .b(gate174inter6), .O(gate174inter12));
  nand2 gate1792(.a(gate174inter12), .b(gate174inter1), .O(G591));

  xor2  gate645(.a(G555), .b(G492), .O(gate175inter0));
  nand2 gate646(.a(gate175inter0), .b(s_14), .O(gate175inter1));
  and2  gate647(.a(G555), .b(G492), .O(gate175inter2));
  inv1  gate648(.a(s_14), .O(gate175inter3));
  inv1  gate649(.a(s_15), .O(gate175inter4));
  nand2 gate650(.a(gate175inter4), .b(gate175inter3), .O(gate175inter5));
  nor2  gate651(.a(gate175inter5), .b(gate175inter2), .O(gate175inter6));
  inv1  gate652(.a(G492), .O(gate175inter7));
  inv1  gate653(.a(G555), .O(gate175inter8));
  nand2 gate654(.a(gate175inter8), .b(gate175inter7), .O(gate175inter9));
  nand2 gate655(.a(s_15), .b(gate175inter3), .O(gate175inter10));
  nor2  gate656(.a(gate175inter10), .b(gate175inter9), .O(gate175inter11));
  nor2  gate657(.a(gate175inter11), .b(gate175inter6), .O(gate175inter12));
  nand2 gate658(.a(gate175inter12), .b(gate175inter1), .O(G592));
nand2 gate176( .a(G495), .b(G555), .O(G593) );
nand2 gate177( .a(G498), .b(G558), .O(G594) );
nand2 gate178( .a(G501), .b(G558), .O(G595) );
nand2 gate179( .a(G504), .b(G561), .O(G596) );

  xor2  gate897(.a(G561), .b(G507), .O(gate180inter0));
  nand2 gate898(.a(gate180inter0), .b(s_50), .O(gate180inter1));
  and2  gate899(.a(G561), .b(G507), .O(gate180inter2));
  inv1  gate900(.a(s_50), .O(gate180inter3));
  inv1  gate901(.a(s_51), .O(gate180inter4));
  nand2 gate902(.a(gate180inter4), .b(gate180inter3), .O(gate180inter5));
  nor2  gate903(.a(gate180inter5), .b(gate180inter2), .O(gate180inter6));
  inv1  gate904(.a(G507), .O(gate180inter7));
  inv1  gate905(.a(G561), .O(gate180inter8));
  nand2 gate906(.a(gate180inter8), .b(gate180inter7), .O(gate180inter9));
  nand2 gate907(.a(s_51), .b(gate180inter3), .O(gate180inter10));
  nor2  gate908(.a(gate180inter10), .b(gate180inter9), .O(gate180inter11));
  nor2  gate909(.a(gate180inter11), .b(gate180inter6), .O(gate180inter12));
  nand2 gate910(.a(gate180inter12), .b(gate180inter1), .O(G597));
nand2 gate181( .a(G510), .b(G564), .O(G598) );
nand2 gate182( .a(G513), .b(G564), .O(G599) );
nand2 gate183( .a(G516), .b(G567), .O(G600) );

  xor2  gate1625(.a(G567), .b(G519), .O(gate184inter0));
  nand2 gate1626(.a(gate184inter0), .b(s_154), .O(gate184inter1));
  and2  gate1627(.a(G567), .b(G519), .O(gate184inter2));
  inv1  gate1628(.a(s_154), .O(gate184inter3));
  inv1  gate1629(.a(s_155), .O(gate184inter4));
  nand2 gate1630(.a(gate184inter4), .b(gate184inter3), .O(gate184inter5));
  nor2  gate1631(.a(gate184inter5), .b(gate184inter2), .O(gate184inter6));
  inv1  gate1632(.a(G519), .O(gate184inter7));
  inv1  gate1633(.a(G567), .O(gate184inter8));
  nand2 gate1634(.a(gate184inter8), .b(gate184inter7), .O(gate184inter9));
  nand2 gate1635(.a(s_155), .b(gate184inter3), .O(gate184inter10));
  nor2  gate1636(.a(gate184inter10), .b(gate184inter9), .O(gate184inter11));
  nor2  gate1637(.a(gate184inter11), .b(gate184inter6), .O(gate184inter12));
  nand2 gate1638(.a(gate184inter12), .b(gate184inter1), .O(G601));
nand2 gate185( .a(G570), .b(G571), .O(G602) );
nand2 gate186( .a(G572), .b(G573), .O(G607) );
nand2 gate187( .a(G574), .b(G575), .O(G612) );
nand2 gate188( .a(G576), .b(G577), .O(G617) );
nand2 gate189( .a(G578), .b(G579), .O(G622) );
nand2 gate190( .a(G580), .b(G581), .O(G627) );

  xor2  gate2409(.a(G583), .b(G582), .O(gate191inter0));
  nand2 gate2410(.a(gate191inter0), .b(s_266), .O(gate191inter1));
  and2  gate2411(.a(G583), .b(G582), .O(gate191inter2));
  inv1  gate2412(.a(s_266), .O(gate191inter3));
  inv1  gate2413(.a(s_267), .O(gate191inter4));
  nand2 gate2414(.a(gate191inter4), .b(gate191inter3), .O(gate191inter5));
  nor2  gate2415(.a(gate191inter5), .b(gate191inter2), .O(gate191inter6));
  inv1  gate2416(.a(G582), .O(gate191inter7));
  inv1  gate2417(.a(G583), .O(gate191inter8));
  nand2 gate2418(.a(gate191inter8), .b(gate191inter7), .O(gate191inter9));
  nand2 gate2419(.a(s_267), .b(gate191inter3), .O(gate191inter10));
  nor2  gate2420(.a(gate191inter10), .b(gate191inter9), .O(gate191inter11));
  nor2  gate2421(.a(gate191inter11), .b(gate191inter6), .O(gate191inter12));
  nand2 gate2422(.a(gate191inter12), .b(gate191inter1), .O(G632));

  xor2  gate1275(.a(G585), .b(G584), .O(gate192inter0));
  nand2 gate1276(.a(gate192inter0), .b(s_104), .O(gate192inter1));
  and2  gate1277(.a(G585), .b(G584), .O(gate192inter2));
  inv1  gate1278(.a(s_104), .O(gate192inter3));
  inv1  gate1279(.a(s_105), .O(gate192inter4));
  nand2 gate1280(.a(gate192inter4), .b(gate192inter3), .O(gate192inter5));
  nor2  gate1281(.a(gate192inter5), .b(gate192inter2), .O(gate192inter6));
  inv1  gate1282(.a(G584), .O(gate192inter7));
  inv1  gate1283(.a(G585), .O(gate192inter8));
  nand2 gate1284(.a(gate192inter8), .b(gate192inter7), .O(gate192inter9));
  nand2 gate1285(.a(s_105), .b(gate192inter3), .O(gate192inter10));
  nor2  gate1286(.a(gate192inter10), .b(gate192inter9), .O(gate192inter11));
  nor2  gate1287(.a(gate192inter11), .b(gate192inter6), .O(gate192inter12));
  nand2 gate1288(.a(gate192inter12), .b(gate192inter1), .O(G637));

  xor2  gate1891(.a(G587), .b(G586), .O(gate193inter0));
  nand2 gate1892(.a(gate193inter0), .b(s_192), .O(gate193inter1));
  and2  gate1893(.a(G587), .b(G586), .O(gate193inter2));
  inv1  gate1894(.a(s_192), .O(gate193inter3));
  inv1  gate1895(.a(s_193), .O(gate193inter4));
  nand2 gate1896(.a(gate193inter4), .b(gate193inter3), .O(gate193inter5));
  nor2  gate1897(.a(gate193inter5), .b(gate193inter2), .O(gate193inter6));
  inv1  gate1898(.a(G586), .O(gate193inter7));
  inv1  gate1899(.a(G587), .O(gate193inter8));
  nand2 gate1900(.a(gate193inter8), .b(gate193inter7), .O(gate193inter9));
  nand2 gate1901(.a(s_193), .b(gate193inter3), .O(gate193inter10));
  nor2  gate1902(.a(gate193inter10), .b(gate193inter9), .O(gate193inter11));
  nor2  gate1903(.a(gate193inter11), .b(gate193inter6), .O(gate193inter12));
  nand2 gate1904(.a(gate193inter12), .b(gate193inter1), .O(G642));
nand2 gate194( .a(G588), .b(G589), .O(G645) );

  xor2  gate995(.a(G591), .b(G590), .O(gate195inter0));
  nand2 gate996(.a(gate195inter0), .b(s_64), .O(gate195inter1));
  and2  gate997(.a(G591), .b(G590), .O(gate195inter2));
  inv1  gate998(.a(s_64), .O(gate195inter3));
  inv1  gate999(.a(s_65), .O(gate195inter4));
  nand2 gate1000(.a(gate195inter4), .b(gate195inter3), .O(gate195inter5));
  nor2  gate1001(.a(gate195inter5), .b(gate195inter2), .O(gate195inter6));
  inv1  gate1002(.a(G590), .O(gate195inter7));
  inv1  gate1003(.a(G591), .O(gate195inter8));
  nand2 gate1004(.a(gate195inter8), .b(gate195inter7), .O(gate195inter9));
  nand2 gate1005(.a(s_65), .b(gate195inter3), .O(gate195inter10));
  nor2  gate1006(.a(gate195inter10), .b(gate195inter9), .O(gate195inter11));
  nor2  gate1007(.a(gate195inter11), .b(gate195inter6), .O(gate195inter12));
  nand2 gate1008(.a(gate195inter12), .b(gate195inter1), .O(G648));
nand2 gate196( .a(G592), .b(G593), .O(G651) );

  xor2  gate1639(.a(G595), .b(G594), .O(gate197inter0));
  nand2 gate1640(.a(gate197inter0), .b(s_156), .O(gate197inter1));
  and2  gate1641(.a(G595), .b(G594), .O(gate197inter2));
  inv1  gate1642(.a(s_156), .O(gate197inter3));
  inv1  gate1643(.a(s_157), .O(gate197inter4));
  nand2 gate1644(.a(gate197inter4), .b(gate197inter3), .O(gate197inter5));
  nor2  gate1645(.a(gate197inter5), .b(gate197inter2), .O(gate197inter6));
  inv1  gate1646(.a(G594), .O(gate197inter7));
  inv1  gate1647(.a(G595), .O(gate197inter8));
  nand2 gate1648(.a(gate197inter8), .b(gate197inter7), .O(gate197inter9));
  nand2 gate1649(.a(s_157), .b(gate197inter3), .O(gate197inter10));
  nor2  gate1650(.a(gate197inter10), .b(gate197inter9), .O(gate197inter11));
  nor2  gate1651(.a(gate197inter11), .b(gate197inter6), .O(gate197inter12));
  nand2 gate1652(.a(gate197inter12), .b(gate197inter1), .O(G654));
nand2 gate198( .a(G596), .b(G597), .O(G657) );
nand2 gate199( .a(G598), .b(G599), .O(G660) );

  xor2  gate2563(.a(G601), .b(G600), .O(gate200inter0));
  nand2 gate2564(.a(gate200inter0), .b(s_288), .O(gate200inter1));
  and2  gate2565(.a(G601), .b(G600), .O(gate200inter2));
  inv1  gate2566(.a(s_288), .O(gate200inter3));
  inv1  gate2567(.a(s_289), .O(gate200inter4));
  nand2 gate2568(.a(gate200inter4), .b(gate200inter3), .O(gate200inter5));
  nor2  gate2569(.a(gate200inter5), .b(gate200inter2), .O(gate200inter6));
  inv1  gate2570(.a(G600), .O(gate200inter7));
  inv1  gate2571(.a(G601), .O(gate200inter8));
  nand2 gate2572(.a(gate200inter8), .b(gate200inter7), .O(gate200inter9));
  nand2 gate2573(.a(s_289), .b(gate200inter3), .O(gate200inter10));
  nor2  gate2574(.a(gate200inter10), .b(gate200inter9), .O(gate200inter11));
  nor2  gate2575(.a(gate200inter11), .b(gate200inter6), .O(gate200inter12));
  nand2 gate2576(.a(gate200inter12), .b(gate200inter1), .O(G663));
nand2 gate201( .a(G602), .b(G607), .O(G666) );

  xor2  gate2129(.a(G617), .b(G612), .O(gate202inter0));
  nand2 gate2130(.a(gate202inter0), .b(s_226), .O(gate202inter1));
  and2  gate2131(.a(G617), .b(G612), .O(gate202inter2));
  inv1  gate2132(.a(s_226), .O(gate202inter3));
  inv1  gate2133(.a(s_227), .O(gate202inter4));
  nand2 gate2134(.a(gate202inter4), .b(gate202inter3), .O(gate202inter5));
  nor2  gate2135(.a(gate202inter5), .b(gate202inter2), .O(gate202inter6));
  inv1  gate2136(.a(G612), .O(gate202inter7));
  inv1  gate2137(.a(G617), .O(gate202inter8));
  nand2 gate2138(.a(gate202inter8), .b(gate202inter7), .O(gate202inter9));
  nand2 gate2139(.a(s_227), .b(gate202inter3), .O(gate202inter10));
  nor2  gate2140(.a(gate202inter10), .b(gate202inter9), .O(gate202inter11));
  nor2  gate2141(.a(gate202inter11), .b(gate202inter6), .O(gate202inter12));
  nand2 gate2142(.a(gate202inter12), .b(gate202inter1), .O(G669));
nand2 gate203( .a(G602), .b(G612), .O(G672) );
nand2 gate204( .a(G607), .b(G617), .O(G675) );

  xor2  gate2059(.a(G627), .b(G622), .O(gate205inter0));
  nand2 gate2060(.a(gate205inter0), .b(s_216), .O(gate205inter1));
  and2  gate2061(.a(G627), .b(G622), .O(gate205inter2));
  inv1  gate2062(.a(s_216), .O(gate205inter3));
  inv1  gate2063(.a(s_217), .O(gate205inter4));
  nand2 gate2064(.a(gate205inter4), .b(gate205inter3), .O(gate205inter5));
  nor2  gate2065(.a(gate205inter5), .b(gate205inter2), .O(gate205inter6));
  inv1  gate2066(.a(G622), .O(gate205inter7));
  inv1  gate2067(.a(G627), .O(gate205inter8));
  nand2 gate2068(.a(gate205inter8), .b(gate205inter7), .O(gate205inter9));
  nand2 gate2069(.a(s_217), .b(gate205inter3), .O(gate205inter10));
  nor2  gate2070(.a(gate205inter10), .b(gate205inter9), .O(gate205inter11));
  nor2  gate2071(.a(gate205inter11), .b(gate205inter6), .O(gate205inter12));
  nand2 gate2072(.a(gate205inter12), .b(gate205inter1), .O(G678));

  xor2  gate1695(.a(G637), .b(G632), .O(gate206inter0));
  nand2 gate1696(.a(gate206inter0), .b(s_164), .O(gate206inter1));
  and2  gate1697(.a(G637), .b(G632), .O(gate206inter2));
  inv1  gate1698(.a(s_164), .O(gate206inter3));
  inv1  gate1699(.a(s_165), .O(gate206inter4));
  nand2 gate1700(.a(gate206inter4), .b(gate206inter3), .O(gate206inter5));
  nor2  gate1701(.a(gate206inter5), .b(gate206inter2), .O(gate206inter6));
  inv1  gate1702(.a(G632), .O(gate206inter7));
  inv1  gate1703(.a(G637), .O(gate206inter8));
  nand2 gate1704(.a(gate206inter8), .b(gate206inter7), .O(gate206inter9));
  nand2 gate1705(.a(s_165), .b(gate206inter3), .O(gate206inter10));
  nor2  gate1706(.a(gate206inter10), .b(gate206inter9), .O(gate206inter11));
  nor2  gate1707(.a(gate206inter11), .b(gate206inter6), .O(gate206inter12));
  nand2 gate1708(.a(gate206inter12), .b(gate206inter1), .O(G681));

  xor2  gate1191(.a(G632), .b(G622), .O(gate207inter0));
  nand2 gate1192(.a(gate207inter0), .b(s_92), .O(gate207inter1));
  and2  gate1193(.a(G632), .b(G622), .O(gate207inter2));
  inv1  gate1194(.a(s_92), .O(gate207inter3));
  inv1  gate1195(.a(s_93), .O(gate207inter4));
  nand2 gate1196(.a(gate207inter4), .b(gate207inter3), .O(gate207inter5));
  nor2  gate1197(.a(gate207inter5), .b(gate207inter2), .O(gate207inter6));
  inv1  gate1198(.a(G622), .O(gate207inter7));
  inv1  gate1199(.a(G632), .O(gate207inter8));
  nand2 gate1200(.a(gate207inter8), .b(gate207inter7), .O(gate207inter9));
  nand2 gate1201(.a(s_93), .b(gate207inter3), .O(gate207inter10));
  nor2  gate1202(.a(gate207inter10), .b(gate207inter9), .O(gate207inter11));
  nor2  gate1203(.a(gate207inter11), .b(gate207inter6), .O(gate207inter12));
  nand2 gate1204(.a(gate207inter12), .b(gate207inter1), .O(G684));

  xor2  gate2507(.a(G637), .b(G627), .O(gate208inter0));
  nand2 gate2508(.a(gate208inter0), .b(s_280), .O(gate208inter1));
  and2  gate2509(.a(G637), .b(G627), .O(gate208inter2));
  inv1  gate2510(.a(s_280), .O(gate208inter3));
  inv1  gate2511(.a(s_281), .O(gate208inter4));
  nand2 gate2512(.a(gate208inter4), .b(gate208inter3), .O(gate208inter5));
  nor2  gate2513(.a(gate208inter5), .b(gate208inter2), .O(gate208inter6));
  inv1  gate2514(.a(G627), .O(gate208inter7));
  inv1  gate2515(.a(G637), .O(gate208inter8));
  nand2 gate2516(.a(gate208inter8), .b(gate208inter7), .O(gate208inter9));
  nand2 gate2517(.a(s_281), .b(gate208inter3), .O(gate208inter10));
  nor2  gate2518(.a(gate208inter10), .b(gate208inter9), .O(gate208inter11));
  nor2  gate2519(.a(gate208inter11), .b(gate208inter6), .O(gate208inter12));
  nand2 gate2520(.a(gate208inter12), .b(gate208inter1), .O(G687));
nand2 gate209( .a(G602), .b(G666), .O(G690) );

  xor2  gate2423(.a(G666), .b(G607), .O(gate210inter0));
  nand2 gate2424(.a(gate210inter0), .b(s_268), .O(gate210inter1));
  and2  gate2425(.a(G666), .b(G607), .O(gate210inter2));
  inv1  gate2426(.a(s_268), .O(gate210inter3));
  inv1  gate2427(.a(s_269), .O(gate210inter4));
  nand2 gate2428(.a(gate210inter4), .b(gate210inter3), .O(gate210inter5));
  nor2  gate2429(.a(gate210inter5), .b(gate210inter2), .O(gate210inter6));
  inv1  gate2430(.a(G607), .O(gate210inter7));
  inv1  gate2431(.a(G666), .O(gate210inter8));
  nand2 gate2432(.a(gate210inter8), .b(gate210inter7), .O(gate210inter9));
  nand2 gate2433(.a(s_269), .b(gate210inter3), .O(gate210inter10));
  nor2  gate2434(.a(gate210inter10), .b(gate210inter9), .O(gate210inter11));
  nor2  gate2435(.a(gate210inter11), .b(gate210inter6), .O(gate210inter12));
  nand2 gate2436(.a(gate210inter12), .b(gate210inter1), .O(G691));

  xor2  gate631(.a(G669), .b(G612), .O(gate211inter0));
  nand2 gate632(.a(gate211inter0), .b(s_12), .O(gate211inter1));
  and2  gate633(.a(G669), .b(G612), .O(gate211inter2));
  inv1  gate634(.a(s_12), .O(gate211inter3));
  inv1  gate635(.a(s_13), .O(gate211inter4));
  nand2 gate636(.a(gate211inter4), .b(gate211inter3), .O(gate211inter5));
  nor2  gate637(.a(gate211inter5), .b(gate211inter2), .O(gate211inter6));
  inv1  gate638(.a(G612), .O(gate211inter7));
  inv1  gate639(.a(G669), .O(gate211inter8));
  nand2 gate640(.a(gate211inter8), .b(gate211inter7), .O(gate211inter9));
  nand2 gate641(.a(s_13), .b(gate211inter3), .O(gate211inter10));
  nor2  gate642(.a(gate211inter10), .b(gate211inter9), .O(gate211inter11));
  nor2  gate643(.a(gate211inter11), .b(gate211inter6), .O(gate211inter12));
  nand2 gate644(.a(gate211inter12), .b(gate211inter1), .O(G692));

  xor2  gate2269(.a(G669), .b(G617), .O(gate212inter0));
  nand2 gate2270(.a(gate212inter0), .b(s_246), .O(gate212inter1));
  and2  gate2271(.a(G669), .b(G617), .O(gate212inter2));
  inv1  gate2272(.a(s_246), .O(gate212inter3));
  inv1  gate2273(.a(s_247), .O(gate212inter4));
  nand2 gate2274(.a(gate212inter4), .b(gate212inter3), .O(gate212inter5));
  nor2  gate2275(.a(gate212inter5), .b(gate212inter2), .O(gate212inter6));
  inv1  gate2276(.a(G617), .O(gate212inter7));
  inv1  gate2277(.a(G669), .O(gate212inter8));
  nand2 gate2278(.a(gate212inter8), .b(gate212inter7), .O(gate212inter9));
  nand2 gate2279(.a(s_247), .b(gate212inter3), .O(gate212inter10));
  nor2  gate2280(.a(gate212inter10), .b(gate212inter9), .O(gate212inter11));
  nor2  gate2281(.a(gate212inter11), .b(gate212inter6), .O(gate212inter12));
  nand2 gate2282(.a(gate212inter12), .b(gate212inter1), .O(G693));
nand2 gate213( .a(G602), .b(G672), .O(G694) );
nand2 gate214( .a(G612), .b(G672), .O(G695) );

  xor2  gate1583(.a(G675), .b(G607), .O(gate215inter0));
  nand2 gate1584(.a(gate215inter0), .b(s_148), .O(gate215inter1));
  and2  gate1585(.a(G675), .b(G607), .O(gate215inter2));
  inv1  gate1586(.a(s_148), .O(gate215inter3));
  inv1  gate1587(.a(s_149), .O(gate215inter4));
  nand2 gate1588(.a(gate215inter4), .b(gate215inter3), .O(gate215inter5));
  nor2  gate1589(.a(gate215inter5), .b(gate215inter2), .O(gate215inter6));
  inv1  gate1590(.a(G607), .O(gate215inter7));
  inv1  gate1591(.a(G675), .O(gate215inter8));
  nand2 gate1592(.a(gate215inter8), .b(gate215inter7), .O(gate215inter9));
  nand2 gate1593(.a(s_149), .b(gate215inter3), .O(gate215inter10));
  nor2  gate1594(.a(gate215inter10), .b(gate215inter9), .O(gate215inter11));
  nor2  gate1595(.a(gate215inter11), .b(gate215inter6), .O(gate215inter12));
  nand2 gate1596(.a(gate215inter12), .b(gate215inter1), .O(G696));

  xor2  gate911(.a(G675), .b(G617), .O(gate216inter0));
  nand2 gate912(.a(gate216inter0), .b(s_52), .O(gate216inter1));
  and2  gate913(.a(G675), .b(G617), .O(gate216inter2));
  inv1  gate914(.a(s_52), .O(gate216inter3));
  inv1  gate915(.a(s_53), .O(gate216inter4));
  nand2 gate916(.a(gate216inter4), .b(gate216inter3), .O(gate216inter5));
  nor2  gate917(.a(gate216inter5), .b(gate216inter2), .O(gate216inter6));
  inv1  gate918(.a(G617), .O(gate216inter7));
  inv1  gate919(.a(G675), .O(gate216inter8));
  nand2 gate920(.a(gate216inter8), .b(gate216inter7), .O(gate216inter9));
  nand2 gate921(.a(s_53), .b(gate216inter3), .O(gate216inter10));
  nor2  gate922(.a(gate216inter10), .b(gate216inter9), .O(gate216inter11));
  nor2  gate923(.a(gate216inter11), .b(gate216inter6), .O(gate216inter12));
  nand2 gate924(.a(gate216inter12), .b(gate216inter1), .O(G697));

  xor2  gate2101(.a(G678), .b(G622), .O(gate217inter0));
  nand2 gate2102(.a(gate217inter0), .b(s_222), .O(gate217inter1));
  and2  gate2103(.a(G678), .b(G622), .O(gate217inter2));
  inv1  gate2104(.a(s_222), .O(gate217inter3));
  inv1  gate2105(.a(s_223), .O(gate217inter4));
  nand2 gate2106(.a(gate217inter4), .b(gate217inter3), .O(gate217inter5));
  nor2  gate2107(.a(gate217inter5), .b(gate217inter2), .O(gate217inter6));
  inv1  gate2108(.a(G622), .O(gate217inter7));
  inv1  gate2109(.a(G678), .O(gate217inter8));
  nand2 gate2110(.a(gate217inter8), .b(gate217inter7), .O(gate217inter9));
  nand2 gate2111(.a(s_223), .b(gate217inter3), .O(gate217inter10));
  nor2  gate2112(.a(gate217inter10), .b(gate217inter9), .O(gate217inter11));
  nor2  gate2113(.a(gate217inter11), .b(gate217inter6), .O(gate217inter12));
  nand2 gate2114(.a(gate217inter12), .b(gate217inter1), .O(G698));
nand2 gate218( .a(G627), .b(G678), .O(G699) );
nand2 gate219( .a(G632), .b(G681), .O(G700) );
nand2 gate220( .a(G637), .b(G681), .O(G701) );
nand2 gate221( .a(G622), .b(G684), .O(G702) );
nand2 gate222( .a(G632), .b(G684), .O(G703) );
nand2 gate223( .a(G627), .b(G687), .O(G704) );

  xor2  gate1611(.a(G687), .b(G637), .O(gate224inter0));
  nand2 gate1612(.a(gate224inter0), .b(s_152), .O(gate224inter1));
  and2  gate1613(.a(G687), .b(G637), .O(gate224inter2));
  inv1  gate1614(.a(s_152), .O(gate224inter3));
  inv1  gate1615(.a(s_153), .O(gate224inter4));
  nand2 gate1616(.a(gate224inter4), .b(gate224inter3), .O(gate224inter5));
  nor2  gate1617(.a(gate224inter5), .b(gate224inter2), .O(gate224inter6));
  inv1  gate1618(.a(G637), .O(gate224inter7));
  inv1  gate1619(.a(G687), .O(gate224inter8));
  nand2 gate1620(.a(gate224inter8), .b(gate224inter7), .O(gate224inter9));
  nand2 gate1621(.a(s_153), .b(gate224inter3), .O(gate224inter10));
  nor2  gate1622(.a(gate224inter10), .b(gate224inter9), .O(gate224inter11));
  nor2  gate1623(.a(gate224inter11), .b(gate224inter6), .O(gate224inter12));
  nand2 gate1624(.a(gate224inter12), .b(gate224inter1), .O(G705));
nand2 gate225( .a(G690), .b(G691), .O(G706) );

  xor2  gate1331(.a(G693), .b(G692), .O(gate226inter0));
  nand2 gate1332(.a(gate226inter0), .b(s_112), .O(gate226inter1));
  and2  gate1333(.a(G693), .b(G692), .O(gate226inter2));
  inv1  gate1334(.a(s_112), .O(gate226inter3));
  inv1  gate1335(.a(s_113), .O(gate226inter4));
  nand2 gate1336(.a(gate226inter4), .b(gate226inter3), .O(gate226inter5));
  nor2  gate1337(.a(gate226inter5), .b(gate226inter2), .O(gate226inter6));
  inv1  gate1338(.a(G692), .O(gate226inter7));
  inv1  gate1339(.a(G693), .O(gate226inter8));
  nand2 gate1340(.a(gate226inter8), .b(gate226inter7), .O(gate226inter9));
  nand2 gate1341(.a(s_113), .b(gate226inter3), .O(gate226inter10));
  nor2  gate1342(.a(gate226inter10), .b(gate226inter9), .O(gate226inter11));
  nor2  gate1343(.a(gate226inter11), .b(gate226inter6), .O(gate226inter12));
  nand2 gate1344(.a(gate226inter12), .b(gate226inter1), .O(G709));
nand2 gate227( .a(G694), .b(G695), .O(G712) );
nand2 gate228( .a(G696), .b(G697), .O(G715) );
nand2 gate229( .a(G698), .b(G699), .O(G718) );
nand2 gate230( .a(G700), .b(G701), .O(G721) );
nand2 gate231( .a(G702), .b(G703), .O(G724) );
nand2 gate232( .a(G704), .b(G705), .O(G727) );
nand2 gate233( .a(G242), .b(G718), .O(G730) );

  xor2  gate1527(.a(G721), .b(G245), .O(gate234inter0));
  nand2 gate1528(.a(gate234inter0), .b(s_140), .O(gate234inter1));
  and2  gate1529(.a(G721), .b(G245), .O(gate234inter2));
  inv1  gate1530(.a(s_140), .O(gate234inter3));
  inv1  gate1531(.a(s_141), .O(gate234inter4));
  nand2 gate1532(.a(gate234inter4), .b(gate234inter3), .O(gate234inter5));
  nor2  gate1533(.a(gate234inter5), .b(gate234inter2), .O(gate234inter6));
  inv1  gate1534(.a(G245), .O(gate234inter7));
  inv1  gate1535(.a(G721), .O(gate234inter8));
  nand2 gate1536(.a(gate234inter8), .b(gate234inter7), .O(gate234inter9));
  nand2 gate1537(.a(s_141), .b(gate234inter3), .O(gate234inter10));
  nor2  gate1538(.a(gate234inter10), .b(gate234inter9), .O(gate234inter11));
  nor2  gate1539(.a(gate234inter11), .b(gate234inter6), .O(gate234inter12));
  nand2 gate1540(.a(gate234inter12), .b(gate234inter1), .O(G733));

  xor2  gate869(.a(G724), .b(G248), .O(gate235inter0));
  nand2 gate870(.a(gate235inter0), .b(s_46), .O(gate235inter1));
  and2  gate871(.a(G724), .b(G248), .O(gate235inter2));
  inv1  gate872(.a(s_46), .O(gate235inter3));
  inv1  gate873(.a(s_47), .O(gate235inter4));
  nand2 gate874(.a(gate235inter4), .b(gate235inter3), .O(gate235inter5));
  nor2  gate875(.a(gate235inter5), .b(gate235inter2), .O(gate235inter6));
  inv1  gate876(.a(G248), .O(gate235inter7));
  inv1  gate877(.a(G724), .O(gate235inter8));
  nand2 gate878(.a(gate235inter8), .b(gate235inter7), .O(gate235inter9));
  nand2 gate879(.a(s_47), .b(gate235inter3), .O(gate235inter10));
  nor2  gate880(.a(gate235inter10), .b(gate235inter9), .O(gate235inter11));
  nor2  gate881(.a(gate235inter11), .b(gate235inter6), .O(gate235inter12));
  nand2 gate882(.a(gate235inter12), .b(gate235inter1), .O(G736));
nand2 gate236( .a(G251), .b(G727), .O(G739) );
nand2 gate237( .a(G254), .b(G706), .O(G742) );
nand2 gate238( .a(G257), .b(G709), .O(G745) );

  xor2  gate2255(.a(G712), .b(G260), .O(gate239inter0));
  nand2 gate2256(.a(gate239inter0), .b(s_244), .O(gate239inter1));
  and2  gate2257(.a(G712), .b(G260), .O(gate239inter2));
  inv1  gate2258(.a(s_244), .O(gate239inter3));
  inv1  gate2259(.a(s_245), .O(gate239inter4));
  nand2 gate2260(.a(gate239inter4), .b(gate239inter3), .O(gate239inter5));
  nor2  gate2261(.a(gate239inter5), .b(gate239inter2), .O(gate239inter6));
  inv1  gate2262(.a(G260), .O(gate239inter7));
  inv1  gate2263(.a(G712), .O(gate239inter8));
  nand2 gate2264(.a(gate239inter8), .b(gate239inter7), .O(gate239inter9));
  nand2 gate2265(.a(s_245), .b(gate239inter3), .O(gate239inter10));
  nor2  gate2266(.a(gate239inter10), .b(gate239inter9), .O(gate239inter11));
  nor2  gate2267(.a(gate239inter11), .b(gate239inter6), .O(gate239inter12));
  nand2 gate2268(.a(gate239inter12), .b(gate239inter1), .O(G748));
nand2 gate240( .a(G263), .b(G715), .O(G751) );

  xor2  gate1135(.a(G730), .b(G242), .O(gate241inter0));
  nand2 gate1136(.a(gate241inter0), .b(s_84), .O(gate241inter1));
  and2  gate1137(.a(G730), .b(G242), .O(gate241inter2));
  inv1  gate1138(.a(s_84), .O(gate241inter3));
  inv1  gate1139(.a(s_85), .O(gate241inter4));
  nand2 gate1140(.a(gate241inter4), .b(gate241inter3), .O(gate241inter5));
  nor2  gate1141(.a(gate241inter5), .b(gate241inter2), .O(gate241inter6));
  inv1  gate1142(.a(G242), .O(gate241inter7));
  inv1  gate1143(.a(G730), .O(gate241inter8));
  nand2 gate1144(.a(gate241inter8), .b(gate241inter7), .O(gate241inter9));
  nand2 gate1145(.a(s_85), .b(gate241inter3), .O(gate241inter10));
  nor2  gate1146(.a(gate241inter10), .b(gate241inter9), .O(gate241inter11));
  nor2  gate1147(.a(gate241inter11), .b(gate241inter6), .O(gate241inter12));
  nand2 gate1148(.a(gate241inter12), .b(gate241inter1), .O(G754));
nand2 gate242( .a(G718), .b(G730), .O(G755) );
nand2 gate243( .a(G245), .b(G733), .O(G756) );

  xor2  gate2759(.a(G733), .b(G721), .O(gate244inter0));
  nand2 gate2760(.a(gate244inter0), .b(s_316), .O(gate244inter1));
  and2  gate2761(.a(G733), .b(G721), .O(gate244inter2));
  inv1  gate2762(.a(s_316), .O(gate244inter3));
  inv1  gate2763(.a(s_317), .O(gate244inter4));
  nand2 gate2764(.a(gate244inter4), .b(gate244inter3), .O(gate244inter5));
  nor2  gate2765(.a(gate244inter5), .b(gate244inter2), .O(gate244inter6));
  inv1  gate2766(.a(G721), .O(gate244inter7));
  inv1  gate2767(.a(G733), .O(gate244inter8));
  nand2 gate2768(.a(gate244inter8), .b(gate244inter7), .O(gate244inter9));
  nand2 gate2769(.a(s_317), .b(gate244inter3), .O(gate244inter10));
  nor2  gate2770(.a(gate244inter10), .b(gate244inter9), .O(gate244inter11));
  nor2  gate2771(.a(gate244inter11), .b(gate244inter6), .O(gate244inter12));
  nand2 gate2772(.a(gate244inter12), .b(gate244inter1), .O(G757));
nand2 gate245( .a(G248), .b(G736), .O(G758) );
nand2 gate246( .a(G724), .b(G736), .O(G759) );
nand2 gate247( .a(G251), .b(G739), .O(G760) );

  xor2  gate953(.a(G739), .b(G727), .O(gate248inter0));
  nand2 gate954(.a(gate248inter0), .b(s_58), .O(gate248inter1));
  and2  gate955(.a(G739), .b(G727), .O(gate248inter2));
  inv1  gate956(.a(s_58), .O(gate248inter3));
  inv1  gate957(.a(s_59), .O(gate248inter4));
  nand2 gate958(.a(gate248inter4), .b(gate248inter3), .O(gate248inter5));
  nor2  gate959(.a(gate248inter5), .b(gate248inter2), .O(gate248inter6));
  inv1  gate960(.a(G727), .O(gate248inter7));
  inv1  gate961(.a(G739), .O(gate248inter8));
  nand2 gate962(.a(gate248inter8), .b(gate248inter7), .O(gate248inter9));
  nand2 gate963(.a(s_59), .b(gate248inter3), .O(gate248inter10));
  nor2  gate964(.a(gate248inter10), .b(gate248inter9), .O(gate248inter11));
  nor2  gate965(.a(gate248inter11), .b(gate248inter6), .O(gate248inter12));
  nand2 gate966(.a(gate248inter12), .b(gate248inter1), .O(G761));

  xor2  gate813(.a(G742), .b(G254), .O(gate249inter0));
  nand2 gate814(.a(gate249inter0), .b(s_38), .O(gate249inter1));
  and2  gate815(.a(G742), .b(G254), .O(gate249inter2));
  inv1  gate816(.a(s_38), .O(gate249inter3));
  inv1  gate817(.a(s_39), .O(gate249inter4));
  nand2 gate818(.a(gate249inter4), .b(gate249inter3), .O(gate249inter5));
  nor2  gate819(.a(gate249inter5), .b(gate249inter2), .O(gate249inter6));
  inv1  gate820(.a(G254), .O(gate249inter7));
  inv1  gate821(.a(G742), .O(gate249inter8));
  nand2 gate822(.a(gate249inter8), .b(gate249inter7), .O(gate249inter9));
  nand2 gate823(.a(s_39), .b(gate249inter3), .O(gate249inter10));
  nor2  gate824(.a(gate249inter10), .b(gate249inter9), .O(gate249inter11));
  nor2  gate825(.a(gate249inter11), .b(gate249inter6), .O(gate249inter12));
  nand2 gate826(.a(gate249inter12), .b(gate249inter1), .O(G762));

  xor2  gate1065(.a(G742), .b(G706), .O(gate250inter0));
  nand2 gate1066(.a(gate250inter0), .b(s_74), .O(gate250inter1));
  and2  gate1067(.a(G742), .b(G706), .O(gate250inter2));
  inv1  gate1068(.a(s_74), .O(gate250inter3));
  inv1  gate1069(.a(s_75), .O(gate250inter4));
  nand2 gate1070(.a(gate250inter4), .b(gate250inter3), .O(gate250inter5));
  nor2  gate1071(.a(gate250inter5), .b(gate250inter2), .O(gate250inter6));
  inv1  gate1072(.a(G706), .O(gate250inter7));
  inv1  gate1073(.a(G742), .O(gate250inter8));
  nand2 gate1074(.a(gate250inter8), .b(gate250inter7), .O(gate250inter9));
  nand2 gate1075(.a(s_75), .b(gate250inter3), .O(gate250inter10));
  nor2  gate1076(.a(gate250inter10), .b(gate250inter9), .O(gate250inter11));
  nor2  gate1077(.a(gate250inter11), .b(gate250inter6), .O(gate250inter12));
  nand2 gate1078(.a(gate250inter12), .b(gate250inter1), .O(G763));
nand2 gate251( .a(G257), .b(G745), .O(G764) );

  xor2  gate2031(.a(G745), .b(G709), .O(gate252inter0));
  nand2 gate2032(.a(gate252inter0), .b(s_212), .O(gate252inter1));
  and2  gate2033(.a(G745), .b(G709), .O(gate252inter2));
  inv1  gate2034(.a(s_212), .O(gate252inter3));
  inv1  gate2035(.a(s_213), .O(gate252inter4));
  nand2 gate2036(.a(gate252inter4), .b(gate252inter3), .O(gate252inter5));
  nor2  gate2037(.a(gate252inter5), .b(gate252inter2), .O(gate252inter6));
  inv1  gate2038(.a(G709), .O(gate252inter7));
  inv1  gate2039(.a(G745), .O(gate252inter8));
  nand2 gate2040(.a(gate252inter8), .b(gate252inter7), .O(gate252inter9));
  nand2 gate2041(.a(s_213), .b(gate252inter3), .O(gate252inter10));
  nor2  gate2042(.a(gate252inter10), .b(gate252inter9), .O(gate252inter11));
  nor2  gate2043(.a(gate252inter11), .b(gate252inter6), .O(gate252inter12));
  nand2 gate2044(.a(gate252inter12), .b(gate252inter1), .O(G765));
nand2 gate253( .a(G260), .b(G748), .O(G766) );
nand2 gate254( .a(G712), .b(G748), .O(G767) );

  xor2  gate1499(.a(G751), .b(G263), .O(gate255inter0));
  nand2 gate1500(.a(gate255inter0), .b(s_136), .O(gate255inter1));
  and2  gate1501(.a(G751), .b(G263), .O(gate255inter2));
  inv1  gate1502(.a(s_136), .O(gate255inter3));
  inv1  gate1503(.a(s_137), .O(gate255inter4));
  nand2 gate1504(.a(gate255inter4), .b(gate255inter3), .O(gate255inter5));
  nor2  gate1505(.a(gate255inter5), .b(gate255inter2), .O(gate255inter6));
  inv1  gate1506(.a(G263), .O(gate255inter7));
  inv1  gate1507(.a(G751), .O(gate255inter8));
  nand2 gate1508(.a(gate255inter8), .b(gate255inter7), .O(gate255inter9));
  nand2 gate1509(.a(s_137), .b(gate255inter3), .O(gate255inter10));
  nor2  gate1510(.a(gate255inter10), .b(gate255inter9), .O(gate255inter11));
  nor2  gate1511(.a(gate255inter11), .b(gate255inter6), .O(gate255inter12));
  nand2 gate1512(.a(gate255inter12), .b(gate255inter1), .O(G768));

  xor2  gate743(.a(G751), .b(G715), .O(gate256inter0));
  nand2 gate744(.a(gate256inter0), .b(s_28), .O(gate256inter1));
  and2  gate745(.a(G751), .b(G715), .O(gate256inter2));
  inv1  gate746(.a(s_28), .O(gate256inter3));
  inv1  gate747(.a(s_29), .O(gate256inter4));
  nand2 gate748(.a(gate256inter4), .b(gate256inter3), .O(gate256inter5));
  nor2  gate749(.a(gate256inter5), .b(gate256inter2), .O(gate256inter6));
  inv1  gate750(.a(G715), .O(gate256inter7));
  inv1  gate751(.a(G751), .O(gate256inter8));
  nand2 gate752(.a(gate256inter8), .b(gate256inter7), .O(gate256inter9));
  nand2 gate753(.a(s_29), .b(gate256inter3), .O(gate256inter10));
  nor2  gate754(.a(gate256inter10), .b(gate256inter9), .O(gate256inter11));
  nor2  gate755(.a(gate256inter11), .b(gate256inter6), .O(gate256inter12));
  nand2 gate756(.a(gate256inter12), .b(gate256inter1), .O(G769));
nand2 gate257( .a(G754), .b(G755), .O(G770) );
nand2 gate258( .a(G756), .b(G757), .O(G773) );
nand2 gate259( .a(G758), .b(G759), .O(G776) );
nand2 gate260( .a(G760), .b(G761), .O(G779) );

  xor2  gate1345(.a(G763), .b(G762), .O(gate261inter0));
  nand2 gate1346(.a(gate261inter0), .b(s_114), .O(gate261inter1));
  and2  gate1347(.a(G763), .b(G762), .O(gate261inter2));
  inv1  gate1348(.a(s_114), .O(gate261inter3));
  inv1  gate1349(.a(s_115), .O(gate261inter4));
  nand2 gate1350(.a(gate261inter4), .b(gate261inter3), .O(gate261inter5));
  nor2  gate1351(.a(gate261inter5), .b(gate261inter2), .O(gate261inter6));
  inv1  gate1352(.a(G762), .O(gate261inter7));
  inv1  gate1353(.a(G763), .O(gate261inter8));
  nand2 gate1354(.a(gate261inter8), .b(gate261inter7), .O(gate261inter9));
  nand2 gate1355(.a(s_115), .b(gate261inter3), .O(gate261inter10));
  nor2  gate1356(.a(gate261inter10), .b(gate261inter9), .O(gate261inter11));
  nor2  gate1357(.a(gate261inter11), .b(gate261inter6), .O(gate261inter12));
  nand2 gate1358(.a(gate261inter12), .b(gate261inter1), .O(G782));
nand2 gate262( .a(G764), .b(G765), .O(G785) );
nand2 gate263( .a(G766), .b(G767), .O(G788) );

  xor2  gate1667(.a(G769), .b(G768), .O(gate264inter0));
  nand2 gate1668(.a(gate264inter0), .b(s_160), .O(gate264inter1));
  and2  gate1669(.a(G769), .b(G768), .O(gate264inter2));
  inv1  gate1670(.a(s_160), .O(gate264inter3));
  inv1  gate1671(.a(s_161), .O(gate264inter4));
  nand2 gate1672(.a(gate264inter4), .b(gate264inter3), .O(gate264inter5));
  nor2  gate1673(.a(gate264inter5), .b(gate264inter2), .O(gate264inter6));
  inv1  gate1674(.a(G768), .O(gate264inter7));
  inv1  gate1675(.a(G769), .O(gate264inter8));
  nand2 gate1676(.a(gate264inter8), .b(gate264inter7), .O(gate264inter9));
  nand2 gate1677(.a(s_161), .b(gate264inter3), .O(gate264inter10));
  nor2  gate1678(.a(gate264inter10), .b(gate264inter9), .O(gate264inter11));
  nor2  gate1679(.a(gate264inter11), .b(gate264inter6), .O(gate264inter12));
  nand2 gate1680(.a(gate264inter12), .b(gate264inter1), .O(G791));
nand2 gate265( .a(G642), .b(G770), .O(G794) );

  xor2  gate1457(.a(G773), .b(G645), .O(gate266inter0));
  nand2 gate1458(.a(gate266inter0), .b(s_130), .O(gate266inter1));
  and2  gate1459(.a(G773), .b(G645), .O(gate266inter2));
  inv1  gate1460(.a(s_130), .O(gate266inter3));
  inv1  gate1461(.a(s_131), .O(gate266inter4));
  nand2 gate1462(.a(gate266inter4), .b(gate266inter3), .O(gate266inter5));
  nor2  gate1463(.a(gate266inter5), .b(gate266inter2), .O(gate266inter6));
  inv1  gate1464(.a(G645), .O(gate266inter7));
  inv1  gate1465(.a(G773), .O(gate266inter8));
  nand2 gate1466(.a(gate266inter8), .b(gate266inter7), .O(gate266inter9));
  nand2 gate1467(.a(s_131), .b(gate266inter3), .O(gate266inter10));
  nor2  gate1468(.a(gate266inter10), .b(gate266inter9), .O(gate266inter11));
  nor2  gate1469(.a(gate266inter11), .b(gate266inter6), .O(gate266inter12));
  nand2 gate1470(.a(gate266inter12), .b(gate266inter1), .O(G797));

  xor2  gate1569(.a(G776), .b(G648), .O(gate267inter0));
  nand2 gate1570(.a(gate267inter0), .b(s_146), .O(gate267inter1));
  and2  gate1571(.a(G776), .b(G648), .O(gate267inter2));
  inv1  gate1572(.a(s_146), .O(gate267inter3));
  inv1  gate1573(.a(s_147), .O(gate267inter4));
  nand2 gate1574(.a(gate267inter4), .b(gate267inter3), .O(gate267inter5));
  nor2  gate1575(.a(gate267inter5), .b(gate267inter2), .O(gate267inter6));
  inv1  gate1576(.a(G648), .O(gate267inter7));
  inv1  gate1577(.a(G776), .O(gate267inter8));
  nand2 gate1578(.a(gate267inter8), .b(gate267inter7), .O(gate267inter9));
  nand2 gate1579(.a(s_147), .b(gate267inter3), .O(gate267inter10));
  nor2  gate1580(.a(gate267inter10), .b(gate267inter9), .O(gate267inter11));
  nor2  gate1581(.a(gate267inter11), .b(gate267inter6), .O(gate267inter12));
  nand2 gate1582(.a(gate267inter12), .b(gate267inter1), .O(G800));
nand2 gate268( .a(G651), .b(G779), .O(G803) );

  xor2  gate1807(.a(G782), .b(G654), .O(gate269inter0));
  nand2 gate1808(.a(gate269inter0), .b(s_180), .O(gate269inter1));
  and2  gate1809(.a(G782), .b(G654), .O(gate269inter2));
  inv1  gate1810(.a(s_180), .O(gate269inter3));
  inv1  gate1811(.a(s_181), .O(gate269inter4));
  nand2 gate1812(.a(gate269inter4), .b(gate269inter3), .O(gate269inter5));
  nor2  gate1813(.a(gate269inter5), .b(gate269inter2), .O(gate269inter6));
  inv1  gate1814(.a(G654), .O(gate269inter7));
  inv1  gate1815(.a(G782), .O(gate269inter8));
  nand2 gate1816(.a(gate269inter8), .b(gate269inter7), .O(gate269inter9));
  nand2 gate1817(.a(s_181), .b(gate269inter3), .O(gate269inter10));
  nor2  gate1818(.a(gate269inter10), .b(gate269inter9), .O(gate269inter11));
  nor2  gate1819(.a(gate269inter11), .b(gate269inter6), .O(gate269inter12));
  nand2 gate1820(.a(gate269inter12), .b(gate269inter1), .O(G806));

  xor2  gate1429(.a(G785), .b(G657), .O(gate270inter0));
  nand2 gate1430(.a(gate270inter0), .b(s_126), .O(gate270inter1));
  and2  gate1431(.a(G785), .b(G657), .O(gate270inter2));
  inv1  gate1432(.a(s_126), .O(gate270inter3));
  inv1  gate1433(.a(s_127), .O(gate270inter4));
  nand2 gate1434(.a(gate270inter4), .b(gate270inter3), .O(gate270inter5));
  nor2  gate1435(.a(gate270inter5), .b(gate270inter2), .O(gate270inter6));
  inv1  gate1436(.a(G657), .O(gate270inter7));
  inv1  gate1437(.a(G785), .O(gate270inter8));
  nand2 gate1438(.a(gate270inter8), .b(gate270inter7), .O(gate270inter9));
  nand2 gate1439(.a(s_127), .b(gate270inter3), .O(gate270inter10));
  nor2  gate1440(.a(gate270inter10), .b(gate270inter9), .O(gate270inter11));
  nor2  gate1441(.a(gate270inter11), .b(gate270inter6), .O(gate270inter12));
  nand2 gate1442(.a(gate270inter12), .b(gate270inter1), .O(G809));

  xor2  gate1093(.a(G788), .b(G660), .O(gate271inter0));
  nand2 gate1094(.a(gate271inter0), .b(s_78), .O(gate271inter1));
  and2  gate1095(.a(G788), .b(G660), .O(gate271inter2));
  inv1  gate1096(.a(s_78), .O(gate271inter3));
  inv1  gate1097(.a(s_79), .O(gate271inter4));
  nand2 gate1098(.a(gate271inter4), .b(gate271inter3), .O(gate271inter5));
  nor2  gate1099(.a(gate271inter5), .b(gate271inter2), .O(gate271inter6));
  inv1  gate1100(.a(G660), .O(gate271inter7));
  inv1  gate1101(.a(G788), .O(gate271inter8));
  nand2 gate1102(.a(gate271inter8), .b(gate271inter7), .O(gate271inter9));
  nand2 gate1103(.a(s_79), .b(gate271inter3), .O(gate271inter10));
  nor2  gate1104(.a(gate271inter10), .b(gate271inter9), .O(gate271inter11));
  nor2  gate1105(.a(gate271inter11), .b(gate271inter6), .O(gate271inter12));
  nand2 gate1106(.a(gate271inter12), .b(gate271inter1), .O(G812));
nand2 gate272( .a(G663), .b(G791), .O(G815) );
nand2 gate273( .a(G642), .b(G794), .O(G818) );

  xor2  gate1681(.a(G794), .b(G770), .O(gate274inter0));
  nand2 gate1682(.a(gate274inter0), .b(s_162), .O(gate274inter1));
  and2  gate1683(.a(G794), .b(G770), .O(gate274inter2));
  inv1  gate1684(.a(s_162), .O(gate274inter3));
  inv1  gate1685(.a(s_163), .O(gate274inter4));
  nand2 gate1686(.a(gate274inter4), .b(gate274inter3), .O(gate274inter5));
  nor2  gate1687(.a(gate274inter5), .b(gate274inter2), .O(gate274inter6));
  inv1  gate1688(.a(G770), .O(gate274inter7));
  inv1  gate1689(.a(G794), .O(gate274inter8));
  nand2 gate1690(.a(gate274inter8), .b(gate274inter7), .O(gate274inter9));
  nand2 gate1691(.a(s_163), .b(gate274inter3), .O(gate274inter10));
  nor2  gate1692(.a(gate274inter10), .b(gate274inter9), .O(gate274inter11));
  nor2  gate1693(.a(gate274inter11), .b(gate274inter6), .O(gate274inter12));
  nand2 gate1694(.a(gate274inter12), .b(gate274inter1), .O(G819));

  xor2  gate701(.a(G797), .b(G645), .O(gate275inter0));
  nand2 gate702(.a(gate275inter0), .b(s_22), .O(gate275inter1));
  and2  gate703(.a(G797), .b(G645), .O(gate275inter2));
  inv1  gate704(.a(s_22), .O(gate275inter3));
  inv1  gate705(.a(s_23), .O(gate275inter4));
  nand2 gate706(.a(gate275inter4), .b(gate275inter3), .O(gate275inter5));
  nor2  gate707(.a(gate275inter5), .b(gate275inter2), .O(gate275inter6));
  inv1  gate708(.a(G645), .O(gate275inter7));
  inv1  gate709(.a(G797), .O(gate275inter8));
  nand2 gate710(.a(gate275inter8), .b(gate275inter7), .O(gate275inter9));
  nand2 gate711(.a(s_23), .b(gate275inter3), .O(gate275inter10));
  nor2  gate712(.a(gate275inter10), .b(gate275inter9), .O(gate275inter11));
  nor2  gate713(.a(gate275inter11), .b(gate275inter6), .O(gate275inter12));
  nand2 gate714(.a(gate275inter12), .b(gate275inter1), .O(G820));

  xor2  gate2451(.a(G797), .b(G773), .O(gate276inter0));
  nand2 gate2452(.a(gate276inter0), .b(s_272), .O(gate276inter1));
  and2  gate2453(.a(G797), .b(G773), .O(gate276inter2));
  inv1  gate2454(.a(s_272), .O(gate276inter3));
  inv1  gate2455(.a(s_273), .O(gate276inter4));
  nand2 gate2456(.a(gate276inter4), .b(gate276inter3), .O(gate276inter5));
  nor2  gate2457(.a(gate276inter5), .b(gate276inter2), .O(gate276inter6));
  inv1  gate2458(.a(G773), .O(gate276inter7));
  inv1  gate2459(.a(G797), .O(gate276inter8));
  nand2 gate2460(.a(gate276inter8), .b(gate276inter7), .O(gate276inter9));
  nand2 gate2461(.a(s_273), .b(gate276inter3), .O(gate276inter10));
  nor2  gate2462(.a(gate276inter10), .b(gate276inter9), .O(gate276inter11));
  nor2  gate2463(.a(gate276inter11), .b(gate276inter6), .O(gate276inter12));
  nand2 gate2464(.a(gate276inter12), .b(gate276inter1), .O(G821));

  xor2  gate1219(.a(G800), .b(G648), .O(gate277inter0));
  nand2 gate1220(.a(gate277inter0), .b(s_96), .O(gate277inter1));
  and2  gate1221(.a(G800), .b(G648), .O(gate277inter2));
  inv1  gate1222(.a(s_96), .O(gate277inter3));
  inv1  gate1223(.a(s_97), .O(gate277inter4));
  nand2 gate1224(.a(gate277inter4), .b(gate277inter3), .O(gate277inter5));
  nor2  gate1225(.a(gate277inter5), .b(gate277inter2), .O(gate277inter6));
  inv1  gate1226(.a(G648), .O(gate277inter7));
  inv1  gate1227(.a(G800), .O(gate277inter8));
  nand2 gate1228(.a(gate277inter8), .b(gate277inter7), .O(gate277inter9));
  nand2 gate1229(.a(s_97), .b(gate277inter3), .O(gate277inter10));
  nor2  gate1230(.a(gate277inter10), .b(gate277inter9), .O(gate277inter11));
  nor2  gate1231(.a(gate277inter11), .b(gate277inter6), .O(gate277inter12));
  nand2 gate1232(.a(gate277inter12), .b(gate277inter1), .O(G822));
nand2 gate278( .a(G776), .b(G800), .O(G823) );

  xor2  gate2731(.a(G803), .b(G651), .O(gate279inter0));
  nand2 gate2732(.a(gate279inter0), .b(s_312), .O(gate279inter1));
  and2  gate2733(.a(G803), .b(G651), .O(gate279inter2));
  inv1  gate2734(.a(s_312), .O(gate279inter3));
  inv1  gate2735(.a(s_313), .O(gate279inter4));
  nand2 gate2736(.a(gate279inter4), .b(gate279inter3), .O(gate279inter5));
  nor2  gate2737(.a(gate279inter5), .b(gate279inter2), .O(gate279inter6));
  inv1  gate2738(.a(G651), .O(gate279inter7));
  inv1  gate2739(.a(G803), .O(gate279inter8));
  nand2 gate2740(.a(gate279inter8), .b(gate279inter7), .O(gate279inter9));
  nand2 gate2741(.a(s_313), .b(gate279inter3), .O(gate279inter10));
  nor2  gate2742(.a(gate279inter10), .b(gate279inter9), .O(gate279inter11));
  nor2  gate2743(.a(gate279inter11), .b(gate279inter6), .O(gate279inter12));
  nand2 gate2744(.a(gate279inter12), .b(gate279inter1), .O(G824));

  xor2  gate1289(.a(G803), .b(G779), .O(gate280inter0));
  nand2 gate1290(.a(gate280inter0), .b(s_106), .O(gate280inter1));
  and2  gate1291(.a(G803), .b(G779), .O(gate280inter2));
  inv1  gate1292(.a(s_106), .O(gate280inter3));
  inv1  gate1293(.a(s_107), .O(gate280inter4));
  nand2 gate1294(.a(gate280inter4), .b(gate280inter3), .O(gate280inter5));
  nor2  gate1295(.a(gate280inter5), .b(gate280inter2), .O(gate280inter6));
  inv1  gate1296(.a(G779), .O(gate280inter7));
  inv1  gate1297(.a(G803), .O(gate280inter8));
  nand2 gate1298(.a(gate280inter8), .b(gate280inter7), .O(gate280inter9));
  nand2 gate1299(.a(s_107), .b(gate280inter3), .O(gate280inter10));
  nor2  gate1300(.a(gate280inter10), .b(gate280inter9), .O(gate280inter11));
  nor2  gate1301(.a(gate280inter11), .b(gate280inter6), .O(gate280inter12));
  nand2 gate1302(.a(gate280inter12), .b(gate280inter1), .O(G825));
nand2 gate281( .a(G654), .b(G806), .O(G826) );
nand2 gate282( .a(G782), .b(G806), .O(G827) );
nand2 gate283( .a(G657), .b(G809), .O(G828) );
nand2 gate284( .a(G785), .b(G809), .O(G829) );
nand2 gate285( .a(G660), .b(G812), .O(G830) );
nand2 gate286( .a(G788), .b(G812), .O(G831) );

  xor2  gate2311(.a(G815), .b(G663), .O(gate287inter0));
  nand2 gate2312(.a(gate287inter0), .b(s_252), .O(gate287inter1));
  and2  gate2313(.a(G815), .b(G663), .O(gate287inter2));
  inv1  gate2314(.a(s_252), .O(gate287inter3));
  inv1  gate2315(.a(s_253), .O(gate287inter4));
  nand2 gate2316(.a(gate287inter4), .b(gate287inter3), .O(gate287inter5));
  nor2  gate2317(.a(gate287inter5), .b(gate287inter2), .O(gate287inter6));
  inv1  gate2318(.a(G663), .O(gate287inter7));
  inv1  gate2319(.a(G815), .O(gate287inter8));
  nand2 gate2320(.a(gate287inter8), .b(gate287inter7), .O(gate287inter9));
  nand2 gate2321(.a(s_253), .b(gate287inter3), .O(gate287inter10));
  nor2  gate2322(.a(gate287inter10), .b(gate287inter9), .O(gate287inter11));
  nor2  gate2323(.a(gate287inter11), .b(gate287inter6), .O(gate287inter12));
  nand2 gate2324(.a(gate287inter12), .b(gate287inter1), .O(G832));
nand2 gate288( .a(G791), .b(G815), .O(G833) );
nand2 gate289( .a(G818), .b(G819), .O(G834) );
nand2 gate290( .a(G820), .b(G821), .O(G847) );

  xor2  gate1359(.a(G823), .b(G822), .O(gate291inter0));
  nand2 gate1360(.a(gate291inter0), .b(s_116), .O(gate291inter1));
  and2  gate1361(.a(G823), .b(G822), .O(gate291inter2));
  inv1  gate1362(.a(s_116), .O(gate291inter3));
  inv1  gate1363(.a(s_117), .O(gate291inter4));
  nand2 gate1364(.a(gate291inter4), .b(gate291inter3), .O(gate291inter5));
  nor2  gate1365(.a(gate291inter5), .b(gate291inter2), .O(gate291inter6));
  inv1  gate1366(.a(G822), .O(gate291inter7));
  inv1  gate1367(.a(G823), .O(gate291inter8));
  nand2 gate1368(.a(gate291inter8), .b(gate291inter7), .O(gate291inter9));
  nand2 gate1369(.a(s_117), .b(gate291inter3), .O(gate291inter10));
  nor2  gate1370(.a(gate291inter10), .b(gate291inter9), .O(gate291inter11));
  nor2  gate1371(.a(gate291inter11), .b(gate291inter6), .O(gate291inter12));
  nand2 gate1372(.a(gate291inter12), .b(gate291inter1), .O(G860));

  xor2  gate785(.a(G825), .b(G824), .O(gate292inter0));
  nand2 gate786(.a(gate292inter0), .b(s_34), .O(gate292inter1));
  and2  gate787(.a(G825), .b(G824), .O(gate292inter2));
  inv1  gate788(.a(s_34), .O(gate292inter3));
  inv1  gate789(.a(s_35), .O(gate292inter4));
  nand2 gate790(.a(gate292inter4), .b(gate292inter3), .O(gate292inter5));
  nor2  gate791(.a(gate292inter5), .b(gate292inter2), .O(gate292inter6));
  inv1  gate792(.a(G824), .O(gate292inter7));
  inv1  gate793(.a(G825), .O(gate292inter8));
  nand2 gate794(.a(gate292inter8), .b(gate292inter7), .O(gate292inter9));
  nand2 gate795(.a(s_35), .b(gate292inter3), .O(gate292inter10));
  nor2  gate796(.a(gate292inter10), .b(gate292inter9), .O(gate292inter11));
  nor2  gate797(.a(gate292inter11), .b(gate292inter6), .O(gate292inter12));
  nand2 gate798(.a(gate292inter12), .b(gate292inter1), .O(G873));

  xor2  gate2717(.a(G829), .b(G828), .O(gate293inter0));
  nand2 gate2718(.a(gate293inter0), .b(s_310), .O(gate293inter1));
  and2  gate2719(.a(G829), .b(G828), .O(gate293inter2));
  inv1  gate2720(.a(s_310), .O(gate293inter3));
  inv1  gate2721(.a(s_311), .O(gate293inter4));
  nand2 gate2722(.a(gate293inter4), .b(gate293inter3), .O(gate293inter5));
  nor2  gate2723(.a(gate293inter5), .b(gate293inter2), .O(gate293inter6));
  inv1  gate2724(.a(G828), .O(gate293inter7));
  inv1  gate2725(.a(G829), .O(gate293inter8));
  nand2 gate2726(.a(gate293inter8), .b(gate293inter7), .O(gate293inter9));
  nand2 gate2727(.a(s_311), .b(gate293inter3), .O(gate293inter10));
  nor2  gate2728(.a(gate293inter10), .b(gate293inter9), .O(gate293inter11));
  nor2  gate2729(.a(gate293inter11), .b(gate293inter6), .O(gate293inter12));
  nand2 gate2730(.a(gate293inter12), .b(gate293inter1), .O(G886));

  xor2  gate2619(.a(G833), .b(G832), .O(gate294inter0));
  nand2 gate2620(.a(gate294inter0), .b(s_296), .O(gate294inter1));
  and2  gate2621(.a(G833), .b(G832), .O(gate294inter2));
  inv1  gate2622(.a(s_296), .O(gate294inter3));
  inv1  gate2623(.a(s_297), .O(gate294inter4));
  nand2 gate2624(.a(gate294inter4), .b(gate294inter3), .O(gate294inter5));
  nor2  gate2625(.a(gate294inter5), .b(gate294inter2), .O(gate294inter6));
  inv1  gate2626(.a(G832), .O(gate294inter7));
  inv1  gate2627(.a(G833), .O(gate294inter8));
  nand2 gate2628(.a(gate294inter8), .b(gate294inter7), .O(gate294inter9));
  nand2 gate2629(.a(s_297), .b(gate294inter3), .O(gate294inter10));
  nor2  gate2630(.a(gate294inter10), .b(gate294inter9), .O(gate294inter11));
  nor2  gate2631(.a(gate294inter11), .b(gate294inter6), .O(gate294inter12));
  nand2 gate2632(.a(gate294inter12), .b(gate294inter1), .O(G899));
nand2 gate295( .a(G830), .b(G831), .O(G912) );

  xor2  gate2913(.a(G827), .b(G826), .O(gate296inter0));
  nand2 gate2914(.a(gate296inter0), .b(s_338), .O(gate296inter1));
  and2  gate2915(.a(G827), .b(G826), .O(gate296inter2));
  inv1  gate2916(.a(s_338), .O(gate296inter3));
  inv1  gate2917(.a(s_339), .O(gate296inter4));
  nand2 gate2918(.a(gate296inter4), .b(gate296inter3), .O(gate296inter5));
  nor2  gate2919(.a(gate296inter5), .b(gate296inter2), .O(gate296inter6));
  inv1  gate2920(.a(G826), .O(gate296inter7));
  inv1  gate2921(.a(G827), .O(gate296inter8));
  nand2 gate2922(.a(gate296inter8), .b(gate296inter7), .O(gate296inter9));
  nand2 gate2923(.a(s_339), .b(gate296inter3), .O(gate296inter10));
  nor2  gate2924(.a(gate296inter10), .b(gate296inter9), .O(gate296inter11));
  nor2  gate2925(.a(gate296inter11), .b(gate296inter6), .O(gate296inter12));
  nand2 gate2926(.a(gate296inter12), .b(gate296inter1), .O(G925));
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );
nand2 gate387( .a(G1), .b(G1036), .O(G1132) );
nand2 gate388( .a(G2), .b(G1039), .O(G1135) );
nand2 gate389( .a(G3), .b(G1042), .O(G1138) );
nand2 gate390( .a(G4), .b(G1045), .O(G1141) );
nand2 gate391( .a(G5), .b(G1048), .O(G1144) );
nand2 gate392( .a(G6), .b(G1051), .O(G1147) );
nand2 gate393( .a(G7), .b(G1054), .O(G1150) );
nand2 gate394( .a(G8), .b(G1057), .O(G1153) );
nand2 gate395( .a(G9), .b(G1060), .O(G1156) );

  xor2  gate757(.a(G1063), .b(G10), .O(gate396inter0));
  nand2 gate758(.a(gate396inter0), .b(s_30), .O(gate396inter1));
  and2  gate759(.a(G1063), .b(G10), .O(gate396inter2));
  inv1  gate760(.a(s_30), .O(gate396inter3));
  inv1  gate761(.a(s_31), .O(gate396inter4));
  nand2 gate762(.a(gate396inter4), .b(gate396inter3), .O(gate396inter5));
  nor2  gate763(.a(gate396inter5), .b(gate396inter2), .O(gate396inter6));
  inv1  gate764(.a(G10), .O(gate396inter7));
  inv1  gate765(.a(G1063), .O(gate396inter8));
  nand2 gate766(.a(gate396inter8), .b(gate396inter7), .O(gate396inter9));
  nand2 gate767(.a(s_31), .b(gate396inter3), .O(gate396inter10));
  nor2  gate768(.a(gate396inter10), .b(gate396inter9), .O(gate396inter11));
  nor2  gate769(.a(gate396inter11), .b(gate396inter6), .O(gate396inter12));
  nand2 gate770(.a(gate396inter12), .b(gate396inter1), .O(G1159));

  xor2  gate1737(.a(G1066), .b(G11), .O(gate397inter0));
  nand2 gate1738(.a(gate397inter0), .b(s_170), .O(gate397inter1));
  and2  gate1739(.a(G1066), .b(G11), .O(gate397inter2));
  inv1  gate1740(.a(s_170), .O(gate397inter3));
  inv1  gate1741(.a(s_171), .O(gate397inter4));
  nand2 gate1742(.a(gate397inter4), .b(gate397inter3), .O(gate397inter5));
  nor2  gate1743(.a(gate397inter5), .b(gate397inter2), .O(gate397inter6));
  inv1  gate1744(.a(G11), .O(gate397inter7));
  inv1  gate1745(.a(G1066), .O(gate397inter8));
  nand2 gate1746(.a(gate397inter8), .b(gate397inter7), .O(gate397inter9));
  nand2 gate1747(.a(s_171), .b(gate397inter3), .O(gate397inter10));
  nor2  gate1748(.a(gate397inter10), .b(gate397inter9), .O(gate397inter11));
  nor2  gate1749(.a(gate397inter11), .b(gate397inter6), .O(gate397inter12));
  nand2 gate1750(.a(gate397inter12), .b(gate397inter1), .O(G1162));

  xor2  gate1471(.a(G1069), .b(G12), .O(gate398inter0));
  nand2 gate1472(.a(gate398inter0), .b(s_132), .O(gate398inter1));
  and2  gate1473(.a(G1069), .b(G12), .O(gate398inter2));
  inv1  gate1474(.a(s_132), .O(gate398inter3));
  inv1  gate1475(.a(s_133), .O(gate398inter4));
  nand2 gate1476(.a(gate398inter4), .b(gate398inter3), .O(gate398inter5));
  nor2  gate1477(.a(gate398inter5), .b(gate398inter2), .O(gate398inter6));
  inv1  gate1478(.a(G12), .O(gate398inter7));
  inv1  gate1479(.a(G1069), .O(gate398inter8));
  nand2 gate1480(.a(gate398inter8), .b(gate398inter7), .O(gate398inter9));
  nand2 gate1481(.a(s_133), .b(gate398inter3), .O(gate398inter10));
  nor2  gate1482(.a(gate398inter10), .b(gate398inter9), .O(gate398inter11));
  nor2  gate1483(.a(gate398inter11), .b(gate398inter6), .O(gate398inter12));
  nand2 gate1484(.a(gate398inter12), .b(gate398inter1), .O(G1165));
nand2 gate399( .a(G13), .b(G1072), .O(G1168) );

  xor2  gate967(.a(G1075), .b(G14), .O(gate400inter0));
  nand2 gate968(.a(gate400inter0), .b(s_60), .O(gate400inter1));
  and2  gate969(.a(G1075), .b(G14), .O(gate400inter2));
  inv1  gate970(.a(s_60), .O(gate400inter3));
  inv1  gate971(.a(s_61), .O(gate400inter4));
  nand2 gate972(.a(gate400inter4), .b(gate400inter3), .O(gate400inter5));
  nor2  gate973(.a(gate400inter5), .b(gate400inter2), .O(gate400inter6));
  inv1  gate974(.a(G14), .O(gate400inter7));
  inv1  gate975(.a(G1075), .O(gate400inter8));
  nand2 gate976(.a(gate400inter8), .b(gate400inter7), .O(gate400inter9));
  nand2 gate977(.a(s_61), .b(gate400inter3), .O(gate400inter10));
  nor2  gate978(.a(gate400inter10), .b(gate400inter9), .O(gate400inter11));
  nor2  gate979(.a(gate400inter11), .b(gate400inter6), .O(gate400inter12));
  nand2 gate980(.a(gate400inter12), .b(gate400inter1), .O(G1171));

  xor2  gate2003(.a(G1078), .b(G15), .O(gate401inter0));
  nand2 gate2004(.a(gate401inter0), .b(s_208), .O(gate401inter1));
  and2  gate2005(.a(G1078), .b(G15), .O(gate401inter2));
  inv1  gate2006(.a(s_208), .O(gate401inter3));
  inv1  gate2007(.a(s_209), .O(gate401inter4));
  nand2 gate2008(.a(gate401inter4), .b(gate401inter3), .O(gate401inter5));
  nor2  gate2009(.a(gate401inter5), .b(gate401inter2), .O(gate401inter6));
  inv1  gate2010(.a(G15), .O(gate401inter7));
  inv1  gate2011(.a(G1078), .O(gate401inter8));
  nand2 gate2012(.a(gate401inter8), .b(gate401inter7), .O(gate401inter9));
  nand2 gate2013(.a(s_209), .b(gate401inter3), .O(gate401inter10));
  nor2  gate2014(.a(gate401inter10), .b(gate401inter9), .O(gate401inter11));
  nor2  gate2015(.a(gate401inter11), .b(gate401inter6), .O(gate401inter12));
  nand2 gate2016(.a(gate401inter12), .b(gate401inter1), .O(G1174));
nand2 gate402( .a(G16), .b(G1081), .O(G1177) );

  xor2  gate1051(.a(G1084), .b(G17), .O(gate403inter0));
  nand2 gate1052(.a(gate403inter0), .b(s_72), .O(gate403inter1));
  and2  gate1053(.a(G1084), .b(G17), .O(gate403inter2));
  inv1  gate1054(.a(s_72), .O(gate403inter3));
  inv1  gate1055(.a(s_73), .O(gate403inter4));
  nand2 gate1056(.a(gate403inter4), .b(gate403inter3), .O(gate403inter5));
  nor2  gate1057(.a(gate403inter5), .b(gate403inter2), .O(gate403inter6));
  inv1  gate1058(.a(G17), .O(gate403inter7));
  inv1  gate1059(.a(G1084), .O(gate403inter8));
  nand2 gate1060(.a(gate403inter8), .b(gate403inter7), .O(gate403inter9));
  nand2 gate1061(.a(s_73), .b(gate403inter3), .O(gate403inter10));
  nor2  gate1062(.a(gate403inter10), .b(gate403inter9), .O(gate403inter11));
  nor2  gate1063(.a(gate403inter11), .b(gate403inter6), .O(gate403inter12));
  nand2 gate1064(.a(gate403inter12), .b(gate403inter1), .O(G1180));
nand2 gate404( .a(G18), .b(G1087), .O(G1183) );
nand2 gate405( .a(G19), .b(G1090), .O(G1186) );

  xor2  gate2339(.a(G1093), .b(G20), .O(gate406inter0));
  nand2 gate2340(.a(gate406inter0), .b(s_256), .O(gate406inter1));
  and2  gate2341(.a(G1093), .b(G20), .O(gate406inter2));
  inv1  gate2342(.a(s_256), .O(gate406inter3));
  inv1  gate2343(.a(s_257), .O(gate406inter4));
  nand2 gate2344(.a(gate406inter4), .b(gate406inter3), .O(gate406inter5));
  nor2  gate2345(.a(gate406inter5), .b(gate406inter2), .O(gate406inter6));
  inv1  gate2346(.a(G20), .O(gate406inter7));
  inv1  gate2347(.a(G1093), .O(gate406inter8));
  nand2 gate2348(.a(gate406inter8), .b(gate406inter7), .O(gate406inter9));
  nand2 gate2349(.a(s_257), .b(gate406inter3), .O(gate406inter10));
  nor2  gate2350(.a(gate406inter10), .b(gate406inter9), .O(gate406inter11));
  nor2  gate2351(.a(gate406inter11), .b(gate406inter6), .O(gate406inter12));
  nand2 gate2352(.a(gate406inter12), .b(gate406inter1), .O(G1189));

  xor2  gate1205(.a(G1096), .b(G21), .O(gate407inter0));
  nand2 gate1206(.a(gate407inter0), .b(s_94), .O(gate407inter1));
  and2  gate1207(.a(G1096), .b(G21), .O(gate407inter2));
  inv1  gate1208(.a(s_94), .O(gate407inter3));
  inv1  gate1209(.a(s_95), .O(gate407inter4));
  nand2 gate1210(.a(gate407inter4), .b(gate407inter3), .O(gate407inter5));
  nor2  gate1211(.a(gate407inter5), .b(gate407inter2), .O(gate407inter6));
  inv1  gate1212(.a(G21), .O(gate407inter7));
  inv1  gate1213(.a(G1096), .O(gate407inter8));
  nand2 gate1214(.a(gate407inter8), .b(gate407inter7), .O(gate407inter9));
  nand2 gate1215(.a(s_95), .b(gate407inter3), .O(gate407inter10));
  nor2  gate1216(.a(gate407inter10), .b(gate407inter9), .O(gate407inter11));
  nor2  gate1217(.a(gate407inter11), .b(gate407inter6), .O(gate407inter12));
  nand2 gate1218(.a(gate407inter12), .b(gate407inter1), .O(G1192));

  xor2  gate1177(.a(G1099), .b(G22), .O(gate408inter0));
  nand2 gate1178(.a(gate408inter0), .b(s_90), .O(gate408inter1));
  and2  gate1179(.a(G1099), .b(G22), .O(gate408inter2));
  inv1  gate1180(.a(s_90), .O(gate408inter3));
  inv1  gate1181(.a(s_91), .O(gate408inter4));
  nand2 gate1182(.a(gate408inter4), .b(gate408inter3), .O(gate408inter5));
  nor2  gate1183(.a(gate408inter5), .b(gate408inter2), .O(gate408inter6));
  inv1  gate1184(.a(G22), .O(gate408inter7));
  inv1  gate1185(.a(G1099), .O(gate408inter8));
  nand2 gate1186(.a(gate408inter8), .b(gate408inter7), .O(gate408inter9));
  nand2 gate1187(.a(s_91), .b(gate408inter3), .O(gate408inter10));
  nor2  gate1188(.a(gate408inter10), .b(gate408inter9), .O(gate408inter11));
  nor2  gate1189(.a(gate408inter11), .b(gate408inter6), .O(gate408inter12));
  nand2 gate1190(.a(gate408inter12), .b(gate408inter1), .O(G1195));
nand2 gate409( .a(G23), .b(G1102), .O(G1198) );
nand2 gate410( .a(G24), .b(G1105), .O(G1201) );

  xor2  gate939(.a(G1108), .b(G25), .O(gate411inter0));
  nand2 gate940(.a(gate411inter0), .b(s_56), .O(gate411inter1));
  and2  gate941(.a(G1108), .b(G25), .O(gate411inter2));
  inv1  gate942(.a(s_56), .O(gate411inter3));
  inv1  gate943(.a(s_57), .O(gate411inter4));
  nand2 gate944(.a(gate411inter4), .b(gate411inter3), .O(gate411inter5));
  nor2  gate945(.a(gate411inter5), .b(gate411inter2), .O(gate411inter6));
  inv1  gate946(.a(G25), .O(gate411inter7));
  inv1  gate947(.a(G1108), .O(gate411inter8));
  nand2 gate948(.a(gate411inter8), .b(gate411inter7), .O(gate411inter9));
  nand2 gate949(.a(s_57), .b(gate411inter3), .O(gate411inter10));
  nor2  gate950(.a(gate411inter10), .b(gate411inter9), .O(gate411inter11));
  nor2  gate951(.a(gate411inter11), .b(gate411inter6), .O(gate411inter12));
  nand2 gate952(.a(gate411inter12), .b(gate411inter1), .O(G1204));
nand2 gate412( .a(G26), .b(G1111), .O(G1207) );

  xor2  gate1821(.a(G1114), .b(G27), .O(gate413inter0));
  nand2 gate1822(.a(gate413inter0), .b(s_182), .O(gate413inter1));
  and2  gate1823(.a(G1114), .b(G27), .O(gate413inter2));
  inv1  gate1824(.a(s_182), .O(gate413inter3));
  inv1  gate1825(.a(s_183), .O(gate413inter4));
  nand2 gate1826(.a(gate413inter4), .b(gate413inter3), .O(gate413inter5));
  nor2  gate1827(.a(gate413inter5), .b(gate413inter2), .O(gate413inter6));
  inv1  gate1828(.a(G27), .O(gate413inter7));
  inv1  gate1829(.a(G1114), .O(gate413inter8));
  nand2 gate1830(.a(gate413inter8), .b(gate413inter7), .O(gate413inter9));
  nand2 gate1831(.a(s_183), .b(gate413inter3), .O(gate413inter10));
  nor2  gate1832(.a(gate413inter10), .b(gate413inter9), .O(gate413inter11));
  nor2  gate1833(.a(gate413inter11), .b(gate413inter6), .O(gate413inter12));
  nand2 gate1834(.a(gate413inter12), .b(gate413inter1), .O(G1210));

  xor2  gate2899(.a(G1117), .b(G28), .O(gate414inter0));
  nand2 gate2900(.a(gate414inter0), .b(s_336), .O(gate414inter1));
  and2  gate2901(.a(G1117), .b(G28), .O(gate414inter2));
  inv1  gate2902(.a(s_336), .O(gate414inter3));
  inv1  gate2903(.a(s_337), .O(gate414inter4));
  nand2 gate2904(.a(gate414inter4), .b(gate414inter3), .O(gate414inter5));
  nor2  gate2905(.a(gate414inter5), .b(gate414inter2), .O(gate414inter6));
  inv1  gate2906(.a(G28), .O(gate414inter7));
  inv1  gate2907(.a(G1117), .O(gate414inter8));
  nand2 gate2908(.a(gate414inter8), .b(gate414inter7), .O(gate414inter9));
  nand2 gate2909(.a(s_337), .b(gate414inter3), .O(gate414inter10));
  nor2  gate2910(.a(gate414inter10), .b(gate414inter9), .O(gate414inter11));
  nor2  gate2911(.a(gate414inter11), .b(gate414inter6), .O(gate414inter12));
  nand2 gate2912(.a(gate414inter12), .b(gate414inter1), .O(G1213));
nand2 gate415( .a(G29), .b(G1120), .O(G1216) );
nand2 gate416( .a(G30), .b(G1123), .O(G1219) );
nand2 gate417( .a(G31), .b(G1126), .O(G1222) );
nand2 gate418( .a(G32), .b(G1129), .O(G1225) );
nand2 gate419( .a(G1), .b(G1132), .O(G1228) );

  xor2  gate2171(.a(G1132), .b(G1036), .O(gate420inter0));
  nand2 gate2172(.a(gate420inter0), .b(s_232), .O(gate420inter1));
  and2  gate2173(.a(G1132), .b(G1036), .O(gate420inter2));
  inv1  gate2174(.a(s_232), .O(gate420inter3));
  inv1  gate2175(.a(s_233), .O(gate420inter4));
  nand2 gate2176(.a(gate420inter4), .b(gate420inter3), .O(gate420inter5));
  nor2  gate2177(.a(gate420inter5), .b(gate420inter2), .O(gate420inter6));
  inv1  gate2178(.a(G1036), .O(gate420inter7));
  inv1  gate2179(.a(G1132), .O(gate420inter8));
  nand2 gate2180(.a(gate420inter8), .b(gate420inter7), .O(gate420inter9));
  nand2 gate2181(.a(s_233), .b(gate420inter3), .O(gate420inter10));
  nor2  gate2182(.a(gate420inter10), .b(gate420inter9), .O(gate420inter11));
  nor2  gate2183(.a(gate420inter11), .b(gate420inter6), .O(gate420inter12));
  nand2 gate2184(.a(gate420inter12), .b(gate420inter1), .O(G1229));

  xor2  gate2367(.a(G1135), .b(G2), .O(gate421inter0));
  nand2 gate2368(.a(gate421inter0), .b(s_260), .O(gate421inter1));
  and2  gate2369(.a(G1135), .b(G2), .O(gate421inter2));
  inv1  gate2370(.a(s_260), .O(gate421inter3));
  inv1  gate2371(.a(s_261), .O(gate421inter4));
  nand2 gate2372(.a(gate421inter4), .b(gate421inter3), .O(gate421inter5));
  nor2  gate2373(.a(gate421inter5), .b(gate421inter2), .O(gate421inter6));
  inv1  gate2374(.a(G2), .O(gate421inter7));
  inv1  gate2375(.a(G1135), .O(gate421inter8));
  nand2 gate2376(.a(gate421inter8), .b(gate421inter7), .O(gate421inter9));
  nand2 gate2377(.a(s_261), .b(gate421inter3), .O(gate421inter10));
  nor2  gate2378(.a(gate421inter10), .b(gate421inter9), .O(gate421inter11));
  nor2  gate2379(.a(gate421inter11), .b(gate421inter6), .O(gate421inter12));
  nand2 gate2380(.a(gate421inter12), .b(gate421inter1), .O(G1230));

  xor2  gate1989(.a(G1135), .b(G1039), .O(gate422inter0));
  nand2 gate1990(.a(gate422inter0), .b(s_206), .O(gate422inter1));
  and2  gate1991(.a(G1135), .b(G1039), .O(gate422inter2));
  inv1  gate1992(.a(s_206), .O(gate422inter3));
  inv1  gate1993(.a(s_207), .O(gate422inter4));
  nand2 gate1994(.a(gate422inter4), .b(gate422inter3), .O(gate422inter5));
  nor2  gate1995(.a(gate422inter5), .b(gate422inter2), .O(gate422inter6));
  inv1  gate1996(.a(G1039), .O(gate422inter7));
  inv1  gate1997(.a(G1135), .O(gate422inter8));
  nand2 gate1998(.a(gate422inter8), .b(gate422inter7), .O(gate422inter9));
  nand2 gate1999(.a(s_207), .b(gate422inter3), .O(gate422inter10));
  nor2  gate2000(.a(gate422inter10), .b(gate422inter9), .O(gate422inter11));
  nor2  gate2001(.a(gate422inter11), .b(gate422inter6), .O(gate422inter12));
  nand2 gate2002(.a(gate422inter12), .b(gate422inter1), .O(G1231));
nand2 gate423( .a(G3), .b(G1138), .O(G1232) );

  xor2  gate1023(.a(G1138), .b(G1042), .O(gate424inter0));
  nand2 gate1024(.a(gate424inter0), .b(s_68), .O(gate424inter1));
  and2  gate1025(.a(G1138), .b(G1042), .O(gate424inter2));
  inv1  gate1026(.a(s_68), .O(gate424inter3));
  inv1  gate1027(.a(s_69), .O(gate424inter4));
  nand2 gate1028(.a(gate424inter4), .b(gate424inter3), .O(gate424inter5));
  nor2  gate1029(.a(gate424inter5), .b(gate424inter2), .O(gate424inter6));
  inv1  gate1030(.a(G1042), .O(gate424inter7));
  inv1  gate1031(.a(G1138), .O(gate424inter8));
  nand2 gate1032(.a(gate424inter8), .b(gate424inter7), .O(gate424inter9));
  nand2 gate1033(.a(s_69), .b(gate424inter3), .O(gate424inter10));
  nor2  gate1034(.a(gate424inter10), .b(gate424inter9), .O(gate424inter11));
  nor2  gate1035(.a(gate424inter11), .b(gate424inter6), .O(gate424inter12));
  nand2 gate1036(.a(gate424inter12), .b(gate424inter1), .O(G1233));
nand2 gate425( .a(G4), .b(G1141), .O(G1234) );
nand2 gate426( .a(G1045), .b(G1141), .O(G1235) );
nand2 gate427( .a(G5), .b(G1144), .O(G1236) );

  xor2  gate2045(.a(G1144), .b(G1048), .O(gate428inter0));
  nand2 gate2046(.a(gate428inter0), .b(s_214), .O(gate428inter1));
  and2  gate2047(.a(G1144), .b(G1048), .O(gate428inter2));
  inv1  gate2048(.a(s_214), .O(gate428inter3));
  inv1  gate2049(.a(s_215), .O(gate428inter4));
  nand2 gate2050(.a(gate428inter4), .b(gate428inter3), .O(gate428inter5));
  nor2  gate2051(.a(gate428inter5), .b(gate428inter2), .O(gate428inter6));
  inv1  gate2052(.a(G1048), .O(gate428inter7));
  inv1  gate2053(.a(G1144), .O(gate428inter8));
  nand2 gate2054(.a(gate428inter8), .b(gate428inter7), .O(gate428inter9));
  nand2 gate2055(.a(s_215), .b(gate428inter3), .O(gate428inter10));
  nor2  gate2056(.a(gate428inter10), .b(gate428inter9), .O(gate428inter11));
  nor2  gate2057(.a(gate428inter11), .b(gate428inter6), .O(gate428inter12));
  nand2 gate2058(.a(gate428inter12), .b(gate428inter1), .O(G1237));

  xor2  gate1163(.a(G1147), .b(G6), .O(gate429inter0));
  nand2 gate1164(.a(gate429inter0), .b(s_88), .O(gate429inter1));
  and2  gate1165(.a(G1147), .b(G6), .O(gate429inter2));
  inv1  gate1166(.a(s_88), .O(gate429inter3));
  inv1  gate1167(.a(s_89), .O(gate429inter4));
  nand2 gate1168(.a(gate429inter4), .b(gate429inter3), .O(gate429inter5));
  nor2  gate1169(.a(gate429inter5), .b(gate429inter2), .O(gate429inter6));
  inv1  gate1170(.a(G6), .O(gate429inter7));
  inv1  gate1171(.a(G1147), .O(gate429inter8));
  nand2 gate1172(.a(gate429inter8), .b(gate429inter7), .O(gate429inter9));
  nand2 gate1173(.a(s_89), .b(gate429inter3), .O(gate429inter10));
  nor2  gate1174(.a(gate429inter10), .b(gate429inter9), .O(gate429inter11));
  nor2  gate1175(.a(gate429inter11), .b(gate429inter6), .O(gate429inter12));
  nand2 gate1176(.a(gate429inter12), .b(gate429inter1), .O(G1238));
nand2 gate430( .a(G1051), .b(G1147), .O(G1239) );
nand2 gate431( .a(G7), .b(G1150), .O(G1240) );
nand2 gate432( .a(G1054), .b(G1150), .O(G1241) );

  xor2  gate2591(.a(G1153), .b(G8), .O(gate433inter0));
  nand2 gate2592(.a(gate433inter0), .b(s_292), .O(gate433inter1));
  and2  gate2593(.a(G1153), .b(G8), .O(gate433inter2));
  inv1  gate2594(.a(s_292), .O(gate433inter3));
  inv1  gate2595(.a(s_293), .O(gate433inter4));
  nand2 gate2596(.a(gate433inter4), .b(gate433inter3), .O(gate433inter5));
  nor2  gate2597(.a(gate433inter5), .b(gate433inter2), .O(gate433inter6));
  inv1  gate2598(.a(G8), .O(gate433inter7));
  inv1  gate2599(.a(G1153), .O(gate433inter8));
  nand2 gate2600(.a(gate433inter8), .b(gate433inter7), .O(gate433inter9));
  nand2 gate2601(.a(s_293), .b(gate433inter3), .O(gate433inter10));
  nor2  gate2602(.a(gate433inter10), .b(gate433inter9), .O(gate433inter11));
  nor2  gate2603(.a(gate433inter11), .b(gate433inter6), .O(gate433inter12));
  nand2 gate2604(.a(gate433inter12), .b(gate433inter1), .O(G1242));

  xor2  gate2353(.a(G1153), .b(G1057), .O(gate434inter0));
  nand2 gate2354(.a(gate434inter0), .b(s_258), .O(gate434inter1));
  and2  gate2355(.a(G1153), .b(G1057), .O(gate434inter2));
  inv1  gate2356(.a(s_258), .O(gate434inter3));
  inv1  gate2357(.a(s_259), .O(gate434inter4));
  nand2 gate2358(.a(gate434inter4), .b(gate434inter3), .O(gate434inter5));
  nor2  gate2359(.a(gate434inter5), .b(gate434inter2), .O(gate434inter6));
  inv1  gate2360(.a(G1057), .O(gate434inter7));
  inv1  gate2361(.a(G1153), .O(gate434inter8));
  nand2 gate2362(.a(gate434inter8), .b(gate434inter7), .O(gate434inter9));
  nand2 gate2363(.a(s_259), .b(gate434inter3), .O(gate434inter10));
  nor2  gate2364(.a(gate434inter10), .b(gate434inter9), .O(gate434inter11));
  nor2  gate2365(.a(gate434inter11), .b(gate434inter6), .O(gate434inter12));
  nand2 gate2366(.a(gate434inter12), .b(gate434inter1), .O(G1243));
nand2 gate435( .a(G9), .b(G1156), .O(G1244) );
nand2 gate436( .a(G1060), .b(G1156), .O(G1245) );
nand2 gate437( .a(G10), .b(G1159), .O(G1246) );
nand2 gate438( .a(G1063), .b(G1159), .O(G1247) );
nand2 gate439( .a(G11), .b(G1162), .O(G1248) );
nand2 gate440( .a(G1066), .b(G1162), .O(G1249) );
nand2 gate441( .a(G12), .b(G1165), .O(G1250) );

  xor2  gate1149(.a(G1165), .b(G1069), .O(gate442inter0));
  nand2 gate1150(.a(gate442inter0), .b(s_86), .O(gate442inter1));
  and2  gate1151(.a(G1165), .b(G1069), .O(gate442inter2));
  inv1  gate1152(.a(s_86), .O(gate442inter3));
  inv1  gate1153(.a(s_87), .O(gate442inter4));
  nand2 gate1154(.a(gate442inter4), .b(gate442inter3), .O(gate442inter5));
  nor2  gate1155(.a(gate442inter5), .b(gate442inter2), .O(gate442inter6));
  inv1  gate1156(.a(G1069), .O(gate442inter7));
  inv1  gate1157(.a(G1165), .O(gate442inter8));
  nand2 gate1158(.a(gate442inter8), .b(gate442inter7), .O(gate442inter9));
  nand2 gate1159(.a(s_87), .b(gate442inter3), .O(gate442inter10));
  nor2  gate1160(.a(gate442inter10), .b(gate442inter9), .O(gate442inter11));
  nor2  gate1161(.a(gate442inter11), .b(gate442inter6), .O(gate442inter12));
  nand2 gate1162(.a(gate442inter12), .b(gate442inter1), .O(G1251));
nand2 gate443( .a(G13), .b(G1168), .O(G1252) );

  xor2  gate2871(.a(G1168), .b(G1072), .O(gate444inter0));
  nand2 gate2872(.a(gate444inter0), .b(s_332), .O(gate444inter1));
  and2  gate2873(.a(G1168), .b(G1072), .O(gate444inter2));
  inv1  gate2874(.a(s_332), .O(gate444inter3));
  inv1  gate2875(.a(s_333), .O(gate444inter4));
  nand2 gate2876(.a(gate444inter4), .b(gate444inter3), .O(gate444inter5));
  nor2  gate2877(.a(gate444inter5), .b(gate444inter2), .O(gate444inter6));
  inv1  gate2878(.a(G1072), .O(gate444inter7));
  inv1  gate2879(.a(G1168), .O(gate444inter8));
  nand2 gate2880(.a(gate444inter8), .b(gate444inter7), .O(gate444inter9));
  nand2 gate2881(.a(s_333), .b(gate444inter3), .O(gate444inter10));
  nor2  gate2882(.a(gate444inter10), .b(gate444inter9), .O(gate444inter11));
  nor2  gate2883(.a(gate444inter11), .b(gate444inter6), .O(gate444inter12));
  nand2 gate2884(.a(gate444inter12), .b(gate444inter1), .O(G1253));
nand2 gate445( .a(G14), .b(G1171), .O(G1254) );
nand2 gate446( .a(G1075), .b(G1171), .O(G1255) );

  xor2  gate841(.a(G1174), .b(G15), .O(gate447inter0));
  nand2 gate842(.a(gate447inter0), .b(s_42), .O(gate447inter1));
  and2  gate843(.a(G1174), .b(G15), .O(gate447inter2));
  inv1  gate844(.a(s_42), .O(gate447inter3));
  inv1  gate845(.a(s_43), .O(gate447inter4));
  nand2 gate846(.a(gate447inter4), .b(gate447inter3), .O(gate447inter5));
  nor2  gate847(.a(gate447inter5), .b(gate447inter2), .O(gate447inter6));
  inv1  gate848(.a(G15), .O(gate447inter7));
  inv1  gate849(.a(G1174), .O(gate447inter8));
  nand2 gate850(.a(gate447inter8), .b(gate447inter7), .O(gate447inter9));
  nand2 gate851(.a(s_43), .b(gate447inter3), .O(gate447inter10));
  nor2  gate852(.a(gate447inter10), .b(gate447inter9), .O(gate447inter11));
  nor2  gate853(.a(gate447inter11), .b(gate447inter6), .O(gate447inter12));
  nand2 gate854(.a(gate447inter12), .b(gate447inter1), .O(G1256));

  xor2  gate2493(.a(G1174), .b(G1078), .O(gate448inter0));
  nand2 gate2494(.a(gate448inter0), .b(s_278), .O(gate448inter1));
  and2  gate2495(.a(G1174), .b(G1078), .O(gate448inter2));
  inv1  gate2496(.a(s_278), .O(gate448inter3));
  inv1  gate2497(.a(s_279), .O(gate448inter4));
  nand2 gate2498(.a(gate448inter4), .b(gate448inter3), .O(gate448inter5));
  nor2  gate2499(.a(gate448inter5), .b(gate448inter2), .O(gate448inter6));
  inv1  gate2500(.a(G1078), .O(gate448inter7));
  inv1  gate2501(.a(G1174), .O(gate448inter8));
  nand2 gate2502(.a(gate448inter8), .b(gate448inter7), .O(gate448inter9));
  nand2 gate2503(.a(s_279), .b(gate448inter3), .O(gate448inter10));
  nor2  gate2504(.a(gate448inter10), .b(gate448inter9), .O(gate448inter11));
  nor2  gate2505(.a(gate448inter11), .b(gate448inter6), .O(gate448inter12));
  nand2 gate2506(.a(gate448inter12), .b(gate448inter1), .O(G1257));

  xor2  gate2787(.a(G1177), .b(G16), .O(gate449inter0));
  nand2 gate2788(.a(gate449inter0), .b(s_320), .O(gate449inter1));
  and2  gate2789(.a(G1177), .b(G16), .O(gate449inter2));
  inv1  gate2790(.a(s_320), .O(gate449inter3));
  inv1  gate2791(.a(s_321), .O(gate449inter4));
  nand2 gate2792(.a(gate449inter4), .b(gate449inter3), .O(gate449inter5));
  nor2  gate2793(.a(gate449inter5), .b(gate449inter2), .O(gate449inter6));
  inv1  gate2794(.a(G16), .O(gate449inter7));
  inv1  gate2795(.a(G1177), .O(gate449inter8));
  nand2 gate2796(.a(gate449inter8), .b(gate449inter7), .O(gate449inter9));
  nand2 gate2797(.a(s_321), .b(gate449inter3), .O(gate449inter10));
  nor2  gate2798(.a(gate449inter10), .b(gate449inter9), .O(gate449inter11));
  nor2  gate2799(.a(gate449inter11), .b(gate449inter6), .O(gate449inter12));
  nand2 gate2800(.a(gate449inter12), .b(gate449inter1), .O(G1258));
nand2 gate450( .a(G1081), .b(G1177), .O(G1259) );
nand2 gate451( .a(G17), .b(G1180), .O(G1260) );

  xor2  gate1877(.a(G1180), .b(G1084), .O(gate452inter0));
  nand2 gate1878(.a(gate452inter0), .b(s_190), .O(gate452inter1));
  and2  gate1879(.a(G1180), .b(G1084), .O(gate452inter2));
  inv1  gate1880(.a(s_190), .O(gate452inter3));
  inv1  gate1881(.a(s_191), .O(gate452inter4));
  nand2 gate1882(.a(gate452inter4), .b(gate452inter3), .O(gate452inter5));
  nor2  gate1883(.a(gate452inter5), .b(gate452inter2), .O(gate452inter6));
  inv1  gate1884(.a(G1084), .O(gate452inter7));
  inv1  gate1885(.a(G1180), .O(gate452inter8));
  nand2 gate1886(.a(gate452inter8), .b(gate452inter7), .O(gate452inter9));
  nand2 gate1887(.a(s_191), .b(gate452inter3), .O(gate452inter10));
  nor2  gate1888(.a(gate452inter10), .b(gate452inter9), .O(gate452inter11));
  nor2  gate1889(.a(gate452inter11), .b(gate452inter6), .O(gate452inter12));
  nand2 gate1890(.a(gate452inter12), .b(gate452inter1), .O(G1261));

  xor2  gate561(.a(G1183), .b(G18), .O(gate453inter0));
  nand2 gate562(.a(gate453inter0), .b(s_2), .O(gate453inter1));
  and2  gate563(.a(G1183), .b(G18), .O(gate453inter2));
  inv1  gate564(.a(s_2), .O(gate453inter3));
  inv1  gate565(.a(s_3), .O(gate453inter4));
  nand2 gate566(.a(gate453inter4), .b(gate453inter3), .O(gate453inter5));
  nor2  gate567(.a(gate453inter5), .b(gate453inter2), .O(gate453inter6));
  inv1  gate568(.a(G18), .O(gate453inter7));
  inv1  gate569(.a(G1183), .O(gate453inter8));
  nand2 gate570(.a(gate453inter8), .b(gate453inter7), .O(gate453inter9));
  nand2 gate571(.a(s_3), .b(gate453inter3), .O(gate453inter10));
  nor2  gate572(.a(gate453inter10), .b(gate453inter9), .O(gate453inter11));
  nor2  gate573(.a(gate453inter11), .b(gate453inter6), .O(gate453inter12));
  nand2 gate574(.a(gate453inter12), .b(gate453inter1), .O(G1262));

  xor2  gate799(.a(G1183), .b(G1087), .O(gate454inter0));
  nand2 gate800(.a(gate454inter0), .b(s_36), .O(gate454inter1));
  and2  gate801(.a(G1183), .b(G1087), .O(gate454inter2));
  inv1  gate802(.a(s_36), .O(gate454inter3));
  inv1  gate803(.a(s_37), .O(gate454inter4));
  nand2 gate804(.a(gate454inter4), .b(gate454inter3), .O(gate454inter5));
  nor2  gate805(.a(gate454inter5), .b(gate454inter2), .O(gate454inter6));
  inv1  gate806(.a(G1087), .O(gate454inter7));
  inv1  gate807(.a(G1183), .O(gate454inter8));
  nand2 gate808(.a(gate454inter8), .b(gate454inter7), .O(gate454inter9));
  nand2 gate809(.a(s_37), .b(gate454inter3), .O(gate454inter10));
  nor2  gate810(.a(gate454inter10), .b(gate454inter9), .O(gate454inter11));
  nor2  gate811(.a(gate454inter11), .b(gate454inter6), .O(gate454inter12));
  nand2 gate812(.a(gate454inter12), .b(gate454inter1), .O(G1263));
nand2 gate455( .a(G19), .b(G1186), .O(G1264) );
nand2 gate456( .a(G1090), .b(G1186), .O(G1265) );
nand2 gate457( .a(G20), .b(G1189), .O(G1266) );
nand2 gate458( .a(G1093), .b(G1189), .O(G1267) );
nand2 gate459( .a(G21), .b(G1192), .O(G1268) );
nand2 gate460( .a(G1096), .b(G1192), .O(G1269) );
nand2 gate461( .a(G22), .b(G1195), .O(G1270) );
nand2 gate462( .a(G1099), .b(G1195), .O(G1271) );
nand2 gate463( .a(G23), .b(G1198), .O(G1272) );
nand2 gate464( .a(G1102), .b(G1198), .O(G1273) );
nand2 gate465( .a(G24), .b(G1201), .O(G1274) );
nand2 gate466( .a(G1105), .b(G1201), .O(G1275) );

  xor2  gate2087(.a(G1204), .b(G25), .O(gate467inter0));
  nand2 gate2088(.a(gate467inter0), .b(s_220), .O(gate467inter1));
  and2  gate2089(.a(G1204), .b(G25), .O(gate467inter2));
  inv1  gate2090(.a(s_220), .O(gate467inter3));
  inv1  gate2091(.a(s_221), .O(gate467inter4));
  nand2 gate2092(.a(gate467inter4), .b(gate467inter3), .O(gate467inter5));
  nor2  gate2093(.a(gate467inter5), .b(gate467inter2), .O(gate467inter6));
  inv1  gate2094(.a(G25), .O(gate467inter7));
  inv1  gate2095(.a(G1204), .O(gate467inter8));
  nand2 gate2096(.a(gate467inter8), .b(gate467inter7), .O(gate467inter9));
  nand2 gate2097(.a(s_221), .b(gate467inter3), .O(gate467inter10));
  nor2  gate2098(.a(gate467inter10), .b(gate467inter9), .O(gate467inter11));
  nor2  gate2099(.a(gate467inter11), .b(gate467inter6), .O(gate467inter12));
  nand2 gate2100(.a(gate467inter12), .b(gate467inter1), .O(G1276));
nand2 gate468( .a(G1108), .b(G1204), .O(G1277) );

  xor2  gate2577(.a(G1207), .b(G26), .O(gate469inter0));
  nand2 gate2578(.a(gate469inter0), .b(s_290), .O(gate469inter1));
  and2  gate2579(.a(G1207), .b(G26), .O(gate469inter2));
  inv1  gate2580(.a(s_290), .O(gate469inter3));
  inv1  gate2581(.a(s_291), .O(gate469inter4));
  nand2 gate2582(.a(gate469inter4), .b(gate469inter3), .O(gate469inter5));
  nor2  gate2583(.a(gate469inter5), .b(gate469inter2), .O(gate469inter6));
  inv1  gate2584(.a(G26), .O(gate469inter7));
  inv1  gate2585(.a(G1207), .O(gate469inter8));
  nand2 gate2586(.a(gate469inter8), .b(gate469inter7), .O(gate469inter9));
  nand2 gate2587(.a(s_291), .b(gate469inter3), .O(gate469inter10));
  nor2  gate2588(.a(gate469inter10), .b(gate469inter9), .O(gate469inter11));
  nor2  gate2589(.a(gate469inter11), .b(gate469inter6), .O(gate469inter12));
  nand2 gate2590(.a(gate469inter12), .b(gate469inter1), .O(G1278));

  xor2  gate2115(.a(G1207), .b(G1111), .O(gate470inter0));
  nand2 gate2116(.a(gate470inter0), .b(s_224), .O(gate470inter1));
  and2  gate2117(.a(G1207), .b(G1111), .O(gate470inter2));
  inv1  gate2118(.a(s_224), .O(gate470inter3));
  inv1  gate2119(.a(s_225), .O(gate470inter4));
  nand2 gate2120(.a(gate470inter4), .b(gate470inter3), .O(gate470inter5));
  nor2  gate2121(.a(gate470inter5), .b(gate470inter2), .O(gate470inter6));
  inv1  gate2122(.a(G1111), .O(gate470inter7));
  inv1  gate2123(.a(G1207), .O(gate470inter8));
  nand2 gate2124(.a(gate470inter8), .b(gate470inter7), .O(gate470inter9));
  nand2 gate2125(.a(s_225), .b(gate470inter3), .O(gate470inter10));
  nor2  gate2126(.a(gate470inter10), .b(gate470inter9), .O(gate470inter11));
  nor2  gate2127(.a(gate470inter11), .b(gate470inter6), .O(gate470inter12));
  nand2 gate2128(.a(gate470inter12), .b(gate470inter1), .O(G1279));
nand2 gate471( .a(G27), .b(G1210), .O(G1280) );
nand2 gate472( .a(G1114), .b(G1210), .O(G1281) );
nand2 gate473( .a(G28), .b(G1213), .O(G1282) );
nand2 gate474( .a(G1117), .b(G1213), .O(G1283) );
nand2 gate475( .a(G29), .b(G1216), .O(G1284) );
nand2 gate476( .a(G1120), .b(G1216), .O(G1285) );

  xor2  gate1765(.a(G1219), .b(G30), .O(gate477inter0));
  nand2 gate1766(.a(gate477inter0), .b(s_174), .O(gate477inter1));
  and2  gate1767(.a(G1219), .b(G30), .O(gate477inter2));
  inv1  gate1768(.a(s_174), .O(gate477inter3));
  inv1  gate1769(.a(s_175), .O(gate477inter4));
  nand2 gate1770(.a(gate477inter4), .b(gate477inter3), .O(gate477inter5));
  nor2  gate1771(.a(gate477inter5), .b(gate477inter2), .O(gate477inter6));
  inv1  gate1772(.a(G30), .O(gate477inter7));
  inv1  gate1773(.a(G1219), .O(gate477inter8));
  nand2 gate1774(.a(gate477inter8), .b(gate477inter7), .O(gate477inter9));
  nand2 gate1775(.a(s_175), .b(gate477inter3), .O(gate477inter10));
  nor2  gate1776(.a(gate477inter10), .b(gate477inter9), .O(gate477inter11));
  nor2  gate1777(.a(gate477inter11), .b(gate477inter6), .O(gate477inter12));
  nand2 gate1778(.a(gate477inter12), .b(gate477inter1), .O(G1286));
nand2 gate478( .a(G1123), .b(G1219), .O(G1287) );

  xor2  gate1849(.a(G1222), .b(G31), .O(gate479inter0));
  nand2 gate1850(.a(gate479inter0), .b(s_186), .O(gate479inter1));
  and2  gate1851(.a(G1222), .b(G31), .O(gate479inter2));
  inv1  gate1852(.a(s_186), .O(gate479inter3));
  inv1  gate1853(.a(s_187), .O(gate479inter4));
  nand2 gate1854(.a(gate479inter4), .b(gate479inter3), .O(gate479inter5));
  nor2  gate1855(.a(gate479inter5), .b(gate479inter2), .O(gate479inter6));
  inv1  gate1856(.a(G31), .O(gate479inter7));
  inv1  gate1857(.a(G1222), .O(gate479inter8));
  nand2 gate1858(.a(gate479inter8), .b(gate479inter7), .O(gate479inter9));
  nand2 gate1859(.a(s_187), .b(gate479inter3), .O(gate479inter10));
  nor2  gate1860(.a(gate479inter10), .b(gate479inter9), .O(gate479inter11));
  nor2  gate1861(.a(gate479inter11), .b(gate479inter6), .O(gate479inter12));
  nand2 gate1862(.a(gate479inter12), .b(gate479inter1), .O(G1288));
nand2 gate480( .a(G1126), .b(G1222), .O(G1289) );

  xor2  gate1261(.a(G1225), .b(G32), .O(gate481inter0));
  nand2 gate1262(.a(gate481inter0), .b(s_102), .O(gate481inter1));
  and2  gate1263(.a(G1225), .b(G32), .O(gate481inter2));
  inv1  gate1264(.a(s_102), .O(gate481inter3));
  inv1  gate1265(.a(s_103), .O(gate481inter4));
  nand2 gate1266(.a(gate481inter4), .b(gate481inter3), .O(gate481inter5));
  nor2  gate1267(.a(gate481inter5), .b(gate481inter2), .O(gate481inter6));
  inv1  gate1268(.a(G32), .O(gate481inter7));
  inv1  gate1269(.a(G1225), .O(gate481inter8));
  nand2 gate1270(.a(gate481inter8), .b(gate481inter7), .O(gate481inter9));
  nand2 gate1271(.a(s_103), .b(gate481inter3), .O(gate481inter10));
  nor2  gate1272(.a(gate481inter10), .b(gate481inter9), .O(gate481inter11));
  nor2  gate1273(.a(gate481inter11), .b(gate481inter6), .O(gate481inter12));
  nand2 gate1274(.a(gate481inter12), .b(gate481inter1), .O(G1290));

  xor2  gate2857(.a(G1225), .b(G1129), .O(gate482inter0));
  nand2 gate2858(.a(gate482inter0), .b(s_330), .O(gate482inter1));
  and2  gate2859(.a(G1225), .b(G1129), .O(gate482inter2));
  inv1  gate2860(.a(s_330), .O(gate482inter3));
  inv1  gate2861(.a(s_331), .O(gate482inter4));
  nand2 gate2862(.a(gate482inter4), .b(gate482inter3), .O(gate482inter5));
  nor2  gate2863(.a(gate482inter5), .b(gate482inter2), .O(gate482inter6));
  inv1  gate2864(.a(G1129), .O(gate482inter7));
  inv1  gate2865(.a(G1225), .O(gate482inter8));
  nand2 gate2866(.a(gate482inter8), .b(gate482inter7), .O(gate482inter9));
  nand2 gate2867(.a(s_331), .b(gate482inter3), .O(gate482inter10));
  nor2  gate2868(.a(gate482inter10), .b(gate482inter9), .O(gate482inter11));
  nor2  gate2869(.a(gate482inter11), .b(gate482inter6), .O(gate482inter12));
  nand2 gate2870(.a(gate482inter12), .b(gate482inter1), .O(G1291));

  xor2  gate925(.a(G1229), .b(G1228), .O(gate483inter0));
  nand2 gate926(.a(gate483inter0), .b(s_54), .O(gate483inter1));
  and2  gate927(.a(G1229), .b(G1228), .O(gate483inter2));
  inv1  gate928(.a(s_54), .O(gate483inter3));
  inv1  gate929(.a(s_55), .O(gate483inter4));
  nand2 gate930(.a(gate483inter4), .b(gate483inter3), .O(gate483inter5));
  nor2  gate931(.a(gate483inter5), .b(gate483inter2), .O(gate483inter6));
  inv1  gate932(.a(G1228), .O(gate483inter7));
  inv1  gate933(.a(G1229), .O(gate483inter8));
  nand2 gate934(.a(gate483inter8), .b(gate483inter7), .O(gate483inter9));
  nand2 gate935(.a(s_55), .b(gate483inter3), .O(gate483inter10));
  nor2  gate936(.a(gate483inter10), .b(gate483inter9), .O(gate483inter11));
  nor2  gate937(.a(gate483inter11), .b(gate483inter6), .O(gate483inter12));
  nand2 gate938(.a(gate483inter12), .b(gate483inter1), .O(G1292));

  xor2  gate1975(.a(G1231), .b(G1230), .O(gate484inter0));
  nand2 gate1976(.a(gate484inter0), .b(s_204), .O(gate484inter1));
  and2  gate1977(.a(G1231), .b(G1230), .O(gate484inter2));
  inv1  gate1978(.a(s_204), .O(gate484inter3));
  inv1  gate1979(.a(s_205), .O(gate484inter4));
  nand2 gate1980(.a(gate484inter4), .b(gate484inter3), .O(gate484inter5));
  nor2  gate1981(.a(gate484inter5), .b(gate484inter2), .O(gate484inter6));
  inv1  gate1982(.a(G1230), .O(gate484inter7));
  inv1  gate1983(.a(G1231), .O(gate484inter8));
  nand2 gate1984(.a(gate484inter8), .b(gate484inter7), .O(gate484inter9));
  nand2 gate1985(.a(s_205), .b(gate484inter3), .O(gate484inter10));
  nor2  gate1986(.a(gate484inter10), .b(gate484inter9), .O(gate484inter11));
  nor2  gate1987(.a(gate484inter11), .b(gate484inter6), .O(gate484inter12));
  nand2 gate1988(.a(gate484inter12), .b(gate484inter1), .O(G1293));

  xor2  gate2437(.a(G1233), .b(G1232), .O(gate485inter0));
  nand2 gate2438(.a(gate485inter0), .b(s_270), .O(gate485inter1));
  and2  gate2439(.a(G1233), .b(G1232), .O(gate485inter2));
  inv1  gate2440(.a(s_270), .O(gate485inter3));
  inv1  gate2441(.a(s_271), .O(gate485inter4));
  nand2 gate2442(.a(gate485inter4), .b(gate485inter3), .O(gate485inter5));
  nor2  gate2443(.a(gate485inter5), .b(gate485inter2), .O(gate485inter6));
  inv1  gate2444(.a(G1232), .O(gate485inter7));
  inv1  gate2445(.a(G1233), .O(gate485inter8));
  nand2 gate2446(.a(gate485inter8), .b(gate485inter7), .O(gate485inter9));
  nand2 gate2447(.a(s_271), .b(gate485inter3), .O(gate485inter10));
  nor2  gate2448(.a(gate485inter10), .b(gate485inter9), .O(gate485inter11));
  nor2  gate2449(.a(gate485inter11), .b(gate485inter6), .O(gate485inter12));
  nand2 gate2450(.a(gate485inter12), .b(gate485inter1), .O(G1294));
nand2 gate486( .a(G1234), .b(G1235), .O(G1295) );

  xor2  gate1513(.a(G1237), .b(G1236), .O(gate487inter0));
  nand2 gate1514(.a(gate487inter0), .b(s_138), .O(gate487inter1));
  and2  gate1515(.a(G1237), .b(G1236), .O(gate487inter2));
  inv1  gate1516(.a(s_138), .O(gate487inter3));
  inv1  gate1517(.a(s_139), .O(gate487inter4));
  nand2 gate1518(.a(gate487inter4), .b(gate487inter3), .O(gate487inter5));
  nor2  gate1519(.a(gate487inter5), .b(gate487inter2), .O(gate487inter6));
  inv1  gate1520(.a(G1236), .O(gate487inter7));
  inv1  gate1521(.a(G1237), .O(gate487inter8));
  nand2 gate1522(.a(gate487inter8), .b(gate487inter7), .O(gate487inter9));
  nand2 gate1523(.a(s_139), .b(gate487inter3), .O(gate487inter10));
  nor2  gate1524(.a(gate487inter10), .b(gate487inter9), .O(gate487inter11));
  nor2  gate1525(.a(gate487inter11), .b(gate487inter6), .O(gate487inter12));
  nand2 gate1526(.a(gate487inter12), .b(gate487inter1), .O(G1296));
nand2 gate488( .a(G1238), .b(G1239), .O(G1297) );
nand2 gate489( .a(G1240), .b(G1241), .O(G1298) );
nand2 gate490( .a(G1242), .b(G1243), .O(G1299) );

  xor2  gate617(.a(G1245), .b(G1244), .O(gate491inter0));
  nand2 gate618(.a(gate491inter0), .b(s_10), .O(gate491inter1));
  and2  gate619(.a(G1245), .b(G1244), .O(gate491inter2));
  inv1  gate620(.a(s_10), .O(gate491inter3));
  inv1  gate621(.a(s_11), .O(gate491inter4));
  nand2 gate622(.a(gate491inter4), .b(gate491inter3), .O(gate491inter5));
  nor2  gate623(.a(gate491inter5), .b(gate491inter2), .O(gate491inter6));
  inv1  gate624(.a(G1244), .O(gate491inter7));
  inv1  gate625(.a(G1245), .O(gate491inter8));
  nand2 gate626(.a(gate491inter8), .b(gate491inter7), .O(gate491inter9));
  nand2 gate627(.a(s_11), .b(gate491inter3), .O(gate491inter10));
  nor2  gate628(.a(gate491inter10), .b(gate491inter9), .O(gate491inter11));
  nor2  gate629(.a(gate491inter11), .b(gate491inter6), .O(gate491inter12));
  nand2 gate630(.a(gate491inter12), .b(gate491inter1), .O(G1300));
nand2 gate492( .a(G1246), .b(G1247), .O(G1301) );

  xor2  gate1947(.a(G1249), .b(G1248), .O(gate493inter0));
  nand2 gate1948(.a(gate493inter0), .b(s_200), .O(gate493inter1));
  and2  gate1949(.a(G1249), .b(G1248), .O(gate493inter2));
  inv1  gate1950(.a(s_200), .O(gate493inter3));
  inv1  gate1951(.a(s_201), .O(gate493inter4));
  nand2 gate1952(.a(gate493inter4), .b(gate493inter3), .O(gate493inter5));
  nor2  gate1953(.a(gate493inter5), .b(gate493inter2), .O(gate493inter6));
  inv1  gate1954(.a(G1248), .O(gate493inter7));
  inv1  gate1955(.a(G1249), .O(gate493inter8));
  nand2 gate1956(.a(gate493inter8), .b(gate493inter7), .O(gate493inter9));
  nand2 gate1957(.a(s_201), .b(gate493inter3), .O(gate493inter10));
  nor2  gate1958(.a(gate493inter10), .b(gate493inter9), .O(gate493inter11));
  nor2  gate1959(.a(gate493inter11), .b(gate493inter6), .O(gate493inter12));
  nand2 gate1960(.a(gate493inter12), .b(gate493inter1), .O(G1302));
nand2 gate494( .a(G1250), .b(G1251), .O(G1303) );

  xor2  gate1933(.a(G1253), .b(G1252), .O(gate495inter0));
  nand2 gate1934(.a(gate495inter0), .b(s_198), .O(gate495inter1));
  and2  gate1935(.a(G1253), .b(G1252), .O(gate495inter2));
  inv1  gate1936(.a(s_198), .O(gate495inter3));
  inv1  gate1937(.a(s_199), .O(gate495inter4));
  nand2 gate1938(.a(gate495inter4), .b(gate495inter3), .O(gate495inter5));
  nor2  gate1939(.a(gate495inter5), .b(gate495inter2), .O(gate495inter6));
  inv1  gate1940(.a(G1252), .O(gate495inter7));
  inv1  gate1941(.a(G1253), .O(gate495inter8));
  nand2 gate1942(.a(gate495inter8), .b(gate495inter7), .O(gate495inter9));
  nand2 gate1943(.a(s_199), .b(gate495inter3), .O(gate495inter10));
  nor2  gate1944(.a(gate495inter10), .b(gate495inter9), .O(gate495inter11));
  nor2  gate1945(.a(gate495inter11), .b(gate495inter6), .O(gate495inter12));
  nand2 gate1946(.a(gate495inter12), .b(gate495inter1), .O(G1304));
nand2 gate496( .a(G1254), .b(G1255), .O(G1305) );
nand2 gate497( .a(G1256), .b(G1257), .O(G1306) );
nand2 gate498( .a(G1258), .b(G1259), .O(G1307) );
nand2 gate499( .a(G1260), .b(G1261), .O(G1308) );
nand2 gate500( .a(G1262), .b(G1263), .O(G1309) );
nand2 gate501( .a(G1264), .b(G1265), .O(G1310) );

  xor2  gate673(.a(G1267), .b(G1266), .O(gate502inter0));
  nand2 gate674(.a(gate502inter0), .b(s_18), .O(gate502inter1));
  and2  gate675(.a(G1267), .b(G1266), .O(gate502inter2));
  inv1  gate676(.a(s_18), .O(gate502inter3));
  inv1  gate677(.a(s_19), .O(gate502inter4));
  nand2 gate678(.a(gate502inter4), .b(gate502inter3), .O(gate502inter5));
  nor2  gate679(.a(gate502inter5), .b(gate502inter2), .O(gate502inter6));
  inv1  gate680(.a(G1266), .O(gate502inter7));
  inv1  gate681(.a(G1267), .O(gate502inter8));
  nand2 gate682(.a(gate502inter8), .b(gate502inter7), .O(gate502inter9));
  nand2 gate683(.a(s_19), .b(gate502inter3), .O(gate502inter10));
  nor2  gate684(.a(gate502inter10), .b(gate502inter9), .O(gate502inter11));
  nor2  gate685(.a(gate502inter11), .b(gate502inter6), .O(gate502inter12));
  nand2 gate686(.a(gate502inter12), .b(gate502inter1), .O(G1311));
nand2 gate503( .a(G1268), .b(G1269), .O(G1312) );
nand2 gate504( .a(G1270), .b(G1271), .O(G1313) );
nand2 gate505( .a(G1272), .b(G1273), .O(G1314) );

  xor2  gate2465(.a(G1275), .b(G1274), .O(gate506inter0));
  nand2 gate2466(.a(gate506inter0), .b(s_274), .O(gate506inter1));
  and2  gate2467(.a(G1275), .b(G1274), .O(gate506inter2));
  inv1  gate2468(.a(s_274), .O(gate506inter3));
  inv1  gate2469(.a(s_275), .O(gate506inter4));
  nand2 gate2470(.a(gate506inter4), .b(gate506inter3), .O(gate506inter5));
  nor2  gate2471(.a(gate506inter5), .b(gate506inter2), .O(gate506inter6));
  inv1  gate2472(.a(G1274), .O(gate506inter7));
  inv1  gate2473(.a(G1275), .O(gate506inter8));
  nand2 gate2474(.a(gate506inter8), .b(gate506inter7), .O(gate506inter9));
  nand2 gate2475(.a(s_275), .b(gate506inter3), .O(gate506inter10));
  nor2  gate2476(.a(gate506inter10), .b(gate506inter9), .O(gate506inter11));
  nor2  gate2477(.a(gate506inter11), .b(gate506inter6), .O(gate506inter12));
  nand2 gate2478(.a(gate506inter12), .b(gate506inter1), .O(G1315));

  xor2  gate715(.a(G1277), .b(G1276), .O(gate507inter0));
  nand2 gate716(.a(gate507inter0), .b(s_24), .O(gate507inter1));
  and2  gate717(.a(G1277), .b(G1276), .O(gate507inter2));
  inv1  gate718(.a(s_24), .O(gate507inter3));
  inv1  gate719(.a(s_25), .O(gate507inter4));
  nand2 gate720(.a(gate507inter4), .b(gate507inter3), .O(gate507inter5));
  nor2  gate721(.a(gate507inter5), .b(gate507inter2), .O(gate507inter6));
  inv1  gate722(.a(G1276), .O(gate507inter7));
  inv1  gate723(.a(G1277), .O(gate507inter8));
  nand2 gate724(.a(gate507inter8), .b(gate507inter7), .O(gate507inter9));
  nand2 gate725(.a(s_25), .b(gate507inter3), .O(gate507inter10));
  nor2  gate726(.a(gate507inter10), .b(gate507inter9), .O(gate507inter11));
  nor2  gate727(.a(gate507inter11), .b(gate507inter6), .O(gate507inter12));
  nand2 gate728(.a(gate507inter12), .b(gate507inter1), .O(G1316));
nand2 gate508( .a(G1278), .b(G1279), .O(G1317) );
nand2 gate509( .a(G1280), .b(G1281), .O(G1318) );
nand2 gate510( .a(G1282), .b(G1283), .O(G1319) );

  xor2  gate1597(.a(G1285), .b(G1284), .O(gate511inter0));
  nand2 gate1598(.a(gate511inter0), .b(s_150), .O(gate511inter1));
  and2  gate1599(.a(G1285), .b(G1284), .O(gate511inter2));
  inv1  gate1600(.a(s_150), .O(gate511inter3));
  inv1  gate1601(.a(s_151), .O(gate511inter4));
  nand2 gate1602(.a(gate511inter4), .b(gate511inter3), .O(gate511inter5));
  nor2  gate1603(.a(gate511inter5), .b(gate511inter2), .O(gate511inter6));
  inv1  gate1604(.a(G1284), .O(gate511inter7));
  inv1  gate1605(.a(G1285), .O(gate511inter8));
  nand2 gate1606(.a(gate511inter8), .b(gate511inter7), .O(gate511inter9));
  nand2 gate1607(.a(s_151), .b(gate511inter3), .O(gate511inter10));
  nor2  gate1608(.a(gate511inter10), .b(gate511inter9), .O(gate511inter11));
  nor2  gate1609(.a(gate511inter11), .b(gate511inter6), .O(gate511inter12));
  nand2 gate1610(.a(gate511inter12), .b(gate511inter1), .O(G1320));
nand2 gate512( .a(G1286), .b(G1287), .O(G1321) );
nand2 gate513( .a(G1288), .b(G1289), .O(G1322) );
nand2 gate514( .a(G1290), .b(G1291), .O(G1323) );
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule