module c1908 (N1,N4,N7,N10,N13,N16,N19,N22,N25,N28,
              N31,N34,N37,N40,N43,N46,N49,N53,N56,N60,
              N63,N66,N69,N72,N76,N79,N82,N85,N88,N91,
              N94,N99,N104,N2753,N2754,N2755,N2756,N2762,N2767,N2768,
              N2779,N2780,N2781,N2782,N2783,N2784,N2785,N2786,N2787,N2811,
              N2886,N2887,N2888,N2889,N2890,N2891,N2892,N2899);
input N1,N4,N7,N10,N13,N16,N19,N22,N25,N28,
      N31,N34,N37,N40,N43,N46,N49,N53,N56,N60,
      N63,N66,N69,N72,N76,N79,N82,N85,N88,N91,
      N94,N99,N104;
  input s_0, s_1, s_2, s_3, s_4, s_5, s_6, s_7, s_8, s_9, s_10, s_11, s_12, s_13, s_14, s_15, s_16, s_17, s_18, s_19, s_20, s_21, s_22, s_23, s_24, s_25, s_26, s_27, s_28, s_29, s_30, s_31, s_32, s_33, s_34, s_35, s_36, s_37, s_38, s_39, s_40, s_41, s_42, s_43, s_44, s_45, s_46, s_47, s_48, s_49, s_50, s_51, s_52, s_53, s_54, s_55, s_56, s_57, s_58, s_59, s_60, s_61, s_62, s_63, s_64, s_65, s_66, s_67, s_68, s_69, s_70, s_71;
output N2753,N2754,N2755,N2756,N2762,N2767,N2768,N2779,N2780,N2781,
       N2782,N2783,N2784,N2785,N2786,N2787,N2811,N2886,N2887,N2888,
       N2889,N2890,N2891,N2892,N2899;
wire N190,N194,N197,N201,N206,N209,N212,N216,N220,N225,
     N229,N232,N235,N239,N243,N247,N251,N252,N253,N256,
     N257,N260,N263,N266,N269,N272,N275,N276,N277,N280,
     N283,N290,N297,N300,N303,N306,N313,N316,N319,N326,
     N331,N338,N343,N346,N349,N352,N355,N358,N361,N364,
     N367,N370,N373,N376,N379,N382,N385,N388,N534,N535,
     N536,N537,N538,N539,N540,N541,N542,N543,N544,N545,
     N546,N547,N548,N549,N550,N551,N552,N553,N554,N555,
     N556,N559,N562,N565,N568,N571,N574,N577,N580,N583,
     N586,N589,N592,N595,N598,N601,N602,N603,N608,N612,
     N616,N619,N622,N625,N628,N631,N634,N637,N640,N643,
     N646,N649,N652,N655,N658,N661,N664,N667,N670,N673,
     N676,N679,N682,N685,N688,N691,N694,N697,N700,N703,
     N706,N709,N712,N715,N718,N721,N724,N727,N730,N733,
     N736,N739,N742,N745,N748,N751,N886,N887,N888,N889,
     N890,N891,N892,N893,N894,N895,N896,N897,N898,N899,
     N903,N907,N910,N913,N914,N915,N916,N917,N918,N919,
     N920,N921,N922,N923,N926,N935,N938,N939,N942,N943,
     N946,N947,N950,N951,N954,N955,N958,N959,N962,N965,
     N968,N969,N972,N973,N976,N977,N980,N981,N984,N985,
     N988,N989,N990,N991,N992,N993,N994,N997,N998,N1001,
     N1002,N1003,N1004,N1005,N1006,N1007,N1008,N1009,N1010,N1013,
     N1016,N1019,N1022,N1025,N1028,N1031,N1034,N1037,N1040,N1043,
     N1046,N1049,N1054,N1055,N1063,N1064,N1067,N1068,N1119,N1120,
     N1121,N1122,N1128,N1129,N1130,N1131,N1132,N1133,N1148,N1149,
     N1150,N1151,N1152,N1153,N1154,N1155,N1156,N1157,N1158,N1159,
     N1160,N1161,N1162,N1163,N1164,N1167,N1168,N1171,N1188,N1205,
     N1206,N1207,N1208,N1209,N1210,N1211,N1212,N1213,N1214,N1215,
     N1216,N1217,N1218,N1219,N1220,N1221,N1222,N1223,N1224,N1225,
     N1226,N1227,N1228,N1229,N1230,N1231,N1232,N1235,N1238,N1239,
     N1240,N1241,N1242,N1243,N1246,N1249,N1252,N1255,N1258,N1261,
     N1264,N1267,N1309,N1310,N1311,N1312,N1313,N1314,N1315,N1316,
     N1317,N1318,N1319,N1322,N1327,N1328,N1334,N1344,N1345,N1346,
     N1348,N1349,N1350,N1351,N1352,N1355,N1358,N1361,N1364,N1367,
     N1370,N1373,N1376,N1379,N1383,N1386,N1387,N1388,N1389,N1390,
     N1393,N1396,N1397,N1398,N1399,N1409,N1412,N1413,N1416,N1419,
     N1433,N1434,N1438,N1439,N1440,N1443,N1444,N1445,N1446,N1447,
     N1448,N1451,N1452,N1453,N1454,N1455,N1456,N1457,N1458,N1459,
     N1460,N1461,N1462,N1463,N1464,N1468,N1469,N1470,N1471,N1472,
     N1475,N1476,N1478,N1481,N1484,N1487,N1488,N1489,N1490,N1491,
     N1492,N1493,N1494,N1495,N1496,N1498,N1499,N1500,N1501,N1504,
     N1510,N1513,N1514,N1517,N1520,N1521,N1522,N1526,N1527,N1528,
     N1529,N1530,N1531,N1532,N1534,N1537,N1540,N1546,N1554,N1557,
     N1561,N1567,N1568,N1569,N1571,N1576,N1588,N1591,N1593,N1594,
     N1595,N1596,N1600,N1603,N1606,N1609,N1612,N1615,N1620,N1623,
     N1635,N1636,N1638,N1639,N1640,N1643,N1647,N1651,N1658,N1661,
     N1664,N1671,N1672,N1675,N1677,N1678,N1679,N1680,N1681,N1682,
     N1683,N1685,N1688,N1697,N1701,N1706,N1707,N1708,N1709,N1710,
     N1711,N1712,N1713,N1714,N1717,N1720,N1721,N1723,N1727,N1728,
     N1730,N1731,N1734,N1740,N1741,N1742,N1746,N1747,N1748,N1751,
     N1759,N1761,N1762,N1763,N1764,N1768,N1769,N1772,N1773,N1774,
     N1777,N1783,N1784,N1785,N1786,N1787,N1788,N1791,N1792,N1795,
     N1796,N1798,N1801,N1802,N1807,N1808,N1809,N1810,N1812,N1815,
     N1818,N1821,N1822,N1823,N1824,N1825,N1826,N1827,N1830,N1837,
     N1838,N1841,N1848,N1849,N1850,N1852,N1855,N1856,N1857,N1858,
     N1864,N1865,N1866,N1869,N1872,N1875,N1878,N1879,N1882,N1883,
     N1884,N1885,N1889,N1895,N1896,N1897,N1898,N1902,N1910,N1911,
     N1912,N1913,N1915,N1919,N1920,N1921,N1922,N1923,N1924,N1927,
     N1930,N1933,N1936,N1937,N1938,N1941,N1942,N1944,N1947,N1950,
     N1953,N1958,N1961,N1965,N1968,N1975,N1976,N1977,N1978,N1979,
     N1980,N1985,N1987,N1999,N2000,N2002,N2003,N2004,N2005,N2006,
     N2007,N2008,N2009,N2012,N2013,N2014,N2015,N2016,N2018,N2019,
     N2020,N2021,N2022,N2023,N2024,N2025,N2026,N2027,N2030,N2033,
     N2036,N2037,N2038,N2039,N2040,N2041,N2042,N2047,N2052,N2055,
     N2060,N2061,N2062,N2067,N2068,N2071,N2076,N2077,N2078,N2081,
     N2086,N2089,N2104,N2119,N2129,N2143,N2148,N2151,N2196,N2199,
     N2202,N2205,N2214,N2215,N2216,N2217,N2222,N2223,N2224,N2225,
     N2226,N2227,N2228,N2229,N2230,N2231,N2232,N2233,N2234,N2235,
     N2236,N2237,N2240,N2241,N2244,N2245,N2250,N2253,N2256,N2257,
     N2260,N2263,N2266,N2269,N2272,N2279,N2286,N2297,N2315,N2326,
     N2340,N2353,N2361,N2375,N2384,N2385,N2386,N2426,N2427,N2537,
     N2540,N2543,N2546,N2549,N2552,N2555,N2558,N2561,N2564,N2567,
     N2570,N2573,N2576,N2594,N2597,N2600,N2603,N2606,N2611,N2614,
     N2617,N2620,N2627,N2628,N2629,N2630,N2631,N2632,N2633,N2634,
     N2639,N2642,N2645,N2648,N2651,N2655,N2658,N2661,N2664,N2669,
     N2670,N2671,N2672,N2673,N2674,N2675,N2676,N2682,N2683,N2688,
     N2689,N2690,N2691,N2710,N2720,N2721,N2722,N2723,N2724,N2725,
     N2726,N2727,N2728,N2729,N2730,N2731,N2732,N2733,N2734,N2735,
     N2736,N2737,N2738,N2739,N2740,N2741,N2742,N2743,N2744,N2745,
     N2746,N2747,N2750,N2757,N2758,N2759,N2760,N2761,N2763,N2764,
     N2765,N2766,N2773,N2776,N2788,N2789,N2800,N2807,N2808,N2809,
     N2810,N2812,N2815,N2818,N2821,N2824,N2827,N2828,N2829,N2843,
     N2846,N2850,N2851,N2852,N2853,N2854,N2857,N2858,N2859,N2860,
     N2861,N2862,N2863,N2866,N2867,N2868,N2869,N2870,N2871,N2872,
     N2873,N2874,N2875,N2876,N2877,N2878,N2879,N2880,N2881,N2882,
     N2883,N2895,N2896,N2897,N2898, gate532inter0, gate532inter1, gate532inter2, gate532inter3, gate532inter4, gate532inter5, gate532inter6, gate532inter7, gate532inter8, gate532inter9, gate532inter10, gate532inter11, gate532inter12, gate336inter0, gate336inter1, gate336inter2, gate336inter3, gate336inter4, gate336inter5, gate336inter6, gate336inter7, gate336inter8, gate336inter9, gate336inter10, gate336inter11, gate336inter12, gate866inter0, gate866inter1, gate866inter2, gate866inter3, gate866inter4, gate866inter5, gate866inter6, gate866inter7, gate866inter8, gate866inter9, gate866inter10, gate866inter11, gate866inter12, gate503inter0, gate503inter1, gate503inter2, gate503inter3, gate503inter4, gate503inter5, gate503inter6, gate503inter7, gate503inter8, gate503inter9, gate503inter10, gate503inter11, gate503inter12, gate784inter0, gate784inter1, gate784inter2, gate784inter3, gate784inter4, gate784inter5, gate784inter6, gate784inter7, gate784inter8, gate784inter9, gate784inter10, gate784inter11, gate784inter12, gate817inter0, gate817inter1, gate817inter2, gate817inter3, gate817inter4, gate817inter5, gate817inter6, gate817inter7, gate817inter8, gate817inter9, gate817inter10, gate817inter11, gate817inter12, gate633inter0, gate633inter1, gate633inter2, gate633inter3, gate633inter4, gate633inter5, gate633inter6, gate633inter7, gate633inter8, gate633inter9, gate633inter10, gate633inter11, gate633inter12, gate762inter0, gate762inter1, gate762inter2, gate762inter3, gate762inter4, gate762inter5, gate762inter6, gate762inter7, gate762inter8, gate762inter9, gate762inter10, gate762inter11, gate762inter12, gate482inter0, gate482inter1, gate482inter2, gate482inter3, gate482inter4, gate482inter5, gate482inter6, gate482inter7, gate482inter8, gate482inter9, gate482inter10, gate482inter11, gate482inter12, gate574inter0, gate574inter1, gate574inter2, gate574inter3, gate574inter4, gate574inter5, gate574inter6, gate574inter7, gate574inter8, gate574inter9, gate574inter10, gate574inter11, gate574inter12, gate304inter0, gate304inter1, gate304inter2, gate304inter3, gate304inter4, gate304inter5, gate304inter6, gate304inter7, gate304inter8, gate304inter9, gate304inter10, gate304inter11, gate304inter12, gate97inter0, gate97inter1, gate97inter2, gate97inter3, gate97inter4, gate97inter5, gate97inter6, gate97inter7, gate97inter8, gate97inter9, gate97inter10, gate97inter11, gate97inter12, gate563inter0, gate563inter1, gate563inter2, gate563inter3, gate563inter4, gate563inter5, gate563inter6, gate563inter7, gate563inter8, gate563inter9, gate563inter10, gate563inter11, gate563inter12, gate843inter0, gate843inter1, gate843inter2, gate843inter3, gate843inter4, gate843inter5, gate843inter6, gate843inter7, gate843inter8, gate843inter9, gate843inter10, gate843inter11, gate843inter12, gate752inter0, gate752inter1, gate752inter2, gate752inter3, gate752inter4, gate752inter5, gate752inter6, gate752inter7, gate752inter8, gate752inter9, gate752inter10, gate752inter11, gate752inter12, gate756inter0, gate756inter1, gate756inter2, gate756inter3, gate756inter4, gate756inter5, gate756inter6, gate756inter7, gate756inter8, gate756inter9, gate756inter10, gate756inter11, gate756inter12, gate351inter0, gate351inter1, gate351inter2, gate351inter3, gate351inter4, gate351inter5, gate351inter6, gate351inter7, gate351inter8, gate351inter9, gate351inter10, gate351inter11, gate351inter12, gate289inter0, gate289inter1, gate289inter2, gate289inter3, gate289inter4, gate289inter5, gate289inter6, gate289inter7, gate289inter8, gate289inter9, gate289inter10, gate289inter11, gate289inter12, gate858inter0, gate858inter1, gate858inter2, gate858inter3, gate858inter4, gate858inter5, gate858inter6, gate858inter7, gate858inter8, gate858inter9, gate858inter10, gate858inter11, gate858inter12, gate559inter0, gate559inter1, gate559inter2, gate559inter3, gate559inter4, gate559inter5, gate559inter6, gate559inter7, gate559inter8, gate559inter9, gate559inter10, gate559inter11, gate559inter12, gate163inter0, gate163inter1, gate163inter2, gate163inter3, gate163inter4, gate163inter5, gate163inter6, gate163inter7, gate163inter8, gate163inter9, gate163inter10, gate163inter11, gate163inter12, gate279inter0, gate279inter1, gate279inter2, gate279inter3, gate279inter4, gate279inter5, gate279inter6, gate279inter7, gate279inter8, gate279inter9, gate279inter10, gate279inter11, gate279inter12, gate676inter0, gate676inter1, gate676inter2, gate676inter3, gate676inter4, gate676inter5, gate676inter6, gate676inter7, gate676inter8, gate676inter9, gate676inter10, gate676inter11, gate676inter12, gate393inter0, gate393inter1, gate393inter2, gate393inter3, gate393inter4, gate393inter5, gate393inter6, gate393inter7, gate393inter8, gate393inter9, gate393inter10, gate393inter11, gate393inter12, gate513inter0, gate513inter1, gate513inter2, gate513inter3, gate513inter4, gate513inter5, gate513inter6, gate513inter7, gate513inter8, gate513inter9, gate513inter10, gate513inter11, gate513inter12, gate497inter0, gate497inter1, gate497inter2, gate497inter3, gate497inter4, gate497inter5, gate497inter6, gate497inter7, gate497inter8, gate497inter9, gate497inter10, gate497inter11, gate497inter12, gate499inter0, gate499inter1, gate499inter2, gate499inter3, gate499inter4, gate499inter5, gate499inter6, gate499inter7, gate499inter8, gate499inter9, gate499inter10, gate499inter11, gate499inter12, gate683inter0, gate683inter1, gate683inter2, gate683inter3, gate683inter4, gate683inter5, gate683inter6, gate683inter7, gate683inter8, gate683inter9, gate683inter10, gate683inter11, gate683inter12, gate416inter0, gate416inter1, gate416inter2, gate416inter3, gate416inter4, gate416inter5, gate416inter6, gate416inter7, gate416inter8, gate416inter9, gate416inter10, gate416inter11, gate416inter12, gate596inter0, gate596inter1, gate596inter2, gate596inter3, gate596inter4, gate596inter5, gate596inter6, gate596inter7, gate596inter8, gate596inter9, gate596inter10, gate596inter11, gate596inter12, gate839inter0, gate839inter1, gate839inter2, gate839inter3, gate839inter4, gate839inter5, gate839inter6, gate839inter7, gate839inter8, gate839inter9, gate839inter10, gate839inter11, gate839inter12, gate627inter0, gate627inter1, gate627inter2, gate627inter3, gate627inter4, gate627inter5, gate627inter6, gate627inter7, gate627inter8, gate627inter9, gate627inter10, gate627inter11, gate627inter12, gate418inter0, gate418inter1, gate418inter2, gate418inter3, gate418inter4, gate418inter5, gate418inter6, gate418inter7, gate418inter8, gate418inter9, gate418inter10, gate418inter11, gate418inter12, gate806inter0, gate806inter1, gate806inter2, gate806inter3, gate806inter4, gate806inter5, gate806inter6, gate806inter7, gate806inter8, gate806inter9, gate806inter10, gate806inter11, gate806inter12, gate389inter0, gate389inter1, gate389inter2, gate389inter3, gate389inter4, gate389inter5, gate389inter6, gate389inter7, gate389inter8, gate389inter9, gate389inter10, gate389inter11, gate389inter12, gate760inter0, gate760inter1, gate760inter2, gate760inter3, gate760inter4, gate760inter5, gate760inter6, gate760inter7, gate760inter8, gate760inter9, gate760inter10, gate760inter11, gate760inter12;


inv1 gate1( .a(N1), .O(N190) );
inv1 gate2( .a(N4), .O(N194) );
inv1 gate3( .a(N7), .O(N197) );
inv1 gate4( .a(N10), .O(N201) );
inv1 gate5( .a(N13), .O(N206) );
inv1 gate6( .a(N16), .O(N209) );
inv1 gate7( .a(N19), .O(N212) );
inv1 gate8( .a(N22), .O(N216) );
inv1 gate9( .a(N25), .O(N220) );
inv1 gate10( .a(N28), .O(N225) );
inv1 gate11( .a(N31), .O(N229) );
inv1 gate12( .a(N34), .O(N232) );
inv1 gate13( .a(N37), .O(N235) );
inv1 gate14( .a(N40), .O(N239) );
inv1 gate15( .a(N43), .O(N243) );
inv1 gate16( .a(N46), .O(N247) );
nand2 gate17( .a(N63), .b(N88), .O(N251) );
nand2 gate18( .a(N66), .b(N91), .O(N252) );
inv1 gate19( .a(N72), .O(N253) );
inv1 gate20( .a(N72), .O(N256) );
buf1 gate21( .a(N69), .O(N257) );
buf1 gate22( .a(N69), .O(N260) );
inv1 gate23( .a(N76), .O(N263) );
inv1 gate24( .a(N79), .O(N266) );
inv1 gate25( .a(N82), .O(N269) );
inv1 gate26( .a(N85), .O(N272) );
inv1 gate27( .a(N104), .O(N275) );
inv1 gate28( .a(N104), .O(N276) );
inv1 gate29( .a(N88), .O(N277) );
inv1 gate30( .a(N91), .O(N280) );
buf1 gate31( .a(N94), .O(N283) );
inv1 gate32( .a(N94), .O(N290) );
buf1 gate33( .a(N94), .O(N297) );
inv1 gate34( .a(N94), .O(N300) );
buf1 gate35( .a(N99), .O(N303) );
inv1 gate36( .a(N99), .O(N306) );
inv1 gate37( .a(N99), .O(N313) );
buf1 gate38( .a(N104), .O(N316) );
inv1 gate39( .a(N104), .O(N319) );
buf1 gate40( .a(N104), .O(N326) );
buf1 gate41( .a(N104), .O(N331) );
inv1 gate42( .a(N104), .O(N338) );
buf1 gate43( .a(N1), .O(N343) );
buf1 gate44( .a(N4), .O(N346) );
buf1 gate45( .a(N7), .O(N349) );
buf1 gate46( .a(N10), .O(N352) );
buf1 gate47( .a(N13), .O(N355) );
buf1 gate48( .a(N16), .O(N358) );
buf1 gate49( .a(N19), .O(N361) );
buf1 gate50( .a(N22), .O(N364) );
buf1 gate51( .a(N25), .O(N367) );
buf1 gate52( .a(N28), .O(N370) );
buf1 gate53( .a(N31), .O(N373) );
buf1 gate54( .a(N34), .O(N376) );
buf1 gate55( .a(N37), .O(N379) );
buf1 gate56( .a(N40), .O(N382) );
buf1 gate57( .a(N43), .O(N385) );
buf1 gate58( .a(N46), .O(N388) );
inv1 gate59( .a(N343), .O(N534) );
inv1 gate60( .a(N346), .O(N535) );
inv1 gate61( .a(N349), .O(N536) );
inv1 gate62( .a(N352), .O(N537) );
inv1 gate63( .a(N355), .O(N538) );
inv1 gate64( .a(N358), .O(N539) );
inv1 gate65( .a(N361), .O(N540) );
inv1 gate66( .a(N364), .O(N541) );
inv1 gate67( .a(N367), .O(N542) );
inv1 gate68( .a(N370), .O(N543) );
inv1 gate69( .a(N373), .O(N544) );
inv1 gate70( .a(N376), .O(N545) );
inv1 gate71( .a(N379), .O(N546) );
inv1 gate72( .a(N382), .O(N547) );
inv1 gate73( .a(N385), .O(N548) );
inv1 gate74( .a(N388), .O(N549) );
nand2 gate75( .a(N306), .b(N331), .O(N550) );
nand2 gate76( .a(N306), .b(N331), .O(N551) );
nand2 gate77( .a(N306), .b(N331), .O(N552) );
nand2 gate78( .a(N306), .b(N331), .O(N553) );
nand2 gate79( .a(N306), .b(N331), .O(N554) );
nand2 gate80( .a(N306), .b(N331), .O(N555) );
buf1 gate81( .a(N190), .O(N556) );
buf1 gate82( .a(N194), .O(N559) );
buf1 gate83( .a(N206), .O(N562) );
buf1 gate84( .a(N209), .O(N565) );
buf1 gate85( .a(N225), .O(N568) );
buf1 gate86( .a(N243), .O(N571) );
and2 gate87( .a(N63), .b(N319), .O(N574) );
buf1 gate88( .a(N220), .O(N577) );
buf1 gate89( .a(N229), .O(N580) );
buf1 gate90( .a(N232), .O(N583) );
and2 gate91( .a(N66), .b(N319), .O(N586) );
buf1 gate92( .a(N239), .O(N589) );
and3 gate93( .a(N49), .b(N253), .c(N319), .O(N592) );
buf1 gate94( .a(N247), .O(N595) );
buf1 gate95( .a(N239), .O(N598) );
nand2 gate96( .a(N326), .b(N277), .O(N601) );

  xor2  gate1035(.a(N280), .b(N326), .O(gate97inter0));
  nand2 gate1036(.a(gate97inter0), .b(s_22), .O(gate97inter1));
  and2  gate1037(.a(N280), .b(N326), .O(gate97inter2));
  inv1  gate1038(.a(s_22), .O(gate97inter3));
  inv1  gate1039(.a(s_23), .O(gate97inter4));
  nand2 gate1040(.a(gate97inter4), .b(gate97inter3), .O(gate97inter5));
  nor2  gate1041(.a(gate97inter5), .b(gate97inter2), .O(gate97inter6));
  inv1  gate1042(.a(N326), .O(gate97inter7));
  inv1  gate1043(.a(N280), .O(gate97inter8));
  nand2 gate1044(.a(gate97inter8), .b(gate97inter7), .O(gate97inter9));
  nand2 gate1045(.a(s_23), .b(gate97inter3), .O(gate97inter10));
  nor2  gate1046(.a(gate97inter10), .b(gate97inter9), .O(gate97inter11));
  nor2  gate1047(.a(gate97inter11), .b(gate97inter6), .O(gate97inter12));
  nand2 gate1048(.a(gate97inter12), .b(gate97inter1), .O(N602));
nand2 gate98( .a(N260), .b(N72), .O(N603) );
nand2 gate99( .a(N260), .b(N300), .O(N608) );
nand2 gate100( .a(N256), .b(N300), .O(N612) );
buf1 gate101( .a(N201), .O(N616) );
buf1 gate102( .a(N216), .O(N619) );
buf1 gate103( .a(N220), .O(N622) );
buf1 gate104( .a(N239), .O(N625) );
buf1 gate105( .a(N190), .O(N628) );
buf1 gate106( .a(N190), .O(N631) );
buf1 gate107( .a(N194), .O(N634) );
buf1 gate108( .a(N229), .O(N637) );
buf1 gate109( .a(N197), .O(N640) );
and3 gate110( .a(N56), .b(N257), .c(N319), .O(N643) );
buf1 gate111( .a(N232), .O(N646) );
buf1 gate112( .a(N201), .O(N649) );
buf1 gate113( .a(N235), .O(N652) );
and3 gate114( .a(N60), .b(N257), .c(N319), .O(N655) );
buf1 gate115( .a(N263), .O(N658) );
buf1 gate116( .a(N263), .O(N661) );
buf1 gate117( .a(N266), .O(N664) );
buf1 gate118( .a(N266), .O(N667) );
buf1 gate119( .a(N269), .O(N670) );
buf1 gate120( .a(N269), .O(N673) );
buf1 gate121( .a(N272), .O(N676) );
buf1 gate122( .a(N272), .O(N679) );
and2 gate123( .a(N251), .b(N316), .O(N682) );
and2 gate124( .a(N252), .b(N316), .O(N685) );
buf1 gate125( .a(N197), .O(N688) );
buf1 gate126( .a(N197), .O(N691) );
buf1 gate127( .a(N212), .O(N694) );
buf1 gate128( .a(N212), .O(N697) );
buf1 gate129( .a(N247), .O(N700) );
buf1 gate130( .a(N247), .O(N703) );
buf1 gate131( .a(N235), .O(N706) );
buf1 gate132( .a(N235), .O(N709) );
buf1 gate133( .a(N201), .O(N712) );
buf1 gate134( .a(N201), .O(N715) );
buf1 gate135( .a(N206), .O(N718) );
buf1 gate136( .a(N216), .O(N721) );
and3 gate137( .a(N53), .b(N253), .c(N319), .O(N724) );
buf1 gate138( .a(N243), .O(N727) );
buf1 gate139( .a(N220), .O(N730) );
buf1 gate140( .a(N220), .O(N733) );
buf1 gate141( .a(N209), .O(N736) );
buf1 gate142( .a(N216), .O(N739) );
buf1 gate143( .a(N225), .O(N742) );
buf1 gate144( .a(N243), .O(N745) );
buf1 gate145( .a(N212), .O(N748) );
buf1 gate146( .a(N225), .O(N751) );
inv1 gate147( .a(N682), .O(N886) );
inv1 gate148( .a(N685), .O(N887) );
inv1 gate149( .a(N616), .O(N888) );
inv1 gate150( .a(N619), .O(N889) );
inv1 gate151( .a(N622), .O(N890) );
inv1 gate152( .a(N625), .O(N891) );
inv1 gate153( .a(N631), .O(N892) );
inv1 gate154( .a(N643), .O(N893) );
inv1 gate155( .a(N649), .O(N894) );
inv1 gate156( .a(N652), .O(N895) );
inv1 gate157( .a(N655), .O(N896) );
and2 gate158( .a(N49), .b(N612), .O(N897) );
and2 gate159( .a(N56), .b(N608), .O(N898) );
nand2 gate160( .a(N53), .b(N612), .O(N899) );
nand2 gate161( .a(N60), .b(N608), .O(N903) );
nand2 gate162( .a(N49), .b(N612), .O(N907) );

  xor2  gate1161(.a(N608), .b(N56), .O(gate163inter0));
  nand2 gate1162(.a(gate163inter0), .b(s_40), .O(gate163inter1));
  and2  gate1163(.a(N608), .b(N56), .O(gate163inter2));
  inv1  gate1164(.a(s_40), .O(gate163inter3));
  inv1  gate1165(.a(s_41), .O(gate163inter4));
  nand2 gate1166(.a(gate163inter4), .b(gate163inter3), .O(gate163inter5));
  nor2  gate1167(.a(gate163inter5), .b(gate163inter2), .O(gate163inter6));
  inv1  gate1168(.a(N56), .O(gate163inter7));
  inv1  gate1169(.a(N608), .O(gate163inter8));
  nand2 gate1170(.a(gate163inter8), .b(gate163inter7), .O(gate163inter9));
  nand2 gate1171(.a(s_41), .b(gate163inter3), .O(gate163inter10));
  nor2  gate1172(.a(gate163inter10), .b(gate163inter9), .O(gate163inter11));
  nor2  gate1173(.a(gate163inter11), .b(gate163inter6), .O(gate163inter12));
  nand2 gate1174(.a(gate163inter12), .b(gate163inter1), .O(N910));
inv1 gate164( .a(N661), .O(N913) );
inv1 gate165( .a(N658), .O(N914) );
inv1 gate166( .a(N667), .O(N915) );
inv1 gate167( .a(N664), .O(N916) );
inv1 gate168( .a(N673), .O(N917) );
inv1 gate169( .a(N670), .O(N918) );
inv1 gate170( .a(N679), .O(N919) );
inv1 gate171( .a(N676), .O(N920) );
nand4 gate172( .a(N277), .b(N297), .c(N326), .d(N603), .O(N921) );
nand4 gate173( .a(N280), .b(N297), .c(N326), .d(N603), .O(N922) );
nand3 gate174( .a(N303), .b(N338), .c(N603), .O(N923) );
and3 gate175( .a(N303), .b(N338), .c(N603), .O(N926) );
buf1 gate176( .a(N556), .O(N935) );
inv1 gate177( .a(N688), .O(N938) );
buf1 gate178( .a(N556), .O(N939) );
inv1 gate179( .a(N691), .O(N942) );
buf1 gate180( .a(N562), .O(N943) );
inv1 gate181( .a(N694), .O(N946) );
buf1 gate182( .a(N562), .O(N947) );
inv1 gate183( .a(N697), .O(N950) );
buf1 gate184( .a(N568), .O(N951) );
inv1 gate185( .a(N700), .O(N954) );
buf1 gate186( .a(N568), .O(N955) );
inv1 gate187( .a(N703), .O(N958) );
buf1 gate188( .a(N574), .O(N959) );
buf1 gate189( .a(N574), .O(N962) );
buf1 gate190( .a(N580), .O(N965) );
inv1 gate191( .a(N706), .O(N968) );
buf1 gate192( .a(N580), .O(N969) );
inv1 gate193( .a(N709), .O(N972) );
buf1 gate194( .a(N586), .O(N973) );
inv1 gate195( .a(N712), .O(N976) );
buf1 gate196( .a(N586), .O(N977) );
inv1 gate197( .a(N715), .O(N980) );
buf1 gate198( .a(N592), .O(N981) );
inv1 gate199( .a(N628), .O(N984) );
buf1 gate200( .a(N592), .O(N985) );
inv1 gate201( .a(N718), .O(N988) );
inv1 gate202( .a(N721), .O(N989) );
inv1 gate203( .a(N634), .O(N990) );
inv1 gate204( .a(N724), .O(N991) );
inv1 gate205( .a(N727), .O(N992) );
inv1 gate206( .a(N637), .O(N993) );
buf1 gate207( .a(N595), .O(N994) );
inv1 gate208( .a(N730), .O(N997) );
buf1 gate209( .a(N595), .O(N998) );
inv1 gate210( .a(N733), .O(N1001) );
inv1 gate211( .a(N736), .O(N1002) );
inv1 gate212( .a(N739), .O(N1003) );
inv1 gate213( .a(N640), .O(N1004) );
inv1 gate214( .a(N742), .O(N1005) );
inv1 gate215( .a(N745), .O(N1006) );
inv1 gate216( .a(N646), .O(N1007) );
inv1 gate217( .a(N748), .O(N1008) );
inv1 gate218( .a(N751), .O(N1009) );
buf1 gate219( .a(N559), .O(N1010) );
buf1 gate220( .a(N559), .O(N1013) );
buf1 gate221( .a(N565), .O(N1016) );
buf1 gate222( .a(N565), .O(N1019) );
buf1 gate223( .a(N571), .O(N1022) );
buf1 gate224( .a(N571), .O(N1025) );
buf1 gate225( .a(N577), .O(N1028) );
buf1 gate226( .a(N577), .O(N1031) );
buf1 gate227( .a(N583), .O(N1034) );
buf1 gate228( .a(N583), .O(N1037) );
buf1 gate229( .a(N589), .O(N1040) );
buf1 gate230( .a(N589), .O(N1043) );
buf1 gate231( .a(N598), .O(N1046) );
buf1 gate232( .a(N598), .O(N1049) );
nand2 gate233( .a(N619), .b(N888), .O(N1054) );
nand2 gate234( .a(N616), .b(N889), .O(N1055) );
nand2 gate235( .a(N625), .b(N890), .O(N1063) );
nand2 gate236( .a(N622), .b(N891), .O(N1064) );
nand2 gate237( .a(N655), .b(N895), .O(N1067) );
nand2 gate238( .a(N652), .b(N896), .O(N1068) );
nand2 gate239( .a(N721), .b(N988), .O(N1119) );
nand2 gate240( .a(N718), .b(N989), .O(N1120) );
nand2 gate241( .a(N727), .b(N991), .O(N1121) );
nand2 gate242( .a(N724), .b(N992), .O(N1122) );
nand2 gate243( .a(N739), .b(N1002), .O(N1128) );
nand2 gate244( .a(N736), .b(N1003), .O(N1129) );
nand2 gate245( .a(N745), .b(N1005), .O(N1130) );
nand2 gate246( .a(N742), .b(N1006), .O(N1131) );
nand2 gate247( .a(N751), .b(N1008), .O(N1132) );
nand2 gate248( .a(N748), .b(N1009), .O(N1133) );
inv1 gate249( .a(N939), .O(N1148) );
inv1 gate250( .a(N935), .O(N1149) );
nand2 gate251( .a(N1054), .b(N1055), .O(N1150) );
inv1 gate252( .a(N943), .O(N1151) );
inv1 gate253( .a(N947), .O(N1152) );
inv1 gate254( .a(N955), .O(N1153) );
inv1 gate255( .a(N951), .O(N1154) );
inv1 gate256( .a(N962), .O(N1155) );
inv1 gate257( .a(N969), .O(N1156) );
inv1 gate258( .a(N977), .O(N1157) );
nand2 gate259( .a(N1063), .b(N1064), .O(N1158) );
inv1 gate260( .a(N985), .O(N1159) );
nand2 gate261( .a(N985), .b(N892), .O(N1160) );
inv1 gate262( .a(N998), .O(N1161) );
nand2 gate263( .a(N1067), .b(N1068), .O(N1162) );
inv1 gate264( .a(N899), .O(N1163) );
buf1 gate265( .a(N899), .O(N1164) );
inv1 gate266( .a(N903), .O(N1167) );
buf1 gate267( .a(N903), .O(N1168) );
nand2 gate268( .a(N921), .b(N923), .O(N1171) );
nand2 gate269( .a(N922), .b(N923), .O(N1188) );
inv1 gate270( .a(N1010), .O(N1205) );
nand2 gate271( .a(N1010), .b(N938), .O(N1206) );
inv1 gate272( .a(N1013), .O(N1207) );
nand2 gate273( .a(N1013), .b(N942), .O(N1208) );
inv1 gate274( .a(N1016), .O(N1209) );
nand2 gate275( .a(N1016), .b(N946), .O(N1210) );
inv1 gate276( .a(N1019), .O(N1211) );
nand2 gate277( .a(N1019), .b(N950), .O(N1212) );
inv1 gate278( .a(N1022), .O(N1213) );

  xor2  gate1175(.a(N954), .b(N1022), .O(gate279inter0));
  nand2 gate1176(.a(gate279inter0), .b(s_42), .O(gate279inter1));
  and2  gate1177(.a(N954), .b(N1022), .O(gate279inter2));
  inv1  gate1178(.a(s_42), .O(gate279inter3));
  inv1  gate1179(.a(s_43), .O(gate279inter4));
  nand2 gate1180(.a(gate279inter4), .b(gate279inter3), .O(gate279inter5));
  nor2  gate1181(.a(gate279inter5), .b(gate279inter2), .O(gate279inter6));
  inv1  gate1182(.a(N1022), .O(gate279inter7));
  inv1  gate1183(.a(N954), .O(gate279inter8));
  nand2 gate1184(.a(gate279inter8), .b(gate279inter7), .O(gate279inter9));
  nand2 gate1185(.a(s_43), .b(gate279inter3), .O(gate279inter10));
  nor2  gate1186(.a(gate279inter10), .b(gate279inter9), .O(gate279inter11));
  nor2  gate1187(.a(gate279inter11), .b(gate279inter6), .O(gate279inter12));
  nand2 gate1188(.a(gate279inter12), .b(gate279inter1), .O(N1214));
inv1 gate280( .a(N1025), .O(N1215) );
nand2 gate281( .a(N1025), .b(N958), .O(N1216) );
inv1 gate282( .a(N1028), .O(N1217) );
inv1 gate283( .a(N959), .O(N1218) );
inv1 gate284( .a(N1031), .O(N1219) );
inv1 gate285( .a(N1034), .O(N1220) );
nand2 gate286( .a(N1034), .b(N968), .O(N1221) );
inv1 gate287( .a(N965), .O(N1222) );
inv1 gate288( .a(N1037), .O(N1223) );

  xor2  gate1119(.a(N972), .b(N1037), .O(gate289inter0));
  nand2 gate1120(.a(gate289inter0), .b(s_34), .O(gate289inter1));
  and2  gate1121(.a(N972), .b(N1037), .O(gate289inter2));
  inv1  gate1122(.a(s_34), .O(gate289inter3));
  inv1  gate1123(.a(s_35), .O(gate289inter4));
  nand2 gate1124(.a(gate289inter4), .b(gate289inter3), .O(gate289inter5));
  nor2  gate1125(.a(gate289inter5), .b(gate289inter2), .O(gate289inter6));
  inv1  gate1126(.a(N1037), .O(gate289inter7));
  inv1  gate1127(.a(N972), .O(gate289inter8));
  nand2 gate1128(.a(gate289inter8), .b(gate289inter7), .O(gate289inter9));
  nand2 gate1129(.a(s_35), .b(gate289inter3), .O(gate289inter10));
  nor2  gate1130(.a(gate289inter10), .b(gate289inter9), .O(gate289inter11));
  nor2  gate1131(.a(gate289inter11), .b(gate289inter6), .O(gate289inter12));
  nand2 gate1132(.a(gate289inter12), .b(gate289inter1), .O(N1224));
inv1 gate290( .a(N1040), .O(N1225) );
nand2 gate291( .a(N1040), .b(N976), .O(N1226) );
inv1 gate292( .a(N973), .O(N1227) );
inv1 gate293( .a(N1043), .O(N1228) );
nand2 gate294( .a(N1043), .b(N980), .O(N1229) );
inv1 gate295( .a(N981), .O(N1230) );
nand2 gate296( .a(N981), .b(N984), .O(N1231) );
nand2 gate297( .a(N1119), .b(N1120), .O(N1232) );
nand2 gate298( .a(N1121), .b(N1122), .O(N1235) );
inv1 gate299( .a(N1046), .O(N1238) );
nand2 gate300( .a(N1046), .b(N997), .O(N1239) );
inv1 gate301( .a(N994), .O(N1240) );
inv1 gate302( .a(N1049), .O(N1241) );
nand2 gate303( .a(N1049), .b(N1001), .O(N1242) );

  xor2  gate1021(.a(N1129), .b(N1128), .O(gate304inter0));
  nand2 gate1022(.a(gate304inter0), .b(s_20), .O(gate304inter1));
  and2  gate1023(.a(N1129), .b(N1128), .O(gate304inter2));
  inv1  gate1024(.a(s_20), .O(gate304inter3));
  inv1  gate1025(.a(s_21), .O(gate304inter4));
  nand2 gate1026(.a(gate304inter4), .b(gate304inter3), .O(gate304inter5));
  nor2  gate1027(.a(gate304inter5), .b(gate304inter2), .O(gate304inter6));
  inv1  gate1028(.a(N1128), .O(gate304inter7));
  inv1  gate1029(.a(N1129), .O(gate304inter8));
  nand2 gate1030(.a(gate304inter8), .b(gate304inter7), .O(gate304inter9));
  nand2 gate1031(.a(s_21), .b(gate304inter3), .O(gate304inter10));
  nor2  gate1032(.a(gate304inter10), .b(gate304inter9), .O(gate304inter11));
  nor2  gate1033(.a(gate304inter11), .b(gate304inter6), .O(gate304inter12));
  nand2 gate1034(.a(gate304inter12), .b(gate304inter1), .O(N1243));
nand2 gate305( .a(N1130), .b(N1131), .O(N1246) );
nand2 gate306( .a(N1132), .b(N1133), .O(N1249) );
buf1 gate307( .a(N907), .O(N1252) );
buf1 gate308( .a(N907), .O(N1255) );
buf1 gate309( .a(N910), .O(N1258) );
buf1 gate310( .a(N910), .O(N1261) );
inv1 gate311( .a(N1150), .O(N1264) );
nand2 gate312( .a(N631), .b(N1159), .O(N1267) );
nand2 gate313( .a(N688), .b(N1205), .O(N1309) );
nand2 gate314( .a(N691), .b(N1207), .O(N1310) );
nand2 gate315( .a(N694), .b(N1209), .O(N1311) );
nand2 gate316( .a(N697), .b(N1211), .O(N1312) );
nand2 gate317( .a(N700), .b(N1213), .O(N1313) );
nand2 gate318( .a(N703), .b(N1215), .O(N1314) );
nand2 gate319( .a(N706), .b(N1220), .O(N1315) );
nand2 gate320( .a(N709), .b(N1223), .O(N1316) );
nand2 gate321( .a(N712), .b(N1225), .O(N1317) );
nand2 gate322( .a(N715), .b(N1228), .O(N1318) );
inv1 gate323( .a(N1158), .O(N1319) );
nand2 gate324( .a(N628), .b(N1230), .O(N1322) );
nand2 gate325( .a(N730), .b(N1238), .O(N1327) );
nand2 gate326( .a(N733), .b(N1241), .O(N1328) );
inv1 gate327( .a(N1162), .O(N1334) );
nand2 gate328( .a(N1267), .b(N1160), .O(N1344) );
nand2 gate329( .a(N1249), .b(N894), .O(N1345) );
inv1 gate330( .a(N1249), .O(N1346) );
inv1 gate331( .a(N1255), .O(N1348) );
inv1 gate332( .a(N1252), .O(N1349) );
inv1 gate333( .a(N1261), .O(N1350) );
inv1 gate334( .a(N1258), .O(N1351) );
nand2 gate335( .a(N1309), .b(N1206), .O(N1352) );

  xor2  gate895(.a(N1208), .b(N1310), .O(gate336inter0));
  nand2 gate896(.a(gate336inter0), .b(s_2), .O(gate336inter1));
  and2  gate897(.a(N1208), .b(N1310), .O(gate336inter2));
  inv1  gate898(.a(s_2), .O(gate336inter3));
  inv1  gate899(.a(s_3), .O(gate336inter4));
  nand2 gate900(.a(gate336inter4), .b(gate336inter3), .O(gate336inter5));
  nor2  gate901(.a(gate336inter5), .b(gate336inter2), .O(gate336inter6));
  inv1  gate902(.a(N1310), .O(gate336inter7));
  inv1  gate903(.a(N1208), .O(gate336inter8));
  nand2 gate904(.a(gate336inter8), .b(gate336inter7), .O(gate336inter9));
  nand2 gate905(.a(s_3), .b(gate336inter3), .O(gate336inter10));
  nor2  gate906(.a(gate336inter10), .b(gate336inter9), .O(gate336inter11));
  nor2  gate907(.a(gate336inter11), .b(gate336inter6), .O(gate336inter12));
  nand2 gate908(.a(gate336inter12), .b(gate336inter1), .O(N1355));
nand2 gate337( .a(N1311), .b(N1210), .O(N1358) );
nand2 gate338( .a(N1312), .b(N1212), .O(N1361) );
nand2 gate339( .a(N1313), .b(N1214), .O(N1364) );
nand2 gate340( .a(N1314), .b(N1216), .O(N1367) );
nand2 gate341( .a(N1315), .b(N1221), .O(N1370) );
nand2 gate342( .a(N1316), .b(N1224), .O(N1373) );
nand2 gate343( .a(N1317), .b(N1226), .O(N1376) );
nand2 gate344( .a(N1318), .b(N1229), .O(N1379) );
nand2 gate345( .a(N1322), .b(N1231), .O(N1383) );
inv1 gate346( .a(N1232), .O(N1386) );
nand2 gate347( .a(N1232), .b(N990), .O(N1387) );
inv1 gate348( .a(N1235), .O(N1388) );
nand2 gate349( .a(N1235), .b(N993), .O(N1389) );
nand2 gate350( .a(N1327), .b(N1239), .O(N1390) );

  xor2  gate1105(.a(N1242), .b(N1328), .O(gate351inter0));
  nand2 gate1106(.a(gate351inter0), .b(s_32), .O(gate351inter1));
  and2  gate1107(.a(N1242), .b(N1328), .O(gate351inter2));
  inv1  gate1108(.a(s_32), .O(gate351inter3));
  inv1  gate1109(.a(s_33), .O(gate351inter4));
  nand2 gate1110(.a(gate351inter4), .b(gate351inter3), .O(gate351inter5));
  nor2  gate1111(.a(gate351inter5), .b(gate351inter2), .O(gate351inter6));
  inv1  gate1112(.a(N1328), .O(gate351inter7));
  inv1  gate1113(.a(N1242), .O(gate351inter8));
  nand2 gate1114(.a(gate351inter8), .b(gate351inter7), .O(gate351inter9));
  nand2 gate1115(.a(s_33), .b(gate351inter3), .O(gate351inter10));
  nor2  gate1116(.a(gate351inter10), .b(gate351inter9), .O(gate351inter11));
  nor2  gate1117(.a(gate351inter11), .b(gate351inter6), .O(gate351inter12));
  nand2 gate1118(.a(gate351inter12), .b(gate351inter1), .O(N1393));
inv1 gate352( .a(N1243), .O(N1396) );
nand2 gate353( .a(N1243), .b(N1004), .O(N1397) );
inv1 gate354( .a(N1246), .O(N1398) );
nand2 gate355( .a(N1246), .b(N1007), .O(N1399) );
inv1 gate356( .a(N1319), .O(N1409) );
nand2 gate357( .a(N649), .b(N1346), .O(N1412) );
inv1 gate358( .a(N1334), .O(N1413) );
buf1 gate359( .a(N1264), .O(N1416) );
buf1 gate360( .a(N1264), .O(N1419) );
nand2 gate361( .a(N634), .b(N1386), .O(N1433) );
nand2 gate362( .a(N637), .b(N1388), .O(N1434) );
nand2 gate363( .a(N640), .b(N1396), .O(N1438) );
nand2 gate364( .a(N646), .b(N1398), .O(N1439) );
inv1 gate365( .a(N1344), .O(N1440) );
nand2 gate366( .a(N1355), .b(N1148), .O(N1443) );
inv1 gate367( .a(N1355), .O(N1444) );
nand2 gate368( .a(N1352), .b(N1149), .O(N1445) );
inv1 gate369( .a(N1352), .O(N1446) );
nand2 gate370( .a(N1358), .b(N1151), .O(N1447) );
inv1 gate371( .a(N1358), .O(N1448) );
nand2 gate372( .a(N1361), .b(N1152), .O(N1451) );
inv1 gate373( .a(N1361), .O(N1452) );
nand2 gate374( .a(N1367), .b(N1153), .O(N1453) );
inv1 gate375( .a(N1367), .O(N1454) );
nand2 gate376( .a(N1364), .b(N1154), .O(N1455) );
inv1 gate377( .a(N1364), .O(N1456) );
nand2 gate378( .a(N1373), .b(N1156), .O(N1457) );
inv1 gate379( .a(N1373), .O(N1458) );
nand2 gate380( .a(N1379), .b(N1157), .O(N1459) );
inv1 gate381( .a(N1379), .O(N1460) );
inv1 gate382( .a(N1383), .O(N1461) );
nand2 gate383( .a(N1393), .b(N1161), .O(N1462) );
inv1 gate384( .a(N1393), .O(N1463) );
nand2 gate385( .a(N1345), .b(N1412), .O(N1464) );
inv1 gate386( .a(N1370), .O(N1468) );
nand2 gate387( .a(N1370), .b(N1222), .O(N1469) );
inv1 gate388( .a(N1376), .O(N1470) );

  xor2  gate1357(.a(N1227), .b(N1376), .O(gate389inter0));
  nand2 gate1358(.a(gate389inter0), .b(s_68), .O(gate389inter1));
  and2  gate1359(.a(N1227), .b(N1376), .O(gate389inter2));
  inv1  gate1360(.a(s_68), .O(gate389inter3));
  inv1  gate1361(.a(s_69), .O(gate389inter4));
  nand2 gate1362(.a(gate389inter4), .b(gate389inter3), .O(gate389inter5));
  nor2  gate1363(.a(gate389inter5), .b(gate389inter2), .O(gate389inter6));
  inv1  gate1364(.a(N1376), .O(gate389inter7));
  inv1  gate1365(.a(N1227), .O(gate389inter8));
  nand2 gate1366(.a(gate389inter8), .b(gate389inter7), .O(gate389inter9));
  nand2 gate1367(.a(s_69), .b(gate389inter3), .O(gate389inter10));
  nor2  gate1368(.a(gate389inter10), .b(gate389inter9), .O(gate389inter11));
  nor2  gate1369(.a(gate389inter11), .b(gate389inter6), .O(gate389inter12));
  nand2 gate1370(.a(gate389inter12), .b(gate389inter1), .O(N1471));
nand2 gate390( .a(N1387), .b(N1433), .O(N1472) );
inv1 gate391( .a(N1390), .O(N1475) );
nand2 gate392( .a(N1390), .b(N1240), .O(N1476) );

  xor2  gate1203(.a(N1434), .b(N1389), .O(gate393inter0));
  nand2 gate1204(.a(gate393inter0), .b(s_46), .O(gate393inter1));
  and2  gate1205(.a(N1434), .b(N1389), .O(gate393inter2));
  inv1  gate1206(.a(s_46), .O(gate393inter3));
  inv1  gate1207(.a(s_47), .O(gate393inter4));
  nand2 gate1208(.a(gate393inter4), .b(gate393inter3), .O(gate393inter5));
  nor2  gate1209(.a(gate393inter5), .b(gate393inter2), .O(gate393inter6));
  inv1  gate1210(.a(N1389), .O(gate393inter7));
  inv1  gate1211(.a(N1434), .O(gate393inter8));
  nand2 gate1212(.a(gate393inter8), .b(gate393inter7), .O(gate393inter9));
  nand2 gate1213(.a(s_47), .b(gate393inter3), .O(gate393inter10));
  nor2  gate1214(.a(gate393inter10), .b(gate393inter9), .O(gate393inter11));
  nor2  gate1215(.a(gate393inter11), .b(gate393inter6), .O(gate393inter12));
  nand2 gate1216(.a(gate393inter12), .b(gate393inter1), .O(N1478));
nand2 gate394( .a(N1399), .b(N1439), .O(N1481) );
nand2 gate395( .a(N1397), .b(N1438), .O(N1484) );
nand2 gate396( .a(N939), .b(N1444), .O(N1487) );
nand2 gate397( .a(N935), .b(N1446), .O(N1488) );
nand2 gate398( .a(N943), .b(N1448), .O(N1489) );
inv1 gate399( .a(N1419), .O(N1490) );
inv1 gate400( .a(N1416), .O(N1491) );
nand2 gate401( .a(N947), .b(N1452), .O(N1492) );
nand2 gate402( .a(N955), .b(N1454), .O(N1493) );
nand2 gate403( .a(N951), .b(N1456), .O(N1494) );
nand2 gate404( .a(N969), .b(N1458), .O(N1495) );
nand2 gate405( .a(N977), .b(N1460), .O(N1496) );
nand2 gate406( .a(N998), .b(N1463), .O(N1498) );
inv1 gate407( .a(N1440), .O(N1499) );
nand2 gate408( .a(N965), .b(N1468), .O(N1500) );
nand2 gate409( .a(N973), .b(N1470), .O(N1501) );
nand2 gate410( .a(N994), .b(N1475), .O(N1504) );
inv1 gate411( .a(N1464), .O(N1510) );
nand2 gate412( .a(N1443), .b(N1487), .O(N1513) );
nand2 gate413( .a(N1445), .b(N1488), .O(N1514) );
nand2 gate414( .a(N1447), .b(N1489), .O(N1517) );
nand2 gate415( .a(N1451), .b(N1492), .O(N1520) );

  xor2  gate1273(.a(N1493), .b(N1453), .O(gate416inter0));
  nand2 gate1274(.a(gate416inter0), .b(s_56), .O(gate416inter1));
  and2  gate1275(.a(N1493), .b(N1453), .O(gate416inter2));
  inv1  gate1276(.a(s_56), .O(gate416inter3));
  inv1  gate1277(.a(s_57), .O(gate416inter4));
  nand2 gate1278(.a(gate416inter4), .b(gate416inter3), .O(gate416inter5));
  nor2  gate1279(.a(gate416inter5), .b(gate416inter2), .O(gate416inter6));
  inv1  gate1280(.a(N1453), .O(gate416inter7));
  inv1  gate1281(.a(N1493), .O(gate416inter8));
  nand2 gate1282(.a(gate416inter8), .b(gate416inter7), .O(gate416inter9));
  nand2 gate1283(.a(s_57), .b(gate416inter3), .O(gate416inter10));
  nor2  gate1284(.a(gate416inter10), .b(gate416inter9), .O(gate416inter11));
  nor2  gate1285(.a(gate416inter11), .b(gate416inter6), .O(gate416inter12));
  nand2 gate1286(.a(gate416inter12), .b(gate416inter1), .O(N1521));
nand2 gate417( .a(N1455), .b(N1494), .O(N1522) );

  xor2  gate1329(.a(N1495), .b(N1457), .O(gate418inter0));
  nand2 gate1330(.a(gate418inter0), .b(s_64), .O(gate418inter1));
  and2  gate1331(.a(N1495), .b(N1457), .O(gate418inter2));
  inv1  gate1332(.a(s_64), .O(gate418inter3));
  inv1  gate1333(.a(s_65), .O(gate418inter4));
  nand2 gate1334(.a(gate418inter4), .b(gate418inter3), .O(gate418inter5));
  nor2  gate1335(.a(gate418inter5), .b(gate418inter2), .O(gate418inter6));
  inv1  gate1336(.a(N1457), .O(gate418inter7));
  inv1  gate1337(.a(N1495), .O(gate418inter8));
  nand2 gate1338(.a(gate418inter8), .b(gate418inter7), .O(gate418inter9));
  nand2 gate1339(.a(s_65), .b(gate418inter3), .O(gate418inter10));
  nor2  gate1340(.a(gate418inter10), .b(gate418inter9), .O(gate418inter11));
  nor2  gate1341(.a(gate418inter11), .b(gate418inter6), .O(gate418inter12));
  nand2 gate1342(.a(gate418inter12), .b(gate418inter1), .O(N1526));
nand2 gate419( .a(N1459), .b(N1496), .O(N1527) );
inv1 gate420( .a(N1472), .O(N1528) );
nand2 gate421( .a(N1462), .b(N1498), .O(N1529) );
inv1 gate422( .a(N1478), .O(N1530) );
inv1 gate423( .a(N1481), .O(N1531) );
inv1 gate424( .a(N1484), .O(N1532) );
nand2 gate425( .a(N1471), .b(N1501), .O(N1534) );
nand2 gate426( .a(N1469), .b(N1500), .O(N1537) );
nand2 gate427( .a(N1476), .b(N1504), .O(N1540) );
inv1 gate428( .a(N1513), .O(N1546) );
inv1 gate429( .a(N1521), .O(N1554) );
inv1 gate430( .a(N1526), .O(N1557) );
inv1 gate431( .a(N1520), .O(N1561) );
nand2 gate432( .a(N1484), .b(N1531), .O(N1567) );
nand2 gate433( .a(N1481), .b(N1532), .O(N1568) );
inv1 gate434( .a(N1510), .O(N1569) );
inv1 gate435( .a(N1527), .O(N1571) );
inv1 gate436( .a(N1529), .O(N1576) );
buf1 gate437( .a(N1522), .O(N1588) );
inv1 gate438( .a(N1534), .O(N1591) );
inv1 gate439( .a(N1537), .O(N1593) );
nand2 gate440( .a(N1540), .b(N1530), .O(N1594) );
inv1 gate441( .a(N1540), .O(N1595) );
nand2 gate442( .a(N1567), .b(N1568), .O(N1596) );
buf1 gate443( .a(N1517), .O(N1600) );
buf1 gate444( .a(N1517), .O(N1603) );
buf1 gate445( .a(N1522), .O(N1606) );
buf1 gate446( .a(N1522), .O(N1609) );
buf1 gate447( .a(N1514), .O(N1612) );
buf1 gate448( .a(N1514), .O(N1615) );
buf1 gate449( .a(N1557), .O(N1620) );
buf1 gate450( .a(N1554), .O(N1623) );
inv1 gate451( .a(N1571), .O(N1635) );
nand2 gate452( .a(N1478), .b(N1595), .O(N1636) );
nand2 gate453( .a(N1576), .b(N1569), .O(N1638) );
inv1 gate454( .a(N1576), .O(N1639) );
buf1 gate455( .a(N1561), .O(N1640) );
buf1 gate456( .a(N1561), .O(N1643) );
buf1 gate457( .a(N1546), .O(N1647) );
buf1 gate458( .a(N1546), .O(N1651) );
buf1 gate459( .a(N1554), .O(N1658) );
buf1 gate460( .a(N1557), .O(N1661) );
buf1 gate461( .a(N1557), .O(N1664) );
nand2 gate462( .a(N1596), .b(N893), .O(N1671) );
inv1 gate463( .a(N1596), .O(N1672) );
inv1 gate464( .a(N1600), .O(N1675) );
inv1 gate465( .a(N1603), .O(N1677) );
nand2 gate466( .a(N1606), .b(N1217), .O(N1678) );
inv1 gate467( .a(N1606), .O(N1679) );
nand2 gate468( .a(N1609), .b(N1219), .O(N1680) );
inv1 gate469( .a(N1609), .O(N1681) );
inv1 gate470( .a(N1612), .O(N1682) );
inv1 gate471( .a(N1615), .O(N1683) );
nand2 gate472( .a(N1594), .b(N1636), .O(N1685) );
nand2 gate473( .a(N1510), .b(N1639), .O(N1688) );
buf1 gate474( .a(N1588), .O(N1697) );
buf1 gate475( .a(N1588), .O(N1701) );
nand2 gate476( .a(N643), .b(N1672), .O(N1706) );
inv1 gate477( .a(N1643), .O(N1707) );
nand2 gate478( .a(N1647), .b(N1675), .O(N1708) );
inv1 gate479( .a(N1647), .O(N1709) );
nand2 gate480( .a(N1651), .b(N1677), .O(N1710) );
inv1 gate481( .a(N1651), .O(N1711) );

  xor2  gate993(.a(N1679), .b(N1028), .O(gate482inter0));
  nand2 gate994(.a(gate482inter0), .b(s_16), .O(gate482inter1));
  and2  gate995(.a(N1679), .b(N1028), .O(gate482inter2));
  inv1  gate996(.a(s_16), .O(gate482inter3));
  inv1  gate997(.a(s_17), .O(gate482inter4));
  nand2 gate998(.a(gate482inter4), .b(gate482inter3), .O(gate482inter5));
  nor2  gate999(.a(gate482inter5), .b(gate482inter2), .O(gate482inter6));
  inv1  gate1000(.a(N1028), .O(gate482inter7));
  inv1  gate1001(.a(N1679), .O(gate482inter8));
  nand2 gate1002(.a(gate482inter8), .b(gate482inter7), .O(gate482inter9));
  nand2 gate1003(.a(s_17), .b(gate482inter3), .O(gate482inter10));
  nor2  gate1004(.a(gate482inter10), .b(gate482inter9), .O(gate482inter11));
  nor2  gate1005(.a(gate482inter11), .b(gate482inter6), .O(gate482inter12));
  nand2 gate1006(.a(gate482inter12), .b(gate482inter1), .O(N1712));
nand2 gate483( .a(N1031), .b(N1681), .O(N1713) );
buf1 gate484( .a(N1620), .O(N1714) );
buf1 gate485( .a(N1620), .O(N1717) );
nand2 gate486( .a(N1658), .b(N1593), .O(N1720) );
inv1 gate487( .a(N1658), .O(N1721) );
nand2 gate488( .a(N1638), .b(N1688), .O(N1723) );
inv1 gate489( .a(N1661), .O(N1727) );
inv1 gate490( .a(N1640), .O(N1728) );
inv1 gate491( .a(N1664), .O(N1730) );
buf1 gate492( .a(N1623), .O(N1731) );
buf1 gate493( .a(N1623), .O(N1734) );
nand2 gate494( .a(N1685), .b(N1528), .O(N1740) );
inv1 gate495( .a(N1685), .O(N1741) );
nand2 gate496( .a(N1671), .b(N1706), .O(N1742) );

  xor2  gate1231(.a(N1709), .b(N1600), .O(gate497inter0));
  nand2 gate1232(.a(gate497inter0), .b(s_50), .O(gate497inter1));
  and2  gate1233(.a(N1709), .b(N1600), .O(gate497inter2));
  inv1  gate1234(.a(s_50), .O(gate497inter3));
  inv1  gate1235(.a(s_51), .O(gate497inter4));
  nand2 gate1236(.a(gate497inter4), .b(gate497inter3), .O(gate497inter5));
  nor2  gate1237(.a(gate497inter5), .b(gate497inter2), .O(gate497inter6));
  inv1  gate1238(.a(N1600), .O(gate497inter7));
  inv1  gate1239(.a(N1709), .O(gate497inter8));
  nand2 gate1240(.a(gate497inter8), .b(gate497inter7), .O(gate497inter9));
  nand2 gate1241(.a(s_51), .b(gate497inter3), .O(gate497inter10));
  nor2  gate1242(.a(gate497inter10), .b(gate497inter9), .O(gate497inter11));
  nor2  gate1243(.a(gate497inter11), .b(gate497inter6), .O(gate497inter12));
  nand2 gate1244(.a(gate497inter12), .b(gate497inter1), .O(N1746));
nand2 gate498( .a(N1603), .b(N1711), .O(N1747) );

  xor2  gate1245(.a(N1712), .b(N1678), .O(gate499inter0));
  nand2 gate1246(.a(gate499inter0), .b(s_52), .O(gate499inter1));
  and2  gate1247(.a(N1712), .b(N1678), .O(gate499inter2));
  inv1  gate1248(.a(s_52), .O(gate499inter3));
  inv1  gate1249(.a(s_53), .O(gate499inter4));
  nand2 gate1250(.a(gate499inter4), .b(gate499inter3), .O(gate499inter5));
  nor2  gate1251(.a(gate499inter5), .b(gate499inter2), .O(gate499inter6));
  inv1  gate1252(.a(N1678), .O(gate499inter7));
  inv1  gate1253(.a(N1712), .O(gate499inter8));
  nand2 gate1254(.a(gate499inter8), .b(gate499inter7), .O(gate499inter9));
  nand2 gate1255(.a(s_53), .b(gate499inter3), .O(gate499inter10));
  nor2  gate1256(.a(gate499inter10), .b(gate499inter9), .O(gate499inter11));
  nor2  gate1257(.a(gate499inter11), .b(gate499inter6), .O(gate499inter12));
  nand2 gate1258(.a(gate499inter12), .b(gate499inter1), .O(N1748));
nand2 gate500( .a(N1680), .b(N1713), .O(N1751) );
nand2 gate501( .a(N1537), .b(N1721), .O(N1759) );
inv1 gate502( .a(N1697), .O(N1761) );

  xor2  gate923(.a(N1727), .b(N1697), .O(gate503inter0));
  nand2 gate924(.a(gate503inter0), .b(s_6), .O(gate503inter1));
  and2  gate925(.a(N1727), .b(N1697), .O(gate503inter2));
  inv1  gate926(.a(s_6), .O(gate503inter3));
  inv1  gate927(.a(s_7), .O(gate503inter4));
  nand2 gate928(.a(gate503inter4), .b(gate503inter3), .O(gate503inter5));
  nor2  gate929(.a(gate503inter5), .b(gate503inter2), .O(gate503inter6));
  inv1  gate930(.a(N1697), .O(gate503inter7));
  inv1  gate931(.a(N1727), .O(gate503inter8));
  nand2 gate932(.a(gate503inter8), .b(gate503inter7), .O(gate503inter9));
  nand2 gate933(.a(s_7), .b(gate503inter3), .O(gate503inter10));
  nor2  gate934(.a(gate503inter10), .b(gate503inter9), .O(gate503inter11));
  nor2  gate935(.a(gate503inter11), .b(gate503inter6), .O(gate503inter12));
  nand2 gate936(.a(gate503inter12), .b(gate503inter1), .O(N1762));
inv1 gate504( .a(N1701), .O(N1763) );
nand2 gate505( .a(N1701), .b(N1730), .O(N1764) );
inv1 gate506( .a(N1717), .O(N1768) );
nand2 gate507( .a(N1472), .b(N1741), .O(N1769) );
nand2 gate508( .a(N1723), .b(N1413), .O(N1772) );
inv1 gate509( .a(N1723), .O(N1773) );
nand2 gate510( .a(N1708), .b(N1746), .O(N1774) );
nand2 gate511( .a(N1710), .b(N1747), .O(N1777) );
inv1 gate512( .a(N1731), .O(N1783) );

  xor2  gate1217(.a(N1682), .b(N1731), .O(gate513inter0));
  nand2 gate1218(.a(gate513inter0), .b(s_48), .O(gate513inter1));
  and2  gate1219(.a(N1682), .b(N1731), .O(gate513inter2));
  inv1  gate1220(.a(s_48), .O(gate513inter3));
  inv1  gate1221(.a(s_49), .O(gate513inter4));
  nand2 gate1222(.a(gate513inter4), .b(gate513inter3), .O(gate513inter5));
  nor2  gate1223(.a(gate513inter5), .b(gate513inter2), .O(gate513inter6));
  inv1  gate1224(.a(N1731), .O(gate513inter7));
  inv1  gate1225(.a(N1682), .O(gate513inter8));
  nand2 gate1226(.a(gate513inter8), .b(gate513inter7), .O(gate513inter9));
  nand2 gate1227(.a(s_49), .b(gate513inter3), .O(gate513inter10));
  nor2  gate1228(.a(gate513inter10), .b(gate513inter9), .O(gate513inter11));
  nor2  gate1229(.a(gate513inter11), .b(gate513inter6), .O(gate513inter12));
  nand2 gate1230(.a(gate513inter12), .b(gate513inter1), .O(N1784));
inv1 gate514( .a(N1714), .O(N1785) );
inv1 gate515( .a(N1734), .O(N1786) );
nand2 gate516( .a(N1734), .b(N1683), .O(N1787) );
nand2 gate517( .a(N1720), .b(N1759), .O(N1788) );
nand2 gate518( .a(N1661), .b(N1761), .O(N1791) );
nand2 gate519( .a(N1664), .b(N1763), .O(N1792) );
nand2 gate520( .a(N1751), .b(N1155), .O(N1795) );
inv1 gate521( .a(N1751), .O(N1796) );
nand2 gate522( .a(N1740), .b(N1769), .O(N1798) );
nand2 gate523( .a(N1334), .b(N1773), .O(N1801) );
nand2 gate524( .a(N1742), .b(N290), .O(N1802) );
inv1 gate525( .a(N1748), .O(N1807) );
nand2 gate526( .a(N1748), .b(N1218), .O(N1808) );
nand2 gate527( .a(N1612), .b(N1783), .O(N1809) );
nand2 gate528( .a(N1615), .b(N1786), .O(N1810) );
nand2 gate529( .a(N1791), .b(N1762), .O(N1812) );
nand2 gate530( .a(N1792), .b(N1764), .O(N1815) );
buf1 gate531( .a(N1742), .O(N1818) );

  xor2  gate881(.a(N1490), .b(N1777), .O(gate532inter0));
  nand2 gate882(.a(gate532inter0), .b(s_0), .O(gate532inter1));
  and2  gate883(.a(N1490), .b(N1777), .O(gate532inter2));
  inv1  gate884(.a(s_0), .O(gate532inter3));
  inv1  gate885(.a(s_1), .O(gate532inter4));
  nand2 gate886(.a(gate532inter4), .b(gate532inter3), .O(gate532inter5));
  nor2  gate887(.a(gate532inter5), .b(gate532inter2), .O(gate532inter6));
  inv1  gate888(.a(N1777), .O(gate532inter7));
  inv1  gate889(.a(N1490), .O(gate532inter8));
  nand2 gate890(.a(gate532inter8), .b(gate532inter7), .O(gate532inter9));
  nand2 gate891(.a(s_1), .b(gate532inter3), .O(gate532inter10));
  nor2  gate892(.a(gate532inter10), .b(gate532inter9), .O(gate532inter11));
  nor2  gate893(.a(gate532inter11), .b(gate532inter6), .O(gate532inter12));
  nand2 gate894(.a(gate532inter12), .b(gate532inter1), .O(N1821));
inv1 gate533( .a(N1777), .O(N1822) );
nand2 gate534( .a(N1774), .b(N1491), .O(N1823) );
inv1 gate535( .a(N1774), .O(N1824) );
nand2 gate536( .a(N962), .b(N1796), .O(N1825) );
nand2 gate537( .a(N1788), .b(N1409), .O(N1826) );
inv1 gate538( .a(N1788), .O(N1827) );
nand2 gate539( .a(N1772), .b(N1801), .O(N1830) );
nand2 gate540( .a(N959), .b(N1807), .O(N1837) );
nand2 gate541( .a(N1809), .b(N1784), .O(N1838) );
nand2 gate542( .a(N1810), .b(N1787), .O(N1841) );
nand2 gate543( .a(N1419), .b(N1822), .O(N1848) );
nand2 gate544( .a(N1416), .b(N1824), .O(N1849) );
nand2 gate545( .a(N1795), .b(N1825), .O(N1850) );
nand2 gate546( .a(N1319), .b(N1827), .O(N1852) );
nand2 gate547( .a(N1815), .b(N1707), .O(N1855) );
inv1 gate548( .a(N1815), .O(N1856) );
inv1 gate549( .a(N1818), .O(N1857) );
nand2 gate550( .a(N1798), .b(N290), .O(N1858) );
inv1 gate551( .a(N1812), .O(N1864) );
nand2 gate552( .a(N1812), .b(N1728), .O(N1865) );
buf1 gate553( .a(N1798), .O(N1866) );
buf1 gate554( .a(N1802), .O(N1869) );
buf1 gate555( .a(N1802), .O(N1872) );
nand2 gate556( .a(N1808), .b(N1837), .O(N1875) );
nand2 gate557( .a(N1821), .b(N1848), .O(N1878) );
nand2 gate558( .a(N1823), .b(N1849), .O(N1879) );

  xor2  gate1147(.a(N1768), .b(N1841), .O(gate559inter0));
  nand2 gate1148(.a(gate559inter0), .b(s_38), .O(gate559inter1));
  and2  gate1149(.a(N1768), .b(N1841), .O(gate559inter2));
  inv1  gate1150(.a(s_38), .O(gate559inter3));
  inv1  gate1151(.a(s_39), .O(gate559inter4));
  nand2 gate1152(.a(gate559inter4), .b(gate559inter3), .O(gate559inter5));
  nor2  gate1153(.a(gate559inter5), .b(gate559inter2), .O(gate559inter6));
  inv1  gate1154(.a(N1841), .O(gate559inter7));
  inv1  gate1155(.a(N1768), .O(gate559inter8));
  nand2 gate1156(.a(gate559inter8), .b(gate559inter7), .O(gate559inter9));
  nand2 gate1157(.a(s_39), .b(gate559inter3), .O(gate559inter10));
  nor2  gate1158(.a(gate559inter10), .b(gate559inter9), .O(gate559inter11));
  nor2  gate1159(.a(gate559inter11), .b(gate559inter6), .O(gate559inter12));
  nand2 gate1160(.a(gate559inter12), .b(gate559inter1), .O(N1882));
inv1 gate560( .a(N1841), .O(N1883) );
nand2 gate561( .a(N1826), .b(N1852), .O(N1884) );
nand2 gate562( .a(N1643), .b(N1856), .O(N1885) );

  xor2  gate1049(.a(N290), .b(N1830), .O(gate563inter0));
  nand2 gate1050(.a(gate563inter0), .b(s_24), .O(gate563inter1));
  and2  gate1051(.a(N290), .b(N1830), .O(gate563inter2));
  inv1  gate1052(.a(s_24), .O(gate563inter3));
  inv1  gate1053(.a(s_25), .O(gate563inter4));
  nand2 gate1054(.a(gate563inter4), .b(gate563inter3), .O(gate563inter5));
  nor2  gate1055(.a(gate563inter5), .b(gate563inter2), .O(gate563inter6));
  inv1  gate1056(.a(N1830), .O(gate563inter7));
  inv1  gate1057(.a(N290), .O(gate563inter8));
  nand2 gate1058(.a(gate563inter8), .b(gate563inter7), .O(gate563inter9));
  nand2 gate1059(.a(s_25), .b(gate563inter3), .O(gate563inter10));
  nor2  gate1060(.a(gate563inter10), .b(gate563inter9), .O(gate563inter11));
  nor2  gate1061(.a(gate563inter11), .b(gate563inter6), .O(gate563inter12));
  nand2 gate1062(.a(gate563inter12), .b(gate563inter1), .O(N1889));
inv1 gate564( .a(N1838), .O(N1895) );
nand2 gate565( .a(N1838), .b(N1785), .O(N1896) );
nand2 gate566( .a(N1640), .b(N1864), .O(N1897) );
inv1 gate567( .a(N1850), .O(N1898) );
buf1 gate568( .a(N1830), .O(N1902) );
inv1 gate569( .a(N1878), .O(N1910) );
nand2 gate570( .a(N1717), .b(N1883), .O(N1911) );
inv1 gate571( .a(N1884), .O(N1912) );
nand2 gate572( .a(N1855), .b(N1885), .O(N1913) );
inv1 gate573( .a(N1866), .O(N1915) );

  xor2  gate1007(.a(N919), .b(N1872), .O(gate574inter0));
  nand2 gate1008(.a(gate574inter0), .b(s_18), .O(gate574inter1));
  and2  gate1009(.a(N919), .b(N1872), .O(gate574inter2));
  inv1  gate1010(.a(s_18), .O(gate574inter3));
  inv1  gate1011(.a(s_19), .O(gate574inter4));
  nand2 gate1012(.a(gate574inter4), .b(gate574inter3), .O(gate574inter5));
  nor2  gate1013(.a(gate574inter5), .b(gate574inter2), .O(gate574inter6));
  inv1  gate1014(.a(N1872), .O(gate574inter7));
  inv1  gate1015(.a(N919), .O(gate574inter8));
  nand2 gate1016(.a(gate574inter8), .b(gate574inter7), .O(gate574inter9));
  nand2 gate1017(.a(s_19), .b(gate574inter3), .O(gate574inter10));
  nor2  gate1018(.a(gate574inter10), .b(gate574inter9), .O(gate574inter11));
  nor2  gate1019(.a(gate574inter11), .b(gate574inter6), .O(gate574inter12));
  nand2 gate1020(.a(gate574inter12), .b(gate574inter1), .O(N1919));
inv1 gate575( .a(N1872), .O(N1920) );
nand2 gate576( .a(N1869), .b(N920), .O(N1921) );
inv1 gate577( .a(N1869), .O(N1922) );
inv1 gate578( .a(N1875), .O(N1923) );
nand2 gate579( .a(N1714), .b(N1895), .O(N1924) );
buf1 gate580( .a(N1858), .O(N1927) );
buf1 gate581( .a(N1858), .O(N1930) );
nand2 gate582( .a(N1865), .b(N1897), .O(N1933) );
nand2 gate583( .a(N1882), .b(N1911), .O(N1936) );
inv1 gate584( .a(N1898), .O(N1937) );
inv1 gate585( .a(N1902), .O(N1938) );
nand2 gate586( .a(N679), .b(N1920), .O(N1941) );
nand2 gate587( .a(N676), .b(N1922), .O(N1942) );
buf1 gate588( .a(N1879), .O(N1944) );
inv1 gate589( .a(N1913), .O(N1947) );
buf1 gate590( .a(N1889), .O(N1950) );
buf1 gate591( .a(N1889), .O(N1953) );
buf1 gate592( .a(N1879), .O(N1958) );
nand2 gate593( .a(N1896), .b(N1924), .O(N1961) );
and2 gate594( .a(N1910), .b(N601), .O(N1965) );
and2 gate595( .a(N602), .b(N1912), .O(N1968) );

  xor2  gate1287(.a(N917), .b(N1930), .O(gate596inter0));
  nand2 gate1288(.a(gate596inter0), .b(s_58), .O(gate596inter1));
  and2  gate1289(.a(N917), .b(N1930), .O(gate596inter2));
  inv1  gate1290(.a(s_58), .O(gate596inter3));
  inv1  gate1291(.a(s_59), .O(gate596inter4));
  nand2 gate1292(.a(gate596inter4), .b(gate596inter3), .O(gate596inter5));
  nor2  gate1293(.a(gate596inter5), .b(gate596inter2), .O(gate596inter6));
  inv1  gate1294(.a(N1930), .O(gate596inter7));
  inv1  gate1295(.a(N917), .O(gate596inter8));
  nand2 gate1296(.a(gate596inter8), .b(gate596inter7), .O(gate596inter9));
  nand2 gate1297(.a(s_59), .b(gate596inter3), .O(gate596inter10));
  nor2  gate1298(.a(gate596inter10), .b(gate596inter9), .O(gate596inter11));
  nor2  gate1299(.a(gate596inter11), .b(gate596inter6), .O(gate596inter12));
  nand2 gate1300(.a(gate596inter12), .b(gate596inter1), .O(N1975));
inv1 gate597( .a(N1930), .O(N1976) );
nand2 gate598( .a(N1927), .b(N918), .O(N1977) );
inv1 gate599( .a(N1927), .O(N1978) );
nand2 gate600( .a(N1919), .b(N1941), .O(N1979) );
nand2 gate601( .a(N1921), .b(N1942), .O(N1980) );
inv1 gate602( .a(N1933), .O(N1985) );
inv1 gate603( .a(N1936), .O(N1987) );
inv1 gate604( .a(N1944), .O(N1999) );
nand2 gate605( .a(N1944), .b(N1937), .O(N2000) );
inv1 gate606( .a(N1947), .O(N2002) );
nand2 gate607( .a(N1947), .b(N1499), .O(N2003) );
nand2 gate608( .a(N1953), .b(N1350), .O(N2004) );
inv1 gate609( .a(N1953), .O(N2005) );
nand2 gate610( .a(N1950), .b(N1351), .O(N2006) );
inv1 gate611( .a(N1950), .O(N2007) );
nand2 gate612( .a(N673), .b(N1976), .O(N2008) );
nand2 gate613( .a(N670), .b(N1978), .O(N2009) );
inv1 gate614( .a(N1979), .O(N2012) );
inv1 gate615( .a(N1958), .O(N2013) );
nand2 gate616( .a(N1958), .b(N1923), .O(N2014) );
inv1 gate617( .a(N1961), .O(N2015) );
nand2 gate618( .a(N1961), .b(N1635), .O(N2016) );
inv1 gate619( .a(N1965), .O(N2018) );
inv1 gate620( .a(N1968), .O(N2019) );
nand2 gate621( .a(N1898), .b(N1999), .O(N2020) );
inv1 gate622( .a(N1987), .O(N2021) );
nand2 gate623( .a(N1987), .b(N1591), .O(N2022) );
nand2 gate624( .a(N1440), .b(N2002), .O(N2023) );
nand2 gate625( .a(N1261), .b(N2005), .O(N2024) );
nand2 gate626( .a(N1258), .b(N2007), .O(N2025) );

  xor2  gate1315(.a(N2008), .b(N1975), .O(gate627inter0));
  nand2 gate1316(.a(gate627inter0), .b(s_62), .O(gate627inter1));
  and2  gate1317(.a(N2008), .b(N1975), .O(gate627inter2));
  inv1  gate1318(.a(s_62), .O(gate627inter3));
  inv1  gate1319(.a(s_63), .O(gate627inter4));
  nand2 gate1320(.a(gate627inter4), .b(gate627inter3), .O(gate627inter5));
  nor2  gate1321(.a(gate627inter5), .b(gate627inter2), .O(gate627inter6));
  inv1  gate1322(.a(N1975), .O(gate627inter7));
  inv1  gate1323(.a(N2008), .O(gate627inter8));
  nand2 gate1324(.a(gate627inter8), .b(gate627inter7), .O(gate627inter9));
  nand2 gate1325(.a(s_63), .b(gate627inter3), .O(gate627inter10));
  nor2  gate1326(.a(gate627inter10), .b(gate627inter9), .O(gate627inter11));
  nor2  gate1327(.a(gate627inter11), .b(gate627inter6), .O(gate627inter12));
  nand2 gate1328(.a(gate627inter12), .b(gate627inter1), .O(N2026));
nand2 gate628( .a(N1977), .b(N2009), .O(N2027) );
inv1 gate629( .a(N1980), .O(N2030) );
buf1 gate630( .a(N1980), .O(N2033) );
nand2 gate631( .a(N1875), .b(N2013), .O(N2036) );
nand2 gate632( .a(N1571), .b(N2015), .O(N2037) );

  xor2  gate965(.a(N2000), .b(N2020), .O(gate633inter0));
  nand2 gate966(.a(gate633inter0), .b(s_12), .O(gate633inter1));
  and2  gate967(.a(N2000), .b(N2020), .O(gate633inter2));
  inv1  gate968(.a(s_12), .O(gate633inter3));
  inv1  gate969(.a(s_13), .O(gate633inter4));
  nand2 gate970(.a(gate633inter4), .b(gate633inter3), .O(gate633inter5));
  nor2  gate971(.a(gate633inter5), .b(gate633inter2), .O(gate633inter6));
  inv1  gate972(.a(N2020), .O(gate633inter7));
  inv1  gate973(.a(N2000), .O(gate633inter8));
  nand2 gate974(.a(gate633inter8), .b(gate633inter7), .O(gate633inter9));
  nand2 gate975(.a(s_13), .b(gate633inter3), .O(gate633inter10));
  nor2  gate976(.a(gate633inter10), .b(gate633inter9), .O(gate633inter11));
  nor2  gate977(.a(gate633inter11), .b(gate633inter6), .O(gate633inter12));
  nand2 gate978(.a(gate633inter12), .b(gate633inter1), .O(N2038));
nand2 gate634( .a(N1534), .b(N2021), .O(N2039) );
nand2 gate635( .a(N2023), .b(N2003), .O(N2040) );
nand2 gate636( .a(N2004), .b(N2024), .O(N2041) );
nand2 gate637( .a(N2006), .b(N2025), .O(N2042) );
inv1 gate638( .a(N2026), .O(N2047) );
nand2 gate639( .a(N2036), .b(N2014), .O(N2052) );
nand2 gate640( .a(N2037), .b(N2016), .O(N2055) );
inv1 gate641( .a(N2038), .O(N2060) );
nand2 gate642( .a(N2039), .b(N2022), .O(N2061) );
nand2 gate643( .a(N2040), .b(N290), .O(N2062) );
inv1 gate644( .a(N2041), .O(N2067) );
inv1 gate645( .a(N2027), .O(N2068) );
buf1 gate646( .a(N2027), .O(N2071) );
inv1 gate647( .a(N2052), .O(N2076) );
inv1 gate648( .a(N2055), .O(N2077) );
nand2 gate649( .a(N2060), .b(N290), .O(N2078) );
nand2 gate650( .a(N2061), .b(N290), .O(N2081) );
inv1 gate651( .a(N2042), .O(N2086) );
buf1 gate652( .a(N2042), .O(N2089) );
and2 gate653( .a(N2030), .b(N2068), .O(N2104) );
and2 gate654( .a(N2033), .b(N2068), .O(N2119) );
and2 gate655( .a(N2030), .b(N2071), .O(N2129) );
and2 gate656( .a(N2033), .b(N2071), .O(N2143) );
buf1 gate657( .a(N2062), .O(N2148) );
buf1 gate658( .a(N2062), .O(N2151) );
buf1 gate659( .a(N2078), .O(N2196) );
buf1 gate660( .a(N2078), .O(N2199) );
buf1 gate661( .a(N2081), .O(N2202) );
buf1 gate662( .a(N2081), .O(N2205) );
nand2 gate663( .a(N2151), .b(N915), .O(N2214) );
inv1 gate664( .a(N2151), .O(N2215) );
nand2 gate665( .a(N2148), .b(N916), .O(N2216) );
inv1 gate666( .a(N2148), .O(N2217) );
nand2 gate667( .a(N2199), .b(N1348), .O(N2222) );
inv1 gate668( .a(N2199), .O(N2223) );
nand2 gate669( .a(N2196), .b(N1349), .O(N2224) );
inv1 gate670( .a(N2196), .O(N2225) );
nand2 gate671( .a(N2205), .b(N913), .O(N2226) );
inv1 gate672( .a(N2205), .O(N2227) );
nand2 gate673( .a(N2202), .b(N914), .O(N2228) );
inv1 gate674( .a(N2202), .O(N2229) );
nand2 gate675( .a(N667), .b(N2215), .O(N2230) );

  xor2  gate1189(.a(N2217), .b(N664), .O(gate676inter0));
  nand2 gate1190(.a(gate676inter0), .b(s_44), .O(gate676inter1));
  and2  gate1191(.a(N2217), .b(N664), .O(gate676inter2));
  inv1  gate1192(.a(s_44), .O(gate676inter3));
  inv1  gate1193(.a(s_45), .O(gate676inter4));
  nand2 gate1194(.a(gate676inter4), .b(gate676inter3), .O(gate676inter5));
  nor2  gate1195(.a(gate676inter5), .b(gate676inter2), .O(gate676inter6));
  inv1  gate1196(.a(N664), .O(gate676inter7));
  inv1  gate1197(.a(N2217), .O(gate676inter8));
  nand2 gate1198(.a(gate676inter8), .b(gate676inter7), .O(gate676inter9));
  nand2 gate1199(.a(s_45), .b(gate676inter3), .O(gate676inter10));
  nor2  gate1200(.a(gate676inter10), .b(gate676inter9), .O(gate676inter11));
  nor2  gate1201(.a(gate676inter11), .b(gate676inter6), .O(gate676inter12));
  nand2 gate1202(.a(gate676inter12), .b(gate676inter1), .O(N2231));
nand2 gate677( .a(N1255), .b(N2223), .O(N2232) );
nand2 gate678( .a(N1252), .b(N2225), .O(N2233) );
nand2 gate679( .a(N661), .b(N2227), .O(N2234) );
nand2 gate680( .a(N658), .b(N2229), .O(N2235) );
nand2 gate681( .a(N2214), .b(N2230), .O(N2236) );
nand2 gate682( .a(N2216), .b(N2231), .O(N2237) );

  xor2  gate1259(.a(N2232), .b(N2222), .O(gate683inter0));
  nand2 gate1260(.a(gate683inter0), .b(s_54), .O(gate683inter1));
  and2  gate1261(.a(N2232), .b(N2222), .O(gate683inter2));
  inv1  gate1262(.a(s_54), .O(gate683inter3));
  inv1  gate1263(.a(s_55), .O(gate683inter4));
  nand2 gate1264(.a(gate683inter4), .b(gate683inter3), .O(gate683inter5));
  nor2  gate1265(.a(gate683inter5), .b(gate683inter2), .O(gate683inter6));
  inv1  gate1266(.a(N2222), .O(gate683inter7));
  inv1  gate1267(.a(N2232), .O(gate683inter8));
  nand2 gate1268(.a(gate683inter8), .b(gate683inter7), .O(gate683inter9));
  nand2 gate1269(.a(s_55), .b(gate683inter3), .O(gate683inter10));
  nor2  gate1270(.a(gate683inter10), .b(gate683inter9), .O(gate683inter11));
  nor2  gate1271(.a(gate683inter11), .b(gate683inter6), .O(gate683inter12));
  nand2 gate1272(.a(gate683inter12), .b(gate683inter1), .O(N2240));
nand2 gate684( .a(N2224), .b(N2233), .O(N2241) );
nand2 gate685( .a(N2226), .b(N2234), .O(N2244) );
nand2 gate686( .a(N2228), .b(N2235), .O(N2245) );
inv1 gate687( .a(N2236), .O(N2250) );
inv1 gate688( .a(N2240), .O(N2253) );
inv1 gate689( .a(N2244), .O(N2256) );
inv1 gate690( .a(N2237), .O(N2257) );
buf1 gate691( .a(N2237), .O(N2260) );
inv1 gate692( .a(N2241), .O(N2263) );
and2 gate693( .a(N1164), .b(N2241), .O(N2266) );
inv1 gate694( .a(N2245), .O(N2269) );
and2 gate695( .a(N1168), .b(N2245), .O(N2272) );
nand8 gate696( .a(N2067), .b(N2012), .c(N2047), .d(N2250), .e(N899), .f(N2256), .g(N2253), .h(N903), .O(N2279) );
buf1 gate697( .a(N2266), .O(N2286) );
buf1 gate698( .a(N2266), .O(N2297) );
buf1 gate699( .a(N2272), .O(N2315) );
buf1 gate700( .a(N2272), .O(N2326) );
and2 gate701( .a(N2086), .b(N2257), .O(N2340) );
and2 gate702( .a(N2089), .b(N2257), .O(N2353) );
and2 gate703( .a(N2086), .b(N2260), .O(N2361) );
and2 gate704( .a(N2089), .b(N2260), .O(N2375) );
and4 gate705( .a(N338), .b(N2279), .c(N313), .d(N313), .O(N2384) );
and2 gate706( .a(N1163), .b(N2263), .O(N2385) );
and2 gate707( .a(N1164), .b(N2263), .O(N2386) );
and2 gate708( .a(N1167), .b(N2269), .O(N2426) );
and2 gate709( .a(N1168), .b(N2269), .O(N2427) );
nand5 gate710( .a(N2286), .b(N2315), .c(N2361), .d(N2104), .e(N1171), .O(N2537) );
nand5 gate711( .a(N2286), .b(N2315), .c(N2340), .d(N2129), .e(N1171), .O(N2540) );
nand5 gate712( .a(N2286), .b(N2315), .c(N2340), .d(N2119), .e(N1171), .O(N2543) );
nand5 gate713( .a(N2286), .b(N2315), .c(N2353), .d(N2104), .e(N1171), .O(N2546) );
nand5 gate714( .a(N2297), .b(N2315), .c(N2375), .d(N2119), .e(N1188), .O(N2549) );
nand5 gate715( .a(N2297), .b(N2326), .c(N2361), .d(N2143), .e(N1188), .O(N2552) );
nand5 gate716( .a(N2297), .b(N2326), .c(N2375), .d(N2129), .e(N1188), .O(N2555) );
and5 gate717( .a(N2286), .b(N2315), .c(N2361), .d(N2104), .e(N1171), .O(N2558) );
and5 gate718( .a(N2286), .b(N2315), .c(N2340), .d(N2129), .e(N1171), .O(N2561) );
and5 gate719( .a(N2286), .b(N2315), .c(N2340), .d(N2119), .e(N1171), .O(N2564) );
and5 gate720( .a(N2286), .b(N2315), .c(N2353), .d(N2104), .e(N1171), .O(N2567) );
and5 gate721( .a(N2297), .b(N2315), .c(N2375), .d(N2119), .e(N1188), .O(N2570) );
and5 gate722( .a(N2297), .b(N2326), .c(N2361), .d(N2143), .e(N1188), .O(N2573) );
and5 gate723( .a(N2297), .b(N2326), .c(N2375), .d(N2129), .e(N1188), .O(N2576) );
nand5 gate724( .a(N2286), .b(N2427), .c(N2361), .d(N2129), .e(N1171), .O(N2594) );
nand5 gate725( .a(N2297), .b(N2427), .c(N2361), .d(N2119), .e(N1171), .O(N2597) );
nand5 gate726( .a(N2297), .b(N2427), .c(N2375), .d(N2104), .e(N1171), .O(N2600) );
nand5 gate727( .a(N2297), .b(N2427), .c(N2340), .d(N2143), .e(N1171), .O(N2603) );
nand5 gate728( .a(N2297), .b(N2427), .c(N2353), .d(N2129), .e(N1188), .O(N2606) );
nand5 gate729( .a(N2386), .b(N2326), .c(N2361), .d(N2129), .e(N1188), .O(N2611) );
nand5 gate730( .a(N2386), .b(N2326), .c(N2361), .d(N2119), .e(N1188), .O(N2614) );
nand5 gate731( .a(N2386), .b(N2326), .c(N2375), .d(N2104), .e(N1188), .O(N2617) );
nand5 gate732( .a(N2386), .b(N2326), .c(N2353), .d(N2129), .e(N1188), .O(N2620) );
nand5 gate733( .a(N2297), .b(N2427), .c(N2340), .d(N2104), .e(N926), .O(N2627) );
nand5 gate734( .a(N2386), .b(N2326), .c(N2340), .d(N2104), .e(N926), .O(N2628) );
nand5 gate735( .a(N2386), .b(N2427), .c(N2361), .d(N2104), .e(N926), .O(N2629) );
nand5 gate736( .a(N2386), .b(N2427), .c(N2340), .d(N2129), .e(N926), .O(N2630) );
nand5 gate737( .a(N2386), .b(N2427), .c(N2340), .d(N2119), .e(N926), .O(N2631) );
nand5 gate738( .a(N2386), .b(N2427), .c(N2353), .d(N2104), .e(N926), .O(N2632) );
nand5 gate739( .a(N2386), .b(N2426), .c(N2340), .d(N2104), .e(N926), .O(N2633) );
nand5 gate740( .a(N2385), .b(N2427), .c(N2340), .d(N2104), .e(N926), .O(N2634) );
and5 gate741( .a(N2286), .b(N2427), .c(N2361), .d(N2129), .e(N1171), .O(N2639) );
and5 gate742( .a(N2297), .b(N2427), .c(N2361), .d(N2119), .e(N1171), .O(N2642) );
and5 gate743( .a(N2297), .b(N2427), .c(N2375), .d(N2104), .e(N1171), .O(N2645) );
and5 gate744( .a(N2297), .b(N2427), .c(N2340), .d(N2143), .e(N1171), .O(N2648) );
and5 gate745( .a(N2297), .b(N2427), .c(N2353), .d(N2129), .e(N1188), .O(N2651) );
and5 gate746( .a(N2386), .b(N2326), .c(N2361), .d(N2129), .e(N1188), .O(N2655) );
and5 gate747( .a(N2386), .b(N2326), .c(N2361), .d(N2119), .e(N1188), .O(N2658) );
and5 gate748( .a(N2386), .b(N2326), .c(N2375), .d(N2104), .e(N1188), .O(N2661) );
and5 gate749( .a(N2386), .b(N2326), .c(N2353), .d(N2129), .e(N1188), .O(N2664) );
nand2 gate750( .a(N2558), .b(N534), .O(N2669) );
inv1 gate751( .a(N2558), .O(N2670) );

  xor2  gate1077(.a(N535), .b(N2561), .O(gate752inter0));
  nand2 gate1078(.a(gate752inter0), .b(s_28), .O(gate752inter1));
  and2  gate1079(.a(N535), .b(N2561), .O(gate752inter2));
  inv1  gate1080(.a(s_28), .O(gate752inter3));
  inv1  gate1081(.a(s_29), .O(gate752inter4));
  nand2 gate1082(.a(gate752inter4), .b(gate752inter3), .O(gate752inter5));
  nor2  gate1083(.a(gate752inter5), .b(gate752inter2), .O(gate752inter6));
  inv1  gate1084(.a(N2561), .O(gate752inter7));
  inv1  gate1085(.a(N535), .O(gate752inter8));
  nand2 gate1086(.a(gate752inter8), .b(gate752inter7), .O(gate752inter9));
  nand2 gate1087(.a(s_29), .b(gate752inter3), .O(gate752inter10));
  nor2  gate1088(.a(gate752inter10), .b(gate752inter9), .O(gate752inter11));
  nor2  gate1089(.a(gate752inter11), .b(gate752inter6), .O(gate752inter12));
  nand2 gate1090(.a(gate752inter12), .b(gate752inter1), .O(N2671));
inv1 gate753( .a(N2561), .O(N2672) );
nand2 gate754( .a(N2564), .b(N536), .O(N2673) );
inv1 gate755( .a(N2564), .O(N2674) );

  xor2  gate1091(.a(N537), .b(N2567), .O(gate756inter0));
  nand2 gate1092(.a(gate756inter0), .b(s_30), .O(gate756inter1));
  and2  gate1093(.a(N537), .b(N2567), .O(gate756inter2));
  inv1  gate1094(.a(s_30), .O(gate756inter3));
  inv1  gate1095(.a(s_31), .O(gate756inter4));
  nand2 gate1096(.a(gate756inter4), .b(gate756inter3), .O(gate756inter5));
  nor2  gate1097(.a(gate756inter5), .b(gate756inter2), .O(gate756inter6));
  inv1  gate1098(.a(N2567), .O(gate756inter7));
  inv1  gate1099(.a(N537), .O(gate756inter8));
  nand2 gate1100(.a(gate756inter8), .b(gate756inter7), .O(gate756inter9));
  nand2 gate1101(.a(s_31), .b(gate756inter3), .O(gate756inter10));
  nor2  gate1102(.a(gate756inter10), .b(gate756inter9), .O(gate756inter11));
  nor2  gate1103(.a(gate756inter11), .b(gate756inter6), .O(gate756inter12));
  nand2 gate1104(.a(gate756inter12), .b(gate756inter1), .O(N2675));
inv1 gate757( .a(N2567), .O(N2676) );
nand2 gate758( .a(N2570), .b(N543), .O(N2682) );
inv1 gate759( .a(N2570), .O(N2683) );

  xor2  gate1371(.a(N548), .b(N2573), .O(gate760inter0));
  nand2 gate1372(.a(gate760inter0), .b(s_70), .O(gate760inter1));
  and2  gate1373(.a(N548), .b(N2573), .O(gate760inter2));
  inv1  gate1374(.a(s_70), .O(gate760inter3));
  inv1  gate1375(.a(s_71), .O(gate760inter4));
  nand2 gate1376(.a(gate760inter4), .b(gate760inter3), .O(gate760inter5));
  nor2  gate1377(.a(gate760inter5), .b(gate760inter2), .O(gate760inter6));
  inv1  gate1378(.a(N2573), .O(gate760inter7));
  inv1  gate1379(.a(N548), .O(gate760inter8));
  nand2 gate1380(.a(gate760inter8), .b(gate760inter7), .O(gate760inter9));
  nand2 gate1381(.a(s_71), .b(gate760inter3), .O(gate760inter10));
  nor2  gate1382(.a(gate760inter10), .b(gate760inter9), .O(gate760inter11));
  nor2  gate1383(.a(gate760inter11), .b(gate760inter6), .O(gate760inter12));
  nand2 gate1384(.a(gate760inter12), .b(gate760inter1), .O(N2688));
inv1 gate761( .a(N2573), .O(N2689) );

  xor2  gate979(.a(N549), .b(N2576), .O(gate762inter0));
  nand2 gate980(.a(gate762inter0), .b(s_14), .O(gate762inter1));
  and2  gate981(.a(N549), .b(N2576), .O(gate762inter2));
  inv1  gate982(.a(s_14), .O(gate762inter3));
  inv1  gate983(.a(s_15), .O(gate762inter4));
  nand2 gate984(.a(gate762inter4), .b(gate762inter3), .O(gate762inter5));
  nor2  gate985(.a(gate762inter5), .b(gate762inter2), .O(gate762inter6));
  inv1  gate986(.a(N2576), .O(gate762inter7));
  inv1  gate987(.a(N549), .O(gate762inter8));
  nand2 gate988(.a(gate762inter8), .b(gate762inter7), .O(gate762inter9));
  nand2 gate989(.a(s_15), .b(gate762inter3), .O(gate762inter10));
  nor2  gate990(.a(gate762inter10), .b(gate762inter9), .O(gate762inter11));
  nor2  gate991(.a(gate762inter11), .b(gate762inter6), .O(gate762inter12));
  nand2 gate992(.a(gate762inter12), .b(gate762inter1), .O(N2690));
inv1 gate763( .a(N2576), .O(N2691) );
and8 gate764( .a(N2627), .b(N2628), .c(N2629), .d(N2630), .e(N2631), .f(N2632), .g(N2633), .h(N2634), .O(N2710) );
nand2 gate765( .a(N343), .b(N2670), .O(N2720) );
nand2 gate766( .a(N346), .b(N2672), .O(N2721) );
nand2 gate767( .a(N349), .b(N2674), .O(N2722) );
nand2 gate768( .a(N352), .b(N2676), .O(N2723) );
nand2 gate769( .a(N2639), .b(N538), .O(N2724) );
inv1 gate770( .a(N2639), .O(N2725) );
nand2 gate771( .a(N2642), .b(N539), .O(N2726) );
inv1 gate772( .a(N2642), .O(N2727) );
nand2 gate773( .a(N2645), .b(N540), .O(N2728) );
inv1 gate774( .a(N2645), .O(N2729) );
nand2 gate775( .a(N2648), .b(N541), .O(N2730) );
inv1 gate776( .a(N2648), .O(N2731) );
nand2 gate777( .a(N2651), .b(N542), .O(N2732) );
inv1 gate778( .a(N2651), .O(N2733) );
nand2 gate779( .a(N370), .b(N2683), .O(N2734) );
nand2 gate780( .a(N2655), .b(N544), .O(N2735) );
inv1 gate781( .a(N2655), .O(N2736) );
nand2 gate782( .a(N2658), .b(N545), .O(N2737) );
inv1 gate783( .a(N2658), .O(N2738) );

  xor2  gate937(.a(N546), .b(N2661), .O(gate784inter0));
  nand2 gate938(.a(gate784inter0), .b(s_8), .O(gate784inter1));
  and2  gate939(.a(N546), .b(N2661), .O(gate784inter2));
  inv1  gate940(.a(s_8), .O(gate784inter3));
  inv1  gate941(.a(s_9), .O(gate784inter4));
  nand2 gate942(.a(gate784inter4), .b(gate784inter3), .O(gate784inter5));
  nor2  gate943(.a(gate784inter5), .b(gate784inter2), .O(gate784inter6));
  inv1  gate944(.a(N2661), .O(gate784inter7));
  inv1  gate945(.a(N546), .O(gate784inter8));
  nand2 gate946(.a(gate784inter8), .b(gate784inter7), .O(gate784inter9));
  nand2 gate947(.a(s_9), .b(gate784inter3), .O(gate784inter10));
  nor2  gate948(.a(gate784inter10), .b(gate784inter9), .O(gate784inter11));
  nor2  gate949(.a(gate784inter11), .b(gate784inter6), .O(gate784inter12));
  nand2 gate950(.a(gate784inter12), .b(gate784inter1), .O(N2739));
inv1 gate785( .a(N2661), .O(N2740) );
nand2 gate786( .a(N2664), .b(N547), .O(N2741) );
inv1 gate787( .a(N2664), .O(N2742) );
nand2 gate788( .a(N385), .b(N2689), .O(N2743) );
nand2 gate789( .a(N388), .b(N2691), .O(N2744) );
nand8 gate790( .a(N2537), .b(N2540), .c(N2543), .d(N2546), .e(N2594), .f(N2597), .g(N2600), .h(N2603), .O(N2745) );
nand8 gate791( .a(N2606), .b(N2549), .c(N2611), .d(N2614), .e(N2617), .f(N2620), .g(N2552), .h(N2555), .O(N2746) );
and8 gate792( .a(N2537), .b(N2540), .c(N2543), .d(N2546), .e(N2594), .f(N2597), .g(N2600), .h(N2603), .O(N2747) );
and8 gate793( .a(N2606), .b(N2549), .c(N2611), .d(N2614), .e(N2617), .f(N2620), .g(N2552), .h(N2555), .O(N2750) );
nand2 gate794( .a(N2669), .b(N2720), .O(N2753) );
nand2 gate795( .a(N2671), .b(N2721), .O(N2754) );
nand2 gate796( .a(N2673), .b(N2722), .O(N2755) );
nand2 gate797( .a(N2675), .b(N2723), .O(N2756) );
nand2 gate798( .a(N355), .b(N2725), .O(N2757) );
nand2 gate799( .a(N358), .b(N2727), .O(N2758) );
nand2 gate800( .a(N361), .b(N2729), .O(N2759) );
nand2 gate801( .a(N364), .b(N2731), .O(N2760) );
nand2 gate802( .a(N367), .b(N2733), .O(N2761) );
nand2 gate803( .a(N2682), .b(N2734), .O(N2762) );
nand2 gate804( .a(N373), .b(N2736), .O(N2763) );
nand2 gate805( .a(N376), .b(N2738), .O(N2764) );

  xor2  gate1343(.a(N2740), .b(N379), .O(gate806inter0));
  nand2 gate1344(.a(gate806inter0), .b(s_66), .O(gate806inter1));
  and2  gate1345(.a(N2740), .b(N379), .O(gate806inter2));
  inv1  gate1346(.a(s_66), .O(gate806inter3));
  inv1  gate1347(.a(s_67), .O(gate806inter4));
  nand2 gate1348(.a(gate806inter4), .b(gate806inter3), .O(gate806inter5));
  nor2  gate1349(.a(gate806inter5), .b(gate806inter2), .O(gate806inter6));
  inv1  gate1350(.a(N379), .O(gate806inter7));
  inv1  gate1351(.a(N2740), .O(gate806inter8));
  nand2 gate1352(.a(gate806inter8), .b(gate806inter7), .O(gate806inter9));
  nand2 gate1353(.a(s_67), .b(gate806inter3), .O(gate806inter10));
  nor2  gate1354(.a(gate806inter10), .b(gate806inter9), .O(gate806inter11));
  nor2  gate1355(.a(gate806inter11), .b(gate806inter6), .O(gate806inter12));
  nand2 gate1356(.a(gate806inter12), .b(gate806inter1), .O(N2765));
nand2 gate807( .a(N382), .b(N2742), .O(N2766) );
nand2 gate808( .a(N2688), .b(N2743), .O(N2767) );
nand2 gate809( .a(N2690), .b(N2744), .O(N2768) );
and2 gate810( .a(N2745), .b(N275), .O(N2773) );
and2 gate811( .a(N2746), .b(N276), .O(N2776) );
nand2 gate812( .a(N2724), .b(N2757), .O(N2779) );
nand2 gate813( .a(N2726), .b(N2758), .O(N2780) );
nand2 gate814( .a(N2728), .b(N2759), .O(N2781) );
nand2 gate815( .a(N2730), .b(N2760), .O(N2782) );
nand2 gate816( .a(N2732), .b(N2761), .O(N2783) );

  xor2  gate951(.a(N2763), .b(N2735), .O(gate817inter0));
  nand2 gate952(.a(gate817inter0), .b(s_10), .O(gate817inter1));
  and2  gate953(.a(N2763), .b(N2735), .O(gate817inter2));
  inv1  gate954(.a(s_10), .O(gate817inter3));
  inv1  gate955(.a(s_11), .O(gate817inter4));
  nand2 gate956(.a(gate817inter4), .b(gate817inter3), .O(gate817inter5));
  nor2  gate957(.a(gate817inter5), .b(gate817inter2), .O(gate817inter6));
  inv1  gate958(.a(N2735), .O(gate817inter7));
  inv1  gate959(.a(N2763), .O(gate817inter8));
  nand2 gate960(.a(gate817inter8), .b(gate817inter7), .O(gate817inter9));
  nand2 gate961(.a(s_11), .b(gate817inter3), .O(gate817inter10));
  nor2  gate962(.a(gate817inter10), .b(gate817inter9), .O(gate817inter11));
  nor2  gate963(.a(gate817inter11), .b(gate817inter6), .O(gate817inter12));
  nand2 gate964(.a(gate817inter12), .b(gate817inter1), .O(N2784));
nand2 gate818( .a(N2737), .b(N2764), .O(N2785) );
nand2 gate819( .a(N2739), .b(N2765), .O(N2786) );
nand2 gate820( .a(N2741), .b(N2766), .O(N2787) );
and3 gate821( .a(N2747), .b(N2750), .c(N2710), .O(N2788) );
nand2 gate822( .a(N2747), .b(N2750), .O(N2789) );
and4 gate823( .a(N338), .b(N2279), .c(N99), .d(N2788), .O(N2800) );
nand2 gate824( .a(N2773), .b(N2018), .O(N2807) );
inv1 gate825( .a(N2773), .O(N2808) );
nand2 gate826( .a(N2776), .b(N2019), .O(N2809) );
inv1 gate827( .a(N2776), .O(N2810) );
nor2 gate828( .a(N2384), .b(N2800), .O(N2811) );
and3 gate829( .a(N897), .b(N283), .c(N2789), .O(N2812) );
and3 gate830( .a(N76), .b(N283), .c(N2789), .O(N2815) );
and3 gate831( .a(N82), .b(N283), .c(N2789), .O(N2818) );
and3 gate832( .a(N85), .b(N283), .c(N2789), .O(N2821) );
and3 gate833( .a(N898), .b(N283), .c(N2789), .O(N2824) );
nand2 gate834( .a(N1965), .b(N2808), .O(N2827) );
nand2 gate835( .a(N1968), .b(N2810), .O(N2828) );
and3 gate836( .a(N79), .b(N283), .c(N2789), .O(N2829) );
nand2 gate837( .a(N2807), .b(N2827), .O(N2843) );
nand2 gate838( .a(N2809), .b(N2828), .O(N2846) );

  xor2  gate1301(.a(N2076), .b(N2812), .O(gate839inter0));
  nand2 gate1302(.a(gate839inter0), .b(s_60), .O(gate839inter1));
  and2  gate1303(.a(N2076), .b(N2812), .O(gate839inter2));
  inv1  gate1304(.a(s_60), .O(gate839inter3));
  inv1  gate1305(.a(s_61), .O(gate839inter4));
  nand2 gate1306(.a(gate839inter4), .b(gate839inter3), .O(gate839inter5));
  nor2  gate1307(.a(gate839inter5), .b(gate839inter2), .O(gate839inter6));
  inv1  gate1308(.a(N2812), .O(gate839inter7));
  inv1  gate1309(.a(N2076), .O(gate839inter8));
  nand2 gate1310(.a(gate839inter8), .b(gate839inter7), .O(gate839inter9));
  nand2 gate1311(.a(s_61), .b(gate839inter3), .O(gate839inter10));
  nor2  gate1312(.a(gate839inter10), .b(gate839inter9), .O(gate839inter11));
  nor2  gate1313(.a(gate839inter11), .b(gate839inter6), .O(gate839inter12));
  nand2 gate1314(.a(gate839inter12), .b(gate839inter1), .O(N2850));
nand2 gate840( .a(N2815), .b(N2077), .O(N2851) );
nand2 gate841( .a(N2818), .b(N1915), .O(N2852) );
nand2 gate842( .a(N2821), .b(N1857), .O(N2853) );

  xor2  gate1063(.a(N1938), .b(N2824), .O(gate843inter0));
  nand2 gate1064(.a(gate843inter0), .b(s_26), .O(gate843inter1));
  and2  gate1065(.a(N1938), .b(N2824), .O(gate843inter2));
  inv1  gate1066(.a(s_26), .O(gate843inter3));
  inv1  gate1067(.a(s_27), .O(gate843inter4));
  nand2 gate1068(.a(gate843inter4), .b(gate843inter3), .O(gate843inter5));
  nor2  gate1069(.a(gate843inter5), .b(gate843inter2), .O(gate843inter6));
  inv1  gate1070(.a(N2824), .O(gate843inter7));
  inv1  gate1071(.a(N1938), .O(gate843inter8));
  nand2 gate1072(.a(gate843inter8), .b(gate843inter7), .O(gate843inter9));
  nand2 gate1073(.a(s_27), .b(gate843inter3), .O(gate843inter10));
  nor2  gate1074(.a(gate843inter10), .b(gate843inter9), .O(gate843inter11));
  nor2  gate1075(.a(gate843inter11), .b(gate843inter6), .O(gate843inter12));
  nand2 gate1076(.a(gate843inter12), .b(gate843inter1), .O(N2854));
inv1 gate844( .a(N2812), .O(N2857) );
inv1 gate845( .a(N2815), .O(N2858) );
inv1 gate846( .a(N2818), .O(N2859) );
inv1 gate847( .a(N2821), .O(N2860) );
inv1 gate848( .a(N2824), .O(N2861) );
inv1 gate849( .a(N2829), .O(N2862) );
nand2 gate850( .a(N2829), .b(N1985), .O(N2863) );
nand2 gate851( .a(N2052), .b(N2857), .O(N2866) );
nand2 gate852( .a(N2055), .b(N2858), .O(N2867) );
nand2 gate853( .a(N1866), .b(N2859), .O(N2868) );
nand2 gate854( .a(N1818), .b(N2860), .O(N2869) );
nand2 gate855( .a(N1902), .b(N2861), .O(N2870) );
nand2 gate856( .a(N2843), .b(N886), .O(N2871) );
inv1 gate857( .a(N2843), .O(N2872) );

  xor2  gate1133(.a(N887), .b(N2846), .O(gate858inter0));
  nand2 gate1134(.a(gate858inter0), .b(s_36), .O(gate858inter1));
  and2  gate1135(.a(N887), .b(N2846), .O(gate858inter2));
  inv1  gate1136(.a(s_36), .O(gate858inter3));
  inv1  gate1137(.a(s_37), .O(gate858inter4));
  nand2 gate1138(.a(gate858inter4), .b(gate858inter3), .O(gate858inter5));
  nor2  gate1139(.a(gate858inter5), .b(gate858inter2), .O(gate858inter6));
  inv1  gate1140(.a(N2846), .O(gate858inter7));
  inv1  gate1141(.a(N887), .O(gate858inter8));
  nand2 gate1142(.a(gate858inter8), .b(gate858inter7), .O(gate858inter9));
  nand2 gate1143(.a(s_37), .b(gate858inter3), .O(gate858inter10));
  nor2  gate1144(.a(gate858inter10), .b(gate858inter9), .O(gate858inter11));
  nor2  gate1145(.a(gate858inter11), .b(gate858inter6), .O(gate858inter12));
  nand2 gate1146(.a(gate858inter12), .b(gate858inter1), .O(N2873));
inv1 gate859( .a(N2846), .O(N2874) );
nand2 gate860( .a(N1933), .b(N2862), .O(N2875) );
nand2 gate861( .a(N2866), .b(N2850), .O(N2876) );
nand2 gate862( .a(N2867), .b(N2851), .O(N2877) );
nand2 gate863( .a(N2868), .b(N2852), .O(N2878) );
nand2 gate864( .a(N2869), .b(N2853), .O(N2879) );
nand2 gate865( .a(N2870), .b(N2854), .O(N2880) );

  xor2  gate909(.a(N2872), .b(N682), .O(gate866inter0));
  nand2 gate910(.a(gate866inter0), .b(s_4), .O(gate866inter1));
  and2  gate911(.a(N2872), .b(N682), .O(gate866inter2));
  inv1  gate912(.a(s_4), .O(gate866inter3));
  inv1  gate913(.a(s_5), .O(gate866inter4));
  nand2 gate914(.a(gate866inter4), .b(gate866inter3), .O(gate866inter5));
  nor2  gate915(.a(gate866inter5), .b(gate866inter2), .O(gate866inter6));
  inv1  gate916(.a(N682), .O(gate866inter7));
  inv1  gate917(.a(N2872), .O(gate866inter8));
  nand2 gate918(.a(gate866inter8), .b(gate866inter7), .O(gate866inter9));
  nand2 gate919(.a(s_5), .b(gate866inter3), .O(gate866inter10));
  nor2  gate920(.a(gate866inter10), .b(gate866inter9), .O(gate866inter11));
  nor2  gate921(.a(gate866inter11), .b(gate866inter6), .O(gate866inter12));
  nand2 gate922(.a(gate866inter12), .b(gate866inter1), .O(N2881));
nand2 gate867( .a(N685), .b(N2874), .O(N2882) );
nand2 gate868( .a(N2875), .b(N2863), .O(N2883) );
and2 gate869( .a(N2876), .b(N550), .O(N2886) );
and2 gate870( .a(N551), .b(N2877), .O(N2887) );
and2 gate871( .a(N553), .b(N2878), .O(N2888) );
and2 gate872( .a(N2879), .b(N554), .O(N2889) );
and2 gate873( .a(N555), .b(N2880), .O(N2890) );
nand2 gate874( .a(N2871), .b(N2881), .O(N2891) );
nand2 gate875( .a(N2873), .b(N2882), .O(N2892) );
nand2 gate876( .a(N2883), .b(N1461), .O(N2895) );
inv1 gate877( .a(N2883), .O(N2896) );
nand2 gate878( .a(N1383), .b(N2896), .O(N2897) );
nand2 gate879( .a(N2895), .b(N2897), .O(N2898) );
and2 gate880( .a(N2898), .b(N552), .O(N2899) );

endmodule