module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);

input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;//RE__PI;

input s_0,s_1;//RE__ALLOW(00,01,10,11);
input s_2,s_3;//RE__ALLOW(00,01,10,11);
input s_4,s_5;//RE__ALLOW(00,01,10,11);
input s_6,s_7;//RE__ALLOW(00,01,10,11);
input s_8,s_9;//RE__ALLOW(00,01,10,11);
input s_10,s_11;//RE__ALLOW(00,01,10,11);
input s_12,s_13;//RE__ALLOW(00,01,10,11);
input s_14,s_15;//RE__ALLOW(00,01,10,11);
input s_16,s_17;//RE__ALLOW(00,01,10,11);
input s_18,s_19;//RE__ALLOW(00,01,10,11);
input s_20,s_21;//RE__ALLOW(00,01,10,11);
input s_22,s_23;//RE__ALLOW(00,01,10,11);
input s_24,s_25;//RE__ALLOW(00,01,10,11);
input s_26,s_27;//RE__ALLOW(00,01,10,11);
input s_28,s_29;//RE__ALLOW(00,01,10,11);
input s_30,s_31;//RE__ALLOW(00,01,10,11);
input s_32,s_33;//RE__ALLOW(00,01,10,11);
input s_34,s_35;//RE__ALLOW(00,01,10,11);
input s_36,s_37;//RE__ALLOW(00,01,10,11);
input s_38,s_39;//RE__ALLOW(00,01,10,11);
input s_40,s_41;//RE__ALLOW(00,01,10,11);
input s_42,s_43;//RE__ALLOW(00,01,10,11);
input s_44,s_45;//RE__ALLOW(00,01,10,11);
input s_46,s_47;//RE__ALLOW(00,01,10,11);
input s_48,s_49;//RE__ALLOW(00,01,10,11);
input s_50,s_51;//RE__ALLOW(00,01,10,11);
input s_52,s_53;//RE__ALLOW(00,01,10,11);
input s_54,s_55;//RE__ALLOW(00,01,10,11);
input s_56,s_57;//RE__ALLOW(00,01,10,11);
input s_58,s_59;//RE__ALLOW(00,01,10,11);
input s_60,s_61;//RE__ALLOW(00,01,10,11);
input s_62,s_63;//RE__ALLOW(00,01,10,11);
input s_64,s_65;//RE__ALLOW(00,01,10,11);
input s_66,s_67;//RE__ALLOW(00,01,10,11);
input s_68,s_69;//RE__ALLOW(00,01,10,11);
input s_70,s_71;//RE__ALLOW(00,01,10,11);
input s_72,s_73;//RE__ALLOW(00,01,10,11);
input s_74,s_75;//RE__ALLOW(00,01,10,11);
input s_76,s_77;//RE__ALLOW(00,01,10,11);
input s_78,s_79;//RE__ALLOW(00,01,10,11);
input s_80,s_81;//RE__ALLOW(00,01,10,11);
input s_82,s_83;//RE__ALLOW(00,01,10,11);
input s_84,s_85;//RE__ALLOW(00,01,10,11);
input s_86,s_87;//RE__ALLOW(00,01,10,11);
input s_88,s_89;//RE__ALLOW(00,01,10,11);
input s_90,s_91;//RE__ALLOW(00,01,10,11);
input s_92,s_93;//RE__ALLOW(00,01,10,11);
input s_94,s_95;//RE__ALLOW(00,01,10,11);
input s_96,s_97;//RE__ALLOW(00,01,10,11);
input s_98,s_99;//RE__ALLOW(00,01,10,11);
input s_100,s_101;//RE__ALLOW(00,01,10,11);
input s_102,s_103;//RE__ALLOW(00,01,10,11);
input s_104,s_105;//RE__ALLOW(00,01,10,11);
input s_106,s_107;//RE__ALLOW(00,01,10,11);
input s_108,s_109;//RE__ALLOW(00,01,10,11);
input s_110,s_111;//RE__ALLOW(00,01,10,11);
input s_112,s_113;//RE__ALLOW(00,01,10,11);
input s_114,s_115;//RE__ALLOW(00,01,10,11);
input s_116,s_117;//RE__ALLOW(00,01,10,11);
input s_118,s_119;//RE__ALLOW(00,01,10,11);
input s_120,s_121;//RE__ALLOW(00,01,10,11);
input s_122,s_123;//RE__ALLOW(00,01,10,11);
input s_124,s_125;//RE__ALLOW(00,01,10,11);
input s_126,s_127;//RE__ALLOW(00,01,10,11);
input s_128,s_129;//RE__ALLOW(00,01,10,11);
input s_130,s_131;//RE__ALLOW(00,01,10,11);
input s_132,s_133;//RE__ALLOW(00,01,10,11);
input s_134,s_135;//RE__ALLOW(00,01,10,11);
input s_136,s_137;//RE__ALLOW(00,01,10,11);
input s_138,s_139;//RE__ALLOW(00,01,10,11);
input s_140,s_141;//RE__ALLOW(00,01,10,11);
input s_142,s_143;//RE__ALLOW(00,01,10,11);
input s_144,s_145;//RE__ALLOW(00,01,10,11);
input s_146,s_147;//RE__ALLOW(00,01,10,11);
input s_148,s_149;//RE__ALLOW(00,01,10,11);
input s_150,s_151;//RE__ALLOW(00,01,10,11);
input s_152,s_153;//RE__ALLOW(00,01,10,11);
input s_154,s_155;//RE__ALLOW(00,01,10,11);
input s_156,s_157;//RE__ALLOW(00,01,10,11);
input s_158,s_159;//RE__ALLOW(00,01,10,11);
input s_160,s_161;//RE__ALLOW(00,01,10,11);
input s_162,s_163;//RE__ALLOW(00,01,10,11);
input s_164,s_165;//RE__ALLOW(00,01,10,11);
input s_166,s_167;//RE__ALLOW(00,01,10,11);
input s_168,s_169;//RE__ALLOW(00,01,10,11);
input s_170,s_171;//RE__ALLOW(00,01,10,11);
input s_172,s_173;//RE__ALLOW(00,01,10,11);
input s_174,s_175;//RE__ALLOW(00,01,10,11);
input s_176,s_177;//RE__ALLOW(00,01,10,11);
input s_178,s_179;//RE__ALLOW(00,01,10,11);
input s_180,s_181;//RE__ALLOW(00,01,10,11);
input s_182,s_183;//RE__ALLOW(00,01,10,11);
input s_184,s_185;//RE__ALLOW(00,01,10,11);
input s_186,s_187;//RE__ALLOW(00,01,10,11);
input s_188,s_189;//RE__ALLOW(00,01,10,11);
input s_190,s_191;//RE__ALLOW(00,01,10,11);
input s_192,s_193;//RE__ALLOW(00,01,10,11);
input s_194,s_195;//RE__ALLOW(00,01,10,11);
input s_196,s_197;//RE__ALLOW(00,01,10,11);
input s_198,s_199;//RE__ALLOW(00,01,10,11);
input s_200,s_201;//RE__ALLOW(00,01,10,11);
input s_202,s_203;//RE__ALLOW(00,01,10,11);
input s_204,s_205;//RE__ALLOW(00,01,10,11);
input s_206,s_207;//RE__ALLOW(00,01,10,11);
input s_208,s_209;//RE__ALLOW(00,01,10,11);
input s_210,s_211;//RE__ALLOW(00,01,10,11);
input s_212,s_213;//RE__ALLOW(00,01,10,11);
input s_214,s_215;//RE__ALLOW(00,01,10,11);
input s_216,s_217;//RE__ALLOW(00,01,10,11);
input s_218,s_219;//RE__ALLOW(00,01,10,11);
input s_220,s_221;//RE__ALLOW(00,01,10,11);
input s_222,s_223;//RE__ALLOW(00,01,10,11);
input s_224,s_225;//RE__ALLOW(00,01,10,11);
input s_226,s_227;//RE__ALLOW(00,01,10,11);
input s_228,s_229;//RE__ALLOW(00,01,10,11);
input s_230,s_231;//RE__ALLOW(00,01,10,11);
input s_232,s_233;//RE__ALLOW(00,01,10,11);
input s_234,s_235;//RE__ALLOW(00,01,10,11);
input s_236,s_237;//RE__ALLOW(00,01,10,11);
input s_238,s_239;//RE__ALLOW(00,01,10,11);
input s_240,s_241;//RE__ALLOW(00,01,10,11);
input s_242,s_243;//RE__ALLOW(00,01,10,11);
input s_244,s_245;//RE__ALLOW(00,01,10,11);
input s_246,s_247;//RE__ALLOW(00,01,10,11);
input s_248,s_249;//RE__ALLOW(00,01,10,11);
input s_250,s_251;//RE__ALLOW(00,01,10,11);
input s_252,s_253;//RE__ALLOW(00,01,10,11);
input s_254,s_255;//RE__ALLOW(00,01,10,11);
input s_256,s_257;//RE__ALLOW(00,01,10,11);
input s_258,s_259;//RE__ALLOW(00,01,10,11);
input s_260,s_261;//RE__ALLOW(00,01,10,11);
input s_262,s_263;//RE__ALLOW(00,01,10,11);
input s_264,s_265;//RE__ALLOW(00,01,10,11);
input s_266,s_267;//RE__ALLOW(00,01,10,11);
input s_268,s_269;//RE__ALLOW(00,01,10,11);
input s_270,s_271;//RE__ALLOW(00,01,10,11);
input s_272,s_273;//RE__ALLOW(00,01,10,11);
input s_274,s_275;//RE__ALLOW(00,01,10,11);
input s_276,s_277;//RE__ALLOW(00,01,10,11);
input s_278,s_279;//RE__ALLOW(00,01,10,11);
input s_280,s_281;//RE__ALLOW(00,01,10,11);
input s_282,s_283;//RE__ALLOW(00,01,10,11);
input s_284,s_285;//RE__ALLOW(00,01,10,11);
input s_286,s_287;//RE__ALLOW(00,01,10,11);
input s_288,s_289;//RE__ALLOW(00,01,10,11);
input s_290,s_291;//RE__ALLOW(00,01,10,11);
input s_292,s_293;//RE__ALLOW(00,01,10,11);
input s_294,s_295;//RE__ALLOW(00,01,10,11);
input s_296,s_297;//RE__ALLOW(00,01,10,11);
input s_298,s_299;//RE__ALLOW(00,01,10,11);
input s_300,s_301;//RE__ALLOW(00,01,10,11);
input s_302,s_303;//RE__ALLOW(00,01,10,11);
input s_304,s_305;//RE__ALLOW(00,01,10,11);
input s_306,s_307;//RE__ALLOW(00,01,10,11);
input s_308,s_309;//RE__ALLOW(00,01,10,11);
input s_310,s_311;//RE__ALLOW(00,01,10,11);
input s_312,s_313;//RE__ALLOW(00,01,10,11);
input s_314,s_315;//RE__ALLOW(00,01,10,11);
input s_316,s_317;//RE__ALLOW(00,01,10,11);
input s_318,s_319;//RE__ALLOW(00,01,10,11);
input s_320,s_321;//RE__ALLOW(00,01,10,11);
input s_322,s_323;//RE__ALLOW(00,01,10,11);
input s_324,s_325;//RE__ALLOW(00,01,10,11);
input s_326,s_327;//RE__ALLOW(00,01,10,11);
input s_328,s_329;//RE__ALLOW(00,01,10,11);
input s_330,s_331;//RE__ALLOW(00,01,10,11);
input s_332,s_333;//RE__ALLOW(00,01,10,11);
input s_334,s_335;//RE__ALLOW(00,01,10,11);
input s_336,s_337;//RE__ALLOW(00,01,10,11);
input s_338,s_339;//RE__ALLOW(00,01,10,11);
input s_340,s_341;//RE__ALLOW(00,01,10,11);
input s_342,s_343;//RE__ALLOW(00,01,10,11);
input s_344,s_345;//RE__ALLOW(00,01,10,11);
input s_346,s_347;//RE__ALLOW(00,01,10,11);
input s_348,s_349;//RE__ALLOW(00,01,10,11);
input s_350,s_351;//RE__ALLOW(00,01,10,11);
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;

  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate392inter0, gate392inter1, gate392inter2, gate392inter3, gate392inter4, gate392inter5, gate392inter6, gate392inter7, gate392inter8, gate392inter9, gate392inter10, gate392inter11, gate392inter12, gate44inter0, gate44inter1, gate44inter2, gate44inter3, gate44inter4, gate44inter5, gate44inter6, gate44inter7, gate44inter8, gate44inter9, gate44inter10, gate44inter11, gate44inter12, gate225inter0, gate225inter1, gate225inter2, gate225inter3, gate225inter4, gate225inter5, gate225inter6, gate225inter7, gate225inter8, gate225inter9, gate225inter10, gate225inter11, gate225inter12, gate228inter0, gate228inter1, gate228inter2, gate228inter3, gate228inter4, gate228inter5, gate228inter6, gate228inter7, gate228inter8, gate228inter9, gate228inter10, gate228inter11, gate228inter12, gate117inter0, gate117inter1, gate117inter2, gate117inter3, gate117inter4, gate117inter5, gate117inter6, gate117inter7, gate117inter8, gate117inter9, gate117inter10, gate117inter11, gate117inter12, gate180inter0, gate180inter1, gate180inter2, gate180inter3, gate180inter4, gate180inter5, gate180inter6, gate180inter7, gate180inter8, gate180inter9, gate180inter10, gate180inter11, gate180inter12, gate236inter0, gate236inter1, gate236inter2, gate236inter3, gate236inter4, gate236inter5, gate236inter6, gate236inter7, gate236inter8, gate236inter9, gate236inter10, gate236inter11, gate236inter12, gate198inter0, gate198inter1, gate198inter2, gate198inter3, gate198inter4, gate198inter5, gate198inter6, gate198inter7, gate198inter8, gate198inter9, gate198inter10, gate198inter11, gate198inter12, gate101inter0, gate101inter1, gate101inter2, gate101inter3, gate101inter4, gate101inter5, gate101inter6, gate101inter7, gate101inter8, gate101inter9, gate101inter10, gate101inter11, gate101inter12, gate145inter0, gate145inter1, gate145inter2, gate145inter3, gate145inter4, gate145inter5, gate145inter6, gate145inter7, gate145inter8, gate145inter9, gate145inter10, gate145inter11, gate145inter12, gate291inter0, gate291inter1, gate291inter2, gate291inter3, gate291inter4, gate291inter5, gate291inter6, gate291inter7, gate291inter8, gate291inter9, gate291inter10, gate291inter11, gate291inter12, gate427inter0, gate427inter1, gate427inter2, gate427inter3, gate427inter4, gate427inter5, gate427inter6, gate427inter7, gate427inter8, gate427inter9, gate427inter10, gate427inter11, gate427inter12, gate221inter0, gate221inter1, gate221inter2, gate221inter3, gate221inter4, gate221inter5, gate221inter6, gate221inter7, gate221inter8, gate221inter9, gate221inter10, gate221inter11, gate221inter12, gate100inter0, gate100inter1, gate100inter2, gate100inter3, gate100inter4, gate100inter5, gate100inter6, gate100inter7, gate100inter8, gate100inter9, gate100inter10, gate100inter11, gate100inter12, gate25inter0, gate25inter1, gate25inter2, gate25inter3, gate25inter4, gate25inter5, gate25inter6, gate25inter7, gate25inter8, gate25inter9, gate25inter10, gate25inter11, gate25inter12, gate494inter0, gate494inter1, gate494inter2, gate494inter3, gate494inter4, gate494inter5, gate494inter6, gate494inter7, gate494inter8, gate494inter9, gate494inter10, gate494inter11, gate494inter12, gate63inter0, gate63inter1, gate63inter2, gate63inter3, gate63inter4, gate63inter5, gate63inter6, gate63inter7, gate63inter8, gate63inter9, gate63inter10, gate63inter11, gate63inter12, gate492inter0, gate492inter1, gate492inter2, gate492inter3, gate492inter4, gate492inter5, gate492inter6, gate492inter7, gate492inter8, gate492inter9, gate492inter10, gate492inter11, gate492inter12, gate474inter0, gate474inter1, gate474inter2, gate474inter3, gate474inter4, gate474inter5, gate474inter6, gate474inter7, gate474inter8, gate474inter9, gate474inter10, gate474inter11, gate474inter12, gate169inter0, gate169inter1, gate169inter2, gate169inter3, gate169inter4, gate169inter5, gate169inter6, gate169inter7, gate169inter8, gate169inter9, gate169inter10, gate169inter11, gate169inter12, gate399inter0, gate399inter1, gate399inter2, gate399inter3, gate399inter4, gate399inter5, gate399inter6, gate399inter7, gate399inter8, gate399inter9, gate399inter10, gate399inter11, gate399inter12, gate452inter0, gate452inter1, gate452inter2, gate452inter3, gate452inter4, gate452inter5, gate452inter6, gate452inter7, gate452inter8, gate452inter9, gate452inter10, gate452inter11, gate452inter12, gate128inter0, gate128inter1, gate128inter2, gate128inter3, gate128inter4, gate128inter5, gate128inter6, gate128inter7, gate128inter8, gate128inter9, gate128inter10, gate128inter11, gate128inter12, gate414inter0, gate414inter1, gate414inter2, gate414inter3, gate414inter4, gate414inter5, gate414inter6, gate414inter7, gate414inter8, gate414inter9, gate414inter10, gate414inter11, gate414inter12, gate49inter0, gate49inter1, gate49inter2, gate49inter3, gate49inter4, gate49inter5, gate49inter6, gate49inter7, gate49inter8, gate49inter9, gate49inter10, gate49inter11, gate49inter12, gate274inter0, gate274inter1, gate274inter2, gate274inter3, gate274inter4, gate274inter5, gate274inter6, gate274inter7, gate274inter8, gate274inter9, gate274inter10, gate274inter11, gate274inter12, gate58inter0, gate58inter1, gate58inter2, gate58inter3, gate58inter4, gate58inter5, gate58inter6, gate58inter7, gate58inter8, gate58inter9, gate58inter10, gate58inter11, gate58inter12, gate209inter0, gate209inter1, gate209inter2, gate209inter3, gate209inter4, gate209inter5, gate209inter6, gate209inter7, gate209inter8, gate209inter9, gate209inter10, gate209inter11, gate209inter12, gate95inter0, gate95inter1, gate95inter2, gate95inter3, gate95inter4, gate95inter5, gate95inter6, gate95inter7, gate95inter8, gate95inter9, gate95inter10, gate95inter11, gate95inter12, gate9inter0, gate9inter1, gate9inter2, gate9inter3, gate9inter4, gate9inter5, gate9inter6, gate9inter7, gate9inter8, gate9inter9, gate9inter10, gate9inter11, gate9inter12, gate290inter0, gate290inter1, gate290inter2, gate290inter3, gate290inter4, gate290inter5, gate290inter6, gate290inter7, gate290inter8, gate290inter9, gate290inter10, gate290inter11, gate290inter12, gate449inter0, gate449inter1, gate449inter2, gate449inter3, gate449inter4, gate449inter5, gate449inter6, gate449inter7, gate449inter8, gate449inter9, gate449inter10, gate449inter11, gate449inter12, gate233inter0, gate233inter1, gate233inter2, gate233inter3, gate233inter4, gate233inter5, gate233inter6, gate233inter7, gate233inter8, gate233inter9, gate233inter10, gate233inter11, gate233inter12, gate514inter0, gate514inter1, gate514inter2, gate514inter3, gate514inter4, gate514inter5, gate514inter6, gate514inter7, gate514inter8, gate514inter9, gate514inter10, gate514inter11, gate514inter12, gate388inter0, gate388inter1, gate388inter2, gate388inter3, gate388inter4, gate388inter5, gate388inter6, gate388inter7, gate388inter8, gate388inter9, gate388inter10, gate388inter11, gate388inter12, gate17inter0, gate17inter1, gate17inter2, gate17inter3, gate17inter4, gate17inter5, gate17inter6, gate17inter7, gate17inter8, gate17inter9, gate17inter10, gate17inter11, gate17inter12, gate458inter0, gate458inter1, gate458inter2, gate458inter3, gate458inter4, gate458inter5, gate458inter6, gate458inter7, gate458inter8, gate458inter9, gate458inter10, gate458inter11, gate458inter12, gate477inter0, gate477inter1, gate477inter2, gate477inter3, gate477inter4, gate477inter5, gate477inter6, gate477inter7, gate477inter8, gate477inter9, gate477inter10, gate477inter11, gate477inter12, gate207inter0, gate207inter1, gate207inter2, gate207inter3, gate207inter4, gate207inter5, gate207inter6, gate207inter7, gate207inter8, gate207inter9, gate207inter10, gate207inter11, gate207inter12, gate451inter0, gate451inter1, gate451inter2, gate451inter3, gate451inter4, gate451inter5, gate451inter6, gate451inter7, gate451inter8, gate451inter9, gate451inter10, gate451inter11, gate451inter12, gate475inter0, gate475inter1, gate475inter2, gate475inter3, gate475inter4, gate475inter5, gate475inter6, gate475inter7, gate475inter8, gate475inter9, gate475inter10, gate475inter11, gate475inter12, gate490inter0, gate490inter1, gate490inter2, gate490inter3, gate490inter4, gate490inter5, gate490inter6, gate490inter7, gate490inter8, gate490inter9, gate490inter10, gate490inter11, gate490inter12, gate420inter0, gate420inter1, gate420inter2, gate420inter3, gate420inter4, gate420inter5, gate420inter6, gate420inter7, gate420inter8, gate420inter9, gate420inter10, gate420inter11, gate420inter12, gate16inter0, gate16inter1, gate16inter2, gate16inter3, gate16inter4, gate16inter5, gate16inter6, gate16inter7, gate16inter8, gate16inter9, gate16inter10, gate16inter11, gate16inter12, gate442inter0, gate442inter1, gate442inter2, gate442inter3, gate442inter4, gate442inter5, gate442inter6, gate442inter7, gate442inter8, gate442inter9, gate442inter10, gate442inter11, gate442inter12, gate288inter0, gate288inter1, gate288inter2, gate288inter3, gate288inter4, gate288inter5, gate288inter6, gate288inter7, gate288inter8, gate288inter9, gate288inter10, gate288inter11, gate288inter12, gate467inter0, gate467inter1, gate467inter2, gate467inter3, gate467inter4, gate467inter5, gate467inter6, gate467inter7, gate467inter8, gate467inter9, gate467inter10, gate467inter11, gate467inter12, gate157inter0, gate157inter1, gate157inter2, gate157inter3, gate157inter4, gate157inter5, gate157inter6, gate157inter7, gate157inter8, gate157inter9, gate157inter10, gate157inter11, gate157inter12, gate126inter0, gate126inter1, gate126inter2, gate126inter3, gate126inter4, gate126inter5, gate126inter6, gate126inter7, gate126inter8, gate126inter9, gate126inter10, gate126inter11, gate126inter12, gate11inter0, gate11inter1, gate11inter2, gate11inter3, gate11inter4, gate11inter5, gate11inter6, gate11inter7, gate11inter8, gate11inter9, gate11inter10, gate11inter11, gate11inter12, gate202inter0, gate202inter1, gate202inter2, gate202inter3, gate202inter4, gate202inter5, gate202inter6, gate202inter7, gate202inter8, gate202inter9, gate202inter10, gate202inter11, gate202inter12, gate97inter0, gate97inter1, gate97inter2, gate97inter3, gate97inter4, gate97inter5, gate97inter6, gate97inter7, gate97inter8, gate97inter9, gate97inter10, gate97inter11, gate97inter12, gate77inter0, gate77inter1, gate77inter2, gate77inter3, gate77inter4, gate77inter5, gate77inter6, gate77inter7, gate77inter8, gate77inter9, gate77inter10, gate77inter11, gate77inter12, gate144inter0, gate144inter1, gate144inter2, gate144inter3, gate144inter4, gate144inter5, gate144inter6, gate144inter7, gate144inter8, gate144inter9, gate144inter10, gate144inter11, gate144inter12, gate224inter0, gate224inter1, gate224inter2, gate224inter3, gate224inter4, gate224inter5, gate224inter6, gate224inter7, gate224inter8, gate224inter9, gate224inter10, gate224inter11, gate224inter12, gate80inter0, gate80inter1, gate80inter2, gate80inter3, gate80inter4, gate80inter5, gate80inter6, gate80inter7, gate80inter8, gate80inter9, gate80inter10, gate80inter11, gate80inter12, gate113inter0, gate113inter1, gate113inter2, gate113inter3, gate113inter4, gate113inter5, gate113inter6, gate113inter7, gate113inter8, gate113inter9, gate113inter10, gate113inter11, gate113inter12, gate102inter0, gate102inter1, gate102inter2, gate102inter3, gate102inter4, gate102inter5, gate102inter6, gate102inter7, gate102inter8, gate102inter9, gate102inter10, gate102inter11, gate102inter12, gate255inter0, gate255inter1, gate255inter2, gate255inter3, gate255inter4, gate255inter5, gate255inter6, gate255inter7, gate255inter8, gate255inter9, gate255inter10, gate255inter11, gate255inter12, gate162inter0, gate162inter1, gate162inter2, gate162inter3, gate162inter4, gate162inter5, gate162inter6, gate162inter7, gate162inter8, gate162inter9, gate162inter10, gate162inter11, gate162inter12, gate407inter0, gate407inter1, gate407inter2, gate407inter3, gate407inter4, gate407inter5, gate407inter6, gate407inter7, gate407inter8, gate407inter9, gate407inter10, gate407inter11, gate407inter12, gate283inter0, gate283inter1, gate283inter2, gate283inter3, gate283inter4, gate283inter5, gate283inter6, gate283inter7, gate283inter8, gate283inter9, gate283inter10, gate283inter11, gate283inter12, gate253inter0, gate253inter1, gate253inter2, gate253inter3, gate253inter4, gate253inter5, gate253inter6, gate253inter7, gate253inter8, gate253inter9, gate253inter10, gate253inter11, gate253inter12, gate447inter0, gate447inter1, gate447inter2, gate447inter3, gate447inter4, gate447inter5, gate447inter6, gate447inter7, gate447inter8, gate447inter9, gate447inter10, gate447inter11, gate447inter12, gate455inter0, gate455inter1, gate455inter2, gate455inter3, gate455inter4, gate455inter5, gate455inter6, gate455inter7, gate455inter8, gate455inter9, gate455inter10, gate455inter11, gate455inter12, gate250inter0, gate250inter1, gate250inter2, gate250inter3, gate250inter4, gate250inter5, gate250inter6, gate250inter7, gate250inter8, gate250inter9, gate250inter10, gate250inter11, gate250inter12, gate120inter0, gate120inter1, gate120inter2, gate120inter3, gate120inter4, gate120inter5, gate120inter6, gate120inter7, gate120inter8, gate120inter9, gate120inter10, gate120inter11, gate120inter12, gate287inter0, gate287inter1, gate287inter2, gate287inter3, gate287inter4, gate287inter5, gate287inter6, gate287inter7, gate287inter8, gate287inter9, gate287inter10, gate287inter11, gate287inter12, gate421inter0, gate421inter1, gate421inter2, gate421inter3, gate421inter4, gate421inter5, gate421inter6, gate421inter7, gate421inter8, gate421inter9, gate421inter10, gate421inter11, gate421inter12, gate29inter0, gate29inter1, gate29inter2, gate29inter3, gate29inter4, gate29inter5, gate29inter6, gate29inter7, gate29inter8, gate29inter9, gate29inter10, gate29inter11, gate29inter12, gate460inter0, gate460inter1, gate460inter2, gate460inter3, gate460inter4, gate460inter5, gate460inter6, gate460inter7, gate460inter8, gate460inter9, gate460inter10, gate460inter11, gate460inter12, gate35inter0, gate35inter1, gate35inter2, gate35inter3, gate35inter4, gate35inter5, gate35inter6, gate35inter7, gate35inter8, gate35inter9, gate35inter10, gate35inter11, gate35inter12, gate395inter0, gate395inter1, gate395inter2, gate395inter3, gate395inter4, gate395inter5, gate395inter6, gate395inter7, gate395inter8, gate395inter9, gate395inter10, gate395inter11, gate395inter12, gate462inter0, gate462inter1, gate462inter2, gate462inter3, gate462inter4, gate462inter5, gate462inter6, gate462inter7, gate462inter8, gate462inter9, gate462inter10, gate462inter11, gate462inter12, gate406inter0, gate406inter1, gate406inter2, gate406inter3, gate406inter4, gate406inter5, gate406inter6, gate406inter7, gate406inter8, gate406inter9, gate406inter10, gate406inter11, gate406inter12, gate179inter0, gate179inter1, gate179inter2, gate179inter3, gate179inter4, gate179inter5, gate179inter6, gate179inter7, gate179inter8, gate179inter9, gate179inter10, gate179inter11, gate179inter12, gate178inter0, gate178inter1, gate178inter2, gate178inter3, gate178inter4, gate178inter5, gate178inter6, gate178inter7, gate178inter8, gate178inter9, gate178inter10, gate178inter11, gate178inter12, gate24inter0, gate24inter1, gate24inter2, gate24inter3, gate24inter4, gate24inter5, gate24inter6, gate24inter7, gate24inter8, gate24inter9, gate24inter10, gate24inter11, gate24inter12, gate497inter0, gate497inter1, gate497inter2, gate497inter3, gate497inter4, gate497inter5, gate497inter6, gate497inter7, gate497inter8, gate497inter9, gate497inter10, gate497inter11, gate497inter12, gate160inter0, gate160inter1, gate160inter2, gate160inter3, gate160inter4, gate160inter5, gate160inter6, gate160inter7, gate160inter8, gate160inter9, gate160inter10, gate160inter11, gate160inter12, gate513inter0, gate513inter1, gate513inter2, gate513inter3, gate513inter4, gate513inter5, gate513inter6, gate513inter7, gate513inter8, gate513inter9, gate513inter10, gate513inter11, gate513inter12, gate165inter0, gate165inter1, gate165inter2, gate165inter3, gate165inter4, gate165inter5, gate165inter6, gate165inter7, gate165inter8, gate165inter9, gate165inter10, gate165inter11, gate165inter12, gate143inter0, gate143inter1, gate143inter2, gate143inter3, gate143inter4, gate143inter5, gate143inter6, gate143inter7, gate143inter8, gate143inter9, gate143inter10, gate143inter11, gate143inter12, gate419inter0, gate419inter1, gate419inter2, gate419inter3, gate419inter4, gate419inter5, gate419inter6, gate419inter7, gate419inter8, gate419inter9, gate419inter10, gate419inter11, gate419inter12, gate230inter0, gate230inter1, gate230inter2, gate230inter3, gate230inter4, gate230inter5, gate230inter6, gate230inter7, gate230inter8, gate230inter9, gate230inter10, gate230inter11, gate230inter12, gate409inter0, gate409inter1, gate409inter2, gate409inter3, gate409inter4, gate409inter5, gate409inter6, gate409inter7, gate409inter8, gate409inter9, gate409inter10, gate409inter11, gate409inter12, gate166inter0, gate166inter1, gate166inter2, gate166inter3, gate166inter4, gate166inter5, gate166inter6, gate166inter7, gate166inter8, gate166inter9, gate166inter10, gate166inter11, gate166inter12, gate161inter0, gate161inter1, gate161inter2, gate161inter3, gate161inter4, gate161inter5, gate161inter6, gate161inter7, gate161inter8, gate161inter9, gate161inter10, gate161inter11, gate161inter12, gate507inter0, gate507inter1, gate507inter2, gate507inter3, gate507inter4, gate507inter5, gate507inter6, gate507inter7, gate507inter8, gate507inter9, gate507inter10, gate507inter11, gate507inter12, gate272inter0, gate272inter1, gate272inter2, gate272inter3, gate272inter4, gate272inter5, gate272inter6, gate272inter7, gate272inter8, gate272inter9, gate272inter10, gate272inter11, gate272inter12, gate26inter0, gate26inter1, gate26inter2, gate26inter3, gate26inter4, gate26inter5, gate26inter6, gate26inter7, gate26inter8, gate26inter9, gate26inter10, gate26inter11, gate26inter12, gate511inter0, gate511inter1, gate511inter2, gate511inter3, gate511inter4, gate511inter5, gate511inter6, gate511inter7, gate511inter8, gate511inter9, gate511inter10, gate511inter11, gate511inter12, gate67inter0, gate67inter1, gate67inter2, gate67inter3, gate67inter4, gate67inter5, gate67inter6, gate67inter7, gate67inter8, gate67inter9, gate67inter10, gate67inter11, gate67inter12, gate401inter0, gate401inter1, gate401inter2, gate401inter3, gate401inter4, gate401inter5, gate401inter6, gate401inter7, gate401inter8, gate401inter9, gate401inter10, gate401inter11, gate401inter12, gate448inter0, gate448inter1, gate448inter2, gate448inter3, gate448inter4, gate448inter5, gate448inter6, gate448inter7, gate448inter8, gate448inter9, gate448inter10, gate448inter11, gate448inter12, gate485inter0, gate485inter1, gate485inter2, gate485inter3, gate485inter4, gate485inter5, gate485inter6, gate485inter7, gate485inter8, gate485inter9, gate485inter10, gate485inter11, gate485inter12, gate33inter0, gate33inter1, gate33inter2, gate33inter3, gate33inter4, gate33inter5, gate33inter6, gate33inter7, gate33inter8, gate33inter9, gate33inter10, gate33inter11, gate33inter12, gate139inter0, gate139inter1, gate139inter2, gate139inter3, gate139inter4, gate139inter5, gate139inter6, gate139inter7, gate139inter8, gate139inter9, gate139inter10, gate139inter11, gate139inter12, gate53inter0, gate53inter1, gate53inter2, gate53inter3, gate53inter4, gate53inter5, gate53inter6, gate53inter7, gate53inter8, gate53inter9, gate53inter10, gate53inter11, gate53inter12, gate400inter0, gate400inter1, gate400inter2, gate400inter3, gate400inter4, gate400inter5, gate400inter6, gate400inter7, gate400inter8, gate400inter9, gate400inter10, gate400inter11, gate400inter12, gate47inter0, gate47inter1, gate47inter2, gate47inter3, gate47inter4, gate47inter5, gate47inter6, gate47inter7, gate47inter8, gate47inter9, gate47inter10, gate47inter11, gate47inter12, gate13inter0, gate13inter1, gate13inter2, gate13inter3, gate13inter4, gate13inter5, gate13inter6, gate13inter7, gate13inter8, gate13inter9, gate13inter10, gate13inter11, gate13inter12, gate436inter0, gate436inter1, gate436inter2, gate436inter3, gate436inter4, gate436inter5, gate436inter6, gate436inter7, gate436inter8, gate436inter9, gate436inter10, gate436inter11, gate436inter12, gate147inter0, gate147inter1, gate147inter2, gate147inter3, gate147inter4, gate147inter5, gate147inter6, gate147inter7, gate147inter8, gate147inter9, gate147inter10, gate147inter11, gate147inter12, gate503inter0, gate503inter1, gate503inter2, gate503inter3, gate503inter4, gate503inter5, gate503inter6, gate503inter7, gate503inter8, gate503inter9, gate503inter10, gate503inter11, gate503inter12, gate190inter0, gate190inter1, gate190inter2, gate190inter3, gate190inter4, gate190inter5, gate190inter6, gate190inter7, gate190inter8, gate190inter9, gate190inter10, gate190inter11, gate190inter12, gate261inter0, gate261inter1, gate261inter2, gate261inter3, gate261inter4, gate261inter5, gate261inter6, gate261inter7, gate261inter8, gate261inter9, gate261inter10, gate261inter11, gate261inter12, gate239inter0, gate239inter1, gate239inter2, gate239inter3, gate239inter4, gate239inter5, gate239inter6, gate239inter7, gate239inter8, gate239inter9, gate239inter10, gate239inter11, gate239inter12, gate232inter0, gate232inter1, gate232inter2, gate232inter3, gate232inter4, gate232inter5, gate232inter6, gate232inter7, gate232inter8, gate232inter9, gate232inter10, gate232inter11, gate232inter12, gate72inter0, gate72inter1, gate72inter2, gate72inter3, gate72inter4, gate72inter5, gate72inter6, gate72inter7, gate72inter8, gate72inter9, gate72inter10, gate72inter11, gate72inter12, gate499inter0, gate499inter1, gate499inter2, gate499inter3, gate499inter4, gate499inter5, gate499inter6, gate499inter7, gate499inter8, gate499inter9, gate499inter10, gate499inter11, gate499inter12, gate217inter0, gate217inter1, gate217inter2, gate217inter3, gate217inter4, gate217inter5, gate217inter6, gate217inter7, gate217inter8, gate217inter9, gate217inter10, gate217inter11, gate217inter12, gate294inter0, gate294inter1, gate294inter2, gate294inter3, gate294inter4, gate294inter5, gate294inter6, gate294inter7, gate294inter8, gate294inter9, gate294inter10, gate294inter11, gate294inter12, gate210inter0, gate210inter1, gate210inter2, gate210inter3, gate210inter4, gate210inter5, gate210inter6, gate210inter7, gate210inter8, gate210inter9, gate210inter10, gate210inter11, gate210inter12, gate238inter0, gate238inter1, gate238inter2, gate238inter3, gate238inter4, gate238inter5, gate238inter6, gate238inter7, gate238inter8, gate238inter9, gate238inter10, gate238inter11, gate238inter12, gate276inter0, gate276inter1, gate276inter2, gate276inter3, gate276inter4, gate276inter5, gate276inter6, gate276inter7, gate276inter8, gate276inter9, gate276inter10, gate276inter11, gate276inter12, gate416inter0, gate416inter1, gate416inter2, gate416inter3, gate416inter4, gate416inter5, gate416inter6, gate416inter7, gate416inter8, gate416inter9, gate416inter10, gate416inter11, gate416inter12, gate295inter0, gate295inter1, gate295inter2, gate295inter3, gate295inter4, gate295inter5, gate295inter6, gate295inter7, gate295inter8, gate295inter9, gate295inter10, gate295inter11, gate295inter12, gate42inter0, gate42inter1, gate42inter2, gate42inter3, gate42inter4, gate42inter5, gate42inter6, gate42inter7, gate42inter8, gate42inter9, gate42inter10, gate42inter11, gate42inter12, gate123inter0, gate123inter1, gate123inter2, gate123inter3, gate123inter4, gate123inter5, gate123inter6, gate123inter7, gate123inter8, gate123inter9, gate123inter10, gate123inter11, gate123inter12, gate435inter0, gate435inter1, gate435inter2, gate435inter3, gate435inter4, gate435inter5, gate435inter6, gate435inter7, gate435inter8, gate435inter9, gate435inter10, gate435inter11, gate435inter12, gate170inter0, gate170inter1, gate170inter2, gate170inter3, gate170inter4, gate170inter5, gate170inter6, gate170inter7, gate170inter8, gate170inter9, gate170inter10, gate170inter11, gate170inter12, gate439inter0, gate439inter1, gate439inter2, gate439inter3, gate439inter4, gate439inter5, gate439inter6, gate439inter7, gate439inter8, gate439inter9, gate439inter10, gate439inter11, gate439inter12, gate398inter0, gate398inter1, gate398inter2, gate398inter3, gate398inter4, gate398inter5, gate398inter6, gate398inter7, gate398inter8, gate398inter9, gate398inter10, gate398inter11, gate398inter12, gate243inter0, gate243inter1, gate243inter2, gate243inter3, gate243inter4, gate243inter5, gate243inter6, gate243inter7, gate243inter8, gate243inter9, gate243inter10, gate243inter11, gate243inter12, gate446inter0, gate446inter1, gate446inter2, gate446inter3, gate446inter4, gate446inter5, gate446inter6, gate446inter7, gate446inter8, gate446inter9, gate446inter10, gate446inter11, gate446inter12, gate408inter0, gate408inter1, gate408inter2, gate408inter3, gate408inter4, gate408inter5, gate408inter6, gate408inter7, gate408inter8, gate408inter9, gate408inter10, gate408inter11, gate408inter12, gate175inter0, gate175inter1, gate175inter2, gate175inter3, gate175inter4, gate175inter5, gate175inter6, gate175inter7, gate175inter8, gate175inter9, gate175inter10, gate175inter11, gate175inter12, gate171inter0, gate171inter1, gate171inter2, gate171inter3, gate171inter4, gate171inter5, gate171inter6, gate171inter7, gate171inter8, gate171inter9, gate171inter10, gate171inter11, gate171inter12, gate48inter0, gate48inter1, gate48inter2, gate48inter3, gate48inter4, gate48inter5, gate48inter6, gate48inter7, gate48inter8, gate48inter9, gate48inter10, gate48inter11, gate48inter12, gate88inter0, gate88inter1, gate88inter2, gate88inter3, gate88inter4, gate88inter5, gate88inter6, gate88inter7, gate88inter8, gate88inter9, gate88inter10, gate88inter11, gate88inter12, gate19inter0, gate19inter1, gate19inter2, gate19inter3, gate19inter4, gate19inter5, gate19inter6, gate19inter7, gate19inter8, gate19inter9, gate19inter10, gate19inter11, gate19inter12, gate129inter0, gate129inter1, gate129inter2, gate129inter3, gate129inter4, gate129inter5, gate129inter6, gate129inter7, gate129inter8, gate129inter9, gate129inter10, gate129inter11, gate129inter12, gate218inter0, gate218inter1, gate218inter2, gate218inter3, gate218inter4, gate218inter5, gate218inter6, gate218inter7, gate218inter8, gate218inter9, gate218inter10, gate218inter11, gate218inter12, gate111inter0, gate111inter1, gate111inter2, gate111inter3, gate111inter4, gate111inter5, gate111inter6, gate111inter7, gate111inter8, gate111inter9, gate111inter10, gate111inter11, gate111inter12, gate12inter0, gate12inter1, gate12inter2, gate12inter3, gate12inter4, gate12inter5, gate12inter6, gate12inter7, gate12inter8, gate12inter9, gate12inter10, gate12inter11, gate12inter12, gate193inter0, gate193inter1, gate193inter2, gate193inter3, gate193inter4, gate193inter5, gate193inter6, gate193inter7, gate193inter8, gate193inter9, gate193inter10, gate193inter11, gate193inter12, gate251inter0, gate251inter1, gate251inter2, gate251inter3, gate251inter4, gate251inter5, gate251inter6, gate251inter7, gate251inter8, gate251inter9, gate251inter10, gate251inter11, gate251inter12, gate264inter0, gate264inter1, gate264inter2, gate264inter3, gate264inter4, gate264inter5, gate264inter6, gate264inter7, gate264inter8, gate264inter9, gate264inter10, gate264inter11, gate264inter12, gate212inter0, gate212inter1, gate212inter2, gate212inter3, gate212inter4, gate212inter5, gate212inter6, gate212inter7, gate212inter8, gate212inter9, gate212inter10, gate212inter11, gate212inter12, gate159inter0, gate159inter1, gate159inter2, gate159inter3, gate159inter4, gate159inter5, gate159inter6, gate159inter7, gate159inter8, gate159inter9, gate159inter10, gate159inter11, gate159inter12, gate277inter0, gate277inter1, gate277inter2, gate277inter3, gate277inter4, gate277inter5, gate277inter6, gate277inter7, gate277inter8, gate277inter9, gate277inter10, gate277inter11, gate277inter12, gate205inter0, gate205inter1, gate205inter2, gate205inter3, gate205inter4, gate205inter5, gate205inter6, gate205inter7, gate205inter8, gate205inter9, gate205inter10, gate205inter11, gate205inter12, gate254inter0, gate254inter1, gate254inter2, gate254inter3, gate254inter4, gate254inter5, gate254inter6, gate254inter7, gate254inter8, gate254inter9, gate254inter10, gate254inter11, gate254inter12, gate32inter0, gate32inter1, gate32inter2, gate32inter3, gate32inter4, gate32inter5, gate32inter6, gate32inter7, gate32inter8, gate32inter9, gate32inter10, gate32inter11, gate32inter12, gate52inter0, gate52inter1, gate52inter2, gate52inter3, gate52inter4, gate52inter5, gate52inter6, gate52inter7, gate52inter8, gate52inter9, gate52inter10, gate52inter11, gate52inter12, gate71inter0, gate71inter1, gate71inter2, gate71inter3, gate71inter4, gate71inter5, gate71inter6, gate71inter7, gate71inter8, gate71inter9, gate71inter10, gate71inter11, gate71inter12, gate131inter0, gate131inter1, gate131inter2, gate131inter3, gate131inter4, gate131inter5, gate131inter6, gate131inter7, gate131inter8, gate131inter9, gate131inter10, gate131inter11, gate131inter12, gate456inter0, gate456inter1, gate456inter2, gate456inter3, gate456inter4, gate456inter5, gate456inter6, gate456inter7, gate456inter8, gate456inter9, gate456inter10, gate456inter11, gate456inter12, gate98inter0, gate98inter1, gate98inter2, gate98inter3, gate98inter4, gate98inter5, gate98inter6, gate98inter7, gate98inter8, gate98inter9, gate98inter10, gate98inter11, gate98inter12, gate121inter0, gate121inter1, gate121inter2, gate121inter3, gate121inter4, gate121inter5, gate121inter6, gate121inter7, gate121inter8, gate121inter9, gate121inter10, gate121inter11, gate121inter12, gate176inter0, gate176inter1, gate176inter2, gate176inter3, gate176inter4, gate176inter5, gate176inter6, gate176inter7, gate176inter8, gate176inter9, gate176inter10, gate176inter11, gate176inter12, gate437inter0, gate437inter1, gate437inter2, gate437inter3, gate437inter4, gate437inter5, gate437inter6, gate437inter7, gate437inter8, gate437inter9, gate437inter10, gate437inter11, gate437inter12, gate20inter0, gate20inter1, gate20inter2, gate20inter3, gate20inter4, gate20inter5, gate20inter6, gate20inter7, gate20inter8, gate20inter9, gate20inter10, gate20inter11, gate20inter12, gate216inter0, gate216inter1, gate216inter2, gate216inter3, gate216inter4, gate216inter5, gate216inter6, gate216inter7, gate216inter8, gate216inter9, gate216inter10, gate216inter11, gate216inter12, gate262inter0, gate262inter1, gate262inter2, gate262inter3, gate262inter4, gate262inter5, gate262inter6, gate262inter7, gate262inter8, gate262inter9, gate262inter10, gate262inter11, gate262inter12, gate135inter0, gate135inter1, gate135inter2, gate135inter3, gate135inter4, gate135inter5, gate135inter6, gate135inter7, gate135inter8, gate135inter9, gate135inter10, gate135inter11, gate135inter12, gate508inter0, gate508inter1, gate508inter2, gate508inter3, gate508inter4, gate508inter5, gate508inter6, gate508inter7, gate508inter8, gate508inter9, gate508inter10, gate508inter11, gate508inter12, gate22inter0, gate22inter1, gate22inter2, gate22inter3, gate22inter4, gate22inter5, gate22inter6, gate22inter7, gate22inter8, gate22inter9, gate22inter10, gate22inter11, gate22inter12, gate85inter0, gate85inter1, gate85inter2, gate85inter3, gate85inter4, gate85inter5, gate85inter6, gate85inter7, gate85inter8, gate85inter9, gate85inter10, gate85inter11, gate85inter12, gate222inter0, gate222inter1, gate222inter2, gate222inter3, gate222inter4, gate222inter5, gate222inter6, gate222inter7, gate222inter8, gate222inter9, gate222inter10, gate222inter11, gate222inter12, gate496inter0, gate496inter1, gate496inter2, gate496inter3, gate496inter4, gate496inter5, gate496inter6, gate496inter7, gate496inter8, gate496inter9, gate496inter10, gate496inter11, gate496inter12, gate116inter0, gate116inter1, gate116inter2, gate116inter3, gate116inter4, gate116inter5, gate116inter6, gate116inter7, gate116inter8, gate116inter9, gate116inter10, gate116inter11, gate116inter12, gate219inter0, gate219inter1, gate219inter2, gate219inter3, gate219inter4, gate219inter5, gate219inter6, gate219inter7, gate219inter8, gate219inter9, gate219inter10, gate219inter11, gate219inter12, gate15inter0, gate15inter1, gate15inter2, gate15inter3, gate15inter4, gate15inter5, gate15inter6, gate15inter7, gate15inter8, gate15inter9, gate15inter10, gate15inter11, gate15inter12, gate201inter0, gate201inter1, gate201inter2, gate201inter3, gate201inter4, gate201inter5, gate201inter6, gate201inter7, gate201inter8, gate201inter9, gate201inter10, gate201inter11, gate201inter12, gate61inter0, gate61inter1, gate61inter2, gate61inter3, gate61inter4, gate61inter5, gate61inter6, gate61inter7, gate61inter8, gate61inter9, gate61inter10, gate61inter11, gate61inter12, gate174inter0, gate174inter1, gate174inter2, gate174inter3, gate174inter4, gate174inter5, gate174inter6, gate174inter7, gate174inter8, gate174inter9, gate174inter10, gate174inter11, gate174inter12, gate43inter0, gate43inter1, gate43inter2, gate43inter3, gate43inter4, gate43inter5, gate43inter6, gate43inter7, gate43inter8, gate43inter9, gate43inter10, gate43inter11, gate43inter12, gate96inter0, gate96inter1, gate96inter2, gate96inter3, gate96inter4, gate96inter5, gate96inter6, gate96inter7, gate96inter8, gate96inter9, gate96inter10, gate96inter11, gate96inter12, gate267inter0, gate267inter1, gate267inter2, gate267inter3, gate267inter4, gate267inter5, gate267inter6, gate267inter7, gate267inter8, gate267inter9, gate267inter10, gate267inter11, gate267inter12, gate142inter0, gate142inter1, gate142inter2, gate142inter3, gate142inter4, gate142inter5, gate142inter6, gate142inter7, gate142inter8, gate142inter9, gate142inter10, gate142inter11, gate142inter12, gate124inter0, gate124inter1, gate124inter2, gate124inter3, gate124inter4, gate124inter5, gate124inter6, gate124inter7, gate124inter8, gate124inter9, gate124inter10, gate124inter11, gate124inter12, gate185inter0, gate185inter1, gate185inter2, gate185inter3, gate185inter4, gate185inter5, gate185inter6, gate185inter7, gate185inter8, gate185inter9, gate185inter10, gate185inter11, gate185inter12, gate82inter0, gate82inter1, gate82inter2, gate82inter3, gate82inter4, gate82inter5, gate82inter6, gate82inter7, gate82inter8, gate82inter9, gate82inter10, gate82inter11, gate82inter12, gate119inter0, gate119inter1, gate119inter2, gate119inter3, gate119inter4, gate119inter5, gate119inter6, gate119inter7, gate119inter8, gate119inter9, gate119inter10, gate119inter11, gate119inter12;



and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );

  xor2  gate953(.a(G2), .b(G1), .O(gate9inter0));
  nand2 gate954(.a(gate9inter0), .b(s_58), .O(gate9inter1));
  and2  gate955(.a(G2), .b(G1), .O(gate9inter2));
  inv1  gate956(.a(s_58), .O(gate9inter3));
  inv1  gate957(.a(s_59), .O(gate9inter4));
  nand2 gate958(.a(gate9inter4), .b(gate9inter3), .O(gate9inter5));
  nor2  gate959(.a(gate9inter5), .b(gate9inter2), .O(gate9inter6));
  inv1  gate960(.a(G1), .O(gate9inter7));
  inv1  gate961(.a(G2), .O(gate9inter8));
  nand2 gate962(.a(gate9inter8), .b(gate9inter7), .O(gate9inter9));
  nand2 gate963(.a(s_59), .b(gate9inter3), .O(gate9inter10));
  nor2  gate964(.a(gate9inter10), .b(gate9inter9), .O(gate9inter11));
  nor2  gate965(.a(gate9inter11), .b(gate9inter6), .O(gate9inter12));
  nand2 gate966(.a(gate9inter12), .b(gate9inter1), .O(G266));
nand2 gate10( .a(G3), .b(G4), .O(G269) );

  xor2  gate1233(.a(G6), .b(G5), .O(gate11inter0));
  nand2 gate1234(.a(gate11inter0), .b(s_98), .O(gate11inter1));
  and2  gate1235(.a(G6), .b(G5), .O(gate11inter2));
  inv1  gate1236(.a(s_98), .O(gate11inter3));
  inv1  gate1237(.a(s_99), .O(gate11inter4));
  nand2 gate1238(.a(gate11inter4), .b(gate11inter3), .O(gate11inter5));
  nor2  gate1239(.a(gate11inter5), .b(gate11inter2), .O(gate11inter6));
  inv1  gate1240(.a(G5), .O(gate11inter7));
  inv1  gate1241(.a(G6), .O(gate11inter8));
  nand2 gate1242(.a(gate11inter8), .b(gate11inter7), .O(gate11inter9));
  nand2 gate1243(.a(s_99), .b(gate11inter3), .O(gate11inter10));
  nor2  gate1244(.a(gate11inter10), .b(gate11inter9), .O(gate11inter11));
  nor2  gate1245(.a(gate11inter11), .b(gate11inter6), .O(gate11inter12));
  nand2 gate1246(.a(gate11inter12), .b(gate11inter1), .O(G272));

  xor2  gate2437(.a(G8), .b(G7), .O(gate12inter0));
  nand2 gate2438(.a(gate12inter0), .b(s_270), .O(gate12inter1));
  and2  gate2439(.a(G8), .b(G7), .O(gate12inter2));
  inv1  gate2440(.a(s_270), .O(gate12inter3));
  inv1  gate2441(.a(s_271), .O(gate12inter4));
  nand2 gate2442(.a(gate12inter4), .b(gate12inter3), .O(gate12inter5));
  nor2  gate2443(.a(gate12inter5), .b(gate12inter2), .O(gate12inter6));
  inv1  gate2444(.a(G7), .O(gate12inter7));
  inv1  gate2445(.a(G8), .O(gate12inter8));
  nand2 gate2446(.a(gate12inter8), .b(gate12inter7), .O(gate12inter9));
  nand2 gate2447(.a(s_271), .b(gate12inter3), .O(gate12inter10));
  nor2  gate2448(.a(gate12inter10), .b(gate12inter9), .O(gate12inter11));
  nor2  gate2449(.a(gate12inter11), .b(gate12inter6), .O(gate12inter12));
  nand2 gate2450(.a(gate12inter12), .b(gate12inter1), .O(G275));

  xor2  gate1961(.a(G10), .b(G9), .O(gate13inter0));
  nand2 gate1962(.a(gate13inter0), .b(s_202), .O(gate13inter1));
  and2  gate1963(.a(G10), .b(G9), .O(gate13inter2));
  inv1  gate1964(.a(s_202), .O(gate13inter3));
  inv1  gate1965(.a(s_203), .O(gate13inter4));
  nand2 gate1966(.a(gate13inter4), .b(gate13inter3), .O(gate13inter5));
  nor2  gate1967(.a(gate13inter5), .b(gate13inter2), .O(gate13inter6));
  inv1  gate1968(.a(G9), .O(gate13inter7));
  inv1  gate1969(.a(G10), .O(gate13inter8));
  nand2 gate1970(.a(gate13inter8), .b(gate13inter7), .O(gate13inter9));
  nand2 gate1971(.a(s_203), .b(gate13inter3), .O(gate13inter10));
  nor2  gate1972(.a(gate13inter10), .b(gate13inter9), .O(gate13inter11));
  nor2  gate1973(.a(gate13inter11), .b(gate13inter6), .O(gate13inter12));
  nand2 gate1974(.a(gate13inter12), .b(gate13inter1), .O(G278));
nand2 gate14( .a(G11), .b(G12), .O(G281) );

  xor2  gate2843(.a(G14), .b(G13), .O(gate15inter0));
  nand2 gate2844(.a(gate15inter0), .b(s_328), .O(gate15inter1));
  and2  gate2845(.a(G14), .b(G13), .O(gate15inter2));
  inv1  gate2846(.a(s_328), .O(gate15inter3));
  inv1  gate2847(.a(s_329), .O(gate15inter4));
  nand2 gate2848(.a(gate15inter4), .b(gate15inter3), .O(gate15inter5));
  nor2  gate2849(.a(gate15inter5), .b(gate15inter2), .O(gate15inter6));
  inv1  gate2850(.a(G13), .O(gate15inter7));
  inv1  gate2851(.a(G14), .O(gate15inter8));
  nand2 gate2852(.a(gate15inter8), .b(gate15inter7), .O(gate15inter9));
  nand2 gate2853(.a(s_329), .b(gate15inter3), .O(gate15inter10));
  nor2  gate2854(.a(gate15inter10), .b(gate15inter9), .O(gate15inter11));
  nor2  gate2855(.a(gate15inter11), .b(gate15inter6), .O(gate15inter12));
  nand2 gate2856(.a(gate15inter12), .b(gate15inter1), .O(G284));

  xor2  gate1149(.a(G16), .b(G15), .O(gate16inter0));
  nand2 gate1150(.a(gate16inter0), .b(s_86), .O(gate16inter1));
  and2  gate1151(.a(G16), .b(G15), .O(gate16inter2));
  inv1  gate1152(.a(s_86), .O(gate16inter3));
  inv1  gate1153(.a(s_87), .O(gate16inter4));
  nand2 gate1154(.a(gate16inter4), .b(gate16inter3), .O(gate16inter5));
  nor2  gate1155(.a(gate16inter5), .b(gate16inter2), .O(gate16inter6));
  inv1  gate1156(.a(G15), .O(gate16inter7));
  inv1  gate1157(.a(G16), .O(gate16inter8));
  nand2 gate1158(.a(gate16inter8), .b(gate16inter7), .O(gate16inter9));
  nand2 gate1159(.a(s_87), .b(gate16inter3), .O(gate16inter10));
  nor2  gate1160(.a(gate16inter10), .b(gate16inter9), .O(gate16inter11));
  nor2  gate1161(.a(gate16inter11), .b(gate16inter6), .O(gate16inter12));
  nand2 gate1162(.a(gate16inter12), .b(gate16inter1), .O(G287));

  xor2  gate1037(.a(G18), .b(G17), .O(gate17inter0));
  nand2 gate1038(.a(gate17inter0), .b(s_70), .O(gate17inter1));
  and2  gate1039(.a(G18), .b(G17), .O(gate17inter2));
  inv1  gate1040(.a(s_70), .O(gate17inter3));
  inv1  gate1041(.a(s_71), .O(gate17inter4));
  nand2 gate1042(.a(gate17inter4), .b(gate17inter3), .O(gate17inter5));
  nor2  gate1043(.a(gate17inter5), .b(gate17inter2), .O(gate17inter6));
  inv1  gate1044(.a(G17), .O(gate17inter7));
  inv1  gate1045(.a(G18), .O(gate17inter8));
  nand2 gate1046(.a(gate17inter8), .b(gate17inter7), .O(gate17inter9));
  nand2 gate1047(.a(s_71), .b(gate17inter3), .O(gate17inter10));
  nor2  gate1048(.a(gate17inter10), .b(gate17inter9), .O(gate17inter11));
  nor2  gate1049(.a(gate17inter11), .b(gate17inter6), .O(gate17inter12));
  nand2 gate1050(.a(gate17inter12), .b(gate17inter1), .O(G290));
nand2 gate18( .a(G19), .b(G20), .O(G293) );

  xor2  gate2381(.a(G22), .b(G21), .O(gate19inter0));
  nand2 gate2382(.a(gate19inter0), .b(s_262), .O(gate19inter1));
  and2  gate2383(.a(G22), .b(G21), .O(gate19inter2));
  inv1  gate2384(.a(s_262), .O(gate19inter3));
  inv1  gate2385(.a(s_263), .O(gate19inter4));
  nand2 gate2386(.a(gate19inter4), .b(gate19inter3), .O(gate19inter5));
  nor2  gate2387(.a(gate19inter5), .b(gate19inter2), .O(gate19inter6));
  inv1  gate2388(.a(G21), .O(gate19inter7));
  inv1  gate2389(.a(G22), .O(gate19inter8));
  nand2 gate2390(.a(gate19inter8), .b(gate19inter7), .O(gate19inter9));
  nand2 gate2391(.a(s_263), .b(gate19inter3), .O(gate19inter10));
  nor2  gate2392(.a(gate19inter10), .b(gate19inter9), .O(gate19inter11));
  nor2  gate2393(.a(gate19inter11), .b(gate19inter6), .O(gate19inter12));
  nand2 gate2394(.a(gate19inter12), .b(gate19inter1), .O(G296));

  xor2  gate2689(.a(G24), .b(G23), .O(gate20inter0));
  nand2 gate2690(.a(gate20inter0), .b(s_306), .O(gate20inter1));
  and2  gate2691(.a(G24), .b(G23), .O(gate20inter2));
  inv1  gate2692(.a(s_306), .O(gate20inter3));
  inv1  gate2693(.a(s_307), .O(gate20inter4));
  nand2 gate2694(.a(gate20inter4), .b(gate20inter3), .O(gate20inter5));
  nor2  gate2695(.a(gate20inter5), .b(gate20inter2), .O(gate20inter6));
  inv1  gate2696(.a(G23), .O(gate20inter7));
  inv1  gate2697(.a(G24), .O(gate20inter8));
  nand2 gate2698(.a(gate20inter8), .b(gate20inter7), .O(gate20inter9));
  nand2 gate2699(.a(s_307), .b(gate20inter3), .O(gate20inter10));
  nor2  gate2700(.a(gate20inter10), .b(gate20inter9), .O(gate20inter11));
  nor2  gate2701(.a(gate20inter11), .b(gate20inter6), .O(gate20inter12));
  nand2 gate2702(.a(gate20inter12), .b(gate20inter1), .O(G299));
nand2 gate21( .a(G25), .b(G26), .O(G302) );

  xor2  gate2759(.a(G28), .b(G27), .O(gate22inter0));
  nand2 gate2760(.a(gate22inter0), .b(s_316), .O(gate22inter1));
  and2  gate2761(.a(G28), .b(G27), .O(gate22inter2));
  inv1  gate2762(.a(s_316), .O(gate22inter3));
  inv1  gate2763(.a(s_317), .O(gate22inter4));
  nand2 gate2764(.a(gate22inter4), .b(gate22inter3), .O(gate22inter5));
  nor2  gate2765(.a(gate22inter5), .b(gate22inter2), .O(gate22inter6));
  inv1  gate2766(.a(G27), .O(gate22inter7));
  inv1  gate2767(.a(G28), .O(gate22inter8));
  nand2 gate2768(.a(gate22inter8), .b(gate22inter7), .O(gate22inter9));
  nand2 gate2769(.a(s_317), .b(gate22inter3), .O(gate22inter10));
  nor2  gate2770(.a(gate22inter10), .b(gate22inter9), .O(gate22inter11));
  nor2  gate2771(.a(gate22inter11), .b(gate22inter6), .O(gate22inter12));
  nand2 gate2772(.a(gate22inter12), .b(gate22inter1), .O(G305));
nand2 gate23( .a(G29), .b(G30), .O(G308) );

  xor2  gate1625(.a(G32), .b(G31), .O(gate24inter0));
  nand2 gate1626(.a(gate24inter0), .b(s_154), .O(gate24inter1));
  and2  gate1627(.a(G32), .b(G31), .O(gate24inter2));
  inv1  gate1628(.a(s_154), .O(gate24inter3));
  inv1  gate1629(.a(s_155), .O(gate24inter4));
  nand2 gate1630(.a(gate24inter4), .b(gate24inter3), .O(gate24inter5));
  nor2  gate1631(.a(gate24inter5), .b(gate24inter2), .O(gate24inter6));
  inv1  gate1632(.a(G31), .O(gate24inter7));
  inv1  gate1633(.a(G32), .O(gate24inter8));
  nand2 gate1634(.a(gate24inter8), .b(gate24inter7), .O(gate24inter9));
  nand2 gate1635(.a(s_155), .b(gate24inter3), .O(gate24inter10));
  nor2  gate1636(.a(gate24inter10), .b(gate24inter9), .O(gate24inter11));
  nor2  gate1637(.a(gate24inter11), .b(gate24inter6), .O(gate24inter12));
  nand2 gate1638(.a(gate24inter12), .b(gate24inter1), .O(G311));

  xor2  gate743(.a(G5), .b(G1), .O(gate25inter0));
  nand2 gate744(.a(gate25inter0), .b(s_28), .O(gate25inter1));
  and2  gate745(.a(G5), .b(G1), .O(gate25inter2));
  inv1  gate746(.a(s_28), .O(gate25inter3));
  inv1  gate747(.a(s_29), .O(gate25inter4));
  nand2 gate748(.a(gate25inter4), .b(gate25inter3), .O(gate25inter5));
  nor2  gate749(.a(gate25inter5), .b(gate25inter2), .O(gate25inter6));
  inv1  gate750(.a(G1), .O(gate25inter7));
  inv1  gate751(.a(G5), .O(gate25inter8));
  nand2 gate752(.a(gate25inter8), .b(gate25inter7), .O(gate25inter9));
  nand2 gate753(.a(s_29), .b(gate25inter3), .O(gate25inter10));
  nor2  gate754(.a(gate25inter10), .b(gate25inter9), .O(gate25inter11));
  nor2  gate755(.a(gate25inter11), .b(gate25inter6), .O(gate25inter12));
  nand2 gate756(.a(gate25inter12), .b(gate25inter1), .O(G314));

  xor2  gate1807(.a(G13), .b(G9), .O(gate26inter0));
  nand2 gate1808(.a(gate26inter0), .b(s_180), .O(gate26inter1));
  and2  gate1809(.a(G13), .b(G9), .O(gate26inter2));
  inv1  gate1810(.a(s_180), .O(gate26inter3));
  inv1  gate1811(.a(s_181), .O(gate26inter4));
  nand2 gate1812(.a(gate26inter4), .b(gate26inter3), .O(gate26inter5));
  nor2  gate1813(.a(gate26inter5), .b(gate26inter2), .O(gate26inter6));
  inv1  gate1814(.a(G9), .O(gate26inter7));
  inv1  gate1815(.a(G13), .O(gate26inter8));
  nand2 gate1816(.a(gate26inter8), .b(gate26inter7), .O(gate26inter9));
  nand2 gate1817(.a(s_181), .b(gate26inter3), .O(gate26inter10));
  nor2  gate1818(.a(gate26inter10), .b(gate26inter9), .O(gate26inter11));
  nor2  gate1819(.a(gate26inter11), .b(gate26inter6), .O(gate26inter12));
  nand2 gate1820(.a(gate26inter12), .b(gate26inter1), .O(G317));
nand2 gate27( .a(G2), .b(G6), .O(G320) );
nand2 gate28( .a(G10), .b(G14), .O(G323) );

  xor2  gate1513(.a(G7), .b(G3), .O(gate29inter0));
  nand2 gate1514(.a(gate29inter0), .b(s_138), .O(gate29inter1));
  and2  gate1515(.a(G7), .b(G3), .O(gate29inter2));
  inv1  gate1516(.a(s_138), .O(gate29inter3));
  inv1  gate1517(.a(s_139), .O(gate29inter4));
  nand2 gate1518(.a(gate29inter4), .b(gate29inter3), .O(gate29inter5));
  nor2  gate1519(.a(gate29inter5), .b(gate29inter2), .O(gate29inter6));
  inv1  gate1520(.a(G3), .O(gate29inter7));
  inv1  gate1521(.a(G7), .O(gate29inter8));
  nand2 gate1522(.a(gate29inter8), .b(gate29inter7), .O(gate29inter9));
  nand2 gate1523(.a(s_139), .b(gate29inter3), .O(gate29inter10));
  nor2  gate1524(.a(gate29inter10), .b(gate29inter9), .O(gate29inter11));
  nor2  gate1525(.a(gate29inter11), .b(gate29inter6), .O(gate29inter12));
  nand2 gate1526(.a(gate29inter12), .b(gate29inter1), .O(G326));
nand2 gate30( .a(G11), .b(G15), .O(G329) );
nand2 gate31( .a(G4), .b(G8), .O(G332) );

  xor2  gate2563(.a(G16), .b(G12), .O(gate32inter0));
  nand2 gate2564(.a(gate32inter0), .b(s_288), .O(gate32inter1));
  and2  gate2565(.a(G16), .b(G12), .O(gate32inter2));
  inv1  gate2566(.a(s_288), .O(gate32inter3));
  inv1  gate2567(.a(s_289), .O(gate32inter4));
  nand2 gate2568(.a(gate32inter4), .b(gate32inter3), .O(gate32inter5));
  nor2  gate2569(.a(gate32inter5), .b(gate32inter2), .O(gate32inter6));
  inv1  gate2570(.a(G12), .O(gate32inter7));
  inv1  gate2571(.a(G16), .O(gate32inter8));
  nand2 gate2572(.a(gate32inter8), .b(gate32inter7), .O(gate32inter9));
  nand2 gate2573(.a(s_289), .b(gate32inter3), .O(gate32inter10));
  nor2  gate2574(.a(gate32inter10), .b(gate32inter9), .O(gate32inter11));
  nor2  gate2575(.a(gate32inter11), .b(gate32inter6), .O(gate32inter12));
  nand2 gate2576(.a(gate32inter12), .b(gate32inter1), .O(G335));

  xor2  gate1891(.a(G21), .b(G17), .O(gate33inter0));
  nand2 gate1892(.a(gate33inter0), .b(s_192), .O(gate33inter1));
  and2  gate1893(.a(G21), .b(G17), .O(gate33inter2));
  inv1  gate1894(.a(s_192), .O(gate33inter3));
  inv1  gate1895(.a(s_193), .O(gate33inter4));
  nand2 gate1896(.a(gate33inter4), .b(gate33inter3), .O(gate33inter5));
  nor2  gate1897(.a(gate33inter5), .b(gate33inter2), .O(gate33inter6));
  inv1  gate1898(.a(G17), .O(gate33inter7));
  inv1  gate1899(.a(G21), .O(gate33inter8));
  nand2 gate1900(.a(gate33inter8), .b(gate33inter7), .O(gate33inter9));
  nand2 gate1901(.a(s_193), .b(gate33inter3), .O(gate33inter10));
  nor2  gate1902(.a(gate33inter10), .b(gate33inter9), .O(gate33inter11));
  nor2  gate1903(.a(gate33inter11), .b(gate33inter6), .O(gate33inter12));
  nand2 gate1904(.a(gate33inter12), .b(gate33inter1), .O(G338));
nand2 gate34( .a(G25), .b(G29), .O(G341) );

  xor2  gate1541(.a(G22), .b(G18), .O(gate35inter0));
  nand2 gate1542(.a(gate35inter0), .b(s_142), .O(gate35inter1));
  and2  gate1543(.a(G22), .b(G18), .O(gate35inter2));
  inv1  gate1544(.a(s_142), .O(gate35inter3));
  inv1  gate1545(.a(s_143), .O(gate35inter4));
  nand2 gate1546(.a(gate35inter4), .b(gate35inter3), .O(gate35inter5));
  nor2  gate1547(.a(gate35inter5), .b(gate35inter2), .O(gate35inter6));
  inv1  gate1548(.a(G18), .O(gate35inter7));
  inv1  gate1549(.a(G22), .O(gate35inter8));
  nand2 gate1550(.a(gate35inter8), .b(gate35inter7), .O(gate35inter9));
  nand2 gate1551(.a(s_143), .b(gate35inter3), .O(gate35inter10));
  nor2  gate1552(.a(gate35inter10), .b(gate35inter9), .O(gate35inter11));
  nor2  gate1553(.a(gate35inter11), .b(gate35inter6), .O(gate35inter12));
  nand2 gate1554(.a(gate35inter12), .b(gate35inter1), .O(G344));
nand2 gate36( .a(G26), .b(G30), .O(G347) );
nand2 gate37( .a(G19), .b(G23), .O(G350) );
nand2 gate38( .a(G27), .b(G31), .O(G353) );
nand2 gate39( .a(G20), .b(G24), .O(G356) );
nand2 gate40( .a(G28), .b(G32), .O(G359) );
nand2 gate41( .a(G1), .b(G266), .O(G362) );

  xor2  gate2199(.a(G266), .b(G2), .O(gate42inter0));
  nand2 gate2200(.a(gate42inter0), .b(s_236), .O(gate42inter1));
  and2  gate2201(.a(G266), .b(G2), .O(gate42inter2));
  inv1  gate2202(.a(s_236), .O(gate42inter3));
  inv1  gate2203(.a(s_237), .O(gate42inter4));
  nand2 gate2204(.a(gate42inter4), .b(gate42inter3), .O(gate42inter5));
  nor2  gate2205(.a(gate42inter5), .b(gate42inter2), .O(gate42inter6));
  inv1  gate2206(.a(G2), .O(gate42inter7));
  inv1  gate2207(.a(G266), .O(gate42inter8));
  nand2 gate2208(.a(gate42inter8), .b(gate42inter7), .O(gate42inter9));
  nand2 gate2209(.a(s_237), .b(gate42inter3), .O(gate42inter10));
  nor2  gate2210(.a(gate42inter10), .b(gate42inter9), .O(gate42inter11));
  nor2  gate2211(.a(gate42inter11), .b(gate42inter6), .O(gate42inter12));
  nand2 gate2212(.a(gate42inter12), .b(gate42inter1), .O(G363));

  xor2  gate2899(.a(G269), .b(G3), .O(gate43inter0));
  nand2 gate2900(.a(gate43inter0), .b(s_336), .O(gate43inter1));
  and2  gate2901(.a(G269), .b(G3), .O(gate43inter2));
  inv1  gate2902(.a(s_336), .O(gate43inter3));
  inv1  gate2903(.a(s_337), .O(gate43inter4));
  nand2 gate2904(.a(gate43inter4), .b(gate43inter3), .O(gate43inter5));
  nor2  gate2905(.a(gate43inter5), .b(gate43inter2), .O(gate43inter6));
  inv1  gate2906(.a(G3), .O(gate43inter7));
  inv1  gate2907(.a(G269), .O(gate43inter8));
  nand2 gate2908(.a(gate43inter8), .b(gate43inter7), .O(gate43inter9));
  nand2 gate2909(.a(s_337), .b(gate43inter3), .O(gate43inter10));
  nor2  gate2910(.a(gate43inter10), .b(gate43inter9), .O(gate43inter11));
  nor2  gate2911(.a(gate43inter11), .b(gate43inter6), .O(gate43inter12));
  nand2 gate2912(.a(gate43inter12), .b(gate43inter1), .O(G364));

  xor2  gate561(.a(G269), .b(G4), .O(gate44inter0));
  nand2 gate562(.a(gate44inter0), .b(s_2), .O(gate44inter1));
  and2  gate563(.a(G269), .b(G4), .O(gate44inter2));
  inv1  gate564(.a(s_2), .O(gate44inter3));
  inv1  gate565(.a(s_3), .O(gate44inter4));
  nand2 gate566(.a(gate44inter4), .b(gate44inter3), .O(gate44inter5));
  nor2  gate567(.a(gate44inter5), .b(gate44inter2), .O(gate44inter6));
  inv1  gate568(.a(G4), .O(gate44inter7));
  inv1  gate569(.a(G269), .O(gate44inter8));
  nand2 gate570(.a(gate44inter8), .b(gate44inter7), .O(gate44inter9));
  nand2 gate571(.a(s_3), .b(gate44inter3), .O(gate44inter10));
  nor2  gate572(.a(gate44inter10), .b(gate44inter9), .O(gate44inter11));
  nor2  gate573(.a(gate44inter11), .b(gate44inter6), .O(gate44inter12));
  nand2 gate574(.a(gate44inter12), .b(gate44inter1), .O(G365));
nand2 gate45( .a(G5), .b(G272), .O(G366) );
nand2 gate46( .a(G6), .b(G272), .O(G367) );

  xor2  gate1947(.a(G275), .b(G7), .O(gate47inter0));
  nand2 gate1948(.a(gate47inter0), .b(s_200), .O(gate47inter1));
  and2  gate1949(.a(G275), .b(G7), .O(gate47inter2));
  inv1  gate1950(.a(s_200), .O(gate47inter3));
  inv1  gate1951(.a(s_201), .O(gate47inter4));
  nand2 gate1952(.a(gate47inter4), .b(gate47inter3), .O(gate47inter5));
  nor2  gate1953(.a(gate47inter5), .b(gate47inter2), .O(gate47inter6));
  inv1  gate1954(.a(G7), .O(gate47inter7));
  inv1  gate1955(.a(G275), .O(gate47inter8));
  nand2 gate1956(.a(gate47inter8), .b(gate47inter7), .O(gate47inter9));
  nand2 gate1957(.a(s_201), .b(gate47inter3), .O(gate47inter10));
  nor2  gate1958(.a(gate47inter10), .b(gate47inter9), .O(gate47inter11));
  nor2  gate1959(.a(gate47inter11), .b(gate47inter6), .O(gate47inter12));
  nand2 gate1960(.a(gate47inter12), .b(gate47inter1), .O(G368));

  xor2  gate2353(.a(G275), .b(G8), .O(gate48inter0));
  nand2 gate2354(.a(gate48inter0), .b(s_258), .O(gate48inter1));
  and2  gate2355(.a(G275), .b(G8), .O(gate48inter2));
  inv1  gate2356(.a(s_258), .O(gate48inter3));
  inv1  gate2357(.a(s_259), .O(gate48inter4));
  nand2 gate2358(.a(gate48inter4), .b(gate48inter3), .O(gate48inter5));
  nor2  gate2359(.a(gate48inter5), .b(gate48inter2), .O(gate48inter6));
  inv1  gate2360(.a(G8), .O(gate48inter7));
  inv1  gate2361(.a(G275), .O(gate48inter8));
  nand2 gate2362(.a(gate48inter8), .b(gate48inter7), .O(gate48inter9));
  nand2 gate2363(.a(s_259), .b(gate48inter3), .O(gate48inter10));
  nor2  gate2364(.a(gate48inter10), .b(gate48inter9), .O(gate48inter11));
  nor2  gate2365(.a(gate48inter11), .b(gate48inter6), .O(gate48inter12));
  nand2 gate2366(.a(gate48inter12), .b(gate48inter1), .O(G369));

  xor2  gate883(.a(G278), .b(G9), .O(gate49inter0));
  nand2 gate884(.a(gate49inter0), .b(s_48), .O(gate49inter1));
  and2  gate885(.a(G278), .b(G9), .O(gate49inter2));
  inv1  gate886(.a(s_48), .O(gate49inter3));
  inv1  gate887(.a(s_49), .O(gate49inter4));
  nand2 gate888(.a(gate49inter4), .b(gate49inter3), .O(gate49inter5));
  nor2  gate889(.a(gate49inter5), .b(gate49inter2), .O(gate49inter6));
  inv1  gate890(.a(G9), .O(gate49inter7));
  inv1  gate891(.a(G278), .O(gate49inter8));
  nand2 gate892(.a(gate49inter8), .b(gate49inter7), .O(gate49inter9));
  nand2 gate893(.a(s_49), .b(gate49inter3), .O(gate49inter10));
  nor2  gate894(.a(gate49inter10), .b(gate49inter9), .O(gate49inter11));
  nor2  gate895(.a(gate49inter11), .b(gate49inter6), .O(gate49inter12));
  nand2 gate896(.a(gate49inter12), .b(gate49inter1), .O(G370));
nand2 gate50( .a(G10), .b(G278), .O(G371) );
nand2 gate51( .a(G11), .b(G281), .O(G372) );

  xor2  gate2577(.a(G281), .b(G12), .O(gate52inter0));
  nand2 gate2578(.a(gate52inter0), .b(s_290), .O(gate52inter1));
  and2  gate2579(.a(G281), .b(G12), .O(gate52inter2));
  inv1  gate2580(.a(s_290), .O(gate52inter3));
  inv1  gate2581(.a(s_291), .O(gate52inter4));
  nand2 gate2582(.a(gate52inter4), .b(gate52inter3), .O(gate52inter5));
  nor2  gate2583(.a(gate52inter5), .b(gate52inter2), .O(gate52inter6));
  inv1  gate2584(.a(G12), .O(gate52inter7));
  inv1  gate2585(.a(G281), .O(gate52inter8));
  nand2 gate2586(.a(gate52inter8), .b(gate52inter7), .O(gate52inter9));
  nand2 gate2587(.a(s_291), .b(gate52inter3), .O(gate52inter10));
  nor2  gate2588(.a(gate52inter10), .b(gate52inter9), .O(gate52inter11));
  nor2  gate2589(.a(gate52inter11), .b(gate52inter6), .O(gate52inter12));
  nand2 gate2590(.a(gate52inter12), .b(gate52inter1), .O(G373));

  xor2  gate1919(.a(G284), .b(G13), .O(gate53inter0));
  nand2 gate1920(.a(gate53inter0), .b(s_196), .O(gate53inter1));
  and2  gate1921(.a(G284), .b(G13), .O(gate53inter2));
  inv1  gate1922(.a(s_196), .O(gate53inter3));
  inv1  gate1923(.a(s_197), .O(gate53inter4));
  nand2 gate1924(.a(gate53inter4), .b(gate53inter3), .O(gate53inter5));
  nor2  gate1925(.a(gate53inter5), .b(gate53inter2), .O(gate53inter6));
  inv1  gate1926(.a(G13), .O(gate53inter7));
  inv1  gate1927(.a(G284), .O(gate53inter8));
  nand2 gate1928(.a(gate53inter8), .b(gate53inter7), .O(gate53inter9));
  nand2 gate1929(.a(s_197), .b(gate53inter3), .O(gate53inter10));
  nor2  gate1930(.a(gate53inter10), .b(gate53inter9), .O(gate53inter11));
  nor2  gate1931(.a(gate53inter11), .b(gate53inter6), .O(gate53inter12));
  nand2 gate1932(.a(gate53inter12), .b(gate53inter1), .O(G374));
nand2 gate54( .a(G14), .b(G284), .O(G375) );
nand2 gate55( .a(G15), .b(G287), .O(G376) );
nand2 gate56( .a(G16), .b(G287), .O(G377) );
nand2 gate57( .a(G17), .b(G290), .O(G378) );

  xor2  gate911(.a(G290), .b(G18), .O(gate58inter0));
  nand2 gate912(.a(gate58inter0), .b(s_52), .O(gate58inter1));
  and2  gate913(.a(G290), .b(G18), .O(gate58inter2));
  inv1  gate914(.a(s_52), .O(gate58inter3));
  inv1  gate915(.a(s_53), .O(gate58inter4));
  nand2 gate916(.a(gate58inter4), .b(gate58inter3), .O(gate58inter5));
  nor2  gate917(.a(gate58inter5), .b(gate58inter2), .O(gate58inter6));
  inv1  gate918(.a(G18), .O(gate58inter7));
  inv1  gate919(.a(G290), .O(gate58inter8));
  nand2 gate920(.a(gate58inter8), .b(gate58inter7), .O(gate58inter9));
  nand2 gate921(.a(s_53), .b(gate58inter3), .O(gate58inter10));
  nor2  gate922(.a(gate58inter10), .b(gate58inter9), .O(gate58inter11));
  nor2  gate923(.a(gate58inter11), .b(gate58inter6), .O(gate58inter12));
  nand2 gate924(.a(gate58inter12), .b(gate58inter1), .O(G379));
nand2 gate59( .a(G19), .b(G293), .O(G380) );
nand2 gate60( .a(G20), .b(G293), .O(G381) );

  xor2  gate2871(.a(G296), .b(G21), .O(gate61inter0));
  nand2 gate2872(.a(gate61inter0), .b(s_332), .O(gate61inter1));
  and2  gate2873(.a(G296), .b(G21), .O(gate61inter2));
  inv1  gate2874(.a(s_332), .O(gate61inter3));
  inv1  gate2875(.a(s_333), .O(gate61inter4));
  nand2 gate2876(.a(gate61inter4), .b(gate61inter3), .O(gate61inter5));
  nor2  gate2877(.a(gate61inter5), .b(gate61inter2), .O(gate61inter6));
  inv1  gate2878(.a(G21), .O(gate61inter7));
  inv1  gate2879(.a(G296), .O(gate61inter8));
  nand2 gate2880(.a(gate61inter8), .b(gate61inter7), .O(gate61inter9));
  nand2 gate2881(.a(s_333), .b(gate61inter3), .O(gate61inter10));
  nor2  gate2882(.a(gate61inter10), .b(gate61inter9), .O(gate61inter11));
  nor2  gate2883(.a(gate61inter11), .b(gate61inter6), .O(gate61inter12));
  nand2 gate2884(.a(gate61inter12), .b(gate61inter1), .O(G382));
nand2 gate62( .a(G22), .b(G296), .O(G383) );

  xor2  gate771(.a(G299), .b(G23), .O(gate63inter0));
  nand2 gate772(.a(gate63inter0), .b(s_32), .O(gate63inter1));
  and2  gate773(.a(G299), .b(G23), .O(gate63inter2));
  inv1  gate774(.a(s_32), .O(gate63inter3));
  inv1  gate775(.a(s_33), .O(gate63inter4));
  nand2 gate776(.a(gate63inter4), .b(gate63inter3), .O(gate63inter5));
  nor2  gate777(.a(gate63inter5), .b(gate63inter2), .O(gate63inter6));
  inv1  gate778(.a(G23), .O(gate63inter7));
  inv1  gate779(.a(G299), .O(gate63inter8));
  nand2 gate780(.a(gate63inter8), .b(gate63inter7), .O(gate63inter9));
  nand2 gate781(.a(s_33), .b(gate63inter3), .O(gate63inter10));
  nor2  gate782(.a(gate63inter10), .b(gate63inter9), .O(gate63inter11));
  nor2  gate783(.a(gate63inter11), .b(gate63inter6), .O(gate63inter12));
  nand2 gate784(.a(gate63inter12), .b(gate63inter1), .O(G384));
nand2 gate64( .a(G24), .b(G299), .O(G385) );
nand2 gate65( .a(G25), .b(G302), .O(G386) );
nand2 gate66( .a(G26), .b(G302), .O(G387) );

  xor2  gate1835(.a(G305), .b(G27), .O(gate67inter0));
  nand2 gate1836(.a(gate67inter0), .b(s_184), .O(gate67inter1));
  and2  gate1837(.a(G305), .b(G27), .O(gate67inter2));
  inv1  gate1838(.a(s_184), .O(gate67inter3));
  inv1  gate1839(.a(s_185), .O(gate67inter4));
  nand2 gate1840(.a(gate67inter4), .b(gate67inter3), .O(gate67inter5));
  nor2  gate1841(.a(gate67inter5), .b(gate67inter2), .O(gate67inter6));
  inv1  gate1842(.a(G27), .O(gate67inter7));
  inv1  gate1843(.a(G305), .O(gate67inter8));
  nand2 gate1844(.a(gate67inter8), .b(gate67inter7), .O(gate67inter9));
  nand2 gate1845(.a(s_185), .b(gate67inter3), .O(gate67inter10));
  nor2  gate1846(.a(gate67inter10), .b(gate67inter9), .O(gate67inter11));
  nor2  gate1847(.a(gate67inter11), .b(gate67inter6), .O(gate67inter12));
  nand2 gate1848(.a(gate67inter12), .b(gate67inter1), .O(G388));
nand2 gate68( .a(G28), .b(G305), .O(G389) );
nand2 gate69( .a(G29), .b(G308), .O(G390) );
nand2 gate70( .a(G30), .b(G308), .O(G391) );

  xor2  gate2591(.a(G311), .b(G31), .O(gate71inter0));
  nand2 gate2592(.a(gate71inter0), .b(s_292), .O(gate71inter1));
  and2  gate2593(.a(G311), .b(G31), .O(gate71inter2));
  inv1  gate2594(.a(s_292), .O(gate71inter3));
  inv1  gate2595(.a(s_293), .O(gate71inter4));
  nand2 gate2596(.a(gate71inter4), .b(gate71inter3), .O(gate71inter5));
  nor2  gate2597(.a(gate71inter5), .b(gate71inter2), .O(gate71inter6));
  inv1  gate2598(.a(G31), .O(gate71inter7));
  inv1  gate2599(.a(G311), .O(gate71inter8));
  nand2 gate2600(.a(gate71inter8), .b(gate71inter7), .O(gate71inter9));
  nand2 gate2601(.a(s_293), .b(gate71inter3), .O(gate71inter10));
  nor2  gate2602(.a(gate71inter10), .b(gate71inter9), .O(gate71inter11));
  nor2  gate2603(.a(gate71inter11), .b(gate71inter6), .O(gate71inter12));
  nand2 gate2604(.a(gate71inter12), .b(gate71inter1), .O(G392));

  xor2  gate2073(.a(G311), .b(G32), .O(gate72inter0));
  nand2 gate2074(.a(gate72inter0), .b(s_218), .O(gate72inter1));
  and2  gate2075(.a(G311), .b(G32), .O(gate72inter2));
  inv1  gate2076(.a(s_218), .O(gate72inter3));
  inv1  gate2077(.a(s_219), .O(gate72inter4));
  nand2 gate2078(.a(gate72inter4), .b(gate72inter3), .O(gate72inter5));
  nor2  gate2079(.a(gate72inter5), .b(gate72inter2), .O(gate72inter6));
  inv1  gate2080(.a(G32), .O(gate72inter7));
  inv1  gate2081(.a(G311), .O(gate72inter8));
  nand2 gate2082(.a(gate72inter8), .b(gate72inter7), .O(gate72inter9));
  nand2 gate2083(.a(s_219), .b(gate72inter3), .O(gate72inter10));
  nor2  gate2084(.a(gate72inter10), .b(gate72inter9), .O(gate72inter11));
  nor2  gate2085(.a(gate72inter11), .b(gate72inter6), .O(gate72inter12));
  nand2 gate2086(.a(gate72inter12), .b(gate72inter1), .O(G393));
nand2 gate73( .a(G1), .b(G314), .O(G394) );
nand2 gate74( .a(G5), .b(G314), .O(G395) );
nand2 gate75( .a(G9), .b(G317), .O(G396) );
nand2 gate76( .a(G13), .b(G317), .O(G397) );

  xor2  gate1275(.a(G320), .b(G2), .O(gate77inter0));
  nand2 gate1276(.a(gate77inter0), .b(s_104), .O(gate77inter1));
  and2  gate1277(.a(G320), .b(G2), .O(gate77inter2));
  inv1  gate1278(.a(s_104), .O(gate77inter3));
  inv1  gate1279(.a(s_105), .O(gate77inter4));
  nand2 gate1280(.a(gate77inter4), .b(gate77inter3), .O(gate77inter5));
  nor2  gate1281(.a(gate77inter5), .b(gate77inter2), .O(gate77inter6));
  inv1  gate1282(.a(G2), .O(gate77inter7));
  inv1  gate1283(.a(G320), .O(gate77inter8));
  nand2 gate1284(.a(gate77inter8), .b(gate77inter7), .O(gate77inter9));
  nand2 gate1285(.a(s_105), .b(gate77inter3), .O(gate77inter10));
  nor2  gate1286(.a(gate77inter10), .b(gate77inter9), .O(gate77inter11));
  nor2  gate1287(.a(gate77inter11), .b(gate77inter6), .O(gate77inter12));
  nand2 gate1288(.a(gate77inter12), .b(gate77inter1), .O(G398));
nand2 gate78( .a(G6), .b(G320), .O(G399) );
nand2 gate79( .a(G10), .b(G323), .O(G400) );

  xor2  gate1317(.a(G323), .b(G14), .O(gate80inter0));
  nand2 gate1318(.a(gate80inter0), .b(s_110), .O(gate80inter1));
  and2  gate1319(.a(G323), .b(G14), .O(gate80inter2));
  inv1  gate1320(.a(s_110), .O(gate80inter3));
  inv1  gate1321(.a(s_111), .O(gate80inter4));
  nand2 gate1322(.a(gate80inter4), .b(gate80inter3), .O(gate80inter5));
  nor2  gate1323(.a(gate80inter5), .b(gate80inter2), .O(gate80inter6));
  inv1  gate1324(.a(G14), .O(gate80inter7));
  inv1  gate1325(.a(G323), .O(gate80inter8));
  nand2 gate1326(.a(gate80inter8), .b(gate80inter7), .O(gate80inter9));
  nand2 gate1327(.a(s_111), .b(gate80inter3), .O(gate80inter10));
  nor2  gate1328(.a(gate80inter10), .b(gate80inter9), .O(gate80inter11));
  nor2  gate1329(.a(gate80inter11), .b(gate80inter6), .O(gate80inter12));
  nand2 gate1330(.a(gate80inter12), .b(gate80inter1), .O(G401));
nand2 gate81( .a(G3), .b(G326), .O(G402) );

  xor2  gate2983(.a(G326), .b(G7), .O(gate82inter0));
  nand2 gate2984(.a(gate82inter0), .b(s_348), .O(gate82inter1));
  and2  gate2985(.a(G326), .b(G7), .O(gate82inter2));
  inv1  gate2986(.a(s_348), .O(gate82inter3));
  inv1  gate2987(.a(s_349), .O(gate82inter4));
  nand2 gate2988(.a(gate82inter4), .b(gate82inter3), .O(gate82inter5));
  nor2  gate2989(.a(gate82inter5), .b(gate82inter2), .O(gate82inter6));
  inv1  gate2990(.a(G7), .O(gate82inter7));
  inv1  gate2991(.a(G326), .O(gate82inter8));
  nand2 gate2992(.a(gate82inter8), .b(gate82inter7), .O(gate82inter9));
  nand2 gate2993(.a(s_349), .b(gate82inter3), .O(gate82inter10));
  nor2  gate2994(.a(gate82inter10), .b(gate82inter9), .O(gate82inter11));
  nor2  gate2995(.a(gate82inter11), .b(gate82inter6), .O(gate82inter12));
  nand2 gate2996(.a(gate82inter12), .b(gate82inter1), .O(G403));
nand2 gate83( .a(G11), .b(G329), .O(G404) );
nand2 gate84( .a(G15), .b(G329), .O(G405) );

  xor2  gate2773(.a(G332), .b(G4), .O(gate85inter0));
  nand2 gate2774(.a(gate85inter0), .b(s_318), .O(gate85inter1));
  and2  gate2775(.a(G332), .b(G4), .O(gate85inter2));
  inv1  gate2776(.a(s_318), .O(gate85inter3));
  inv1  gate2777(.a(s_319), .O(gate85inter4));
  nand2 gate2778(.a(gate85inter4), .b(gate85inter3), .O(gate85inter5));
  nor2  gate2779(.a(gate85inter5), .b(gate85inter2), .O(gate85inter6));
  inv1  gate2780(.a(G4), .O(gate85inter7));
  inv1  gate2781(.a(G332), .O(gate85inter8));
  nand2 gate2782(.a(gate85inter8), .b(gate85inter7), .O(gate85inter9));
  nand2 gate2783(.a(s_319), .b(gate85inter3), .O(gate85inter10));
  nor2  gate2784(.a(gate85inter10), .b(gate85inter9), .O(gate85inter11));
  nor2  gate2785(.a(gate85inter11), .b(gate85inter6), .O(gate85inter12));
  nand2 gate2786(.a(gate85inter12), .b(gate85inter1), .O(G406));
nand2 gate86( .a(G8), .b(G332), .O(G407) );
nand2 gate87( .a(G12), .b(G335), .O(G408) );

  xor2  gate2367(.a(G335), .b(G16), .O(gate88inter0));
  nand2 gate2368(.a(gate88inter0), .b(s_260), .O(gate88inter1));
  and2  gate2369(.a(G335), .b(G16), .O(gate88inter2));
  inv1  gate2370(.a(s_260), .O(gate88inter3));
  inv1  gate2371(.a(s_261), .O(gate88inter4));
  nand2 gate2372(.a(gate88inter4), .b(gate88inter3), .O(gate88inter5));
  nor2  gate2373(.a(gate88inter5), .b(gate88inter2), .O(gate88inter6));
  inv1  gate2374(.a(G16), .O(gate88inter7));
  inv1  gate2375(.a(G335), .O(gate88inter8));
  nand2 gate2376(.a(gate88inter8), .b(gate88inter7), .O(gate88inter9));
  nand2 gate2377(.a(s_261), .b(gate88inter3), .O(gate88inter10));
  nor2  gate2378(.a(gate88inter10), .b(gate88inter9), .O(gate88inter11));
  nor2  gate2379(.a(gate88inter11), .b(gate88inter6), .O(gate88inter12));
  nand2 gate2380(.a(gate88inter12), .b(gate88inter1), .O(G409));
nand2 gate89( .a(G17), .b(G338), .O(G410) );
nand2 gate90( .a(G21), .b(G338), .O(G411) );
nand2 gate91( .a(G25), .b(G341), .O(G412) );
nand2 gate92( .a(G29), .b(G341), .O(G413) );
nand2 gate93( .a(G18), .b(G344), .O(G414) );
nand2 gate94( .a(G22), .b(G344), .O(G415) );

  xor2  gate939(.a(G347), .b(G26), .O(gate95inter0));
  nand2 gate940(.a(gate95inter0), .b(s_56), .O(gate95inter1));
  and2  gate941(.a(G347), .b(G26), .O(gate95inter2));
  inv1  gate942(.a(s_56), .O(gate95inter3));
  inv1  gate943(.a(s_57), .O(gate95inter4));
  nand2 gate944(.a(gate95inter4), .b(gate95inter3), .O(gate95inter5));
  nor2  gate945(.a(gate95inter5), .b(gate95inter2), .O(gate95inter6));
  inv1  gate946(.a(G26), .O(gate95inter7));
  inv1  gate947(.a(G347), .O(gate95inter8));
  nand2 gate948(.a(gate95inter8), .b(gate95inter7), .O(gate95inter9));
  nand2 gate949(.a(s_57), .b(gate95inter3), .O(gate95inter10));
  nor2  gate950(.a(gate95inter10), .b(gate95inter9), .O(gate95inter11));
  nor2  gate951(.a(gate95inter11), .b(gate95inter6), .O(gate95inter12));
  nand2 gate952(.a(gate95inter12), .b(gate95inter1), .O(G416));

  xor2  gate2913(.a(G347), .b(G30), .O(gate96inter0));
  nand2 gate2914(.a(gate96inter0), .b(s_338), .O(gate96inter1));
  and2  gate2915(.a(G347), .b(G30), .O(gate96inter2));
  inv1  gate2916(.a(s_338), .O(gate96inter3));
  inv1  gate2917(.a(s_339), .O(gate96inter4));
  nand2 gate2918(.a(gate96inter4), .b(gate96inter3), .O(gate96inter5));
  nor2  gate2919(.a(gate96inter5), .b(gate96inter2), .O(gate96inter6));
  inv1  gate2920(.a(G30), .O(gate96inter7));
  inv1  gate2921(.a(G347), .O(gate96inter8));
  nand2 gate2922(.a(gate96inter8), .b(gate96inter7), .O(gate96inter9));
  nand2 gate2923(.a(s_339), .b(gate96inter3), .O(gate96inter10));
  nor2  gate2924(.a(gate96inter10), .b(gate96inter9), .O(gate96inter11));
  nor2  gate2925(.a(gate96inter11), .b(gate96inter6), .O(gate96inter12));
  nand2 gate2926(.a(gate96inter12), .b(gate96inter1), .O(G417));

  xor2  gate1261(.a(G350), .b(G19), .O(gate97inter0));
  nand2 gate1262(.a(gate97inter0), .b(s_102), .O(gate97inter1));
  and2  gate1263(.a(G350), .b(G19), .O(gate97inter2));
  inv1  gate1264(.a(s_102), .O(gate97inter3));
  inv1  gate1265(.a(s_103), .O(gate97inter4));
  nand2 gate1266(.a(gate97inter4), .b(gate97inter3), .O(gate97inter5));
  nor2  gate1267(.a(gate97inter5), .b(gate97inter2), .O(gate97inter6));
  inv1  gate1268(.a(G19), .O(gate97inter7));
  inv1  gate1269(.a(G350), .O(gate97inter8));
  nand2 gate1270(.a(gate97inter8), .b(gate97inter7), .O(gate97inter9));
  nand2 gate1271(.a(s_103), .b(gate97inter3), .O(gate97inter10));
  nor2  gate1272(.a(gate97inter10), .b(gate97inter9), .O(gate97inter11));
  nor2  gate1273(.a(gate97inter11), .b(gate97inter6), .O(gate97inter12));
  nand2 gate1274(.a(gate97inter12), .b(gate97inter1), .O(G418));

  xor2  gate2633(.a(G350), .b(G23), .O(gate98inter0));
  nand2 gate2634(.a(gate98inter0), .b(s_298), .O(gate98inter1));
  and2  gate2635(.a(G350), .b(G23), .O(gate98inter2));
  inv1  gate2636(.a(s_298), .O(gate98inter3));
  inv1  gate2637(.a(s_299), .O(gate98inter4));
  nand2 gate2638(.a(gate98inter4), .b(gate98inter3), .O(gate98inter5));
  nor2  gate2639(.a(gate98inter5), .b(gate98inter2), .O(gate98inter6));
  inv1  gate2640(.a(G23), .O(gate98inter7));
  inv1  gate2641(.a(G350), .O(gate98inter8));
  nand2 gate2642(.a(gate98inter8), .b(gate98inter7), .O(gate98inter9));
  nand2 gate2643(.a(s_299), .b(gate98inter3), .O(gate98inter10));
  nor2  gate2644(.a(gate98inter10), .b(gate98inter9), .O(gate98inter11));
  nor2  gate2645(.a(gate98inter11), .b(gate98inter6), .O(gate98inter12));
  nand2 gate2646(.a(gate98inter12), .b(gate98inter1), .O(G419));
nand2 gate99( .a(G27), .b(G353), .O(G420) );

  xor2  gate729(.a(G353), .b(G31), .O(gate100inter0));
  nand2 gate730(.a(gate100inter0), .b(s_26), .O(gate100inter1));
  and2  gate731(.a(G353), .b(G31), .O(gate100inter2));
  inv1  gate732(.a(s_26), .O(gate100inter3));
  inv1  gate733(.a(s_27), .O(gate100inter4));
  nand2 gate734(.a(gate100inter4), .b(gate100inter3), .O(gate100inter5));
  nor2  gate735(.a(gate100inter5), .b(gate100inter2), .O(gate100inter6));
  inv1  gate736(.a(G31), .O(gate100inter7));
  inv1  gate737(.a(G353), .O(gate100inter8));
  nand2 gate738(.a(gate100inter8), .b(gate100inter7), .O(gate100inter9));
  nand2 gate739(.a(s_27), .b(gate100inter3), .O(gate100inter10));
  nor2  gate740(.a(gate100inter10), .b(gate100inter9), .O(gate100inter11));
  nor2  gate741(.a(gate100inter11), .b(gate100inter6), .O(gate100inter12));
  nand2 gate742(.a(gate100inter12), .b(gate100inter1), .O(G421));

  xor2  gate659(.a(G356), .b(G20), .O(gate101inter0));
  nand2 gate660(.a(gate101inter0), .b(s_16), .O(gate101inter1));
  and2  gate661(.a(G356), .b(G20), .O(gate101inter2));
  inv1  gate662(.a(s_16), .O(gate101inter3));
  inv1  gate663(.a(s_17), .O(gate101inter4));
  nand2 gate664(.a(gate101inter4), .b(gate101inter3), .O(gate101inter5));
  nor2  gate665(.a(gate101inter5), .b(gate101inter2), .O(gate101inter6));
  inv1  gate666(.a(G20), .O(gate101inter7));
  inv1  gate667(.a(G356), .O(gate101inter8));
  nand2 gate668(.a(gate101inter8), .b(gate101inter7), .O(gate101inter9));
  nand2 gate669(.a(s_17), .b(gate101inter3), .O(gate101inter10));
  nor2  gate670(.a(gate101inter10), .b(gate101inter9), .O(gate101inter11));
  nor2  gate671(.a(gate101inter11), .b(gate101inter6), .O(gate101inter12));
  nand2 gate672(.a(gate101inter12), .b(gate101inter1), .O(G422));

  xor2  gate1345(.a(G356), .b(G24), .O(gate102inter0));
  nand2 gate1346(.a(gate102inter0), .b(s_114), .O(gate102inter1));
  and2  gate1347(.a(G356), .b(G24), .O(gate102inter2));
  inv1  gate1348(.a(s_114), .O(gate102inter3));
  inv1  gate1349(.a(s_115), .O(gate102inter4));
  nand2 gate1350(.a(gate102inter4), .b(gate102inter3), .O(gate102inter5));
  nor2  gate1351(.a(gate102inter5), .b(gate102inter2), .O(gate102inter6));
  inv1  gate1352(.a(G24), .O(gate102inter7));
  inv1  gate1353(.a(G356), .O(gate102inter8));
  nand2 gate1354(.a(gate102inter8), .b(gate102inter7), .O(gate102inter9));
  nand2 gate1355(.a(s_115), .b(gate102inter3), .O(gate102inter10));
  nor2  gate1356(.a(gate102inter10), .b(gate102inter9), .O(gate102inter11));
  nor2  gate1357(.a(gate102inter11), .b(gate102inter6), .O(gate102inter12));
  nand2 gate1358(.a(gate102inter12), .b(gate102inter1), .O(G423));
nand2 gate103( .a(G28), .b(G359), .O(G424) );
nand2 gate104( .a(G32), .b(G359), .O(G425) );
nand2 gate105( .a(G362), .b(G363), .O(G426) );
nand2 gate106( .a(G364), .b(G365), .O(G429) );
nand2 gate107( .a(G366), .b(G367), .O(G432) );
nand2 gate108( .a(G368), .b(G369), .O(G435) );
nand2 gate109( .a(G370), .b(G371), .O(G438) );
nand2 gate110( .a(G372), .b(G373), .O(G441) );

  xor2  gate2423(.a(G375), .b(G374), .O(gate111inter0));
  nand2 gate2424(.a(gate111inter0), .b(s_268), .O(gate111inter1));
  and2  gate2425(.a(G375), .b(G374), .O(gate111inter2));
  inv1  gate2426(.a(s_268), .O(gate111inter3));
  inv1  gate2427(.a(s_269), .O(gate111inter4));
  nand2 gate2428(.a(gate111inter4), .b(gate111inter3), .O(gate111inter5));
  nor2  gate2429(.a(gate111inter5), .b(gate111inter2), .O(gate111inter6));
  inv1  gate2430(.a(G374), .O(gate111inter7));
  inv1  gate2431(.a(G375), .O(gate111inter8));
  nand2 gate2432(.a(gate111inter8), .b(gate111inter7), .O(gate111inter9));
  nand2 gate2433(.a(s_269), .b(gate111inter3), .O(gate111inter10));
  nor2  gate2434(.a(gate111inter10), .b(gate111inter9), .O(gate111inter11));
  nor2  gate2435(.a(gate111inter11), .b(gate111inter6), .O(gate111inter12));
  nand2 gate2436(.a(gate111inter12), .b(gate111inter1), .O(G444));
nand2 gate112( .a(G376), .b(G377), .O(G447) );

  xor2  gate1331(.a(G379), .b(G378), .O(gate113inter0));
  nand2 gate1332(.a(gate113inter0), .b(s_112), .O(gate113inter1));
  and2  gate1333(.a(G379), .b(G378), .O(gate113inter2));
  inv1  gate1334(.a(s_112), .O(gate113inter3));
  inv1  gate1335(.a(s_113), .O(gate113inter4));
  nand2 gate1336(.a(gate113inter4), .b(gate113inter3), .O(gate113inter5));
  nor2  gate1337(.a(gate113inter5), .b(gate113inter2), .O(gate113inter6));
  inv1  gate1338(.a(G378), .O(gate113inter7));
  inv1  gate1339(.a(G379), .O(gate113inter8));
  nand2 gate1340(.a(gate113inter8), .b(gate113inter7), .O(gate113inter9));
  nand2 gate1341(.a(s_113), .b(gate113inter3), .O(gate113inter10));
  nor2  gate1342(.a(gate113inter10), .b(gate113inter9), .O(gate113inter11));
  nor2  gate1343(.a(gate113inter11), .b(gate113inter6), .O(gate113inter12));
  nand2 gate1344(.a(gate113inter12), .b(gate113inter1), .O(G450));
nand2 gate114( .a(G380), .b(G381), .O(G453) );
nand2 gate115( .a(G382), .b(G383), .O(G456) );

  xor2  gate2815(.a(G385), .b(G384), .O(gate116inter0));
  nand2 gate2816(.a(gate116inter0), .b(s_324), .O(gate116inter1));
  and2  gate2817(.a(G385), .b(G384), .O(gate116inter2));
  inv1  gate2818(.a(s_324), .O(gate116inter3));
  inv1  gate2819(.a(s_325), .O(gate116inter4));
  nand2 gate2820(.a(gate116inter4), .b(gate116inter3), .O(gate116inter5));
  nor2  gate2821(.a(gate116inter5), .b(gate116inter2), .O(gate116inter6));
  inv1  gate2822(.a(G384), .O(gate116inter7));
  inv1  gate2823(.a(G385), .O(gate116inter8));
  nand2 gate2824(.a(gate116inter8), .b(gate116inter7), .O(gate116inter9));
  nand2 gate2825(.a(s_325), .b(gate116inter3), .O(gate116inter10));
  nor2  gate2826(.a(gate116inter10), .b(gate116inter9), .O(gate116inter11));
  nor2  gate2827(.a(gate116inter11), .b(gate116inter6), .O(gate116inter12));
  nand2 gate2828(.a(gate116inter12), .b(gate116inter1), .O(G459));

  xor2  gate603(.a(G387), .b(G386), .O(gate117inter0));
  nand2 gate604(.a(gate117inter0), .b(s_8), .O(gate117inter1));
  and2  gate605(.a(G387), .b(G386), .O(gate117inter2));
  inv1  gate606(.a(s_8), .O(gate117inter3));
  inv1  gate607(.a(s_9), .O(gate117inter4));
  nand2 gate608(.a(gate117inter4), .b(gate117inter3), .O(gate117inter5));
  nor2  gate609(.a(gate117inter5), .b(gate117inter2), .O(gate117inter6));
  inv1  gate610(.a(G386), .O(gate117inter7));
  inv1  gate611(.a(G387), .O(gate117inter8));
  nand2 gate612(.a(gate117inter8), .b(gate117inter7), .O(gate117inter9));
  nand2 gate613(.a(s_9), .b(gate117inter3), .O(gate117inter10));
  nor2  gate614(.a(gate117inter10), .b(gate117inter9), .O(gate117inter11));
  nor2  gate615(.a(gate117inter11), .b(gate117inter6), .O(gate117inter12));
  nand2 gate616(.a(gate117inter12), .b(gate117inter1), .O(G462));
nand2 gate118( .a(G388), .b(G389), .O(G465) );

  xor2  gate2997(.a(G391), .b(G390), .O(gate119inter0));
  nand2 gate2998(.a(gate119inter0), .b(s_350), .O(gate119inter1));
  and2  gate2999(.a(G391), .b(G390), .O(gate119inter2));
  inv1  gate3000(.a(s_350), .O(gate119inter3));
  inv1  gate3001(.a(s_351), .O(gate119inter4));
  nand2 gate3002(.a(gate119inter4), .b(gate119inter3), .O(gate119inter5));
  nor2  gate3003(.a(gate119inter5), .b(gate119inter2), .O(gate119inter6));
  inv1  gate3004(.a(G390), .O(gate119inter7));
  inv1  gate3005(.a(G391), .O(gate119inter8));
  nand2 gate3006(.a(gate119inter8), .b(gate119inter7), .O(gate119inter9));
  nand2 gate3007(.a(s_351), .b(gate119inter3), .O(gate119inter10));
  nor2  gate3008(.a(gate119inter10), .b(gate119inter9), .O(gate119inter11));
  nor2  gate3009(.a(gate119inter11), .b(gate119inter6), .O(gate119inter12));
  nand2 gate3010(.a(gate119inter12), .b(gate119inter1), .O(G468));

  xor2  gate1471(.a(G393), .b(G392), .O(gate120inter0));
  nand2 gate1472(.a(gate120inter0), .b(s_132), .O(gate120inter1));
  and2  gate1473(.a(G393), .b(G392), .O(gate120inter2));
  inv1  gate1474(.a(s_132), .O(gate120inter3));
  inv1  gate1475(.a(s_133), .O(gate120inter4));
  nand2 gate1476(.a(gate120inter4), .b(gate120inter3), .O(gate120inter5));
  nor2  gate1477(.a(gate120inter5), .b(gate120inter2), .O(gate120inter6));
  inv1  gate1478(.a(G392), .O(gate120inter7));
  inv1  gate1479(.a(G393), .O(gate120inter8));
  nand2 gate1480(.a(gate120inter8), .b(gate120inter7), .O(gate120inter9));
  nand2 gate1481(.a(s_133), .b(gate120inter3), .O(gate120inter10));
  nor2  gate1482(.a(gate120inter10), .b(gate120inter9), .O(gate120inter11));
  nor2  gate1483(.a(gate120inter11), .b(gate120inter6), .O(gate120inter12));
  nand2 gate1484(.a(gate120inter12), .b(gate120inter1), .O(G471));

  xor2  gate2647(.a(G395), .b(G394), .O(gate121inter0));
  nand2 gate2648(.a(gate121inter0), .b(s_300), .O(gate121inter1));
  and2  gate2649(.a(G395), .b(G394), .O(gate121inter2));
  inv1  gate2650(.a(s_300), .O(gate121inter3));
  inv1  gate2651(.a(s_301), .O(gate121inter4));
  nand2 gate2652(.a(gate121inter4), .b(gate121inter3), .O(gate121inter5));
  nor2  gate2653(.a(gate121inter5), .b(gate121inter2), .O(gate121inter6));
  inv1  gate2654(.a(G394), .O(gate121inter7));
  inv1  gate2655(.a(G395), .O(gate121inter8));
  nand2 gate2656(.a(gate121inter8), .b(gate121inter7), .O(gate121inter9));
  nand2 gate2657(.a(s_301), .b(gate121inter3), .O(gate121inter10));
  nor2  gate2658(.a(gate121inter10), .b(gate121inter9), .O(gate121inter11));
  nor2  gate2659(.a(gate121inter11), .b(gate121inter6), .O(gate121inter12));
  nand2 gate2660(.a(gate121inter12), .b(gate121inter1), .O(G474));
nand2 gate122( .a(G396), .b(G397), .O(G477) );

  xor2  gate2213(.a(G399), .b(G398), .O(gate123inter0));
  nand2 gate2214(.a(gate123inter0), .b(s_238), .O(gate123inter1));
  and2  gate2215(.a(G399), .b(G398), .O(gate123inter2));
  inv1  gate2216(.a(s_238), .O(gate123inter3));
  inv1  gate2217(.a(s_239), .O(gate123inter4));
  nand2 gate2218(.a(gate123inter4), .b(gate123inter3), .O(gate123inter5));
  nor2  gate2219(.a(gate123inter5), .b(gate123inter2), .O(gate123inter6));
  inv1  gate2220(.a(G398), .O(gate123inter7));
  inv1  gate2221(.a(G399), .O(gate123inter8));
  nand2 gate2222(.a(gate123inter8), .b(gate123inter7), .O(gate123inter9));
  nand2 gate2223(.a(s_239), .b(gate123inter3), .O(gate123inter10));
  nor2  gate2224(.a(gate123inter10), .b(gate123inter9), .O(gate123inter11));
  nor2  gate2225(.a(gate123inter11), .b(gate123inter6), .O(gate123inter12));
  nand2 gate2226(.a(gate123inter12), .b(gate123inter1), .O(G480));

  xor2  gate2955(.a(G401), .b(G400), .O(gate124inter0));
  nand2 gate2956(.a(gate124inter0), .b(s_344), .O(gate124inter1));
  and2  gate2957(.a(G401), .b(G400), .O(gate124inter2));
  inv1  gate2958(.a(s_344), .O(gate124inter3));
  inv1  gate2959(.a(s_345), .O(gate124inter4));
  nand2 gate2960(.a(gate124inter4), .b(gate124inter3), .O(gate124inter5));
  nor2  gate2961(.a(gate124inter5), .b(gate124inter2), .O(gate124inter6));
  inv1  gate2962(.a(G400), .O(gate124inter7));
  inv1  gate2963(.a(G401), .O(gate124inter8));
  nand2 gate2964(.a(gate124inter8), .b(gate124inter7), .O(gate124inter9));
  nand2 gate2965(.a(s_345), .b(gate124inter3), .O(gate124inter10));
  nor2  gate2966(.a(gate124inter10), .b(gate124inter9), .O(gate124inter11));
  nor2  gate2967(.a(gate124inter11), .b(gate124inter6), .O(gate124inter12));
  nand2 gate2968(.a(gate124inter12), .b(gate124inter1), .O(G483));
nand2 gate125( .a(G402), .b(G403), .O(G486) );

  xor2  gate1219(.a(G405), .b(G404), .O(gate126inter0));
  nand2 gate1220(.a(gate126inter0), .b(s_96), .O(gate126inter1));
  and2  gate1221(.a(G405), .b(G404), .O(gate126inter2));
  inv1  gate1222(.a(s_96), .O(gate126inter3));
  inv1  gate1223(.a(s_97), .O(gate126inter4));
  nand2 gate1224(.a(gate126inter4), .b(gate126inter3), .O(gate126inter5));
  nor2  gate1225(.a(gate126inter5), .b(gate126inter2), .O(gate126inter6));
  inv1  gate1226(.a(G404), .O(gate126inter7));
  inv1  gate1227(.a(G405), .O(gate126inter8));
  nand2 gate1228(.a(gate126inter8), .b(gate126inter7), .O(gate126inter9));
  nand2 gate1229(.a(s_97), .b(gate126inter3), .O(gate126inter10));
  nor2  gate1230(.a(gate126inter10), .b(gate126inter9), .O(gate126inter11));
  nor2  gate1231(.a(gate126inter11), .b(gate126inter6), .O(gate126inter12));
  nand2 gate1232(.a(gate126inter12), .b(gate126inter1), .O(G489));
nand2 gate127( .a(G406), .b(G407), .O(G492) );

  xor2  gate855(.a(G409), .b(G408), .O(gate128inter0));
  nand2 gate856(.a(gate128inter0), .b(s_44), .O(gate128inter1));
  and2  gate857(.a(G409), .b(G408), .O(gate128inter2));
  inv1  gate858(.a(s_44), .O(gate128inter3));
  inv1  gate859(.a(s_45), .O(gate128inter4));
  nand2 gate860(.a(gate128inter4), .b(gate128inter3), .O(gate128inter5));
  nor2  gate861(.a(gate128inter5), .b(gate128inter2), .O(gate128inter6));
  inv1  gate862(.a(G408), .O(gate128inter7));
  inv1  gate863(.a(G409), .O(gate128inter8));
  nand2 gate864(.a(gate128inter8), .b(gate128inter7), .O(gate128inter9));
  nand2 gate865(.a(s_45), .b(gate128inter3), .O(gate128inter10));
  nor2  gate866(.a(gate128inter10), .b(gate128inter9), .O(gate128inter11));
  nor2  gate867(.a(gate128inter11), .b(gate128inter6), .O(gate128inter12));
  nand2 gate868(.a(gate128inter12), .b(gate128inter1), .O(G495));

  xor2  gate2395(.a(G411), .b(G410), .O(gate129inter0));
  nand2 gate2396(.a(gate129inter0), .b(s_264), .O(gate129inter1));
  and2  gate2397(.a(G411), .b(G410), .O(gate129inter2));
  inv1  gate2398(.a(s_264), .O(gate129inter3));
  inv1  gate2399(.a(s_265), .O(gate129inter4));
  nand2 gate2400(.a(gate129inter4), .b(gate129inter3), .O(gate129inter5));
  nor2  gate2401(.a(gate129inter5), .b(gate129inter2), .O(gate129inter6));
  inv1  gate2402(.a(G410), .O(gate129inter7));
  inv1  gate2403(.a(G411), .O(gate129inter8));
  nand2 gate2404(.a(gate129inter8), .b(gate129inter7), .O(gate129inter9));
  nand2 gate2405(.a(s_265), .b(gate129inter3), .O(gate129inter10));
  nor2  gate2406(.a(gate129inter10), .b(gate129inter9), .O(gate129inter11));
  nor2  gate2407(.a(gate129inter11), .b(gate129inter6), .O(gate129inter12));
  nand2 gate2408(.a(gate129inter12), .b(gate129inter1), .O(G498));
nand2 gate130( .a(G412), .b(G413), .O(G501) );

  xor2  gate2605(.a(G415), .b(G414), .O(gate131inter0));
  nand2 gate2606(.a(gate131inter0), .b(s_294), .O(gate131inter1));
  and2  gate2607(.a(G415), .b(G414), .O(gate131inter2));
  inv1  gate2608(.a(s_294), .O(gate131inter3));
  inv1  gate2609(.a(s_295), .O(gate131inter4));
  nand2 gate2610(.a(gate131inter4), .b(gate131inter3), .O(gate131inter5));
  nor2  gate2611(.a(gate131inter5), .b(gate131inter2), .O(gate131inter6));
  inv1  gate2612(.a(G414), .O(gate131inter7));
  inv1  gate2613(.a(G415), .O(gate131inter8));
  nand2 gate2614(.a(gate131inter8), .b(gate131inter7), .O(gate131inter9));
  nand2 gate2615(.a(s_295), .b(gate131inter3), .O(gate131inter10));
  nor2  gate2616(.a(gate131inter10), .b(gate131inter9), .O(gate131inter11));
  nor2  gate2617(.a(gate131inter11), .b(gate131inter6), .O(gate131inter12));
  nand2 gate2618(.a(gate131inter12), .b(gate131inter1), .O(G504));
nand2 gate132( .a(G416), .b(G417), .O(G507) );
nand2 gate133( .a(G418), .b(G419), .O(G510) );
nand2 gate134( .a(G420), .b(G421), .O(G513) );

  xor2  gate2731(.a(G423), .b(G422), .O(gate135inter0));
  nand2 gate2732(.a(gate135inter0), .b(s_312), .O(gate135inter1));
  and2  gate2733(.a(G423), .b(G422), .O(gate135inter2));
  inv1  gate2734(.a(s_312), .O(gate135inter3));
  inv1  gate2735(.a(s_313), .O(gate135inter4));
  nand2 gate2736(.a(gate135inter4), .b(gate135inter3), .O(gate135inter5));
  nor2  gate2737(.a(gate135inter5), .b(gate135inter2), .O(gate135inter6));
  inv1  gate2738(.a(G422), .O(gate135inter7));
  inv1  gate2739(.a(G423), .O(gate135inter8));
  nand2 gate2740(.a(gate135inter8), .b(gate135inter7), .O(gate135inter9));
  nand2 gate2741(.a(s_313), .b(gate135inter3), .O(gate135inter10));
  nor2  gate2742(.a(gate135inter10), .b(gate135inter9), .O(gate135inter11));
  nor2  gate2743(.a(gate135inter11), .b(gate135inter6), .O(gate135inter12));
  nand2 gate2744(.a(gate135inter12), .b(gate135inter1), .O(G516));
nand2 gate136( .a(G424), .b(G425), .O(G519) );
nand2 gate137( .a(G426), .b(G429), .O(G522) );
nand2 gate138( .a(G432), .b(G435), .O(G525) );

  xor2  gate1905(.a(G441), .b(G438), .O(gate139inter0));
  nand2 gate1906(.a(gate139inter0), .b(s_194), .O(gate139inter1));
  and2  gate1907(.a(G441), .b(G438), .O(gate139inter2));
  inv1  gate1908(.a(s_194), .O(gate139inter3));
  inv1  gate1909(.a(s_195), .O(gate139inter4));
  nand2 gate1910(.a(gate139inter4), .b(gate139inter3), .O(gate139inter5));
  nor2  gate1911(.a(gate139inter5), .b(gate139inter2), .O(gate139inter6));
  inv1  gate1912(.a(G438), .O(gate139inter7));
  inv1  gate1913(.a(G441), .O(gate139inter8));
  nand2 gate1914(.a(gate139inter8), .b(gate139inter7), .O(gate139inter9));
  nand2 gate1915(.a(s_195), .b(gate139inter3), .O(gate139inter10));
  nor2  gate1916(.a(gate139inter10), .b(gate139inter9), .O(gate139inter11));
  nor2  gate1917(.a(gate139inter11), .b(gate139inter6), .O(gate139inter12));
  nand2 gate1918(.a(gate139inter12), .b(gate139inter1), .O(G528));
nand2 gate140( .a(G444), .b(G447), .O(G531) );
nand2 gate141( .a(G450), .b(G453), .O(G534) );

  xor2  gate2941(.a(G459), .b(G456), .O(gate142inter0));
  nand2 gate2942(.a(gate142inter0), .b(s_342), .O(gate142inter1));
  and2  gate2943(.a(G459), .b(G456), .O(gate142inter2));
  inv1  gate2944(.a(s_342), .O(gate142inter3));
  inv1  gate2945(.a(s_343), .O(gate142inter4));
  nand2 gate2946(.a(gate142inter4), .b(gate142inter3), .O(gate142inter5));
  nor2  gate2947(.a(gate142inter5), .b(gate142inter2), .O(gate142inter6));
  inv1  gate2948(.a(G456), .O(gate142inter7));
  inv1  gate2949(.a(G459), .O(gate142inter8));
  nand2 gate2950(.a(gate142inter8), .b(gate142inter7), .O(gate142inter9));
  nand2 gate2951(.a(s_343), .b(gate142inter3), .O(gate142inter10));
  nor2  gate2952(.a(gate142inter10), .b(gate142inter9), .O(gate142inter11));
  nor2  gate2953(.a(gate142inter11), .b(gate142inter6), .O(gate142inter12));
  nand2 gate2954(.a(gate142inter12), .b(gate142inter1), .O(G537));

  xor2  gate1695(.a(G465), .b(G462), .O(gate143inter0));
  nand2 gate1696(.a(gate143inter0), .b(s_164), .O(gate143inter1));
  and2  gate1697(.a(G465), .b(G462), .O(gate143inter2));
  inv1  gate1698(.a(s_164), .O(gate143inter3));
  inv1  gate1699(.a(s_165), .O(gate143inter4));
  nand2 gate1700(.a(gate143inter4), .b(gate143inter3), .O(gate143inter5));
  nor2  gate1701(.a(gate143inter5), .b(gate143inter2), .O(gate143inter6));
  inv1  gate1702(.a(G462), .O(gate143inter7));
  inv1  gate1703(.a(G465), .O(gate143inter8));
  nand2 gate1704(.a(gate143inter8), .b(gate143inter7), .O(gate143inter9));
  nand2 gate1705(.a(s_165), .b(gate143inter3), .O(gate143inter10));
  nor2  gate1706(.a(gate143inter10), .b(gate143inter9), .O(gate143inter11));
  nor2  gate1707(.a(gate143inter11), .b(gate143inter6), .O(gate143inter12));
  nand2 gate1708(.a(gate143inter12), .b(gate143inter1), .O(G540));

  xor2  gate1289(.a(G471), .b(G468), .O(gate144inter0));
  nand2 gate1290(.a(gate144inter0), .b(s_106), .O(gate144inter1));
  and2  gate1291(.a(G471), .b(G468), .O(gate144inter2));
  inv1  gate1292(.a(s_106), .O(gate144inter3));
  inv1  gate1293(.a(s_107), .O(gate144inter4));
  nand2 gate1294(.a(gate144inter4), .b(gate144inter3), .O(gate144inter5));
  nor2  gate1295(.a(gate144inter5), .b(gate144inter2), .O(gate144inter6));
  inv1  gate1296(.a(G468), .O(gate144inter7));
  inv1  gate1297(.a(G471), .O(gate144inter8));
  nand2 gate1298(.a(gate144inter8), .b(gate144inter7), .O(gate144inter9));
  nand2 gate1299(.a(s_107), .b(gate144inter3), .O(gate144inter10));
  nor2  gate1300(.a(gate144inter10), .b(gate144inter9), .O(gate144inter11));
  nor2  gate1301(.a(gate144inter11), .b(gate144inter6), .O(gate144inter12));
  nand2 gate1302(.a(gate144inter12), .b(gate144inter1), .O(G543));

  xor2  gate673(.a(G477), .b(G474), .O(gate145inter0));
  nand2 gate674(.a(gate145inter0), .b(s_18), .O(gate145inter1));
  and2  gate675(.a(G477), .b(G474), .O(gate145inter2));
  inv1  gate676(.a(s_18), .O(gate145inter3));
  inv1  gate677(.a(s_19), .O(gate145inter4));
  nand2 gate678(.a(gate145inter4), .b(gate145inter3), .O(gate145inter5));
  nor2  gate679(.a(gate145inter5), .b(gate145inter2), .O(gate145inter6));
  inv1  gate680(.a(G474), .O(gate145inter7));
  inv1  gate681(.a(G477), .O(gate145inter8));
  nand2 gate682(.a(gate145inter8), .b(gate145inter7), .O(gate145inter9));
  nand2 gate683(.a(s_19), .b(gate145inter3), .O(gate145inter10));
  nor2  gate684(.a(gate145inter10), .b(gate145inter9), .O(gate145inter11));
  nor2  gate685(.a(gate145inter11), .b(gate145inter6), .O(gate145inter12));
  nand2 gate686(.a(gate145inter12), .b(gate145inter1), .O(G546));
nand2 gate146( .a(G480), .b(G483), .O(G549) );

  xor2  gate1989(.a(G489), .b(G486), .O(gate147inter0));
  nand2 gate1990(.a(gate147inter0), .b(s_206), .O(gate147inter1));
  and2  gate1991(.a(G489), .b(G486), .O(gate147inter2));
  inv1  gate1992(.a(s_206), .O(gate147inter3));
  inv1  gate1993(.a(s_207), .O(gate147inter4));
  nand2 gate1994(.a(gate147inter4), .b(gate147inter3), .O(gate147inter5));
  nor2  gate1995(.a(gate147inter5), .b(gate147inter2), .O(gate147inter6));
  inv1  gate1996(.a(G486), .O(gate147inter7));
  inv1  gate1997(.a(G489), .O(gate147inter8));
  nand2 gate1998(.a(gate147inter8), .b(gate147inter7), .O(gate147inter9));
  nand2 gate1999(.a(s_207), .b(gate147inter3), .O(gate147inter10));
  nor2  gate2000(.a(gate147inter10), .b(gate147inter9), .O(gate147inter11));
  nor2  gate2001(.a(gate147inter11), .b(gate147inter6), .O(gate147inter12));
  nand2 gate2002(.a(gate147inter12), .b(gate147inter1), .O(G552));
nand2 gate148( .a(G492), .b(G495), .O(G555) );
nand2 gate149( .a(G498), .b(G501), .O(G558) );
nand2 gate150( .a(G504), .b(G507), .O(G561) );
nand2 gate151( .a(G510), .b(G513), .O(G564) );
nand2 gate152( .a(G516), .b(G519), .O(G567) );
nand2 gate153( .a(G426), .b(G522), .O(G570) );
nand2 gate154( .a(G429), .b(G522), .O(G571) );
nand2 gate155( .a(G432), .b(G525), .O(G572) );
nand2 gate156( .a(G435), .b(G525), .O(G573) );

  xor2  gate1205(.a(G528), .b(G438), .O(gate157inter0));
  nand2 gate1206(.a(gate157inter0), .b(s_94), .O(gate157inter1));
  and2  gate1207(.a(G528), .b(G438), .O(gate157inter2));
  inv1  gate1208(.a(s_94), .O(gate157inter3));
  inv1  gate1209(.a(s_95), .O(gate157inter4));
  nand2 gate1210(.a(gate157inter4), .b(gate157inter3), .O(gate157inter5));
  nor2  gate1211(.a(gate157inter5), .b(gate157inter2), .O(gate157inter6));
  inv1  gate1212(.a(G438), .O(gate157inter7));
  inv1  gate1213(.a(G528), .O(gate157inter8));
  nand2 gate1214(.a(gate157inter8), .b(gate157inter7), .O(gate157inter9));
  nand2 gate1215(.a(s_95), .b(gate157inter3), .O(gate157inter10));
  nor2  gate1216(.a(gate157inter10), .b(gate157inter9), .O(gate157inter11));
  nor2  gate1217(.a(gate157inter11), .b(gate157inter6), .O(gate157inter12));
  nand2 gate1218(.a(gate157inter12), .b(gate157inter1), .O(G574));
nand2 gate158( .a(G441), .b(G528), .O(G575) );

  xor2  gate2507(.a(G531), .b(G444), .O(gate159inter0));
  nand2 gate2508(.a(gate159inter0), .b(s_280), .O(gate159inter1));
  and2  gate2509(.a(G531), .b(G444), .O(gate159inter2));
  inv1  gate2510(.a(s_280), .O(gate159inter3));
  inv1  gate2511(.a(s_281), .O(gate159inter4));
  nand2 gate2512(.a(gate159inter4), .b(gate159inter3), .O(gate159inter5));
  nor2  gate2513(.a(gate159inter5), .b(gate159inter2), .O(gate159inter6));
  inv1  gate2514(.a(G444), .O(gate159inter7));
  inv1  gate2515(.a(G531), .O(gate159inter8));
  nand2 gate2516(.a(gate159inter8), .b(gate159inter7), .O(gate159inter9));
  nand2 gate2517(.a(s_281), .b(gate159inter3), .O(gate159inter10));
  nor2  gate2518(.a(gate159inter10), .b(gate159inter9), .O(gate159inter11));
  nor2  gate2519(.a(gate159inter11), .b(gate159inter6), .O(gate159inter12));
  nand2 gate2520(.a(gate159inter12), .b(gate159inter1), .O(G576));

  xor2  gate1653(.a(G531), .b(G447), .O(gate160inter0));
  nand2 gate1654(.a(gate160inter0), .b(s_158), .O(gate160inter1));
  and2  gate1655(.a(G531), .b(G447), .O(gate160inter2));
  inv1  gate1656(.a(s_158), .O(gate160inter3));
  inv1  gate1657(.a(s_159), .O(gate160inter4));
  nand2 gate1658(.a(gate160inter4), .b(gate160inter3), .O(gate160inter5));
  nor2  gate1659(.a(gate160inter5), .b(gate160inter2), .O(gate160inter6));
  inv1  gate1660(.a(G447), .O(gate160inter7));
  inv1  gate1661(.a(G531), .O(gate160inter8));
  nand2 gate1662(.a(gate160inter8), .b(gate160inter7), .O(gate160inter9));
  nand2 gate1663(.a(s_159), .b(gate160inter3), .O(gate160inter10));
  nor2  gate1664(.a(gate160inter10), .b(gate160inter9), .O(gate160inter11));
  nor2  gate1665(.a(gate160inter11), .b(gate160inter6), .O(gate160inter12));
  nand2 gate1666(.a(gate160inter12), .b(gate160inter1), .O(G577));

  xor2  gate1765(.a(G534), .b(G450), .O(gate161inter0));
  nand2 gate1766(.a(gate161inter0), .b(s_174), .O(gate161inter1));
  and2  gate1767(.a(G534), .b(G450), .O(gate161inter2));
  inv1  gate1768(.a(s_174), .O(gate161inter3));
  inv1  gate1769(.a(s_175), .O(gate161inter4));
  nand2 gate1770(.a(gate161inter4), .b(gate161inter3), .O(gate161inter5));
  nor2  gate1771(.a(gate161inter5), .b(gate161inter2), .O(gate161inter6));
  inv1  gate1772(.a(G450), .O(gate161inter7));
  inv1  gate1773(.a(G534), .O(gate161inter8));
  nand2 gate1774(.a(gate161inter8), .b(gate161inter7), .O(gate161inter9));
  nand2 gate1775(.a(s_175), .b(gate161inter3), .O(gate161inter10));
  nor2  gate1776(.a(gate161inter10), .b(gate161inter9), .O(gate161inter11));
  nor2  gate1777(.a(gate161inter11), .b(gate161inter6), .O(gate161inter12));
  nand2 gate1778(.a(gate161inter12), .b(gate161inter1), .O(G578));

  xor2  gate1373(.a(G534), .b(G453), .O(gate162inter0));
  nand2 gate1374(.a(gate162inter0), .b(s_118), .O(gate162inter1));
  and2  gate1375(.a(G534), .b(G453), .O(gate162inter2));
  inv1  gate1376(.a(s_118), .O(gate162inter3));
  inv1  gate1377(.a(s_119), .O(gate162inter4));
  nand2 gate1378(.a(gate162inter4), .b(gate162inter3), .O(gate162inter5));
  nor2  gate1379(.a(gate162inter5), .b(gate162inter2), .O(gate162inter6));
  inv1  gate1380(.a(G453), .O(gate162inter7));
  inv1  gate1381(.a(G534), .O(gate162inter8));
  nand2 gate1382(.a(gate162inter8), .b(gate162inter7), .O(gate162inter9));
  nand2 gate1383(.a(s_119), .b(gate162inter3), .O(gate162inter10));
  nor2  gate1384(.a(gate162inter10), .b(gate162inter9), .O(gate162inter11));
  nor2  gate1385(.a(gate162inter11), .b(gate162inter6), .O(gate162inter12));
  nand2 gate1386(.a(gate162inter12), .b(gate162inter1), .O(G579));
nand2 gate163( .a(G456), .b(G537), .O(G580) );
nand2 gate164( .a(G459), .b(G537), .O(G581) );

  xor2  gate1681(.a(G540), .b(G462), .O(gate165inter0));
  nand2 gate1682(.a(gate165inter0), .b(s_162), .O(gate165inter1));
  and2  gate1683(.a(G540), .b(G462), .O(gate165inter2));
  inv1  gate1684(.a(s_162), .O(gate165inter3));
  inv1  gate1685(.a(s_163), .O(gate165inter4));
  nand2 gate1686(.a(gate165inter4), .b(gate165inter3), .O(gate165inter5));
  nor2  gate1687(.a(gate165inter5), .b(gate165inter2), .O(gate165inter6));
  inv1  gate1688(.a(G462), .O(gate165inter7));
  inv1  gate1689(.a(G540), .O(gate165inter8));
  nand2 gate1690(.a(gate165inter8), .b(gate165inter7), .O(gate165inter9));
  nand2 gate1691(.a(s_163), .b(gate165inter3), .O(gate165inter10));
  nor2  gate1692(.a(gate165inter10), .b(gate165inter9), .O(gate165inter11));
  nor2  gate1693(.a(gate165inter11), .b(gate165inter6), .O(gate165inter12));
  nand2 gate1694(.a(gate165inter12), .b(gate165inter1), .O(G582));

  xor2  gate1751(.a(G540), .b(G465), .O(gate166inter0));
  nand2 gate1752(.a(gate166inter0), .b(s_172), .O(gate166inter1));
  and2  gate1753(.a(G540), .b(G465), .O(gate166inter2));
  inv1  gate1754(.a(s_172), .O(gate166inter3));
  inv1  gate1755(.a(s_173), .O(gate166inter4));
  nand2 gate1756(.a(gate166inter4), .b(gate166inter3), .O(gate166inter5));
  nor2  gate1757(.a(gate166inter5), .b(gate166inter2), .O(gate166inter6));
  inv1  gate1758(.a(G465), .O(gate166inter7));
  inv1  gate1759(.a(G540), .O(gate166inter8));
  nand2 gate1760(.a(gate166inter8), .b(gate166inter7), .O(gate166inter9));
  nand2 gate1761(.a(s_173), .b(gate166inter3), .O(gate166inter10));
  nor2  gate1762(.a(gate166inter10), .b(gate166inter9), .O(gate166inter11));
  nor2  gate1763(.a(gate166inter11), .b(gate166inter6), .O(gate166inter12));
  nand2 gate1764(.a(gate166inter12), .b(gate166inter1), .O(G583));
nand2 gate167( .a(G468), .b(G543), .O(G584) );
nand2 gate168( .a(G471), .b(G543), .O(G585) );

  xor2  gate813(.a(G546), .b(G474), .O(gate169inter0));
  nand2 gate814(.a(gate169inter0), .b(s_38), .O(gate169inter1));
  and2  gate815(.a(G546), .b(G474), .O(gate169inter2));
  inv1  gate816(.a(s_38), .O(gate169inter3));
  inv1  gate817(.a(s_39), .O(gate169inter4));
  nand2 gate818(.a(gate169inter4), .b(gate169inter3), .O(gate169inter5));
  nor2  gate819(.a(gate169inter5), .b(gate169inter2), .O(gate169inter6));
  inv1  gate820(.a(G474), .O(gate169inter7));
  inv1  gate821(.a(G546), .O(gate169inter8));
  nand2 gate822(.a(gate169inter8), .b(gate169inter7), .O(gate169inter9));
  nand2 gate823(.a(s_39), .b(gate169inter3), .O(gate169inter10));
  nor2  gate824(.a(gate169inter10), .b(gate169inter9), .O(gate169inter11));
  nor2  gate825(.a(gate169inter11), .b(gate169inter6), .O(gate169inter12));
  nand2 gate826(.a(gate169inter12), .b(gate169inter1), .O(G586));

  xor2  gate2241(.a(G546), .b(G477), .O(gate170inter0));
  nand2 gate2242(.a(gate170inter0), .b(s_242), .O(gate170inter1));
  and2  gate2243(.a(G546), .b(G477), .O(gate170inter2));
  inv1  gate2244(.a(s_242), .O(gate170inter3));
  inv1  gate2245(.a(s_243), .O(gate170inter4));
  nand2 gate2246(.a(gate170inter4), .b(gate170inter3), .O(gate170inter5));
  nor2  gate2247(.a(gate170inter5), .b(gate170inter2), .O(gate170inter6));
  inv1  gate2248(.a(G477), .O(gate170inter7));
  inv1  gate2249(.a(G546), .O(gate170inter8));
  nand2 gate2250(.a(gate170inter8), .b(gate170inter7), .O(gate170inter9));
  nand2 gate2251(.a(s_243), .b(gate170inter3), .O(gate170inter10));
  nor2  gate2252(.a(gate170inter10), .b(gate170inter9), .O(gate170inter11));
  nor2  gate2253(.a(gate170inter11), .b(gate170inter6), .O(gate170inter12));
  nand2 gate2254(.a(gate170inter12), .b(gate170inter1), .O(G587));

  xor2  gate2339(.a(G549), .b(G480), .O(gate171inter0));
  nand2 gate2340(.a(gate171inter0), .b(s_256), .O(gate171inter1));
  and2  gate2341(.a(G549), .b(G480), .O(gate171inter2));
  inv1  gate2342(.a(s_256), .O(gate171inter3));
  inv1  gate2343(.a(s_257), .O(gate171inter4));
  nand2 gate2344(.a(gate171inter4), .b(gate171inter3), .O(gate171inter5));
  nor2  gate2345(.a(gate171inter5), .b(gate171inter2), .O(gate171inter6));
  inv1  gate2346(.a(G480), .O(gate171inter7));
  inv1  gate2347(.a(G549), .O(gate171inter8));
  nand2 gate2348(.a(gate171inter8), .b(gate171inter7), .O(gate171inter9));
  nand2 gate2349(.a(s_257), .b(gate171inter3), .O(gate171inter10));
  nor2  gate2350(.a(gate171inter10), .b(gate171inter9), .O(gate171inter11));
  nor2  gate2351(.a(gate171inter11), .b(gate171inter6), .O(gate171inter12));
  nand2 gate2352(.a(gate171inter12), .b(gate171inter1), .O(G588));
nand2 gate172( .a(G483), .b(G549), .O(G589) );
nand2 gate173( .a(G486), .b(G552), .O(G590) );

  xor2  gate2885(.a(G552), .b(G489), .O(gate174inter0));
  nand2 gate2886(.a(gate174inter0), .b(s_334), .O(gate174inter1));
  and2  gate2887(.a(G552), .b(G489), .O(gate174inter2));
  inv1  gate2888(.a(s_334), .O(gate174inter3));
  inv1  gate2889(.a(s_335), .O(gate174inter4));
  nand2 gate2890(.a(gate174inter4), .b(gate174inter3), .O(gate174inter5));
  nor2  gate2891(.a(gate174inter5), .b(gate174inter2), .O(gate174inter6));
  inv1  gate2892(.a(G489), .O(gate174inter7));
  inv1  gate2893(.a(G552), .O(gate174inter8));
  nand2 gate2894(.a(gate174inter8), .b(gate174inter7), .O(gate174inter9));
  nand2 gate2895(.a(s_335), .b(gate174inter3), .O(gate174inter10));
  nor2  gate2896(.a(gate174inter10), .b(gate174inter9), .O(gate174inter11));
  nor2  gate2897(.a(gate174inter11), .b(gate174inter6), .O(gate174inter12));
  nand2 gate2898(.a(gate174inter12), .b(gate174inter1), .O(G591));

  xor2  gate2325(.a(G555), .b(G492), .O(gate175inter0));
  nand2 gate2326(.a(gate175inter0), .b(s_254), .O(gate175inter1));
  and2  gate2327(.a(G555), .b(G492), .O(gate175inter2));
  inv1  gate2328(.a(s_254), .O(gate175inter3));
  inv1  gate2329(.a(s_255), .O(gate175inter4));
  nand2 gate2330(.a(gate175inter4), .b(gate175inter3), .O(gate175inter5));
  nor2  gate2331(.a(gate175inter5), .b(gate175inter2), .O(gate175inter6));
  inv1  gate2332(.a(G492), .O(gate175inter7));
  inv1  gate2333(.a(G555), .O(gate175inter8));
  nand2 gate2334(.a(gate175inter8), .b(gate175inter7), .O(gate175inter9));
  nand2 gate2335(.a(s_255), .b(gate175inter3), .O(gate175inter10));
  nor2  gate2336(.a(gate175inter10), .b(gate175inter9), .O(gate175inter11));
  nor2  gate2337(.a(gate175inter11), .b(gate175inter6), .O(gate175inter12));
  nand2 gate2338(.a(gate175inter12), .b(gate175inter1), .O(G592));

  xor2  gate2661(.a(G555), .b(G495), .O(gate176inter0));
  nand2 gate2662(.a(gate176inter0), .b(s_302), .O(gate176inter1));
  and2  gate2663(.a(G555), .b(G495), .O(gate176inter2));
  inv1  gate2664(.a(s_302), .O(gate176inter3));
  inv1  gate2665(.a(s_303), .O(gate176inter4));
  nand2 gate2666(.a(gate176inter4), .b(gate176inter3), .O(gate176inter5));
  nor2  gate2667(.a(gate176inter5), .b(gate176inter2), .O(gate176inter6));
  inv1  gate2668(.a(G495), .O(gate176inter7));
  inv1  gate2669(.a(G555), .O(gate176inter8));
  nand2 gate2670(.a(gate176inter8), .b(gate176inter7), .O(gate176inter9));
  nand2 gate2671(.a(s_303), .b(gate176inter3), .O(gate176inter10));
  nor2  gate2672(.a(gate176inter10), .b(gate176inter9), .O(gate176inter11));
  nor2  gate2673(.a(gate176inter11), .b(gate176inter6), .O(gate176inter12));
  nand2 gate2674(.a(gate176inter12), .b(gate176inter1), .O(G593));
nand2 gate177( .a(G498), .b(G558), .O(G594) );

  xor2  gate1611(.a(G558), .b(G501), .O(gate178inter0));
  nand2 gate1612(.a(gate178inter0), .b(s_152), .O(gate178inter1));
  and2  gate1613(.a(G558), .b(G501), .O(gate178inter2));
  inv1  gate1614(.a(s_152), .O(gate178inter3));
  inv1  gate1615(.a(s_153), .O(gate178inter4));
  nand2 gate1616(.a(gate178inter4), .b(gate178inter3), .O(gate178inter5));
  nor2  gate1617(.a(gate178inter5), .b(gate178inter2), .O(gate178inter6));
  inv1  gate1618(.a(G501), .O(gate178inter7));
  inv1  gate1619(.a(G558), .O(gate178inter8));
  nand2 gate1620(.a(gate178inter8), .b(gate178inter7), .O(gate178inter9));
  nand2 gate1621(.a(s_153), .b(gate178inter3), .O(gate178inter10));
  nor2  gate1622(.a(gate178inter10), .b(gate178inter9), .O(gate178inter11));
  nor2  gate1623(.a(gate178inter11), .b(gate178inter6), .O(gate178inter12));
  nand2 gate1624(.a(gate178inter12), .b(gate178inter1), .O(G595));

  xor2  gate1597(.a(G561), .b(G504), .O(gate179inter0));
  nand2 gate1598(.a(gate179inter0), .b(s_150), .O(gate179inter1));
  and2  gate1599(.a(G561), .b(G504), .O(gate179inter2));
  inv1  gate1600(.a(s_150), .O(gate179inter3));
  inv1  gate1601(.a(s_151), .O(gate179inter4));
  nand2 gate1602(.a(gate179inter4), .b(gate179inter3), .O(gate179inter5));
  nor2  gate1603(.a(gate179inter5), .b(gate179inter2), .O(gate179inter6));
  inv1  gate1604(.a(G504), .O(gate179inter7));
  inv1  gate1605(.a(G561), .O(gate179inter8));
  nand2 gate1606(.a(gate179inter8), .b(gate179inter7), .O(gate179inter9));
  nand2 gate1607(.a(s_151), .b(gate179inter3), .O(gate179inter10));
  nor2  gate1608(.a(gate179inter10), .b(gate179inter9), .O(gate179inter11));
  nor2  gate1609(.a(gate179inter11), .b(gate179inter6), .O(gate179inter12));
  nand2 gate1610(.a(gate179inter12), .b(gate179inter1), .O(G596));

  xor2  gate617(.a(G561), .b(G507), .O(gate180inter0));
  nand2 gate618(.a(gate180inter0), .b(s_10), .O(gate180inter1));
  and2  gate619(.a(G561), .b(G507), .O(gate180inter2));
  inv1  gate620(.a(s_10), .O(gate180inter3));
  inv1  gate621(.a(s_11), .O(gate180inter4));
  nand2 gate622(.a(gate180inter4), .b(gate180inter3), .O(gate180inter5));
  nor2  gate623(.a(gate180inter5), .b(gate180inter2), .O(gate180inter6));
  inv1  gate624(.a(G507), .O(gate180inter7));
  inv1  gate625(.a(G561), .O(gate180inter8));
  nand2 gate626(.a(gate180inter8), .b(gate180inter7), .O(gate180inter9));
  nand2 gate627(.a(s_11), .b(gate180inter3), .O(gate180inter10));
  nor2  gate628(.a(gate180inter10), .b(gate180inter9), .O(gate180inter11));
  nor2  gate629(.a(gate180inter11), .b(gate180inter6), .O(gate180inter12));
  nand2 gate630(.a(gate180inter12), .b(gate180inter1), .O(G597));
nand2 gate181( .a(G510), .b(G564), .O(G598) );
nand2 gate182( .a(G513), .b(G564), .O(G599) );
nand2 gate183( .a(G516), .b(G567), .O(G600) );
nand2 gate184( .a(G519), .b(G567), .O(G601) );

  xor2  gate2969(.a(G571), .b(G570), .O(gate185inter0));
  nand2 gate2970(.a(gate185inter0), .b(s_346), .O(gate185inter1));
  and2  gate2971(.a(G571), .b(G570), .O(gate185inter2));
  inv1  gate2972(.a(s_346), .O(gate185inter3));
  inv1  gate2973(.a(s_347), .O(gate185inter4));
  nand2 gate2974(.a(gate185inter4), .b(gate185inter3), .O(gate185inter5));
  nor2  gate2975(.a(gate185inter5), .b(gate185inter2), .O(gate185inter6));
  inv1  gate2976(.a(G570), .O(gate185inter7));
  inv1  gate2977(.a(G571), .O(gate185inter8));
  nand2 gate2978(.a(gate185inter8), .b(gate185inter7), .O(gate185inter9));
  nand2 gate2979(.a(s_347), .b(gate185inter3), .O(gate185inter10));
  nor2  gate2980(.a(gate185inter10), .b(gate185inter9), .O(gate185inter11));
  nor2  gate2981(.a(gate185inter11), .b(gate185inter6), .O(gate185inter12));
  nand2 gate2982(.a(gate185inter12), .b(gate185inter1), .O(G602));
nand2 gate186( .a(G572), .b(G573), .O(G607) );
nand2 gate187( .a(G574), .b(G575), .O(G612) );
nand2 gate188( .a(G576), .b(G577), .O(G617) );
nand2 gate189( .a(G578), .b(G579), .O(G622) );

  xor2  gate2017(.a(G581), .b(G580), .O(gate190inter0));
  nand2 gate2018(.a(gate190inter0), .b(s_210), .O(gate190inter1));
  and2  gate2019(.a(G581), .b(G580), .O(gate190inter2));
  inv1  gate2020(.a(s_210), .O(gate190inter3));
  inv1  gate2021(.a(s_211), .O(gate190inter4));
  nand2 gate2022(.a(gate190inter4), .b(gate190inter3), .O(gate190inter5));
  nor2  gate2023(.a(gate190inter5), .b(gate190inter2), .O(gate190inter6));
  inv1  gate2024(.a(G580), .O(gate190inter7));
  inv1  gate2025(.a(G581), .O(gate190inter8));
  nand2 gate2026(.a(gate190inter8), .b(gate190inter7), .O(gate190inter9));
  nand2 gate2027(.a(s_211), .b(gate190inter3), .O(gate190inter10));
  nor2  gate2028(.a(gate190inter10), .b(gate190inter9), .O(gate190inter11));
  nor2  gate2029(.a(gate190inter11), .b(gate190inter6), .O(gate190inter12));
  nand2 gate2030(.a(gate190inter12), .b(gate190inter1), .O(G627));
nand2 gate191( .a(G582), .b(G583), .O(G632) );
nand2 gate192( .a(G584), .b(G585), .O(G637) );

  xor2  gate2451(.a(G587), .b(G586), .O(gate193inter0));
  nand2 gate2452(.a(gate193inter0), .b(s_272), .O(gate193inter1));
  and2  gate2453(.a(G587), .b(G586), .O(gate193inter2));
  inv1  gate2454(.a(s_272), .O(gate193inter3));
  inv1  gate2455(.a(s_273), .O(gate193inter4));
  nand2 gate2456(.a(gate193inter4), .b(gate193inter3), .O(gate193inter5));
  nor2  gate2457(.a(gate193inter5), .b(gate193inter2), .O(gate193inter6));
  inv1  gate2458(.a(G586), .O(gate193inter7));
  inv1  gate2459(.a(G587), .O(gate193inter8));
  nand2 gate2460(.a(gate193inter8), .b(gate193inter7), .O(gate193inter9));
  nand2 gate2461(.a(s_273), .b(gate193inter3), .O(gate193inter10));
  nor2  gate2462(.a(gate193inter10), .b(gate193inter9), .O(gate193inter11));
  nor2  gate2463(.a(gate193inter11), .b(gate193inter6), .O(gate193inter12));
  nand2 gate2464(.a(gate193inter12), .b(gate193inter1), .O(G642));
nand2 gate194( .a(G588), .b(G589), .O(G645) );
nand2 gate195( .a(G590), .b(G591), .O(G648) );
nand2 gate196( .a(G592), .b(G593), .O(G651) );
nand2 gate197( .a(G594), .b(G595), .O(G654) );

  xor2  gate645(.a(G597), .b(G596), .O(gate198inter0));
  nand2 gate646(.a(gate198inter0), .b(s_14), .O(gate198inter1));
  and2  gate647(.a(G597), .b(G596), .O(gate198inter2));
  inv1  gate648(.a(s_14), .O(gate198inter3));
  inv1  gate649(.a(s_15), .O(gate198inter4));
  nand2 gate650(.a(gate198inter4), .b(gate198inter3), .O(gate198inter5));
  nor2  gate651(.a(gate198inter5), .b(gate198inter2), .O(gate198inter6));
  inv1  gate652(.a(G596), .O(gate198inter7));
  inv1  gate653(.a(G597), .O(gate198inter8));
  nand2 gate654(.a(gate198inter8), .b(gate198inter7), .O(gate198inter9));
  nand2 gate655(.a(s_15), .b(gate198inter3), .O(gate198inter10));
  nor2  gate656(.a(gate198inter10), .b(gate198inter9), .O(gate198inter11));
  nor2  gate657(.a(gate198inter11), .b(gate198inter6), .O(gate198inter12));
  nand2 gate658(.a(gate198inter12), .b(gate198inter1), .O(G657));
nand2 gate199( .a(G598), .b(G599), .O(G660) );
nand2 gate200( .a(G600), .b(G601), .O(G663) );

  xor2  gate2857(.a(G607), .b(G602), .O(gate201inter0));
  nand2 gate2858(.a(gate201inter0), .b(s_330), .O(gate201inter1));
  and2  gate2859(.a(G607), .b(G602), .O(gate201inter2));
  inv1  gate2860(.a(s_330), .O(gate201inter3));
  inv1  gate2861(.a(s_331), .O(gate201inter4));
  nand2 gate2862(.a(gate201inter4), .b(gate201inter3), .O(gate201inter5));
  nor2  gate2863(.a(gate201inter5), .b(gate201inter2), .O(gate201inter6));
  inv1  gate2864(.a(G602), .O(gate201inter7));
  inv1  gate2865(.a(G607), .O(gate201inter8));
  nand2 gate2866(.a(gate201inter8), .b(gate201inter7), .O(gate201inter9));
  nand2 gate2867(.a(s_331), .b(gate201inter3), .O(gate201inter10));
  nor2  gate2868(.a(gate201inter10), .b(gate201inter9), .O(gate201inter11));
  nor2  gate2869(.a(gate201inter11), .b(gate201inter6), .O(gate201inter12));
  nand2 gate2870(.a(gate201inter12), .b(gate201inter1), .O(G666));

  xor2  gate1247(.a(G617), .b(G612), .O(gate202inter0));
  nand2 gate1248(.a(gate202inter0), .b(s_100), .O(gate202inter1));
  and2  gate1249(.a(G617), .b(G612), .O(gate202inter2));
  inv1  gate1250(.a(s_100), .O(gate202inter3));
  inv1  gate1251(.a(s_101), .O(gate202inter4));
  nand2 gate1252(.a(gate202inter4), .b(gate202inter3), .O(gate202inter5));
  nor2  gate1253(.a(gate202inter5), .b(gate202inter2), .O(gate202inter6));
  inv1  gate1254(.a(G612), .O(gate202inter7));
  inv1  gate1255(.a(G617), .O(gate202inter8));
  nand2 gate1256(.a(gate202inter8), .b(gate202inter7), .O(gate202inter9));
  nand2 gate1257(.a(s_101), .b(gate202inter3), .O(gate202inter10));
  nor2  gate1258(.a(gate202inter10), .b(gate202inter9), .O(gate202inter11));
  nor2  gate1259(.a(gate202inter11), .b(gate202inter6), .O(gate202inter12));
  nand2 gate1260(.a(gate202inter12), .b(gate202inter1), .O(G669));
nand2 gate203( .a(G602), .b(G612), .O(G672) );
nand2 gate204( .a(G607), .b(G617), .O(G675) );

  xor2  gate2535(.a(G627), .b(G622), .O(gate205inter0));
  nand2 gate2536(.a(gate205inter0), .b(s_284), .O(gate205inter1));
  and2  gate2537(.a(G627), .b(G622), .O(gate205inter2));
  inv1  gate2538(.a(s_284), .O(gate205inter3));
  inv1  gate2539(.a(s_285), .O(gate205inter4));
  nand2 gate2540(.a(gate205inter4), .b(gate205inter3), .O(gate205inter5));
  nor2  gate2541(.a(gate205inter5), .b(gate205inter2), .O(gate205inter6));
  inv1  gate2542(.a(G622), .O(gate205inter7));
  inv1  gate2543(.a(G627), .O(gate205inter8));
  nand2 gate2544(.a(gate205inter8), .b(gate205inter7), .O(gate205inter9));
  nand2 gate2545(.a(s_285), .b(gate205inter3), .O(gate205inter10));
  nor2  gate2546(.a(gate205inter10), .b(gate205inter9), .O(gate205inter11));
  nor2  gate2547(.a(gate205inter11), .b(gate205inter6), .O(gate205inter12));
  nand2 gate2548(.a(gate205inter12), .b(gate205inter1), .O(G678));
nand2 gate206( .a(G632), .b(G637), .O(G681) );

  xor2  gate1079(.a(G632), .b(G622), .O(gate207inter0));
  nand2 gate1080(.a(gate207inter0), .b(s_76), .O(gate207inter1));
  and2  gate1081(.a(G632), .b(G622), .O(gate207inter2));
  inv1  gate1082(.a(s_76), .O(gate207inter3));
  inv1  gate1083(.a(s_77), .O(gate207inter4));
  nand2 gate1084(.a(gate207inter4), .b(gate207inter3), .O(gate207inter5));
  nor2  gate1085(.a(gate207inter5), .b(gate207inter2), .O(gate207inter6));
  inv1  gate1086(.a(G622), .O(gate207inter7));
  inv1  gate1087(.a(G632), .O(gate207inter8));
  nand2 gate1088(.a(gate207inter8), .b(gate207inter7), .O(gate207inter9));
  nand2 gate1089(.a(s_77), .b(gate207inter3), .O(gate207inter10));
  nor2  gate1090(.a(gate207inter10), .b(gate207inter9), .O(gate207inter11));
  nor2  gate1091(.a(gate207inter11), .b(gate207inter6), .O(gate207inter12));
  nand2 gate1092(.a(gate207inter12), .b(gate207inter1), .O(G684));
nand2 gate208( .a(G627), .b(G637), .O(G687) );

  xor2  gate925(.a(G666), .b(G602), .O(gate209inter0));
  nand2 gate926(.a(gate209inter0), .b(s_54), .O(gate209inter1));
  and2  gate927(.a(G666), .b(G602), .O(gate209inter2));
  inv1  gate928(.a(s_54), .O(gate209inter3));
  inv1  gate929(.a(s_55), .O(gate209inter4));
  nand2 gate930(.a(gate209inter4), .b(gate209inter3), .O(gate209inter5));
  nor2  gate931(.a(gate209inter5), .b(gate209inter2), .O(gate209inter6));
  inv1  gate932(.a(G602), .O(gate209inter7));
  inv1  gate933(.a(G666), .O(gate209inter8));
  nand2 gate934(.a(gate209inter8), .b(gate209inter7), .O(gate209inter9));
  nand2 gate935(.a(s_55), .b(gate209inter3), .O(gate209inter10));
  nor2  gate936(.a(gate209inter10), .b(gate209inter9), .O(gate209inter11));
  nor2  gate937(.a(gate209inter11), .b(gate209inter6), .O(gate209inter12));
  nand2 gate938(.a(gate209inter12), .b(gate209inter1), .O(G690));

  xor2  gate2129(.a(G666), .b(G607), .O(gate210inter0));
  nand2 gate2130(.a(gate210inter0), .b(s_226), .O(gate210inter1));
  and2  gate2131(.a(G666), .b(G607), .O(gate210inter2));
  inv1  gate2132(.a(s_226), .O(gate210inter3));
  inv1  gate2133(.a(s_227), .O(gate210inter4));
  nand2 gate2134(.a(gate210inter4), .b(gate210inter3), .O(gate210inter5));
  nor2  gate2135(.a(gate210inter5), .b(gate210inter2), .O(gate210inter6));
  inv1  gate2136(.a(G607), .O(gate210inter7));
  inv1  gate2137(.a(G666), .O(gate210inter8));
  nand2 gate2138(.a(gate210inter8), .b(gate210inter7), .O(gate210inter9));
  nand2 gate2139(.a(s_227), .b(gate210inter3), .O(gate210inter10));
  nor2  gate2140(.a(gate210inter10), .b(gate210inter9), .O(gate210inter11));
  nor2  gate2141(.a(gate210inter11), .b(gate210inter6), .O(gate210inter12));
  nand2 gate2142(.a(gate210inter12), .b(gate210inter1), .O(G691));
nand2 gate211( .a(G612), .b(G669), .O(G692) );

  xor2  gate2493(.a(G669), .b(G617), .O(gate212inter0));
  nand2 gate2494(.a(gate212inter0), .b(s_278), .O(gate212inter1));
  and2  gate2495(.a(G669), .b(G617), .O(gate212inter2));
  inv1  gate2496(.a(s_278), .O(gate212inter3));
  inv1  gate2497(.a(s_279), .O(gate212inter4));
  nand2 gate2498(.a(gate212inter4), .b(gate212inter3), .O(gate212inter5));
  nor2  gate2499(.a(gate212inter5), .b(gate212inter2), .O(gate212inter6));
  inv1  gate2500(.a(G617), .O(gate212inter7));
  inv1  gate2501(.a(G669), .O(gate212inter8));
  nand2 gate2502(.a(gate212inter8), .b(gate212inter7), .O(gate212inter9));
  nand2 gate2503(.a(s_279), .b(gate212inter3), .O(gate212inter10));
  nor2  gate2504(.a(gate212inter10), .b(gate212inter9), .O(gate212inter11));
  nor2  gate2505(.a(gate212inter11), .b(gate212inter6), .O(gate212inter12));
  nand2 gate2506(.a(gate212inter12), .b(gate212inter1), .O(G693));
nand2 gate213( .a(G602), .b(G672), .O(G694) );
nand2 gate214( .a(G612), .b(G672), .O(G695) );
nand2 gate215( .a(G607), .b(G675), .O(G696) );

  xor2  gate2703(.a(G675), .b(G617), .O(gate216inter0));
  nand2 gate2704(.a(gate216inter0), .b(s_308), .O(gate216inter1));
  and2  gate2705(.a(G675), .b(G617), .O(gate216inter2));
  inv1  gate2706(.a(s_308), .O(gate216inter3));
  inv1  gate2707(.a(s_309), .O(gate216inter4));
  nand2 gate2708(.a(gate216inter4), .b(gate216inter3), .O(gate216inter5));
  nor2  gate2709(.a(gate216inter5), .b(gate216inter2), .O(gate216inter6));
  inv1  gate2710(.a(G617), .O(gate216inter7));
  inv1  gate2711(.a(G675), .O(gate216inter8));
  nand2 gate2712(.a(gate216inter8), .b(gate216inter7), .O(gate216inter9));
  nand2 gate2713(.a(s_309), .b(gate216inter3), .O(gate216inter10));
  nor2  gate2714(.a(gate216inter10), .b(gate216inter9), .O(gate216inter11));
  nor2  gate2715(.a(gate216inter11), .b(gate216inter6), .O(gate216inter12));
  nand2 gate2716(.a(gate216inter12), .b(gate216inter1), .O(G697));

  xor2  gate2101(.a(G678), .b(G622), .O(gate217inter0));
  nand2 gate2102(.a(gate217inter0), .b(s_222), .O(gate217inter1));
  and2  gate2103(.a(G678), .b(G622), .O(gate217inter2));
  inv1  gate2104(.a(s_222), .O(gate217inter3));
  inv1  gate2105(.a(s_223), .O(gate217inter4));
  nand2 gate2106(.a(gate217inter4), .b(gate217inter3), .O(gate217inter5));
  nor2  gate2107(.a(gate217inter5), .b(gate217inter2), .O(gate217inter6));
  inv1  gate2108(.a(G622), .O(gate217inter7));
  inv1  gate2109(.a(G678), .O(gate217inter8));
  nand2 gate2110(.a(gate217inter8), .b(gate217inter7), .O(gate217inter9));
  nand2 gate2111(.a(s_223), .b(gate217inter3), .O(gate217inter10));
  nor2  gate2112(.a(gate217inter10), .b(gate217inter9), .O(gate217inter11));
  nor2  gate2113(.a(gate217inter11), .b(gate217inter6), .O(gate217inter12));
  nand2 gate2114(.a(gate217inter12), .b(gate217inter1), .O(G698));

  xor2  gate2409(.a(G678), .b(G627), .O(gate218inter0));
  nand2 gate2410(.a(gate218inter0), .b(s_266), .O(gate218inter1));
  and2  gate2411(.a(G678), .b(G627), .O(gate218inter2));
  inv1  gate2412(.a(s_266), .O(gate218inter3));
  inv1  gate2413(.a(s_267), .O(gate218inter4));
  nand2 gate2414(.a(gate218inter4), .b(gate218inter3), .O(gate218inter5));
  nor2  gate2415(.a(gate218inter5), .b(gate218inter2), .O(gate218inter6));
  inv1  gate2416(.a(G627), .O(gate218inter7));
  inv1  gate2417(.a(G678), .O(gate218inter8));
  nand2 gate2418(.a(gate218inter8), .b(gate218inter7), .O(gate218inter9));
  nand2 gate2419(.a(s_267), .b(gate218inter3), .O(gate218inter10));
  nor2  gate2420(.a(gate218inter10), .b(gate218inter9), .O(gate218inter11));
  nor2  gate2421(.a(gate218inter11), .b(gate218inter6), .O(gate218inter12));
  nand2 gate2422(.a(gate218inter12), .b(gate218inter1), .O(G699));

  xor2  gate2829(.a(G681), .b(G632), .O(gate219inter0));
  nand2 gate2830(.a(gate219inter0), .b(s_326), .O(gate219inter1));
  and2  gate2831(.a(G681), .b(G632), .O(gate219inter2));
  inv1  gate2832(.a(s_326), .O(gate219inter3));
  inv1  gate2833(.a(s_327), .O(gate219inter4));
  nand2 gate2834(.a(gate219inter4), .b(gate219inter3), .O(gate219inter5));
  nor2  gate2835(.a(gate219inter5), .b(gate219inter2), .O(gate219inter6));
  inv1  gate2836(.a(G632), .O(gate219inter7));
  inv1  gate2837(.a(G681), .O(gate219inter8));
  nand2 gate2838(.a(gate219inter8), .b(gate219inter7), .O(gate219inter9));
  nand2 gate2839(.a(s_327), .b(gate219inter3), .O(gate219inter10));
  nor2  gate2840(.a(gate219inter10), .b(gate219inter9), .O(gate219inter11));
  nor2  gate2841(.a(gate219inter11), .b(gate219inter6), .O(gate219inter12));
  nand2 gate2842(.a(gate219inter12), .b(gate219inter1), .O(G700));
nand2 gate220( .a(G637), .b(G681), .O(G701) );

  xor2  gate715(.a(G684), .b(G622), .O(gate221inter0));
  nand2 gate716(.a(gate221inter0), .b(s_24), .O(gate221inter1));
  and2  gate717(.a(G684), .b(G622), .O(gate221inter2));
  inv1  gate718(.a(s_24), .O(gate221inter3));
  inv1  gate719(.a(s_25), .O(gate221inter4));
  nand2 gate720(.a(gate221inter4), .b(gate221inter3), .O(gate221inter5));
  nor2  gate721(.a(gate221inter5), .b(gate221inter2), .O(gate221inter6));
  inv1  gate722(.a(G622), .O(gate221inter7));
  inv1  gate723(.a(G684), .O(gate221inter8));
  nand2 gate724(.a(gate221inter8), .b(gate221inter7), .O(gate221inter9));
  nand2 gate725(.a(s_25), .b(gate221inter3), .O(gate221inter10));
  nor2  gate726(.a(gate221inter10), .b(gate221inter9), .O(gate221inter11));
  nor2  gate727(.a(gate221inter11), .b(gate221inter6), .O(gate221inter12));
  nand2 gate728(.a(gate221inter12), .b(gate221inter1), .O(G702));

  xor2  gate2787(.a(G684), .b(G632), .O(gate222inter0));
  nand2 gate2788(.a(gate222inter0), .b(s_320), .O(gate222inter1));
  and2  gate2789(.a(G684), .b(G632), .O(gate222inter2));
  inv1  gate2790(.a(s_320), .O(gate222inter3));
  inv1  gate2791(.a(s_321), .O(gate222inter4));
  nand2 gate2792(.a(gate222inter4), .b(gate222inter3), .O(gate222inter5));
  nor2  gate2793(.a(gate222inter5), .b(gate222inter2), .O(gate222inter6));
  inv1  gate2794(.a(G632), .O(gate222inter7));
  inv1  gate2795(.a(G684), .O(gate222inter8));
  nand2 gate2796(.a(gate222inter8), .b(gate222inter7), .O(gate222inter9));
  nand2 gate2797(.a(s_321), .b(gate222inter3), .O(gate222inter10));
  nor2  gate2798(.a(gate222inter10), .b(gate222inter9), .O(gate222inter11));
  nor2  gate2799(.a(gate222inter11), .b(gate222inter6), .O(gate222inter12));
  nand2 gate2800(.a(gate222inter12), .b(gate222inter1), .O(G703));
nand2 gate223( .a(G627), .b(G687), .O(G704) );

  xor2  gate1303(.a(G687), .b(G637), .O(gate224inter0));
  nand2 gate1304(.a(gate224inter0), .b(s_108), .O(gate224inter1));
  and2  gate1305(.a(G687), .b(G637), .O(gate224inter2));
  inv1  gate1306(.a(s_108), .O(gate224inter3));
  inv1  gate1307(.a(s_109), .O(gate224inter4));
  nand2 gate1308(.a(gate224inter4), .b(gate224inter3), .O(gate224inter5));
  nor2  gate1309(.a(gate224inter5), .b(gate224inter2), .O(gate224inter6));
  inv1  gate1310(.a(G637), .O(gate224inter7));
  inv1  gate1311(.a(G687), .O(gate224inter8));
  nand2 gate1312(.a(gate224inter8), .b(gate224inter7), .O(gate224inter9));
  nand2 gate1313(.a(s_109), .b(gate224inter3), .O(gate224inter10));
  nor2  gate1314(.a(gate224inter10), .b(gate224inter9), .O(gate224inter11));
  nor2  gate1315(.a(gate224inter11), .b(gate224inter6), .O(gate224inter12));
  nand2 gate1316(.a(gate224inter12), .b(gate224inter1), .O(G705));

  xor2  gate575(.a(G691), .b(G690), .O(gate225inter0));
  nand2 gate576(.a(gate225inter0), .b(s_4), .O(gate225inter1));
  and2  gate577(.a(G691), .b(G690), .O(gate225inter2));
  inv1  gate578(.a(s_4), .O(gate225inter3));
  inv1  gate579(.a(s_5), .O(gate225inter4));
  nand2 gate580(.a(gate225inter4), .b(gate225inter3), .O(gate225inter5));
  nor2  gate581(.a(gate225inter5), .b(gate225inter2), .O(gate225inter6));
  inv1  gate582(.a(G690), .O(gate225inter7));
  inv1  gate583(.a(G691), .O(gate225inter8));
  nand2 gate584(.a(gate225inter8), .b(gate225inter7), .O(gate225inter9));
  nand2 gate585(.a(s_5), .b(gate225inter3), .O(gate225inter10));
  nor2  gate586(.a(gate225inter10), .b(gate225inter9), .O(gate225inter11));
  nor2  gate587(.a(gate225inter11), .b(gate225inter6), .O(gate225inter12));
  nand2 gate588(.a(gate225inter12), .b(gate225inter1), .O(G706));
nand2 gate226( .a(G692), .b(G693), .O(G709) );
nand2 gate227( .a(G694), .b(G695), .O(G712) );

  xor2  gate589(.a(G697), .b(G696), .O(gate228inter0));
  nand2 gate590(.a(gate228inter0), .b(s_6), .O(gate228inter1));
  and2  gate591(.a(G697), .b(G696), .O(gate228inter2));
  inv1  gate592(.a(s_6), .O(gate228inter3));
  inv1  gate593(.a(s_7), .O(gate228inter4));
  nand2 gate594(.a(gate228inter4), .b(gate228inter3), .O(gate228inter5));
  nor2  gate595(.a(gate228inter5), .b(gate228inter2), .O(gate228inter6));
  inv1  gate596(.a(G696), .O(gate228inter7));
  inv1  gate597(.a(G697), .O(gate228inter8));
  nand2 gate598(.a(gate228inter8), .b(gate228inter7), .O(gate228inter9));
  nand2 gate599(.a(s_7), .b(gate228inter3), .O(gate228inter10));
  nor2  gate600(.a(gate228inter10), .b(gate228inter9), .O(gate228inter11));
  nor2  gate601(.a(gate228inter11), .b(gate228inter6), .O(gate228inter12));
  nand2 gate602(.a(gate228inter12), .b(gate228inter1), .O(G715));
nand2 gate229( .a(G698), .b(G699), .O(G718) );

  xor2  gate1723(.a(G701), .b(G700), .O(gate230inter0));
  nand2 gate1724(.a(gate230inter0), .b(s_168), .O(gate230inter1));
  and2  gate1725(.a(G701), .b(G700), .O(gate230inter2));
  inv1  gate1726(.a(s_168), .O(gate230inter3));
  inv1  gate1727(.a(s_169), .O(gate230inter4));
  nand2 gate1728(.a(gate230inter4), .b(gate230inter3), .O(gate230inter5));
  nor2  gate1729(.a(gate230inter5), .b(gate230inter2), .O(gate230inter6));
  inv1  gate1730(.a(G700), .O(gate230inter7));
  inv1  gate1731(.a(G701), .O(gate230inter8));
  nand2 gate1732(.a(gate230inter8), .b(gate230inter7), .O(gate230inter9));
  nand2 gate1733(.a(s_169), .b(gate230inter3), .O(gate230inter10));
  nor2  gate1734(.a(gate230inter10), .b(gate230inter9), .O(gate230inter11));
  nor2  gate1735(.a(gate230inter11), .b(gate230inter6), .O(gate230inter12));
  nand2 gate1736(.a(gate230inter12), .b(gate230inter1), .O(G721));
nand2 gate231( .a(G702), .b(G703), .O(G724) );

  xor2  gate2059(.a(G705), .b(G704), .O(gate232inter0));
  nand2 gate2060(.a(gate232inter0), .b(s_216), .O(gate232inter1));
  and2  gate2061(.a(G705), .b(G704), .O(gate232inter2));
  inv1  gate2062(.a(s_216), .O(gate232inter3));
  inv1  gate2063(.a(s_217), .O(gate232inter4));
  nand2 gate2064(.a(gate232inter4), .b(gate232inter3), .O(gate232inter5));
  nor2  gate2065(.a(gate232inter5), .b(gate232inter2), .O(gate232inter6));
  inv1  gate2066(.a(G704), .O(gate232inter7));
  inv1  gate2067(.a(G705), .O(gate232inter8));
  nand2 gate2068(.a(gate232inter8), .b(gate232inter7), .O(gate232inter9));
  nand2 gate2069(.a(s_217), .b(gate232inter3), .O(gate232inter10));
  nor2  gate2070(.a(gate232inter10), .b(gate232inter9), .O(gate232inter11));
  nor2  gate2071(.a(gate232inter11), .b(gate232inter6), .O(gate232inter12));
  nand2 gate2072(.a(gate232inter12), .b(gate232inter1), .O(G727));

  xor2  gate995(.a(G718), .b(G242), .O(gate233inter0));
  nand2 gate996(.a(gate233inter0), .b(s_64), .O(gate233inter1));
  and2  gate997(.a(G718), .b(G242), .O(gate233inter2));
  inv1  gate998(.a(s_64), .O(gate233inter3));
  inv1  gate999(.a(s_65), .O(gate233inter4));
  nand2 gate1000(.a(gate233inter4), .b(gate233inter3), .O(gate233inter5));
  nor2  gate1001(.a(gate233inter5), .b(gate233inter2), .O(gate233inter6));
  inv1  gate1002(.a(G242), .O(gate233inter7));
  inv1  gate1003(.a(G718), .O(gate233inter8));
  nand2 gate1004(.a(gate233inter8), .b(gate233inter7), .O(gate233inter9));
  nand2 gate1005(.a(s_65), .b(gate233inter3), .O(gate233inter10));
  nor2  gate1006(.a(gate233inter10), .b(gate233inter9), .O(gate233inter11));
  nor2  gate1007(.a(gate233inter11), .b(gate233inter6), .O(gate233inter12));
  nand2 gate1008(.a(gate233inter12), .b(gate233inter1), .O(G730));
nand2 gate234( .a(G245), .b(G721), .O(G733) );
nand2 gate235( .a(G248), .b(G724), .O(G736) );

  xor2  gate631(.a(G727), .b(G251), .O(gate236inter0));
  nand2 gate632(.a(gate236inter0), .b(s_12), .O(gate236inter1));
  and2  gate633(.a(G727), .b(G251), .O(gate236inter2));
  inv1  gate634(.a(s_12), .O(gate236inter3));
  inv1  gate635(.a(s_13), .O(gate236inter4));
  nand2 gate636(.a(gate236inter4), .b(gate236inter3), .O(gate236inter5));
  nor2  gate637(.a(gate236inter5), .b(gate236inter2), .O(gate236inter6));
  inv1  gate638(.a(G251), .O(gate236inter7));
  inv1  gate639(.a(G727), .O(gate236inter8));
  nand2 gate640(.a(gate236inter8), .b(gate236inter7), .O(gate236inter9));
  nand2 gate641(.a(s_13), .b(gate236inter3), .O(gate236inter10));
  nor2  gate642(.a(gate236inter10), .b(gate236inter9), .O(gate236inter11));
  nor2  gate643(.a(gate236inter11), .b(gate236inter6), .O(gate236inter12));
  nand2 gate644(.a(gate236inter12), .b(gate236inter1), .O(G739));
nand2 gate237( .a(G254), .b(G706), .O(G742) );

  xor2  gate2143(.a(G709), .b(G257), .O(gate238inter0));
  nand2 gate2144(.a(gate238inter0), .b(s_228), .O(gate238inter1));
  and2  gate2145(.a(G709), .b(G257), .O(gate238inter2));
  inv1  gate2146(.a(s_228), .O(gate238inter3));
  inv1  gate2147(.a(s_229), .O(gate238inter4));
  nand2 gate2148(.a(gate238inter4), .b(gate238inter3), .O(gate238inter5));
  nor2  gate2149(.a(gate238inter5), .b(gate238inter2), .O(gate238inter6));
  inv1  gate2150(.a(G257), .O(gate238inter7));
  inv1  gate2151(.a(G709), .O(gate238inter8));
  nand2 gate2152(.a(gate238inter8), .b(gate238inter7), .O(gate238inter9));
  nand2 gate2153(.a(s_229), .b(gate238inter3), .O(gate238inter10));
  nor2  gate2154(.a(gate238inter10), .b(gate238inter9), .O(gate238inter11));
  nor2  gate2155(.a(gate238inter11), .b(gate238inter6), .O(gate238inter12));
  nand2 gate2156(.a(gate238inter12), .b(gate238inter1), .O(G745));

  xor2  gate2045(.a(G712), .b(G260), .O(gate239inter0));
  nand2 gate2046(.a(gate239inter0), .b(s_214), .O(gate239inter1));
  and2  gate2047(.a(G712), .b(G260), .O(gate239inter2));
  inv1  gate2048(.a(s_214), .O(gate239inter3));
  inv1  gate2049(.a(s_215), .O(gate239inter4));
  nand2 gate2050(.a(gate239inter4), .b(gate239inter3), .O(gate239inter5));
  nor2  gate2051(.a(gate239inter5), .b(gate239inter2), .O(gate239inter6));
  inv1  gate2052(.a(G260), .O(gate239inter7));
  inv1  gate2053(.a(G712), .O(gate239inter8));
  nand2 gate2054(.a(gate239inter8), .b(gate239inter7), .O(gate239inter9));
  nand2 gate2055(.a(s_215), .b(gate239inter3), .O(gate239inter10));
  nor2  gate2056(.a(gate239inter10), .b(gate239inter9), .O(gate239inter11));
  nor2  gate2057(.a(gate239inter11), .b(gate239inter6), .O(gate239inter12));
  nand2 gate2058(.a(gate239inter12), .b(gate239inter1), .O(G748));
nand2 gate240( .a(G263), .b(G715), .O(G751) );
nand2 gate241( .a(G242), .b(G730), .O(G754) );
nand2 gate242( .a(G718), .b(G730), .O(G755) );

  xor2  gate2283(.a(G733), .b(G245), .O(gate243inter0));
  nand2 gate2284(.a(gate243inter0), .b(s_248), .O(gate243inter1));
  and2  gate2285(.a(G733), .b(G245), .O(gate243inter2));
  inv1  gate2286(.a(s_248), .O(gate243inter3));
  inv1  gate2287(.a(s_249), .O(gate243inter4));
  nand2 gate2288(.a(gate243inter4), .b(gate243inter3), .O(gate243inter5));
  nor2  gate2289(.a(gate243inter5), .b(gate243inter2), .O(gate243inter6));
  inv1  gate2290(.a(G245), .O(gate243inter7));
  inv1  gate2291(.a(G733), .O(gate243inter8));
  nand2 gate2292(.a(gate243inter8), .b(gate243inter7), .O(gate243inter9));
  nand2 gate2293(.a(s_249), .b(gate243inter3), .O(gate243inter10));
  nor2  gate2294(.a(gate243inter10), .b(gate243inter9), .O(gate243inter11));
  nor2  gate2295(.a(gate243inter11), .b(gate243inter6), .O(gate243inter12));
  nand2 gate2296(.a(gate243inter12), .b(gate243inter1), .O(G756));
nand2 gate244( .a(G721), .b(G733), .O(G757) );
nand2 gate245( .a(G248), .b(G736), .O(G758) );
nand2 gate246( .a(G724), .b(G736), .O(G759) );
nand2 gate247( .a(G251), .b(G739), .O(G760) );
nand2 gate248( .a(G727), .b(G739), .O(G761) );
nand2 gate249( .a(G254), .b(G742), .O(G762) );

  xor2  gate1457(.a(G742), .b(G706), .O(gate250inter0));
  nand2 gate1458(.a(gate250inter0), .b(s_130), .O(gate250inter1));
  and2  gate1459(.a(G742), .b(G706), .O(gate250inter2));
  inv1  gate1460(.a(s_130), .O(gate250inter3));
  inv1  gate1461(.a(s_131), .O(gate250inter4));
  nand2 gate1462(.a(gate250inter4), .b(gate250inter3), .O(gate250inter5));
  nor2  gate1463(.a(gate250inter5), .b(gate250inter2), .O(gate250inter6));
  inv1  gate1464(.a(G706), .O(gate250inter7));
  inv1  gate1465(.a(G742), .O(gate250inter8));
  nand2 gate1466(.a(gate250inter8), .b(gate250inter7), .O(gate250inter9));
  nand2 gate1467(.a(s_131), .b(gate250inter3), .O(gate250inter10));
  nor2  gate1468(.a(gate250inter10), .b(gate250inter9), .O(gate250inter11));
  nor2  gate1469(.a(gate250inter11), .b(gate250inter6), .O(gate250inter12));
  nand2 gate1470(.a(gate250inter12), .b(gate250inter1), .O(G763));

  xor2  gate2465(.a(G745), .b(G257), .O(gate251inter0));
  nand2 gate2466(.a(gate251inter0), .b(s_274), .O(gate251inter1));
  and2  gate2467(.a(G745), .b(G257), .O(gate251inter2));
  inv1  gate2468(.a(s_274), .O(gate251inter3));
  inv1  gate2469(.a(s_275), .O(gate251inter4));
  nand2 gate2470(.a(gate251inter4), .b(gate251inter3), .O(gate251inter5));
  nor2  gate2471(.a(gate251inter5), .b(gate251inter2), .O(gate251inter6));
  inv1  gate2472(.a(G257), .O(gate251inter7));
  inv1  gate2473(.a(G745), .O(gate251inter8));
  nand2 gate2474(.a(gate251inter8), .b(gate251inter7), .O(gate251inter9));
  nand2 gate2475(.a(s_275), .b(gate251inter3), .O(gate251inter10));
  nor2  gate2476(.a(gate251inter10), .b(gate251inter9), .O(gate251inter11));
  nor2  gate2477(.a(gate251inter11), .b(gate251inter6), .O(gate251inter12));
  nand2 gate2478(.a(gate251inter12), .b(gate251inter1), .O(G764));
nand2 gate252( .a(G709), .b(G745), .O(G765) );

  xor2  gate1415(.a(G748), .b(G260), .O(gate253inter0));
  nand2 gate1416(.a(gate253inter0), .b(s_124), .O(gate253inter1));
  and2  gate1417(.a(G748), .b(G260), .O(gate253inter2));
  inv1  gate1418(.a(s_124), .O(gate253inter3));
  inv1  gate1419(.a(s_125), .O(gate253inter4));
  nand2 gate1420(.a(gate253inter4), .b(gate253inter3), .O(gate253inter5));
  nor2  gate1421(.a(gate253inter5), .b(gate253inter2), .O(gate253inter6));
  inv1  gate1422(.a(G260), .O(gate253inter7));
  inv1  gate1423(.a(G748), .O(gate253inter8));
  nand2 gate1424(.a(gate253inter8), .b(gate253inter7), .O(gate253inter9));
  nand2 gate1425(.a(s_125), .b(gate253inter3), .O(gate253inter10));
  nor2  gate1426(.a(gate253inter10), .b(gate253inter9), .O(gate253inter11));
  nor2  gate1427(.a(gate253inter11), .b(gate253inter6), .O(gate253inter12));
  nand2 gate1428(.a(gate253inter12), .b(gate253inter1), .O(G766));

  xor2  gate2549(.a(G748), .b(G712), .O(gate254inter0));
  nand2 gate2550(.a(gate254inter0), .b(s_286), .O(gate254inter1));
  and2  gate2551(.a(G748), .b(G712), .O(gate254inter2));
  inv1  gate2552(.a(s_286), .O(gate254inter3));
  inv1  gate2553(.a(s_287), .O(gate254inter4));
  nand2 gate2554(.a(gate254inter4), .b(gate254inter3), .O(gate254inter5));
  nor2  gate2555(.a(gate254inter5), .b(gate254inter2), .O(gate254inter6));
  inv1  gate2556(.a(G712), .O(gate254inter7));
  inv1  gate2557(.a(G748), .O(gate254inter8));
  nand2 gate2558(.a(gate254inter8), .b(gate254inter7), .O(gate254inter9));
  nand2 gate2559(.a(s_287), .b(gate254inter3), .O(gate254inter10));
  nor2  gate2560(.a(gate254inter10), .b(gate254inter9), .O(gate254inter11));
  nor2  gate2561(.a(gate254inter11), .b(gate254inter6), .O(gate254inter12));
  nand2 gate2562(.a(gate254inter12), .b(gate254inter1), .O(G767));

  xor2  gate1359(.a(G751), .b(G263), .O(gate255inter0));
  nand2 gate1360(.a(gate255inter0), .b(s_116), .O(gate255inter1));
  and2  gate1361(.a(G751), .b(G263), .O(gate255inter2));
  inv1  gate1362(.a(s_116), .O(gate255inter3));
  inv1  gate1363(.a(s_117), .O(gate255inter4));
  nand2 gate1364(.a(gate255inter4), .b(gate255inter3), .O(gate255inter5));
  nor2  gate1365(.a(gate255inter5), .b(gate255inter2), .O(gate255inter6));
  inv1  gate1366(.a(G263), .O(gate255inter7));
  inv1  gate1367(.a(G751), .O(gate255inter8));
  nand2 gate1368(.a(gate255inter8), .b(gate255inter7), .O(gate255inter9));
  nand2 gate1369(.a(s_117), .b(gate255inter3), .O(gate255inter10));
  nor2  gate1370(.a(gate255inter10), .b(gate255inter9), .O(gate255inter11));
  nor2  gate1371(.a(gate255inter11), .b(gate255inter6), .O(gate255inter12));
  nand2 gate1372(.a(gate255inter12), .b(gate255inter1), .O(G768));
nand2 gate256( .a(G715), .b(G751), .O(G769) );
nand2 gate257( .a(G754), .b(G755), .O(G770) );
nand2 gate258( .a(G756), .b(G757), .O(G773) );
nand2 gate259( .a(G758), .b(G759), .O(G776) );
nand2 gate260( .a(G760), .b(G761), .O(G779) );

  xor2  gate2031(.a(G763), .b(G762), .O(gate261inter0));
  nand2 gate2032(.a(gate261inter0), .b(s_212), .O(gate261inter1));
  and2  gate2033(.a(G763), .b(G762), .O(gate261inter2));
  inv1  gate2034(.a(s_212), .O(gate261inter3));
  inv1  gate2035(.a(s_213), .O(gate261inter4));
  nand2 gate2036(.a(gate261inter4), .b(gate261inter3), .O(gate261inter5));
  nor2  gate2037(.a(gate261inter5), .b(gate261inter2), .O(gate261inter6));
  inv1  gate2038(.a(G762), .O(gate261inter7));
  inv1  gate2039(.a(G763), .O(gate261inter8));
  nand2 gate2040(.a(gate261inter8), .b(gate261inter7), .O(gate261inter9));
  nand2 gate2041(.a(s_213), .b(gate261inter3), .O(gate261inter10));
  nor2  gate2042(.a(gate261inter10), .b(gate261inter9), .O(gate261inter11));
  nor2  gate2043(.a(gate261inter11), .b(gate261inter6), .O(gate261inter12));
  nand2 gate2044(.a(gate261inter12), .b(gate261inter1), .O(G782));

  xor2  gate2717(.a(G765), .b(G764), .O(gate262inter0));
  nand2 gate2718(.a(gate262inter0), .b(s_310), .O(gate262inter1));
  and2  gate2719(.a(G765), .b(G764), .O(gate262inter2));
  inv1  gate2720(.a(s_310), .O(gate262inter3));
  inv1  gate2721(.a(s_311), .O(gate262inter4));
  nand2 gate2722(.a(gate262inter4), .b(gate262inter3), .O(gate262inter5));
  nor2  gate2723(.a(gate262inter5), .b(gate262inter2), .O(gate262inter6));
  inv1  gate2724(.a(G764), .O(gate262inter7));
  inv1  gate2725(.a(G765), .O(gate262inter8));
  nand2 gate2726(.a(gate262inter8), .b(gate262inter7), .O(gate262inter9));
  nand2 gate2727(.a(s_311), .b(gate262inter3), .O(gate262inter10));
  nor2  gate2728(.a(gate262inter10), .b(gate262inter9), .O(gate262inter11));
  nor2  gate2729(.a(gate262inter11), .b(gate262inter6), .O(gate262inter12));
  nand2 gate2730(.a(gate262inter12), .b(gate262inter1), .O(G785));
nand2 gate263( .a(G766), .b(G767), .O(G788) );

  xor2  gate2479(.a(G769), .b(G768), .O(gate264inter0));
  nand2 gate2480(.a(gate264inter0), .b(s_276), .O(gate264inter1));
  and2  gate2481(.a(G769), .b(G768), .O(gate264inter2));
  inv1  gate2482(.a(s_276), .O(gate264inter3));
  inv1  gate2483(.a(s_277), .O(gate264inter4));
  nand2 gate2484(.a(gate264inter4), .b(gate264inter3), .O(gate264inter5));
  nor2  gate2485(.a(gate264inter5), .b(gate264inter2), .O(gate264inter6));
  inv1  gate2486(.a(G768), .O(gate264inter7));
  inv1  gate2487(.a(G769), .O(gate264inter8));
  nand2 gate2488(.a(gate264inter8), .b(gate264inter7), .O(gate264inter9));
  nand2 gate2489(.a(s_277), .b(gate264inter3), .O(gate264inter10));
  nor2  gate2490(.a(gate264inter10), .b(gate264inter9), .O(gate264inter11));
  nor2  gate2491(.a(gate264inter11), .b(gate264inter6), .O(gate264inter12));
  nand2 gate2492(.a(gate264inter12), .b(gate264inter1), .O(G791));
nand2 gate265( .a(G642), .b(G770), .O(G794) );
nand2 gate266( .a(G645), .b(G773), .O(G797) );

  xor2  gate2927(.a(G776), .b(G648), .O(gate267inter0));
  nand2 gate2928(.a(gate267inter0), .b(s_340), .O(gate267inter1));
  and2  gate2929(.a(G776), .b(G648), .O(gate267inter2));
  inv1  gate2930(.a(s_340), .O(gate267inter3));
  inv1  gate2931(.a(s_341), .O(gate267inter4));
  nand2 gate2932(.a(gate267inter4), .b(gate267inter3), .O(gate267inter5));
  nor2  gate2933(.a(gate267inter5), .b(gate267inter2), .O(gate267inter6));
  inv1  gate2934(.a(G648), .O(gate267inter7));
  inv1  gate2935(.a(G776), .O(gate267inter8));
  nand2 gate2936(.a(gate267inter8), .b(gate267inter7), .O(gate267inter9));
  nand2 gate2937(.a(s_341), .b(gate267inter3), .O(gate267inter10));
  nor2  gate2938(.a(gate267inter10), .b(gate267inter9), .O(gate267inter11));
  nor2  gate2939(.a(gate267inter11), .b(gate267inter6), .O(gate267inter12));
  nand2 gate2940(.a(gate267inter12), .b(gate267inter1), .O(G800));
nand2 gate268( .a(G651), .b(G779), .O(G803) );
nand2 gate269( .a(G654), .b(G782), .O(G806) );
nand2 gate270( .a(G657), .b(G785), .O(G809) );
nand2 gate271( .a(G660), .b(G788), .O(G812) );

  xor2  gate1793(.a(G791), .b(G663), .O(gate272inter0));
  nand2 gate1794(.a(gate272inter0), .b(s_178), .O(gate272inter1));
  and2  gate1795(.a(G791), .b(G663), .O(gate272inter2));
  inv1  gate1796(.a(s_178), .O(gate272inter3));
  inv1  gate1797(.a(s_179), .O(gate272inter4));
  nand2 gate1798(.a(gate272inter4), .b(gate272inter3), .O(gate272inter5));
  nor2  gate1799(.a(gate272inter5), .b(gate272inter2), .O(gate272inter6));
  inv1  gate1800(.a(G663), .O(gate272inter7));
  inv1  gate1801(.a(G791), .O(gate272inter8));
  nand2 gate1802(.a(gate272inter8), .b(gate272inter7), .O(gate272inter9));
  nand2 gate1803(.a(s_179), .b(gate272inter3), .O(gate272inter10));
  nor2  gate1804(.a(gate272inter10), .b(gate272inter9), .O(gate272inter11));
  nor2  gate1805(.a(gate272inter11), .b(gate272inter6), .O(gate272inter12));
  nand2 gate1806(.a(gate272inter12), .b(gate272inter1), .O(G815));
nand2 gate273( .a(G642), .b(G794), .O(G818) );

  xor2  gate897(.a(G794), .b(G770), .O(gate274inter0));
  nand2 gate898(.a(gate274inter0), .b(s_50), .O(gate274inter1));
  and2  gate899(.a(G794), .b(G770), .O(gate274inter2));
  inv1  gate900(.a(s_50), .O(gate274inter3));
  inv1  gate901(.a(s_51), .O(gate274inter4));
  nand2 gate902(.a(gate274inter4), .b(gate274inter3), .O(gate274inter5));
  nor2  gate903(.a(gate274inter5), .b(gate274inter2), .O(gate274inter6));
  inv1  gate904(.a(G770), .O(gate274inter7));
  inv1  gate905(.a(G794), .O(gate274inter8));
  nand2 gate906(.a(gate274inter8), .b(gate274inter7), .O(gate274inter9));
  nand2 gate907(.a(s_51), .b(gate274inter3), .O(gate274inter10));
  nor2  gate908(.a(gate274inter10), .b(gate274inter9), .O(gate274inter11));
  nor2  gate909(.a(gate274inter11), .b(gate274inter6), .O(gate274inter12));
  nand2 gate910(.a(gate274inter12), .b(gate274inter1), .O(G819));
nand2 gate275( .a(G645), .b(G797), .O(G820) );

  xor2  gate2157(.a(G797), .b(G773), .O(gate276inter0));
  nand2 gate2158(.a(gate276inter0), .b(s_230), .O(gate276inter1));
  and2  gate2159(.a(G797), .b(G773), .O(gate276inter2));
  inv1  gate2160(.a(s_230), .O(gate276inter3));
  inv1  gate2161(.a(s_231), .O(gate276inter4));
  nand2 gate2162(.a(gate276inter4), .b(gate276inter3), .O(gate276inter5));
  nor2  gate2163(.a(gate276inter5), .b(gate276inter2), .O(gate276inter6));
  inv1  gate2164(.a(G773), .O(gate276inter7));
  inv1  gate2165(.a(G797), .O(gate276inter8));
  nand2 gate2166(.a(gate276inter8), .b(gate276inter7), .O(gate276inter9));
  nand2 gate2167(.a(s_231), .b(gate276inter3), .O(gate276inter10));
  nor2  gate2168(.a(gate276inter10), .b(gate276inter9), .O(gate276inter11));
  nor2  gate2169(.a(gate276inter11), .b(gate276inter6), .O(gate276inter12));
  nand2 gate2170(.a(gate276inter12), .b(gate276inter1), .O(G821));

  xor2  gate2521(.a(G800), .b(G648), .O(gate277inter0));
  nand2 gate2522(.a(gate277inter0), .b(s_282), .O(gate277inter1));
  and2  gate2523(.a(G800), .b(G648), .O(gate277inter2));
  inv1  gate2524(.a(s_282), .O(gate277inter3));
  inv1  gate2525(.a(s_283), .O(gate277inter4));
  nand2 gate2526(.a(gate277inter4), .b(gate277inter3), .O(gate277inter5));
  nor2  gate2527(.a(gate277inter5), .b(gate277inter2), .O(gate277inter6));
  inv1  gate2528(.a(G648), .O(gate277inter7));
  inv1  gate2529(.a(G800), .O(gate277inter8));
  nand2 gate2530(.a(gate277inter8), .b(gate277inter7), .O(gate277inter9));
  nand2 gate2531(.a(s_283), .b(gate277inter3), .O(gate277inter10));
  nor2  gate2532(.a(gate277inter10), .b(gate277inter9), .O(gate277inter11));
  nor2  gate2533(.a(gate277inter11), .b(gate277inter6), .O(gate277inter12));
  nand2 gate2534(.a(gate277inter12), .b(gate277inter1), .O(G822));
nand2 gate278( .a(G776), .b(G800), .O(G823) );
nand2 gate279( .a(G651), .b(G803), .O(G824) );
nand2 gate280( .a(G779), .b(G803), .O(G825) );
nand2 gate281( .a(G654), .b(G806), .O(G826) );
nand2 gate282( .a(G782), .b(G806), .O(G827) );

  xor2  gate1401(.a(G809), .b(G657), .O(gate283inter0));
  nand2 gate1402(.a(gate283inter0), .b(s_122), .O(gate283inter1));
  and2  gate1403(.a(G809), .b(G657), .O(gate283inter2));
  inv1  gate1404(.a(s_122), .O(gate283inter3));
  inv1  gate1405(.a(s_123), .O(gate283inter4));
  nand2 gate1406(.a(gate283inter4), .b(gate283inter3), .O(gate283inter5));
  nor2  gate1407(.a(gate283inter5), .b(gate283inter2), .O(gate283inter6));
  inv1  gate1408(.a(G657), .O(gate283inter7));
  inv1  gate1409(.a(G809), .O(gate283inter8));
  nand2 gate1410(.a(gate283inter8), .b(gate283inter7), .O(gate283inter9));
  nand2 gate1411(.a(s_123), .b(gate283inter3), .O(gate283inter10));
  nor2  gate1412(.a(gate283inter10), .b(gate283inter9), .O(gate283inter11));
  nor2  gate1413(.a(gate283inter11), .b(gate283inter6), .O(gate283inter12));
  nand2 gate1414(.a(gate283inter12), .b(gate283inter1), .O(G828));
nand2 gate284( .a(G785), .b(G809), .O(G829) );
nand2 gate285( .a(G660), .b(G812), .O(G830) );
nand2 gate286( .a(G788), .b(G812), .O(G831) );

  xor2  gate1485(.a(G815), .b(G663), .O(gate287inter0));
  nand2 gate1486(.a(gate287inter0), .b(s_134), .O(gate287inter1));
  and2  gate1487(.a(G815), .b(G663), .O(gate287inter2));
  inv1  gate1488(.a(s_134), .O(gate287inter3));
  inv1  gate1489(.a(s_135), .O(gate287inter4));
  nand2 gate1490(.a(gate287inter4), .b(gate287inter3), .O(gate287inter5));
  nor2  gate1491(.a(gate287inter5), .b(gate287inter2), .O(gate287inter6));
  inv1  gate1492(.a(G663), .O(gate287inter7));
  inv1  gate1493(.a(G815), .O(gate287inter8));
  nand2 gate1494(.a(gate287inter8), .b(gate287inter7), .O(gate287inter9));
  nand2 gate1495(.a(s_135), .b(gate287inter3), .O(gate287inter10));
  nor2  gate1496(.a(gate287inter10), .b(gate287inter9), .O(gate287inter11));
  nor2  gate1497(.a(gate287inter11), .b(gate287inter6), .O(gate287inter12));
  nand2 gate1498(.a(gate287inter12), .b(gate287inter1), .O(G832));

  xor2  gate1177(.a(G815), .b(G791), .O(gate288inter0));
  nand2 gate1178(.a(gate288inter0), .b(s_90), .O(gate288inter1));
  and2  gate1179(.a(G815), .b(G791), .O(gate288inter2));
  inv1  gate1180(.a(s_90), .O(gate288inter3));
  inv1  gate1181(.a(s_91), .O(gate288inter4));
  nand2 gate1182(.a(gate288inter4), .b(gate288inter3), .O(gate288inter5));
  nor2  gate1183(.a(gate288inter5), .b(gate288inter2), .O(gate288inter6));
  inv1  gate1184(.a(G791), .O(gate288inter7));
  inv1  gate1185(.a(G815), .O(gate288inter8));
  nand2 gate1186(.a(gate288inter8), .b(gate288inter7), .O(gate288inter9));
  nand2 gate1187(.a(s_91), .b(gate288inter3), .O(gate288inter10));
  nor2  gate1188(.a(gate288inter10), .b(gate288inter9), .O(gate288inter11));
  nor2  gate1189(.a(gate288inter11), .b(gate288inter6), .O(gate288inter12));
  nand2 gate1190(.a(gate288inter12), .b(gate288inter1), .O(G833));
nand2 gate289( .a(G818), .b(G819), .O(G834) );

  xor2  gate967(.a(G821), .b(G820), .O(gate290inter0));
  nand2 gate968(.a(gate290inter0), .b(s_60), .O(gate290inter1));
  and2  gate969(.a(G821), .b(G820), .O(gate290inter2));
  inv1  gate970(.a(s_60), .O(gate290inter3));
  inv1  gate971(.a(s_61), .O(gate290inter4));
  nand2 gate972(.a(gate290inter4), .b(gate290inter3), .O(gate290inter5));
  nor2  gate973(.a(gate290inter5), .b(gate290inter2), .O(gate290inter6));
  inv1  gate974(.a(G820), .O(gate290inter7));
  inv1  gate975(.a(G821), .O(gate290inter8));
  nand2 gate976(.a(gate290inter8), .b(gate290inter7), .O(gate290inter9));
  nand2 gate977(.a(s_61), .b(gate290inter3), .O(gate290inter10));
  nor2  gate978(.a(gate290inter10), .b(gate290inter9), .O(gate290inter11));
  nor2  gate979(.a(gate290inter11), .b(gate290inter6), .O(gate290inter12));
  nand2 gate980(.a(gate290inter12), .b(gate290inter1), .O(G847));

  xor2  gate687(.a(G823), .b(G822), .O(gate291inter0));
  nand2 gate688(.a(gate291inter0), .b(s_20), .O(gate291inter1));
  and2  gate689(.a(G823), .b(G822), .O(gate291inter2));
  inv1  gate690(.a(s_20), .O(gate291inter3));
  inv1  gate691(.a(s_21), .O(gate291inter4));
  nand2 gate692(.a(gate291inter4), .b(gate291inter3), .O(gate291inter5));
  nor2  gate693(.a(gate291inter5), .b(gate291inter2), .O(gate291inter6));
  inv1  gate694(.a(G822), .O(gate291inter7));
  inv1  gate695(.a(G823), .O(gate291inter8));
  nand2 gate696(.a(gate291inter8), .b(gate291inter7), .O(gate291inter9));
  nand2 gate697(.a(s_21), .b(gate291inter3), .O(gate291inter10));
  nor2  gate698(.a(gate291inter10), .b(gate291inter9), .O(gate291inter11));
  nor2  gate699(.a(gate291inter11), .b(gate291inter6), .O(gate291inter12));
  nand2 gate700(.a(gate291inter12), .b(gate291inter1), .O(G860));
nand2 gate292( .a(G824), .b(G825), .O(G873) );
nand2 gate293( .a(G828), .b(G829), .O(G886) );

  xor2  gate2115(.a(G833), .b(G832), .O(gate294inter0));
  nand2 gate2116(.a(gate294inter0), .b(s_224), .O(gate294inter1));
  and2  gate2117(.a(G833), .b(G832), .O(gate294inter2));
  inv1  gate2118(.a(s_224), .O(gate294inter3));
  inv1  gate2119(.a(s_225), .O(gate294inter4));
  nand2 gate2120(.a(gate294inter4), .b(gate294inter3), .O(gate294inter5));
  nor2  gate2121(.a(gate294inter5), .b(gate294inter2), .O(gate294inter6));
  inv1  gate2122(.a(G832), .O(gate294inter7));
  inv1  gate2123(.a(G833), .O(gate294inter8));
  nand2 gate2124(.a(gate294inter8), .b(gate294inter7), .O(gate294inter9));
  nand2 gate2125(.a(s_225), .b(gate294inter3), .O(gate294inter10));
  nor2  gate2126(.a(gate294inter10), .b(gate294inter9), .O(gate294inter11));
  nor2  gate2127(.a(gate294inter11), .b(gate294inter6), .O(gate294inter12));
  nand2 gate2128(.a(gate294inter12), .b(gate294inter1), .O(G899));

  xor2  gate2185(.a(G831), .b(G830), .O(gate295inter0));
  nand2 gate2186(.a(gate295inter0), .b(s_234), .O(gate295inter1));
  and2  gate2187(.a(G831), .b(G830), .O(gate295inter2));
  inv1  gate2188(.a(s_234), .O(gate295inter3));
  inv1  gate2189(.a(s_235), .O(gate295inter4));
  nand2 gate2190(.a(gate295inter4), .b(gate295inter3), .O(gate295inter5));
  nor2  gate2191(.a(gate295inter5), .b(gate295inter2), .O(gate295inter6));
  inv1  gate2192(.a(G830), .O(gate295inter7));
  inv1  gate2193(.a(G831), .O(gate295inter8));
  nand2 gate2194(.a(gate295inter8), .b(gate295inter7), .O(gate295inter9));
  nand2 gate2195(.a(s_235), .b(gate295inter3), .O(gate295inter10));
  nor2  gate2196(.a(gate295inter10), .b(gate295inter9), .O(gate295inter11));
  nor2  gate2197(.a(gate295inter11), .b(gate295inter6), .O(gate295inter12));
  nand2 gate2198(.a(gate295inter12), .b(gate295inter1), .O(G912));
nand2 gate296( .a(G826), .b(G827), .O(G925) );
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );
nand2 gate387( .a(G1), .b(G1036), .O(G1132) );

  xor2  gate1023(.a(G1039), .b(G2), .O(gate388inter0));
  nand2 gate1024(.a(gate388inter0), .b(s_68), .O(gate388inter1));
  and2  gate1025(.a(G1039), .b(G2), .O(gate388inter2));
  inv1  gate1026(.a(s_68), .O(gate388inter3));
  inv1  gate1027(.a(s_69), .O(gate388inter4));
  nand2 gate1028(.a(gate388inter4), .b(gate388inter3), .O(gate388inter5));
  nor2  gate1029(.a(gate388inter5), .b(gate388inter2), .O(gate388inter6));
  inv1  gate1030(.a(G2), .O(gate388inter7));
  inv1  gate1031(.a(G1039), .O(gate388inter8));
  nand2 gate1032(.a(gate388inter8), .b(gate388inter7), .O(gate388inter9));
  nand2 gate1033(.a(s_69), .b(gate388inter3), .O(gate388inter10));
  nor2  gate1034(.a(gate388inter10), .b(gate388inter9), .O(gate388inter11));
  nor2  gate1035(.a(gate388inter11), .b(gate388inter6), .O(gate388inter12));
  nand2 gate1036(.a(gate388inter12), .b(gate388inter1), .O(G1135));
nand2 gate389( .a(G3), .b(G1042), .O(G1138) );
nand2 gate390( .a(G4), .b(G1045), .O(G1141) );
nand2 gate391( .a(G5), .b(G1048), .O(G1144) );

  xor2  gate547(.a(G1051), .b(G6), .O(gate392inter0));
  nand2 gate548(.a(gate392inter0), .b(s_0), .O(gate392inter1));
  and2  gate549(.a(G1051), .b(G6), .O(gate392inter2));
  inv1  gate550(.a(s_0), .O(gate392inter3));
  inv1  gate551(.a(s_1), .O(gate392inter4));
  nand2 gate552(.a(gate392inter4), .b(gate392inter3), .O(gate392inter5));
  nor2  gate553(.a(gate392inter5), .b(gate392inter2), .O(gate392inter6));
  inv1  gate554(.a(G6), .O(gate392inter7));
  inv1  gate555(.a(G1051), .O(gate392inter8));
  nand2 gate556(.a(gate392inter8), .b(gate392inter7), .O(gate392inter9));
  nand2 gate557(.a(s_1), .b(gate392inter3), .O(gate392inter10));
  nor2  gate558(.a(gate392inter10), .b(gate392inter9), .O(gate392inter11));
  nor2  gate559(.a(gate392inter11), .b(gate392inter6), .O(gate392inter12));
  nand2 gate560(.a(gate392inter12), .b(gate392inter1), .O(G1147));
nand2 gate393( .a(G7), .b(G1054), .O(G1150) );
nand2 gate394( .a(G8), .b(G1057), .O(G1153) );

  xor2  gate1555(.a(G1060), .b(G9), .O(gate395inter0));
  nand2 gate1556(.a(gate395inter0), .b(s_144), .O(gate395inter1));
  and2  gate1557(.a(G1060), .b(G9), .O(gate395inter2));
  inv1  gate1558(.a(s_144), .O(gate395inter3));
  inv1  gate1559(.a(s_145), .O(gate395inter4));
  nand2 gate1560(.a(gate395inter4), .b(gate395inter3), .O(gate395inter5));
  nor2  gate1561(.a(gate395inter5), .b(gate395inter2), .O(gate395inter6));
  inv1  gate1562(.a(G9), .O(gate395inter7));
  inv1  gate1563(.a(G1060), .O(gate395inter8));
  nand2 gate1564(.a(gate395inter8), .b(gate395inter7), .O(gate395inter9));
  nand2 gate1565(.a(s_145), .b(gate395inter3), .O(gate395inter10));
  nor2  gate1566(.a(gate395inter10), .b(gate395inter9), .O(gate395inter11));
  nor2  gate1567(.a(gate395inter11), .b(gate395inter6), .O(gate395inter12));
  nand2 gate1568(.a(gate395inter12), .b(gate395inter1), .O(G1156));
nand2 gate396( .a(G10), .b(G1063), .O(G1159) );
nand2 gate397( .a(G11), .b(G1066), .O(G1162) );

  xor2  gate2269(.a(G1069), .b(G12), .O(gate398inter0));
  nand2 gate2270(.a(gate398inter0), .b(s_246), .O(gate398inter1));
  and2  gate2271(.a(G1069), .b(G12), .O(gate398inter2));
  inv1  gate2272(.a(s_246), .O(gate398inter3));
  inv1  gate2273(.a(s_247), .O(gate398inter4));
  nand2 gate2274(.a(gate398inter4), .b(gate398inter3), .O(gate398inter5));
  nor2  gate2275(.a(gate398inter5), .b(gate398inter2), .O(gate398inter6));
  inv1  gate2276(.a(G12), .O(gate398inter7));
  inv1  gate2277(.a(G1069), .O(gate398inter8));
  nand2 gate2278(.a(gate398inter8), .b(gate398inter7), .O(gate398inter9));
  nand2 gate2279(.a(s_247), .b(gate398inter3), .O(gate398inter10));
  nor2  gate2280(.a(gate398inter10), .b(gate398inter9), .O(gate398inter11));
  nor2  gate2281(.a(gate398inter11), .b(gate398inter6), .O(gate398inter12));
  nand2 gate2282(.a(gate398inter12), .b(gate398inter1), .O(G1165));

  xor2  gate827(.a(G1072), .b(G13), .O(gate399inter0));
  nand2 gate828(.a(gate399inter0), .b(s_40), .O(gate399inter1));
  and2  gate829(.a(G1072), .b(G13), .O(gate399inter2));
  inv1  gate830(.a(s_40), .O(gate399inter3));
  inv1  gate831(.a(s_41), .O(gate399inter4));
  nand2 gate832(.a(gate399inter4), .b(gate399inter3), .O(gate399inter5));
  nor2  gate833(.a(gate399inter5), .b(gate399inter2), .O(gate399inter6));
  inv1  gate834(.a(G13), .O(gate399inter7));
  inv1  gate835(.a(G1072), .O(gate399inter8));
  nand2 gate836(.a(gate399inter8), .b(gate399inter7), .O(gate399inter9));
  nand2 gate837(.a(s_41), .b(gate399inter3), .O(gate399inter10));
  nor2  gate838(.a(gate399inter10), .b(gate399inter9), .O(gate399inter11));
  nor2  gate839(.a(gate399inter11), .b(gate399inter6), .O(gate399inter12));
  nand2 gate840(.a(gate399inter12), .b(gate399inter1), .O(G1168));

  xor2  gate1933(.a(G1075), .b(G14), .O(gate400inter0));
  nand2 gate1934(.a(gate400inter0), .b(s_198), .O(gate400inter1));
  and2  gate1935(.a(G1075), .b(G14), .O(gate400inter2));
  inv1  gate1936(.a(s_198), .O(gate400inter3));
  inv1  gate1937(.a(s_199), .O(gate400inter4));
  nand2 gate1938(.a(gate400inter4), .b(gate400inter3), .O(gate400inter5));
  nor2  gate1939(.a(gate400inter5), .b(gate400inter2), .O(gate400inter6));
  inv1  gate1940(.a(G14), .O(gate400inter7));
  inv1  gate1941(.a(G1075), .O(gate400inter8));
  nand2 gate1942(.a(gate400inter8), .b(gate400inter7), .O(gate400inter9));
  nand2 gate1943(.a(s_199), .b(gate400inter3), .O(gate400inter10));
  nor2  gate1944(.a(gate400inter10), .b(gate400inter9), .O(gate400inter11));
  nor2  gate1945(.a(gate400inter11), .b(gate400inter6), .O(gate400inter12));
  nand2 gate1946(.a(gate400inter12), .b(gate400inter1), .O(G1171));

  xor2  gate1849(.a(G1078), .b(G15), .O(gate401inter0));
  nand2 gate1850(.a(gate401inter0), .b(s_186), .O(gate401inter1));
  and2  gate1851(.a(G1078), .b(G15), .O(gate401inter2));
  inv1  gate1852(.a(s_186), .O(gate401inter3));
  inv1  gate1853(.a(s_187), .O(gate401inter4));
  nand2 gate1854(.a(gate401inter4), .b(gate401inter3), .O(gate401inter5));
  nor2  gate1855(.a(gate401inter5), .b(gate401inter2), .O(gate401inter6));
  inv1  gate1856(.a(G15), .O(gate401inter7));
  inv1  gate1857(.a(G1078), .O(gate401inter8));
  nand2 gate1858(.a(gate401inter8), .b(gate401inter7), .O(gate401inter9));
  nand2 gate1859(.a(s_187), .b(gate401inter3), .O(gate401inter10));
  nor2  gate1860(.a(gate401inter10), .b(gate401inter9), .O(gate401inter11));
  nor2  gate1861(.a(gate401inter11), .b(gate401inter6), .O(gate401inter12));
  nand2 gate1862(.a(gate401inter12), .b(gate401inter1), .O(G1174));
nand2 gate402( .a(G16), .b(G1081), .O(G1177) );
nand2 gate403( .a(G17), .b(G1084), .O(G1180) );
nand2 gate404( .a(G18), .b(G1087), .O(G1183) );
nand2 gate405( .a(G19), .b(G1090), .O(G1186) );

  xor2  gate1583(.a(G1093), .b(G20), .O(gate406inter0));
  nand2 gate1584(.a(gate406inter0), .b(s_148), .O(gate406inter1));
  and2  gate1585(.a(G1093), .b(G20), .O(gate406inter2));
  inv1  gate1586(.a(s_148), .O(gate406inter3));
  inv1  gate1587(.a(s_149), .O(gate406inter4));
  nand2 gate1588(.a(gate406inter4), .b(gate406inter3), .O(gate406inter5));
  nor2  gate1589(.a(gate406inter5), .b(gate406inter2), .O(gate406inter6));
  inv1  gate1590(.a(G20), .O(gate406inter7));
  inv1  gate1591(.a(G1093), .O(gate406inter8));
  nand2 gate1592(.a(gate406inter8), .b(gate406inter7), .O(gate406inter9));
  nand2 gate1593(.a(s_149), .b(gate406inter3), .O(gate406inter10));
  nor2  gate1594(.a(gate406inter10), .b(gate406inter9), .O(gate406inter11));
  nor2  gate1595(.a(gate406inter11), .b(gate406inter6), .O(gate406inter12));
  nand2 gate1596(.a(gate406inter12), .b(gate406inter1), .O(G1189));

  xor2  gate1387(.a(G1096), .b(G21), .O(gate407inter0));
  nand2 gate1388(.a(gate407inter0), .b(s_120), .O(gate407inter1));
  and2  gate1389(.a(G1096), .b(G21), .O(gate407inter2));
  inv1  gate1390(.a(s_120), .O(gate407inter3));
  inv1  gate1391(.a(s_121), .O(gate407inter4));
  nand2 gate1392(.a(gate407inter4), .b(gate407inter3), .O(gate407inter5));
  nor2  gate1393(.a(gate407inter5), .b(gate407inter2), .O(gate407inter6));
  inv1  gate1394(.a(G21), .O(gate407inter7));
  inv1  gate1395(.a(G1096), .O(gate407inter8));
  nand2 gate1396(.a(gate407inter8), .b(gate407inter7), .O(gate407inter9));
  nand2 gate1397(.a(s_121), .b(gate407inter3), .O(gate407inter10));
  nor2  gate1398(.a(gate407inter10), .b(gate407inter9), .O(gate407inter11));
  nor2  gate1399(.a(gate407inter11), .b(gate407inter6), .O(gate407inter12));
  nand2 gate1400(.a(gate407inter12), .b(gate407inter1), .O(G1192));

  xor2  gate2311(.a(G1099), .b(G22), .O(gate408inter0));
  nand2 gate2312(.a(gate408inter0), .b(s_252), .O(gate408inter1));
  and2  gate2313(.a(G1099), .b(G22), .O(gate408inter2));
  inv1  gate2314(.a(s_252), .O(gate408inter3));
  inv1  gate2315(.a(s_253), .O(gate408inter4));
  nand2 gate2316(.a(gate408inter4), .b(gate408inter3), .O(gate408inter5));
  nor2  gate2317(.a(gate408inter5), .b(gate408inter2), .O(gate408inter6));
  inv1  gate2318(.a(G22), .O(gate408inter7));
  inv1  gate2319(.a(G1099), .O(gate408inter8));
  nand2 gate2320(.a(gate408inter8), .b(gate408inter7), .O(gate408inter9));
  nand2 gate2321(.a(s_253), .b(gate408inter3), .O(gate408inter10));
  nor2  gate2322(.a(gate408inter10), .b(gate408inter9), .O(gate408inter11));
  nor2  gate2323(.a(gate408inter11), .b(gate408inter6), .O(gate408inter12));
  nand2 gate2324(.a(gate408inter12), .b(gate408inter1), .O(G1195));

  xor2  gate1737(.a(G1102), .b(G23), .O(gate409inter0));
  nand2 gate1738(.a(gate409inter0), .b(s_170), .O(gate409inter1));
  and2  gate1739(.a(G1102), .b(G23), .O(gate409inter2));
  inv1  gate1740(.a(s_170), .O(gate409inter3));
  inv1  gate1741(.a(s_171), .O(gate409inter4));
  nand2 gate1742(.a(gate409inter4), .b(gate409inter3), .O(gate409inter5));
  nor2  gate1743(.a(gate409inter5), .b(gate409inter2), .O(gate409inter6));
  inv1  gate1744(.a(G23), .O(gate409inter7));
  inv1  gate1745(.a(G1102), .O(gate409inter8));
  nand2 gate1746(.a(gate409inter8), .b(gate409inter7), .O(gate409inter9));
  nand2 gate1747(.a(s_171), .b(gate409inter3), .O(gate409inter10));
  nor2  gate1748(.a(gate409inter10), .b(gate409inter9), .O(gate409inter11));
  nor2  gate1749(.a(gate409inter11), .b(gate409inter6), .O(gate409inter12));
  nand2 gate1750(.a(gate409inter12), .b(gate409inter1), .O(G1198));
nand2 gate410( .a(G24), .b(G1105), .O(G1201) );
nand2 gate411( .a(G25), .b(G1108), .O(G1204) );
nand2 gate412( .a(G26), .b(G1111), .O(G1207) );
nand2 gate413( .a(G27), .b(G1114), .O(G1210) );

  xor2  gate869(.a(G1117), .b(G28), .O(gate414inter0));
  nand2 gate870(.a(gate414inter0), .b(s_46), .O(gate414inter1));
  and2  gate871(.a(G1117), .b(G28), .O(gate414inter2));
  inv1  gate872(.a(s_46), .O(gate414inter3));
  inv1  gate873(.a(s_47), .O(gate414inter4));
  nand2 gate874(.a(gate414inter4), .b(gate414inter3), .O(gate414inter5));
  nor2  gate875(.a(gate414inter5), .b(gate414inter2), .O(gate414inter6));
  inv1  gate876(.a(G28), .O(gate414inter7));
  inv1  gate877(.a(G1117), .O(gate414inter8));
  nand2 gate878(.a(gate414inter8), .b(gate414inter7), .O(gate414inter9));
  nand2 gate879(.a(s_47), .b(gate414inter3), .O(gate414inter10));
  nor2  gate880(.a(gate414inter10), .b(gate414inter9), .O(gate414inter11));
  nor2  gate881(.a(gate414inter11), .b(gate414inter6), .O(gate414inter12));
  nand2 gate882(.a(gate414inter12), .b(gate414inter1), .O(G1213));
nand2 gate415( .a(G29), .b(G1120), .O(G1216) );

  xor2  gate2171(.a(G1123), .b(G30), .O(gate416inter0));
  nand2 gate2172(.a(gate416inter0), .b(s_232), .O(gate416inter1));
  and2  gate2173(.a(G1123), .b(G30), .O(gate416inter2));
  inv1  gate2174(.a(s_232), .O(gate416inter3));
  inv1  gate2175(.a(s_233), .O(gate416inter4));
  nand2 gate2176(.a(gate416inter4), .b(gate416inter3), .O(gate416inter5));
  nor2  gate2177(.a(gate416inter5), .b(gate416inter2), .O(gate416inter6));
  inv1  gate2178(.a(G30), .O(gate416inter7));
  inv1  gate2179(.a(G1123), .O(gate416inter8));
  nand2 gate2180(.a(gate416inter8), .b(gate416inter7), .O(gate416inter9));
  nand2 gate2181(.a(s_233), .b(gate416inter3), .O(gate416inter10));
  nor2  gate2182(.a(gate416inter10), .b(gate416inter9), .O(gate416inter11));
  nor2  gate2183(.a(gate416inter11), .b(gate416inter6), .O(gate416inter12));
  nand2 gate2184(.a(gate416inter12), .b(gate416inter1), .O(G1219));
nand2 gate417( .a(G31), .b(G1126), .O(G1222) );
nand2 gate418( .a(G32), .b(G1129), .O(G1225) );

  xor2  gate1709(.a(G1132), .b(G1), .O(gate419inter0));
  nand2 gate1710(.a(gate419inter0), .b(s_166), .O(gate419inter1));
  and2  gate1711(.a(G1132), .b(G1), .O(gate419inter2));
  inv1  gate1712(.a(s_166), .O(gate419inter3));
  inv1  gate1713(.a(s_167), .O(gate419inter4));
  nand2 gate1714(.a(gate419inter4), .b(gate419inter3), .O(gate419inter5));
  nor2  gate1715(.a(gate419inter5), .b(gate419inter2), .O(gate419inter6));
  inv1  gate1716(.a(G1), .O(gate419inter7));
  inv1  gate1717(.a(G1132), .O(gate419inter8));
  nand2 gate1718(.a(gate419inter8), .b(gate419inter7), .O(gate419inter9));
  nand2 gate1719(.a(s_167), .b(gate419inter3), .O(gate419inter10));
  nor2  gate1720(.a(gate419inter10), .b(gate419inter9), .O(gate419inter11));
  nor2  gate1721(.a(gate419inter11), .b(gate419inter6), .O(gate419inter12));
  nand2 gate1722(.a(gate419inter12), .b(gate419inter1), .O(G1228));

  xor2  gate1135(.a(G1132), .b(G1036), .O(gate420inter0));
  nand2 gate1136(.a(gate420inter0), .b(s_84), .O(gate420inter1));
  and2  gate1137(.a(G1132), .b(G1036), .O(gate420inter2));
  inv1  gate1138(.a(s_84), .O(gate420inter3));
  inv1  gate1139(.a(s_85), .O(gate420inter4));
  nand2 gate1140(.a(gate420inter4), .b(gate420inter3), .O(gate420inter5));
  nor2  gate1141(.a(gate420inter5), .b(gate420inter2), .O(gate420inter6));
  inv1  gate1142(.a(G1036), .O(gate420inter7));
  inv1  gate1143(.a(G1132), .O(gate420inter8));
  nand2 gate1144(.a(gate420inter8), .b(gate420inter7), .O(gate420inter9));
  nand2 gate1145(.a(s_85), .b(gate420inter3), .O(gate420inter10));
  nor2  gate1146(.a(gate420inter10), .b(gate420inter9), .O(gate420inter11));
  nor2  gate1147(.a(gate420inter11), .b(gate420inter6), .O(gate420inter12));
  nand2 gate1148(.a(gate420inter12), .b(gate420inter1), .O(G1229));

  xor2  gate1499(.a(G1135), .b(G2), .O(gate421inter0));
  nand2 gate1500(.a(gate421inter0), .b(s_136), .O(gate421inter1));
  and2  gate1501(.a(G1135), .b(G2), .O(gate421inter2));
  inv1  gate1502(.a(s_136), .O(gate421inter3));
  inv1  gate1503(.a(s_137), .O(gate421inter4));
  nand2 gate1504(.a(gate421inter4), .b(gate421inter3), .O(gate421inter5));
  nor2  gate1505(.a(gate421inter5), .b(gate421inter2), .O(gate421inter6));
  inv1  gate1506(.a(G2), .O(gate421inter7));
  inv1  gate1507(.a(G1135), .O(gate421inter8));
  nand2 gate1508(.a(gate421inter8), .b(gate421inter7), .O(gate421inter9));
  nand2 gate1509(.a(s_137), .b(gate421inter3), .O(gate421inter10));
  nor2  gate1510(.a(gate421inter10), .b(gate421inter9), .O(gate421inter11));
  nor2  gate1511(.a(gate421inter11), .b(gate421inter6), .O(gate421inter12));
  nand2 gate1512(.a(gate421inter12), .b(gate421inter1), .O(G1230));
nand2 gate422( .a(G1039), .b(G1135), .O(G1231) );
nand2 gate423( .a(G3), .b(G1138), .O(G1232) );
nand2 gate424( .a(G1042), .b(G1138), .O(G1233) );
nand2 gate425( .a(G4), .b(G1141), .O(G1234) );
nand2 gate426( .a(G1045), .b(G1141), .O(G1235) );

  xor2  gate701(.a(G1144), .b(G5), .O(gate427inter0));
  nand2 gate702(.a(gate427inter0), .b(s_22), .O(gate427inter1));
  and2  gate703(.a(G1144), .b(G5), .O(gate427inter2));
  inv1  gate704(.a(s_22), .O(gate427inter3));
  inv1  gate705(.a(s_23), .O(gate427inter4));
  nand2 gate706(.a(gate427inter4), .b(gate427inter3), .O(gate427inter5));
  nor2  gate707(.a(gate427inter5), .b(gate427inter2), .O(gate427inter6));
  inv1  gate708(.a(G5), .O(gate427inter7));
  inv1  gate709(.a(G1144), .O(gate427inter8));
  nand2 gate710(.a(gate427inter8), .b(gate427inter7), .O(gate427inter9));
  nand2 gate711(.a(s_23), .b(gate427inter3), .O(gate427inter10));
  nor2  gate712(.a(gate427inter10), .b(gate427inter9), .O(gate427inter11));
  nor2  gate713(.a(gate427inter11), .b(gate427inter6), .O(gate427inter12));
  nand2 gate714(.a(gate427inter12), .b(gate427inter1), .O(G1236));
nand2 gate428( .a(G1048), .b(G1144), .O(G1237) );
nand2 gate429( .a(G6), .b(G1147), .O(G1238) );
nand2 gate430( .a(G1051), .b(G1147), .O(G1239) );
nand2 gate431( .a(G7), .b(G1150), .O(G1240) );
nand2 gate432( .a(G1054), .b(G1150), .O(G1241) );
nand2 gate433( .a(G8), .b(G1153), .O(G1242) );
nand2 gate434( .a(G1057), .b(G1153), .O(G1243) );

  xor2  gate2227(.a(G1156), .b(G9), .O(gate435inter0));
  nand2 gate2228(.a(gate435inter0), .b(s_240), .O(gate435inter1));
  and2  gate2229(.a(G1156), .b(G9), .O(gate435inter2));
  inv1  gate2230(.a(s_240), .O(gate435inter3));
  inv1  gate2231(.a(s_241), .O(gate435inter4));
  nand2 gate2232(.a(gate435inter4), .b(gate435inter3), .O(gate435inter5));
  nor2  gate2233(.a(gate435inter5), .b(gate435inter2), .O(gate435inter6));
  inv1  gate2234(.a(G9), .O(gate435inter7));
  inv1  gate2235(.a(G1156), .O(gate435inter8));
  nand2 gate2236(.a(gate435inter8), .b(gate435inter7), .O(gate435inter9));
  nand2 gate2237(.a(s_241), .b(gate435inter3), .O(gate435inter10));
  nor2  gate2238(.a(gate435inter10), .b(gate435inter9), .O(gate435inter11));
  nor2  gate2239(.a(gate435inter11), .b(gate435inter6), .O(gate435inter12));
  nand2 gate2240(.a(gate435inter12), .b(gate435inter1), .O(G1244));

  xor2  gate1975(.a(G1156), .b(G1060), .O(gate436inter0));
  nand2 gate1976(.a(gate436inter0), .b(s_204), .O(gate436inter1));
  and2  gate1977(.a(G1156), .b(G1060), .O(gate436inter2));
  inv1  gate1978(.a(s_204), .O(gate436inter3));
  inv1  gate1979(.a(s_205), .O(gate436inter4));
  nand2 gate1980(.a(gate436inter4), .b(gate436inter3), .O(gate436inter5));
  nor2  gate1981(.a(gate436inter5), .b(gate436inter2), .O(gate436inter6));
  inv1  gate1982(.a(G1060), .O(gate436inter7));
  inv1  gate1983(.a(G1156), .O(gate436inter8));
  nand2 gate1984(.a(gate436inter8), .b(gate436inter7), .O(gate436inter9));
  nand2 gate1985(.a(s_205), .b(gate436inter3), .O(gate436inter10));
  nor2  gate1986(.a(gate436inter10), .b(gate436inter9), .O(gate436inter11));
  nor2  gate1987(.a(gate436inter11), .b(gate436inter6), .O(gate436inter12));
  nand2 gate1988(.a(gate436inter12), .b(gate436inter1), .O(G1245));

  xor2  gate2675(.a(G1159), .b(G10), .O(gate437inter0));
  nand2 gate2676(.a(gate437inter0), .b(s_304), .O(gate437inter1));
  and2  gate2677(.a(G1159), .b(G10), .O(gate437inter2));
  inv1  gate2678(.a(s_304), .O(gate437inter3));
  inv1  gate2679(.a(s_305), .O(gate437inter4));
  nand2 gate2680(.a(gate437inter4), .b(gate437inter3), .O(gate437inter5));
  nor2  gate2681(.a(gate437inter5), .b(gate437inter2), .O(gate437inter6));
  inv1  gate2682(.a(G10), .O(gate437inter7));
  inv1  gate2683(.a(G1159), .O(gate437inter8));
  nand2 gate2684(.a(gate437inter8), .b(gate437inter7), .O(gate437inter9));
  nand2 gate2685(.a(s_305), .b(gate437inter3), .O(gate437inter10));
  nor2  gate2686(.a(gate437inter10), .b(gate437inter9), .O(gate437inter11));
  nor2  gate2687(.a(gate437inter11), .b(gate437inter6), .O(gate437inter12));
  nand2 gate2688(.a(gate437inter12), .b(gate437inter1), .O(G1246));
nand2 gate438( .a(G1063), .b(G1159), .O(G1247) );

  xor2  gate2255(.a(G1162), .b(G11), .O(gate439inter0));
  nand2 gate2256(.a(gate439inter0), .b(s_244), .O(gate439inter1));
  and2  gate2257(.a(G1162), .b(G11), .O(gate439inter2));
  inv1  gate2258(.a(s_244), .O(gate439inter3));
  inv1  gate2259(.a(s_245), .O(gate439inter4));
  nand2 gate2260(.a(gate439inter4), .b(gate439inter3), .O(gate439inter5));
  nor2  gate2261(.a(gate439inter5), .b(gate439inter2), .O(gate439inter6));
  inv1  gate2262(.a(G11), .O(gate439inter7));
  inv1  gate2263(.a(G1162), .O(gate439inter8));
  nand2 gate2264(.a(gate439inter8), .b(gate439inter7), .O(gate439inter9));
  nand2 gate2265(.a(s_245), .b(gate439inter3), .O(gate439inter10));
  nor2  gate2266(.a(gate439inter10), .b(gate439inter9), .O(gate439inter11));
  nor2  gate2267(.a(gate439inter11), .b(gate439inter6), .O(gate439inter12));
  nand2 gate2268(.a(gate439inter12), .b(gate439inter1), .O(G1248));
nand2 gate440( .a(G1066), .b(G1162), .O(G1249) );
nand2 gate441( .a(G12), .b(G1165), .O(G1250) );

  xor2  gate1163(.a(G1165), .b(G1069), .O(gate442inter0));
  nand2 gate1164(.a(gate442inter0), .b(s_88), .O(gate442inter1));
  and2  gate1165(.a(G1165), .b(G1069), .O(gate442inter2));
  inv1  gate1166(.a(s_88), .O(gate442inter3));
  inv1  gate1167(.a(s_89), .O(gate442inter4));
  nand2 gate1168(.a(gate442inter4), .b(gate442inter3), .O(gate442inter5));
  nor2  gate1169(.a(gate442inter5), .b(gate442inter2), .O(gate442inter6));
  inv1  gate1170(.a(G1069), .O(gate442inter7));
  inv1  gate1171(.a(G1165), .O(gate442inter8));
  nand2 gate1172(.a(gate442inter8), .b(gate442inter7), .O(gate442inter9));
  nand2 gate1173(.a(s_89), .b(gate442inter3), .O(gate442inter10));
  nor2  gate1174(.a(gate442inter10), .b(gate442inter9), .O(gate442inter11));
  nor2  gate1175(.a(gate442inter11), .b(gate442inter6), .O(gate442inter12));
  nand2 gate1176(.a(gate442inter12), .b(gate442inter1), .O(G1251));
nand2 gate443( .a(G13), .b(G1168), .O(G1252) );
nand2 gate444( .a(G1072), .b(G1168), .O(G1253) );
nand2 gate445( .a(G14), .b(G1171), .O(G1254) );

  xor2  gate2297(.a(G1171), .b(G1075), .O(gate446inter0));
  nand2 gate2298(.a(gate446inter0), .b(s_250), .O(gate446inter1));
  and2  gate2299(.a(G1171), .b(G1075), .O(gate446inter2));
  inv1  gate2300(.a(s_250), .O(gate446inter3));
  inv1  gate2301(.a(s_251), .O(gate446inter4));
  nand2 gate2302(.a(gate446inter4), .b(gate446inter3), .O(gate446inter5));
  nor2  gate2303(.a(gate446inter5), .b(gate446inter2), .O(gate446inter6));
  inv1  gate2304(.a(G1075), .O(gate446inter7));
  inv1  gate2305(.a(G1171), .O(gate446inter8));
  nand2 gate2306(.a(gate446inter8), .b(gate446inter7), .O(gate446inter9));
  nand2 gate2307(.a(s_251), .b(gate446inter3), .O(gate446inter10));
  nor2  gate2308(.a(gate446inter10), .b(gate446inter9), .O(gate446inter11));
  nor2  gate2309(.a(gate446inter11), .b(gate446inter6), .O(gate446inter12));
  nand2 gate2310(.a(gate446inter12), .b(gate446inter1), .O(G1255));

  xor2  gate1429(.a(G1174), .b(G15), .O(gate447inter0));
  nand2 gate1430(.a(gate447inter0), .b(s_126), .O(gate447inter1));
  and2  gate1431(.a(G1174), .b(G15), .O(gate447inter2));
  inv1  gate1432(.a(s_126), .O(gate447inter3));
  inv1  gate1433(.a(s_127), .O(gate447inter4));
  nand2 gate1434(.a(gate447inter4), .b(gate447inter3), .O(gate447inter5));
  nor2  gate1435(.a(gate447inter5), .b(gate447inter2), .O(gate447inter6));
  inv1  gate1436(.a(G15), .O(gate447inter7));
  inv1  gate1437(.a(G1174), .O(gate447inter8));
  nand2 gate1438(.a(gate447inter8), .b(gate447inter7), .O(gate447inter9));
  nand2 gate1439(.a(s_127), .b(gate447inter3), .O(gate447inter10));
  nor2  gate1440(.a(gate447inter10), .b(gate447inter9), .O(gate447inter11));
  nor2  gate1441(.a(gate447inter11), .b(gate447inter6), .O(gate447inter12));
  nand2 gate1442(.a(gate447inter12), .b(gate447inter1), .O(G1256));

  xor2  gate1863(.a(G1174), .b(G1078), .O(gate448inter0));
  nand2 gate1864(.a(gate448inter0), .b(s_188), .O(gate448inter1));
  and2  gate1865(.a(G1174), .b(G1078), .O(gate448inter2));
  inv1  gate1866(.a(s_188), .O(gate448inter3));
  inv1  gate1867(.a(s_189), .O(gate448inter4));
  nand2 gate1868(.a(gate448inter4), .b(gate448inter3), .O(gate448inter5));
  nor2  gate1869(.a(gate448inter5), .b(gate448inter2), .O(gate448inter6));
  inv1  gate1870(.a(G1078), .O(gate448inter7));
  inv1  gate1871(.a(G1174), .O(gate448inter8));
  nand2 gate1872(.a(gate448inter8), .b(gate448inter7), .O(gate448inter9));
  nand2 gate1873(.a(s_189), .b(gate448inter3), .O(gate448inter10));
  nor2  gate1874(.a(gate448inter10), .b(gate448inter9), .O(gate448inter11));
  nor2  gate1875(.a(gate448inter11), .b(gate448inter6), .O(gate448inter12));
  nand2 gate1876(.a(gate448inter12), .b(gate448inter1), .O(G1257));

  xor2  gate981(.a(G1177), .b(G16), .O(gate449inter0));
  nand2 gate982(.a(gate449inter0), .b(s_62), .O(gate449inter1));
  and2  gate983(.a(G1177), .b(G16), .O(gate449inter2));
  inv1  gate984(.a(s_62), .O(gate449inter3));
  inv1  gate985(.a(s_63), .O(gate449inter4));
  nand2 gate986(.a(gate449inter4), .b(gate449inter3), .O(gate449inter5));
  nor2  gate987(.a(gate449inter5), .b(gate449inter2), .O(gate449inter6));
  inv1  gate988(.a(G16), .O(gate449inter7));
  inv1  gate989(.a(G1177), .O(gate449inter8));
  nand2 gate990(.a(gate449inter8), .b(gate449inter7), .O(gate449inter9));
  nand2 gate991(.a(s_63), .b(gate449inter3), .O(gate449inter10));
  nor2  gate992(.a(gate449inter10), .b(gate449inter9), .O(gate449inter11));
  nor2  gate993(.a(gate449inter11), .b(gate449inter6), .O(gate449inter12));
  nand2 gate994(.a(gate449inter12), .b(gate449inter1), .O(G1258));
nand2 gate450( .a(G1081), .b(G1177), .O(G1259) );

  xor2  gate1093(.a(G1180), .b(G17), .O(gate451inter0));
  nand2 gate1094(.a(gate451inter0), .b(s_78), .O(gate451inter1));
  and2  gate1095(.a(G1180), .b(G17), .O(gate451inter2));
  inv1  gate1096(.a(s_78), .O(gate451inter3));
  inv1  gate1097(.a(s_79), .O(gate451inter4));
  nand2 gate1098(.a(gate451inter4), .b(gate451inter3), .O(gate451inter5));
  nor2  gate1099(.a(gate451inter5), .b(gate451inter2), .O(gate451inter6));
  inv1  gate1100(.a(G17), .O(gate451inter7));
  inv1  gate1101(.a(G1180), .O(gate451inter8));
  nand2 gate1102(.a(gate451inter8), .b(gate451inter7), .O(gate451inter9));
  nand2 gate1103(.a(s_79), .b(gate451inter3), .O(gate451inter10));
  nor2  gate1104(.a(gate451inter10), .b(gate451inter9), .O(gate451inter11));
  nor2  gate1105(.a(gate451inter11), .b(gate451inter6), .O(gate451inter12));
  nand2 gate1106(.a(gate451inter12), .b(gate451inter1), .O(G1260));

  xor2  gate841(.a(G1180), .b(G1084), .O(gate452inter0));
  nand2 gate842(.a(gate452inter0), .b(s_42), .O(gate452inter1));
  and2  gate843(.a(G1180), .b(G1084), .O(gate452inter2));
  inv1  gate844(.a(s_42), .O(gate452inter3));
  inv1  gate845(.a(s_43), .O(gate452inter4));
  nand2 gate846(.a(gate452inter4), .b(gate452inter3), .O(gate452inter5));
  nor2  gate847(.a(gate452inter5), .b(gate452inter2), .O(gate452inter6));
  inv1  gate848(.a(G1084), .O(gate452inter7));
  inv1  gate849(.a(G1180), .O(gate452inter8));
  nand2 gate850(.a(gate452inter8), .b(gate452inter7), .O(gate452inter9));
  nand2 gate851(.a(s_43), .b(gate452inter3), .O(gate452inter10));
  nor2  gate852(.a(gate452inter10), .b(gate452inter9), .O(gate452inter11));
  nor2  gate853(.a(gate452inter11), .b(gate452inter6), .O(gate452inter12));
  nand2 gate854(.a(gate452inter12), .b(gate452inter1), .O(G1261));
nand2 gate453( .a(G18), .b(G1183), .O(G1262) );
nand2 gate454( .a(G1087), .b(G1183), .O(G1263) );

  xor2  gate1443(.a(G1186), .b(G19), .O(gate455inter0));
  nand2 gate1444(.a(gate455inter0), .b(s_128), .O(gate455inter1));
  and2  gate1445(.a(G1186), .b(G19), .O(gate455inter2));
  inv1  gate1446(.a(s_128), .O(gate455inter3));
  inv1  gate1447(.a(s_129), .O(gate455inter4));
  nand2 gate1448(.a(gate455inter4), .b(gate455inter3), .O(gate455inter5));
  nor2  gate1449(.a(gate455inter5), .b(gate455inter2), .O(gate455inter6));
  inv1  gate1450(.a(G19), .O(gate455inter7));
  inv1  gate1451(.a(G1186), .O(gate455inter8));
  nand2 gate1452(.a(gate455inter8), .b(gate455inter7), .O(gate455inter9));
  nand2 gate1453(.a(s_129), .b(gate455inter3), .O(gate455inter10));
  nor2  gate1454(.a(gate455inter10), .b(gate455inter9), .O(gate455inter11));
  nor2  gate1455(.a(gate455inter11), .b(gate455inter6), .O(gate455inter12));
  nand2 gate1456(.a(gate455inter12), .b(gate455inter1), .O(G1264));

  xor2  gate2619(.a(G1186), .b(G1090), .O(gate456inter0));
  nand2 gate2620(.a(gate456inter0), .b(s_296), .O(gate456inter1));
  and2  gate2621(.a(G1186), .b(G1090), .O(gate456inter2));
  inv1  gate2622(.a(s_296), .O(gate456inter3));
  inv1  gate2623(.a(s_297), .O(gate456inter4));
  nand2 gate2624(.a(gate456inter4), .b(gate456inter3), .O(gate456inter5));
  nor2  gate2625(.a(gate456inter5), .b(gate456inter2), .O(gate456inter6));
  inv1  gate2626(.a(G1090), .O(gate456inter7));
  inv1  gate2627(.a(G1186), .O(gate456inter8));
  nand2 gate2628(.a(gate456inter8), .b(gate456inter7), .O(gate456inter9));
  nand2 gate2629(.a(s_297), .b(gate456inter3), .O(gate456inter10));
  nor2  gate2630(.a(gate456inter10), .b(gate456inter9), .O(gate456inter11));
  nor2  gate2631(.a(gate456inter11), .b(gate456inter6), .O(gate456inter12));
  nand2 gate2632(.a(gate456inter12), .b(gate456inter1), .O(G1265));
nand2 gate457( .a(G20), .b(G1189), .O(G1266) );

  xor2  gate1051(.a(G1189), .b(G1093), .O(gate458inter0));
  nand2 gate1052(.a(gate458inter0), .b(s_72), .O(gate458inter1));
  and2  gate1053(.a(G1189), .b(G1093), .O(gate458inter2));
  inv1  gate1054(.a(s_72), .O(gate458inter3));
  inv1  gate1055(.a(s_73), .O(gate458inter4));
  nand2 gate1056(.a(gate458inter4), .b(gate458inter3), .O(gate458inter5));
  nor2  gate1057(.a(gate458inter5), .b(gate458inter2), .O(gate458inter6));
  inv1  gate1058(.a(G1093), .O(gate458inter7));
  inv1  gate1059(.a(G1189), .O(gate458inter8));
  nand2 gate1060(.a(gate458inter8), .b(gate458inter7), .O(gate458inter9));
  nand2 gate1061(.a(s_73), .b(gate458inter3), .O(gate458inter10));
  nor2  gate1062(.a(gate458inter10), .b(gate458inter9), .O(gate458inter11));
  nor2  gate1063(.a(gate458inter11), .b(gate458inter6), .O(gate458inter12));
  nand2 gate1064(.a(gate458inter12), .b(gate458inter1), .O(G1267));
nand2 gate459( .a(G21), .b(G1192), .O(G1268) );

  xor2  gate1527(.a(G1192), .b(G1096), .O(gate460inter0));
  nand2 gate1528(.a(gate460inter0), .b(s_140), .O(gate460inter1));
  and2  gate1529(.a(G1192), .b(G1096), .O(gate460inter2));
  inv1  gate1530(.a(s_140), .O(gate460inter3));
  inv1  gate1531(.a(s_141), .O(gate460inter4));
  nand2 gate1532(.a(gate460inter4), .b(gate460inter3), .O(gate460inter5));
  nor2  gate1533(.a(gate460inter5), .b(gate460inter2), .O(gate460inter6));
  inv1  gate1534(.a(G1096), .O(gate460inter7));
  inv1  gate1535(.a(G1192), .O(gate460inter8));
  nand2 gate1536(.a(gate460inter8), .b(gate460inter7), .O(gate460inter9));
  nand2 gate1537(.a(s_141), .b(gate460inter3), .O(gate460inter10));
  nor2  gate1538(.a(gate460inter10), .b(gate460inter9), .O(gate460inter11));
  nor2  gate1539(.a(gate460inter11), .b(gate460inter6), .O(gate460inter12));
  nand2 gate1540(.a(gate460inter12), .b(gate460inter1), .O(G1269));
nand2 gate461( .a(G22), .b(G1195), .O(G1270) );

  xor2  gate1569(.a(G1195), .b(G1099), .O(gate462inter0));
  nand2 gate1570(.a(gate462inter0), .b(s_146), .O(gate462inter1));
  and2  gate1571(.a(G1195), .b(G1099), .O(gate462inter2));
  inv1  gate1572(.a(s_146), .O(gate462inter3));
  inv1  gate1573(.a(s_147), .O(gate462inter4));
  nand2 gate1574(.a(gate462inter4), .b(gate462inter3), .O(gate462inter5));
  nor2  gate1575(.a(gate462inter5), .b(gate462inter2), .O(gate462inter6));
  inv1  gate1576(.a(G1099), .O(gate462inter7));
  inv1  gate1577(.a(G1195), .O(gate462inter8));
  nand2 gate1578(.a(gate462inter8), .b(gate462inter7), .O(gate462inter9));
  nand2 gate1579(.a(s_147), .b(gate462inter3), .O(gate462inter10));
  nor2  gate1580(.a(gate462inter10), .b(gate462inter9), .O(gate462inter11));
  nor2  gate1581(.a(gate462inter11), .b(gate462inter6), .O(gate462inter12));
  nand2 gate1582(.a(gate462inter12), .b(gate462inter1), .O(G1271));
nand2 gate463( .a(G23), .b(G1198), .O(G1272) );
nand2 gate464( .a(G1102), .b(G1198), .O(G1273) );
nand2 gate465( .a(G24), .b(G1201), .O(G1274) );
nand2 gate466( .a(G1105), .b(G1201), .O(G1275) );

  xor2  gate1191(.a(G1204), .b(G25), .O(gate467inter0));
  nand2 gate1192(.a(gate467inter0), .b(s_92), .O(gate467inter1));
  and2  gate1193(.a(G1204), .b(G25), .O(gate467inter2));
  inv1  gate1194(.a(s_92), .O(gate467inter3));
  inv1  gate1195(.a(s_93), .O(gate467inter4));
  nand2 gate1196(.a(gate467inter4), .b(gate467inter3), .O(gate467inter5));
  nor2  gate1197(.a(gate467inter5), .b(gate467inter2), .O(gate467inter6));
  inv1  gate1198(.a(G25), .O(gate467inter7));
  inv1  gate1199(.a(G1204), .O(gate467inter8));
  nand2 gate1200(.a(gate467inter8), .b(gate467inter7), .O(gate467inter9));
  nand2 gate1201(.a(s_93), .b(gate467inter3), .O(gate467inter10));
  nor2  gate1202(.a(gate467inter10), .b(gate467inter9), .O(gate467inter11));
  nor2  gate1203(.a(gate467inter11), .b(gate467inter6), .O(gate467inter12));
  nand2 gate1204(.a(gate467inter12), .b(gate467inter1), .O(G1276));
nand2 gate468( .a(G1108), .b(G1204), .O(G1277) );
nand2 gate469( .a(G26), .b(G1207), .O(G1278) );
nand2 gate470( .a(G1111), .b(G1207), .O(G1279) );
nand2 gate471( .a(G27), .b(G1210), .O(G1280) );
nand2 gate472( .a(G1114), .b(G1210), .O(G1281) );
nand2 gate473( .a(G28), .b(G1213), .O(G1282) );

  xor2  gate799(.a(G1213), .b(G1117), .O(gate474inter0));
  nand2 gate800(.a(gate474inter0), .b(s_36), .O(gate474inter1));
  and2  gate801(.a(G1213), .b(G1117), .O(gate474inter2));
  inv1  gate802(.a(s_36), .O(gate474inter3));
  inv1  gate803(.a(s_37), .O(gate474inter4));
  nand2 gate804(.a(gate474inter4), .b(gate474inter3), .O(gate474inter5));
  nor2  gate805(.a(gate474inter5), .b(gate474inter2), .O(gate474inter6));
  inv1  gate806(.a(G1117), .O(gate474inter7));
  inv1  gate807(.a(G1213), .O(gate474inter8));
  nand2 gate808(.a(gate474inter8), .b(gate474inter7), .O(gate474inter9));
  nand2 gate809(.a(s_37), .b(gate474inter3), .O(gate474inter10));
  nor2  gate810(.a(gate474inter10), .b(gate474inter9), .O(gate474inter11));
  nor2  gate811(.a(gate474inter11), .b(gate474inter6), .O(gate474inter12));
  nand2 gate812(.a(gate474inter12), .b(gate474inter1), .O(G1283));

  xor2  gate1107(.a(G1216), .b(G29), .O(gate475inter0));
  nand2 gate1108(.a(gate475inter0), .b(s_80), .O(gate475inter1));
  and2  gate1109(.a(G1216), .b(G29), .O(gate475inter2));
  inv1  gate1110(.a(s_80), .O(gate475inter3));
  inv1  gate1111(.a(s_81), .O(gate475inter4));
  nand2 gate1112(.a(gate475inter4), .b(gate475inter3), .O(gate475inter5));
  nor2  gate1113(.a(gate475inter5), .b(gate475inter2), .O(gate475inter6));
  inv1  gate1114(.a(G29), .O(gate475inter7));
  inv1  gate1115(.a(G1216), .O(gate475inter8));
  nand2 gate1116(.a(gate475inter8), .b(gate475inter7), .O(gate475inter9));
  nand2 gate1117(.a(s_81), .b(gate475inter3), .O(gate475inter10));
  nor2  gate1118(.a(gate475inter10), .b(gate475inter9), .O(gate475inter11));
  nor2  gate1119(.a(gate475inter11), .b(gate475inter6), .O(gate475inter12));
  nand2 gate1120(.a(gate475inter12), .b(gate475inter1), .O(G1284));
nand2 gate476( .a(G1120), .b(G1216), .O(G1285) );

  xor2  gate1065(.a(G1219), .b(G30), .O(gate477inter0));
  nand2 gate1066(.a(gate477inter0), .b(s_74), .O(gate477inter1));
  and2  gate1067(.a(G1219), .b(G30), .O(gate477inter2));
  inv1  gate1068(.a(s_74), .O(gate477inter3));
  inv1  gate1069(.a(s_75), .O(gate477inter4));
  nand2 gate1070(.a(gate477inter4), .b(gate477inter3), .O(gate477inter5));
  nor2  gate1071(.a(gate477inter5), .b(gate477inter2), .O(gate477inter6));
  inv1  gate1072(.a(G30), .O(gate477inter7));
  inv1  gate1073(.a(G1219), .O(gate477inter8));
  nand2 gate1074(.a(gate477inter8), .b(gate477inter7), .O(gate477inter9));
  nand2 gate1075(.a(s_75), .b(gate477inter3), .O(gate477inter10));
  nor2  gate1076(.a(gate477inter10), .b(gate477inter9), .O(gate477inter11));
  nor2  gate1077(.a(gate477inter11), .b(gate477inter6), .O(gate477inter12));
  nand2 gate1078(.a(gate477inter12), .b(gate477inter1), .O(G1286));
nand2 gate478( .a(G1123), .b(G1219), .O(G1287) );
nand2 gate479( .a(G31), .b(G1222), .O(G1288) );
nand2 gate480( .a(G1126), .b(G1222), .O(G1289) );
nand2 gate481( .a(G32), .b(G1225), .O(G1290) );
nand2 gate482( .a(G1129), .b(G1225), .O(G1291) );
nand2 gate483( .a(G1228), .b(G1229), .O(G1292) );
nand2 gate484( .a(G1230), .b(G1231), .O(G1293) );

  xor2  gate1877(.a(G1233), .b(G1232), .O(gate485inter0));
  nand2 gate1878(.a(gate485inter0), .b(s_190), .O(gate485inter1));
  and2  gate1879(.a(G1233), .b(G1232), .O(gate485inter2));
  inv1  gate1880(.a(s_190), .O(gate485inter3));
  inv1  gate1881(.a(s_191), .O(gate485inter4));
  nand2 gate1882(.a(gate485inter4), .b(gate485inter3), .O(gate485inter5));
  nor2  gate1883(.a(gate485inter5), .b(gate485inter2), .O(gate485inter6));
  inv1  gate1884(.a(G1232), .O(gate485inter7));
  inv1  gate1885(.a(G1233), .O(gate485inter8));
  nand2 gate1886(.a(gate485inter8), .b(gate485inter7), .O(gate485inter9));
  nand2 gate1887(.a(s_191), .b(gate485inter3), .O(gate485inter10));
  nor2  gate1888(.a(gate485inter10), .b(gate485inter9), .O(gate485inter11));
  nor2  gate1889(.a(gate485inter11), .b(gate485inter6), .O(gate485inter12));
  nand2 gate1890(.a(gate485inter12), .b(gate485inter1), .O(G1294));
nand2 gate486( .a(G1234), .b(G1235), .O(G1295) );
nand2 gate487( .a(G1236), .b(G1237), .O(G1296) );
nand2 gate488( .a(G1238), .b(G1239), .O(G1297) );
nand2 gate489( .a(G1240), .b(G1241), .O(G1298) );

  xor2  gate1121(.a(G1243), .b(G1242), .O(gate490inter0));
  nand2 gate1122(.a(gate490inter0), .b(s_82), .O(gate490inter1));
  and2  gate1123(.a(G1243), .b(G1242), .O(gate490inter2));
  inv1  gate1124(.a(s_82), .O(gate490inter3));
  inv1  gate1125(.a(s_83), .O(gate490inter4));
  nand2 gate1126(.a(gate490inter4), .b(gate490inter3), .O(gate490inter5));
  nor2  gate1127(.a(gate490inter5), .b(gate490inter2), .O(gate490inter6));
  inv1  gate1128(.a(G1242), .O(gate490inter7));
  inv1  gate1129(.a(G1243), .O(gate490inter8));
  nand2 gate1130(.a(gate490inter8), .b(gate490inter7), .O(gate490inter9));
  nand2 gate1131(.a(s_83), .b(gate490inter3), .O(gate490inter10));
  nor2  gate1132(.a(gate490inter10), .b(gate490inter9), .O(gate490inter11));
  nor2  gate1133(.a(gate490inter11), .b(gate490inter6), .O(gate490inter12));
  nand2 gate1134(.a(gate490inter12), .b(gate490inter1), .O(G1299));
nand2 gate491( .a(G1244), .b(G1245), .O(G1300) );

  xor2  gate785(.a(G1247), .b(G1246), .O(gate492inter0));
  nand2 gate786(.a(gate492inter0), .b(s_34), .O(gate492inter1));
  and2  gate787(.a(G1247), .b(G1246), .O(gate492inter2));
  inv1  gate788(.a(s_34), .O(gate492inter3));
  inv1  gate789(.a(s_35), .O(gate492inter4));
  nand2 gate790(.a(gate492inter4), .b(gate492inter3), .O(gate492inter5));
  nor2  gate791(.a(gate492inter5), .b(gate492inter2), .O(gate492inter6));
  inv1  gate792(.a(G1246), .O(gate492inter7));
  inv1  gate793(.a(G1247), .O(gate492inter8));
  nand2 gate794(.a(gate492inter8), .b(gate492inter7), .O(gate492inter9));
  nand2 gate795(.a(s_35), .b(gate492inter3), .O(gate492inter10));
  nor2  gate796(.a(gate492inter10), .b(gate492inter9), .O(gate492inter11));
  nor2  gate797(.a(gate492inter11), .b(gate492inter6), .O(gate492inter12));
  nand2 gate798(.a(gate492inter12), .b(gate492inter1), .O(G1301));
nand2 gate493( .a(G1248), .b(G1249), .O(G1302) );

  xor2  gate757(.a(G1251), .b(G1250), .O(gate494inter0));
  nand2 gate758(.a(gate494inter0), .b(s_30), .O(gate494inter1));
  and2  gate759(.a(G1251), .b(G1250), .O(gate494inter2));
  inv1  gate760(.a(s_30), .O(gate494inter3));
  inv1  gate761(.a(s_31), .O(gate494inter4));
  nand2 gate762(.a(gate494inter4), .b(gate494inter3), .O(gate494inter5));
  nor2  gate763(.a(gate494inter5), .b(gate494inter2), .O(gate494inter6));
  inv1  gate764(.a(G1250), .O(gate494inter7));
  inv1  gate765(.a(G1251), .O(gate494inter8));
  nand2 gate766(.a(gate494inter8), .b(gate494inter7), .O(gate494inter9));
  nand2 gate767(.a(s_31), .b(gate494inter3), .O(gate494inter10));
  nor2  gate768(.a(gate494inter10), .b(gate494inter9), .O(gate494inter11));
  nor2  gate769(.a(gate494inter11), .b(gate494inter6), .O(gate494inter12));
  nand2 gate770(.a(gate494inter12), .b(gate494inter1), .O(G1303));
nand2 gate495( .a(G1252), .b(G1253), .O(G1304) );

  xor2  gate2801(.a(G1255), .b(G1254), .O(gate496inter0));
  nand2 gate2802(.a(gate496inter0), .b(s_322), .O(gate496inter1));
  and2  gate2803(.a(G1255), .b(G1254), .O(gate496inter2));
  inv1  gate2804(.a(s_322), .O(gate496inter3));
  inv1  gate2805(.a(s_323), .O(gate496inter4));
  nand2 gate2806(.a(gate496inter4), .b(gate496inter3), .O(gate496inter5));
  nor2  gate2807(.a(gate496inter5), .b(gate496inter2), .O(gate496inter6));
  inv1  gate2808(.a(G1254), .O(gate496inter7));
  inv1  gate2809(.a(G1255), .O(gate496inter8));
  nand2 gate2810(.a(gate496inter8), .b(gate496inter7), .O(gate496inter9));
  nand2 gate2811(.a(s_323), .b(gate496inter3), .O(gate496inter10));
  nor2  gate2812(.a(gate496inter10), .b(gate496inter9), .O(gate496inter11));
  nor2  gate2813(.a(gate496inter11), .b(gate496inter6), .O(gate496inter12));
  nand2 gate2814(.a(gate496inter12), .b(gate496inter1), .O(G1305));

  xor2  gate1639(.a(G1257), .b(G1256), .O(gate497inter0));
  nand2 gate1640(.a(gate497inter0), .b(s_156), .O(gate497inter1));
  and2  gate1641(.a(G1257), .b(G1256), .O(gate497inter2));
  inv1  gate1642(.a(s_156), .O(gate497inter3));
  inv1  gate1643(.a(s_157), .O(gate497inter4));
  nand2 gate1644(.a(gate497inter4), .b(gate497inter3), .O(gate497inter5));
  nor2  gate1645(.a(gate497inter5), .b(gate497inter2), .O(gate497inter6));
  inv1  gate1646(.a(G1256), .O(gate497inter7));
  inv1  gate1647(.a(G1257), .O(gate497inter8));
  nand2 gate1648(.a(gate497inter8), .b(gate497inter7), .O(gate497inter9));
  nand2 gate1649(.a(s_157), .b(gate497inter3), .O(gate497inter10));
  nor2  gate1650(.a(gate497inter10), .b(gate497inter9), .O(gate497inter11));
  nor2  gate1651(.a(gate497inter11), .b(gate497inter6), .O(gate497inter12));
  nand2 gate1652(.a(gate497inter12), .b(gate497inter1), .O(G1306));
nand2 gate498( .a(G1258), .b(G1259), .O(G1307) );

  xor2  gate2087(.a(G1261), .b(G1260), .O(gate499inter0));
  nand2 gate2088(.a(gate499inter0), .b(s_220), .O(gate499inter1));
  and2  gate2089(.a(G1261), .b(G1260), .O(gate499inter2));
  inv1  gate2090(.a(s_220), .O(gate499inter3));
  inv1  gate2091(.a(s_221), .O(gate499inter4));
  nand2 gate2092(.a(gate499inter4), .b(gate499inter3), .O(gate499inter5));
  nor2  gate2093(.a(gate499inter5), .b(gate499inter2), .O(gate499inter6));
  inv1  gate2094(.a(G1260), .O(gate499inter7));
  inv1  gate2095(.a(G1261), .O(gate499inter8));
  nand2 gate2096(.a(gate499inter8), .b(gate499inter7), .O(gate499inter9));
  nand2 gate2097(.a(s_221), .b(gate499inter3), .O(gate499inter10));
  nor2  gate2098(.a(gate499inter10), .b(gate499inter9), .O(gate499inter11));
  nor2  gate2099(.a(gate499inter11), .b(gate499inter6), .O(gate499inter12));
  nand2 gate2100(.a(gate499inter12), .b(gate499inter1), .O(G1308));
nand2 gate500( .a(G1262), .b(G1263), .O(G1309) );
nand2 gate501( .a(G1264), .b(G1265), .O(G1310) );
nand2 gate502( .a(G1266), .b(G1267), .O(G1311) );

  xor2  gate2003(.a(G1269), .b(G1268), .O(gate503inter0));
  nand2 gate2004(.a(gate503inter0), .b(s_208), .O(gate503inter1));
  and2  gate2005(.a(G1269), .b(G1268), .O(gate503inter2));
  inv1  gate2006(.a(s_208), .O(gate503inter3));
  inv1  gate2007(.a(s_209), .O(gate503inter4));
  nand2 gate2008(.a(gate503inter4), .b(gate503inter3), .O(gate503inter5));
  nor2  gate2009(.a(gate503inter5), .b(gate503inter2), .O(gate503inter6));
  inv1  gate2010(.a(G1268), .O(gate503inter7));
  inv1  gate2011(.a(G1269), .O(gate503inter8));
  nand2 gate2012(.a(gate503inter8), .b(gate503inter7), .O(gate503inter9));
  nand2 gate2013(.a(s_209), .b(gate503inter3), .O(gate503inter10));
  nor2  gate2014(.a(gate503inter10), .b(gate503inter9), .O(gate503inter11));
  nor2  gate2015(.a(gate503inter11), .b(gate503inter6), .O(gate503inter12));
  nand2 gate2016(.a(gate503inter12), .b(gate503inter1), .O(G1312));
nand2 gate504( .a(G1270), .b(G1271), .O(G1313) );
nand2 gate505( .a(G1272), .b(G1273), .O(G1314) );
nand2 gate506( .a(G1274), .b(G1275), .O(G1315) );

  xor2  gate1779(.a(G1277), .b(G1276), .O(gate507inter0));
  nand2 gate1780(.a(gate507inter0), .b(s_176), .O(gate507inter1));
  and2  gate1781(.a(G1277), .b(G1276), .O(gate507inter2));
  inv1  gate1782(.a(s_176), .O(gate507inter3));
  inv1  gate1783(.a(s_177), .O(gate507inter4));
  nand2 gate1784(.a(gate507inter4), .b(gate507inter3), .O(gate507inter5));
  nor2  gate1785(.a(gate507inter5), .b(gate507inter2), .O(gate507inter6));
  inv1  gate1786(.a(G1276), .O(gate507inter7));
  inv1  gate1787(.a(G1277), .O(gate507inter8));
  nand2 gate1788(.a(gate507inter8), .b(gate507inter7), .O(gate507inter9));
  nand2 gate1789(.a(s_177), .b(gate507inter3), .O(gate507inter10));
  nor2  gate1790(.a(gate507inter10), .b(gate507inter9), .O(gate507inter11));
  nor2  gate1791(.a(gate507inter11), .b(gate507inter6), .O(gate507inter12));
  nand2 gate1792(.a(gate507inter12), .b(gate507inter1), .O(G1316));

  xor2  gate2745(.a(G1279), .b(G1278), .O(gate508inter0));
  nand2 gate2746(.a(gate508inter0), .b(s_314), .O(gate508inter1));
  and2  gate2747(.a(G1279), .b(G1278), .O(gate508inter2));
  inv1  gate2748(.a(s_314), .O(gate508inter3));
  inv1  gate2749(.a(s_315), .O(gate508inter4));
  nand2 gate2750(.a(gate508inter4), .b(gate508inter3), .O(gate508inter5));
  nor2  gate2751(.a(gate508inter5), .b(gate508inter2), .O(gate508inter6));
  inv1  gate2752(.a(G1278), .O(gate508inter7));
  inv1  gate2753(.a(G1279), .O(gate508inter8));
  nand2 gate2754(.a(gate508inter8), .b(gate508inter7), .O(gate508inter9));
  nand2 gate2755(.a(s_315), .b(gate508inter3), .O(gate508inter10));
  nor2  gate2756(.a(gate508inter10), .b(gate508inter9), .O(gate508inter11));
  nor2  gate2757(.a(gate508inter11), .b(gate508inter6), .O(gate508inter12));
  nand2 gate2758(.a(gate508inter12), .b(gate508inter1), .O(G1317));
nand2 gate509( .a(G1280), .b(G1281), .O(G1318) );
nand2 gate510( .a(G1282), .b(G1283), .O(G1319) );

  xor2  gate1821(.a(G1285), .b(G1284), .O(gate511inter0));
  nand2 gate1822(.a(gate511inter0), .b(s_182), .O(gate511inter1));
  and2  gate1823(.a(G1285), .b(G1284), .O(gate511inter2));
  inv1  gate1824(.a(s_182), .O(gate511inter3));
  inv1  gate1825(.a(s_183), .O(gate511inter4));
  nand2 gate1826(.a(gate511inter4), .b(gate511inter3), .O(gate511inter5));
  nor2  gate1827(.a(gate511inter5), .b(gate511inter2), .O(gate511inter6));
  inv1  gate1828(.a(G1284), .O(gate511inter7));
  inv1  gate1829(.a(G1285), .O(gate511inter8));
  nand2 gate1830(.a(gate511inter8), .b(gate511inter7), .O(gate511inter9));
  nand2 gate1831(.a(s_183), .b(gate511inter3), .O(gate511inter10));
  nor2  gate1832(.a(gate511inter10), .b(gate511inter9), .O(gate511inter11));
  nor2  gate1833(.a(gate511inter11), .b(gate511inter6), .O(gate511inter12));
  nand2 gate1834(.a(gate511inter12), .b(gate511inter1), .O(G1320));
nand2 gate512( .a(G1286), .b(G1287), .O(G1321) );

  xor2  gate1667(.a(G1289), .b(G1288), .O(gate513inter0));
  nand2 gate1668(.a(gate513inter0), .b(s_160), .O(gate513inter1));
  and2  gate1669(.a(G1289), .b(G1288), .O(gate513inter2));
  inv1  gate1670(.a(s_160), .O(gate513inter3));
  inv1  gate1671(.a(s_161), .O(gate513inter4));
  nand2 gate1672(.a(gate513inter4), .b(gate513inter3), .O(gate513inter5));
  nor2  gate1673(.a(gate513inter5), .b(gate513inter2), .O(gate513inter6));
  inv1  gate1674(.a(G1288), .O(gate513inter7));
  inv1  gate1675(.a(G1289), .O(gate513inter8));
  nand2 gate1676(.a(gate513inter8), .b(gate513inter7), .O(gate513inter9));
  nand2 gate1677(.a(s_161), .b(gate513inter3), .O(gate513inter10));
  nor2  gate1678(.a(gate513inter10), .b(gate513inter9), .O(gate513inter11));
  nor2  gate1679(.a(gate513inter11), .b(gate513inter6), .O(gate513inter12));
  nand2 gate1680(.a(gate513inter12), .b(gate513inter1), .O(G1322));

  xor2  gate1009(.a(G1291), .b(G1290), .O(gate514inter0));
  nand2 gate1010(.a(gate514inter0), .b(s_66), .O(gate514inter1));
  and2  gate1011(.a(G1291), .b(G1290), .O(gate514inter2));
  inv1  gate1012(.a(s_66), .O(gate514inter3));
  inv1  gate1013(.a(s_67), .O(gate514inter4));
  nand2 gate1014(.a(gate514inter4), .b(gate514inter3), .O(gate514inter5));
  nor2  gate1015(.a(gate514inter5), .b(gate514inter2), .O(gate514inter6));
  inv1  gate1016(.a(G1290), .O(gate514inter7));
  inv1  gate1017(.a(G1291), .O(gate514inter8));
  nand2 gate1018(.a(gate514inter8), .b(gate514inter7), .O(gate514inter9));
  nand2 gate1019(.a(s_67), .b(gate514inter3), .O(gate514inter10));
  nor2  gate1020(.a(gate514inter10), .b(gate514inter9), .O(gate514inter11));
  nor2  gate1021(.a(gate514inter11), .b(gate514inter6), .O(gate514inter12));
  nand2 gate1022(.a(gate514inter12), .b(gate514inter1), .O(G1323));
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule