module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);

input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;//RE__PI;

input s_0,s_1;//RE__ALLOW(00,01,10,11);
input s_2,s_3;//RE__ALLOW(00,01,10,11);
input s_4,s_5;//RE__ALLOW(00,01,10,11);
input s_6,s_7;//RE__ALLOW(00,01,10,11);
input s_8,s_9;//RE__ALLOW(00,01,10,11);
input s_10,s_11;//RE__ALLOW(00,01,10,11);
input s_12,s_13;//RE__ALLOW(00,01,10,11);
input s_14,s_15;//RE__ALLOW(00,01,10,11);
input s_16,s_17;//RE__ALLOW(00,01,10,11);
input s_18,s_19;//RE__ALLOW(00,01,10,11);
input s_20,s_21;//RE__ALLOW(00,01,10,11);
input s_22,s_23;//RE__ALLOW(00,01,10,11);
input s_24,s_25;//RE__ALLOW(00,01,10,11);
input s_26,s_27;//RE__ALLOW(00,01,10,11);
input s_28,s_29;//RE__ALLOW(00,01,10,11);
input s_30,s_31;//RE__ALLOW(00,01,10,11);
input s_32,s_33;//RE__ALLOW(00,01,10,11);
input s_34,s_35;//RE__ALLOW(00,01,10,11);
input s_36,s_37;//RE__ALLOW(00,01,10,11);
input s_38,s_39;//RE__ALLOW(00,01,10,11);
input s_40,s_41;//RE__ALLOW(00,01,10,11);
input s_42,s_43;//RE__ALLOW(00,01,10,11);
input s_44,s_45;//RE__ALLOW(00,01,10,11);
input s_46,s_47;//RE__ALLOW(00,01,10,11);
input s_48,s_49;//RE__ALLOW(00,01,10,11);
input s_50,s_51;//RE__ALLOW(00,01,10,11);
input s_52,s_53;//RE__ALLOW(00,01,10,11);
input s_54,s_55;//RE__ALLOW(00,01,10,11);
input s_56,s_57;//RE__ALLOW(00,01,10,11);
input s_58,s_59;//RE__ALLOW(00,01,10,11);
input s_60,s_61;//RE__ALLOW(00,01,10,11);
input s_62,s_63;//RE__ALLOW(00,01,10,11);
input s_64,s_65;//RE__ALLOW(00,01,10,11);
input s_66,s_67;//RE__ALLOW(00,01,10,11);
input s_68,s_69;//RE__ALLOW(00,01,10,11);
input s_70,s_71;//RE__ALLOW(00,01,10,11);
input s_72,s_73;//RE__ALLOW(00,01,10,11);
input s_74,s_75;//RE__ALLOW(00,01,10,11);
input s_76,s_77;//RE__ALLOW(00,01,10,11);
input s_78,s_79;//RE__ALLOW(00,01,10,11);
input s_80,s_81;//RE__ALLOW(00,01,10,11);
input s_82,s_83;//RE__ALLOW(00,01,10,11);
input s_84,s_85;//RE__ALLOW(00,01,10,11);
input s_86,s_87;//RE__ALLOW(00,01,10,11);
input s_88,s_89;//RE__ALLOW(00,01,10,11);
input s_90,s_91;//RE__ALLOW(00,01,10,11);
input s_92,s_93;//RE__ALLOW(00,01,10,11);
input s_94,s_95;//RE__ALLOW(00,01,10,11);
input s_96,s_97;//RE__ALLOW(00,01,10,11);
input s_98,s_99;//RE__ALLOW(00,01,10,11);
input s_100,s_101;//RE__ALLOW(00,01,10,11);
input s_102,s_103;//RE__ALLOW(00,01,10,11);
input s_104,s_105;//RE__ALLOW(00,01,10,11);
input s_106,s_107;//RE__ALLOW(00,01,10,11);
input s_108,s_109;//RE__ALLOW(00,01,10,11);
input s_110,s_111;//RE__ALLOW(00,01,10,11);
input s_112,s_113;//RE__ALLOW(00,01,10,11);
input s_114,s_115;//RE__ALLOW(00,01,10,11);
input s_116,s_117;//RE__ALLOW(00,01,10,11);
input s_118,s_119;//RE__ALLOW(00,01,10,11);
input s_120,s_121;//RE__ALLOW(00,01,10,11);
input s_122,s_123;//RE__ALLOW(00,01,10,11);
input s_124,s_125;//RE__ALLOW(00,01,10,11);
input s_126,s_127;//RE__ALLOW(00,01,10,11);
input s_128,s_129;//RE__ALLOW(00,01,10,11);
input s_130,s_131;//RE__ALLOW(00,01,10,11);
input s_132,s_133;//RE__ALLOW(00,01,10,11);
input s_134,s_135;//RE__ALLOW(00,01,10,11);
input s_136,s_137;//RE__ALLOW(00,01,10,11);
input s_138,s_139;//RE__ALLOW(00,01,10,11);
input s_140,s_141;//RE__ALLOW(00,01,10,11);
input s_142,s_143;//RE__ALLOW(00,01,10,11);
input s_144,s_145;//RE__ALLOW(00,01,10,11);
input s_146,s_147;//RE__ALLOW(00,01,10,11);
input s_148,s_149;//RE__ALLOW(00,01,10,11);
input s_150,s_151;//RE__ALLOW(00,01,10,11);
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;

  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate242inter0, gate242inter1, gate242inter2, gate242inter3, gate242inter4, gate242inter5, gate242inter6, gate242inter7, gate242inter8, gate242inter9, gate242inter10, gate242inter11, gate242inter12, gate243inter0, gate243inter1, gate243inter2, gate243inter3, gate243inter4, gate243inter5, gate243inter6, gate243inter7, gate243inter8, gate243inter9, gate243inter10, gate243inter11, gate243inter12, gate249inter0, gate249inter1, gate249inter2, gate249inter3, gate249inter4, gate249inter5, gate249inter6, gate249inter7, gate249inter8, gate249inter9, gate249inter10, gate249inter11, gate249inter12, gate466inter0, gate466inter1, gate466inter2, gate466inter3, gate466inter4, gate466inter5, gate466inter6, gate466inter7, gate466inter8, gate466inter9, gate466inter10, gate466inter11, gate466inter12, gate20inter0, gate20inter1, gate20inter2, gate20inter3, gate20inter4, gate20inter5, gate20inter6, gate20inter7, gate20inter8, gate20inter9, gate20inter10, gate20inter11, gate20inter12, gate70inter0, gate70inter1, gate70inter2, gate70inter3, gate70inter4, gate70inter5, gate70inter6, gate70inter7, gate70inter8, gate70inter9, gate70inter10, gate70inter11, gate70inter12, gate229inter0, gate229inter1, gate229inter2, gate229inter3, gate229inter4, gate229inter5, gate229inter6, gate229inter7, gate229inter8, gate229inter9, gate229inter10, gate229inter11, gate229inter12, gate53inter0, gate53inter1, gate53inter2, gate53inter3, gate53inter4, gate53inter5, gate53inter6, gate53inter7, gate53inter8, gate53inter9, gate53inter10, gate53inter11, gate53inter12, gate95inter0, gate95inter1, gate95inter2, gate95inter3, gate95inter4, gate95inter5, gate95inter6, gate95inter7, gate95inter8, gate95inter9, gate95inter10, gate95inter11, gate95inter12, gate454inter0, gate454inter1, gate454inter2, gate454inter3, gate454inter4, gate454inter5, gate454inter6, gate454inter7, gate454inter8, gate454inter9, gate454inter10, gate454inter11, gate454inter12, gate83inter0, gate83inter1, gate83inter2, gate83inter3, gate83inter4, gate83inter5, gate83inter6, gate83inter7, gate83inter8, gate83inter9, gate83inter10, gate83inter11, gate83inter12, gate190inter0, gate190inter1, gate190inter2, gate190inter3, gate190inter4, gate190inter5, gate190inter6, gate190inter7, gate190inter8, gate190inter9, gate190inter10, gate190inter11, gate190inter12, gate461inter0, gate461inter1, gate461inter2, gate461inter3, gate461inter4, gate461inter5, gate461inter6, gate461inter7, gate461inter8, gate461inter9, gate461inter10, gate461inter11, gate461inter12, gate69inter0, gate69inter1, gate69inter2, gate69inter3, gate69inter4, gate69inter5, gate69inter6, gate69inter7, gate69inter8, gate69inter9, gate69inter10, gate69inter11, gate69inter12, gate215inter0, gate215inter1, gate215inter2, gate215inter3, gate215inter4, gate215inter5, gate215inter6, gate215inter7, gate215inter8, gate215inter9, gate215inter10, gate215inter11, gate215inter12, gate121inter0, gate121inter1, gate121inter2, gate121inter3, gate121inter4, gate121inter5, gate121inter6, gate121inter7, gate121inter8, gate121inter9, gate121inter10, gate121inter11, gate121inter12, gate225inter0, gate225inter1, gate225inter2, gate225inter3, gate225inter4, gate225inter5, gate225inter6, gate225inter7, gate225inter8, gate225inter9, gate225inter10, gate225inter11, gate225inter12, gate129inter0, gate129inter1, gate129inter2, gate129inter3, gate129inter4, gate129inter5, gate129inter6, gate129inter7, gate129inter8, gate129inter9, gate129inter10, gate129inter11, gate129inter12, gate452inter0, gate452inter1, gate452inter2, gate452inter3, gate452inter4, gate452inter5, gate452inter6, gate452inter7, gate452inter8, gate452inter9, gate452inter10, gate452inter11, gate452inter12, gate504inter0, gate504inter1, gate504inter2, gate504inter3, gate504inter4, gate504inter5, gate504inter6, gate504inter7, gate504inter8, gate504inter9, gate504inter10, gate504inter11, gate504inter12, gate151inter0, gate151inter1, gate151inter2, gate151inter3, gate151inter4, gate151inter5, gate151inter6, gate151inter7, gate151inter8, gate151inter9, gate151inter10, gate151inter11, gate151inter12, gate217inter0, gate217inter1, gate217inter2, gate217inter3, gate217inter4, gate217inter5, gate217inter6, gate217inter7, gate217inter8, gate217inter9, gate217inter10, gate217inter11, gate217inter12, gate196inter0, gate196inter1, gate196inter2, gate196inter3, gate196inter4, gate196inter5, gate196inter6, gate196inter7, gate196inter8, gate196inter9, gate196inter10, gate196inter11, gate196inter12, gate231inter0, gate231inter1, gate231inter2, gate231inter3, gate231inter4, gate231inter5, gate231inter6, gate231inter7, gate231inter8, gate231inter9, gate231inter10, gate231inter11, gate231inter12, gate60inter0, gate60inter1, gate60inter2, gate60inter3, gate60inter4, gate60inter5, gate60inter6, gate60inter7, gate60inter8, gate60inter9, gate60inter10, gate60inter11, gate60inter12, gate76inter0, gate76inter1, gate76inter2, gate76inter3, gate76inter4, gate76inter5, gate76inter6, gate76inter7, gate76inter8, gate76inter9, gate76inter10, gate76inter11, gate76inter12, gate489inter0, gate489inter1, gate489inter2, gate489inter3, gate489inter4, gate489inter5, gate489inter6, gate489inter7, gate489inter8, gate489inter9, gate489inter10, gate489inter11, gate489inter12, gate482inter0, gate482inter1, gate482inter2, gate482inter3, gate482inter4, gate482inter5, gate482inter6, gate482inter7, gate482inter8, gate482inter9, gate482inter10, gate482inter11, gate482inter12, gate67inter0, gate67inter1, gate67inter2, gate67inter3, gate67inter4, gate67inter5, gate67inter6, gate67inter7, gate67inter8, gate67inter9, gate67inter10, gate67inter11, gate67inter12, gate93inter0, gate93inter1, gate93inter2, gate93inter3, gate93inter4, gate93inter5, gate93inter6, gate93inter7, gate93inter8, gate93inter9, gate93inter10, gate93inter11, gate93inter12, gate43inter0, gate43inter1, gate43inter2, gate43inter3, gate43inter4, gate43inter5, gate43inter6, gate43inter7, gate43inter8, gate43inter9, gate43inter10, gate43inter11, gate43inter12, gate423inter0, gate423inter1, gate423inter2, gate423inter3, gate423inter4, gate423inter5, gate423inter6, gate423inter7, gate423inter8, gate423inter9, gate423inter10, gate423inter11, gate423inter12, gate475inter0, gate475inter1, gate475inter2, gate475inter3, gate475inter4, gate475inter5, gate475inter6, gate475inter7, gate475inter8, gate475inter9, gate475inter10, gate475inter11, gate475inter12, gate98inter0, gate98inter1, gate98inter2, gate98inter3, gate98inter4, gate98inter5, gate98inter6, gate98inter7, gate98inter8, gate98inter9, gate98inter10, gate98inter11, gate98inter12, gate390inter0, gate390inter1, gate390inter2, gate390inter3, gate390inter4, gate390inter5, gate390inter6, gate390inter7, gate390inter8, gate390inter9, gate390inter10, gate390inter11, gate390inter12, gate459inter0, gate459inter1, gate459inter2, gate459inter3, gate459inter4, gate459inter5, gate459inter6, gate459inter7, gate459inter8, gate459inter9, gate459inter10, gate459inter11, gate459inter12, gate228inter0, gate228inter1, gate228inter2, gate228inter3, gate228inter4, gate228inter5, gate228inter6, gate228inter7, gate228inter8, gate228inter9, gate228inter10, gate228inter11, gate228inter12, gate471inter0, gate471inter1, gate471inter2, gate471inter3, gate471inter4, gate471inter5, gate471inter6, gate471inter7, gate471inter8, gate471inter9, gate471inter10, gate471inter11, gate471inter12, gate485inter0, gate485inter1, gate485inter2, gate485inter3, gate485inter4, gate485inter5, gate485inter6, gate485inter7, gate485inter8, gate485inter9, gate485inter10, gate485inter11, gate485inter12, gate124inter0, gate124inter1, gate124inter2, gate124inter3, gate124inter4, gate124inter5, gate124inter6, gate124inter7, gate124inter8, gate124inter9, gate124inter10, gate124inter11, gate124inter12, gate61inter0, gate61inter1, gate61inter2, gate61inter3, gate61inter4, gate61inter5, gate61inter6, gate61inter7, gate61inter8, gate61inter9, gate61inter10, gate61inter11, gate61inter12, gate269inter0, gate269inter1, gate269inter2, gate269inter3, gate269inter4, gate269inter5, gate269inter6, gate269inter7, gate269inter8, gate269inter9, gate269inter10, gate269inter11, gate269inter12, gate415inter0, gate415inter1, gate415inter2, gate415inter3, gate415inter4, gate415inter5, gate415inter6, gate415inter7, gate415inter8, gate415inter9, gate415inter10, gate415inter11, gate415inter12, gate444inter0, gate444inter1, gate444inter2, gate444inter3, gate444inter4, gate444inter5, gate444inter6, gate444inter7, gate444inter8, gate444inter9, gate444inter10, gate444inter11, gate444inter12, gate211inter0, gate211inter1, gate211inter2, gate211inter3, gate211inter4, gate211inter5, gate211inter6, gate211inter7, gate211inter8, gate211inter9, gate211inter10, gate211inter11, gate211inter12, gate511inter0, gate511inter1, gate511inter2, gate511inter3, gate511inter4, gate511inter5, gate511inter6, gate511inter7, gate511inter8, gate511inter9, gate511inter10, gate511inter11, gate511inter12, gate189inter0, gate189inter1, gate189inter2, gate189inter3, gate189inter4, gate189inter5, gate189inter6, gate189inter7, gate189inter8, gate189inter9, gate189inter10, gate189inter11, gate189inter12, gate82inter0, gate82inter1, gate82inter2, gate82inter3, gate82inter4, gate82inter5, gate82inter6, gate82inter7, gate82inter8, gate82inter9, gate82inter10, gate82inter11, gate82inter12, gate88inter0, gate88inter1, gate88inter2, gate88inter3, gate88inter4, gate88inter5, gate88inter6, gate88inter7, gate88inter8, gate88inter9, gate88inter10, gate88inter11, gate88inter12, gate64inter0, gate64inter1, gate64inter2, gate64inter3, gate64inter4, gate64inter5, gate64inter6, gate64inter7, gate64inter8, gate64inter9, gate64inter10, gate64inter11, gate64inter12, gate458inter0, gate458inter1, gate458inter2, gate458inter3, gate458inter4, gate458inter5, gate458inter6, gate458inter7, gate458inter8, gate458inter9, gate458inter10, gate458inter11, gate458inter12, gate30inter0, gate30inter1, gate30inter2, gate30inter3, gate30inter4, gate30inter5, gate30inter6, gate30inter7, gate30inter8, gate30inter9, gate30inter10, gate30inter11, gate30inter12, gate167inter0, gate167inter1, gate167inter2, gate167inter3, gate167inter4, gate167inter5, gate167inter6, gate167inter7, gate167inter8, gate167inter9, gate167inter10, gate167inter11, gate167inter12, gate230inter0, gate230inter1, gate230inter2, gate230inter3, gate230inter4, gate230inter5, gate230inter6, gate230inter7, gate230inter8, gate230inter9, gate230inter10, gate230inter11, gate230inter12, gate185inter0, gate185inter1, gate185inter2, gate185inter3, gate185inter4, gate185inter5, gate185inter6, gate185inter7, gate185inter8, gate185inter9, gate185inter10, gate185inter11, gate185inter12, gate497inter0, gate497inter1, gate497inter2, gate497inter3, gate497inter4, gate497inter5, gate497inter6, gate497inter7, gate497inter8, gate497inter9, gate497inter10, gate497inter11, gate497inter12, gate114inter0, gate114inter1, gate114inter2, gate114inter3, gate114inter4, gate114inter5, gate114inter6, gate114inter7, gate114inter8, gate114inter9, gate114inter10, gate114inter11, gate114inter12, gate28inter0, gate28inter1, gate28inter2, gate28inter3, gate28inter4, gate28inter5, gate28inter6, gate28inter7, gate28inter8, gate28inter9, gate28inter10, gate28inter11, gate28inter12, gate130inter0, gate130inter1, gate130inter2, gate130inter3, gate130inter4, gate130inter5, gate130inter6, gate130inter7, gate130inter8, gate130inter9, gate130inter10, gate130inter11, gate130inter12, gate166inter0, gate166inter1, gate166inter2, gate166inter3, gate166inter4, gate166inter5, gate166inter6, gate166inter7, gate166inter8, gate166inter9, gate166inter10, gate166inter11, gate166inter12, gate110inter0, gate110inter1, gate110inter2, gate110inter3, gate110inter4, gate110inter5, gate110inter6, gate110inter7, gate110inter8, gate110inter9, gate110inter10, gate110inter11, gate110inter12, gate14inter0, gate14inter1, gate14inter2, gate14inter3, gate14inter4, gate14inter5, gate14inter6, gate14inter7, gate14inter8, gate14inter9, gate14inter10, gate14inter11, gate14inter12, gate455inter0, gate455inter1, gate455inter2, gate455inter3, gate455inter4, gate455inter5, gate455inter6, gate455inter7, gate455inter8, gate455inter9, gate455inter10, gate455inter11, gate455inter12, gate11inter0, gate11inter1, gate11inter2, gate11inter3, gate11inter4, gate11inter5, gate11inter6, gate11inter7, gate11inter8, gate11inter9, gate11inter10, gate11inter11, gate11inter12, gate125inter0, gate125inter1, gate125inter2, gate125inter3, gate125inter4, gate125inter5, gate125inter6, gate125inter7, gate125inter8, gate125inter9, gate125inter10, gate125inter11, gate125inter12, gate126inter0, gate126inter1, gate126inter2, gate126inter3, gate126inter4, gate126inter5, gate126inter6, gate126inter7, gate126inter8, gate126inter9, gate126inter10, gate126inter11, gate126inter12, gate441inter0, gate441inter1, gate441inter2, gate441inter3, gate441inter4, gate441inter5, gate441inter6, gate441inter7, gate441inter8, gate441inter9, gate441inter10, gate441inter11, gate441inter12, gate120inter0, gate120inter1, gate120inter2, gate120inter3, gate120inter4, gate120inter5, gate120inter6, gate120inter7, gate120inter8, gate120inter9, gate120inter10, gate120inter11, gate120inter12, gate434inter0, gate434inter1, gate434inter2, gate434inter3, gate434inter4, gate434inter5, gate434inter6, gate434inter7, gate434inter8, gate434inter9, gate434inter10, gate434inter11, gate434inter12, gate96inter0, gate96inter1, gate96inter2, gate96inter3, gate96inter4, gate96inter5, gate96inter6, gate96inter7, gate96inter8, gate96inter9, gate96inter10, gate96inter11, gate96inter12, gate46inter0, gate46inter1, gate46inter2, gate46inter3, gate46inter4, gate46inter5, gate46inter6, gate46inter7, gate46inter8, gate46inter9, gate46inter10, gate46inter11, gate46inter12, gate72inter0, gate72inter1, gate72inter2, gate72inter3, gate72inter4, gate72inter5, gate72inter6, gate72inter7, gate72inter8, gate72inter9, gate72inter10, gate72inter11, gate72inter12, gate140inter0, gate140inter1, gate140inter2, gate140inter3, gate140inter4, gate140inter5, gate140inter6, gate140inter7, gate140inter8, gate140inter9, gate140inter10, gate140inter11, gate140inter12, gate481inter0, gate481inter1, gate481inter2, gate481inter3, gate481inter4, gate481inter5, gate481inter6, gate481inter7, gate481inter8, gate481inter9, gate481inter10, gate481inter11, gate481inter12, gate24inter0, gate24inter1, gate24inter2, gate24inter3, gate24inter4, gate24inter5, gate24inter6, gate24inter7, gate24inter8, gate24inter9, gate24inter10, gate24inter11, gate24inter12, gate387inter0, gate387inter1, gate387inter2, gate387inter3, gate387inter4, gate387inter5, gate387inter6, gate387inter7, gate387inter8, gate387inter9, gate387inter10, gate387inter11, gate387inter12;



and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );
nand2 gate9( .a(G1), .b(G2), .O(G266) );
nand2 gate10( .a(G3), .b(G4), .O(G269) );

  xor2  gate1429(.a(G6), .b(G5), .O(gate11inter0));
  nand2 gate1430(.a(gate11inter0), .b(s_126), .O(gate11inter1));
  and2  gate1431(.a(G6), .b(G5), .O(gate11inter2));
  inv1  gate1432(.a(s_126), .O(gate11inter3));
  inv1  gate1433(.a(s_127), .O(gate11inter4));
  nand2 gate1434(.a(gate11inter4), .b(gate11inter3), .O(gate11inter5));
  nor2  gate1435(.a(gate11inter5), .b(gate11inter2), .O(gate11inter6));
  inv1  gate1436(.a(G5), .O(gate11inter7));
  inv1  gate1437(.a(G6), .O(gate11inter8));
  nand2 gate1438(.a(gate11inter8), .b(gate11inter7), .O(gate11inter9));
  nand2 gate1439(.a(s_127), .b(gate11inter3), .O(gate11inter10));
  nor2  gate1440(.a(gate11inter10), .b(gate11inter9), .O(gate11inter11));
  nor2  gate1441(.a(gate11inter11), .b(gate11inter6), .O(gate11inter12));
  nand2 gate1442(.a(gate11inter12), .b(gate11inter1), .O(G272));
nand2 gate12( .a(G7), .b(G8), .O(G275) );
nand2 gate13( .a(G9), .b(G10), .O(G278) );

  xor2  gate1401(.a(G12), .b(G11), .O(gate14inter0));
  nand2 gate1402(.a(gate14inter0), .b(s_122), .O(gate14inter1));
  and2  gate1403(.a(G12), .b(G11), .O(gate14inter2));
  inv1  gate1404(.a(s_122), .O(gate14inter3));
  inv1  gate1405(.a(s_123), .O(gate14inter4));
  nand2 gate1406(.a(gate14inter4), .b(gate14inter3), .O(gate14inter5));
  nor2  gate1407(.a(gate14inter5), .b(gate14inter2), .O(gate14inter6));
  inv1  gate1408(.a(G11), .O(gate14inter7));
  inv1  gate1409(.a(G12), .O(gate14inter8));
  nand2 gate1410(.a(gate14inter8), .b(gate14inter7), .O(gate14inter9));
  nand2 gate1411(.a(s_123), .b(gate14inter3), .O(gate14inter10));
  nor2  gate1412(.a(gate14inter10), .b(gate14inter9), .O(gate14inter11));
  nor2  gate1413(.a(gate14inter11), .b(gate14inter6), .O(gate14inter12));
  nand2 gate1414(.a(gate14inter12), .b(gate14inter1), .O(G281));
nand2 gate15( .a(G13), .b(G14), .O(G284) );
nand2 gate16( .a(G15), .b(G16), .O(G287) );
nand2 gate17( .a(G17), .b(G18), .O(G290) );
nand2 gate18( .a(G19), .b(G20), .O(G293) );
nand2 gate19( .a(G21), .b(G22), .O(G296) );

  xor2  gate603(.a(G24), .b(G23), .O(gate20inter0));
  nand2 gate604(.a(gate20inter0), .b(s_8), .O(gate20inter1));
  and2  gate605(.a(G24), .b(G23), .O(gate20inter2));
  inv1  gate606(.a(s_8), .O(gate20inter3));
  inv1  gate607(.a(s_9), .O(gate20inter4));
  nand2 gate608(.a(gate20inter4), .b(gate20inter3), .O(gate20inter5));
  nor2  gate609(.a(gate20inter5), .b(gate20inter2), .O(gate20inter6));
  inv1  gate610(.a(G23), .O(gate20inter7));
  inv1  gate611(.a(G24), .O(gate20inter8));
  nand2 gate612(.a(gate20inter8), .b(gate20inter7), .O(gate20inter9));
  nand2 gate613(.a(s_9), .b(gate20inter3), .O(gate20inter10));
  nor2  gate614(.a(gate20inter10), .b(gate20inter9), .O(gate20inter11));
  nor2  gate615(.a(gate20inter11), .b(gate20inter6), .O(gate20inter12));
  nand2 gate616(.a(gate20inter12), .b(gate20inter1), .O(G299));
nand2 gate21( .a(G25), .b(G26), .O(G302) );
nand2 gate22( .a(G27), .b(G28), .O(G305) );
nand2 gate23( .a(G29), .b(G30), .O(G308) );

  xor2  gate1583(.a(G32), .b(G31), .O(gate24inter0));
  nand2 gate1584(.a(gate24inter0), .b(s_148), .O(gate24inter1));
  and2  gate1585(.a(G32), .b(G31), .O(gate24inter2));
  inv1  gate1586(.a(s_148), .O(gate24inter3));
  inv1  gate1587(.a(s_149), .O(gate24inter4));
  nand2 gate1588(.a(gate24inter4), .b(gate24inter3), .O(gate24inter5));
  nor2  gate1589(.a(gate24inter5), .b(gate24inter2), .O(gate24inter6));
  inv1  gate1590(.a(G31), .O(gate24inter7));
  inv1  gate1591(.a(G32), .O(gate24inter8));
  nand2 gate1592(.a(gate24inter8), .b(gate24inter7), .O(gate24inter9));
  nand2 gate1593(.a(s_149), .b(gate24inter3), .O(gate24inter10));
  nor2  gate1594(.a(gate24inter10), .b(gate24inter9), .O(gate24inter11));
  nor2  gate1595(.a(gate24inter11), .b(gate24inter6), .O(gate24inter12));
  nand2 gate1596(.a(gate24inter12), .b(gate24inter1), .O(G311));
nand2 gate25( .a(G1), .b(G5), .O(G314) );
nand2 gate26( .a(G9), .b(G13), .O(G317) );
nand2 gate27( .a(G2), .b(G6), .O(G320) );

  xor2  gate1345(.a(G14), .b(G10), .O(gate28inter0));
  nand2 gate1346(.a(gate28inter0), .b(s_114), .O(gate28inter1));
  and2  gate1347(.a(G14), .b(G10), .O(gate28inter2));
  inv1  gate1348(.a(s_114), .O(gate28inter3));
  inv1  gate1349(.a(s_115), .O(gate28inter4));
  nand2 gate1350(.a(gate28inter4), .b(gate28inter3), .O(gate28inter5));
  nor2  gate1351(.a(gate28inter5), .b(gate28inter2), .O(gate28inter6));
  inv1  gate1352(.a(G10), .O(gate28inter7));
  inv1  gate1353(.a(G14), .O(gate28inter8));
  nand2 gate1354(.a(gate28inter8), .b(gate28inter7), .O(gate28inter9));
  nand2 gate1355(.a(s_115), .b(gate28inter3), .O(gate28inter10));
  nor2  gate1356(.a(gate28inter10), .b(gate28inter9), .O(gate28inter11));
  nor2  gate1357(.a(gate28inter11), .b(gate28inter6), .O(gate28inter12));
  nand2 gate1358(.a(gate28inter12), .b(gate28inter1), .O(G323));
nand2 gate29( .a(G3), .b(G7), .O(G326) );

  xor2  gate1261(.a(G15), .b(G11), .O(gate30inter0));
  nand2 gate1262(.a(gate30inter0), .b(s_102), .O(gate30inter1));
  and2  gate1263(.a(G15), .b(G11), .O(gate30inter2));
  inv1  gate1264(.a(s_102), .O(gate30inter3));
  inv1  gate1265(.a(s_103), .O(gate30inter4));
  nand2 gate1266(.a(gate30inter4), .b(gate30inter3), .O(gate30inter5));
  nor2  gate1267(.a(gate30inter5), .b(gate30inter2), .O(gate30inter6));
  inv1  gate1268(.a(G11), .O(gate30inter7));
  inv1  gate1269(.a(G15), .O(gate30inter8));
  nand2 gate1270(.a(gate30inter8), .b(gate30inter7), .O(gate30inter9));
  nand2 gate1271(.a(s_103), .b(gate30inter3), .O(gate30inter10));
  nor2  gate1272(.a(gate30inter10), .b(gate30inter9), .O(gate30inter11));
  nor2  gate1273(.a(gate30inter11), .b(gate30inter6), .O(gate30inter12));
  nand2 gate1274(.a(gate30inter12), .b(gate30inter1), .O(G329));
nand2 gate31( .a(G4), .b(G8), .O(G332) );
nand2 gate32( .a(G12), .b(G16), .O(G335) );
nand2 gate33( .a(G17), .b(G21), .O(G338) );
nand2 gate34( .a(G25), .b(G29), .O(G341) );
nand2 gate35( .a(G18), .b(G22), .O(G344) );
nand2 gate36( .a(G26), .b(G30), .O(G347) );
nand2 gate37( .a(G19), .b(G23), .O(G350) );
nand2 gate38( .a(G27), .b(G31), .O(G353) );
nand2 gate39( .a(G20), .b(G24), .O(G356) );
nand2 gate40( .a(G28), .b(G32), .O(G359) );
nand2 gate41( .a(G1), .b(G266), .O(G362) );
nand2 gate42( .a(G2), .b(G266), .O(G363) );

  xor2  gate967(.a(G269), .b(G3), .O(gate43inter0));
  nand2 gate968(.a(gate43inter0), .b(s_60), .O(gate43inter1));
  and2  gate969(.a(G269), .b(G3), .O(gate43inter2));
  inv1  gate970(.a(s_60), .O(gate43inter3));
  inv1  gate971(.a(s_61), .O(gate43inter4));
  nand2 gate972(.a(gate43inter4), .b(gate43inter3), .O(gate43inter5));
  nor2  gate973(.a(gate43inter5), .b(gate43inter2), .O(gate43inter6));
  inv1  gate974(.a(G3), .O(gate43inter7));
  inv1  gate975(.a(G269), .O(gate43inter8));
  nand2 gate976(.a(gate43inter8), .b(gate43inter7), .O(gate43inter9));
  nand2 gate977(.a(s_61), .b(gate43inter3), .O(gate43inter10));
  nor2  gate978(.a(gate43inter10), .b(gate43inter9), .O(gate43inter11));
  nor2  gate979(.a(gate43inter11), .b(gate43inter6), .O(gate43inter12));
  nand2 gate980(.a(gate43inter12), .b(gate43inter1), .O(G364));
nand2 gate44( .a(G4), .b(G269), .O(G365) );
nand2 gate45( .a(G5), .b(G272), .O(G366) );

  xor2  gate1527(.a(G272), .b(G6), .O(gate46inter0));
  nand2 gate1528(.a(gate46inter0), .b(s_140), .O(gate46inter1));
  and2  gate1529(.a(G272), .b(G6), .O(gate46inter2));
  inv1  gate1530(.a(s_140), .O(gate46inter3));
  inv1  gate1531(.a(s_141), .O(gate46inter4));
  nand2 gate1532(.a(gate46inter4), .b(gate46inter3), .O(gate46inter5));
  nor2  gate1533(.a(gate46inter5), .b(gate46inter2), .O(gate46inter6));
  inv1  gate1534(.a(G6), .O(gate46inter7));
  inv1  gate1535(.a(G272), .O(gate46inter8));
  nand2 gate1536(.a(gate46inter8), .b(gate46inter7), .O(gate46inter9));
  nand2 gate1537(.a(s_141), .b(gate46inter3), .O(gate46inter10));
  nor2  gate1538(.a(gate46inter10), .b(gate46inter9), .O(gate46inter11));
  nor2  gate1539(.a(gate46inter11), .b(gate46inter6), .O(gate46inter12));
  nand2 gate1540(.a(gate46inter12), .b(gate46inter1), .O(G367));
nand2 gate47( .a(G7), .b(G275), .O(G368) );
nand2 gate48( .a(G8), .b(G275), .O(G369) );
nand2 gate49( .a(G9), .b(G278), .O(G370) );
nand2 gate50( .a(G10), .b(G278), .O(G371) );
nand2 gate51( .a(G11), .b(G281), .O(G372) );
nand2 gate52( .a(G12), .b(G281), .O(G373) );

  xor2  gate645(.a(G284), .b(G13), .O(gate53inter0));
  nand2 gate646(.a(gate53inter0), .b(s_14), .O(gate53inter1));
  and2  gate647(.a(G284), .b(G13), .O(gate53inter2));
  inv1  gate648(.a(s_14), .O(gate53inter3));
  inv1  gate649(.a(s_15), .O(gate53inter4));
  nand2 gate650(.a(gate53inter4), .b(gate53inter3), .O(gate53inter5));
  nor2  gate651(.a(gate53inter5), .b(gate53inter2), .O(gate53inter6));
  inv1  gate652(.a(G13), .O(gate53inter7));
  inv1  gate653(.a(G284), .O(gate53inter8));
  nand2 gate654(.a(gate53inter8), .b(gate53inter7), .O(gate53inter9));
  nand2 gate655(.a(s_15), .b(gate53inter3), .O(gate53inter10));
  nor2  gate656(.a(gate53inter10), .b(gate53inter9), .O(gate53inter11));
  nor2  gate657(.a(gate53inter11), .b(gate53inter6), .O(gate53inter12));
  nand2 gate658(.a(gate53inter12), .b(gate53inter1), .O(G374));
nand2 gate54( .a(G14), .b(G284), .O(G375) );
nand2 gate55( .a(G15), .b(G287), .O(G376) );
nand2 gate56( .a(G16), .b(G287), .O(G377) );
nand2 gate57( .a(G17), .b(G290), .O(G378) );
nand2 gate58( .a(G18), .b(G290), .O(G379) );
nand2 gate59( .a(G19), .b(G293), .O(G380) );

  xor2  gate883(.a(G293), .b(G20), .O(gate60inter0));
  nand2 gate884(.a(gate60inter0), .b(s_48), .O(gate60inter1));
  and2  gate885(.a(G293), .b(G20), .O(gate60inter2));
  inv1  gate886(.a(s_48), .O(gate60inter3));
  inv1  gate887(.a(s_49), .O(gate60inter4));
  nand2 gate888(.a(gate60inter4), .b(gate60inter3), .O(gate60inter5));
  nor2  gate889(.a(gate60inter5), .b(gate60inter2), .O(gate60inter6));
  inv1  gate890(.a(G20), .O(gate60inter7));
  inv1  gate891(.a(G293), .O(gate60inter8));
  nand2 gate892(.a(gate60inter8), .b(gate60inter7), .O(gate60inter9));
  nand2 gate893(.a(s_49), .b(gate60inter3), .O(gate60inter10));
  nor2  gate894(.a(gate60inter10), .b(gate60inter9), .O(gate60inter11));
  nor2  gate895(.a(gate60inter11), .b(gate60inter6), .O(gate60inter12));
  nand2 gate896(.a(gate60inter12), .b(gate60inter1), .O(G381));

  xor2  gate1107(.a(G296), .b(G21), .O(gate61inter0));
  nand2 gate1108(.a(gate61inter0), .b(s_80), .O(gate61inter1));
  and2  gate1109(.a(G296), .b(G21), .O(gate61inter2));
  inv1  gate1110(.a(s_80), .O(gate61inter3));
  inv1  gate1111(.a(s_81), .O(gate61inter4));
  nand2 gate1112(.a(gate61inter4), .b(gate61inter3), .O(gate61inter5));
  nor2  gate1113(.a(gate61inter5), .b(gate61inter2), .O(gate61inter6));
  inv1  gate1114(.a(G21), .O(gate61inter7));
  inv1  gate1115(.a(G296), .O(gate61inter8));
  nand2 gate1116(.a(gate61inter8), .b(gate61inter7), .O(gate61inter9));
  nand2 gate1117(.a(s_81), .b(gate61inter3), .O(gate61inter10));
  nor2  gate1118(.a(gate61inter10), .b(gate61inter9), .O(gate61inter11));
  nor2  gate1119(.a(gate61inter11), .b(gate61inter6), .O(gate61inter12));
  nand2 gate1120(.a(gate61inter12), .b(gate61inter1), .O(G382));
nand2 gate62( .a(G22), .b(G296), .O(G383) );
nand2 gate63( .a(G23), .b(G299), .O(G384) );

  xor2  gate1233(.a(G299), .b(G24), .O(gate64inter0));
  nand2 gate1234(.a(gate64inter0), .b(s_98), .O(gate64inter1));
  and2  gate1235(.a(G299), .b(G24), .O(gate64inter2));
  inv1  gate1236(.a(s_98), .O(gate64inter3));
  inv1  gate1237(.a(s_99), .O(gate64inter4));
  nand2 gate1238(.a(gate64inter4), .b(gate64inter3), .O(gate64inter5));
  nor2  gate1239(.a(gate64inter5), .b(gate64inter2), .O(gate64inter6));
  inv1  gate1240(.a(G24), .O(gate64inter7));
  inv1  gate1241(.a(G299), .O(gate64inter8));
  nand2 gate1242(.a(gate64inter8), .b(gate64inter7), .O(gate64inter9));
  nand2 gate1243(.a(s_99), .b(gate64inter3), .O(gate64inter10));
  nor2  gate1244(.a(gate64inter10), .b(gate64inter9), .O(gate64inter11));
  nor2  gate1245(.a(gate64inter11), .b(gate64inter6), .O(gate64inter12));
  nand2 gate1246(.a(gate64inter12), .b(gate64inter1), .O(G385));
nand2 gate65( .a(G25), .b(G302), .O(G386) );
nand2 gate66( .a(G26), .b(G302), .O(G387) );

  xor2  gate939(.a(G305), .b(G27), .O(gate67inter0));
  nand2 gate940(.a(gate67inter0), .b(s_56), .O(gate67inter1));
  and2  gate941(.a(G305), .b(G27), .O(gate67inter2));
  inv1  gate942(.a(s_56), .O(gate67inter3));
  inv1  gate943(.a(s_57), .O(gate67inter4));
  nand2 gate944(.a(gate67inter4), .b(gate67inter3), .O(gate67inter5));
  nor2  gate945(.a(gate67inter5), .b(gate67inter2), .O(gate67inter6));
  inv1  gate946(.a(G27), .O(gate67inter7));
  inv1  gate947(.a(G305), .O(gate67inter8));
  nand2 gate948(.a(gate67inter8), .b(gate67inter7), .O(gate67inter9));
  nand2 gate949(.a(s_57), .b(gate67inter3), .O(gate67inter10));
  nor2  gate950(.a(gate67inter10), .b(gate67inter9), .O(gate67inter11));
  nor2  gate951(.a(gate67inter11), .b(gate67inter6), .O(gate67inter12));
  nand2 gate952(.a(gate67inter12), .b(gate67inter1), .O(G388));
nand2 gate68( .a(G28), .b(G305), .O(G389) );

  xor2  gate729(.a(G308), .b(G29), .O(gate69inter0));
  nand2 gate730(.a(gate69inter0), .b(s_26), .O(gate69inter1));
  and2  gate731(.a(G308), .b(G29), .O(gate69inter2));
  inv1  gate732(.a(s_26), .O(gate69inter3));
  inv1  gate733(.a(s_27), .O(gate69inter4));
  nand2 gate734(.a(gate69inter4), .b(gate69inter3), .O(gate69inter5));
  nor2  gate735(.a(gate69inter5), .b(gate69inter2), .O(gate69inter6));
  inv1  gate736(.a(G29), .O(gate69inter7));
  inv1  gate737(.a(G308), .O(gate69inter8));
  nand2 gate738(.a(gate69inter8), .b(gate69inter7), .O(gate69inter9));
  nand2 gate739(.a(s_27), .b(gate69inter3), .O(gate69inter10));
  nor2  gate740(.a(gate69inter10), .b(gate69inter9), .O(gate69inter11));
  nor2  gate741(.a(gate69inter11), .b(gate69inter6), .O(gate69inter12));
  nand2 gate742(.a(gate69inter12), .b(gate69inter1), .O(G390));

  xor2  gate617(.a(G308), .b(G30), .O(gate70inter0));
  nand2 gate618(.a(gate70inter0), .b(s_10), .O(gate70inter1));
  and2  gate619(.a(G308), .b(G30), .O(gate70inter2));
  inv1  gate620(.a(s_10), .O(gate70inter3));
  inv1  gate621(.a(s_11), .O(gate70inter4));
  nand2 gate622(.a(gate70inter4), .b(gate70inter3), .O(gate70inter5));
  nor2  gate623(.a(gate70inter5), .b(gate70inter2), .O(gate70inter6));
  inv1  gate624(.a(G30), .O(gate70inter7));
  inv1  gate625(.a(G308), .O(gate70inter8));
  nand2 gate626(.a(gate70inter8), .b(gate70inter7), .O(gate70inter9));
  nand2 gate627(.a(s_11), .b(gate70inter3), .O(gate70inter10));
  nor2  gate628(.a(gate70inter10), .b(gate70inter9), .O(gate70inter11));
  nor2  gate629(.a(gate70inter11), .b(gate70inter6), .O(gate70inter12));
  nand2 gate630(.a(gate70inter12), .b(gate70inter1), .O(G391));
nand2 gate71( .a(G31), .b(G311), .O(G392) );

  xor2  gate1541(.a(G311), .b(G32), .O(gate72inter0));
  nand2 gate1542(.a(gate72inter0), .b(s_142), .O(gate72inter1));
  and2  gate1543(.a(G311), .b(G32), .O(gate72inter2));
  inv1  gate1544(.a(s_142), .O(gate72inter3));
  inv1  gate1545(.a(s_143), .O(gate72inter4));
  nand2 gate1546(.a(gate72inter4), .b(gate72inter3), .O(gate72inter5));
  nor2  gate1547(.a(gate72inter5), .b(gate72inter2), .O(gate72inter6));
  inv1  gate1548(.a(G32), .O(gate72inter7));
  inv1  gate1549(.a(G311), .O(gate72inter8));
  nand2 gate1550(.a(gate72inter8), .b(gate72inter7), .O(gate72inter9));
  nand2 gate1551(.a(s_143), .b(gate72inter3), .O(gate72inter10));
  nor2  gate1552(.a(gate72inter10), .b(gate72inter9), .O(gate72inter11));
  nor2  gate1553(.a(gate72inter11), .b(gate72inter6), .O(gate72inter12));
  nand2 gate1554(.a(gate72inter12), .b(gate72inter1), .O(G393));
nand2 gate73( .a(G1), .b(G314), .O(G394) );
nand2 gate74( .a(G5), .b(G314), .O(G395) );
nand2 gate75( .a(G9), .b(G317), .O(G396) );

  xor2  gate897(.a(G317), .b(G13), .O(gate76inter0));
  nand2 gate898(.a(gate76inter0), .b(s_50), .O(gate76inter1));
  and2  gate899(.a(G317), .b(G13), .O(gate76inter2));
  inv1  gate900(.a(s_50), .O(gate76inter3));
  inv1  gate901(.a(s_51), .O(gate76inter4));
  nand2 gate902(.a(gate76inter4), .b(gate76inter3), .O(gate76inter5));
  nor2  gate903(.a(gate76inter5), .b(gate76inter2), .O(gate76inter6));
  inv1  gate904(.a(G13), .O(gate76inter7));
  inv1  gate905(.a(G317), .O(gate76inter8));
  nand2 gate906(.a(gate76inter8), .b(gate76inter7), .O(gate76inter9));
  nand2 gate907(.a(s_51), .b(gate76inter3), .O(gate76inter10));
  nor2  gate908(.a(gate76inter10), .b(gate76inter9), .O(gate76inter11));
  nor2  gate909(.a(gate76inter11), .b(gate76inter6), .O(gate76inter12));
  nand2 gate910(.a(gate76inter12), .b(gate76inter1), .O(G397));
nand2 gate77( .a(G2), .b(G320), .O(G398) );
nand2 gate78( .a(G6), .b(G320), .O(G399) );
nand2 gate79( .a(G10), .b(G323), .O(G400) );
nand2 gate80( .a(G14), .b(G323), .O(G401) );
nand2 gate81( .a(G3), .b(G326), .O(G402) );

  xor2  gate1205(.a(G326), .b(G7), .O(gate82inter0));
  nand2 gate1206(.a(gate82inter0), .b(s_94), .O(gate82inter1));
  and2  gate1207(.a(G326), .b(G7), .O(gate82inter2));
  inv1  gate1208(.a(s_94), .O(gate82inter3));
  inv1  gate1209(.a(s_95), .O(gate82inter4));
  nand2 gate1210(.a(gate82inter4), .b(gate82inter3), .O(gate82inter5));
  nor2  gate1211(.a(gate82inter5), .b(gate82inter2), .O(gate82inter6));
  inv1  gate1212(.a(G7), .O(gate82inter7));
  inv1  gate1213(.a(G326), .O(gate82inter8));
  nand2 gate1214(.a(gate82inter8), .b(gate82inter7), .O(gate82inter9));
  nand2 gate1215(.a(s_95), .b(gate82inter3), .O(gate82inter10));
  nor2  gate1216(.a(gate82inter10), .b(gate82inter9), .O(gate82inter11));
  nor2  gate1217(.a(gate82inter11), .b(gate82inter6), .O(gate82inter12));
  nand2 gate1218(.a(gate82inter12), .b(gate82inter1), .O(G403));

  xor2  gate687(.a(G329), .b(G11), .O(gate83inter0));
  nand2 gate688(.a(gate83inter0), .b(s_20), .O(gate83inter1));
  and2  gate689(.a(G329), .b(G11), .O(gate83inter2));
  inv1  gate690(.a(s_20), .O(gate83inter3));
  inv1  gate691(.a(s_21), .O(gate83inter4));
  nand2 gate692(.a(gate83inter4), .b(gate83inter3), .O(gate83inter5));
  nor2  gate693(.a(gate83inter5), .b(gate83inter2), .O(gate83inter6));
  inv1  gate694(.a(G11), .O(gate83inter7));
  inv1  gate695(.a(G329), .O(gate83inter8));
  nand2 gate696(.a(gate83inter8), .b(gate83inter7), .O(gate83inter9));
  nand2 gate697(.a(s_21), .b(gate83inter3), .O(gate83inter10));
  nor2  gate698(.a(gate83inter10), .b(gate83inter9), .O(gate83inter11));
  nor2  gate699(.a(gate83inter11), .b(gate83inter6), .O(gate83inter12));
  nand2 gate700(.a(gate83inter12), .b(gate83inter1), .O(G404));
nand2 gate84( .a(G15), .b(G329), .O(G405) );
nand2 gate85( .a(G4), .b(G332), .O(G406) );
nand2 gate86( .a(G8), .b(G332), .O(G407) );
nand2 gate87( .a(G12), .b(G335), .O(G408) );

  xor2  gate1219(.a(G335), .b(G16), .O(gate88inter0));
  nand2 gate1220(.a(gate88inter0), .b(s_96), .O(gate88inter1));
  and2  gate1221(.a(G335), .b(G16), .O(gate88inter2));
  inv1  gate1222(.a(s_96), .O(gate88inter3));
  inv1  gate1223(.a(s_97), .O(gate88inter4));
  nand2 gate1224(.a(gate88inter4), .b(gate88inter3), .O(gate88inter5));
  nor2  gate1225(.a(gate88inter5), .b(gate88inter2), .O(gate88inter6));
  inv1  gate1226(.a(G16), .O(gate88inter7));
  inv1  gate1227(.a(G335), .O(gate88inter8));
  nand2 gate1228(.a(gate88inter8), .b(gate88inter7), .O(gate88inter9));
  nand2 gate1229(.a(s_97), .b(gate88inter3), .O(gate88inter10));
  nor2  gate1230(.a(gate88inter10), .b(gate88inter9), .O(gate88inter11));
  nor2  gate1231(.a(gate88inter11), .b(gate88inter6), .O(gate88inter12));
  nand2 gate1232(.a(gate88inter12), .b(gate88inter1), .O(G409));
nand2 gate89( .a(G17), .b(G338), .O(G410) );
nand2 gate90( .a(G21), .b(G338), .O(G411) );
nand2 gate91( .a(G25), .b(G341), .O(G412) );
nand2 gate92( .a(G29), .b(G341), .O(G413) );

  xor2  gate953(.a(G344), .b(G18), .O(gate93inter0));
  nand2 gate954(.a(gate93inter0), .b(s_58), .O(gate93inter1));
  and2  gate955(.a(G344), .b(G18), .O(gate93inter2));
  inv1  gate956(.a(s_58), .O(gate93inter3));
  inv1  gate957(.a(s_59), .O(gate93inter4));
  nand2 gate958(.a(gate93inter4), .b(gate93inter3), .O(gate93inter5));
  nor2  gate959(.a(gate93inter5), .b(gate93inter2), .O(gate93inter6));
  inv1  gate960(.a(G18), .O(gate93inter7));
  inv1  gate961(.a(G344), .O(gate93inter8));
  nand2 gate962(.a(gate93inter8), .b(gate93inter7), .O(gate93inter9));
  nand2 gate963(.a(s_59), .b(gate93inter3), .O(gate93inter10));
  nor2  gate964(.a(gate93inter10), .b(gate93inter9), .O(gate93inter11));
  nor2  gate965(.a(gate93inter11), .b(gate93inter6), .O(gate93inter12));
  nand2 gate966(.a(gate93inter12), .b(gate93inter1), .O(G414));
nand2 gate94( .a(G22), .b(G344), .O(G415) );

  xor2  gate659(.a(G347), .b(G26), .O(gate95inter0));
  nand2 gate660(.a(gate95inter0), .b(s_16), .O(gate95inter1));
  and2  gate661(.a(G347), .b(G26), .O(gate95inter2));
  inv1  gate662(.a(s_16), .O(gate95inter3));
  inv1  gate663(.a(s_17), .O(gate95inter4));
  nand2 gate664(.a(gate95inter4), .b(gate95inter3), .O(gate95inter5));
  nor2  gate665(.a(gate95inter5), .b(gate95inter2), .O(gate95inter6));
  inv1  gate666(.a(G26), .O(gate95inter7));
  inv1  gate667(.a(G347), .O(gate95inter8));
  nand2 gate668(.a(gate95inter8), .b(gate95inter7), .O(gate95inter9));
  nand2 gate669(.a(s_17), .b(gate95inter3), .O(gate95inter10));
  nor2  gate670(.a(gate95inter10), .b(gate95inter9), .O(gate95inter11));
  nor2  gate671(.a(gate95inter11), .b(gate95inter6), .O(gate95inter12));
  nand2 gate672(.a(gate95inter12), .b(gate95inter1), .O(G416));

  xor2  gate1513(.a(G347), .b(G30), .O(gate96inter0));
  nand2 gate1514(.a(gate96inter0), .b(s_138), .O(gate96inter1));
  and2  gate1515(.a(G347), .b(G30), .O(gate96inter2));
  inv1  gate1516(.a(s_138), .O(gate96inter3));
  inv1  gate1517(.a(s_139), .O(gate96inter4));
  nand2 gate1518(.a(gate96inter4), .b(gate96inter3), .O(gate96inter5));
  nor2  gate1519(.a(gate96inter5), .b(gate96inter2), .O(gate96inter6));
  inv1  gate1520(.a(G30), .O(gate96inter7));
  inv1  gate1521(.a(G347), .O(gate96inter8));
  nand2 gate1522(.a(gate96inter8), .b(gate96inter7), .O(gate96inter9));
  nand2 gate1523(.a(s_139), .b(gate96inter3), .O(gate96inter10));
  nor2  gate1524(.a(gate96inter10), .b(gate96inter9), .O(gate96inter11));
  nor2  gate1525(.a(gate96inter11), .b(gate96inter6), .O(gate96inter12));
  nand2 gate1526(.a(gate96inter12), .b(gate96inter1), .O(G417));
nand2 gate97( .a(G19), .b(G350), .O(G418) );

  xor2  gate1009(.a(G350), .b(G23), .O(gate98inter0));
  nand2 gate1010(.a(gate98inter0), .b(s_66), .O(gate98inter1));
  and2  gate1011(.a(G350), .b(G23), .O(gate98inter2));
  inv1  gate1012(.a(s_66), .O(gate98inter3));
  inv1  gate1013(.a(s_67), .O(gate98inter4));
  nand2 gate1014(.a(gate98inter4), .b(gate98inter3), .O(gate98inter5));
  nor2  gate1015(.a(gate98inter5), .b(gate98inter2), .O(gate98inter6));
  inv1  gate1016(.a(G23), .O(gate98inter7));
  inv1  gate1017(.a(G350), .O(gate98inter8));
  nand2 gate1018(.a(gate98inter8), .b(gate98inter7), .O(gate98inter9));
  nand2 gate1019(.a(s_67), .b(gate98inter3), .O(gate98inter10));
  nor2  gate1020(.a(gate98inter10), .b(gate98inter9), .O(gate98inter11));
  nor2  gate1021(.a(gate98inter11), .b(gate98inter6), .O(gate98inter12));
  nand2 gate1022(.a(gate98inter12), .b(gate98inter1), .O(G419));
nand2 gate99( .a(G27), .b(G353), .O(G420) );
nand2 gate100( .a(G31), .b(G353), .O(G421) );
nand2 gate101( .a(G20), .b(G356), .O(G422) );
nand2 gate102( .a(G24), .b(G356), .O(G423) );
nand2 gate103( .a(G28), .b(G359), .O(G424) );
nand2 gate104( .a(G32), .b(G359), .O(G425) );
nand2 gate105( .a(G362), .b(G363), .O(G426) );
nand2 gate106( .a(G364), .b(G365), .O(G429) );
nand2 gate107( .a(G366), .b(G367), .O(G432) );
nand2 gate108( .a(G368), .b(G369), .O(G435) );
nand2 gate109( .a(G370), .b(G371), .O(G438) );

  xor2  gate1387(.a(G373), .b(G372), .O(gate110inter0));
  nand2 gate1388(.a(gate110inter0), .b(s_120), .O(gate110inter1));
  and2  gate1389(.a(G373), .b(G372), .O(gate110inter2));
  inv1  gate1390(.a(s_120), .O(gate110inter3));
  inv1  gate1391(.a(s_121), .O(gate110inter4));
  nand2 gate1392(.a(gate110inter4), .b(gate110inter3), .O(gate110inter5));
  nor2  gate1393(.a(gate110inter5), .b(gate110inter2), .O(gate110inter6));
  inv1  gate1394(.a(G372), .O(gate110inter7));
  inv1  gate1395(.a(G373), .O(gate110inter8));
  nand2 gate1396(.a(gate110inter8), .b(gate110inter7), .O(gate110inter9));
  nand2 gate1397(.a(s_121), .b(gate110inter3), .O(gate110inter10));
  nor2  gate1398(.a(gate110inter10), .b(gate110inter9), .O(gate110inter11));
  nor2  gate1399(.a(gate110inter11), .b(gate110inter6), .O(gate110inter12));
  nand2 gate1400(.a(gate110inter12), .b(gate110inter1), .O(G441));
nand2 gate111( .a(G374), .b(G375), .O(G444) );
nand2 gate112( .a(G376), .b(G377), .O(G447) );
nand2 gate113( .a(G378), .b(G379), .O(G450) );

  xor2  gate1331(.a(G381), .b(G380), .O(gate114inter0));
  nand2 gate1332(.a(gate114inter0), .b(s_112), .O(gate114inter1));
  and2  gate1333(.a(G381), .b(G380), .O(gate114inter2));
  inv1  gate1334(.a(s_112), .O(gate114inter3));
  inv1  gate1335(.a(s_113), .O(gate114inter4));
  nand2 gate1336(.a(gate114inter4), .b(gate114inter3), .O(gate114inter5));
  nor2  gate1337(.a(gate114inter5), .b(gate114inter2), .O(gate114inter6));
  inv1  gate1338(.a(G380), .O(gate114inter7));
  inv1  gate1339(.a(G381), .O(gate114inter8));
  nand2 gate1340(.a(gate114inter8), .b(gate114inter7), .O(gate114inter9));
  nand2 gate1341(.a(s_113), .b(gate114inter3), .O(gate114inter10));
  nor2  gate1342(.a(gate114inter10), .b(gate114inter9), .O(gate114inter11));
  nor2  gate1343(.a(gate114inter11), .b(gate114inter6), .O(gate114inter12));
  nand2 gate1344(.a(gate114inter12), .b(gate114inter1), .O(G453));
nand2 gate115( .a(G382), .b(G383), .O(G456) );
nand2 gate116( .a(G384), .b(G385), .O(G459) );
nand2 gate117( .a(G386), .b(G387), .O(G462) );
nand2 gate118( .a(G388), .b(G389), .O(G465) );
nand2 gate119( .a(G390), .b(G391), .O(G468) );

  xor2  gate1485(.a(G393), .b(G392), .O(gate120inter0));
  nand2 gate1486(.a(gate120inter0), .b(s_134), .O(gate120inter1));
  and2  gate1487(.a(G393), .b(G392), .O(gate120inter2));
  inv1  gate1488(.a(s_134), .O(gate120inter3));
  inv1  gate1489(.a(s_135), .O(gate120inter4));
  nand2 gate1490(.a(gate120inter4), .b(gate120inter3), .O(gate120inter5));
  nor2  gate1491(.a(gate120inter5), .b(gate120inter2), .O(gate120inter6));
  inv1  gate1492(.a(G392), .O(gate120inter7));
  inv1  gate1493(.a(G393), .O(gate120inter8));
  nand2 gate1494(.a(gate120inter8), .b(gate120inter7), .O(gate120inter9));
  nand2 gate1495(.a(s_135), .b(gate120inter3), .O(gate120inter10));
  nor2  gate1496(.a(gate120inter10), .b(gate120inter9), .O(gate120inter11));
  nor2  gate1497(.a(gate120inter11), .b(gate120inter6), .O(gate120inter12));
  nand2 gate1498(.a(gate120inter12), .b(gate120inter1), .O(G471));

  xor2  gate757(.a(G395), .b(G394), .O(gate121inter0));
  nand2 gate758(.a(gate121inter0), .b(s_30), .O(gate121inter1));
  and2  gate759(.a(G395), .b(G394), .O(gate121inter2));
  inv1  gate760(.a(s_30), .O(gate121inter3));
  inv1  gate761(.a(s_31), .O(gate121inter4));
  nand2 gate762(.a(gate121inter4), .b(gate121inter3), .O(gate121inter5));
  nor2  gate763(.a(gate121inter5), .b(gate121inter2), .O(gate121inter6));
  inv1  gate764(.a(G394), .O(gate121inter7));
  inv1  gate765(.a(G395), .O(gate121inter8));
  nand2 gate766(.a(gate121inter8), .b(gate121inter7), .O(gate121inter9));
  nand2 gate767(.a(s_31), .b(gate121inter3), .O(gate121inter10));
  nor2  gate768(.a(gate121inter10), .b(gate121inter9), .O(gate121inter11));
  nor2  gate769(.a(gate121inter11), .b(gate121inter6), .O(gate121inter12));
  nand2 gate770(.a(gate121inter12), .b(gate121inter1), .O(G474));
nand2 gate122( .a(G396), .b(G397), .O(G477) );
nand2 gate123( .a(G398), .b(G399), .O(G480) );

  xor2  gate1093(.a(G401), .b(G400), .O(gate124inter0));
  nand2 gate1094(.a(gate124inter0), .b(s_78), .O(gate124inter1));
  and2  gate1095(.a(G401), .b(G400), .O(gate124inter2));
  inv1  gate1096(.a(s_78), .O(gate124inter3));
  inv1  gate1097(.a(s_79), .O(gate124inter4));
  nand2 gate1098(.a(gate124inter4), .b(gate124inter3), .O(gate124inter5));
  nor2  gate1099(.a(gate124inter5), .b(gate124inter2), .O(gate124inter6));
  inv1  gate1100(.a(G400), .O(gate124inter7));
  inv1  gate1101(.a(G401), .O(gate124inter8));
  nand2 gate1102(.a(gate124inter8), .b(gate124inter7), .O(gate124inter9));
  nand2 gate1103(.a(s_79), .b(gate124inter3), .O(gate124inter10));
  nor2  gate1104(.a(gate124inter10), .b(gate124inter9), .O(gate124inter11));
  nor2  gate1105(.a(gate124inter11), .b(gate124inter6), .O(gate124inter12));
  nand2 gate1106(.a(gate124inter12), .b(gate124inter1), .O(G483));

  xor2  gate1443(.a(G403), .b(G402), .O(gate125inter0));
  nand2 gate1444(.a(gate125inter0), .b(s_128), .O(gate125inter1));
  and2  gate1445(.a(G403), .b(G402), .O(gate125inter2));
  inv1  gate1446(.a(s_128), .O(gate125inter3));
  inv1  gate1447(.a(s_129), .O(gate125inter4));
  nand2 gate1448(.a(gate125inter4), .b(gate125inter3), .O(gate125inter5));
  nor2  gate1449(.a(gate125inter5), .b(gate125inter2), .O(gate125inter6));
  inv1  gate1450(.a(G402), .O(gate125inter7));
  inv1  gate1451(.a(G403), .O(gate125inter8));
  nand2 gate1452(.a(gate125inter8), .b(gate125inter7), .O(gate125inter9));
  nand2 gate1453(.a(s_129), .b(gate125inter3), .O(gate125inter10));
  nor2  gate1454(.a(gate125inter10), .b(gate125inter9), .O(gate125inter11));
  nor2  gate1455(.a(gate125inter11), .b(gate125inter6), .O(gate125inter12));
  nand2 gate1456(.a(gate125inter12), .b(gate125inter1), .O(G486));

  xor2  gate1457(.a(G405), .b(G404), .O(gate126inter0));
  nand2 gate1458(.a(gate126inter0), .b(s_130), .O(gate126inter1));
  and2  gate1459(.a(G405), .b(G404), .O(gate126inter2));
  inv1  gate1460(.a(s_130), .O(gate126inter3));
  inv1  gate1461(.a(s_131), .O(gate126inter4));
  nand2 gate1462(.a(gate126inter4), .b(gate126inter3), .O(gate126inter5));
  nor2  gate1463(.a(gate126inter5), .b(gate126inter2), .O(gate126inter6));
  inv1  gate1464(.a(G404), .O(gate126inter7));
  inv1  gate1465(.a(G405), .O(gate126inter8));
  nand2 gate1466(.a(gate126inter8), .b(gate126inter7), .O(gate126inter9));
  nand2 gate1467(.a(s_131), .b(gate126inter3), .O(gate126inter10));
  nor2  gate1468(.a(gate126inter10), .b(gate126inter9), .O(gate126inter11));
  nor2  gate1469(.a(gate126inter11), .b(gate126inter6), .O(gate126inter12));
  nand2 gate1470(.a(gate126inter12), .b(gate126inter1), .O(G489));
nand2 gate127( .a(G406), .b(G407), .O(G492) );
nand2 gate128( .a(G408), .b(G409), .O(G495) );

  xor2  gate785(.a(G411), .b(G410), .O(gate129inter0));
  nand2 gate786(.a(gate129inter0), .b(s_34), .O(gate129inter1));
  and2  gate787(.a(G411), .b(G410), .O(gate129inter2));
  inv1  gate788(.a(s_34), .O(gate129inter3));
  inv1  gate789(.a(s_35), .O(gate129inter4));
  nand2 gate790(.a(gate129inter4), .b(gate129inter3), .O(gate129inter5));
  nor2  gate791(.a(gate129inter5), .b(gate129inter2), .O(gate129inter6));
  inv1  gate792(.a(G410), .O(gate129inter7));
  inv1  gate793(.a(G411), .O(gate129inter8));
  nand2 gate794(.a(gate129inter8), .b(gate129inter7), .O(gate129inter9));
  nand2 gate795(.a(s_35), .b(gate129inter3), .O(gate129inter10));
  nor2  gate796(.a(gate129inter10), .b(gate129inter9), .O(gate129inter11));
  nor2  gate797(.a(gate129inter11), .b(gate129inter6), .O(gate129inter12));
  nand2 gate798(.a(gate129inter12), .b(gate129inter1), .O(G498));

  xor2  gate1359(.a(G413), .b(G412), .O(gate130inter0));
  nand2 gate1360(.a(gate130inter0), .b(s_116), .O(gate130inter1));
  and2  gate1361(.a(G413), .b(G412), .O(gate130inter2));
  inv1  gate1362(.a(s_116), .O(gate130inter3));
  inv1  gate1363(.a(s_117), .O(gate130inter4));
  nand2 gate1364(.a(gate130inter4), .b(gate130inter3), .O(gate130inter5));
  nor2  gate1365(.a(gate130inter5), .b(gate130inter2), .O(gate130inter6));
  inv1  gate1366(.a(G412), .O(gate130inter7));
  inv1  gate1367(.a(G413), .O(gate130inter8));
  nand2 gate1368(.a(gate130inter8), .b(gate130inter7), .O(gate130inter9));
  nand2 gate1369(.a(s_117), .b(gate130inter3), .O(gate130inter10));
  nor2  gate1370(.a(gate130inter10), .b(gate130inter9), .O(gate130inter11));
  nor2  gate1371(.a(gate130inter11), .b(gate130inter6), .O(gate130inter12));
  nand2 gate1372(.a(gate130inter12), .b(gate130inter1), .O(G501));
nand2 gate131( .a(G414), .b(G415), .O(G504) );
nand2 gate132( .a(G416), .b(G417), .O(G507) );
nand2 gate133( .a(G418), .b(G419), .O(G510) );
nand2 gate134( .a(G420), .b(G421), .O(G513) );
nand2 gate135( .a(G422), .b(G423), .O(G516) );
nand2 gate136( .a(G424), .b(G425), .O(G519) );
nand2 gate137( .a(G426), .b(G429), .O(G522) );
nand2 gate138( .a(G432), .b(G435), .O(G525) );
nand2 gate139( .a(G438), .b(G441), .O(G528) );

  xor2  gate1555(.a(G447), .b(G444), .O(gate140inter0));
  nand2 gate1556(.a(gate140inter0), .b(s_144), .O(gate140inter1));
  and2  gate1557(.a(G447), .b(G444), .O(gate140inter2));
  inv1  gate1558(.a(s_144), .O(gate140inter3));
  inv1  gate1559(.a(s_145), .O(gate140inter4));
  nand2 gate1560(.a(gate140inter4), .b(gate140inter3), .O(gate140inter5));
  nor2  gate1561(.a(gate140inter5), .b(gate140inter2), .O(gate140inter6));
  inv1  gate1562(.a(G444), .O(gate140inter7));
  inv1  gate1563(.a(G447), .O(gate140inter8));
  nand2 gate1564(.a(gate140inter8), .b(gate140inter7), .O(gate140inter9));
  nand2 gate1565(.a(s_145), .b(gate140inter3), .O(gate140inter10));
  nor2  gate1566(.a(gate140inter10), .b(gate140inter9), .O(gate140inter11));
  nor2  gate1567(.a(gate140inter11), .b(gate140inter6), .O(gate140inter12));
  nand2 gate1568(.a(gate140inter12), .b(gate140inter1), .O(G531));
nand2 gate141( .a(G450), .b(G453), .O(G534) );
nand2 gate142( .a(G456), .b(G459), .O(G537) );
nand2 gate143( .a(G462), .b(G465), .O(G540) );
nand2 gate144( .a(G468), .b(G471), .O(G543) );
nand2 gate145( .a(G474), .b(G477), .O(G546) );
nand2 gate146( .a(G480), .b(G483), .O(G549) );
nand2 gate147( .a(G486), .b(G489), .O(G552) );
nand2 gate148( .a(G492), .b(G495), .O(G555) );
nand2 gate149( .a(G498), .b(G501), .O(G558) );
nand2 gate150( .a(G504), .b(G507), .O(G561) );

  xor2  gate827(.a(G513), .b(G510), .O(gate151inter0));
  nand2 gate828(.a(gate151inter0), .b(s_40), .O(gate151inter1));
  and2  gate829(.a(G513), .b(G510), .O(gate151inter2));
  inv1  gate830(.a(s_40), .O(gate151inter3));
  inv1  gate831(.a(s_41), .O(gate151inter4));
  nand2 gate832(.a(gate151inter4), .b(gate151inter3), .O(gate151inter5));
  nor2  gate833(.a(gate151inter5), .b(gate151inter2), .O(gate151inter6));
  inv1  gate834(.a(G510), .O(gate151inter7));
  inv1  gate835(.a(G513), .O(gate151inter8));
  nand2 gate836(.a(gate151inter8), .b(gate151inter7), .O(gate151inter9));
  nand2 gate837(.a(s_41), .b(gate151inter3), .O(gate151inter10));
  nor2  gate838(.a(gate151inter10), .b(gate151inter9), .O(gate151inter11));
  nor2  gate839(.a(gate151inter11), .b(gate151inter6), .O(gate151inter12));
  nand2 gate840(.a(gate151inter12), .b(gate151inter1), .O(G564));
nand2 gate152( .a(G516), .b(G519), .O(G567) );
nand2 gate153( .a(G426), .b(G522), .O(G570) );
nand2 gate154( .a(G429), .b(G522), .O(G571) );
nand2 gate155( .a(G432), .b(G525), .O(G572) );
nand2 gate156( .a(G435), .b(G525), .O(G573) );
nand2 gate157( .a(G438), .b(G528), .O(G574) );
nand2 gate158( .a(G441), .b(G528), .O(G575) );
nand2 gate159( .a(G444), .b(G531), .O(G576) );
nand2 gate160( .a(G447), .b(G531), .O(G577) );
nand2 gate161( .a(G450), .b(G534), .O(G578) );
nand2 gate162( .a(G453), .b(G534), .O(G579) );
nand2 gate163( .a(G456), .b(G537), .O(G580) );
nand2 gate164( .a(G459), .b(G537), .O(G581) );
nand2 gate165( .a(G462), .b(G540), .O(G582) );

  xor2  gate1373(.a(G540), .b(G465), .O(gate166inter0));
  nand2 gate1374(.a(gate166inter0), .b(s_118), .O(gate166inter1));
  and2  gate1375(.a(G540), .b(G465), .O(gate166inter2));
  inv1  gate1376(.a(s_118), .O(gate166inter3));
  inv1  gate1377(.a(s_119), .O(gate166inter4));
  nand2 gate1378(.a(gate166inter4), .b(gate166inter3), .O(gate166inter5));
  nor2  gate1379(.a(gate166inter5), .b(gate166inter2), .O(gate166inter6));
  inv1  gate1380(.a(G465), .O(gate166inter7));
  inv1  gate1381(.a(G540), .O(gate166inter8));
  nand2 gate1382(.a(gate166inter8), .b(gate166inter7), .O(gate166inter9));
  nand2 gate1383(.a(s_119), .b(gate166inter3), .O(gate166inter10));
  nor2  gate1384(.a(gate166inter10), .b(gate166inter9), .O(gate166inter11));
  nor2  gate1385(.a(gate166inter11), .b(gate166inter6), .O(gate166inter12));
  nand2 gate1386(.a(gate166inter12), .b(gate166inter1), .O(G583));

  xor2  gate1275(.a(G543), .b(G468), .O(gate167inter0));
  nand2 gate1276(.a(gate167inter0), .b(s_104), .O(gate167inter1));
  and2  gate1277(.a(G543), .b(G468), .O(gate167inter2));
  inv1  gate1278(.a(s_104), .O(gate167inter3));
  inv1  gate1279(.a(s_105), .O(gate167inter4));
  nand2 gate1280(.a(gate167inter4), .b(gate167inter3), .O(gate167inter5));
  nor2  gate1281(.a(gate167inter5), .b(gate167inter2), .O(gate167inter6));
  inv1  gate1282(.a(G468), .O(gate167inter7));
  inv1  gate1283(.a(G543), .O(gate167inter8));
  nand2 gate1284(.a(gate167inter8), .b(gate167inter7), .O(gate167inter9));
  nand2 gate1285(.a(s_105), .b(gate167inter3), .O(gate167inter10));
  nor2  gate1286(.a(gate167inter10), .b(gate167inter9), .O(gate167inter11));
  nor2  gate1287(.a(gate167inter11), .b(gate167inter6), .O(gate167inter12));
  nand2 gate1288(.a(gate167inter12), .b(gate167inter1), .O(G584));
nand2 gate168( .a(G471), .b(G543), .O(G585) );
nand2 gate169( .a(G474), .b(G546), .O(G586) );
nand2 gate170( .a(G477), .b(G546), .O(G587) );
nand2 gate171( .a(G480), .b(G549), .O(G588) );
nand2 gate172( .a(G483), .b(G549), .O(G589) );
nand2 gate173( .a(G486), .b(G552), .O(G590) );
nand2 gate174( .a(G489), .b(G552), .O(G591) );
nand2 gate175( .a(G492), .b(G555), .O(G592) );
nand2 gate176( .a(G495), .b(G555), .O(G593) );
nand2 gate177( .a(G498), .b(G558), .O(G594) );
nand2 gate178( .a(G501), .b(G558), .O(G595) );
nand2 gate179( .a(G504), .b(G561), .O(G596) );
nand2 gate180( .a(G507), .b(G561), .O(G597) );
nand2 gate181( .a(G510), .b(G564), .O(G598) );
nand2 gate182( .a(G513), .b(G564), .O(G599) );
nand2 gate183( .a(G516), .b(G567), .O(G600) );
nand2 gate184( .a(G519), .b(G567), .O(G601) );

  xor2  gate1303(.a(G571), .b(G570), .O(gate185inter0));
  nand2 gate1304(.a(gate185inter0), .b(s_108), .O(gate185inter1));
  and2  gate1305(.a(G571), .b(G570), .O(gate185inter2));
  inv1  gate1306(.a(s_108), .O(gate185inter3));
  inv1  gate1307(.a(s_109), .O(gate185inter4));
  nand2 gate1308(.a(gate185inter4), .b(gate185inter3), .O(gate185inter5));
  nor2  gate1309(.a(gate185inter5), .b(gate185inter2), .O(gate185inter6));
  inv1  gate1310(.a(G570), .O(gate185inter7));
  inv1  gate1311(.a(G571), .O(gate185inter8));
  nand2 gate1312(.a(gate185inter8), .b(gate185inter7), .O(gate185inter9));
  nand2 gate1313(.a(s_109), .b(gate185inter3), .O(gate185inter10));
  nor2  gate1314(.a(gate185inter10), .b(gate185inter9), .O(gate185inter11));
  nor2  gate1315(.a(gate185inter11), .b(gate185inter6), .O(gate185inter12));
  nand2 gate1316(.a(gate185inter12), .b(gate185inter1), .O(G602));
nand2 gate186( .a(G572), .b(G573), .O(G607) );
nand2 gate187( .a(G574), .b(G575), .O(G612) );
nand2 gate188( .a(G576), .b(G577), .O(G617) );

  xor2  gate1191(.a(G579), .b(G578), .O(gate189inter0));
  nand2 gate1192(.a(gate189inter0), .b(s_92), .O(gate189inter1));
  and2  gate1193(.a(G579), .b(G578), .O(gate189inter2));
  inv1  gate1194(.a(s_92), .O(gate189inter3));
  inv1  gate1195(.a(s_93), .O(gate189inter4));
  nand2 gate1196(.a(gate189inter4), .b(gate189inter3), .O(gate189inter5));
  nor2  gate1197(.a(gate189inter5), .b(gate189inter2), .O(gate189inter6));
  inv1  gate1198(.a(G578), .O(gate189inter7));
  inv1  gate1199(.a(G579), .O(gate189inter8));
  nand2 gate1200(.a(gate189inter8), .b(gate189inter7), .O(gate189inter9));
  nand2 gate1201(.a(s_93), .b(gate189inter3), .O(gate189inter10));
  nor2  gate1202(.a(gate189inter10), .b(gate189inter9), .O(gate189inter11));
  nor2  gate1203(.a(gate189inter11), .b(gate189inter6), .O(gate189inter12));
  nand2 gate1204(.a(gate189inter12), .b(gate189inter1), .O(G622));

  xor2  gate701(.a(G581), .b(G580), .O(gate190inter0));
  nand2 gate702(.a(gate190inter0), .b(s_22), .O(gate190inter1));
  and2  gate703(.a(G581), .b(G580), .O(gate190inter2));
  inv1  gate704(.a(s_22), .O(gate190inter3));
  inv1  gate705(.a(s_23), .O(gate190inter4));
  nand2 gate706(.a(gate190inter4), .b(gate190inter3), .O(gate190inter5));
  nor2  gate707(.a(gate190inter5), .b(gate190inter2), .O(gate190inter6));
  inv1  gate708(.a(G580), .O(gate190inter7));
  inv1  gate709(.a(G581), .O(gate190inter8));
  nand2 gate710(.a(gate190inter8), .b(gate190inter7), .O(gate190inter9));
  nand2 gate711(.a(s_23), .b(gate190inter3), .O(gate190inter10));
  nor2  gate712(.a(gate190inter10), .b(gate190inter9), .O(gate190inter11));
  nor2  gate713(.a(gate190inter11), .b(gate190inter6), .O(gate190inter12));
  nand2 gate714(.a(gate190inter12), .b(gate190inter1), .O(G627));
nand2 gate191( .a(G582), .b(G583), .O(G632) );
nand2 gate192( .a(G584), .b(G585), .O(G637) );
nand2 gate193( .a(G586), .b(G587), .O(G642) );
nand2 gate194( .a(G588), .b(G589), .O(G645) );
nand2 gate195( .a(G590), .b(G591), .O(G648) );

  xor2  gate855(.a(G593), .b(G592), .O(gate196inter0));
  nand2 gate856(.a(gate196inter0), .b(s_44), .O(gate196inter1));
  and2  gate857(.a(G593), .b(G592), .O(gate196inter2));
  inv1  gate858(.a(s_44), .O(gate196inter3));
  inv1  gate859(.a(s_45), .O(gate196inter4));
  nand2 gate860(.a(gate196inter4), .b(gate196inter3), .O(gate196inter5));
  nor2  gate861(.a(gate196inter5), .b(gate196inter2), .O(gate196inter6));
  inv1  gate862(.a(G592), .O(gate196inter7));
  inv1  gate863(.a(G593), .O(gate196inter8));
  nand2 gate864(.a(gate196inter8), .b(gate196inter7), .O(gate196inter9));
  nand2 gate865(.a(s_45), .b(gate196inter3), .O(gate196inter10));
  nor2  gate866(.a(gate196inter10), .b(gate196inter9), .O(gate196inter11));
  nor2  gate867(.a(gate196inter11), .b(gate196inter6), .O(gate196inter12));
  nand2 gate868(.a(gate196inter12), .b(gate196inter1), .O(G651));
nand2 gate197( .a(G594), .b(G595), .O(G654) );
nand2 gate198( .a(G596), .b(G597), .O(G657) );
nand2 gate199( .a(G598), .b(G599), .O(G660) );
nand2 gate200( .a(G600), .b(G601), .O(G663) );
nand2 gate201( .a(G602), .b(G607), .O(G666) );
nand2 gate202( .a(G612), .b(G617), .O(G669) );
nand2 gate203( .a(G602), .b(G612), .O(G672) );
nand2 gate204( .a(G607), .b(G617), .O(G675) );
nand2 gate205( .a(G622), .b(G627), .O(G678) );
nand2 gate206( .a(G632), .b(G637), .O(G681) );
nand2 gate207( .a(G622), .b(G632), .O(G684) );
nand2 gate208( .a(G627), .b(G637), .O(G687) );
nand2 gate209( .a(G602), .b(G666), .O(G690) );
nand2 gate210( .a(G607), .b(G666), .O(G691) );

  xor2  gate1163(.a(G669), .b(G612), .O(gate211inter0));
  nand2 gate1164(.a(gate211inter0), .b(s_88), .O(gate211inter1));
  and2  gate1165(.a(G669), .b(G612), .O(gate211inter2));
  inv1  gate1166(.a(s_88), .O(gate211inter3));
  inv1  gate1167(.a(s_89), .O(gate211inter4));
  nand2 gate1168(.a(gate211inter4), .b(gate211inter3), .O(gate211inter5));
  nor2  gate1169(.a(gate211inter5), .b(gate211inter2), .O(gate211inter6));
  inv1  gate1170(.a(G612), .O(gate211inter7));
  inv1  gate1171(.a(G669), .O(gate211inter8));
  nand2 gate1172(.a(gate211inter8), .b(gate211inter7), .O(gate211inter9));
  nand2 gate1173(.a(s_89), .b(gate211inter3), .O(gate211inter10));
  nor2  gate1174(.a(gate211inter10), .b(gate211inter9), .O(gate211inter11));
  nor2  gate1175(.a(gate211inter11), .b(gate211inter6), .O(gate211inter12));
  nand2 gate1176(.a(gate211inter12), .b(gate211inter1), .O(G692));
nand2 gate212( .a(G617), .b(G669), .O(G693) );
nand2 gate213( .a(G602), .b(G672), .O(G694) );
nand2 gate214( .a(G612), .b(G672), .O(G695) );

  xor2  gate743(.a(G675), .b(G607), .O(gate215inter0));
  nand2 gate744(.a(gate215inter0), .b(s_28), .O(gate215inter1));
  and2  gate745(.a(G675), .b(G607), .O(gate215inter2));
  inv1  gate746(.a(s_28), .O(gate215inter3));
  inv1  gate747(.a(s_29), .O(gate215inter4));
  nand2 gate748(.a(gate215inter4), .b(gate215inter3), .O(gate215inter5));
  nor2  gate749(.a(gate215inter5), .b(gate215inter2), .O(gate215inter6));
  inv1  gate750(.a(G607), .O(gate215inter7));
  inv1  gate751(.a(G675), .O(gate215inter8));
  nand2 gate752(.a(gate215inter8), .b(gate215inter7), .O(gate215inter9));
  nand2 gate753(.a(s_29), .b(gate215inter3), .O(gate215inter10));
  nor2  gate754(.a(gate215inter10), .b(gate215inter9), .O(gate215inter11));
  nor2  gate755(.a(gate215inter11), .b(gate215inter6), .O(gate215inter12));
  nand2 gate756(.a(gate215inter12), .b(gate215inter1), .O(G696));
nand2 gate216( .a(G617), .b(G675), .O(G697) );

  xor2  gate841(.a(G678), .b(G622), .O(gate217inter0));
  nand2 gate842(.a(gate217inter0), .b(s_42), .O(gate217inter1));
  and2  gate843(.a(G678), .b(G622), .O(gate217inter2));
  inv1  gate844(.a(s_42), .O(gate217inter3));
  inv1  gate845(.a(s_43), .O(gate217inter4));
  nand2 gate846(.a(gate217inter4), .b(gate217inter3), .O(gate217inter5));
  nor2  gate847(.a(gate217inter5), .b(gate217inter2), .O(gate217inter6));
  inv1  gate848(.a(G622), .O(gate217inter7));
  inv1  gate849(.a(G678), .O(gate217inter8));
  nand2 gate850(.a(gate217inter8), .b(gate217inter7), .O(gate217inter9));
  nand2 gate851(.a(s_43), .b(gate217inter3), .O(gate217inter10));
  nor2  gate852(.a(gate217inter10), .b(gate217inter9), .O(gate217inter11));
  nor2  gate853(.a(gate217inter11), .b(gate217inter6), .O(gate217inter12));
  nand2 gate854(.a(gate217inter12), .b(gate217inter1), .O(G698));
nand2 gate218( .a(G627), .b(G678), .O(G699) );
nand2 gate219( .a(G632), .b(G681), .O(G700) );
nand2 gate220( .a(G637), .b(G681), .O(G701) );
nand2 gate221( .a(G622), .b(G684), .O(G702) );
nand2 gate222( .a(G632), .b(G684), .O(G703) );
nand2 gate223( .a(G627), .b(G687), .O(G704) );
nand2 gate224( .a(G637), .b(G687), .O(G705) );

  xor2  gate771(.a(G691), .b(G690), .O(gate225inter0));
  nand2 gate772(.a(gate225inter0), .b(s_32), .O(gate225inter1));
  and2  gate773(.a(G691), .b(G690), .O(gate225inter2));
  inv1  gate774(.a(s_32), .O(gate225inter3));
  inv1  gate775(.a(s_33), .O(gate225inter4));
  nand2 gate776(.a(gate225inter4), .b(gate225inter3), .O(gate225inter5));
  nor2  gate777(.a(gate225inter5), .b(gate225inter2), .O(gate225inter6));
  inv1  gate778(.a(G690), .O(gate225inter7));
  inv1  gate779(.a(G691), .O(gate225inter8));
  nand2 gate780(.a(gate225inter8), .b(gate225inter7), .O(gate225inter9));
  nand2 gate781(.a(s_33), .b(gate225inter3), .O(gate225inter10));
  nor2  gate782(.a(gate225inter10), .b(gate225inter9), .O(gate225inter11));
  nor2  gate783(.a(gate225inter11), .b(gate225inter6), .O(gate225inter12));
  nand2 gate784(.a(gate225inter12), .b(gate225inter1), .O(G706));
nand2 gate226( .a(G692), .b(G693), .O(G709) );
nand2 gate227( .a(G694), .b(G695), .O(G712) );

  xor2  gate1051(.a(G697), .b(G696), .O(gate228inter0));
  nand2 gate1052(.a(gate228inter0), .b(s_72), .O(gate228inter1));
  and2  gate1053(.a(G697), .b(G696), .O(gate228inter2));
  inv1  gate1054(.a(s_72), .O(gate228inter3));
  inv1  gate1055(.a(s_73), .O(gate228inter4));
  nand2 gate1056(.a(gate228inter4), .b(gate228inter3), .O(gate228inter5));
  nor2  gate1057(.a(gate228inter5), .b(gate228inter2), .O(gate228inter6));
  inv1  gate1058(.a(G696), .O(gate228inter7));
  inv1  gate1059(.a(G697), .O(gate228inter8));
  nand2 gate1060(.a(gate228inter8), .b(gate228inter7), .O(gate228inter9));
  nand2 gate1061(.a(s_73), .b(gate228inter3), .O(gate228inter10));
  nor2  gate1062(.a(gate228inter10), .b(gate228inter9), .O(gate228inter11));
  nor2  gate1063(.a(gate228inter11), .b(gate228inter6), .O(gate228inter12));
  nand2 gate1064(.a(gate228inter12), .b(gate228inter1), .O(G715));

  xor2  gate631(.a(G699), .b(G698), .O(gate229inter0));
  nand2 gate632(.a(gate229inter0), .b(s_12), .O(gate229inter1));
  and2  gate633(.a(G699), .b(G698), .O(gate229inter2));
  inv1  gate634(.a(s_12), .O(gate229inter3));
  inv1  gate635(.a(s_13), .O(gate229inter4));
  nand2 gate636(.a(gate229inter4), .b(gate229inter3), .O(gate229inter5));
  nor2  gate637(.a(gate229inter5), .b(gate229inter2), .O(gate229inter6));
  inv1  gate638(.a(G698), .O(gate229inter7));
  inv1  gate639(.a(G699), .O(gate229inter8));
  nand2 gate640(.a(gate229inter8), .b(gate229inter7), .O(gate229inter9));
  nand2 gate641(.a(s_13), .b(gate229inter3), .O(gate229inter10));
  nor2  gate642(.a(gate229inter10), .b(gate229inter9), .O(gate229inter11));
  nor2  gate643(.a(gate229inter11), .b(gate229inter6), .O(gate229inter12));
  nand2 gate644(.a(gate229inter12), .b(gate229inter1), .O(G718));

  xor2  gate1289(.a(G701), .b(G700), .O(gate230inter0));
  nand2 gate1290(.a(gate230inter0), .b(s_106), .O(gate230inter1));
  and2  gate1291(.a(G701), .b(G700), .O(gate230inter2));
  inv1  gate1292(.a(s_106), .O(gate230inter3));
  inv1  gate1293(.a(s_107), .O(gate230inter4));
  nand2 gate1294(.a(gate230inter4), .b(gate230inter3), .O(gate230inter5));
  nor2  gate1295(.a(gate230inter5), .b(gate230inter2), .O(gate230inter6));
  inv1  gate1296(.a(G700), .O(gate230inter7));
  inv1  gate1297(.a(G701), .O(gate230inter8));
  nand2 gate1298(.a(gate230inter8), .b(gate230inter7), .O(gate230inter9));
  nand2 gate1299(.a(s_107), .b(gate230inter3), .O(gate230inter10));
  nor2  gate1300(.a(gate230inter10), .b(gate230inter9), .O(gate230inter11));
  nor2  gate1301(.a(gate230inter11), .b(gate230inter6), .O(gate230inter12));
  nand2 gate1302(.a(gate230inter12), .b(gate230inter1), .O(G721));

  xor2  gate869(.a(G703), .b(G702), .O(gate231inter0));
  nand2 gate870(.a(gate231inter0), .b(s_46), .O(gate231inter1));
  and2  gate871(.a(G703), .b(G702), .O(gate231inter2));
  inv1  gate872(.a(s_46), .O(gate231inter3));
  inv1  gate873(.a(s_47), .O(gate231inter4));
  nand2 gate874(.a(gate231inter4), .b(gate231inter3), .O(gate231inter5));
  nor2  gate875(.a(gate231inter5), .b(gate231inter2), .O(gate231inter6));
  inv1  gate876(.a(G702), .O(gate231inter7));
  inv1  gate877(.a(G703), .O(gate231inter8));
  nand2 gate878(.a(gate231inter8), .b(gate231inter7), .O(gate231inter9));
  nand2 gate879(.a(s_47), .b(gate231inter3), .O(gate231inter10));
  nor2  gate880(.a(gate231inter10), .b(gate231inter9), .O(gate231inter11));
  nor2  gate881(.a(gate231inter11), .b(gate231inter6), .O(gate231inter12));
  nand2 gate882(.a(gate231inter12), .b(gate231inter1), .O(G724));
nand2 gate232( .a(G704), .b(G705), .O(G727) );
nand2 gate233( .a(G242), .b(G718), .O(G730) );
nand2 gate234( .a(G245), .b(G721), .O(G733) );
nand2 gate235( .a(G248), .b(G724), .O(G736) );
nand2 gate236( .a(G251), .b(G727), .O(G739) );
nand2 gate237( .a(G254), .b(G706), .O(G742) );
nand2 gate238( .a(G257), .b(G709), .O(G745) );
nand2 gate239( .a(G260), .b(G712), .O(G748) );
nand2 gate240( .a(G263), .b(G715), .O(G751) );
nand2 gate241( .a(G242), .b(G730), .O(G754) );

  xor2  gate547(.a(G730), .b(G718), .O(gate242inter0));
  nand2 gate548(.a(gate242inter0), .b(s_0), .O(gate242inter1));
  and2  gate549(.a(G730), .b(G718), .O(gate242inter2));
  inv1  gate550(.a(s_0), .O(gate242inter3));
  inv1  gate551(.a(s_1), .O(gate242inter4));
  nand2 gate552(.a(gate242inter4), .b(gate242inter3), .O(gate242inter5));
  nor2  gate553(.a(gate242inter5), .b(gate242inter2), .O(gate242inter6));
  inv1  gate554(.a(G718), .O(gate242inter7));
  inv1  gate555(.a(G730), .O(gate242inter8));
  nand2 gate556(.a(gate242inter8), .b(gate242inter7), .O(gate242inter9));
  nand2 gate557(.a(s_1), .b(gate242inter3), .O(gate242inter10));
  nor2  gate558(.a(gate242inter10), .b(gate242inter9), .O(gate242inter11));
  nor2  gate559(.a(gate242inter11), .b(gate242inter6), .O(gate242inter12));
  nand2 gate560(.a(gate242inter12), .b(gate242inter1), .O(G755));

  xor2  gate561(.a(G733), .b(G245), .O(gate243inter0));
  nand2 gate562(.a(gate243inter0), .b(s_2), .O(gate243inter1));
  and2  gate563(.a(G733), .b(G245), .O(gate243inter2));
  inv1  gate564(.a(s_2), .O(gate243inter3));
  inv1  gate565(.a(s_3), .O(gate243inter4));
  nand2 gate566(.a(gate243inter4), .b(gate243inter3), .O(gate243inter5));
  nor2  gate567(.a(gate243inter5), .b(gate243inter2), .O(gate243inter6));
  inv1  gate568(.a(G245), .O(gate243inter7));
  inv1  gate569(.a(G733), .O(gate243inter8));
  nand2 gate570(.a(gate243inter8), .b(gate243inter7), .O(gate243inter9));
  nand2 gate571(.a(s_3), .b(gate243inter3), .O(gate243inter10));
  nor2  gate572(.a(gate243inter10), .b(gate243inter9), .O(gate243inter11));
  nor2  gate573(.a(gate243inter11), .b(gate243inter6), .O(gate243inter12));
  nand2 gate574(.a(gate243inter12), .b(gate243inter1), .O(G756));
nand2 gate244( .a(G721), .b(G733), .O(G757) );
nand2 gate245( .a(G248), .b(G736), .O(G758) );
nand2 gate246( .a(G724), .b(G736), .O(G759) );
nand2 gate247( .a(G251), .b(G739), .O(G760) );
nand2 gate248( .a(G727), .b(G739), .O(G761) );

  xor2  gate575(.a(G742), .b(G254), .O(gate249inter0));
  nand2 gate576(.a(gate249inter0), .b(s_4), .O(gate249inter1));
  and2  gate577(.a(G742), .b(G254), .O(gate249inter2));
  inv1  gate578(.a(s_4), .O(gate249inter3));
  inv1  gate579(.a(s_5), .O(gate249inter4));
  nand2 gate580(.a(gate249inter4), .b(gate249inter3), .O(gate249inter5));
  nor2  gate581(.a(gate249inter5), .b(gate249inter2), .O(gate249inter6));
  inv1  gate582(.a(G254), .O(gate249inter7));
  inv1  gate583(.a(G742), .O(gate249inter8));
  nand2 gate584(.a(gate249inter8), .b(gate249inter7), .O(gate249inter9));
  nand2 gate585(.a(s_5), .b(gate249inter3), .O(gate249inter10));
  nor2  gate586(.a(gate249inter10), .b(gate249inter9), .O(gate249inter11));
  nor2  gate587(.a(gate249inter11), .b(gate249inter6), .O(gate249inter12));
  nand2 gate588(.a(gate249inter12), .b(gate249inter1), .O(G762));
nand2 gate250( .a(G706), .b(G742), .O(G763) );
nand2 gate251( .a(G257), .b(G745), .O(G764) );
nand2 gate252( .a(G709), .b(G745), .O(G765) );
nand2 gate253( .a(G260), .b(G748), .O(G766) );
nand2 gate254( .a(G712), .b(G748), .O(G767) );
nand2 gate255( .a(G263), .b(G751), .O(G768) );
nand2 gate256( .a(G715), .b(G751), .O(G769) );
nand2 gate257( .a(G754), .b(G755), .O(G770) );
nand2 gate258( .a(G756), .b(G757), .O(G773) );
nand2 gate259( .a(G758), .b(G759), .O(G776) );
nand2 gate260( .a(G760), .b(G761), .O(G779) );
nand2 gate261( .a(G762), .b(G763), .O(G782) );
nand2 gate262( .a(G764), .b(G765), .O(G785) );
nand2 gate263( .a(G766), .b(G767), .O(G788) );
nand2 gate264( .a(G768), .b(G769), .O(G791) );
nand2 gate265( .a(G642), .b(G770), .O(G794) );
nand2 gate266( .a(G645), .b(G773), .O(G797) );
nand2 gate267( .a(G648), .b(G776), .O(G800) );
nand2 gate268( .a(G651), .b(G779), .O(G803) );

  xor2  gate1121(.a(G782), .b(G654), .O(gate269inter0));
  nand2 gate1122(.a(gate269inter0), .b(s_82), .O(gate269inter1));
  and2  gate1123(.a(G782), .b(G654), .O(gate269inter2));
  inv1  gate1124(.a(s_82), .O(gate269inter3));
  inv1  gate1125(.a(s_83), .O(gate269inter4));
  nand2 gate1126(.a(gate269inter4), .b(gate269inter3), .O(gate269inter5));
  nor2  gate1127(.a(gate269inter5), .b(gate269inter2), .O(gate269inter6));
  inv1  gate1128(.a(G654), .O(gate269inter7));
  inv1  gate1129(.a(G782), .O(gate269inter8));
  nand2 gate1130(.a(gate269inter8), .b(gate269inter7), .O(gate269inter9));
  nand2 gate1131(.a(s_83), .b(gate269inter3), .O(gate269inter10));
  nor2  gate1132(.a(gate269inter10), .b(gate269inter9), .O(gate269inter11));
  nor2  gate1133(.a(gate269inter11), .b(gate269inter6), .O(gate269inter12));
  nand2 gate1134(.a(gate269inter12), .b(gate269inter1), .O(G806));
nand2 gate270( .a(G657), .b(G785), .O(G809) );
nand2 gate271( .a(G660), .b(G788), .O(G812) );
nand2 gate272( .a(G663), .b(G791), .O(G815) );
nand2 gate273( .a(G642), .b(G794), .O(G818) );
nand2 gate274( .a(G770), .b(G794), .O(G819) );
nand2 gate275( .a(G645), .b(G797), .O(G820) );
nand2 gate276( .a(G773), .b(G797), .O(G821) );
nand2 gate277( .a(G648), .b(G800), .O(G822) );
nand2 gate278( .a(G776), .b(G800), .O(G823) );
nand2 gate279( .a(G651), .b(G803), .O(G824) );
nand2 gate280( .a(G779), .b(G803), .O(G825) );
nand2 gate281( .a(G654), .b(G806), .O(G826) );
nand2 gate282( .a(G782), .b(G806), .O(G827) );
nand2 gate283( .a(G657), .b(G809), .O(G828) );
nand2 gate284( .a(G785), .b(G809), .O(G829) );
nand2 gate285( .a(G660), .b(G812), .O(G830) );
nand2 gate286( .a(G788), .b(G812), .O(G831) );
nand2 gate287( .a(G663), .b(G815), .O(G832) );
nand2 gate288( .a(G791), .b(G815), .O(G833) );
nand2 gate289( .a(G818), .b(G819), .O(G834) );
nand2 gate290( .a(G820), .b(G821), .O(G847) );
nand2 gate291( .a(G822), .b(G823), .O(G860) );
nand2 gate292( .a(G824), .b(G825), .O(G873) );
nand2 gate293( .a(G828), .b(G829), .O(G886) );
nand2 gate294( .a(G832), .b(G833), .O(G899) );
nand2 gate295( .a(G830), .b(G831), .O(G912) );
nand2 gate296( .a(G826), .b(G827), .O(G925) );
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );

  xor2  gate1597(.a(G1036), .b(G1), .O(gate387inter0));
  nand2 gate1598(.a(gate387inter0), .b(s_150), .O(gate387inter1));
  and2  gate1599(.a(G1036), .b(G1), .O(gate387inter2));
  inv1  gate1600(.a(s_150), .O(gate387inter3));
  inv1  gate1601(.a(s_151), .O(gate387inter4));
  nand2 gate1602(.a(gate387inter4), .b(gate387inter3), .O(gate387inter5));
  nor2  gate1603(.a(gate387inter5), .b(gate387inter2), .O(gate387inter6));
  inv1  gate1604(.a(G1), .O(gate387inter7));
  inv1  gate1605(.a(G1036), .O(gate387inter8));
  nand2 gate1606(.a(gate387inter8), .b(gate387inter7), .O(gate387inter9));
  nand2 gate1607(.a(s_151), .b(gate387inter3), .O(gate387inter10));
  nor2  gate1608(.a(gate387inter10), .b(gate387inter9), .O(gate387inter11));
  nor2  gate1609(.a(gate387inter11), .b(gate387inter6), .O(gate387inter12));
  nand2 gate1610(.a(gate387inter12), .b(gate387inter1), .O(G1132));
nand2 gate388( .a(G2), .b(G1039), .O(G1135) );
nand2 gate389( .a(G3), .b(G1042), .O(G1138) );

  xor2  gate1023(.a(G1045), .b(G4), .O(gate390inter0));
  nand2 gate1024(.a(gate390inter0), .b(s_68), .O(gate390inter1));
  and2  gate1025(.a(G1045), .b(G4), .O(gate390inter2));
  inv1  gate1026(.a(s_68), .O(gate390inter3));
  inv1  gate1027(.a(s_69), .O(gate390inter4));
  nand2 gate1028(.a(gate390inter4), .b(gate390inter3), .O(gate390inter5));
  nor2  gate1029(.a(gate390inter5), .b(gate390inter2), .O(gate390inter6));
  inv1  gate1030(.a(G4), .O(gate390inter7));
  inv1  gate1031(.a(G1045), .O(gate390inter8));
  nand2 gate1032(.a(gate390inter8), .b(gate390inter7), .O(gate390inter9));
  nand2 gate1033(.a(s_69), .b(gate390inter3), .O(gate390inter10));
  nor2  gate1034(.a(gate390inter10), .b(gate390inter9), .O(gate390inter11));
  nor2  gate1035(.a(gate390inter11), .b(gate390inter6), .O(gate390inter12));
  nand2 gate1036(.a(gate390inter12), .b(gate390inter1), .O(G1141));
nand2 gate391( .a(G5), .b(G1048), .O(G1144) );
nand2 gate392( .a(G6), .b(G1051), .O(G1147) );
nand2 gate393( .a(G7), .b(G1054), .O(G1150) );
nand2 gate394( .a(G8), .b(G1057), .O(G1153) );
nand2 gate395( .a(G9), .b(G1060), .O(G1156) );
nand2 gate396( .a(G10), .b(G1063), .O(G1159) );
nand2 gate397( .a(G11), .b(G1066), .O(G1162) );
nand2 gate398( .a(G12), .b(G1069), .O(G1165) );
nand2 gate399( .a(G13), .b(G1072), .O(G1168) );
nand2 gate400( .a(G14), .b(G1075), .O(G1171) );
nand2 gate401( .a(G15), .b(G1078), .O(G1174) );
nand2 gate402( .a(G16), .b(G1081), .O(G1177) );
nand2 gate403( .a(G17), .b(G1084), .O(G1180) );
nand2 gate404( .a(G18), .b(G1087), .O(G1183) );
nand2 gate405( .a(G19), .b(G1090), .O(G1186) );
nand2 gate406( .a(G20), .b(G1093), .O(G1189) );
nand2 gate407( .a(G21), .b(G1096), .O(G1192) );
nand2 gate408( .a(G22), .b(G1099), .O(G1195) );
nand2 gate409( .a(G23), .b(G1102), .O(G1198) );
nand2 gate410( .a(G24), .b(G1105), .O(G1201) );
nand2 gate411( .a(G25), .b(G1108), .O(G1204) );
nand2 gate412( .a(G26), .b(G1111), .O(G1207) );
nand2 gate413( .a(G27), .b(G1114), .O(G1210) );
nand2 gate414( .a(G28), .b(G1117), .O(G1213) );

  xor2  gate1135(.a(G1120), .b(G29), .O(gate415inter0));
  nand2 gate1136(.a(gate415inter0), .b(s_84), .O(gate415inter1));
  and2  gate1137(.a(G1120), .b(G29), .O(gate415inter2));
  inv1  gate1138(.a(s_84), .O(gate415inter3));
  inv1  gate1139(.a(s_85), .O(gate415inter4));
  nand2 gate1140(.a(gate415inter4), .b(gate415inter3), .O(gate415inter5));
  nor2  gate1141(.a(gate415inter5), .b(gate415inter2), .O(gate415inter6));
  inv1  gate1142(.a(G29), .O(gate415inter7));
  inv1  gate1143(.a(G1120), .O(gate415inter8));
  nand2 gate1144(.a(gate415inter8), .b(gate415inter7), .O(gate415inter9));
  nand2 gate1145(.a(s_85), .b(gate415inter3), .O(gate415inter10));
  nor2  gate1146(.a(gate415inter10), .b(gate415inter9), .O(gate415inter11));
  nor2  gate1147(.a(gate415inter11), .b(gate415inter6), .O(gate415inter12));
  nand2 gate1148(.a(gate415inter12), .b(gate415inter1), .O(G1216));
nand2 gate416( .a(G30), .b(G1123), .O(G1219) );
nand2 gate417( .a(G31), .b(G1126), .O(G1222) );
nand2 gate418( .a(G32), .b(G1129), .O(G1225) );
nand2 gate419( .a(G1), .b(G1132), .O(G1228) );
nand2 gate420( .a(G1036), .b(G1132), .O(G1229) );
nand2 gate421( .a(G2), .b(G1135), .O(G1230) );
nand2 gate422( .a(G1039), .b(G1135), .O(G1231) );

  xor2  gate981(.a(G1138), .b(G3), .O(gate423inter0));
  nand2 gate982(.a(gate423inter0), .b(s_62), .O(gate423inter1));
  and2  gate983(.a(G1138), .b(G3), .O(gate423inter2));
  inv1  gate984(.a(s_62), .O(gate423inter3));
  inv1  gate985(.a(s_63), .O(gate423inter4));
  nand2 gate986(.a(gate423inter4), .b(gate423inter3), .O(gate423inter5));
  nor2  gate987(.a(gate423inter5), .b(gate423inter2), .O(gate423inter6));
  inv1  gate988(.a(G3), .O(gate423inter7));
  inv1  gate989(.a(G1138), .O(gate423inter8));
  nand2 gate990(.a(gate423inter8), .b(gate423inter7), .O(gate423inter9));
  nand2 gate991(.a(s_63), .b(gate423inter3), .O(gate423inter10));
  nor2  gate992(.a(gate423inter10), .b(gate423inter9), .O(gate423inter11));
  nor2  gate993(.a(gate423inter11), .b(gate423inter6), .O(gate423inter12));
  nand2 gate994(.a(gate423inter12), .b(gate423inter1), .O(G1232));
nand2 gate424( .a(G1042), .b(G1138), .O(G1233) );
nand2 gate425( .a(G4), .b(G1141), .O(G1234) );
nand2 gate426( .a(G1045), .b(G1141), .O(G1235) );
nand2 gate427( .a(G5), .b(G1144), .O(G1236) );
nand2 gate428( .a(G1048), .b(G1144), .O(G1237) );
nand2 gate429( .a(G6), .b(G1147), .O(G1238) );
nand2 gate430( .a(G1051), .b(G1147), .O(G1239) );
nand2 gate431( .a(G7), .b(G1150), .O(G1240) );
nand2 gate432( .a(G1054), .b(G1150), .O(G1241) );
nand2 gate433( .a(G8), .b(G1153), .O(G1242) );

  xor2  gate1499(.a(G1153), .b(G1057), .O(gate434inter0));
  nand2 gate1500(.a(gate434inter0), .b(s_136), .O(gate434inter1));
  and2  gate1501(.a(G1153), .b(G1057), .O(gate434inter2));
  inv1  gate1502(.a(s_136), .O(gate434inter3));
  inv1  gate1503(.a(s_137), .O(gate434inter4));
  nand2 gate1504(.a(gate434inter4), .b(gate434inter3), .O(gate434inter5));
  nor2  gate1505(.a(gate434inter5), .b(gate434inter2), .O(gate434inter6));
  inv1  gate1506(.a(G1057), .O(gate434inter7));
  inv1  gate1507(.a(G1153), .O(gate434inter8));
  nand2 gate1508(.a(gate434inter8), .b(gate434inter7), .O(gate434inter9));
  nand2 gate1509(.a(s_137), .b(gate434inter3), .O(gate434inter10));
  nor2  gate1510(.a(gate434inter10), .b(gate434inter9), .O(gate434inter11));
  nor2  gate1511(.a(gate434inter11), .b(gate434inter6), .O(gate434inter12));
  nand2 gate1512(.a(gate434inter12), .b(gate434inter1), .O(G1243));
nand2 gate435( .a(G9), .b(G1156), .O(G1244) );
nand2 gate436( .a(G1060), .b(G1156), .O(G1245) );
nand2 gate437( .a(G10), .b(G1159), .O(G1246) );
nand2 gate438( .a(G1063), .b(G1159), .O(G1247) );
nand2 gate439( .a(G11), .b(G1162), .O(G1248) );
nand2 gate440( .a(G1066), .b(G1162), .O(G1249) );

  xor2  gate1471(.a(G1165), .b(G12), .O(gate441inter0));
  nand2 gate1472(.a(gate441inter0), .b(s_132), .O(gate441inter1));
  and2  gate1473(.a(G1165), .b(G12), .O(gate441inter2));
  inv1  gate1474(.a(s_132), .O(gate441inter3));
  inv1  gate1475(.a(s_133), .O(gate441inter4));
  nand2 gate1476(.a(gate441inter4), .b(gate441inter3), .O(gate441inter5));
  nor2  gate1477(.a(gate441inter5), .b(gate441inter2), .O(gate441inter6));
  inv1  gate1478(.a(G12), .O(gate441inter7));
  inv1  gate1479(.a(G1165), .O(gate441inter8));
  nand2 gate1480(.a(gate441inter8), .b(gate441inter7), .O(gate441inter9));
  nand2 gate1481(.a(s_133), .b(gate441inter3), .O(gate441inter10));
  nor2  gate1482(.a(gate441inter10), .b(gate441inter9), .O(gate441inter11));
  nor2  gate1483(.a(gate441inter11), .b(gate441inter6), .O(gate441inter12));
  nand2 gate1484(.a(gate441inter12), .b(gate441inter1), .O(G1250));
nand2 gate442( .a(G1069), .b(G1165), .O(G1251) );
nand2 gate443( .a(G13), .b(G1168), .O(G1252) );

  xor2  gate1149(.a(G1168), .b(G1072), .O(gate444inter0));
  nand2 gate1150(.a(gate444inter0), .b(s_86), .O(gate444inter1));
  and2  gate1151(.a(G1168), .b(G1072), .O(gate444inter2));
  inv1  gate1152(.a(s_86), .O(gate444inter3));
  inv1  gate1153(.a(s_87), .O(gate444inter4));
  nand2 gate1154(.a(gate444inter4), .b(gate444inter3), .O(gate444inter5));
  nor2  gate1155(.a(gate444inter5), .b(gate444inter2), .O(gate444inter6));
  inv1  gate1156(.a(G1072), .O(gate444inter7));
  inv1  gate1157(.a(G1168), .O(gate444inter8));
  nand2 gate1158(.a(gate444inter8), .b(gate444inter7), .O(gate444inter9));
  nand2 gate1159(.a(s_87), .b(gate444inter3), .O(gate444inter10));
  nor2  gate1160(.a(gate444inter10), .b(gate444inter9), .O(gate444inter11));
  nor2  gate1161(.a(gate444inter11), .b(gate444inter6), .O(gate444inter12));
  nand2 gate1162(.a(gate444inter12), .b(gate444inter1), .O(G1253));
nand2 gate445( .a(G14), .b(G1171), .O(G1254) );
nand2 gate446( .a(G1075), .b(G1171), .O(G1255) );
nand2 gate447( .a(G15), .b(G1174), .O(G1256) );
nand2 gate448( .a(G1078), .b(G1174), .O(G1257) );
nand2 gate449( .a(G16), .b(G1177), .O(G1258) );
nand2 gate450( .a(G1081), .b(G1177), .O(G1259) );
nand2 gate451( .a(G17), .b(G1180), .O(G1260) );

  xor2  gate799(.a(G1180), .b(G1084), .O(gate452inter0));
  nand2 gate800(.a(gate452inter0), .b(s_36), .O(gate452inter1));
  and2  gate801(.a(G1180), .b(G1084), .O(gate452inter2));
  inv1  gate802(.a(s_36), .O(gate452inter3));
  inv1  gate803(.a(s_37), .O(gate452inter4));
  nand2 gate804(.a(gate452inter4), .b(gate452inter3), .O(gate452inter5));
  nor2  gate805(.a(gate452inter5), .b(gate452inter2), .O(gate452inter6));
  inv1  gate806(.a(G1084), .O(gate452inter7));
  inv1  gate807(.a(G1180), .O(gate452inter8));
  nand2 gate808(.a(gate452inter8), .b(gate452inter7), .O(gate452inter9));
  nand2 gate809(.a(s_37), .b(gate452inter3), .O(gate452inter10));
  nor2  gate810(.a(gate452inter10), .b(gate452inter9), .O(gate452inter11));
  nor2  gate811(.a(gate452inter11), .b(gate452inter6), .O(gate452inter12));
  nand2 gate812(.a(gate452inter12), .b(gate452inter1), .O(G1261));
nand2 gate453( .a(G18), .b(G1183), .O(G1262) );

  xor2  gate673(.a(G1183), .b(G1087), .O(gate454inter0));
  nand2 gate674(.a(gate454inter0), .b(s_18), .O(gate454inter1));
  and2  gate675(.a(G1183), .b(G1087), .O(gate454inter2));
  inv1  gate676(.a(s_18), .O(gate454inter3));
  inv1  gate677(.a(s_19), .O(gate454inter4));
  nand2 gate678(.a(gate454inter4), .b(gate454inter3), .O(gate454inter5));
  nor2  gate679(.a(gate454inter5), .b(gate454inter2), .O(gate454inter6));
  inv1  gate680(.a(G1087), .O(gate454inter7));
  inv1  gate681(.a(G1183), .O(gate454inter8));
  nand2 gate682(.a(gate454inter8), .b(gate454inter7), .O(gate454inter9));
  nand2 gate683(.a(s_19), .b(gate454inter3), .O(gate454inter10));
  nor2  gate684(.a(gate454inter10), .b(gate454inter9), .O(gate454inter11));
  nor2  gate685(.a(gate454inter11), .b(gate454inter6), .O(gate454inter12));
  nand2 gate686(.a(gate454inter12), .b(gate454inter1), .O(G1263));

  xor2  gate1415(.a(G1186), .b(G19), .O(gate455inter0));
  nand2 gate1416(.a(gate455inter0), .b(s_124), .O(gate455inter1));
  and2  gate1417(.a(G1186), .b(G19), .O(gate455inter2));
  inv1  gate1418(.a(s_124), .O(gate455inter3));
  inv1  gate1419(.a(s_125), .O(gate455inter4));
  nand2 gate1420(.a(gate455inter4), .b(gate455inter3), .O(gate455inter5));
  nor2  gate1421(.a(gate455inter5), .b(gate455inter2), .O(gate455inter6));
  inv1  gate1422(.a(G19), .O(gate455inter7));
  inv1  gate1423(.a(G1186), .O(gate455inter8));
  nand2 gate1424(.a(gate455inter8), .b(gate455inter7), .O(gate455inter9));
  nand2 gate1425(.a(s_125), .b(gate455inter3), .O(gate455inter10));
  nor2  gate1426(.a(gate455inter10), .b(gate455inter9), .O(gate455inter11));
  nor2  gate1427(.a(gate455inter11), .b(gate455inter6), .O(gate455inter12));
  nand2 gate1428(.a(gate455inter12), .b(gate455inter1), .O(G1264));
nand2 gate456( .a(G1090), .b(G1186), .O(G1265) );
nand2 gate457( .a(G20), .b(G1189), .O(G1266) );

  xor2  gate1247(.a(G1189), .b(G1093), .O(gate458inter0));
  nand2 gate1248(.a(gate458inter0), .b(s_100), .O(gate458inter1));
  and2  gate1249(.a(G1189), .b(G1093), .O(gate458inter2));
  inv1  gate1250(.a(s_100), .O(gate458inter3));
  inv1  gate1251(.a(s_101), .O(gate458inter4));
  nand2 gate1252(.a(gate458inter4), .b(gate458inter3), .O(gate458inter5));
  nor2  gate1253(.a(gate458inter5), .b(gate458inter2), .O(gate458inter6));
  inv1  gate1254(.a(G1093), .O(gate458inter7));
  inv1  gate1255(.a(G1189), .O(gate458inter8));
  nand2 gate1256(.a(gate458inter8), .b(gate458inter7), .O(gate458inter9));
  nand2 gate1257(.a(s_101), .b(gate458inter3), .O(gate458inter10));
  nor2  gate1258(.a(gate458inter10), .b(gate458inter9), .O(gate458inter11));
  nor2  gate1259(.a(gate458inter11), .b(gate458inter6), .O(gate458inter12));
  nand2 gate1260(.a(gate458inter12), .b(gate458inter1), .O(G1267));

  xor2  gate1037(.a(G1192), .b(G21), .O(gate459inter0));
  nand2 gate1038(.a(gate459inter0), .b(s_70), .O(gate459inter1));
  and2  gate1039(.a(G1192), .b(G21), .O(gate459inter2));
  inv1  gate1040(.a(s_70), .O(gate459inter3));
  inv1  gate1041(.a(s_71), .O(gate459inter4));
  nand2 gate1042(.a(gate459inter4), .b(gate459inter3), .O(gate459inter5));
  nor2  gate1043(.a(gate459inter5), .b(gate459inter2), .O(gate459inter6));
  inv1  gate1044(.a(G21), .O(gate459inter7));
  inv1  gate1045(.a(G1192), .O(gate459inter8));
  nand2 gate1046(.a(gate459inter8), .b(gate459inter7), .O(gate459inter9));
  nand2 gate1047(.a(s_71), .b(gate459inter3), .O(gate459inter10));
  nor2  gate1048(.a(gate459inter10), .b(gate459inter9), .O(gate459inter11));
  nor2  gate1049(.a(gate459inter11), .b(gate459inter6), .O(gate459inter12));
  nand2 gate1050(.a(gate459inter12), .b(gate459inter1), .O(G1268));
nand2 gate460( .a(G1096), .b(G1192), .O(G1269) );

  xor2  gate715(.a(G1195), .b(G22), .O(gate461inter0));
  nand2 gate716(.a(gate461inter0), .b(s_24), .O(gate461inter1));
  and2  gate717(.a(G1195), .b(G22), .O(gate461inter2));
  inv1  gate718(.a(s_24), .O(gate461inter3));
  inv1  gate719(.a(s_25), .O(gate461inter4));
  nand2 gate720(.a(gate461inter4), .b(gate461inter3), .O(gate461inter5));
  nor2  gate721(.a(gate461inter5), .b(gate461inter2), .O(gate461inter6));
  inv1  gate722(.a(G22), .O(gate461inter7));
  inv1  gate723(.a(G1195), .O(gate461inter8));
  nand2 gate724(.a(gate461inter8), .b(gate461inter7), .O(gate461inter9));
  nand2 gate725(.a(s_25), .b(gate461inter3), .O(gate461inter10));
  nor2  gate726(.a(gate461inter10), .b(gate461inter9), .O(gate461inter11));
  nor2  gate727(.a(gate461inter11), .b(gate461inter6), .O(gate461inter12));
  nand2 gate728(.a(gate461inter12), .b(gate461inter1), .O(G1270));
nand2 gate462( .a(G1099), .b(G1195), .O(G1271) );
nand2 gate463( .a(G23), .b(G1198), .O(G1272) );
nand2 gate464( .a(G1102), .b(G1198), .O(G1273) );
nand2 gate465( .a(G24), .b(G1201), .O(G1274) );

  xor2  gate589(.a(G1201), .b(G1105), .O(gate466inter0));
  nand2 gate590(.a(gate466inter0), .b(s_6), .O(gate466inter1));
  and2  gate591(.a(G1201), .b(G1105), .O(gate466inter2));
  inv1  gate592(.a(s_6), .O(gate466inter3));
  inv1  gate593(.a(s_7), .O(gate466inter4));
  nand2 gate594(.a(gate466inter4), .b(gate466inter3), .O(gate466inter5));
  nor2  gate595(.a(gate466inter5), .b(gate466inter2), .O(gate466inter6));
  inv1  gate596(.a(G1105), .O(gate466inter7));
  inv1  gate597(.a(G1201), .O(gate466inter8));
  nand2 gate598(.a(gate466inter8), .b(gate466inter7), .O(gate466inter9));
  nand2 gate599(.a(s_7), .b(gate466inter3), .O(gate466inter10));
  nor2  gate600(.a(gate466inter10), .b(gate466inter9), .O(gate466inter11));
  nor2  gate601(.a(gate466inter11), .b(gate466inter6), .O(gate466inter12));
  nand2 gate602(.a(gate466inter12), .b(gate466inter1), .O(G1275));
nand2 gate467( .a(G25), .b(G1204), .O(G1276) );
nand2 gate468( .a(G1108), .b(G1204), .O(G1277) );
nand2 gate469( .a(G26), .b(G1207), .O(G1278) );
nand2 gate470( .a(G1111), .b(G1207), .O(G1279) );

  xor2  gate1065(.a(G1210), .b(G27), .O(gate471inter0));
  nand2 gate1066(.a(gate471inter0), .b(s_74), .O(gate471inter1));
  and2  gate1067(.a(G1210), .b(G27), .O(gate471inter2));
  inv1  gate1068(.a(s_74), .O(gate471inter3));
  inv1  gate1069(.a(s_75), .O(gate471inter4));
  nand2 gate1070(.a(gate471inter4), .b(gate471inter3), .O(gate471inter5));
  nor2  gate1071(.a(gate471inter5), .b(gate471inter2), .O(gate471inter6));
  inv1  gate1072(.a(G27), .O(gate471inter7));
  inv1  gate1073(.a(G1210), .O(gate471inter8));
  nand2 gate1074(.a(gate471inter8), .b(gate471inter7), .O(gate471inter9));
  nand2 gate1075(.a(s_75), .b(gate471inter3), .O(gate471inter10));
  nor2  gate1076(.a(gate471inter10), .b(gate471inter9), .O(gate471inter11));
  nor2  gate1077(.a(gate471inter11), .b(gate471inter6), .O(gate471inter12));
  nand2 gate1078(.a(gate471inter12), .b(gate471inter1), .O(G1280));
nand2 gate472( .a(G1114), .b(G1210), .O(G1281) );
nand2 gate473( .a(G28), .b(G1213), .O(G1282) );
nand2 gate474( .a(G1117), .b(G1213), .O(G1283) );

  xor2  gate995(.a(G1216), .b(G29), .O(gate475inter0));
  nand2 gate996(.a(gate475inter0), .b(s_64), .O(gate475inter1));
  and2  gate997(.a(G1216), .b(G29), .O(gate475inter2));
  inv1  gate998(.a(s_64), .O(gate475inter3));
  inv1  gate999(.a(s_65), .O(gate475inter4));
  nand2 gate1000(.a(gate475inter4), .b(gate475inter3), .O(gate475inter5));
  nor2  gate1001(.a(gate475inter5), .b(gate475inter2), .O(gate475inter6));
  inv1  gate1002(.a(G29), .O(gate475inter7));
  inv1  gate1003(.a(G1216), .O(gate475inter8));
  nand2 gate1004(.a(gate475inter8), .b(gate475inter7), .O(gate475inter9));
  nand2 gate1005(.a(s_65), .b(gate475inter3), .O(gate475inter10));
  nor2  gate1006(.a(gate475inter10), .b(gate475inter9), .O(gate475inter11));
  nor2  gate1007(.a(gate475inter11), .b(gate475inter6), .O(gate475inter12));
  nand2 gate1008(.a(gate475inter12), .b(gate475inter1), .O(G1284));
nand2 gate476( .a(G1120), .b(G1216), .O(G1285) );
nand2 gate477( .a(G30), .b(G1219), .O(G1286) );
nand2 gate478( .a(G1123), .b(G1219), .O(G1287) );
nand2 gate479( .a(G31), .b(G1222), .O(G1288) );
nand2 gate480( .a(G1126), .b(G1222), .O(G1289) );

  xor2  gate1569(.a(G1225), .b(G32), .O(gate481inter0));
  nand2 gate1570(.a(gate481inter0), .b(s_146), .O(gate481inter1));
  and2  gate1571(.a(G1225), .b(G32), .O(gate481inter2));
  inv1  gate1572(.a(s_146), .O(gate481inter3));
  inv1  gate1573(.a(s_147), .O(gate481inter4));
  nand2 gate1574(.a(gate481inter4), .b(gate481inter3), .O(gate481inter5));
  nor2  gate1575(.a(gate481inter5), .b(gate481inter2), .O(gate481inter6));
  inv1  gate1576(.a(G32), .O(gate481inter7));
  inv1  gate1577(.a(G1225), .O(gate481inter8));
  nand2 gate1578(.a(gate481inter8), .b(gate481inter7), .O(gate481inter9));
  nand2 gate1579(.a(s_147), .b(gate481inter3), .O(gate481inter10));
  nor2  gate1580(.a(gate481inter10), .b(gate481inter9), .O(gate481inter11));
  nor2  gate1581(.a(gate481inter11), .b(gate481inter6), .O(gate481inter12));
  nand2 gate1582(.a(gate481inter12), .b(gate481inter1), .O(G1290));

  xor2  gate925(.a(G1225), .b(G1129), .O(gate482inter0));
  nand2 gate926(.a(gate482inter0), .b(s_54), .O(gate482inter1));
  and2  gate927(.a(G1225), .b(G1129), .O(gate482inter2));
  inv1  gate928(.a(s_54), .O(gate482inter3));
  inv1  gate929(.a(s_55), .O(gate482inter4));
  nand2 gate930(.a(gate482inter4), .b(gate482inter3), .O(gate482inter5));
  nor2  gate931(.a(gate482inter5), .b(gate482inter2), .O(gate482inter6));
  inv1  gate932(.a(G1129), .O(gate482inter7));
  inv1  gate933(.a(G1225), .O(gate482inter8));
  nand2 gate934(.a(gate482inter8), .b(gate482inter7), .O(gate482inter9));
  nand2 gate935(.a(s_55), .b(gate482inter3), .O(gate482inter10));
  nor2  gate936(.a(gate482inter10), .b(gate482inter9), .O(gate482inter11));
  nor2  gate937(.a(gate482inter11), .b(gate482inter6), .O(gate482inter12));
  nand2 gate938(.a(gate482inter12), .b(gate482inter1), .O(G1291));
nand2 gate483( .a(G1228), .b(G1229), .O(G1292) );
nand2 gate484( .a(G1230), .b(G1231), .O(G1293) );

  xor2  gate1079(.a(G1233), .b(G1232), .O(gate485inter0));
  nand2 gate1080(.a(gate485inter0), .b(s_76), .O(gate485inter1));
  and2  gate1081(.a(G1233), .b(G1232), .O(gate485inter2));
  inv1  gate1082(.a(s_76), .O(gate485inter3));
  inv1  gate1083(.a(s_77), .O(gate485inter4));
  nand2 gate1084(.a(gate485inter4), .b(gate485inter3), .O(gate485inter5));
  nor2  gate1085(.a(gate485inter5), .b(gate485inter2), .O(gate485inter6));
  inv1  gate1086(.a(G1232), .O(gate485inter7));
  inv1  gate1087(.a(G1233), .O(gate485inter8));
  nand2 gate1088(.a(gate485inter8), .b(gate485inter7), .O(gate485inter9));
  nand2 gate1089(.a(s_77), .b(gate485inter3), .O(gate485inter10));
  nor2  gate1090(.a(gate485inter10), .b(gate485inter9), .O(gate485inter11));
  nor2  gate1091(.a(gate485inter11), .b(gate485inter6), .O(gate485inter12));
  nand2 gate1092(.a(gate485inter12), .b(gate485inter1), .O(G1294));
nand2 gate486( .a(G1234), .b(G1235), .O(G1295) );
nand2 gate487( .a(G1236), .b(G1237), .O(G1296) );
nand2 gate488( .a(G1238), .b(G1239), .O(G1297) );

  xor2  gate911(.a(G1241), .b(G1240), .O(gate489inter0));
  nand2 gate912(.a(gate489inter0), .b(s_52), .O(gate489inter1));
  and2  gate913(.a(G1241), .b(G1240), .O(gate489inter2));
  inv1  gate914(.a(s_52), .O(gate489inter3));
  inv1  gate915(.a(s_53), .O(gate489inter4));
  nand2 gate916(.a(gate489inter4), .b(gate489inter3), .O(gate489inter5));
  nor2  gate917(.a(gate489inter5), .b(gate489inter2), .O(gate489inter6));
  inv1  gate918(.a(G1240), .O(gate489inter7));
  inv1  gate919(.a(G1241), .O(gate489inter8));
  nand2 gate920(.a(gate489inter8), .b(gate489inter7), .O(gate489inter9));
  nand2 gate921(.a(s_53), .b(gate489inter3), .O(gate489inter10));
  nor2  gate922(.a(gate489inter10), .b(gate489inter9), .O(gate489inter11));
  nor2  gate923(.a(gate489inter11), .b(gate489inter6), .O(gate489inter12));
  nand2 gate924(.a(gate489inter12), .b(gate489inter1), .O(G1298));
nand2 gate490( .a(G1242), .b(G1243), .O(G1299) );
nand2 gate491( .a(G1244), .b(G1245), .O(G1300) );
nand2 gate492( .a(G1246), .b(G1247), .O(G1301) );
nand2 gate493( .a(G1248), .b(G1249), .O(G1302) );
nand2 gate494( .a(G1250), .b(G1251), .O(G1303) );
nand2 gate495( .a(G1252), .b(G1253), .O(G1304) );
nand2 gate496( .a(G1254), .b(G1255), .O(G1305) );

  xor2  gate1317(.a(G1257), .b(G1256), .O(gate497inter0));
  nand2 gate1318(.a(gate497inter0), .b(s_110), .O(gate497inter1));
  and2  gate1319(.a(G1257), .b(G1256), .O(gate497inter2));
  inv1  gate1320(.a(s_110), .O(gate497inter3));
  inv1  gate1321(.a(s_111), .O(gate497inter4));
  nand2 gate1322(.a(gate497inter4), .b(gate497inter3), .O(gate497inter5));
  nor2  gate1323(.a(gate497inter5), .b(gate497inter2), .O(gate497inter6));
  inv1  gate1324(.a(G1256), .O(gate497inter7));
  inv1  gate1325(.a(G1257), .O(gate497inter8));
  nand2 gate1326(.a(gate497inter8), .b(gate497inter7), .O(gate497inter9));
  nand2 gate1327(.a(s_111), .b(gate497inter3), .O(gate497inter10));
  nor2  gate1328(.a(gate497inter10), .b(gate497inter9), .O(gate497inter11));
  nor2  gate1329(.a(gate497inter11), .b(gate497inter6), .O(gate497inter12));
  nand2 gate1330(.a(gate497inter12), .b(gate497inter1), .O(G1306));
nand2 gate498( .a(G1258), .b(G1259), .O(G1307) );
nand2 gate499( .a(G1260), .b(G1261), .O(G1308) );
nand2 gate500( .a(G1262), .b(G1263), .O(G1309) );
nand2 gate501( .a(G1264), .b(G1265), .O(G1310) );
nand2 gate502( .a(G1266), .b(G1267), .O(G1311) );
nand2 gate503( .a(G1268), .b(G1269), .O(G1312) );

  xor2  gate813(.a(G1271), .b(G1270), .O(gate504inter0));
  nand2 gate814(.a(gate504inter0), .b(s_38), .O(gate504inter1));
  and2  gate815(.a(G1271), .b(G1270), .O(gate504inter2));
  inv1  gate816(.a(s_38), .O(gate504inter3));
  inv1  gate817(.a(s_39), .O(gate504inter4));
  nand2 gate818(.a(gate504inter4), .b(gate504inter3), .O(gate504inter5));
  nor2  gate819(.a(gate504inter5), .b(gate504inter2), .O(gate504inter6));
  inv1  gate820(.a(G1270), .O(gate504inter7));
  inv1  gate821(.a(G1271), .O(gate504inter8));
  nand2 gate822(.a(gate504inter8), .b(gate504inter7), .O(gate504inter9));
  nand2 gate823(.a(s_39), .b(gate504inter3), .O(gate504inter10));
  nor2  gate824(.a(gate504inter10), .b(gate504inter9), .O(gate504inter11));
  nor2  gate825(.a(gate504inter11), .b(gate504inter6), .O(gate504inter12));
  nand2 gate826(.a(gate504inter12), .b(gate504inter1), .O(G1313));
nand2 gate505( .a(G1272), .b(G1273), .O(G1314) );
nand2 gate506( .a(G1274), .b(G1275), .O(G1315) );
nand2 gate507( .a(G1276), .b(G1277), .O(G1316) );
nand2 gate508( .a(G1278), .b(G1279), .O(G1317) );
nand2 gate509( .a(G1280), .b(G1281), .O(G1318) );
nand2 gate510( .a(G1282), .b(G1283), .O(G1319) );

  xor2  gate1177(.a(G1285), .b(G1284), .O(gate511inter0));
  nand2 gate1178(.a(gate511inter0), .b(s_90), .O(gate511inter1));
  and2  gate1179(.a(G1285), .b(G1284), .O(gate511inter2));
  inv1  gate1180(.a(s_90), .O(gate511inter3));
  inv1  gate1181(.a(s_91), .O(gate511inter4));
  nand2 gate1182(.a(gate511inter4), .b(gate511inter3), .O(gate511inter5));
  nor2  gate1183(.a(gate511inter5), .b(gate511inter2), .O(gate511inter6));
  inv1  gate1184(.a(G1284), .O(gate511inter7));
  inv1  gate1185(.a(G1285), .O(gate511inter8));
  nand2 gate1186(.a(gate511inter8), .b(gate511inter7), .O(gate511inter9));
  nand2 gate1187(.a(s_91), .b(gate511inter3), .O(gate511inter10));
  nor2  gate1188(.a(gate511inter10), .b(gate511inter9), .O(gate511inter11));
  nor2  gate1189(.a(gate511inter11), .b(gate511inter6), .O(gate511inter12));
  nand2 gate1190(.a(gate511inter12), .b(gate511inter1), .O(G1320));
nand2 gate512( .a(G1286), .b(G1287), .O(G1321) );
nand2 gate513( .a(G1288), .b(G1289), .O(G1322) );
nand2 gate514( .a(G1290), .b(G1291), .O(G1323) );
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule