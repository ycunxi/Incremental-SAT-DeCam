module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);

input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;//RE__PI;

input s_0,s_1;//RE__ALLOW(00,01,10,11);
input s_2,s_3;//RE__ALLOW(00,01,10,11);
input s_4,s_5;//RE__ALLOW(00,01,10,11);
input s_6,s_7;//RE__ALLOW(00,01,10,11);
input s_8,s_9;//RE__ALLOW(00,01,10,11);
input s_10,s_11;//RE__ALLOW(00,01,10,11);
input s_12,s_13;//RE__ALLOW(00,01,10,11);
input s_14,s_15;//RE__ALLOW(00,01,10,11);
input s_16,s_17;//RE__ALLOW(00,01,10,11);
input s_18,s_19;//RE__ALLOW(00,01,10,11);
input s_20,s_21;//RE__ALLOW(00,01,10,11);
input s_22,s_23;//RE__ALLOW(00,01,10,11);
input s_24,s_25;//RE__ALLOW(00,01,10,11);
input s_26,s_27;//RE__ALLOW(00,01,10,11);
input s_28,s_29;//RE__ALLOW(00,01,10,11);
input s_30,s_31;//RE__ALLOW(00,01,10,11);
input s_32,s_33;//RE__ALLOW(00,01,10,11);
input s_34,s_35;//RE__ALLOW(00,01,10,11);
input s_36,s_37;//RE__ALLOW(00,01,10,11);
input s_38,s_39;//RE__ALLOW(00,01,10,11);
input s_40,s_41;//RE__ALLOW(00,01,10,11);
input s_42,s_43;//RE__ALLOW(00,01,10,11);
input s_44,s_45;//RE__ALLOW(00,01,10,11);
input s_46,s_47;//RE__ALLOW(00,01,10,11);
input s_48,s_49;//RE__ALLOW(00,01,10,11);
input s_50,s_51;//RE__ALLOW(00,01,10,11);
input s_52,s_53;//RE__ALLOW(00,01,10,11);
input s_54,s_55;//RE__ALLOW(00,01,10,11);
input s_56,s_57;//RE__ALLOW(00,01,10,11);
input s_58,s_59;//RE__ALLOW(00,01,10,11);
input s_60,s_61;//RE__ALLOW(00,01,10,11);
input s_62,s_63;//RE__ALLOW(00,01,10,11);
input s_64,s_65;//RE__ALLOW(00,01,10,11);
input s_66,s_67;//RE__ALLOW(00,01,10,11);
input s_68,s_69;//RE__ALLOW(00,01,10,11);
input s_70,s_71;//RE__ALLOW(00,01,10,11);
input s_72,s_73;//RE__ALLOW(00,01,10,11);
input s_74,s_75;//RE__ALLOW(00,01,10,11);
input s_76,s_77;//RE__ALLOW(00,01,10,11);
input s_78,s_79;//RE__ALLOW(00,01,10,11);
input s_80,s_81;//RE__ALLOW(00,01,10,11);
input s_82,s_83;//RE__ALLOW(00,01,10,11);
input s_84,s_85;//RE__ALLOW(00,01,10,11);
input s_86,s_87;//RE__ALLOW(00,01,10,11);
input s_88,s_89;//RE__ALLOW(00,01,10,11);
input s_90,s_91;//RE__ALLOW(00,01,10,11);
input s_92,s_93;//RE__ALLOW(00,01,10,11);
input s_94,s_95;//RE__ALLOW(00,01,10,11);
input s_96,s_97;//RE__ALLOW(00,01,10,11);
input s_98,s_99;//RE__ALLOW(00,01,10,11);
input s_100,s_101;//RE__ALLOW(00,01,10,11);
input s_102,s_103;//RE__ALLOW(00,01,10,11);
input s_104,s_105;//RE__ALLOW(00,01,10,11);
input s_106,s_107;//RE__ALLOW(00,01,10,11);
input s_108,s_109;//RE__ALLOW(00,01,10,11);
input s_110,s_111;//RE__ALLOW(00,01,10,11);
input s_112,s_113;//RE__ALLOW(00,01,10,11);
input s_114,s_115;//RE__ALLOW(00,01,10,11);
input s_116,s_117;//RE__ALLOW(00,01,10,11);
input s_118,s_119;//RE__ALLOW(00,01,10,11);
input s_120,s_121;//RE__ALLOW(00,01,10,11);
input s_122,s_123;//RE__ALLOW(00,01,10,11);
input s_124,s_125;//RE__ALLOW(00,01,10,11);
input s_126,s_127;//RE__ALLOW(00,01,10,11);
input s_128,s_129;//RE__ALLOW(00,01,10,11);
input s_130,s_131;//RE__ALLOW(00,01,10,11);
input s_132,s_133;//RE__ALLOW(00,01,10,11);
input s_134,s_135;//RE__ALLOW(00,01,10,11);
input s_136,s_137;//RE__ALLOW(00,01,10,11);
input s_138,s_139;//RE__ALLOW(00,01,10,11);
input s_140,s_141;//RE__ALLOW(00,01,10,11);
input s_142,s_143;//RE__ALLOW(00,01,10,11);
input s_144,s_145;//RE__ALLOW(00,01,10,11);
input s_146,s_147;//RE__ALLOW(00,01,10,11);
input s_148,s_149;//RE__ALLOW(00,01,10,11);
input s_150,s_151;//RE__ALLOW(00,01,10,11);
input s_152,s_153;//RE__ALLOW(00,01,10,11);
input s_154,s_155;//RE__ALLOW(00,01,10,11);
input s_156,s_157;//RE__ALLOW(00,01,10,11);
input s_158,s_159;//RE__ALLOW(00,01,10,11);
input s_160,s_161;//RE__ALLOW(00,01,10,11);
input s_162,s_163;//RE__ALLOW(00,01,10,11);
input s_164,s_165;//RE__ALLOW(00,01,10,11);
input s_166,s_167;//RE__ALLOW(00,01,10,11);
input s_168,s_169;//RE__ALLOW(00,01,10,11);
input s_170,s_171;//RE__ALLOW(00,01,10,11);
input s_172,s_173;//RE__ALLOW(00,01,10,11);
input s_174,s_175;//RE__ALLOW(00,01,10,11);
input s_176,s_177;//RE__ALLOW(00,01,10,11);
input s_178,s_179;//RE__ALLOW(00,01,10,11);
input s_180,s_181;//RE__ALLOW(00,01,10,11);
input s_182,s_183;//RE__ALLOW(00,01,10,11);
input s_184,s_185;//RE__ALLOW(00,01,10,11);
input s_186,s_187;//RE__ALLOW(00,01,10,11);
input s_188,s_189;//RE__ALLOW(00,01,10,11);
input s_190,s_191;//RE__ALLOW(00,01,10,11);
input s_192,s_193;//RE__ALLOW(00,01,10,11);
input s_194,s_195;//RE__ALLOW(00,01,10,11);
input s_196,s_197;//RE__ALLOW(00,01,10,11);
input s_198,s_199;//RE__ALLOW(00,01,10,11);
input s_200,s_201;//RE__ALLOW(00,01,10,11);
input s_202,s_203;//RE__ALLOW(00,01,10,11);
input s_204,s_205;//RE__ALLOW(00,01,10,11);
input s_206,s_207;//RE__ALLOW(00,01,10,11);
input s_208,s_209;//RE__ALLOW(00,01,10,11);
input s_210,s_211;//RE__ALLOW(00,01,10,11);
input s_212,s_213;//RE__ALLOW(00,01,10,11);
input s_214,s_215;//RE__ALLOW(00,01,10,11);
input s_216,s_217;//RE__ALLOW(00,01,10,11);
input s_218,s_219;//RE__ALLOW(00,01,10,11);
input s_220,s_221;//RE__ALLOW(00,01,10,11);
input s_222,s_223;//RE__ALLOW(00,01,10,11);
input s_224,s_225;//RE__ALLOW(00,01,10,11);
input s_226,s_227;//RE__ALLOW(00,01,10,11);
input s_228,s_229;//RE__ALLOW(00,01,10,11);
input s_230,s_231;//RE__ALLOW(00,01,10,11);
input s_232,s_233;//RE__ALLOW(00,01,10,11);
input s_234,s_235;//RE__ALLOW(00,01,10,11);
input s_236,s_237;//RE__ALLOW(00,01,10,11);
input s_238,s_239;//RE__ALLOW(00,01,10,11);
input s_240,s_241;//RE__ALLOW(00,01,10,11);
input s_242,s_243;//RE__ALLOW(00,01,10,11);
input s_244,s_245;//RE__ALLOW(00,01,10,11);
input s_246,s_247;//RE__ALLOW(00,01,10,11);
input s_248,s_249;//RE__ALLOW(00,01,10,11);
input s_250,s_251;//RE__ALLOW(00,01,10,11);
input s_252,s_253;//RE__ALLOW(00,01,10,11);
input s_254,s_255;//RE__ALLOW(00,01,10,11);
input s_256,s_257;//RE__ALLOW(00,01,10,11);
input s_258,s_259;//RE__ALLOW(00,01,10,11);
input s_260,s_261;//RE__ALLOW(00,01,10,11);
input s_262,s_263;//RE__ALLOW(00,01,10,11);
input s_264,s_265;//RE__ALLOW(00,01,10,11);
input s_266,s_267;//RE__ALLOW(00,01,10,11);
input s_268,s_269;//RE__ALLOW(00,01,10,11);
input s_270,s_271;//RE__ALLOW(00,01,10,11);
input s_272,s_273;//RE__ALLOW(00,01,10,11);
input s_274,s_275;//RE__ALLOW(00,01,10,11);
input s_276,s_277;//RE__ALLOW(00,01,10,11);
input s_278,s_279;//RE__ALLOW(00,01,10,11);
input s_280,s_281;//RE__ALLOW(00,01,10,11);
input s_282,s_283;//RE__ALLOW(00,01,10,11);
input s_284,s_285;//RE__ALLOW(00,01,10,11);
input s_286,s_287;//RE__ALLOW(00,01,10,11);
input s_288,s_289;//RE__ALLOW(00,01,10,11);
input s_290,s_291;//RE__ALLOW(00,01,10,11);
input s_292,s_293;//RE__ALLOW(00,01,10,11);
input s_294,s_295;//RE__ALLOW(00,01,10,11);
input s_296,s_297;//RE__ALLOW(00,01,10,11);
input s_298,s_299;//RE__ALLOW(00,01,10,11);
input s_300,s_301;//RE__ALLOW(00,01,10,11);
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;

  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate100inter0, gate100inter1, gate100inter2, gate100inter3, gate100inter4, gate100inter5, gate100inter6, gate100inter7, gate100inter8, gate100inter9, gate100inter10, gate100inter11, gate100inter12, gate177inter0, gate177inter1, gate177inter2, gate177inter3, gate177inter4, gate177inter5, gate177inter6, gate177inter7, gate177inter8, gate177inter9, gate177inter10, gate177inter11, gate177inter12, gate254inter0, gate254inter1, gate254inter2, gate254inter3, gate254inter4, gate254inter5, gate254inter6, gate254inter7, gate254inter8, gate254inter9, gate254inter10, gate254inter11, gate254inter12, gate101inter0, gate101inter1, gate101inter2, gate101inter3, gate101inter4, gate101inter5, gate101inter6, gate101inter7, gate101inter8, gate101inter9, gate101inter10, gate101inter11, gate101inter12, gate199inter0, gate199inter1, gate199inter2, gate199inter3, gate199inter4, gate199inter5, gate199inter6, gate199inter7, gate199inter8, gate199inter9, gate199inter10, gate199inter11, gate199inter12, gate17inter0, gate17inter1, gate17inter2, gate17inter3, gate17inter4, gate17inter5, gate17inter6, gate17inter7, gate17inter8, gate17inter9, gate17inter10, gate17inter11, gate17inter12, gate85inter0, gate85inter1, gate85inter2, gate85inter3, gate85inter4, gate85inter5, gate85inter6, gate85inter7, gate85inter8, gate85inter9, gate85inter10, gate85inter11, gate85inter12, gate489inter0, gate489inter1, gate489inter2, gate489inter3, gate489inter4, gate489inter5, gate489inter6, gate489inter7, gate489inter8, gate489inter9, gate489inter10, gate489inter11, gate489inter12, gate13inter0, gate13inter1, gate13inter2, gate13inter3, gate13inter4, gate13inter5, gate13inter6, gate13inter7, gate13inter8, gate13inter9, gate13inter10, gate13inter11, gate13inter12, gate408inter0, gate408inter1, gate408inter2, gate408inter3, gate408inter4, gate408inter5, gate408inter6, gate408inter7, gate408inter8, gate408inter9, gate408inter10, gate408inter11, gate408inter12, gate273inter0, gate273inter1, gate273inter2, gate273inter3, gate273inter4, gate273inter5, gate273inter6, gate273inter7, gate273inter8, gate273inter9, gate273inter10, gate273inter11, gate273inter12, gate75inter0, gate75inter1, gate75inter2, gate75inter3, gate75inter4, gate75inter5, gate75inter6, gate75inter7, gate75inter8, gate75inter9, gate75inter10, gate75inter11, gate75inter12, gate65inter0, gate65inter1, gate65inter2, gate65inter3, gate65inter4, gate65inter5, gate65inter6, gate65inter7, gate65inter8, gate65inter9, gate65inter10, gate65inter11, gate65inter12, gate154inter0, gate154inter1, gate154inter2, gate154inter3, gate154inter4, gate154inter5, gate154inter6, gate154inter7, gate154inter8, gate154inter9, gate154inter10, gate154inter11, gate154inter12, gate153inter0, gate153inter1, gate153inter2, gate153inter3, gate153inter4, gate153inter5, gate153inter6, gate153inter7, gate153inter8, gate153inter9, gate153inter10, gate153inter11, gate153inter12, gate132inter0, gate132inter1, gate132inter2, gate132inter3, gate132inter4, gate132inter5, gate132inter6, gate132inter7, gate132inter8, gate132inter9, gate132inter10, gate132inter11, gate132inter12, gate197inter0, gate197inter1, gate197inter2, gate197inter3, gate197inter4, gate197inter5, gate197inter6, gate197inter7, gate197inter8, gate197inter9, gate197inter10, gate197inter11, gate197inter12, gate282inter0, gate282inter1, gate282inter2, gate282inter3, gate282inter4, gate282inter5, gate282inter6, gate282inter7, gate282inter8, gate282inter9, gate282inter10, gate282inter11, gate282inter12, gate391inter0, gate391inter1, gate391inter2, gate391inter3, gate391inter4, gate391inter5, gate391inter6, gate391inter7, gate391inter8, gate391inter9, gate391inter10, gate391inter11, gate391inter12, gate247inter0, gate247inter1, gate247inter2, gate247inter3, gate247inter4, gate247inter5, gate247inter6, gate247inter7, gate247inter8, gate247inter9, gate247inter10, gate247inter11, gate247inter12, gate62inter0, gate62inter1, gate62inter2, gate62inter3, gate62inter4, gate62inter5, gate62inter6, gate62inter7, gate62inter8, gate62inter9, gate62inter10, gate62inter11, gate62inter12, gate22inter0, gate22inter1, gate22inter2, gate22inter3, gate22inter4, gate22inter5, gate22inter6, gate22inter7, gate22inter8, gate22inter9, gate22inter10, gate22inter11, gate22inter12, gate84inter0, gate84inter1, gate84inter2, gate84inter3, gate84inter4, gate84inter5, gate84inter6, gate84inter7, gate84inter8, gate84inter9, gate84inter10, gate84inter11, gate84inter12, gate130inter0, gate130inter1, gate130inter2, gate130inter3, gate130inter4, gate130inter5, gate130inter6, gate130inter7, gate130inter8, gate130inter9, gate130inter10, gate130inter11, gate130inter12, gate92inter0, gate92inter1, gate92inter2, gate92inter3, gate92inter4, gate92inter5, gate92inter6, gate92inter7, gate92inter8, gate92inter9, gate92inter10, gate92inter11, gate92inter12, gate426inter0, gate426inter1, gate426inter2, gate426inter3, gate426inter4, gate426inter5, gate426inter6, gate426inter7, gate426inter8, gate426inter9, gate426inter10, gate426inter11, gate426inter12, gate478inter0, gate478inter1, gate478inter2, gate478inter3, gate478inter4, gate478inter5, gate478inter6, gate478inter7, gate478inter8, gate478inter9, gate478inter10, gate478inter11, gate478inter12, gate461inter0, gate461inter1, gate461inter2, gate461inter3, gate461inter4, gate461inter5, gate461inter6, gate461inter7, gate461inter8, gate461inter9, gate461inter10, gate461inter11, gate461inter12, gate32inter0, gate32inter1, gate32inter2, gate32inter3, gate32inter4, gate32inter5, gate32inter6, gate32inter7, gate32inter8, gate32inter9, gate32inter10, gate32inter11, gate32inter12, gate430inter0, gate430inter1, gate430inter2, gate430inter3, gate430inter4, gate430inter5, gate430inter6, gate430inter7, gate430inter8, gate430inter9, gate430inter10, gate430inter11, gate430inter12, gate509inter0, gate509inter1, gate509inter2, gate509inter3, gate509inter4, gate509inter5, gate509inter6, gate509inter7, gate509inter8, gate509inter9, gate509inter10, gate509inter11, gate509inter12, gate117inter0, gate117inter1, gate117inter2, gate117inter3, gate117inter4, gate117inter5, gate117inter6, gate117inter7, gate117inter8, gate117inter9, gate117inter10, gate117inter11, gate117inter12, gate107inter0, gate107inter1, gate107inter2, gate107inter3, gate107inter4, gate107inter5, gate107inter6, gate107inter7, gate107inter8, gate107inter9, gate107inter10, gate107inter11, gate107inter12, gate163inter0, gate163inter1, gate163inter2, gate163inter3, gate163inter4, gate163inter5, gate163inter6, gate163inter7, gate163inter8, gate163inter9, gate163inter10, gate163inter11, gate163inter12, gate186inter0, gate186inter1, gate186inter2, gate186inter3, gate186inter4, gate186inter5, gate186inter6, gate186inter7, gate186inter8, gate186inter9, gate186inter10, gate186inter11, gate186inter12, gate114inter0, gate114inter1, gate114inter2, gate114inter3, gate114inter4, gate114inter5, gate114inter6, gate114inter7, gate114inter8, gate114inter9, gate114inter10, gate114inter11, gate114inter12, gate233inter0, gate233inter1, gate233inter2, gate233inter3, gate233inter4, gate233inter5, gate233inter6, gate233inter7, gate233inter8, gate233inter9, gate233inter10, gate233inter11, gate233inter12, gate160inter0, gate160inter1, gate160inter2, gate160inter3, gate160inter4, gate160inter5, gate160inter6, gate160inter7, gate160inter8, gate160inter9, gate160inter10, gate160inter11, gate160inter12, gate48inter0, gate48inter1, gate48inter2, gate48inter3, gate48inter4, gate48inter5, gate48inter6, gate48inter7, gate48inter8, gate48inter9, gate48inter10, gate48inter11, gate48inter12, gate494inter0, gate494inter1, gate494inter2, gate494inter3, gate494inter4, gate494inter5, gate494inter6, gate494inter7, gate494inter8, gate494inter9, gate494inter10, gate494inter11, gate494inter12, gate234inter0, gate234inter1, gate234inter2, gate234inter3, gate234inter4, gate234inter5, gate234inter6, gate234inter7, gate234inter8, gate234inter9, gate234inter10, gate234inter11, gate234inter12, gate162inter0, gate162inter1, gate162inter2, gate162inter3, gate162inter4, gate162inter5, gate162inter6, gate162inter7, gate162inter8, gate162inter9, gate162inter10, gate162inter11, gate162inter12, gate460inter0, gate460inter1, gate460inter2, gate460inter3, gate460inter4, gate460inter5, gate460inter6, gate460inter7, gate460inter8, gate460inter9, gate460inter10, gate460inter11, gate460inter12, gate176inter0, gate176inter1, gate176inter2, gate176inter3, gate176inter4, gate176inter5, gate176inter6, gate176inter7, gate176inter8, gate176inter9, gate176inter10, gate176inter11, gate176inter12, gate243inter0, gate243inter1, gate243inter2, gate243inter3, gate243inter4, gate243inter5, gate243inter6, gate243inter7, gate243inter8, gate243inter9, gate243inter10, gate243inter11, gate243inter12, gate501inter0, gate501inter1, gate501inter2, gate501inter3, gate501inter4, gate501inter5, gate501inter6, gate501inter7, gate501inter8, gate501inter9, gate501inter10, gate501inter11, gate501inter12, gate201inter0, gate201inter1, gate201inter2, gate201inter3, gate201inter4, gate201inter5, gate201inter6, gate201inter7, gate201inter8, gate201inter9, gate201inter10, gate201inter11, gate201inter12, gate498inter0, gate498inter1, gate498inter2, gate498inter3, gate498inter4, gate498inter5, gate498inter6, gate498inter7, gate498inter8, gate498inter9, gate498inter10, gate498inter11, gate498inter12, gate152inter0, gate152inter1, gate152inter2, gate152inter3, gate152inter4, gate152inter5, gate152inter6, gate152inter7, gate152inter8, gate152inter9, gate152inter10, gate152inter11, gate152inter12, gate394inter0, gate394inter1, gate394inter2, gate394inter3, gate394inter4, gate394inter5, gate394inter6, gate394inter7, gate394inter8, gate394inter9, gate394inter10, gate394inter11, gate394inter12, gate166inter0, gate166inter1, gate166inter2, gate166inter3, gate166inter4, gate166inter5, gate166inter6, gate166inter7, gate166inter8, gate166inter9, gate166inter10, gate166inter11, gate166inter12, gate35inter0, gate35inter1, gate35inter2, gate35inter3, gate35inter4, gate35inter5, gate35inter6, gate35inter7, gate35inter8, gate35inter9, gate35inter10, gate35inter11, gate35inter12, gate448inter0, gate448inter1, gate448inter2, gate448inter3, gate448inter4, gate448inter5, gate448inter6, gate448inter7, gate448inter8, gate448inter9, gate448inter10, gate448inter11, gate448inter12, gate263inter0, gate263inter1, gate263inter2, gate263inter3, gate263inter4, gate263inter5, gate263inter6, gate263inter7, gate263inter8, gate263inter9, gate263inter10, gate263inter11, gate263inter12, gate60inter0, gate60inter1, gate60inter2, gate60inter3, gate60inter4, gate60inter5, gate60inter6, gate60inter7, gate60inter8, gate60inter9, gate60inter10, gate60inter11, gate60inter12, gate449inter0, gate449inter1, gate449inter2, gate449inter3, gate449inter4, gate449inter5, gate449inter6, gate449inter7, gate449inter8, gate449inter9, gate449inter10, gate449inter11, gate449inter12, gate499inter0, gate499inter1, gate499inter2, gate499inter3, gate499inter4, gate499inter5, gate499inter6, gate499inter7, gate499inter8, gate499inter9, gate499inter10, gate499inter11, gate499inter12, gate95inter0, gate95inter1, gate95inter2, gate95inter3, gate95inter4, gate95inter5, gate95inter6, gate95inter7, gate95inter8, gate95inter9, gate95inter10, gate95inter11, gate95inter12, gate451inter0, gate451inter1, gate451inter2, gate451inter3, gate451inter4, gate451inter5, gate451inter6, gate451inter7, gate451inter8, gate451inter9, gate451inter10, gate451inter11, gate451inter12, gate102inter0, gate102inter1, gate102inter2, gate102inter3, gate102inter4, gate102inter5, gate102inter6, gate102inter7, gate102inter8, gate102inter9, gate102inter10, gate102inter11, gate102inter12, gate278inter0, gate278inter1, gate278inter2, gate278inter3, gate278inter4, gate278inter5, gate278inter6, gate278inter7, gate278inter8, gate278inter9, gate278inter10, gate278inter11, gate278inter12, gate15inter0, gate15inter1, gate15inter2, gate15inter3, gate15inter4, gate15inter5, gate15inter6, gate15inter7, gate15inter8, gate15inter9, gate15inter10, gate15inter11, gate15inter12, gate165inter0, gate165inter1, gate165inter2, gate165inter3, gate165inter4, gate165inter5, gate165inter6, gate165inter7, gate165inter8, gate165inter9, gate165inter10, gate165inter11, gate165inter12, gate445inter0, gate445inter1, gate445inter2, gate445inter3, gate445inter4, gate445inter5, gate445inter6, gate445inter7, gate445inter8, gate445inter9, gate445inter10, gate445inter11, gate445inter12, gate68inter0, gate68inter1, gate68inter2, gate68inter3, gate68inter4, gate68inter5, gate68inter6, gate68inter7, gate68inter8, gate68inter9, gate68inter10, gate68inter11, gate68inter12, gate147inter0, gate147inter1, gate147inter2, gate147inter3, gate147inter4, gate147inter5, gate147inter6, gate147inter7, gate147inter8, gate147inter9, gate147inter10, gate147inter11, gate147inter12, gate137inter0, gate137inter1, gate137inter2, gate137inter3, gate137inter4, gate137inter5, gate137inter6, gate137inter7, gate137inter8, gate137inter9, gate137inter10, gate137inter11, gate137inter12, gate183inter0, gate183inter1, gate183inter2, gate183inter3, gate183inter4, gate183inter5, gate183inter6, gate183inter7, gate183inter8, gate183inter9, gate183inter10, gate183inter11, gate183inter12, gate511inter0, gate511inter1, gate511inter2, gate511inter3, gate511inter4, gate511inter5, gate511inter6, gate511inter7, gate511inter8, gate511inter9, gate511inter10, gate511inter11, gate511inter12, gate239inter0, gate239inter1, gate239inter2, gate239inter3, gate239inter4, gate239inter5, gate239inter6, gate239inter7, gate239inter8, gate239inter9, gate239inter10, gate239inter11, gate239inter12, gate457inter0, gate457inter1, gate457inter2, gate457inter3, gate457inter4, gate457inter5, gate457inter6, gate457inter7, gate457inter8, gate457inter9, gate457inter10, gate457inter11, gate457inter12, gate441inter0, gate441inter1, gate441inter2, gate441inter3, gate441inter4, gate441inter5, gate441inter6, gate441inter7, gate441inter8, gate441inter9, gate441inter10, gate441inter11, gate441inter12, gate476inter0, gate476inter1, gate476inter2, gate476inter3, gate476inter4, gate476inter5, gate476inter6, gate476inter7, gate476inter8, gate476inter9, gate476inter10, gate476inter11, gate476inter12, gate76inter0, gate76inter1, gate76inter2, gate76inter3, gate76inter4, gate76inter5, gate76inter6, gate76inter7, gate76inter8, gate76inter9, gate76inter10, gate76inter11, gate76inter12, gate285inter0, gate285inter1, gate285inter2, gate285inter3, gate285inter4, gate285inter5, gate285inter6, gate285inter7, gate285inter8, gate285inter9, gate285inter10, gate285inter11, gate285inter12, gate482inter0, gate482inter1, gate482inter2, gate482inter3, gate482inter4, gate482inter5, gate482inter6, gate482inter7, gate482inter8, gate482inter9, gate482inter10, gate482inter11, gate482inter12, gate477inter0, gate477inter1, gate477inter2, gate477inter3, gate477inter4, gate477inter5, gate477inter6, gate477inter7, gate477inter8, gate477inter9, gate477inter10, gate477inter11, gate477inter12, gate175inter0, gate175inter1, gate175inter2, gate175inter3, gate175inter4, gate175inter5, gate175inter6, gate175inter7, gate175inter8, gate175inter9, gate175inter10, gate175inter11, gate175inter12, gate463inter0, gate463inter1, gate463inter2, gate463inter3, gate463inter4, gate463inter5, gate463inter6, gate463inter7, gate463inter8, gate463inter9, gate463inter10, gate463inter11, gate463inter12, gate484inter0, gate484inter1, gate484inter2, gate484inter3, gate484inter4, gate484inter5, gate484inter6, gate484inter7, gate484inter8, gate484inter9, gate484inter10, gate484inter11, gate484inter12, gate474inter0, gate474inter1, gate474inter2, gate474inter3, gate474inter4, gate474inter5, gate474inter6, gate474inter7, gate474inter8, gate474inter9, gate474inter10, gate474inter11, gate474inter12, gate294inter0, gate294inter1, gate294inter2, gate294inter3, gate294inter4, gate294inter5, gate294inter6, gate294inter7, gate294inter8, gate294inter9, gate294inter10, gate294inter11, gate294inter12, gate480inter0, gate480inter1, gate480inter2, gate480inter3, gate480inter4, gate480inter5, gate480inter6, gate480inter7, gate480inter8, gate480inter9, gate480inter10, gate480inter11, gate480inter12, gate503inter0, gate503inter1, gate503inter2, gate503inter3, gate503inter4, gate503inter5, gate503inter6, gate503inter7, gate503inter8, gate503inter9, gate503inter10, gate503inter11, gate503inter12, gate245inter0, gate245inter1, gate245inter2, gate245inter3, gate245inter4, gate245inter5, gate245inter6, gate245inter7, gate245inter8, gate245inter9, gate245inter10, gate245inter11, gate245inter12, gate24inter0, gate24inter1, gate24inter2, gate24inter3, gate24inter4, gate24inter5, gate24inter6, gate24inter7, gate24inter8, gate24inter9, gate24inter10, gate24inter11, gate24inter12, gate64inter0, gate64inter1, gate64inter2, gate64inter3, gate64inter4, gate64inter5, gate64inter6, gate64inter7, gate64inter8, gate64inter9, gate64inter10, gate64inter11, gate64inter12, gate82inter0, gate82inter1, gate82inter2, gate82inter3, gate82inter4, gate82inter5, gate82inter6, gate82inter7, gate82inter8, gate82inter9, gate82inter10, gate82inter11, gate82inter12, gate467inter0, gate467inter1, gate467inter2, gate467inter3, gate467inter4, gate467inter5, gate467inter6, gate467inter7, gate467inter8, gate467inter9, gate467inter10, gate467inter11, gate467inter12, gate133inter0, gate133inter1, gate133inter2, gate133inter3, gate133inter4, gate133inter5, gate133inter6, gate133inter7, gate133inter8, gate133inter9, gate133inter10, gate133inter11, gate133inter12, gate284inter0, gate284inter1, gate284inter2, gate284inter3, gate284inter4, gate284inter5, gate284inter6, gate284inter7, gate284inter8, gate284inter9, gate284inter10, gate284inter11, gate284inter12, gate388inter0, gate388inter1, gate388inter2, gate388inter3, gate388inter4, gate388inter5, gate388inter6, gate388inter7, gate388inter8, gate388inter9, gate388inter10, gate388inter11, gate388inter12, gate224inter0, gate224inter1, gate224inter2, gate224inter3, gate224inter4, gate224inter5, gate224inter6, gate224inter7, gate224inter8, gate224inter9, gate224inter10, gate224inter11, gate224inter12, gate401inter0, gate401inter1, gate401inter2, gate401inter3, gate401inter4, gate401inter5, gate401inter6, gate401inter7, gate401inter8, gate401inter9, gate401inter10, gate401inter11, gate401inter12, gate103inter0, gate103inter1, gate103inter2, gate103inter3, gate103inter4, gate103inter5, gate103inter6, gate103inter7, gate103inter8, gate103inter9, gate103inter10, gate103inter11, gate103inter12, gate174inter0, gate174inter1, gate174inter2, gate174inter3, gate174inter4, gate174inter5, gate174inter6, gate174inter7, gate174inter8, gate174inter9, gate174inter10, gate174inter11, gate174inter12, gate402inter0, gate402inter1, gate402inter2, gate402inter3, gate402inter4, gate402inter5, gate402inter6, gate402inter7, gate402inter8, gate402inter9, gate402inter10, gate402inter11, gate402inter12, gate44inter0, gate44inter1, gate44inter2, gate44inter3, gate44inter4, gate44inter5, gate44inter6, gate44inter7, gate44inter8, gate44inter9, gate44inter10, gate44inter11, gate44inter12, gate86inter0, gate86inter1, gate86inter2, gate86inter3, gate86inter4, gate86inter5, gate86inter6, gate86inter7, gate86inter8, gate86inter9, gate86inter10, gate86inter11, gate86inter12, gate410inter0, gate410inter1, gate410inter2, gate410inter3, gate410inter4, gate410inter5, gate410inter6, gate410inter7, gate410inter8, gate410inter9, gate410inter10, gate410inter11, gate410inter12, gate392inter0, gate392inter1, gate392inter2, gate392inter3, gate392inter4, gate392inter5, gate392inter6, gate392inter7, gate392inter8, gate392inter9, gate392inter10, gate392inter11, gate392inter12, gate112inter0, gate112inter1, gate112inter2, gate112inter3, gate112inter4, gate112inter5, gate112inter6, gate112inter7, gate112inter8, gate112inter9, gate112inter10, gate112inter11, gate112inter12, gate231inter0, gate231inter1, gate231inter2, gate231inter3, gate231inter4, gate231inter5, gate231inter6, gate231inter7, gate231inter8, gate231inter9, gate231inter10, gate231inter11, gate231inter12, gate456inter0, gate456inter1, gate456inter2, gate456inter3, gate456inter4, gate456inter5, gate456inter6, gate456inter7, gate456inter8, gate456inter9, gate456inter10, gate456inter11, gate456inter12, gate400inter0, gate400inter1, gate400inter2, gate400inter3, gate400inter4, gate400inter5, gate400inter6, gate400inter7, gate400inter8, gate400inter9, gate400inter10, gate400inter11, gate400inter12, gate397inter0, gate397inter1, gate397inter2, gate397inter3, gate397inter4, gate397inter5, gate397inter6, gate397inter7, gate397inter8, gate397inter9, gate397inter10, gate397inter11, gate397inter12, gate135inter0, gate135inter1, gate135inter2, gate135inter3, gate135inter4, gate135inter5, gate135inter6, gate135inter7, gate135inter8, gate135inter9, gate135inter10, gate135inter11, gate135inter12, gate38inter0, gate38inter1, gate38inter2, gate38inter3, gate38inter4, gate38inter5, gate38inter6, gate38inter7, gate38inter8, gate38inter9, gate38inter10, gate38inter11, gate38inter12, gate447inter0, gate447inter1, gate447inter2, gate447inter3, gate447inter4, gate447inter5, gate447inter6, gate447inter7, gate447inter8, gate447inter9, gate447inter10, gate447inter11, gate447inter12, gate472inter0, gate472inter1, gate472inter2, gate472inter3, gate472inter4, gate472inter5, gate472inter6, gate472inter7, gate472inter8, gate472inter9, gate472inter10, gate472inter11, gate472inter12, gate502inter0, gate502inter1, gate502inter2, gate502inter3, gate502inter4, gate502inter5, gate502inter6, gate502inter7, gate502inter8, gate502inter9, gate502inter10, gate502inter11, gate502inter12, gate161inter0, gate161inter1, gate161inter2, gate161inter3, gate161inter4, gate161inter5, gate161inter6, gate161inter7, gate161inter8, gate161inter9, gate161inter10, gate161inter11, gate161inter12, gate272inter0, gate272inter1, gate272inter2, gate272inter3, gate272inter4, gate272inter5, gate272inter6, gate272inter7, gate272inter8, gate272inter9, gate272inter10, gate272inter11, gate272inter12, gate43inter0, gate43inter1, gate43inter2, gate43inter3, gate43inter4, gate43inter5, gate43inter6, gate43inter7, gate43inter8, gate43inter9, gate43inter10, gate43inter11, gate43inter12, gate90inter0, gate90inter1, gate90inter2, gate90inter3, gate90inter4, gate90inter5, gate90inter6, gate90inter7, gate90inter8, gate90inter9, gate90inter10, gate90inter11, gate90inter12, gate486inter0, gate486inter1, gate486inter2, gate486inter3, gate486inter4, gate486inter5, gate486inter6, gate486inter7, gate486inter8, gate486inter9, gate486inter10, gate486inter11, gate486inter12, gate34inter0, gate34inter1, gate34inter2, gate34inter3, gate34inter4, gate34inter5, gate34inter6, gate34inter7, gate34inter8, gate34inter9, gate34inter10, gate34inter11, gate34inter12, gate264inter0, gate264inter1, gate264inter2, gate264inter3, gate264inter4, gate264inter5, gate264inter6, gate264inter7, gate264inter8, gate264inter9, gate264inter10, gate264inter11, gate264inter12, gate252inter0, gate252inter1, gate252inter2, gate252inter3, gate252inter4, gate252inter5, gate252inter6, gate252inter7, gate252inter8, gate252inter9, gate252inter10, gate252inter11, gate252inter12, gate12inter0, gate12inter1, gate12inter2, gate12inter3, gate12inter4, gate12inter5, gate12inter6, gate12inter7, gate12inter8, gate12inter9, gate12inter10, gate12inter11, gate12inter12, gate190inter0, gate190inter1, gate190inter2, gate190inter3, gate190inter4, gate190inter5, gate190inter6, gate190inter7, gate190inter8, gate190inter9, gate190inter10, gate190inter11, gate190inter12, gate207inter0, gate207inter1, gate207inter2, gate207inter3, gate207inter4, gate207inter5, gate207inter6, gate207inter7, gate207inter8, gate207inter9, gate207inter10, gate207inter11, gate207inter12, gate26inter0, gate26inter1, gate26inter2, gate26inter3, gate26inter4, gate26inter5, gate26inter6, gate26inter7, gate26inter8, gate26inter9, gate26inter10, gate26inter11, gate26inter12, gate131inter0, gate131inter1, gate131inter2, gate131inter3, gate131inter4, gate131inter5, gate131inter6, gate131inter7, gate131inter8, gate131inter9, gate131inter10, gate131inter11, gate131inter12, gate269inter0, gate269inter1, gate269inter2, gate269inter3, gate269inter4, gate269inter5, gate269inter6, gate269inter7, gate269inter8, gate269inter9, gate269inter10, gate269inter11, gate269inter12, gate438inter0, gate438inter1, gate438inter2, gate438inter3, gate438inter4, gate438inter5, gate438inter6, gate438inter7, gate438inter8, gate438inter9, gate438inter10, gate438inter11, gate438inter12, gate143inter0, gate143inter1, gate143inter2, gate143inter3, gate143inter4, gate143inter5, gate143inter6, gate143inter7, gate143inter8, gate143inter9, gate143inter10, gate143inter11, gate143inter12, gate491inter0, gate491inter1, gate491inter2, gate491inter3, gate491inter4, gate491inter5, gate491inter6, gate491inter7, gate491inter8, gate491inter9, gate491inter10, gate491inter11, gate491inter12, gate11inter0, gate11inter1, gate11inter2, gate11inter3, gate11inter4, gate11inter5, gate11inter6, gate11inter7, gate11inter8, gate11inter9, gate11inter10, gate11inter11, gate11inter12, gate265inter0, gate265inter1, gate265inter2, gate265inter3, gate265inter4, gate265inter5, gate265inter6, gate265inter7, gate265inter8, gate265inter9, gate265inter10, gate265inter11, gate265inter12, gate428inter0, gate428inter1, gate428inter2, gate428inter3, gate428inter4, gate428inter5, gate428inter6, gate428inter7, gate428inter8, gate428inter9, gate428inter10, gate428inter11, gate428inter12, gate452inter0, gate452inter1, gate452inter2, gate452inter3, gate452inter4, gate452inter5, gate452inter6, gate452inter7, gate452inter8, gate452inter9, gate452inter10, gate452inter11, gate452inter12, gate57inter0, gate57inter1, gate57inter2, gate57inter3, gate57inter4, gate57inter5, gate57inter6, gate57inter7, gate57inter8, gate57inter9, gate57inter10, gate57inter11, gate57inter12, gate126inter0, gate126inter1, gate126inter2, gate126inter3, gate126inter4, gate126inter5, gate126inter6, gate126inter7, gate126inter8, gate126inter9, gate126inter10, gate126inter11, gate126inter12, gate119inter0, gate119inter1, gate119inter2, gate119inter3, gate119inter4, gate119inter5, gate119inter6, gate119inter7, gate119inter8, gate119inter9, gate119inter10, gate119inter11, gate119inter12, gate232inter0, gate232inter1, gate232inter2, gate232inter3, gate232inter4, gate232inter5, gate232inter6, gate232inter7, gate232inter8, gate232inter9, gate232inter10, gate232inter11, gate232inter12, gate206inter0, gate206inter1, gate206inter2, gate206inter3, gate206inter4, gate206inter5, gate206inter6, gate206inter7, gate206inter8, gate206inter9, gate206inter10, gate206inter11, gate206inter12, gate67inter0, gate67inter1, gate67inter2, gate67inter3, gate67inter4, gate67inter5, gate67inter6, gate67inter7, gate67inter8, gate67inter9, gate67inter10, gate67inter11, gate67inter12, gate473inter0, gate473inter1, gate473inter2, gate473inter3, gate473inter4, gate473inter5, gate473inter6, gate473inter7, gate473inter8, gate473inter9, gate473inter10, gate473inter11, gate473inter12, gate193inter0, gate193inter1, gate193inter2, gate193inter3, gate193inter4, gate193inter5, gate193inter6, gate193inter7, gate193inter8, gate193inter9, gate193inter10, gate193inter11, gate193inter12, gate421inter0, gate421inter1, gate421inter2, gate421inter3, gate421inter4, gate421inter5, gate421inter6, gate421inter7, gate421inter8, gate421inter9, gate421inter10, gate421inter11, gate421inter12, gate226inter0, gate226inter1, gate226inter2, gate226inter3, gate226inter4, gate226inter5, gate226inter6, gate226inter7, gate226inter8, gate226inter9, gate226inter10, gate226inter11, gate226inter12, gate464inter0, gate464inter1, gate464inter2, gate464inter3, gate464inter4, gate464inter5, gate464inter6, gate464inter7, gate464inter8, gate464inter9, gate464inter10, gate464inter11, gate464inter12, gate70inter0, gate70inter1, gate70inter2, gate70inter3, gate70inter4, gate70inter5, gate70inter6, gate70inter7, gate70inter8, gate70inter9, gate70inter10, gate70inter11, gate70inter12, gate274inter0, gate274inter1, gate274inter2, gate274inter3, gate274inter4, gate274inter5, gate274inter6, gate274inter7, gate274inter8, gate274inter9, gate274inter10, gate274inter11, gate274inter12, gate236inter0, gate236inter1, gate236inter2, gate236inter3, gate236inter4, gate236inter5, gate236inter6, gate236inter7, gate236inter8, gate236inter9, gate236inter10, gate236inter11, gate236inter12, gate261inter0, gate261inter1, gate261inter2, gate261inter3, gate261inter4, gate261inter5, gate261inter6, gate261inter7, gate261inter8, gate261inter9, gate261inter10, gate261inter11, gate261inter12, gate195inter0, gate195inter1, gate195inter2, gate195inter3, gate195inter4, gate195inter5, gate195inter6, gate195inter7, gate195inter8, gate195inter9, gate195inter10, gate195inter11, gate195inter12, gate440inter0, gate440inter1, gate440inter2, gate440inter3, gate440inter4, gate440inter5, gate440inter6, gate440inter7, gate440inter8, gate440inter9, gate440inter10, gate440inter11, gate440inter12, gate466inter0, gate466inter1, gate466inter2, gate466inter3, gate466inter4, gate466inter5, gate466inter6, gate466inter7, gate466inter8, gate466inter9, gate466inter10, gate466inter11, gate466inter12, gate495inter0, gate495inter1, gate495inter2, gate495inter3, gate495inter4, gate495inter5, gate495inter6, gate495inter7, gate495inter8, gate495inter9, gate495inter10, gate495inter11, gate495inter12;



and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );
nand2 gate9( .a(G1), .b(G2), .O(G266) );
nand2 gate10( .a(G3), .b(G4), .O(G269) );

  xor2  gate2339(.a(G6), .b(G5), .O(gate11inter0));
  nand2 gate2340(.a(gate11inter0), .b(s_256), .O(gate11inter1));
  and2  gate2341(.a(G6), .b(G5), .O(gate11inter2));
  inv1  gate2342(.a(s_256), .O(gate11inter3));
  inv1  gate2343(.a(s_257), .O(gate11inter4));
  nand2 gate2344(.a(gate11inter4), .b(gate11inter3), .O(gate11inter5));
  nor2  gate2345(.a(gate11inter5), .b(gate11inter2), .O(gate11inter6));
  inv1  gate2346(.a(G5), .O(gate11inter7));
  inv1  gate2347(.a(G6), .O(gate11inter8));
  nand2 gate2348(.a(gate11inter8), .b(gate11inter7), .O(gate11inter9));
  nand2 gate2349(.a(s_257), .b(gate11inter3), .O(gate11inter10));
  nor2  gate2350(.a(gate11inter10), .b(gate11inter9), .O(gate11inter11));
  nor2  gate2351(.a(gate11inter11), .b(gate11inter6), .O(gate11inter12));
  nand2 gate2352(.a(gate11inter12), .b(gate11inter1), .O(G272));

  xor2  gate2213(.a(G8), .b(G7), .O(gate12inter0));
  nand2 gate2214(.a(gate12inter0), .b(s_238), .O(gate12inter1));
  and2  gate2215(.a(G8), .b(G7), .O(gate12inter2));
  inv1  gate2216(.a(s_238), .O(gate12inter3));
  inv1  gate2217(.a(s_239), .O(gate12inter4));
  nand2 gate2218(.a(gate12inter4), .b(gate12inter3), .O(gate12inter5));
  nor2  gate2219(.a(gate12inter5), .b(gate12inter2), .O(gate12inter6));
  inv1  gate2220(.a(G7), .O(gate12inter7));
  inv1  gate2221(.a(G8), .O(gate12inter8));
  nand2 gate2222(.a(gate12inter8), .b(gate12inter7), .O(gate12inter9));
  nand2 gate2223(.a(s_239), .b(gate12inter3), .O(gate12inter10));
  nor2  gate2224(.a(gate12inter10), .b(gate12inter9), .O(gate12inter11));
  nor2  gate2225(.a(gate12inter11), .b(gate12inter6), .O(gate12inter12));
  nand2 gate2226(.a(gate12inter12), .b(gate12inter1), .O(G275));

  xor2  gate659(.a(G10), .b(G9), .O(gate13inter0));
  nand2 gate660(.a(gate13inter0), .b(s_16), .O(gate13inter1));
  and2  gate661(.a(G10), .b(G9), .O(gate13inter2));
  inv1  gate662(.a(s_16), .O(gate13inter3));
  inv1  gate663(.a(s_17), .O(gate13inter4));
  nand2 gate664(.a(gate13inter4), .b(gate13inter3), .O(gate13inter5));
  nor2  gate665(.a(gate13inter5), .b(gate13inter2), .O(gate13inter6));
  inv1  gate666(.a(G9), .O(gate13inter7));
  inv1  gate667(.a(G10), .O(gate13inter8));
  nand2 gate668(.a(gate13inter8), .b(gate13inter7), .O(gate13inter9));
  nand2 gate669(.a(s_17), .b(gate13inter3), .O(gate13inter10));
  nor2  gate670(.a(gate13inter10), .b(gate13inter9), .O(gate13inter11));
  nor2  gate671(.a(gate13inter11), .b(gate13inter6), .O(gate13inter12));
  nand2 gate672(.a(gate13inter12), .b(gate13inter1), .O(G278));
nand2 gate14( .a(G11), .b(G12), .O(G281) );

  xor2  gate1401(.a(G14), .b(G13), .O(gate15inter0));
  nand2 gate1402(.a(gate15inter0), .b(s_122), .O(gate15inter1));
  and2  gate1403(.a(G14), .b(G13), .O(gate15inter2));
  inv1  gate1404(.a(s_122), .O(gate15inter3));
  inv1  gate1405(.a(s_123), .O(gate15inter4));
  nand2 gate1406(.a(gate15inter4), .b(gate15inter3), .O(gate15inter5));
  nor2  gate1407(.a(gate15inter5), .b(gate15inter2), .O(gate15inter6));
  inv1  gate1408(.a(G13), .O(gate15inter7));
  inv1  gate1409(.a(G14), .O(gate15inter8));
  nand2 gate1410(.a(gate15inter8), .b(gate15inter7), .O(gate15inter9));
  nand2 gate1411(.a(s_123), .b(gate15inter3), .O(gate15inter10));
  nor2  gate1412(.a(gate15inter10), .b(gate15inter9), .O(gate15inter11));
  nor2  gate1413(.a(gate15inter11), .b(gate15inter6), .O(gate15inter12));
  nand2 gate1414(.a(gate15inter12), .b(gate15inter1), .O(G284));
nand2 gate16( .a(G15), .b(G16), .O(G287) );

  xor2  gate617(.a(G18), .b(G17), .O(gate17inter0));
  nand2 gate618(.a(gate17inter0), .b(s_10), .O(gate17inter1));
  and2  gate619(.a(G18), .b(G17), .O(gate17inter2));
  inv1  gate620(.a(s_10), .O(gate17inter3));
  inv1  gate621(.a(s_11), .O(gate17inter4));
  nand2 gate622(.a(gate17inter4), .b(gate17inter3), .O(gate17inter5));
  nor2  gate623(.a(gate17inter5), .b(gate17inter2), .O(gate17inter6));
  inv1  gate624(.a(G17), .O(gate17inter7));
  inv1  gate625(.a(G18), .O(gate17inter8));
  nand2 gate626(.a(gate17inter8), .b(gate17inter7), .O(gate17inter9));
  nand2 gate627(.a(s_11), .b(gate17inter3), .O(gate17inter10));
  nor2  gate628(.a(gate17inter10), .b(gate17inter9), .O(gate17inter11));
  nor2  gate629(.a(gate17inter11), .b(gate17inter6), .O(gate17inter12));
  nand2 gate630(.a(gate17inter12), .b(gate17inter1), .O(G290));
nand2 gate18( .a(G19), .b(G20), .O(G293) );
nand2 gate19( .a(G21), .b(G22), .O(G296) );
nand2 gate20( .a(G23), .b(G24), .O(G299) );
nand2 gate21( .a(G25), .b(G26), .O(G302) );

  xor2  gate841(.a(G28), .b(G27), .O(gate22inter0));
  nand2 gate842(.a(gate22inter0), .b(s_42), .O(gate22inter1));
  and2  gate843(.a(G28), .b(G27), .O(gate22inter2));
  inv1  gate844(.a(s_42), .O(gate22inter3));
  inv1  gate845(.a(s_43), .O(gate22inter4));
  nand2 gate846(.a(gate22inter4), .b(gate22inter3), .O(gate22inter5));
  nor2  gate847(.a(gate22inter5), .b(gate22inter2), .O(gate22inter6));
  inv1  gate848(.a(G27), .O(gate22inter7));
  inv1  gate849(.a(G28), .O(gate22inter8));
  nand2 gate850(.a(gate22inter8), .b(gate22inter7), .O(gate22inter9));
  nand2 gate851(.a(s_43), .b(gate22inter3), .O(gate22inter10));
  nor2  gate852(.a(gate22inter10), .b(gate22inter9), .O(gate22inter11));
  nor2  gate853(.a(gate22inter11), .b(gate22inter6), .O(gate22inter12));
  nand2 gate854(.a(gate22inter12), .b(gate22inter1), .O(G305));
nand2 gate23( .a(G29), .b(G30), .O(G308) );

  xor2  gate1737(.a(G32), .b(G31), .O(gate24inter0));
  nand2 gate1738(.a(gate24inter0), .b(s_170), .O(gate24inter1));
  and2  gate1739(.a(G32), .b(G31), .O(gate24inter2));
  inv1  gate1740(.a(s_170), .O(gate24inter3));
  inv1  gate1741(.a(s_171), .O(gate24inter4));
  nand2 gate1742(.a(gate24inter4), .b(gate24inter3), .O(gate24inter5));
  nor2  gate1743(.a(gate24inter5), .b(gate24inter2), .O(gate24inter6));
  inv1  gate1744(.a(G31), .O(gate24inter7));
  inv1  gate1745(.a(G32), .O(gate24inter8));
  nand2 gate1746(.a(gate24inter8), .b(gate24inter7), .O(gate24inter9));
  nand2 gate1747(.a(s_171), .b(gate24inter3), .O(gate24inter10));
  nor2  gate1748(.a(gate24inter10), .b(gate24inter9), .O(gate24inter11));
  nor2  gate1749(.a(gate24inter11), .b(gate24inter6), .O(gate24inter12));
  nand2 gate1750(.a(gate24inter12), .b(gate24inter1), .O(G311));
nand2 gate25( .a(G1), .b(G5), .O(G314) );

  xor2  gate2255(.a(G13), .b(G9), .O(gate26inter0));
  nand2 gate2256(.a(gate26inter0), .b(s_244), .O(gate26inter1));
  and2  gate2257(.a(G13), .b(G9), .O(gate26inter2));
  inv1  gate2258(.a(s_244), .O(gate26inter3));
  inv1  gate2259(.a(s_245), .O(gate26inter4));
  nand2 gate2260(.a(gate26inter4), .b(gate26inter3), .O(gate26inter5));
  nor2  gate2261(.a(gate26inter5), .b(gate26inter2), .O(gate26inter6));
  inv1  gate2262(.a(G9), .O(gate26inter7));
  inv1  gate2263(.a(G13), .O(gate26inter8));
  nand2 gate2264(.a(gate26inter8), .b(gate26inter7), .O(gate26inter9));
  nand2 gate2265(.a(s_245), .b(gate26inter3), .O(gate26inter10));
  nor2  gate2266(.a(gate26inter10), .b(gate26inter9), .O(gate26inter11));
  nor2  gate2267(.a(gate26inter11), .b(gate26inter6), .O(gate26inter12));
  nand2 gate2268(.a(gate26inter12), .b(gate26inter1), .O(G317));
nand2 gate27( .a(G2), .b(G6), .O(G320) );
nand2 gate28( .a(G10), .b(G14), .O(G323) );
nand2 gate29( .a(G3), .b(G7), .O(G326) );
nand2 gate30( .a(G11), .b(G15), .O(G329) );
nand2 gate31( .a(G4), .b(G8), .O(G332) );

  xor2  gate939(.a(G16), .b(G12), .O(gate32inter0));
  nand2 gate940(.a(gate32inter0), .b(s_56), .O(gate32inter1));
  and2  gate941(.a(G16), .b(G12), .O(gate32inter2));
  inv1  gate942(.a(s_56), .O(gate32inter3));
  inv1  gate943(.a(s_57), .O(gate32inter4));
  nand2 gate944(.a(gate32inter4), .b(gate32inter3), .O(gate32inter5));
  nor2  gate945(.a(gate32inter5), .b(gate32inter2), .O(gate32inter6));
  inv1  gate946(.a(G12), .O(gate32inter7));
  inv1  gate947(.a(G16), .O(gate32inter8));
  nand2 gate948(.a(gate32inter8), .b(gate32inter7), .O(gate32inter9));
  nand2 gate949(.a(s_57), .b(gate32inter3), .O(gate32inter10));
  nor2  gate950(.a(gate32inter10), .b(gate32inter9), .O(gate32inter11));
  nor2  gate951(.a(gate32inter11), .b(gate32inter6), .O(gate32inter12));
  nand2 gate952(.a(gate32inter12), .b(gate32inter1), .O(G335));
nand2 gate33( .a(G17), .b(G21), .O(G338) );

  xor2  gate2171(.a(G29), .b(G25), .O(gate34inter0));
  nand2 gate2172(.a(gate34inter0), .b(s_232), .O(gate34inter1));
  and2  gate2173(.a(G29), .b(G25), .O(gate34inter2));
  inv1  gate2174(.a(s_232), .O(gate34inter3));
  inv1  gate2175(.a(s_233), .O(gate34inter4));
  nand2 gate2176(.a(gate34inter4), .b(gate34inter3), .O(gate34inter5));
  nor2  gate2177(.a(gate34inter5), .b(gate34inter2), .O(gate34inter6));
  inv1  gate2178(.a(G25), .O(gate34inter7));
  inv1  gate2179(.a(G29), .O(gate34inter8));
  nand2 gate2180(.a(gate34inter8), .b(gate34inter7), .O(gate34inter9));
  nand2 gate2181(.a(s_233), .b(gate34inter3), .O(gate34inter10));
  nor2  gate2182(.a(gate34inter10), .b(gate34inter9), .O(gate34inter11));
  nor2  gate2183(.a(gate34inter11), .b(gate34inter6), .O(gate34inter12));
  nand2 gate2184(.a(gate34inter12), .b(gate34inter1), .O(G341));

  xor2  gate1261(.a(G22), .b(G18), .O(gate35inter0));
  nand2 gate1262(.a(gate35inter0), .b(s_102), .O(gate35inter1));
  and2  gate1263(.a(G22), .b(G18), .O(gate35inter2));
  inv1  gate1264(.a(s_102), .O(gate35inter3));
  inv1  gate1265(.a(s_103), .O(gate35inter4));
  nand2 gate1266(.a(gate35inter4), .b(gate35inter3), .O(gate35inter5));
  nor2  gate1267(.a(gate35inter5), .b(gate35inter2), .O(gate35inter6));
  inv1  gate1268(.a(G18), .O(gate35inter7));
  inv1  gate1269(.a(G22), .O(gate35inter8));
  nand2 gate1270(.a(gate35inter8), .b(gate35inter7), .O(gate35inter9));
  nand2 gate1271(.a(s_103), .b(gate35inter3), .O(gate35inter10));
  nor2  gate1272(.a(gate35inter10), .b(gate35inter9), .O(gate35inter11));
  nor2  gate1273(.a(gate35inter11), .b(gate35inter6), .O(gate35inter12));
  nand2 gate1274(.a(gate35inter12), .b(gate35inter1), .O(G344));
nand2 gate36( .a(G26), .b(G30), .O(G347) );
nand2 gate37( .a(G19), .b(G23), .O(G350) );

  xor2  gate2045(.a(G31), .b(G27), .O(gate38inter0));
  nand2 gate2046(.a(gate38inter0), .b(s_214), .O(gate38inter1));
  and2  gate2047(.a(G31), .b(G27), .O(gate38inter2));
  inv1  gate2048(.a(s_214), .O(gate38inter3));
  inv1  gate2049(.a(s_215), .O(gate38inter4));
  nand2 gate2050(.a(gate38inter4), .b(gate38inter3), .O(gate38inter5));
  nor2  gate2051(.a(gate38inter5), .b(gate38inter2), .O(gate38inter6));
  inv1  gate2052(.a(G27), .O(gate38inter7));
  inv1  gate2053(.a(G31), .O(gate38inter8));
  nand2 gate2054(.a(gate38inter8), .b(gate38inter7), .O(gate38inter9));
  nand2 gate2055(.a(s_215), .b(gate38inter3), .O(gate38inter10));
  nor2  gate2056(.a(gate38inter10), .b(gate38inter9), .O(gate38inter11));
  nor2  gate2057(.a(gate38inter11), .b(gate38inter6), .O(gate38inter12));
  nand2 gate2058(.a(gate38inter12), .b(gate38inter1), .O(G353));
nand2 gate39( .a(G20), .b(G24), .O(G356) );
nand2 gate40( .a(G28), .b(G32), .O(G359) );
nand2 gate41( .a(G1), .b(G266), .O(G362) );
nand2 gate42( .a(G2), .b(G266), .O(G363) );

  xor2  gate2129(.a(G269), .b(G3), .O(gate43inter0));
  nand2 gate2130(.a(gate43inter0), .b(s_226), .O(gate43inter1));
  and2  gate2131(.a(G269), .b(G3), .O(gate43inter2));
  inv1  gate2132(.a(s_226), .O(gate43inter3));
  inv1  gate2133(.a(s_227), .O(gate43inter4));
  nand2 gate2134(.a(gate43inter4), .b(gate43inter3), .O(gate43inter5));
  nor2  gate2135(.a(gate43inter5), .b(gate43inter2), .O(gate43inter6));
  inv1  gate2136(.a(G3), .O(gate43inter7));
  inv1  gate2137(.a(G269), .O(gate43inter8));
  nand2 gate2138(.a(gate43inter8), .b(gate43inter7), .O(gate43inter9));
  nand2 gate2139(.a(s_227), .b(gate43inter3), .O(gate43inter10));
  nor2  gate2140(.a(gate43inter10), .b(gate43inter9), .O(gate43inter11));
  nor2  gate2141(.a(gate43inter11), .b(gate43inter6), .O(gate43inter12));
  nand2 gate2142(.a(gate43inter12), .b(gate43inter1), .O(G364));

  xor2  gate1905(.a(G269), .b(G4), .O(gate44inter0));
  nand2 gate1906(.a(gate44inter0), .b(s_194), .O(gate44inter1));
  and2  gate1907(.a(G269), .b(G4), .O(gate44inter2));
  inv1  gate1908(.a(s_194), .O(gate44inter3));
  inv1  gate1909(.a(s_195), .O(gate44inter4));
  nand2 gate1910(.a(gate44inter4), .b(gate44inter3), .O(gate44inter5));
  nor2  gate1911(.a(gate44inter5), .b(gate44inter2), .O(gate44inter6));
  inv1  gate1912(.a(G4), .O(gate44inter7));
  inv1  gate1913(.a(G269), .O(gate44inter8));
  nand2 gate1914(.a(gate44inter8), .b(gate44inter7), .O(gate44inter9));
  nand2 gate1915(.a(s_195), .b(gate44inter3), .O(gate44inter10));
  nor2  gate1916(.a(gate44inter10), .b(gate44inter9), .O(gate44inter11));
  nor2  gate1917(.a(gate44inter11), .b(gate44inter6), .O(gate44inter12));
  nand2 gate1918(.a(gate44inter12), .b(gate44inter1), .O(G365));
nand2 gate45( .a(G5), .b(G272), .O(G366) );
nand2 gate46( .a(G6), .b(G272), .O(G367) );
nand2 gate47( .a(G7), .b(G275), .O(G368) );

  xor2  gate1079(.a(G275), .b(G8), .O(gate48inter0));
  nand2 gate1080(.a(gate48inter0), .b(s_76), .O(gate48inter1));
  and2  gate1081(.a(G275), .b(G8), .O(gate48inter2));
  inv1  gate1082(.a(s_76), .O(gate48inter3));
  inv1  gate1083(.a(s_77), .O(gate48inter4));
  nand2 gate1084(.a(gate48inter4), .b(gate48inter3), .O(gate48inter5));
  nor2  gate1085(.a(gate48inter5), .b(gate48inter2), .O(gate48inter6));
  inv1  gate1086(.a(G8), .O(gate48inter7));
  inv1  gate1087(.a(G275), .O(gate48inter8));
  nand2 gate1088(.a(gate48inter8), .b(gate48inter7), .O(gate48inter9));
  nand2 gate1089(.a(s_77), .b(gate48inter3), .O(gate48inter10));
  nor2  gate1090(.a(gate48inter10), .b(gate48inter9), .O(gate48inter11));
  nor2  gate1091(.a(gate48inter11), .b(gate48inter6), .O(gate48inter12));
  nand2 gate1092(.a(gate48inter12), .b(gate48inter1), .O(G369));
nand2 gate49( .a(G9), .b(G278), .O(G370) );
nand2 gate50( .a(G10), .b(G278), .O(G371) );
nand2 gate51( .a(G11), .b(G281), .O(G372) );
nand2 gate52( .a(G12), .b(G281), .O(G373) );
nand2 gate53( .a(G13), .b(G284), .O(G374) );
nand2 gate54( .a(G14), .b(G284), .O(G375) );
nand2 gate55( .a(G15), .b(G287), .O(G376) );
nand2 gate56( .a(G16), .b(G287), .O(G377) );

  xor2  gate2395(.a(G290), .b(G17), .O(gate57inter0));
  nand2 gate2396(.a(gate57inter0), .b(s_264), .O(gate57inter1));
  and2  gate2397(.a(G290), .b(G17), .O(gate57inter2));
  inv1  gate2398(.a(s_264), .O(gate57inter3));
  inv1  gate2399(.a(s_265), .O(gate57inter4));
  nand2 gate2400(.a(gate57inter4), .b(gate57inter3), .O(gate57inter5));
  nor2  gate2401(.a(gate57inter5), .b(gate57inter2), .O(gate57inter6));
  inv1  gate2402(.a(G17), .O(gate57inter7));
  inv1  gate2403(.a(G290), .O(gate57inter8));
  nand2 gate2404(.a(gate57inter8), .b(gate57inter7), .O(gate57inter9));
  nand2 gate2405(.a(s_265), .b(gate57inter3), .O(gate57inter10));
  nor2  gate2406(.a(gate57inter10), .b(gate57inter9), .O(gate57inter11));
  nor2  gate2407(.a(gate57inter11), .b(gate57inter6), .O(gate57inter12));
  nand2 gate2408(.a(gate57inter12), .b(gate57inter1), .O(G378));
nand2 gate58( .a(G18), .b(G290), .O(G379) );
nand2 gate59( .a(G19), .b(G293), .O(G380) );

  xor2  gate1303(.a(G293), .b(G20), .O(gate60inter0));
  nand2 gate1304(.a(gate60inter0), .b(s_108), .O(gate60inter1));
  and2  gate1305(.a(G293), .b(G20), .O(gate60inter2));
  inv1  gate1306(.a(s_108), .O(gate60inter3));
  inv1  gate1307(.a(s_109), .O(gate60inter4));
  nand2 gate1308(.a(gate60inter4), .b(gate60inter3), .O(gate60inter5));
  nor2  gate1309(.a(gate60inter5), .b(gate60inter2), .O(gate60inter6));
  inv1  gate1310(.a(G20), .O(gate60inter7));
  inv1  gate1311(.a(G293), .O(gate60inter8));
  nand2 gate1312(.a(gate60inter8), .b(gate60inter7), .O(gate60inter9));
  nand2 gate1313(.a(s_109), .b(gate60inter3), .O(gate60inter10));
  nor2  gate1314(.a(gate60inter10), .b(gate60inter9), .O(gate60inter11));
  nor2  gate1315(.a(gate60inter11), .b(gate60inter6), .O(gate60inter12));
  nand2 gate1316(.a(gate60inter12), .b(gate60inter1), .O(G381));
nand2 gate61( .a(G21), .b(G296), .O(G382) );

  xor2  gate827(.a(G296), .b(G22), .O(gate62inter0));
  nand2 gate828(.a(gate62inter0), .b(s_40), .O(gate62inter1));
  and2  gate829(.a(G296), .b(G22), .O(gate62inter2));
  inv1  gate830(.a(s_40), .O(gate62inter3));
  inv1  gate831(.a(s_41), .O(gate62inter4));
  nand2 gate832(.a(gate62inter4), .b(gate62inter3), .O(gate62inter5));
  nor2  gate833(.a(gate62inter5), .b(gate62inter2), .O(gate62inter6));
  inv1  gate834(.a(G22), .O(gate62inter7));
  inv1  gate835(.a(G296), .O(gate62inter8));
  nand2 gate836(.a(gate62inter8), .b(gate62inter7), .O(gate62inter9));
  nand2 gate837(.a(s_41), .b(gate62inter3), .O(gate62inter10));
  nor2  gate838(.a(gate62inter10), .b(gate62inter9), .O(gate62inter11));
  nor2  gate839(.a(gate62inter11), .b(gate62inter6), .O(gate62inter12));
  nand2 gate840(.a(gate62inter12), .b(gate62inter1), .O(G383));
nand2 gate63( .a(G23), .b(G299), .O(G384) );

  xor2  gate1751(.a(G299), .b(G24), .O(gate64inter0));
  nand2 gate1752(.a(gate64inter0), .b(s_172), .O(gate64inter1));
  and2  gate1753(.a(G299), .b(G24), .O(gate64inter2));
  inv1  gate1754(.a(s_172), .O(gate64inter3));
  inv1  gate1755(.a(s_173), .O(gate64inter4));
  nand2 gate1756(.a(gate64inter4), .b(gate64inter3), .O(gate64inter5));
  nor2  gate1757(.a(gate64inter5), .b(gate64inter2), .O(gate64inter6));
  inv1  gate1758(.a(G24), .O(gate64inter7));
  inv1  gate1759(.a(G299), .O(gate64inter8));
  nand2 gate1760(.a(gate64inter8), .b(gate64inter7), .O(gate64inter9));
  nand2 gate1761(.a(s_173), .b(gate64inter3), .O(gate64inter10));
  nor2  gate1762(.a(gate64inter10), .b(gate64inter9), .O(gate64inter11));
  nor2  gate1763(.a(gate64inter11), .b(gate64inter6), .O(gate64inter12));
  nand2 gate1764(.a(gate64inter12), .b(gate64inter1), .O(G385));

  xor2  gate715(.a(G302), .b(G25), .O(gate65inter0));
  nand2 gate716(.a(gate65inter0), .b(s_24), .O(gate65inter1));
  and2  gate717(.a(G302), .b(G25), .O(gate65inter2));
  inv1  gate718(.a(s_24), .O(gate65inter3));
  inv1  gate719(.a(s_25), .O(gate65inter4));
  nand2 gate720(.a(gate65inter4), .b(gate65inter3), .O(gate65inter5));
  nor2  gate721(.a(gate65inter5), .b(gate65inter2), .O(gate65inter6));
  inv1  gate722(.a(G25), .O(gate65inter7));
  inv1  gate723(.a(G302), .O(gate65inter8));
  nand2 gate724(.a(gate65inter8), .b(gate65inter7), .O(gate65inter9));
  nand2 gate725(.a(s_25), .b(gate65inter3), .O(gate65inter10));
  nor2  gate726(.a(gate65inter10), .b(gate65inter9), .O(gate65inter11));
  nor2  gate727(.a(gate65inter11), .b(gate65inter6), .O(gate65inter12));
  nand2 gate728(.a(gate65inter12), .b(gate65inter1), .O(G386));
nand2 gate66( .a(G26), .b(G302), .O(G387) );

  xor2  gate2465(.a(G305), .b(G27), .O(gate67inter0));
  nand2 gate2466(.a(gate67inter0), .b(s_274), .O(gate67inter1));
  and2  gate2467(.a(G305), .b(G27), .O(gate67inter2));
  inv1  gate2468(.a(s_274), .O(gate67inter3));
  inv1  gate2469(.a(s_275), .O(gate67inter4));
  nand2 gate2470(.a(gate67inter4), .b(gate67inter3), .O(gate67inter5));
  nor2  gate2471(.a(gate67inter5), .b(gate67inter2), .O(gate67inter6));
  inv1  gate2472(.a(G27), .O(gate67inter7));
  inv1  gate2473(.a(G305), .O(gate67inter8));
  nand2 gate2474(.a(gate67inter8), .b(gate67inter7), .O(gate67inter9));
  nand2 gate2475(.a(s_275), .b(gate67inter3), .O(gate67inter10));
  nor2  gate2476(.a(gate67inter10), .b(gate67inter9), .O(gate67inter11));
  nor2  gate2477(.a(gate67inter11), .b(gate67inter6), .O(gate67inter12));
  nand2 gate2478(.a(gate67inter12), .b(gate67inter1), .O(G388));

  xor2  gate1443(.a(G305), .b(G28), .O(gate68inter0));
  nand2 gate1444(.a(gate68inter0), .b(s_128), .O(gate68inter1));
  and2  gate1445(.a(G305), .b(G28), .O(gate68inter2));
  inv1  gate1446(.a(s_128), .O(gate68inter3));
  inv1  gate1447(.a(s_129), .O(gate68inter4));
  nand2 gate1448(.a(gate68inter4), .b(gate68inter3), .O(gate68inter5));
  nor2  gate1449(.a(gate68inter5), .b(gate68inter2), .O(gate68inter6));
  inv1  gate1450(.a(G28), .O(gate68inter7));
  inv1  gate1451(.a(G305), .O(gate68inter8));
  nand2 gate1452(.a(gate68inter8), .b(gate68inter7), .O(gate68inter9));
  nand2 gate1453(.a(s_129), .b(gate68inter3), .O(gate68inter10));
  nor2  gate1454(.a(gate68inter10), .b(gate68inter9), .O(gate68inter11));
  nor2  gate1455(.a(gate68inter11), .b(gate68inter6), .O(gate68inter12));
  nand2 gate1456(.a(gate68inter12), .b(gate68inter1), .O(G389));
nand2 gate69( .a(G29), .b(G308), .O(G390) );

  xor2  gate2549(.a(G308), .b(G30), .O(gate70inter0));
  nand2 gate2550(.a(gate70inter0), .b(s_286), .O(gate70inter1));
  and2  gate2551(.a(G308), .b(G30), .O(gate70inter2));
  inv1  gate2552(.a(s_286), .O(gate70inter3));
  inv1  gate2553(.a(s_287), .O(gate70inter4));
  nand2 gate2554(.a(gate70inter4), .b(gate70inter3), .O(gate70inter5));
  nor2  gate2555(.a(gate70inter5), .b(gate70inter2), .O(gate70inter6));
  inv1  gate2556(.a(G30), .O(gate70inter7));
  inv1  gate2557(.a(G308), .O(gate70inter8));
  nand2 gate2558(.a(gate70inter8), .b(gate70inter7), .O(gate70inter9));
  nand2 gate2559(.a(s_287), .b(gate70inter3), .O(gate70inter10));
  nor2  gate2560(.a(gate70inter10), .b(gate70inter9), .O(gate70inter11));
  nor2  gate2561(.a(gate70inter11), .b(gate70inter6), .O(gate70inter12));
  nand2 gate2562(.a(gate70inter12), .b(gate70inter1), .O(G391));
nand2 gate71( .a(G31), .b(G311), .O(G392) );
nand2 gate72( .a(G32), .b(G311), .O(G393) );
nand2 gate73( .a(G1), .b(G314), .O(G394) );
nand2 gate74( .a(G5), .b(G314), .O(G395) );

  xor2  gate701(.a(G317), .b(G9), .O(gate75inter0));
  nand2 gate702(.a(gate75inter0), .b(s_22), .O(gate75inter1));
  and2  gate703(.a(G317), .b(G9), .O(gate75inter2));
  inv1  gate704(.a(s_22), .O(gate75inter3));
  inv1  gate705(.a(s_23), .O(gate75inter4));
  nand2 gate706(.a(gate75inter4), .b(gate75inter3), .O(gate75inter5));
  nor2  gate707(.a(gate75inter5), .b(gate75inter2), .O(gate75inter6));
  inv1  gate708(.a(G9), .O(gate75inter7));
  inv1  gate709(.a(G317), .O(gate75inter8));
  nand2 gate710(.a(gate75inter8), .b(gate75inter7), .O(gate75inter9));
  nand2 gate711(.a(s_23), .b(gate75inter3), .O(gate75inter10));
  nor2  gate712(.a(gate75inter10), .b(gate75inter9), .O(gate75inter11));
  nor2  gate713(.a(gate75inter11), .b(gate75inter6), .O(gate75inter12));
  nand2 gate714(.a(gate75inter12), .b(gate75inter1), .O(G396));

  xor2  gate1569(.a(G317), .b(G13), .O(gate76inter0));
  nand2 gate1570(.a(gate76inter0), .b(s_146), .O(gate76inter1));
  and2  gate1571(.a(G317), .b(G13), .O(gate76inter2));
  inv1  gate1572(.a(s_146), .O(gate76inter3));
  inv1  gate1573(.a(s_147), .O(gate76inter4));
  nand2 gate1574(.a(gate76inter4), .b(gate76inter3), .O(gate76inter5));
  nor2  gate1575(.a(gate76inter5), .b(gate76inter2), .O(gate76inter6));
  inv1  gate1576(.a(G13), .O(gate76inter7));
  inv1  gate1577(.a(G317), .O(gate76inter8));
  nand2 gate1578(.a(gate76inter8), .b(gate76inter7), .O(gate76inter9));
  nand2 gate1579(.a(s_147), .b(gate76inter3), .O(gate76inter10));
  nor2  gate1580(.a(gate76inter10), .b(gate76inter9), .O(gate76inter11));
  nor2  gate1581(.a(gate76inter11), .b(gate76inter6), .O(gate76inter12));
  nand2 gate1582(.a(gate76inter12), .b(gate76inter1), .O(G397));
nand2 gate77( .a(G2), .b(G320), .O(G398) );
nand2 gate78( .a(G6), .b(G320), .O(G399) );
nand2 gate79( .a(G10), .b(G323), .O(G400) );
nand2 gate80( .a(G14), .b(G323), .O(G401) );
nand2 gate81( .a(G3), .b(G326), .O(G402) );

  xor2  gate1765(.a(G326), .b(G7), .O(gate82inter0));
  nand2 gate1766(.a(gate82inter0), .b(s_174), .O(gate82inter1));
  and2  gate1767(.a(G326), .b(G7), .O(gate82inter2));
  inv1  gate1768(.a(s_174), .O(gate82inter3));
  inv1  gate1769(.a(s_175), .O(gate82inter4));
  nand2 gate1770(.a(gate82inter4), .b(gate82inter3), .O(gate82inter5));
  nor2  gate1771(.a(gate82inter5), .b(gate82inter2), .O(gate82inter6));
  inv1  gate1772(.a(G7), .O(gate82inter7));
  inv1  gate1773(.a(G326), .O(gate82inter8));
  nand2 gate1774(.a(gate82inter8), .b(gate82inter7), .O(gate82inter9));
  nand2 gate1775(.a(s_175), .b(gate82inter3), .O(gate82inter10));
  nor2  gate1776(.a(gate82inter10), .b(gate82inter9), .O(gate82inter11));
  nor2  gate1777(.a(gate82inter11), .b(gate82inter6), .O(gate82inter12));
  nand2 gate1778(.a(gate82inter12), .b(gate82inter1), .O(G403));
nand2 gate83( .a(G11), .b(G329), .O(G404) );

  xor2  gate855(.a(G329), .b(G15), .O(gate84inter0));
  nand2 gate856(.a(gate84inter0), .b(s_44), .O(gate84inter1));
  and2  gate857(.a(G329), .b(G15), .O(gate84inter2));
  inv1  gate858(.a(s_44), .O(gate84inter3));
  inv1  gate859(.a(s_45), .O(gate84inter4));
  nand2 gate860(.a(gate84inter4), .b(gate84inter3), .O(gate84inter5));
  nor2  gate861(.a(gate84inter5), .b(gate84inter2), .O(gate84inter6));
  inv1  gate862(.a(G15), .O(gate84inter7));
  inv1  gate863(.a(G329), .O(gate84inter8));
  nand2 gate864(.a(gate84inter8), .b(gate84inter7), .O(gate84inter9));
  nand2 gate865(.a(s_45), .b(gate84inter3), .O(gate84inter10));
  nor2  gate866(.a(gate84inter10), .b(gate84inter9), .O(gate84inter11));
  nor2  gate867(.a(gate84inter11), .b(gate84inter6), .O(gate84inter12));
  nand2 gate868(.a(gate84inter12), .b(gate84inter1), .O(G405));

  xor2  gate631(.a(G332), .b(G4), .O(gate85inter0));
  nand2 gate632(.a(gate85inter0), .b(s_12), .O(gate85inter1));
  and2  gate633(.a(G332), .b(G4), .O(gate85inter2));
  inv1  gate634(.a(s_12), .O(gate85inter3));
  inv1  gate635(.a(s_13), .O(gate85inter4));
  nand2 gate636(.a(gate85inter4), .b(gate85inter3), .O(gate85inter5));
  nor2  gate637(.a(gate85inter5), .b(gate85inter2), .O(gate85inter6));
  inv1  gate638(.a(G4), .O(gate85inter7));
  inv1  gate639(.a(G332), .O(gate85inter8));
  nand2 gate640(.a(gate85inter8), .b(gate85inter7), .O(gate85inter9));
  nand2 gate641(.a(s_13), .b(gate85inter3), .O(gate85inter10));
  nor2  gate642(.a(gate85inter10), .b(gate85inter9), .O(gate85inter11));
  nor2  gate643(.a(gate85inter11), .b(gate85inter6), .O(gate85inter12));
  nand2 gate644(.a(gate85inter12), .b(gate85inter1), .O(G406));

  xor2  gate1919(.a(G332), .b(G8), .O(gate86inter0));
  nand2 gate1920(.a(gate86inter0), .b(s_196), .O(gate86inter1));
  and2  gate1921(.a(G332), .b(G8), .O(gate86inter2));
  inv1  gate1922(.a(s_196), .O(gate86inter3));
  inv1  gate1923(.a(s_197), .O(gate86inter4));
  nand2 gate1924(.a(gate86inter4), .b(gate86inter3), .O(gate86inter5));
  nor2  gate1925(.a(gate86inter5), .b(gate86inter2), .O(gate86inter6));
  inv1  gate1926(.a(G8), .O(gate86inter7));
  inv1  gate1927(.a(G332), .O(gate86inter8));
  nand2 gate1928(.a(gate86inter8), .b(gate86inter7), .O(gate86inter9));
  nand2 gate1929(.a(s_197), .b(gate86inter3), .O(gate86inter10));
  nor2  gate1930(.a(gate86inter10), .b(gate86inter9), .O(gate86inter11));
  nor2  gate1931(.a(gate86inter11), .b(gate86inter6), .O(gate86inter12));
  nand2 gate1932(.a(gate86inter12), .b(gate86inter1), .O(G407));
nand2 gate87( .a(G12), .b(G335), .O(G408) );
nand2 gate88( .a(G16), .b(G335), .O(G409) );
nand2 gate89( .a(G17), .b(G338), .O(G410) );

  xor2  gate2143(.a(G338), .b(G21), .O(gate90inter0));
  nand2 gate2144(.a(gate90inter0), .b(s_228), .O(gate90inter1));
  and2  gate2145(.a(G338), .b(G21), .O(gate90inter2));
  inv1  gate2146(.a(s_228), .O(gate90inter3));
  inv1  gate2147(.a(s_229), .O(gate90inter4));
  nand2 gate2148(.a(gate90inter4), .b(gate90inter3), .O(gate90inter5));
  nor2  gate2149(.a(gate90inter5), .b(gate90inter2), .O(gate90inter6));
  inv1  gate2150(.a(G21), .O(gate90inter7));
  inv1  gate2151(.a(G338), .O(gate90inter8));
  nand2 gate2152(.a(gate90inter8), .b(gate90inter7), .O(gate90inter9));
  nand2 gate2153(.a(s_229), .b(gate90inter3), .O(gate90inter10));
  nor2  gate2154(.a(gate90inter10), .b(gate90inter9), .O(gate90inter11));
  nor2  gate2155(.a(gate90inter11), .b(gate90inter6), .O(gate90inter12));
  nand2 gate2156(.a(gate90inter12), .b(gate90inter1), .O(G411));
nand2 gate91( .a(G25), .b(G341), .O(G412) );

  xor2  gate883(.a(G341), .b(G29), .O(gate92inter0));
  nand2 gate884(.a(gate92inter0), .b(s_48), .O(gate92inter1));
  and2  gate885(.a(G341), .b(G29), .O(gate92inter2));
  inv1  gate886(.a(s_48), .O(gate92inter3));
  inv1  gate887(.a(s_49), .O(gate92inter4));
  nand2 gate888(.a(gate92inter4), .b(gate92inter3), .O(gate92inter5));
  nor2  gate889(.a(gate92inter5), .b(gate92inter2), .O(gate92inter6));
  inv1  gate890(.a(G29), .O(gate92inter7));
  inv1  gate891(.a(G341), .O(gate92inter8));
  nand2 gate892(.a(gate92inter8), .b(gate92inter7), .O(gate92inter9));
  nand2 gate893(.a(s_49), .b(gate92inter3), .O(gate92inter10));
  nor2  gate894(.a(gate92inter10), .b(gate92inter9), .O(gate92inter11));
  nor2  gate895(.a(gate92inter11), .b(gate92inter6), .O(gate92inter12));
  nand2 gate896(.a(gate92inter12), .b(gate92inter1), .O(G413));
nand2 gate93( .a(G18), .b(G344), .O(G414) );
nand2 gate94( .a(G22), .b(G344), .O(G415) );

  xor2  gate1345(.a(G347), .b(G26), .O(gate95inter0));
  nand2 gate1346(.a(gate95inter0), .b(s_114), .O(gate95inter1));
  and2  gate1347(.a(G347), .b(G26), .O(gate95inter2));
  inv1  gate1348(.a(s_114), .O(gate95inter3));
  inv1  gate1349(.a(s_115), .O(gate95inter4));
  nand2 gate1350(.a(gate95inter4), .b(gate95inter3), .O(gate95inter5));
  nor2  gate1351(.a(gate95inter5), .b(gate95inter2), .O(gate95inter6));
  inv1  gate1352(.a(G26), .O(gate95inter7));
  inv1  gate1353(.a(G347), .O(gate95inter8));
  nand2 gate1354(.a(gate95inter8), .b(gate95inter7), .O(gate95inter9));
  nand2 gate1355(.a(s_115), .b(gate95inter3), .O(gate95inter10));
  nor2  gate1356(.a(gate95inter10), .b(gate95inter9), .O(gate95inter11));
  nor2  gate1357(.a(gate95inter11), .b(gate95inter6), .O(gate95inter12));
  nand2 gate1358(.a(gate95inter12), .b(gate95inter1), .O(G416));
nand2 gate96( .a(G30), .b(G347), .O(G417) );
nand2 gate97( .a(G19), .b(G350), .O(G418) );
nand2 gate98( .a(G23), .b(G350), .O(G419) );
nand2 gate99( .a(G27), .b(G353), .O(G420) );

  xor2  gate547(.a(G353), .b(G31), .O(gate100inter0));
  nand2 gate548(.a(gate100inter0), .b(s_0), .O(gate100inter1));
  and2  gate549(.a(G353), .b(G31), .O(gate100inter2));
  inv1  gate550(.a(s_0), .O(gate100inter3));
  inv1  gate551(.a(s_1), .O(gate100inter4));
  nand2 gate552(.a(gate100inter4), .b(gate100inter3), .O(gate100inter5));
  nor2  gate553(.a(gate100inter5), .b(gate100inter2), .O(gate100inter6));
  inv1  gate554(.a(G31), .O(gate100inter7));
  inv1  gate555(.a(G353), .O(gate100inter8));
  nand2 gate556(.a(gate100inter8), .b(gate100inter7), .O(gate100inter9));
  nand2 gate557(.a(s_1), .b(gate100inter3), .O(gate100inter10));
  nor2  gate558(.a(gate100inter10), .b(gate100inter9), .O(gate100inter11));
  nor2  gate559(.a(gate100inter11), .b(gate100inter6), .O(gate100inter12));
  nand2 gate560(.a(gate100inter12), .b(gate100inter1), .O(G421));

  xor2  gate589(.a(G356), .b(G20), .O(gate101inter0));
  nand2 gate590(.a(gate101inter0), .b(s_6), .O(gate101inter1));
  and2  gate591(.a(G356), .b(G20), .O(gate101inter2));
  inv1  gate592(.a(s_6), .O(gate101inter3));
  inv1  gate593(.a(s_7), .O(gate101inter4));
  nand2 gate594(.a(gate101inter4), .b(gate101inter3), .O(gate101inter5));
  nor2  gate595(.a(gate101inter5), .b(gate101inter2), .O(gate101inter6));
  inv1  gate596(.a(G20), .O(gate101inter7));
  inv1  gate597(.a(G356), .O(gate101inter8));
  nand2 gate598(.a(gate101inter8), .b(gate101inter7), .O(gate101inter9));
  nand2 gate599(.a(s_7), .b(gate101inter3), .O(gate101inter10));
  nor2  gate600(.a(gate101inter10), .b(gate101inter9), .O(gate101inter11));
  nor2  gate601(.a(gate101inter11), .b(gate101inter6), .O(gate101inter12));
  nand2 gate602(.a(gate101inter12), .b(gate101inter1), .O(G422));

  xor2  gate1373(.a(G356), .b(G24), .O(gate102inter0));
  nand2 gate1374(.a(gate102inter0), .b(s_118), .O(gate102inter1));
  and2  gate1375(.a(G356), .b(G24), .O(gate102inter2));
  inv1  gate1376(.a(s_118), .O(gate102inter3));
  inv1  gate1377(.a(s_119), .O(gate102inter4));
  nand2 gate1378(.a(gate102inter4), .b(gate102inter3), .O(gate102inter5));
  nor2  gate1379(.a(gate102inter5), .b(gate102inter2), .O(gate102inter6));
  inv1  gate1380(.a(G24), .O(gate102inter7));
  inv1  gate1381(.a(G356), .O(gate102inter8));
  nand2 gate1382(.a(gate102inter8), .b(gate102inter7), .O(gate102inter9));
  nand2 gate1383(.a(s_119), .b(gate102inter3), .O(gate102inter10));
  nor2  gate1384(.a(gate102inter10), .b(gate102inter9), .O(gate102inter11));
  nor2  gate1385(.a(gate102inter11), .b(gate102inter6), .O(gate102inter12));
  nand2 gate1386(.a(gate102inter12), .b(gate102inter1), .O(G423));

  xor2  gate1863(.a(G359), .b(G28), .O(gate103inter0));
  nand2 gate1864(.a(gate103inter0), .b(s_188), .O(gate103inter1));
  and2  gate1865(.a(G359), .b(G28), .O(gate103inter2));
  inv1  gate1866(.a(s_188), .O(gate103inter3));
  inv1  gate1867(.a(s_189), .O(gate103inter4));
  nand2 gate1868(.a(gate103inter4), .b(gate103inter3), .O(gate103inter5));
  nor2  gate1869(.a(gate103inter5), .b(gate103inter2), .O(gate103inter6));
  inv1  gate1870(.a(G28), .O(gate103inter7));
  inv1  gate1871(.a(G359), .O(gate103inter8));
  nand2 gate1872(.a(gate103inter8), .b(gate103inter7), .O(gate103inter9));
  nand2 gate1873(.a(s_189), .b(gate103inter3), .O(gate103inter10));
  nor2  gate1874(.a(gate103inter10), .b(gate103inter9), .O(gate103inter11));
  nor2  gate1875(.a(gate103inter11), .b(gate103inter6), .O(gate103inter12));
  nand2 gate1876(.a(gate103inter12), .b(gate103inter1), .O(G424));
nand2 gate104( .a(G32), .b(G359), .O(G425) );
nand2 gate105( .a(G362), .b(G363), .O(G426) );
nand2 gate106( .a(G364), .b(G365), .O(G429) );

  xor2  gate995(.a(G367), .b(G366), .O(gate107inter0));
  nand2 gate996(.a(gate107inter0), .b(s_64), .O(gate107inter1));
  and2  gate997(.a(G367), .b(G366), .O(gate107inter2));
  inv1  gate998(.a(s_64), .O(gate107inter3));
  inv1  gate999(.a(s_65), .O(gate107inter4));
  nand2 gate1000(.a(gate107inter4), .b(gate107inter3), .O(gate107inter5));
  nor2  gate1001(.a(gate107inter5), .b(gate107inter2), .O(gate107inter6));
  inv1  gate1002(.a(G366), .O(gate107inter7));
  inv1  gate1003(.a(G367), .O(gate107inter8));
  nand2 gate1004(.a(gate107inter8), .b(gate107inter7), .O(gate107inter9));
  nand2 gate1005(.a(s_65), .b(gate107inter3), .O(gate107inter10));
  nor2  gate1006(.a(gate107inter10), .b(gate107inter9), .O(gate107inter11));
  nor2  gate1007(.a(gate107inter11), .b(gate107inter6), .O(gate107inter12));
  nand2 gate1008(.a(gate107inter12), .b(gate107inter1), .O(G432));
nand2 gate108( .a(G368), .b(G369), .O(G435) );
nand2 gate109( .a(G370), .b(G371), .O(G438) );
nand2 gate110( .a(G372), .b(G373), .O(G441) );
nand2 gate111( .a(G374), .b(G375), .O(G444) );

  xor2  gate1961(.a(G377), .b(G376), .O(gate112inter0));
  nand2 gate1962(.a(gate112inter0), .b(s_202), .O(gate112inter1));
  and2  gate1963(.a(G377), .b(G376), .O(gate112inter2));
  inv1  gate1964(.a(s_202), .O(gate112inter3));
  inv1  gate1965(.a(s_203), .O(gate112inter4));
  nand2 gate1966(.a(gate112inter4), .b(gate112inter3), .O(gate112inter5));
  nor2  gate1967(.a(gate112inter5), .b(gate112inter2), .O(gate112inter6));
  inv1  gate1968(.a(G376), .O(gate112inter7));
  inv1  gate1969(.a(G377), .O(gate112inter8));
  nand2 gate1970(.a(gate112inter8), .b(gate112inter7), .O(gate112inter9));
  nand2 gate1971(.a(s_203), .b(gate112inter3), .O(gate112inter10));
  nor2  gate1972(.a(gate112inter10), .b(gate112inter9), .O(gate112inter11));
  nor2  gate1973(.a(gate112inter11), .b(gate112inter6), .O(gate112inter12));
  nand2 gate1974(.a(gate112inter12), .b(gate112inter1), .O(G447));
nand2 gate113( .a(G378), .b(G379), .O(G450) );

  xor2  gate1037(.a(G381), .b(G380), .O(gate114inter0));
  nand2 gate1038(.a(gate114inter0), .b(s_70), .O(gate114inter1));
  and2  gate1039(.a(G381), .b(G380), .O(gate114inter2));
  inv1  gate1040(.a(s_70), .O(gate114inter3));
  inv1  gate1041(.a(s_71), .O(gate114inter4));
  nand2 gate1042(.a(gate114inter4), .b(gate114inter3), .O(gate114inter5));
  nor2  gate1043(.a(gate114inter5), .b(gate114inter2), .O(gate114inter6));
  inv1  gate1044(.a(G380), .O(gate114inter7));
  inv1  gate1045(.a(G381), .O(gate114inter8));
  nand2 gate1046(.a(gate114inter8), .b(gate114inter7), .O(gate114inter9));
  nand2 gate1047(.a(s_71), .b(gate114inter3), .O(gate114inter10));
  nor2  gate1048(.a(gate114inter10), .b(gate114inter9), .O(gate114inter11));
  nor2  gate1049(.a(gate114inter11), .b(gate114inter6), .O(gate114inter12));
  nand2 gate1050(.a(gate114inter12), .b(gate114inter1), .O(G453));
nand2 gate115( .a(G382), .b(G383), .O(G456) );
nand2 gate116( .a(G384), .b(G385), .O(G459) );

  xor2  gate981(.a(G387), .b(G386), .O(gate117inter0));
  nand2 gate982(.a(gate117inter0), .b(s_62), .O(gate117inter1));
  and2  gate983(.a(G387), .b(G386), .O(gate117inter2));
  inv1  gate984(.a(s_62), .O(gate117inter3));
  inv1  gate985(.a(s_63), .O(gate117inter4));
  nand2 gate986(.a(gate117inter4), .b(gate117inter3), .O(gate117inter5));
  nor2  gate987(.a(gate117inter5), .b(gate117inter2), .O(gate117inter6));
  inv1  gate988(.a(G386), .O(gate117inter7));
  inv1  gate989(.a(G387), .O(gate117inter8));
  nand2 gate990(.a(gate117inter8), .b(gate117inter7), .O(gate117inter9));
  nand2 gate991(.a(s_63), .b(gate117inter3), .O(gate117inter10));
  nor2  gate992(.a(gate117inter10), .b(gate117inter9), .O(gate117inter11));
  nor2  gate993(.a(gate117inter11), .b(gate117inter6), .O(gate117inter12));
  nand2 gate994(.a(gate117inter12), .b(gate117inter1), .O(G462));
nand2 gate118( .a(G388), .b(G389), .O(G465) );

  xor2  gate2423(.a(G391), .b(G390), .O(gate119inter0));
  nand2 gate2424(.a(gate119inter0), .b(s_268), .O(gate119inter1));
  and2  gate2425(.a(G391), .b(G390), .O(gate119inter2));
  inv1  gate2426(.a(s_268), .O(gate119inter3));
  inv1  gate2427(.a(s_269), .O(gate119inter4));
  nand2 gate2428(.a(gate119inter4), .b(gate119inter3), .O(gate119inter5));
  nor2  gate2429(.a(gate119inter5), .b(gate119inter2), .O(gate119inter6));
  inv1  gate2430(.a(G390), .O(gate119inter7));
  inv1  gate2431(.a(G391), .O(gate119inter8));
  nand2 gate2432(.a(gate119inter8), .b(gate119inter7), .O(gate119inter9));
  nand2 gate2433(.a(s_269), .b(gate119inter3), .O(gate119inter10));
  nor2  gate2434(.a(gate119inter10), .b(gate119inter9), .O(gate119inter11));
  nor2  gate2435(.a(gate119inter11), .b(gate119inter6), .O(gate119inter12));
  nand2 gate2436(.a(gate119inter12), .b(gate119inter1), .O(G468));
nand2 gate120( .a(G392), .b(G393), .O(G471) );
nand2 gate121( .a(G394), .b(G395), .O(G474) );
nand2 gate122( .a(G396), .b(G397), .O(G477) );
nand2 gate123( .a(G398), .b(G399), .O(G480) );
nand2 gate124( .a(G400), .b(G401), .O(G483) );
nand2 gate125( .a(G402), .b(G403), .O(G486) );

  xor2  gate2409(.a(G405), .b(G404), .O(gate126inter0));
  nand2 gate2410(.a(gate126inter0), .b(s_266), .O(gate126inter1));
  and2  gate2411(.a(G405), .b(G404), .O(gate126inter2));
  inv1  gate2412(.a(s_266), .O(gate126inter3));
  inv1  gate2413(.a(s_267), .O(gate126inter4));
  nand2 gate2414(.a(gate126inter4), .b(gate126inter3), .O(gate126inter5));
  nor2  gate2415(.a(gate126inter5), .b(gate126inter2), .O(gate126inter6));
  inv1  gate2416(.a(G404), .O(gate126inter7));
  inv1  gate2417(.a(G405), .O(gate126inter8));
  nand2 gate2418(.a(gate126inter8), .b(gate126inter7), .O(gate126inter9));
  nand2 gate2419(.a(s_267), .b(gate126inter3), .O(gate126inter10));
  nor2  gate2420(.a(gate126inter10), .b(gate126inter9), .O(gate126inter11));
  nor2  gate2421(.a(gate126inter11), .b(gate126inter6), .O(gate126inter12));
  nand2 gate2422(.a(gate126inter12), .b(gate126inter1), .O(G489));
nand2 gate127( .a(G406), .b(G407), .O(G492) );
nand2 gate128( .a(G408), .b(G409), .O(G495) );
nand2 gate129( .a(G410), .b(G411), .O(G498) );

  xor2  gate869(.a(G413), .b(G412), .O(gate130inter0));
  nand2 gate870(.a(gate130inter0), .b(s_46), .O(gate130inter1));
  and2  gate871(.a(G413), .b(G412), .O(gate130inter2));
  inv1  gate872(.a(s_46), .O(gate130inter3));
  inv1  gate873(.a(s_47), .O(gate130inter4));
  nand2 gate874(.a(gate130inter4), .b(gate130inter3), .O(gate130inter5));
  nor2  gate875(.a(gate130inter5), .b(gate130inter2), .O(gate130inter6));
  inv1  gate876(.a(G412), .O(gate130inter7));
  inv1  gate877(.a(G413), .O(gate130inter8));
  nand2 gate878(.a(gate130inter8), .b(gate130inter7), .O(gate130inter9));
  nand2 gate879(.a(s_47), .b(gate130inter3), .O(gate130inter10));
  nor2  gate880(.a(gate130inter10), .b(gate130inter9), .O(gate130inter11));
  nor2  gate881(.a(gate130inter11), .b(gate130inter6), .O(gate130inter12));
  nand2 gate882(.a(gate130inter12), .b(gate130inter1), .O(G501));

  xor2  gate2269(.a(G415), .b(G414), .O(gate131inter0));
  nand2 gate2270(.a(gate131inter0), .b(s_246), .O(gate131inter1));
  and2  gate2271(.a(G415), .b(G414), .O(gate131inter2));
  inv1  gate2272(.a(s_246), .O(gate131inter3));
  inv1  gate2273(.a(s_247), .O(gate131inter4));
  nand2 gate2274(.a(gate131inter4), .b(gate131inter3), .O(gate131inter5));
  nor2  gate2275(.a(gate131inter5), .b(gate131inter2), .O(gate131inter6));
  inv1  gate2276(.a(G414), .O(gate131inter7));
  inv1  gate2277(.a(G415), .O(gate131inter8));
  nand2 gate2278(.a(gate131inter8), .b(gate131inter7), .O(gate131inter9));
  nand2 gate2279(.a(s_247), .b(gate131inter3), .O(gate131inter10));
  nor2  gate2280(.a(gate131inter10), .b(gate131inter9), .O(gate131inter11));
  nor2  gate2281(.a(gate131inter11), .b(gate131inter6), .O(gate131inter12));
  nand2 gate2282(.a(gate131inter12), .b(gate131inter1), .O(G504));

  xor2  gate757(.a(G417), .b(G416), .O(gate132inter0));
  nand2 gate758(.a(gate132inter0), .b(s_30), .O(gate132inter1));
  and2  gate759(.a(G417), .b(G416), .O(gate132inter2));
  inv1  gate760(.a(s_30), .O(gate132inter3));
  inv1  gate761(.a(s_31), .O(gate132inter4));
  nand2 gate762(.a(gate132inter4), .b(gate132inter3), .O(gate132inter5));
  nor2  gate763(.a(gate132inter5), .b(gate132inter2), .O(gate132inter6));
  inv1  gate764(.a(G416), .O(gate132inter7));
  inv1  gate765(.a(G417), .O(gate132inter8));
  nand2 gate766(.a(gate132inter8), .b(gate132inter7), .O(gate132inter9));
  nand2 gate767(.a(s_31), .b(gate132inter3), .O(gate132inter10));
  nor2  gate768(.a(gate132inter10), .b(gate132inter9), .O(gate132inter11));
  nor2  gate769(.a(gate132inter11), .b(gate132inter6), .O(gate132inter12));
  nand2 gate770(.a(gate132inter12), .b(gate132inter1), .O(G507));

  xor2  gate1793(.a(G419), .b(G418), .O(gate133inter0));
  nand2 gate1794(.a(gate133inter0), .b(s_178), .O(gate133inter1));
  and2  gate1795(.a(G419), .b(G418), .O(gate133inter2));
  inv1  gate1796(.a(s_178), .O(gate133inter3));
  inv1  gate1797(.a(s_179), .O(gate133inter4));
  nand2 gate1798(.a(gate133inter4), .b(gate133inter3), .O(gate133inter5));
  nor2  gate1799(.a(gate133inter5), .b(gate133inter2), .O(gate133inter6));
  inv1  gate1800(.a(G418), .O(gate133inter7));
  inv1  gate1801(.a(G419), .O(gate133inter8));
  nand2 gate1802(.a(gate133inter8), .b(gate133inter7), .O(gate133inter9));
  nand2 gate1803(.a(s_179), .b(gate133inter3), .O(gate133inter10));
  nor2  gate1804(.a(gate133inter10), .b(gate133inter9), .O(gate133inter11));
  nor2  gate1805(.a(gate133inter11), .b(gate133inter6), .O(gate133inter12));
  nand2 gate1806(.a(gate133inter12), .b(gate133inter1), .O(G510));
nand2 gate134( .a(G420), .b(G421), .O(G513) );

  xor2  gate2031(.a(G423), .b(G422), .O(gate135inter0));
  nand2 gate2032(.a(gate135inter0), .b(s_212), .O(gate135inter1));
  and2  gate2033(.a(G423), .b(G422), .O(gate135inter2));
  inv1  gate2034(.a(s_212), .O(gate135inter3));
  inv1  gate2035(.a(s_213), .O(gate135inter4));
  nand2 gate2036(.a(gate135inter4), .b(gate135inter3), .O(gate135inter5));
  nor2  gate2037(.a(gate135inter5), .b(gate135inter2), .O(gate135inter6));
  inv1  gate2038(.a(G422), .O(gate135inter7));
  inv1  gate2039(.a(G423), .O(gate135inter8));
  nand2 gate2040(.a(gate135inter8), .b(gate135inter7), .O(gate135inter9));
  nand2 gate2041(.a(s_213), .b(gate135inter3), .O(gate135inter10));
  nor2  gate2042(.a(gate135inter10), .b(gate135inter9), .O(gate135inter11));
  nor2  gate2043(.a(gate135inter11), .b(gate135inter6), .O(gate135inter12));
  nand2 gate2044(.a(gate135inter12), .b(gate135inter1), .O(G516));
nand2 gate136( .a(G424), .b(G425), .O(G519) );

  xor2  gate1471(.a(G429), .b(G426), .O(gate137inter0));
  nand2 gate1472(.a(gate137inter0), .b(s_132), .O(gate137inter1));
  and2  gate1473(.a(G429), .b(G426), .O(gate137inter2));
  inv1  gate1474(.a(s_132), .O(gate137inter3));
  inv1  gate1475(.a(s_133), .O(gate137inter4));
  nand2 gate1476(.a(gate137inter4), .b(gate137inter3), .O(gate137inter5));
  nor2  gate1477(.a(gate137inter5), .b(gate137inter2), .O(gate137inter6));
  inv1  gate1478(.a(G426), .O(gate137inter7));
  inv1  gate1479(.a(G429), .O(gate137inter8));
  nand2 gate1480(.a(gate137inter8), .b(gate137inter7), .O(gate137inter9));
  nand2 gate1481(.a(s_133), .b(gate137inter3), .O(gate137inter10));
  nor2  gate1482(.a(gate137inter10), .b(gate137inter9), .O(gate137inter11));
  nor2  gate1483(.a(gate137inter11), .b(gate137inter6), .O(gate137inter12));
  nand2 gate1484(.a(gate137inter12), .b(gate137inter1), .O(G522));
nand2 gate138( .a(G432), .b(G435), .O(G525) );
nand2 gate139( .a(G438), .b(G441), .O(G528) );
nand2 gate140( .a(G444), .b(G447), .O(G531) );
nand2 gate141( .a(G450), .b(G453), .O(G534) );
nand2 gate142( .a(G456), .b(G459), .O(G537) );

  xor2  gate2311(.a(G465), .b(G462), .O(gate143inter0));
  nand2 gate2312(.a(gate143inter0), .b(s_252), .O(gate143inter1));
  and2  gate2313(.a(G465), .b(G462), .O(gate143inter2));
  inv1  gate2314(.a(s_252), .O(gate143inter3));
  inv1  gate2315(.a(s_253), .O(gate143inter4));
  nand2 gate2316(.a(gate143inter4), .b(gate143inter3), .O(gate143inter5));
  nor2  gate2317(.a(gate143inter5), .b(gate143inter2), .O(gate143inter6));
  inv1  gate2318(.a(G462), .O(gate143inter7));
  inv1  gate2319(.a(G465), .O(gate143inter8));
  nand2 gate2320(.a(gate143inter8), .b(gate143inter7), .O(gate143inter9));
  nand2 gate2321(.a(s_253), .b(gate143inter3), .O(gate143inter10));
  nor2  gate2322(.a(gate143inter10), .b(gate143inter9), .O(gate143inter11));
  nor2  gate2323(.a(gate143inter11), .b(gate143inter6), .O(gate143inter12));
  nand2 gate2324(.a(gate143inter12), .b(gate143inter1), .O(G540));
nand2 gate144( .a(G468), .b(G471), .O(G543) );
nand2 gate145( .a(G474), .b(G477), .O(G546) );
nand2 gate146( .a(G480), .b(G483), .O(G549) );

  xor2  gate1457(.a(G489), .b(G486), .O(gate147inter0));
  nand2 gate1458(.a(gate147inter0), .b(s_130), .O(gate147inter1));
  and2  gate1459(.a(G489), .b(G486), .O(gate147inter2));
  inv1  gate1460(.a(s_130), .O(gate147inter3));
  inv1  gate1461(.a(s_131), .O(gate147inter4));
  nand2 gate1462(.a(gate147inter4), .b(gate147inter3), .O(gate147inter5));
  nor2  gate1463(.a(gate147inter5), .b(gate147inter2), .O(gate147inter6));
  inv1  gate1464(.a(G486), .O(gate147inter7));
  inv1  gate1465(.a(G489), .O(gate147inter8));
  nand2 gate1466(.a(gate147inter8), .b(gate147inter7), .O(gate147inter9));
  nand2 gate1467(.a(s_131), .b(gate147inter3), .O(gate147inter10));
  nor2  gate1468(.a(gate147inter10), .b(gate147inter9), .O(gate147inter11));
  nor2  gate1469(.a(gate147inter11), .b(gate147inter6), .O(gate147inter12));
  nand2 gate1470(.a(gate147inter12), .b(gate147inter1), .O(G552));
nand2 gate148( .a(G492), .b(G495), .O(G555) );
nand2 gate149( .a(G498), .b(G501), .O(G558) );
nand2 gate150( .a(G504), .b(G507), .O(G561) );
nand2 gate151( .a(G510), .b(G513), .O(G564) );

  xor2  gate1219(.a(G519), .b(G516), .O(gate152inter0));
  nand2 gate1220(.a(gate152inter0), .b(s_96), .O(gate152inter1));
  and2  gate1221(.a(G519), .b(G516), .O(gate152inter2));
  inv1  gate1222(.a(s_96), .O(gate152inter3));
  inv1  gate1223(.a(s_97), .O(gate152inter4));
  nand2 gate1224(.a(gate152inter4), .b(gate152inter3), .O(gate152inter5));
  nor2  gate1225(.a(gate152inter5), .b(gate152inter2), .O(gate152inter6));
  inv1  gate1226(.a(G516), .O(gate152inter7));
  inv1  gate1227(.a(G519), .O(gate152inter8));
  nand2 gate1228(.a(gate152inter8), .b(gate152inter7), .O(gate152inter9));
  nand2 gate1229(.a(s_97), .b(gate152inter3), .O(gate152inter10));
  nor2  gate1230(.a(gate152inter10), .b(gate152inter9), .O(gate152inter11));
  nor2  gate1231(.a(gate152inter11), .b(gate152inter6), .O(gate152inter12));
  nand2 gate1232(.a(gate152inter12), .b(gate152inter1), .O(G567));

  xor2  gate743(.a(G522), .b(G426), .O(gate153inter0));
  nand2 gate744(.a(gate153inter0), .b(s_28), .O(gate153inter1));
  and2  gate745(.a(G522), .b(G426), .O(gate153inter2));
  inv1  gate746(.a(s_28), .O(gate153inter3));
  inv1  gate747(.a(s_29), .O(gate153inter4));
  nand2 gate748(.a(gate153inter4), .b(gate153inter3), .O(gate153inter5));
  nor2  gate749(.a(gate153inter5), .b(gate153inter2), .O(gate153inter6));
  inv1  gate750(.a(G426), .O(gate153inter7));
  inv1  gate751(.a(G522), .O(gate153inter8));
  nand2 gate752(.a(gate153inter8), .b(gate153inter7), .O(gate153inter9));
  nand2 gate753(.a(s_29), .b(gate153inter3), .O(gate153inter10));
  nor2  gate754(.a(gate153inter10), .b(gate153inter9), .O(gate153inter11));
  nor2  gate755(.a(gate153inter11), .b(gate153inter6), .O(gate153inter12));
  nand2 gate756(.a(gate153inter12), .b(gate153inter1), .O(G570));

  xor2  gate729(.a(G522), .b(G429), .O(gate154inter0));
  nand2 gate730(.a(gate154inter0), .b(s_26), .O(gate154inter1));
  and2  gate731(.a(G522), .b(G429), .O(gate154inter2));
  inv1  gate732(.a(s_26), .O(gate154inter3));
  inv1  gate733(.a(s_27), .O(gate154inter4));
  nand2 gate734(.a(gate154inter4), .b(gate154inter3), .O(gate154inter5));
  nor2  gate735(.a(gate154inter5), .b(gate154inter2), .O(gate154inter6));
  inv1  gate736(.a(G429), .O(gate154inter7));
  inv1  gate737(.a(G522), .O(gate154inter8));
  nand2 gate738(.a(gate154inter8), .b(gate154inter7), .O(gate154inter9));
  nand2 gate739(.a(s_27), .b(gate154inter3), .O(gate154inter10));
  nor2  gate740(.a(gate154inter10), .b(gate154inter9), .O(gate154inter11));
  nor2  gate741(.a(gate154inter11), .b(gate154inter6), .O(gate154inter12));
  nand2 gate742(.a(gate154inter12), .b(gate154inter1), .O(G571));
nand2 gate155( .a(G432), .b(G525), .O(G572) );
nand2 gate156( .a(G435), .b(G525), .O(G573) );
nand2 gate157( .a(G438), .b(G528), .O(G574) );
nand2 gate158( .a(G441), .b(G528), .O(G575) );
nand2 gate159( .a(G444), .b(G531), .O(G576) );

  xor2  gate1065(.a(G531), .b(G447), .O(gate160inter0));
  nand2 gate1066(.a(gate160inter0), .b(s_74), .O(gate160inter1));
  and2  gate1067(.a(G531), .b(G447), .O(gate160inter2));
  inv1  gate1068(.a(s_74), .O(gate160inter3));
  inv1  gate1069(.a(s_75), .O(gate160inter4));
  nand2 gate1070(.a(gate160inter4), .b(gate160inter3), .O(gate160inter5));
  nor2  gate1071(.a(gate160inter5), .b(gate160inter2), .O(gate160inter6));
  inv1  gate1072(.a(G447), .O(gate160inter7));
  inv1  gate1073(.a(G531), .O(gate160inter8));
  nand2 gate1074(.a(gate160inter8), .b(gate160inter7), .O(gate160inter9));
  nand2 gate1075(.a(s_75), .b(gate160inter3), .O(gate160inter10));
  nor2  gate1076(.a(gate160inter10), .b(gate160inter9), .O(gate160inter11));
  nor2  gate1077(.a(gate160inter11), .b(gate160inter6), .O(gate160inter12));
  nand2 gate1078(.a(gate160inter12), .b(gate160inter1), .O(G577));

  xor2  gate2101(.a(G534), .b(G450), .O(gate161inter0));
  nand2 gate2102(.a(gate161inter0), .b(s_222), .O(gate161inter1));
  and2  gate2103(.a(G534), .b(G450), .O(gate161inter2));
  inv1  gate2104(.a(s_222), .O(gate161inter3));
  inv1  gate2105(.a(s_223), .O(gate161inter4));
  nand2 gate2106(.a(gate161inter4), .b(gate161inter3), .O(gate161inter5));
  nor2  gate2107(.a(gate161inter5), .b(gate161inter2), .O(gate161inter6));
  inv1  gate2108(.a(G450), .O(gate161inter7));
  inv1  gate2109(.a(G534), .O(gate161inter8));
  nand2 gate2110(.a(gate161inter8), .b(gate161inter7), .O(gate161inter9));
  nand2 gate2111(.a(s_223), .b(gate161inter3), .O(gate161inter10));
  nor2  gate2112(.a(gate161inter10), .b(gate161inter9), .O(gate161inter11));
  nor2  gate2113(.a(gate161inter11), .b(gate161inter6), .O(gate161inter12));
  nand2 gate2114(.a(gate161inter12), .b(gate161inter1), .O(G578));

  xor2  gate1121(.a(G534), .b(G453), .O(gate162inter0));
  nand2 gate1122(.a(gate162inter0), .b(s_82), .O(gate162inter1));
  and2  gate1123(.a(G534), .b(G453), .O(gate162inter2));
  inv1  gate1124(.a(s_82), .O(gate162inter3));
  inv1  gate1125(.a(s_83), .O(gate162inter4));
  nand2 gate1126(.a(gate162inter4), .b(gate162inter3), .O(gate162inter5));
  nor2  gate1127(.a(gate162inter5), .b(gate162inter2), .O(gate162inter6));
  inv1  gate1128(.a(G453), .O(gate162inter7));
  inv1  gate1129(.a(G534), .O(gate162inter8));
  nand2 gate1130(.a(gate162inter8), .b(gate162inter7), .O(gate162inter9));
  nand2 gate1131(.a(s_83), .b(gate162inter3), .O(gate162inter10));
  nor2  gate1132(.a(gate162inter10), .b(gate162inter9), .O(gate162inter11));
  nor2  gate1133(.a(gate162inter11), .b(gate162inter6), .O(gate162inter12));
  nand2 gate1134(.a(gate162inter12), .b(gate162inter1), .O(G579));

  xor2  gate1009(.a(G537), .b(G456), .O(gate163inter0));
  nand2 gate1010(.a(gate163inter0), .b(s_66), .O(gate163inter1));
  and2  gate1011(.a(G537), .b(G456), .O(gate163inter2));
  inv1  gate1012(.a(s_66), .O(gate163inter3));
  inv1  gate1013(.a(s_67), .O(gate163inter4));
  nand2 gate1014(.a(gate163inter4), .b(gate163inter3), .O(gate163inter5));
  nor2  gate1015(.a(gate163inter5), .b(gate163inter2), .O(gate163inter6));
  inv1  gate1016(.a(G456), .O(gate163inter7));
  inv1  gate1017(.a(G537), .O(gate163inter8));
  nand2 gate1018(.a(gate163inter8), .b(gate163inter7), .O(gate163inter9));
  nand2 gate1019(.a(s_67), .b(gate163inter3), .O(gate163inter10));
  nor2  gate1020(.a(gate163inter10), .b(gate163inter9), .O(gate163inter11));
  nor2  gate1021(.a(gate163inter11), .b(gate163inter6), .O(gate163inter12));
  nand2 gate1022(.a(gate163inter12), .b(gate163inter1), .O(G580));
nand2 gate164( .a(G459), .b(G537), .O(G581) );

  xor2  gate1415(.a(G540), .b(G462), .O(gate165inter0));
  nand2 gate1416(.a(gate165inter0), .b(s_124), .O(gate165inter1));
  and2  gate1417(.a(G540), .b(G462), .O(gate165inter2));
  inv1  gate1418(.a(s_124), .O(gate165inter3));
  inv1  gate1419(.a(s_125), .O(gate165inter4));
  nand2 gate1420(.a(gate165inter4), .b(gate165inter3), .O(gate165inter5));
  nor2  gate1421(.a(gate165inter5), .b(gate165inter2), .O(gate165inter6));
  inv1  gate1422(.a(G462), .O(gate165inter7));
  inv1  gate1423(.a(G540), .O(gate165inter8));
  nand2 gate1424(.a(gate165inter8), .b(gate165inter7), .O(gate165inter9));
  nand2 gate1425(.a(s_125), .b(gate165inter3), .O(gate165inter10));
  nor2  gate1426(.a(gate165inter10), .b(gate165inter9), .O(gate165inter11));
  nor2  gate1427(.a(gate165inter11), .b(gate165inter6), .O(gate165inter12));
  nand2 gate1428(.a(gate165inter12), .b(gate165inter1), .O(G582));

  xor2  gate1247(.a(G540), .b(G465), .O(gate166inter0));
  nand2 gate1248(.a(gate166inter0), .b(s_100), .O(gate166inter1));
  and2  gate1249(.a(G540), .b(G465), .O(gate166inter2));
  inv1  gate1250(.a(s_100), .O(gate166inter3));
  inv1  gate1251(.a(s_101), .O(gate166inter4));
  nand2 gate1252(.a(gate166inter4), .b(gate166inter3), .O(gate166inter5));
  nor2  gate1253(.a(gate166inter5), .b(gate166inter2), .O(gate166inter6));
  inv1  gate1254(.a(G465), .O(gate166inter7));
  inv1  gate1255(.a(G540), .O(gate166inter8));
  nand2 gate1256(.a(gate166inter8), .b(gate166inter7), .O(gate166inter9));
  nand2 gate1257(.a(s_101), .b(gate166inter3), .O(gate166inter10));
  nor2  gate1258(.a(gate166inter10), .b(gate166inter9), .O(gate166inter11));
  nor2  gate1259(.a(gate166inter11), .b(gate166inter6), .O(gate166inter12));
  nand2 gate1260(.a(gate166inter12), .b(gate166inter1), .O(G583));
nand2 gate167( .a(G468), .b(G543), .O(G584) );
nand2 gate168( .a(G471), .b(G543), .O(G585) );
nand2 gate169( .a(G474), .b(G546), .O(G586) );
nand2 gate170( .a(G477), .b(G546), .O(G587) );
nand2 gate171( .a(G480), .b(G549), .O(G588) );
nand2 gate172( .a(G483), .b(G549), .O(G589) );
nand2 gate173( .a(G486), .b(G552), .O(G590) );

  xor2  gate1877(.a(G552), .b(G489), .O(gate174inter0));
  nand2 gate1878(.a(gate174inter0), .b(s_190), .O(gate174inter1));
  and2  gate1879(.a(G552), .b(G489), .O(gate174inter2));
  inv1  gate1880(.a(s_190), .O(gate174inter3));
  inv1  gate1881(.a(s_191), .O(gate174inter4));
  nand2 gate1882(.a(gate174inter4), .b(gate174inter3), .O(gate174inter5));
  nor2  gate1883(.a(gate174inter5), .b(gate174inter2), .O(gate174inter6));
  inv1  gate1884(.a(G489), .O(gate174inter7));
  inv1  gate1885(.a(G552), .O(gate174inter8));
  nand2 gate1886(.a(gate174inter8), .b(gate174inter7), .O(gate174inter9));
  nand2 gate1887(.a(s_191), .b(gate174inter3), .O(gate174inter10));
  nor2  gate1888(.a(gate174inter10), .b(gate174inter9), .O(gate174inter11));
  nor2  gate1889(.a(gate174inter11), .b(gate174inter6), .O(gate174inter12));
  nand2 gate1890(.a(gate174inter12), .b(gate174inter1), .O(G591));

  xor2  gate1625(.a(G555), .b(G492), .O(gate175inter0));
  nand2 gate1626(.a(gate175inter0), .b(s_154), .O(gate175inter1));
  and2  gate1627(.a(G555), .b(G492), .O(gate175inter2));
  inv1  gate1628(.a(s_154), .O(gate175inter3));
  inv1  gate1629(.a(s_155), .O(gate175inter4));
  nand2 gate1630(.a(gate175inter4), .b(gate175inter3), .O(gate175inter5));
  nor2  gate1631(.a(gate175inter5), .b(gate175inter2), .O(gate175inter6));
  inv1  gate1632(.a(G492), .O(gate175inter7));
  inv1  gate1633(.a(G555), .O(gate175inter8));
  nand2 gate1634(.a(gate175inter8), .b(gate175inter7), .O(gate175inter9));
  nand2 gate1635(.a(s_155), .b(gate175inter3), .O(gate175inter10));
  nor2  gate1636(.a(gate175inter10), .b(gate175inter9), .O(gate175inter11));
  nor2  gate1637(.a(gate175inter11), .b(gate175inter6), .O(gate175inter12));
  nand2 gate1638(.a(gate175inter12), .b(gate175inter1), .O(G592));

  xor2  gate1149(.a(G555), .b(G495), .O(gate176inter0));
  nand2 gate1150(.a(gate176inter0), .b(s_86), .O(gate176inter1));
  and2  gate1151(.a(G555), .b(G495), .O(gate176inter2));
  inv1  gate1152(.a(s_86), .O(gate176inter3));
  inv1  gate1153(.a(s_87), .O(gate176inter4));
  nand2 gate1154(.a(gate176inter4), .b(gate176inter3), .O(gate176inter5));
  nor2  gate1155(.a(gate176inter5), .b(gate176inter2), .O(gate176inter6));
  inv1  gate1156(.a(G495), .O(gate176inter7));
  inv1  gate1157(.a(G555), .O(gate176inter8));
  nand2 gate1158(.a(gate176inter8), .b(gate176inter7), .O(gate176inter9));
  nand2 gate1159(.a(s_87), .b(gate176inter3), .O(gate176inter10));
  nor2  gate1160(.a(gate176inter10), .b(gate176inter9), .O(gate176inter11));
  nor2  gate1161(.a(gate176inter11), .b(gate176inter6), .O(gate176inter12));
  nand2 gate1162(.a(gate176inter12), .b(gate176inter1), .O(G593));

  xor2  gate561(.a(G558), .b(G498), .O(gate177inter0));
  nand2 gate562(.a(gate177inter0), .b(s_2), .O(gate177inter1));
  and2  gate563(.a(G558), .b(G498), .O(gate177inter2));
  inv1  gate564(.a(s_2), .O(gate177inter3));
  inv1  gate565(.a(s_3), .O(gate177inter4));
  nand2 gate566(.a(gate177inter4), .b(gate177inter3), .O(gate177inter5));
  nor2  gate567(.a(gate177inter5), .b(gate177inter2), .O(gate177inter6));
  inv1  gate568(.a(G498), .O(gate177inter7));
  inv1  gate569(.a(G558), .O(gate177inter8));
  nand2 gate570(.a(gate177inter8), .b(gate177inter7), .O(gate177inter9));
  nand2 gate571(.a(s_3), .b(gate177inter3), .O(gate177inter10));
  nor2  gate572(.a(gate177inter10), .b(gate177inter9), .O(gate177inter11));
  nor2  gate573(.a(gate177inter11), .b(gate177inter6), .O(gate177inter12));
  nand2 gate574(.a(gate177inter12), .b(gate177inter1), .O(G594));
nand2 gate178( .a(G501), .b(G558), .O(G595) );
nand2 gate179( .a(G504), .b(G561), .O(G596) );
nand2 gate180( .a(G507), .b(G561), .O(G597) );
nand2 gate181( .a(G510), .b(G564), .O(G598) );
nand2 gate182( .a(G513), .b(G564), .O(G599) );

  xor2  gate1485(.a(G567), .b(G516), .O(gate183inter0));
  nand2 gate1486(.a(gate183inter0), .b(s_134), .O(gate183inter1));
  and2  gate1487(.a(G567), .b(G516), .O(gate183inter2));
  inv1  gate1488(.a(s_134), .O(gate183inter3));
  inv1  gate1489(.a(s_135), .O(gate183inter4));
  nand2 gate1490(.a(gate183inter4), .b(gate183inter3), .O(gate183inter5));
  nor2  gate1491(.a(gate183inter5), .b(gate183inter2), .O(gate183inter6));
  inv1  gate1492(.a(G516), .O(gate183inter7));
  inv1  gate1493(.a(G567), .O(gate183inter8));
  nand2 gate1494(.a(gate183inter8), .b(gate183inter7), .O(gate183inter9));
  nand2 gate1495(.a(s_135), .b(gate183inter3), .O(gate183inter10));
  nor2  gate1496(.a(gate183inter10), .b(gate183inter9), .O(gate183inter11));
  nor2  gate1497(.a(gate183inter11), .b(gate183inter6), .O(gate183inter12));
  nand2 gate1498(.a(gate183inter12), .b(gate183inter1), .O(G600));
nand2 gate184( .a(G519), .b(G567), .O(G601) );
nand2 gate185( .a(G570), .b(G571), .O(G602) );

  xor2  gate1023(.a(G573), .b(G572), .O(gate186inter0));
  nand2 gate1024(.a(gate186inter0), .b(s_68), .O(gate186inter1));
  and2  gate1025(.a(G573), .b(G572), .O(gate186inter2));
  inv1  gate1026(.a(s_68), .O(gate186inter3));
  inv1  gate1027(.a(s_69), .O(gate186inter4));
  nand2 gate1028(.a(gate186inter4), .b(gate186inter3), .O(gate186inter5));
  nor2  gate1029(.a(gate186inter5), .b(gate186inter2), .O(gate186inter6));
  inv1  gate1030(.a(G572), .O(gate186inter7));
  inv1  gate1031(.a(G573), .O(gate186inter8));
  nand2 gate1032(.a(gate186inter8), .b(gate186inter7), .O(gate186inter9));
  nand2 gate1033(.a(s_69), .b(gate186inter3), .O(gate186inter10));
  nor2  gate1034(.a(gate186inter10), .b(gate186inter9), .O(gate186inter11));
  nor2  gate1035(.a(gate186inter11), .b(gate186inter6), .O(gate186inter12));
  nand2 gate1036(.a(gate186inter12), .b(gate186inter1), .O(G607));
nand2 gate187( .a(G574), .b(G575), .O(G612) );
nand2 gate188( .a(G576), .b(G577), .O(G617) );
nand2 gate189( .a(G578), .b(G579), .O(G622) );

  xor2  gate2227(.a(G581), .b(G580), .O(gate190inter0));
  nand2 gate2228(.a(gate190inter0), .b(s_240), .O(gate190inter1));
  and2  gate2229(.a(G581), .b(G580), .O(gate190inter2));
  inv1  gate2230(.a(s_240), .O(gate190inter3));
  inv1  gate2231(.a(s_241), .O(gate190inter4));
  nand2 gate2232(.a(gate190inter4), .b(gate190inter3), .O(gate190inter5));
  nor2  gate2233(.a(gate190inter5), .b(gate190inter2), .O(gate190inter6));
  inv1  gate2234(.a(G580), .O(gate190inter7));
  inv1  gate2235(.a(G581), .O(gate190inter8));
  nand2 gate2236(.a(gate190inter8), .b(gate190inter7), .O(gate190inter9));
  nand2 gate2237(.a(s_241), .b(gate190inter3), .O(gate190inter10));
  nor2  gate2238(.a(gate190inter10), .b(gate190inter9), .O(gate190inter11));
  nor2  gate2239(.a(gate190inter11), .b(gate190inter6), .O(gate190inter12));
  nand2 gate2240(.a(gate190inter12), .b(gate190inter1), .O(G627));
nand2 gate191( .a(G582), .b(G583), .O(G632) );
nand2 gate192( .a(G584), .b(G585), .O(G637) );

  xor2  gate2493(.a(G587), .b(G586), .O(gate193inter0));
  nand2 gate2494(.a(gate193inter0), .b(s_278), .O(gate193inter1));
  and2  gate2495(.a(G587), .b(G586), .O(gate193inter2));
  inv1  gate2496(.a(s_278), .O(gate193inter3));
  inv1  gate2497(.a(s_279), .O(gate193inter4));
  nand2 gate2498(.a(gate193inter4), .b(gate193inter3), .O(gate193inter5));
  nor2  gate2499(.a(gate193inter5), .b(gate193inter2), .O(gate193inter6));
  inv1  gate2500(.a(G586), .O(gate193inter7));
  inv1  gate2501(.a(G587), .O(gate193inter8));
  nand2 gate2502(.a(gate193inter8), .b(gate193inter7), .O(gate193inter9));
  nand2 gate2503(.a(s_279), .b(gate193inter3), .O(gate193inter10));
  nor2  gate2504(.a(gate193inter10), .b(gate193inter9), .O(gate193inter11));
  nor2  gate2505(.a(gate193inter11), .b(gate193inter6), .O(gate193inter12));
  nand2 gate2506(.a(gate193inter12), .b(gate193inter1), .O(G642));
nand2 gate194( .a(G588), .b(G589), .O(G645) );

  xor2  gate2605(.a(G591), .b(G590), .O(gate195inter0));
  nand2 gate2606(.a(gate195inter0), .b(s_294), .O(gate195inter1));
  and2  gate2607(.a(G591), .b(G590), .O(gate195inter2));
  inv1  gate2608(.a(s_294), .O(gate195inter3));
  inv1  gate2609(.a(s_295), .O(gate195inter4));
  nand2 gate2610(.a(gate195inter4), .b(gate195inter3), .O(gate195inter5));
  nor2  gate2611(.a(gate195inter5), .b(gate195inter2), .O(gate195inter6));
  inv1  gate2612(.a(G590), .O(gate195inter7));
  inv1  gate2613(.a(G591), .O(gate195inter8));
  nand2 gate2614(.a(gate195inter8), .b(gate195inter7), .O(gate195inter9));
  nand2 gate2615(.a(s_295), .b(gate195inter3), .O(gate195inter10));
  nor2  gate2616(.a(gate195inter10), .b(gate195inter9), .O(gate195inter11));
  nor2  gate2617(.a(gate195inter11), .b(gate195inter6), .O(gate195inter12));
  nand2 gate2618(.a(gate195inter12), .b(gate195inter1), .O(G648));
nand2 gate196( .a(G592), .b(G593), .O(G651) );

  xor2  gate771(.a(G595), .b(G594), .O(gate197inter0));
  nand2 gate772(.a(gate197inter0), .b(s_32), .O(gate197inter1));
  and2  gate773(.a(G595), .b(G594), .O(gate197inter2));
  inv1  gate774(.a(s_32), .O(gate197inter3));
  inv1  gate775(.a(s_33), .O(gate197inter4));
  nand2 gate776(.a(gate197inter4), .b(gate197inter3), .O(gate197inter5));
  nor2  gate777(.a(gate197inter5), .b(gate197inter2), .O(gate197inter6));
  inv1  gate778(.a(G594), .O(gate197inter7));
  inv1  gate779(.a(G595), .O(gate197inter8));
  nand2 gate780(.a(gate197inter8), .b(gate197inter7), .O(gate197inter9));
  nand2 gate781(.a(s_33), .b(gate197inter3), .O(gate197inter10));
  nor2  gate782(.a(gate197inter10), .b(gate197inter9), .O(gate197inter11));
  nor2  gate783(.a(gate197inter11), .b(gate197inter6), .O(gate197inter12));
  nand2 gate784(.a(gate197inter12), .b(gate197inter1), .O(G654));
nand2 gate198( .a(G596), .b(G597), .O(G657) );

  xor2  gate603(.a(G599), .b(G598), .O(gate199inter0));
  nand2 gate604(.a(gate199inter0), .b(s_8), .O(gate199inter1));
  and2  gate605(.a(G599), .b(G598), .O(gate199inter2));
  inv1  gate606(.a(s_8), .O(gate199inter3));
  inv1  gate607(.a(s_9), .O(gate199inter4));
  nand2 gate608(.a(gate199inter4), .b(gate199inter3), .O(gate199inter5));
  nor2  gate609(.a(gate199inter5), .b(gate199inter2), .O(gate199inter6));
  inv1  gate610(.a(G598), .O(gate199inter7));
  inv1  gate611(.a(G599), .O(gate199inter8));
  nand2 gate612(.a(gate199inter8), .b(gate199inter7), .O(gate199inter9));
  nand2 gate613(.a(s_9), .b(gate199inter3), .O(gate199inter10));
  nor2  gate614(.a(gate199inter10), .b(gate199inter9), .O(gate199inter11));
  nor2  gate615(.a(gate199inter11), .b(gate199inter6), .O(gate199inter12));
  nand2 gate616(.a(gate199inter12), .b(gate199inter1), .O(G660));
nand2 gate200( .a(G600), .b(G601), .O(G663) );

  xor2  gate1191(.a(G607), .b(G602), .O(gate201inter0));
  nand2 gate1192(.a(gate201inter0), .b(s_92), .O(gate201inter1));
  and2  gate1193(.a(G607), .b(G602), .O(gate201inter2));
  inv1  gate1194(.a(s_92), .O(gate201inter3));
  inv1  gate1195(.a(s_93), .O(gate201inter4));
  nand2 gate1196(.a(gate201inter4), .b(gate201inter3), .O(gate201inter5));
  nor2  gate1197(.a(gate201inter5), .b(gate201inter2), .O(gate201inter6));
  inv1  gate1198(.a(G602), .O(gate201inter7));
  inv1  gate1199(.a(G607), .O(gate201inter8));
  nand2 gate1200(.a(gate201inter8), .b(gate201inter7), .O(gate201inter9));
  nand2 gate1201(.a(s_93), .b(gate201inter3), .O(gate201inter10));
  nor2  gate1202(.a(gate201inter10), .b(gate201inter9), .O(gate201inter11));
  nor2  gate1203(.a(gate201inter11), .b(gate201inter6), .O(gate201inter12));
  nand2 gate1204(.a(gate201inter12), .b(gate201inter1), .O(G666));
nand2 gate202( .a(G612), .b(G617), .O(G669) );
nand2 gate203( .a(G602), .b(G612), .O(G672) );
nand2 gate204( .a(G607), .b(G617), .O(G675) );
nand2 gate205( .a(G622), .b(G627), .O(G678) );

  xor2  gate2451(.a(G637), .b(G632), .O(gate206inter0));
  nand2 gate2452(.a(gate206inter0), .b(s_272), .O(gate206inter1));
  and2  gate2453(.a(G637), .b(G632), .O(gate206inter2));
  inv1  gate2454(.a(s_272), .O(gate206inter3));
  inv1  gate2455(.a(s_273), .O(gate206inter4));
  nand2 gate2456(.a(gate206inter4), .b(gate206inter3), .O(gate206inter5));
  nor2  gate2457(.a(gate206inter5), .b(gate206inter2), .O(gate206inter6));
  inv1  gate2458(.a(G632), .O(gate206inter7));
  inv1  gate2459(.a(G637), .O(gate206inter8));
  nand2 gate2460(.a(gate206inter8), .b(gate206inter7), .O(gate206inter9));
  nand2 gate2461(.a(s_273), .b(gate206inter3), .O(gate206inter10));
  nor2  gate2462(.a(gate206inter10), .b(gate206inter9), .O(gate206inter11));
  nor2  gate2463(.a(gate206inter11), .b(gate206inter6), .O(gate206inter12));
  nand2 gate2464(.a(gate206inter12), .b(gate206inter1), .O(G681));

  xor2  gate2241(.a(G632), .b(G622), .O(gate207inter0));
  nand2 gate2242(.a(gate207inter0), .b(s_242), .O(gate207inter1));
  and2  gate2243(.a(G632), .b(G622), .O(gate207inter2));
  inv1  gate2244(.a(s_242), .O(gate207inter3));
  inv1  gate2245(.a(s_243), .O(gate207inter4));
  nand2 gate2246(.a(gate207inter4), .b(gate207inter3), .O(gate207inter5));
  nor2  gate2247(.a(gate207inter5), .b(gate207inter2), .O(gate207inter6));
  inv1  gate2248(.a(G622), .O(gate207inter7));
  inv1  gate2249(.a(G632), .O(gate207inter8));
  nand2 gate2250(.a(gate207inter8), .b(gate207inter7), .O(gate207inter9));
  nand2 gate2251(.a(s_243), .b(gate207inter3), .O(gate207inter10));
  nor2  gate2252(.a(gate207inter10), .b(gate207inter9), .O(gate207inter11));
  nor2  gate2253(.a(gate207inter11), .b(gate207inter6), .O(gate207inter12));
  nand2 gate2254(.a(gate207inter12), .b(gate207inter1), .O(G684));
nand2 gate208( .a(G627), .b(G637), .O(G687) );
nand2 gate209( .a(G602), .b(G666), .O(G690) );
nand2 gate210( .a(G607), .b(G666), .O(G691) );
nand2 gate211( .a(G612), .b(G669), .O(G692) );
nand2 gate212( .a(G617), .b(G669), .O(G693) );
nand2 gate213( .a(G602), .b(G672), .O(G694) );
nand2 gate214( .a(G612), .b(G672), .O(G695) );
nand2 gate215( .a(G607), .b(G675), .O(G696) );
nand2 gate216( .a(G617), .b(G675), .O(G697) );
nand2 gate217( .a(G622), .b(G678), .O(G698) );
nand2 gate218( .a(G627), .b(G678), .O(G699) );
nand2 gate219( .a(G632), .b(G681), .O(G700) );
nand2 gate220( .a(G637), .b(G681), .O(G701) );
nand2 gate221( .a(G622), .b(G684), .O(G702) );
nand2 gate222( .a(G632), .b(G684), .O(G703) );
nand2 gate223( .a(G627), .b(G687), .O(G704) );

  xor2  gate1835(.a(G687), .b(G637), .O(gate224inter0));
  nand2 gate1836(.a(gate224inter0), .b(s_184), .O(gate224inter1));
  and2  gate1837(.a(G687), .b(G637), .O(gate224inter2));
  inv1  gate1838(.a(s_184), .O(gate224inter3));
  inv1  gate1839(.a(s_185), .O(gate224inter4));
  nand2 gate1840(.a(gate224inter4), .b(gate224inter3), .O(gate224inter5));
  nor2  gate1841(.a(gate224inter5), .b(gate224inter2), .O(gate224inter6));
  inv1  gate1842(.a(G637), .O(gate224inter7));
  inv1  gate1843(.a(G687), .O(gate224inter8));
  nand2 gate1844(.a(gate224inter8), .b(gate224inter7), .O(gate224inter9));
  nand2 gate1845(.a(s_185), .b(gate224inter3), .O(gate224inter10));
  nor2  gate1846(.a(gate224inter10), .b(gate224inter9), .O(gate224inter11));
  nor2  gate1847(.a(gate224inter11), .b(gate224inter6), .O(gate224inter12));
  nand2 gate1848(.a(gate224inter12), .b(gate224inter1), .O(G705));
nand2 gate225( .a(G690), .b(G691), .O(G706) );

  xor2  gate2521(.a(G693), .b(G692), .O(gate226inter0));
  nand2 gate2522(.a(gate226inter0), .b(s_282), .O(gate226inter1));
  and2  gate2523(.a(G693), .b(G692), .O(gate226inter2));
  inv1  gate2524(.a(s_282), .O(gate226inter3));
  inv1  gate2525(.a(s_283), .O(gate226inter4));
  nand2 gate2526(.a(gate226inter4), .b(gate226inter3), .O(gate226inter5));
  nor2  gate2527(.a(gate226inter5), .b(gate226inter2), .O(gate226inter6));
  inv1  gate2528(.a(G692), .O(gate226inter7));
  inv1  gate2529(.a(G693), .O(gate226inter8));
  nand2 gate2530(.a(gate226inter8), .b(gate226inter7), .O(gate226inter9));
  nand2 gate2531(.a(s_283), .b(gate226inter3), .O(gate226inter10));
  nor2  gate2532(.a(gate226inter10), .b(gate226inter9), .O(gate226inter11));
  nor2  gate2533(.a(gate226inter11), .b(gate226inter6), .O(gate226inter12));
  nand2 gate2534(.a(gate226inter12), .b(gate226inter1), .O(G709));
nand2 gate227( .a(G694), .b(G695), .O(G712) );
nand2 gate228( .a(G696), .b(G697), .O(G715) );
nand2 gate229( .a(G698), .b(G699), .O(G718) );
nand2 gate230( .a(G700), .b(G701), .O(G721) );

  xor2  gate1975(.a(G703), .b(G702), .O(gate231inter0));
  nand2 gate1976(.a(gate231inter0), .b(s_204), .O(gate231inter1));
  and2  gate1977(.a(G703), .b(G702), .O(gate231inter2));
  inv1  gate1978(.a(s_204), .O(gate231inter3));
  inv1  gate1979(.a(s_205), .O(gate231inter4));
  nand2 gate1980(.a(gate231inter4), .b(gate231inter3), .O(gate231inter5));
  nor2  gate1981(.a(gate231inter5), .b(gate231inter2), .O(gate231inter6));
  inv1  gate1982(.a(G702), .O(gate231inter7));
  inv1  gate1983(.a(G703), .O(gate231inter8));
  nand2 gate1984(.a(gate231inter8), .b(gate231inter7), .O(gate231inter9));
  nand2 gate1985(.a(s_205), .b(gate231inter3), .O(gate231inter10));
  nor2  gate1986(.a(gate231inter10), .b(gate231inter9), .O(gate231inter11));
  nor2  gate1987(.a(gate231inter11), .b(gate231inter6), .O(gate231inter12));
  nand2 gate1988(.a(gate231inter12), .b(gate231inter1), .O(G724));

  xor2  gate2437(.a(G705), .b(G704), .O(gate232inter0));
  nand2 gate2438(.a(gate232inter0), .b(s_270), .O(gate232inter1));
  and2  gate2439(.a(G705), .b(G704), .O(gate232inter2));
  inv1  gate2440(.a(s_270), .O(gate232inter3));
  inv1  gate2441(.a(s_271), .O(gate232inter4));
  nand2 gate2442(.a(gate232inter4), .b(gate232inter3), .O(gate232inter5));
  nor2  gate2443(.a(gate232inter5), .b(gate232inter2), .O(gate232inter6));
  inv1  gate2444(.a(G704), .O(gate232inter7));
  inv1  gate2445(.a(G705), .O(gate232inter8));
  nand2 gate2446(.a(gate232inter8), .b(gate232inter7), .O(gate232inter9));
  nand2 gate2447(.a(s_271), .b(gate232inter3), .O(gate232inter10));
  nor2  gate2448(.a(gate232inter10), .b(gate232inter9), .O(gate232inter11));
  nor2  gate2449(.a(gate232inter11), .b(gate232inter6), .O(gate232inter12));
  nand2 gate2450(.a(gate232inter12), .b(gate232inter1), .O(G727));

  xor2  gate1051(.a(G718), .b(G242), .O(gate233inter0));
  nand2 gate1052(.a(gate233inter0), .b(s_72), .O(gate233inter1));
  and2  gate1053(.a(G718), .b(G242), .O(gate233inter2));
  inv1  gate1054(.a(s_72), .O(gate233inter3));
  inv1  gate1055(.a(s_73), .O(gate233inter4));
  nand2 gate1056(.a(gate233inter4), .b(gate233inter3), .O(gate233inter5));
  nor2  gate1057(.a(gate233inter5), .b(gate233inter2), .O(gate233inter6));
  inv1  gate1058(.a(G242), .O(gate233inter7));
  inv1  gate1059(.a(G718), .O(gate233inter8));
  nand2 gate1060(.a(gate233inter8), .b(gate233inter7), .O(gate233inter9));
  nand2 gate1061(.a(s_73), .b(gate233inter3), .O(gate233inter10));
  nor2  gate1062(.a(gate233inter10), .b(gate233inter9), .O(gate233inter11));
  nor2  gate1063(.a(gate233inter11), .b(gate233inter6), .O(gate233inter12));
  nand2 gate1064(.a(gate233inter12), .b(gate233inter1), .O(G730));

  xor2  gate1107(.a(G721), .b(G245), .O(gate234inter0));
  nand2 gate1108(.a(gate234inter0), .b(s_80), .O(gate234inter1));
  and2  gate1109(.a(G721), .b(G245), .O(gate234inter2));
  inv1  gate1110(.a(s_80), .O(gate234inter3));
  inv1  gate1111(.a(s_81), .O(gate234inter4));
  nand2 gate1112(.a(gate234inter4), .b(gate234inter3), .O(gate234inter5));
  nor2  gate1113(.a(gate234inter5), .b(gate234inter2), .O(gate234inter6));
  inv1  gate1114(.a(G245), .O(gate234inter7));
  inv1  gate1115(.a(G721), .O(gate234inter8));
  nand2 gate1116(.a(gate234inter8), .b(gate234inter7), .O(gate234inter9));
  nand2 gate1117(.a(s_81), .b(gate234inter3), .O(gate234inter10));
  nor2  gate1118(.a(gate234inter10), .b(gate234inter9), .O(gate234inter11));
  nor2  gate1119(.a(gate234inter11), .b(gate234inter6), .O(gate234inter12));
  nand2 gate1120(.a(gate234inter12), .b(gate234inter1), .O(G733));
nand2 gate235( .a(G248), .b(G724), .O(G736) );

  xor2  gate2577(.a(G727), .b(G251), .O(gate236inter0));
  nand2 gate2578(.a(gate236inter0), .b(s_290), .O(gate236inter1));
  and2  gate2579(.a(G727), .b(G251), .O(gate236inter2));
  inv1  gate2580(.a(s_290), .O(gate236inter3));
  inv1  gate2581(.a(s_291), .O(gate236inter4));
  nand2 gate2582(.a(gate236inter4), .b(gate236inter3), .O(gate236inter5));
  nor2  gate2583(.a(gate236inter5), .b(gate236inter2), .O(gate236inter6));
  inv1  gate2584(.a(G251), .O(gate236inter7));
  inv1  gate2585(.a(G727), .O(gate236inter8));
  nand2 gate2586(.a(gate236inter8), .b(gate236inter7), .O(gate236inter9));
  nand2 gate2587(.a(s_291), .b(gate236inter3), .O(gate236inter10));
  nor2  gate2588(.a(gate236inter10), .b(gate236inter9), .O(gate236inter11));
  nor2  gate2589(.a(gate236inter11), .b(gate236inter6), .O(gate236inter12));
  nand2 gate2590(.a(gate236inter12), .b(gate236inter1), .O(G739));
nand2 gate237( .a(G254), .b(G706), .O(G742) );
nand2 gate238( .a(G257), .b(G709), .O(G745) );

  xor2  gate1513(.a(G712), .b(G260), .O(gate239inter0));
  nand2 gate1514(.a(gate239inter0), .b(s_138), .O(gate239inter1));
  and2  gate1515(.a(G712), .b(G260), .O(gate239inter2));
  inv1  gate1516(.a(s_138), .O(gate239inter3));
  inv1  gate1517(.a(s_139), .O(gate239inter4));
  nand2 gate1518(.a(gate239inter4), .b(gate239inter3), .O(gate239inter5));
  nor2  gate1519(.a(gate239inter5), .b(gate239inter2), .O(gate239inter6));
  inv1  gate1520(.a(G260), .O(gate239inter7));
  inv1  gate1521(.a(G712), .O(gate239inter8));
  nand2 gate1522(.a(gate239inter8), .b(gate239inter7), .O(gate239inter9));
  nand2 gate1523(.a(s_139), .b(gate239inter3), .O(gate239inter10));
  nor2  gate1524(.a(gate239inter10), .b(gate239inter9), .O(gate239inter11));
  nor2  gate1525(.a(gate239inter11), .b(gate239inter6), .O(gate239inter12));
  nand2 gate1526(.a(gate239inter12), .b(gate239inter1), .O(G748));
nand2 gate240( .a(G263), .b(G715), .O(G751) );
nand2 gate241( .a(G242), .b(G730), .O(G754) );
nand2 gate242( .a(G718), .b(G730), .O(G755) );

  xor2  gate1163(.a(G733), .b(G245), .O(gate243inter0));
  nand2 gate1164(.a(gate243inter0), .b(s_88), .O(gate243inter1));
  and2  gate1165(.a(G733), .b(G245), .O(gate243inter2));
  inv1  gate1166(.a(s_88), .O(gate243inter3));
  inv1  gate1167(.a(s_89), .O(gate243inter4));
  nand2 gate1168(.a(gate243inter4), .b(gate243inter3), .O(gate243inter5));
  nor2  gate1169(.a(gate243inter5), .b(gate243inter2), .O(gate243inter6));
  inv1  gate1170(.a(G245), .O(gate243inter7));
  inv1  gate1171(.a(G733), .O(gate243inter8));
  nand2 gate1172(.a(gate243inter8), .b(gate243inter7), .O(gate243inter9));
  nand2 gate1173(.a(s_89), .b(gate243inter3), .O(gate243inter10));
  nor2  gate1174(.a(gate243inter10), .b(gate243inter9), .O(gate243inter11));
  nor2  gate1175(.a(gate243inter11), .b(gate243inter6), .O(gate243inter12));
  nand2 gate1176(.a(gate243inter12), .b(gate243inter1), .O(G756));
nand2 gate244( .a(G721), .b(G733), .O(G757) );

  xor2  gate1723(.a(G736), .b(G248), .O(gate245inter0));
  nand2 gate1724(.a(gate245inter0), .b(s_168), .O(gate245inter1));
  and2  gate1725(.a(G736), .b(G248), .O(gate245inter2));
  inv1  gate1726(.a(s_168), .O(gate245inter3));
  inv1  gate1727(.a(s_169), .O(gate245inter4));
  nand2 gate1728(.a(gate245inter4), .b(gate245inter3), .O(gate245inter5));
  nor2  gate1729(.a(gate245inter5), .b(gate245inter2), .O(gate245inter6));
  inv1  gate1730(.a(G248), .O(gate245inter7));
  inv1  gate1731(.a(G736), .O(gate245inter8));
  nand2 gate1732(.a(gate245inter8), .b(gate245inter7), .O(gate245inter9));
  nand2 gate1733(.a(s_169), .b(gate245inter3), .O(gate245inter10));
  nor2  gate1734(.a(gate245inter10), .b(gate245inter9), .O(gate245inter11));
  nor2  gate1735(.a(gate245inter11), .b(gate245inter6), .O(gate245inter12));
  nand2 gate1736(.a(gate245inter12), .b(gate245inter1), .O(G758));
nand2 gate246( .a(G724), .b(G736), .O(G759) );

  xor2  gate813(.a(G739), .b(G251), .O(gate247inter0));
  nand2 gate814(.a(gate247inter0), .b(s_38), .O(gate247inter1));
  and2  gate815(.a(G739), .b(G251), .O(gate247inter2));
  inv1  gate816(.a(s_38), .O(gate247inter3));
  inv1  gate817(.a(s_39), .O(gate247inter4));
  nand2 gate818(.a(gate247inter4), .b(gate247inter3), .O(gate247inter5));
  nor2  gate819(.a(gate247inter5), .b(gate247inter2), .O(gate247inter6));
  inv1  gate820(.a(G251), .O(gate247inter7));
  inv1  gate821(.a(G739), .O(gate247inter8));
  nand2 gate822(.a(gate247inter8), .b(gate247inter7), .O(gate247inter9));
  nand2 gate823(.a(s_39), .b(gate247inter3), .O(gate247inter10));
  nor2  gate824(.a(gate247inter10), .b(gate247inter9), .O(gate247inter11));
  nor2  gate825(.a(gate247inter11), .b(gate247inter6), .O(gate247inter12));
  nand2 gate826(.a(gate247inter12), .b(gate247inter1), .O(G760));
nand2 gate248( .a(G727), .b(G739), .O(G761) );
nand2 gate249( .a(G254), .b(G742), .O(G762) );
nand2 gate250( .a(G706), .b(G742), .O(G763) );
nand2 gate251( .a(G257), .b(G745), .O(G764) );

  xor2  gate2199(.a(G745), .b(G709), .O(gate252inter0));
  nand2 gate2200(.a(gate252inter0), .b(s_236), .O(gate252inter1));
  and2  gate2201(.a(G745), .b(G709), .O(gate252inter2));
  inv1  gate2202(.a(s_236), .O(gate252inter3));
  inv1  gate2203(.a(s_237), .O(gate252inter4));
  nand2 gate2204(.a(gate252inter4), .b(gate252inter3), .O(gate252inter5));
  nor2  gate2205(.a(gate252inter5), .b(gate252inter2), .O(gate252inter6));
  inv1  gate2206(.a(G709), .O(gate252inter7));
  inv1  gate2207(.a(G745), .O(gate252inter8));
  nand2 gate2208(.a(gate252inter8), .b(gate252inter7), .O(gate252inter9));
  nand2 gate2209(.a(s_237), .b(gate252inter3), .O(gate252inter10));
  nor2  gate2210(.a(gate252inter10), .b(gate252inter9), .O(gate252inter11));
  nor2  gate2211(.a(gate252inter11), .b(gate252inter6), .O(gate252inter12));
  nand2 gate2212(.a(gate252inter12), .b(gate252inter1), .O(G765));
nand2 gate253( .a(G260), .b(G748), .O(G766) );

  xor2  gate575(.a(G748), .b(G712), .O(gate254inter0));
  nand2 gate576(.a(gate254inter0), .b(s_4), .O(gate254inter1));
  and2  gate577(.a(G748), .b(G712), .O(gate254inter2));
  inv1  gate578(.a(s_4), .O(gate254inter3));
  inv1  gate579(.a(s_5), .O(gate254inter4));
  nand2 gate580(.a(gate254inter4), .b(gate254inter3), .O(gate254inter5));
  nor2  gate581(.a(gate254inter5), .b(gate254inter2), .O(gate254inter6));
  inv1  gate582(.a(G712), .O(gate254inter7));
  inv1  gate583(.a(G748), .O(gate254inter8));
  nand2 gate584(.a(gate254inter8), .b(gate254inter7), .O(gate254inter9));
  nand2 gate585(.a(s_5), .b(gate254inter3), .O(gate254inter10));
  nor2  gate586(.a(gate254inter10), .b(gate254inter9), .O(gate254inter11));
  nor2  gate587(.a(gate254inter11), .b(gate254inter6), .O(gate254inter12));
  nand2 gate588(.a(gate254inter12), .b(gate254inter1), .O(G767));
nand2 gate255( .a(G263), .b(G751), .O(G768) );
nand2 gate256( .a(G715), .b(G751), .O(G769) );
nand2 gate257( .a(G754), .b(G755), .O(G770) );
nand2 gate258( .a(G756), .b(G757), .O(G773) );
nand2 gate259( .a(G758), .b(G759), .O(G776) );
nand2 gate260( .a(G760), .b(G761), .O(G779) );

  xor2  gate2591(.a(G763), .b(G762), .O(gate261inter0));
  nand2 gate2592(.a(gate261inter0), .b(s_292), .O(gate261inter1));
  and2  gate2593(.a(G763), .b(G762), .O(gate261inter2));
  inv1  gate2594(.a(s_292), .O(gate261inter3));
  inv1  gate2595(.a(s_293), .O(gate261inter4));
  nand2 gate2596(.a(gate261inter4), .b(gate261inter3), .O(gate261inter5));
  nor2  gate2597(.a(gate261inter5), .b(gate261inter2), .O(gate261inter6));
  inv1  gate2598(.a(G762), .O(gate261inter7));
  inv1  gate2599(.a(G763), .O(gate261inter8));
  nand2 gate2600(.a(gate261inter8), .b(gate261inter7), .O(gate261inter9));
  nand2 gate2601(.a(s_293), .b(gate261inter3), .O(gate261inter10));
  nor2  gate2602(.a(gate261inter10), .b(gate261inter9), .O(gate261inter11));
  nor2  gate2603(.a(gate261inter11), .b(gate261inter6), .O(gate261inter12));
  nand2 gate2604(.a(gate261inter12), .b(gate261inter1), .O(G782));
nand2 gate262( .a(G764), .b(G765), .O(G785) );

  xor2  gate1289(.a(G767), .b(G766), .O(gate263inter0));
  nand2 gate1290(.a(gate263inter0), .b(s_106), .O(gate263inter1));
  and2  gate1291(.a(G767), .b(G766), .O(gate263inter2));
  inv1  gate1292(.a(s_106), .O(gate263inter3));
  inv1  gate1293(.a(s_107), .O(gate263inter4));
  nand2 gate1294(.a(gate263inter4), .b(gate263inter3), .O(gate263inter5));
  nor2  gate1295(.a(gate263inter5), .b(gate263inter2), .O(gate263inter6));
  inv1  gate1296(.a(G766), .O(gate263inter7));
  inv1  gate1297(.a(G767), .O(gate263inter8));
  nand2 gate1298(.a(gate263inter8), .b(gate263inter7), .O(gate263inter9));
  nand2 gate1299(.a(s_107), .b(gate263inter3), .O(gate263inter10));
  nor2  gate1300(.a(gate263inter10), .b(gate263inter9), .O(gate263inter11));
  nor2  gate1301(.a(gate263inter11), .b(gate263inter6), .O(gate263inter12));
  nand2 gate1302(.a(gate263inter12), .b(gate263inter1), .O(G788));

  xor2  gate2185(.a(G769), .b(G768), .O(gate264inter0));
  nand2 gate2186(.a(gate264inter0), .b(s_234), .O(gate264inter1));
  and2  gate2187(.a(G769), .b(G768), .O(gate264inter2));
  inv1  gate2188(.a(s_234), .O(gate264inter3));
  inv1  gate2189(.a(s_235), .O(gate264inter4));
  nand2 gate2190(.a(gate264inter4), .b(gate264inter3), .O(gate264inter5));
  nor2  gate2191(.a(gate264inter5), .b(gate264inter2), .O(gate264inter6));
  inv1  gate2192(.a(G768), .O(gate264inter7));
  inv1  gate2193(.a(G769), .O(gate264inter8));
  nand2 gate2194(.a(gate264inter8), .b(gate264inter7), .O(gate264inter9));
  nand2 gate2195(.a(s_235), .b(gate264inter3), .O(gate264inter10));
  nor2  gate2196(.a(gate264inter10), .b(gate264inter9), .O(gate264inter11));
  nor2  gate2197(.a(gate264inter11), .b(gate264inter6), .O(gate264inter12));
  nand2 gate2198(.a(gate264inter12), .b(gate264inter1), .O(G791));

  xor2  gate2353(.a(G770), .b(G642), .O(gate265inter0));
  nand2 gate2354(.a(gate265inter0), .b(s_258), .O(gate265inter1));
  and2  gate2355(.a(G770), .b(G642), .O(gate265inter2));
  inv1  gate2356(.a(s_258), .O(gate265inter3));
  inv1  gate2357(.a(s_259), .O(gate265inter4));
  nand2 gate2358(.a(gate265inter4), .b(gate265inter3), .O(gate265inter5));
  nor2  gate2359(.a(gate265inter5), .b(gate265inter2), .O(gate265inter6));
  inv1  gate2360(.a(G642), .O(gate265inter7));
  inv1  gate2361(.a(G770), .O(gate265inter8));
  nand2 gate2362(.a(gate265inter8), .b(gate265inter7), .O(gate265inter9));
  nand2 gate2363(.a(s_259), .b(gate265inter3), .O(gate265inter10));
  nor2  gate2364(.a(gate265inter10), .b(gate265inter9), .O(gate265inter11));
  nor2  gate2365(.a(gate265inter11), .b(gate265inter6), .O(gate265inter12));
  nand2 gate2366(.a(gate265inter12), .b(gate265inter1), .O(G794));
nand2 gate266( .a(G645), .b(G773), .O(G797) );
nand2 gate267( .a(G648), .b(G776), .O(G800) );
nand2 gate268( .a(G651), .b(G779), .O(G803) );

  xor2  gate2283(.a(G782), .b(G654), .O(gate269inter0));
  nand2 gate2284(.a(gate269inter0), .b(s_248), .O(gate269inter1));
  and2  gate2285(.a(G782), .b(G654), .O(gate269inter2));
  inv1  gate2286(.a(s_248), .O(gate269inter3));
  inv1  gate2287(.a(s_249), .O(gate269inter4));
  nand2 gate2288(.a(gate269inter4), .b(gate269inter3), .O(gate269inter5));
  nor2  gate2289(.a(gate269inter5), .b(gate269inter2), .O(gate269inter6));
  inv1  gate2290(.a(G654), .O(gate269inter7));
  inv1  gate2291(.a(G782), .O(gate269inter8));
  nand2 gate2292(.a(gate269inter8), .b(gate269inter7), .O(gate269inter9));
  nand2 gate2293(.a(s_249), .b(gate269inter3), .O(gate269inter10));
  nor2  gate2294(.a(gate269inter10), .b(gate269inter9), .O(gate269inter11));
  nor2  gate2295(.a(gate269inter11), .b(gate269inter6), .O(gate269inter12));
  nand2 gate2296(.a(gate269inter12), .b(gate269inter1), .O(G806));
nand2 gate270( .a(G657), .b(G785), .O(G809) );
nand2 gate271( .a(G660), .b(G788), .O(G812) );

  xor2  gate2115(.a(G791), .b(G663), .O(gate272inter0));
  nand2 gate2116(.a(gate272inter0), .b(s_224), .O(gate272inter1));
  and2  gate2117(.a(G791), .b(G663), .O(gate272inter2));
  inv1  gate2118(.a(s_224), .O(gate272inter3));
  inv1  gate2119(.a(s_225), .O(gate272inter4));
  nand2 gate2120(.a(gate272inter4), .b(gate272inter3), .O(gate272inter5));
  nor2  gate2121(.a(gate272inter5), .b(gate272inter2), .O(gate272inter6));
  inv1  gate2122(.a(G663), .O(gate272inter7));
  inv1  gate2123(.a(G791), .O(gate272inter8));
  nand2 gate2124(.a(gate272inter8), .b(gate272inter7), .O(gate272inter9));
  nand2 gate2125(.a(s_225), .b(gate272inter3), .O(gate272inter10));
  nor2  gate2126(.a(gate272inter10), .b(gate272inter9), .O(gate272inter11));
  nor2  gate2127(.a(gate272inter11), .b(gate272inter6), .O(gate272inter12));
  nand2 gate2128(.a(gate272inter12), .b(gate272inter1), .O(G815));

  xor2  gate687(.a(G794), .b(G642), .O(gate273inter0));
  nand2 gate688(.a(gate273inter0), .b(s_20), .O(gate273inter1));
  and2  gate689(.a(G794), .b(G642), .O(gate273inter2));
  inv1  gate690(.a(s_20), .O(gate273inter3));
  inv1  gate691(.a(s_21), .O(gate273inter4));
  nand2 gate692(.a(gate273inter4), .b(gate273inter3), .O(gate273inter5));
  nor2  gate693(.a(gate273inter5), .b(gate273inter2), .O(gate273inter6));
  inv1  gate694(.a(G642), .O(gate273inter7));
  inv1  gate695(.a(G794), .O(gate273inter8));
  nand2 gate696(.a(gate273inter8), .b(gate273inter7), .O(gate273inter9));
  nand2 gate697(.a(s_21), .b(gate273inter3), .O(gate273inter10));
  nor2  gate698(.a(gate273inter10), .b(gate273inter9), .O(gate273inter11));
  nor2  gate699(.a(gate273inter11), .b(gate273inter6), .O(gate273inter12));
  nand2 gate700(.a(gate273inter12), .b(gate273inter1), .O(G818));

  xor2  gate2563(.a(G794), .b(G770), .O(gate274inter0));
  nand2 gate2564(.a(gate274inter0), .b(s_288), .O(gate274inter1));
  and2  gate2565(.a(G794), .b(G770), .O(gate274inter2));
  inv1  gate2566(.a(s_288), .O(gate274inter3));
  inv1  gate2567(.a(s_289), .O(gate274inter4));
  nand2 gate2568(.a(gate274inter4), .b(gate274inter3), .O(gate274inter5));
  nor2  gate2569(.a(gate274inter5), .b(gate274inter2), .O(gate274inter6));
  inv1  gate2570(.a(G770), .O(gate274inter7));
  inv1  gate2571(.a(G794), .O(gate274inter8));
  nand2 gate2572(.a(gate274inter8), .b(gate274inter7), .O(gate274inter9));
  nand2 gate2573(.a(s_289), .b(gate274inter3), .O(gate274inter10));
  nor2  gate2574(.a(gate274inter10), .b(gate274inter9), .O(gate274inter11));
  nor2  gate2575(.a(gate274inter11), .b(gate274inter6), .O(gate274inter12));
  nand2 gate2576(.a(gate274inter12), .b(gate274inter1), .O(G819));
nand2 gate275( .a(G645), .b(G797), .O(G820) );
nand2 gate276( .a(G773), .b(G797), .O(G821) );
nand2 gate277( .a(G648), .b(G800), .O(G822) );

  xor2  gate1387(.a(G800), .b(G776), .O(gate278inter0));
  nand2 gate1388(.a(gate278inter0), .b(s_120), .O(gate278inter1));
  and2  gate1389(.a(G800), .b(G776), .O(gate278inter2));
  inv1  gate1390(.a(s_120), .O(gate278inter3));
  inv1  gate1391(.a(s_121), .O(gate278inter4));
  nand2 gate1392(.a(gate278inter4), .b(gate278inter3), .O(gate278inter5));
  nor2  gate1393(.a(gate278inter5), .b(gate278inter2), .O(gate278inter6));
  inv1  gate1394(.a(G776), .O(gate278inter7));
  inv1  gate1395(.a(G800), .O(gate278inter8));
  nand2 gate1396(.a(gate278inter8), .b(gate278inter7), .O(gate278inter9));
  nand2 gate1397(.a(s_121), .b(gate278inter3), .O(gate278inter10));
  nor2  gate1398(.a(gate278inter10), .b(gate278inter9), .O(gate278inter11));
  nor2  gate1399(.a(gate278inter11), .b(gate278inter6), .O(gate278inter12));
  nand2 gate1400(.a(gate278inter12), .b(gate278inter1), .O(G823));
nand2 gate279( .a(G651), .b(G803), .O(G824) );
nand2 gate280( .a(G779), .b(G803), .O(G825) );
nand2 gate281( .a(G654), .b(G806), .O(G826) );

  xor2  gate785(.a(G806), .b(G782), .O(gate282inter0));
  nand2 gate786(.a(gate282inter0), .b(s_34), .O(gate282inter1));
  and2  gate787(.a(G806), .b(G782), .O(gate282inter2));
  inv1  gate788(.a(s_34), .O(gate282inter3));
  inv1  gate789(.a(s_35), .O(gate282inter4));
  nand2 gate790(.a(gate282inter4), .b(gate282inter3), .O(gate282inter5));
  nor2  gate791(.a(gate282inter5), .b(gate282inter2), .O(gate282inter6));
  inv1  gate792(.a(G782), .O(gate282inter7));
  inv1  gate793(.a(G806), .O(gate282inter8));
  nand2 gate794(.a(gate282inter8), .b(gate282inter7), .O(gate282inter9));
  nand2 gate795(.a(s_35), .b(gate282inter3), .O(gate282inter10));
  nor2  gate796(.a(gate282inter10), .b(gate282inter9), .O(gate282inter11));
  nor2  gate797(.a(gate282inter11), .b(gate282inter6), .O(gate282inter12));
  nand2 gate798(.a(gate282inter12), .b(gate282inter1), .O(G827));
nand2 gate283( .a(G657), .b(G809), .O(G828) );

  xor2  gate1807(.a(G809), .b(G785), .O(gate284inter0));
  nand2 gate1808(.a(gate284inter0), .b(s_180), .O(gate284inter1));
  and2  gate1809(.a(G809), .b(G785), .O(gate284inter2));
  inv1  gate1810(.a(s_180), .O(gate284inter3));
  inv1  gate1811(.a(s_181), .O(gate284inter4));
  nand2 gate1812(.a(gate284inter4), .b(gate284inter3), .O(gate284inter5));
  nor2  gate1813(.a(gate284inter5), .b(gate284inter2), .O(gate284inter6));
  inv1  gate1814(.a(G785), .O(gate284inter7));
  inv1  gate1815(.a(G809), .O(gate284inter8));
  nand2 gate1816(.a(gate284inter8), .b(gate284inter7), .O(gate284inter9));
  nand2 gate1817(.a(s_181), .b(gate284inter3), .O(gate284inter10));
  nor2  gate1818(.a(gate284inter10), .b(gate284inter9), .O(gate284inter11));
  nor2  gate1819(.a(gate284inter11), .b(gate284inter6), .O(gate284inter12));
  nand2 gate1820(.a(gate284inter12), .b(gate284inter1), .O(G829));

  xor2  gate1583(.a(G812), .b(G660), .O(gate285inter0));
  nand2 gate1584(.a(gate285inter0), .b(s_148), .O(gate285inter1));
  and2  gate1585(.a(G812), .b(G660), .O(gate285inter2));
  inv1  gate1586(.a(s_148), .O(gate285inter3));
  inv1  gate1587(.a(s_149), .O(gate285inter4));
  nand2 gate1588(.a(gate285inter4), .b(gate285inter3), .O(gate285inter5));
  nor2  gate1589(.a(gate285inter5), .b(gate285inter2), .O(gate285inter6));
  inv1  gate1590(.a(G660), .O(gate285inter7));
  inv1  gate1591(.a(G812), .O(gate285inter8));
  nand2 gate1592(.a(gate285inter8), .b(gate285inter7), .O(gate285inter9));
  nand2 gate1593(.a(s_149), .b(gate285inter3), .O(gate285inter10));
  nor2  gate1594(.a(gate285inter10), .b(gate285inter9), .O(gate285inter11));
  nor2  gate1595(.a(gate285inter11), .b(gate285inter6), .O(gate285inter12));
  nand2 gate1596(.a(gate285inter12), .b(gate285inter1), .O(G830));
nand2 gate286( .a(G788), .b(G812), .O(G831) );
nand2 gate287( .a(G663), .b(G815), .O(G832) );
nand2 gate288( .a(G791), .b(G815), .O(G833) );
nand2 gate289( .a(G818), .b(G819), .O(G834) );
nand2 gate290( .a(G820), .b(G821), .O(G847) );
nand2 gate291( .a(G822), .b(G823), .O(G860) );
nand2 gate292( .a(G824), .b(G825), .O(G873) );
nand2 gate293( .a(G828), .b(G829), .O(G886) );

  xor2  gate1681(.a(G833), .b(G832), .O(gate294inter0));
  nand2 gate1682(.a(gate294inter0), .b(s_162), .O(gate294inter1));
  and2  gate1683(.a(G833), .b(G832), .O(gate294inter2));
  inv1  gate1684(.a(s_162), .O(gate294inter3));
  inv1  gate1685(.a(s_163), .O(gate294inter4));
  nand2 gate1686(.a(gate294inter4), .b(gate294inter3), .O(gate294inter5));
  nor2  gate1687(.a(gate294inter5), .b(gate294inter2), .O(gate294inter6));
  inv1  gate1688(.a(G832), .O(gate294inter7));
  inv1  gate1689(.a(G833), .O(gate294inter8));
  nand2 gate1690(.a(gate294inter8), .b(gate294inter7), .O(gate294inter9));
  nand2 gate1691(.a(s_163), .b(gate294inter3), .O(gate294inter10));
  nor2  gate1692(.a(gate294inter10), .b(gate294inter9), .O(gate294inter11));
  nor2  gate1693(.a(gate294inter11), .b(gate294inter6), .O(gate294inter12));
  nand2 gate1694(.a(gate294inter12), .b(gate294inter1), .O(G899));
nand2 gate295( .a(G830), .b(G831), .O(G912) );
nand2 gate296( .a(G826), .b(G827), .O(G925) );
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );
nand2 gate387( .a(G1), .b(G1036), .O(G1132) );

  xor2  gate1821(.a(G1039), .b(G2), .O(gate388inter0));
  nand2 gate1822(.a(gate388inter0), .b(s_182), .O(gate388inter1));
  and2  gate1823(.a(G1039), .b(G2), .O(gate388inter2));
  inv1  gate1824(.a(s_182), .O(gate388inter3));
  inv1  gate1825(.a(s_183), .O(gate388inter4));
  nand2 gate1826(.a(gate388inter4), .b(gate388inter3), .O(gate388inter5));
  nor2  gate1827(.a(gate388inter5), .b(gate388inter2), .O(gate388inter6));
  inv1  gate1828(.a(G2), .O(gate388inter7));
  inv1  gate1829(.a(G1039), .O(gate388inter8));
  nand2 gate1830(.a(gate388inter8), .b(gate388inter7), .O(gate388inter9));
  nand2 gate1831(.a(s_183), .b(gate388inter3), .O(gate388inter10));
  nor2  gate1832(.a(gate388inter10), .b(gate388inter9), .O(gate388inter11));
  nor2  gate1833(.a(gate388inter11), .b(gate388inter6), .O(gate388inter12));
  nand2 gate1834(.a(gate388inter12), .b(gate388inter1), .O(G1135));
nand2 gate389( .a(G3), .b(G1042), .O(G1138) );
nand2 gate390( .a(G4), .b(G1045), .O(G1141) );

  xor2  gate799(.a(G1048), .b(G5), .O(gate391inter0));
  nand2 gate800(.a(gate391inter0), .b(s_36), .O(gate391inter1));
  and2  gate801(.a(G1048), .b(G5), .O(gate391inter2));
  inv1  gate802(.a(s_36), .O(gate391inter3));
  inv1  gate803(.a(s_37), .O(gate391inter4));
  nand2 gate804(.a(gate391inter4), .b(gate391inter3), .O(gate391inter5));
  nor2  gate805(.a(gate391inter5), .b(gate391inter2), .O(gate391inter6));
  inv1  gate806(.a(G5), .O(gate391inter7));
  inv1  gate807(.a(G1048), .O(gate391inter8));
  nand2 gate808(.a(gate391inter8), .b(gate391inter7), .O(gate391inter9));
  nand2 gate809(.a(s_37), .b(gate391inter3), .O(gate391inter10));
  nor2  gate810(.a(gate391inter10), .b(gate391inter9), .O(gate391inter11));
  nor2  gate811(.a(gate391inter11), .b(gate391inter6), .O(gate391inter12));
  nand2 gate812(.a(gate391inter12), .b(gate391inter1), .O(G1144));

  xor2  gate1947(.a(G1051), .b(G6), .O(gate392inter0));
  nand2 gate1948(.a(gate392inter0), .b(s_200), .O(gate392inter1));
  and2  gate1949(.a(G1051), .b(G6), .O(gate392inter2));
  inv1  gate1950(.a(s_200), .O(gate392inter3));
  inv1  gate1951(.a(s_201), .O(gate392inter4));
  nand2 gate1952(.a(gate392inter4), .b(gate392inter3), .O(gate392inter5));
  nor2  gate1953(.a(gate392inter5), .b(gate392inter2), .O(gate392inter6));
  inv1  gate1954(.a(G6), .O(gate392inter7));
  inv1  gate1955(.a(G1051), .O(gate392inter8));
  nand2 gate1956(.a(gate392inter8), .b(gate392inter7), .O(gate392inter9));
  nand2 gate1957(.a(s_201), .b(gate392inter3), .O(gate392inter10));
  nor2  gate1958(.a(gate392inter10), .b(gate392inter9), .O(gate392inter11));
  nor2  gate1959(.a(gate392inter11), .b(gate392inter6), .O(gate392inter12));
  nand2 gate1960(.a(gate392inter12), .b(gate392inter1), .O(G1147));
nand2 gate393( .a(G7), .b(G1054), .O(G1150) );

  xor2  gate1233(.a(G1057), .b(G8), .O(gate394inter0));
  nand2 gate1234(.a(gate394inter0), .b(s_98), .O(gate394inter1));
  and2  gate1235(.a(G1057), .b(G8), .O(gate394inter2));
  inv1  gate1236(.a(s_98), .O(gate394inter3));
  inv1  gate1237(.a(s_99), .O(gate394inter4));
  nand2 gate1238(.a(gate394inter4), .b(gate394inter3), .O(gate394inter5));
  nor2  gate1239(.a(gate394inter5), .b(gate394inter2), .O(gate394inter6));
  inv1  gate1240(.a(G8), .O(gate394inter7));
  inv1  gate1241(.a(G1057), .O(gate394inter8));
  nand2 gate1242(.a(gate394inter8), .b(gate394inter7), .O(gate394inter9));
  nand2 gate1243(.a(s_99), .b(gate394inter3), .O(gate394inter10));
  nor2  gate1244(.a(gate394inter10), .b(gate394inter9), .O(gate394inter11));
  nor2  gate1245(.a(gate394inter11), .b(gate394inter6), .O(gate394inter12));
  nand2 gate1246(.a(gate394inter12), .b(gate394inter1), .O(G1153));
nand2 gate395( .a(G9), .b(G1060), .O(G1156) );
nand2 gate396( .a(G10), .b(G1063), .O(G1159) );

  xor2  gate2017(.a(G1066), .b(G11), .O(gate397inter0));
  nand2 gate2018(.a(gate397inter0), .b(s_210), .O(gate397inter1));
  and2  gate2019(.a(G1066), .b(G11), .O(gate397inter2));
  inv1  gate2020(.a(s_210), .O(gate397inter3));
  inv1  gate2021(.a(s_211), .O(gate397inter4));
  nand2 gate2022(.a(gate397inter4), .b(gate397inter3), .O(gate397inter5));
  nor2  gate2023(.a(gate397inter5), .b(gate397inter2), .O(gate397inter6));
  inv1  gate2024(.a(G11), .O(gate397inter7));
  inv1  gate2025(.a(G1066), .O(gate397inter8));
  nand2 gate2026(.a(gate397inter8), .b(gate397inter7), .O(gate397inter9));
  nand2 gate2027(.a(s_211), .b(gate397inter3), .O(gate397inter10));
  nor2  gate2028(.a(gate397inter10), .b(gate397inter9), .O(gate397inter11));
  nor2  gate2029(.a(gate397inter11), .b(gate397inter6), .O(gate397inter12));
  nand2 gate2030(.a(gate397inter12), .b(gate397inter1), .O(G1162));
nand2 gate398( .a(G12), .b(G1069), .O(G1165) );
nand2 gate399( .a(G13), .b(G1072), .O(G1168) );

  xor2  gate2003(.a(G1075), .b(G14), .O(gate400inter0));
  nand2 gate2004(.a(gate400inter0), .b(s_208), .O(gate400inter1));
  and2  gate2005(.a(G1075), .b(G14), .O(gate400inter2));
  inv1  gate2006(.a(s_208), .O(gate400inter3));
  inv1  gate2007(.a(s_209), .O(gate400inter4));
  nand2 gate2008(.a(gate400inter4), .b(gate400inter3), .O(gate400inter5));
  nor2  gate2009(.a(gate400inter5), .b(gate400inter2), .O(gate400inter6));
  inv1  gate2010(.a(G14), .O(gate400inter7));
  inv1  gate2011(.a(G1075), .O(gate400inter8));
  nand2 gate2012(.a(gate400inter8), .b(gate400inter7), .O(gate400inter9));
  nand2 gate2013(.a(s_209), .b(gate400inter3), .O(gate400inter10));
  nor2  gate2014(.a(gate400inter10), .b(gate400inter9), .O(gate400inter11));
  nor2  gate2015(.a(gate400inter11), .b(gate400inter6), .O(gate400inter12));
  nand2 gate2016(.a(gate400inter12), .b(gate400inter1), .O(G1171));

  xor2  gate1849(.a(G1078), .b(G15), .O(gate401inter0));
  nand2 gate1850(.a(gate401inter0), .b(s_186), .O(gate401inter1));
  and2  gate1851(.a(G1078), .b(G15), .O(gate401inter2));
  inv1  gate1852(.a(s_186), .O(gate401inter3));
  inv1  gate1853(.a(s_187), .O(gate401inter4));
  nand2 gate1854(.a(gate401inter4), .b(gate401inter3), .O(gate401inter5));
  nor2  gate1855(.a(gate401inter5), .b(gate401inter2), .O(gate401inter6));
  inv1  gate1856(.a(G15), .O(gate401inter7));
  inv1  gate1857(.a(G1078), .O(gate401inter8));
  nand2 gate1858(.a(gate401inter8), .b(gate401inter7), .O(gate401inter9));
  nand2 gate1859(.a(s_187), .b(gate401inter3), .O(gate401inter10));
  nor2  gate1860(.a(gate401inter10), .b(gate401inter9), .O(gate401inter11));
  nor2  gate1861(.a(gate401inter11), .b(gate401inter6), .O(gate401inter12));
  nand2 gate1862(.a(gate401inter12), .b(gate401inter1), .O(G1174));

  xor2  gate1891(.a(G1081), .b(G16), .O(gate402inter0));
  nand2 gate1892(.a(gate402inter0), .b(s_192), .O(gate402inter1));
  and2  gate1893(.a(G1081), .b(G16), .O(gate402inter2));
  inv1  gate1894(.a(s_192), .O(gate402inter3));
  inv1  gate1895(.a(s_193), .O(gate402inter4));
  nand2 gate1896(.a(gate402inter4), .b(gate402inter3), .O(gate402inter5));
  nor2  gate1897(.a(gate402inter5), .b(gate402inter2), .O(gate402inter6));
  inv1  gate1898(.a(G16), .O(gate402inter7));
  inv1  gate1899(.a(G1081), .O(gate402inter8));
  nand2 gate1900(.a(gate402inter8), .b(gate402inter7), .O(gate402inter9));
  nand2 gate1901(.a(s_193), .b(gate402inter3), .O(gate402inter10));
  nor2  gate1902(.a(gate402inter10), .b(gate402inter9), .O(gate402inter11));
  nor2  gate1903(.a(gate402inter11), .b(gate402inter6), .O(gate402inter12));
  nand2 gate1904(.a(gate402inter12), .b(gate402inter1), .O(G1177));
nand2 gate403( .a(G17), .b(G1084), .O(G1180) );
nand2 gate404( .a(G18), .b(G1087), .O(G1183) );
nand2 gate405( .a(G19), .b(G1090), .O(G1186) );
nand2 gate406( .a(G20), .b(G1093), .O(G1189) );
nand2 gate407( .a(G21), .b(G1096), .O(G1192) );

  xor2  gate673(.a(G1099), .b(G22), .O(gate408inter0));
  nand2 gate674(.a(gate408inter0), .b(s_18), .O(gate408inter1));
  and2  gate675(.a(G1099), .b(G22), .O(gate408inter2));
  inv1  gate676(.a(s_18), .O(gate408inter3));
  inv1  gate677(.a(s_19), .O(gate408inter4));
  nand2 gate678(.a(gate408inter4), .b(gate408inter3), .O(gate408inter5));
  nor2  gate679(.a(gate408inter5), .b(gate408inter2), .O(gate408inter6));
  inv1  gate680(.a(G22), .O(gate408inter7));
  inv1  gate681(.a(G1099), .O(gate408inter8));
  nand2 gate682(.a(gate408inter8), .b(gate408inter7), .O(gate408inter9));
  nand2 gate683(.a(s_19), .b(gate408inter3), .O(gate408inter10));
  nor2  gate684(.a(gate408inter10), .b(gate408inter9), .O(gate408inter11));
  nor2  gate685(.a(gate408inter11), .b(gate408inter6), .O(gate408inter12));
  nand2 gate686(.a(gate408inter12), .b(gate408inter1), .O(G1195));
nand2 gate409( .a(G23), .b(G1102), .O(G1198) );

  xor2  gate1933(.a(G1105), .b(G24), .O(gate410inter0));
  nand2 gate1934(.a(gate410inter0), .b(s_198), .O(gate410inter1));
  and2  gate1935(.a(G1105), .b(G24), .O(gate410inter2));
  inv1  gate1936(.a(s_198), .O(gate410inter3));
  inv1  gate1937(.a(s_199), .O(gate410inter4));
  nand2 gate1938(.a(gate410inter4), .b(gate410inter3), .O(gate410inter5));
  nor2  gate1939(.a(gate410inter5), .b(gate410inter2), .O(gate410inter6));
  inv1  gate1940(.a(G24), .O(gate410inter7));
  inv1  gate1941(.a(G1105), .O(gate410inter8));
  nand2 gate1942(.a(gate410inter8), .b(gate410inter7), .O(gate410inter9));
  nand2 gate1943(.a(s_199), .b(gate410inter3), .O(gate410inter10));
  nor2  gate1944(.a(gate410inter10), .b(gate410inter9), .O(gate410inter11));
  nor2  gate1945(.a(gate410inter11), .b(gate410inter6), .O(gate410inter12));
  nand2 gate1946(.a(gate410inter12), .b(gate410inter1), .O(G1201));
nand2 gate411( .a(G25), .b(G1108), .O(G1204) );
nand2 gate412( .a(G26), .b(G1111), .O(G1207) );
nand2 gate413( .a(G27), .b(G1114), .O(G1210) );
nand2 gate414( .a(G28), .b(G1117), .O(G1213) );
nand2 gate415( .a(G29), .b(G1120), .O(G1216) );
nand2 gate416( .a(G30), .b(G1123), .O(G1219) );
nand2 gate417( .a(G31), .b(G1126), .O(G1222) );
nand2 gate418( .a(G32), .b(G1129), .O(G1225) );
nand2 gate419( .a(G1), .b(G1132), .O(G1228) );
nand2 gate420( .a(G1036), .b(G1132), .O(G1229) );

  xor2  gate2507(.a(G1135), .b(G2), .O(gate421inter0));
  nand2 gate2508(.a(gate421inter0), .b(s_280), .O(gate421inter1));
  and2  gate2509(.a(G1135), .b(G2), .O(gate421inter2));
  inv1  gate2510(.a(s_280), .O(gate421inter3));
  inv1  gate2511(.a(s_281), .O(gate421inter4));
  nand2 gate2512(.a(gate421inter4), .b(gate421inter3), .O(gate421inter5));
  nor2  gate2513(.a(gate421inter5), .b(gate421inter2), .O(gate421inter6));
  inv1  gate2514(.a(G2), .O(gate421inter7));
  inv1  gate2515(.a(G1135), .O(gate421inter8));
  nand2 gate2516(.a(gate421inter8), .b(gate421inter7), .O(gate421inter9));
  nand2 gate2517(.a(s_281), .b(gate421inter3), .O(gate421inter10));
  nor2  gate2518(.a(gate421inter10), .b(gate421inter9), .O(gate421inter11));
  nor2  gate2519(.a(gate421inter11), .b(gate421inter6), .O(gate421inter12));
  nand2 gate2520(.a(gate421inter12), .b(gate421inter1), .O(G1230));
nand2 gate422( .a(G1039), .b(G1135), .O(G1231) );
nand2 gate423( .a(G3), .b(G1138), .O(G1232) );
nand2 gate424( .a(G1042), .b(G1138), .O(G1233) );
nand2 gate425( .a(G4), .b(G1141), .O(G1234) );

  xor2  gate897(.a(G1141), .b(G1045), .O(gate426inter0));
  nand2 gate898(.a(gate426inter0), .b(s_50), .O(gate426inter1));
  and2  gate899(.a(G1141), .b(G1045), .O(gate426inter2));
  inv1  gate900(.a(s_50), .O(gate426inter3));
  inv1  gate901(.a(s_51), .O(gate426inter4));
  nand2 gate902(.a(gate426inter4), .b(gate426inter3), .O(gate426inter5));
  nor2  gate903(.a(gate426inter5), .b(gate426inter2), .O(gate426inter6));
  inv1  gate904(.a(G1045), .O(gate426inter7));
  inv1  gate905(.a(G1141), .O(gate426inter8));
  nand2 gate906(.a(gate426inter8), .b(gate426inter7), .O(gate426inter9));
  nand2 gate907(.a(s_51), .b(gate426inter3), .O(gate426inter10));
  nor2  gate908(.a(gate426inter10), .b(gate426inter9), .O(gate426inter11));
  nor2  gate909(.a(gate426inter11), .b(gate426inter6), .O(gate426inter12));
  nand2 gate910(.a(gate426inter12), .b(gate426inter1), .O(G1235));
nand2 gate427( .a(G5), .b(G1144), .O(G1236) );

  xor2  gate2367(.a(G1144), .b(G1048), .O(gate428inter0));
  nand2 gate2368(.a(gate428inter0), .b(s_260), .O(gate428inter1));
  and2  gate2369(.a(G1144), .b(G1048), .O(gate428inter2));
  inv1  gate2370(.a(s_260), .O(gate428inter3));
  inv1  gate2371(.a(s_261), .O(gate428inter4));
  nand2 gate2372(.a(gate428inter4), .b(gate428inter3), .O(gate428inter5));
  nor2  gate2373(.a(gate428inter5), .b(gate428inter2), .O(gate428inter6));
  inv1  gate2374(.a(G1048), .O(gate428inter7));
  inv1  gate2375(.a(G1144), .O(gate428inter8));
  nand2 gate2376(.a(gate428inter8), .b(gate428inter7), .O(gate428inter9));
  nand2 gate2377(.a(s_261), .b(gate428inter3), .O(gate428inter10));
  nor2  gate2378(.a(gate428inter10), .b(gate428inter9), .O(gate428inter11));
  nor2  gate2379(.a(gate428inter11), .b(gate428inter6), .O(gate428inter12));
  nand2 gate2380(.a(gate428inter12), .b(gate428inter1), .O(G1237));
nand2 gate429( .a(G6), .b(G1147), .O(G1238) );

  xor2  gate953(.a(G1147), .b(G1051), .O(gate430inter0));
  nand2 gate954(.a(gate430inter0), .b(s_58), .O(gate430inter1));
  and2  gate955(.a(G1147), .b(G1051), .O(gate430inter2));
  inv1  gate956(.a(s_58), .O(gate430inter3));
  inv1  gate957(.a(s_59), .O(gate430inter4));
  nand2 gate958(.a(gate430inter4), .b(gate430inter3), .O(gate430inter5));
  nor2  gate959(.a(gate430inter5), .b(gate430inter2), .O(gate430inter6));
  inv1  gate960(.a(G1051), .O(gate430inter7));
  inv1  gate961(.a(G1147), .O(gate430inter8));
  nand2 gate962(.a(gate430inter8), .b(gate430inter7), .O(gate430inter9));
  nand2 gate963(.a(s_59), .b(gate430inter3), .O(gate430inter10));
  nor2  gate964(.a(gate430inter10), .b(gate430inter9), .O(gate430inter11));
  nor2  gate965(.a(gate430inter11), .b(gate430inter6), .O(gate430inter12));
  nand2 gate966(.a(gate430inter12), .b(gate430inter1), .O(G1239));
nand2 gate431( .a(G7), .b(G1150), .O(G1240) );
nand2 gate432( .a(G1054), .b(G1150), .O(G1241) );
nand2 gate433( .a(G8), .b(G1153), .O(G1242) );
nand2 gate434( .a(G1057), .b(G1153), .O(G1243) );
nand2 gate435( .a(G9), .b(G1156), .O(G1244) );
nand2 gate436( .a(G1060), .b(G1156), .O(G1245) );
nand2 gate437( .a(G10), .b(G1159), .O(G1246) );

  xor2  gate2297(.a(G1159), .b(G1063), .O(gate438inter0));
  nand2 gate2298(.a(gate438inter0), .b(s_250), .O(gate438inter1));
  and2  gate2299(.a(G1159), .b(G1063), .O(gate438inter2));
  inv1  gate2300(.a(s_250), .O(gate438inter3));
  inv1  gate2301(.a(s_251), .O(gate438inter4));
  nand2 gate2302(.a(gate438inter4), .b(gate438inter3), .O(gate438inter5));
  nor2  gate2303(.a(gate438inter5), .b(gate438inter2), .O(gate438inter6));
  inv1  gate2304(.a(G1063), .O(gate438inter7));
  inv1  gate2305(.a(G1159), .O(gate438inter8));
  nand2 gate2306(.a(gate438inter8), .b(gate438inter7), .O(gate438inter9));
  nand2 gate2307(.a(s_251), .b(gate438inter3), .O(gate438inter10));
  nor2  gate2308(.a(gate438inter10), .b(gate438inter9), .O(gate438inter11));
  nor2  gate2309(.a(gate438inter11), .b(gate438inter6), .O(gate438inter12));
  nand2 gate2310(.a(gate438inter12), .b(gate438inter1), .O(G1247));
nand2 gate439( .a(G11), .b(G1162), .O(G1248) );

  xor2  gate2619(.a(G1162), .b(G1066), .O(gate440inter0));
  nand2 gate2620(.a(gate440inter0), .b(s_296), .O(gate440inter1));
  and2  gate2621(.a(G1162), .b(G1066), .O(gate440inter2));
  inv1  gate2622(.a(s_296), .O(gate440inter3));
  inv1  gate2623(.a(s_297), .O(gate440inter4));
  nand2 gate2624(.a(gate440inter4), .b(gate440inter3), .O(gate440inter5));
  nor2  gate2625(.a(gate440inter5), .b(gate440inter2), .O(gate440inter6));
  inv1  gate2626(.a(G1066), .O(gate440inter7));
  inv1  gate2627(.a(G1162), .O(gate440inter8));
  nand2 gate2628(.a(gate440inter8), .b(gate440inter7), .O(gate440inter9));
  nand2 gate2629(.a(s_297), .b(gate440inter3), .O(gate440inter10));
  nor2  gate2630(.a(gate440inter10), .b(gate440inter9), .O(gate440inter11));
  nor2  gate2631(.a(gate440inter11), .b(gate440inter6), .O(gate440inter12));
  nand2 gate2632(.a(gate440inter12), .b(gate440inter1), .O(G1249));

  xor2  gate1541(.a(G1165), .b(G12), .O(gate441inter0));
  nand2 gate1542(.a(gate441inter0), .b(s_142), .O(gate441inter1));
  and2  gate1543(.a(G1165), .b(G12), .O(gate441inter2));
  inv1  gate1544(.a(s_142), .O(gate441inter3));
  inv1  gate1545(.a(s_143), .O(gate441inter4));
  nand2 gate1546(.a(gate441inter4), .b(gate441inter3), .O(gate441inter5));
  nor2  gate1547(.a(gate441inter5), .b(gate441inter2), .O(gate441inter6));
  inv1  gate1548(.a(G12), .O(gate441inter7));
  inv1  gate1549(.a(G1165), .O(gate441inter8));
  nand2 gate1550(.a(gate441inter8), .b(gate441inter7), .O(gate441inter9));
  nand2 gate1551(.a(s_143), .b(gate441inter3), .O(gate441inter10));
  nor2  gate1552(.a(gate441inter10), .b(gate441inter9), .O(gate441inter11));
  nor2  gate1553(.a(gate441inter11), .b(gate441inter6), .O(gate441inter12));
  nand2 gate1554(.a(gate441inter12), .b(gate441inter1), .O(G1250));
nand2 gate442( .a(G1069), .b(G1165), .O(G1251) );
nand2 gate443( .a(G13), .b(G1168), .O(G1252) );
nand2 gate444( .a(G1072), .b(G1168), .O(G1253) );

  xor2  gate1429(.a(G1171), .b(G14), .O(gate445inter0));
  nand2 gate1430(.a(gate445inter0), .b(s_126), .O(gate445inter1));
  and2  gate1431(.a(G1171), .b(G14), .O(gate445inter2));
  inv1  gate1432(.a(s_126), .O(gate445inter3));
  inv1  gate1433(.a(s_127), .O(gate445inter4));
  nand2 gate1434(.a(gate445inter4), .b(gate445inter3), .O(gate445inter5));
  nor2  gate1435(.a(gate445inter5), .b(gate445inter2), .O(gate445inter6));
  inv1  gate1436(.a(G14), .O(gate445inter7));
  inv1  gate1437(.a(G1171), .O(gate445inter8));
  nand2 gate1438(.a(gate445inter8), .b(gate445inter7), .O(gate445inter9));
  nand2 gate1439(.a(s_127), .b(gate445inter3), .O(gate445inter10));
  nor2  gate1440(.a(gate445inter10), .b(gate445inter9), .O(gate445inter11));
  nor2  gate1441(.a(gate445inter11), .b(gate445inter6), .O(gate445inter12));
  nand2 gate1442(.a(gate445inter12), .b(gate445inter1), .O(G1254));
nand2 gate446( .a(G1075), .b(G1171), .O(G1255) );

  xor2  gate2059(.a(G1174), .b(G15), .O(gate447inter0));
  nand2 gate2060(.a(gate447inter0), .b(s_216), .O(gate447inter1));
  and2  gate2061(.a(G1174), .b(G15), .O(gate447inter2));
  inv1  gate2062(.a(s_216), .O(gate447inter3));
  inv1  gate2063(.a(s_217), .O(gate447inter4));
  nand2 gate2064(.a(gate447inter4), .b(gate447inter3), .O(gate447inter5));
  nor2  gate2065(.a(gate447inter5), .b(gate447inter2), .O(gate447inter6));
  inv1  gate2066(.a(G15), .O(gate447inter7));
  inv1  gate2067(.a(G1174), .O(gate447inter8));
  nand2 gate2068(.a(gate447inter8), .b(gate447inter7), .O(gate447inter9));
  nand2 gate2069(.a(s_217), .b(gate447inter3), .O(gate447inter10));
  nor2  gate2070(.a(gate447inter10), .b(gate447inter9), .O(gate447inter11));
  nor2  gate2071(.a(gate447inter11), .b(gate447inter6), .O(gate447inter12));
  nand2 gate2072(.a(gate447inter12), .b(gate447inter1), .O(G1256));

  xor2  gate1275(.a(G1174), .b(G1078), .O(gate448inter0));
  nand2 gate1276(.a(gate448inter0), .b(s_104), .O(gate448inter1));
  and2  gate1277(.a(G1174), .b(G1078), .O(gate448inter2));
  inv1  gate1278(.a(s_104), .O(gate448inter3));
  inv1  gate1279(.a(s_105), .O(gate448inter4));
  nand2 gate1280(.a(gate448inter4), .b(gate448inter3), .O(gate448inter5));
  nor2  gate1281(.a(gate448inter5), .b(gate448inter2), .O(gate448inter6));
  inv1  gate1282(.a(G1078), .O(gate448inter7));
  inv1  gate1283(.a(G1174), .O(gate448inter8));
  nand2 gate1284(.a(gate448inter8), .b(gate448inter7), .O(gate448inter9));
  nand2 gate1285(.a(s_105), .b(gate448inter3), .O(gate448inter10));
  nor2  gate1286(.a(gate448inter10), .b(gate448inter9), .O(gate448inter11));
  nor2  gate1287(.a(gate448inter11), .b(gate448inter6), .O(gate448inter12));
  nand2 gate1288(.a(gate448inter12), .b(gate448inter1), .O(G1257));

  xor2  gate1317(.a(G1177), .b(G16), .O(gate449inter0));
  nand2 gate1318(.a(gate449inter0), .b(s_110), .O(gate449inter1));
  and2  gate1319(.a(G1177), .b(G16), .O(gate449inter2));
  inv1  gate1320(.a(s_110), .O(gate449inter3));
  inv1  gate1321(.a(s_111), .O(gate449inter4));
  nand2 gate1322(.a(gate449inter4), .b(gate449inter3), .O(gate449inter5));
  nor2  gate1323(.a(gate449inter5), .b(gate449inter2), .O(gate449inter6));
  inv1  gate1324(.a(G16), .O(gate449inter7));
  inv1  gate1325(.a(G1177), .O(gate449inter8));
  nand2 gate1326(.a(gate449inter8), .b(gate449inter7), .O(gate449inter9));
  nand2 gate1327(.a(s_111), .b(gate449inter3), .O(gate449inter10));
  nor2  gate1328(.a(gate449inter10), .b(gate449inter9), .O(gate449inter11));
  nor2  gate1329(.a(gate449inter11), .b(gate449inter6), .O(gate449inter12));
  nand2 gate1330(.a(gate449inter12), .b(gate449inter1), .O(G1258));
nand2 gate450( .a(G1081), .b(G1177), .O(G1259) );

  xor2  gate1359(.a(G1180), .b(G17), .O(gate451inter0));
  nand2 gate1360(.a(gate451inter0), .b(s_116), .O(gate451inter1));
  and2  gate1361(.a(G1180), .b(G17), .O(gate451inter2));
  inv1  gate1362(.a(s_116), .O(gate451inter3));
  inv1  gate1363(.a(s_117), .O(gate451inter4));
  nand2 gate1364(.a(gate451inter4), .b(gate451inter3), .O(gate451inter5));
  nor2  gate1365(.a(gate451inter5), .b(gate451inter2), .O(gate451inter6));
  inv1  gate1366(.a(G17), .O(gate451inter7));
  inv1  gate1367(.a(G1180), .O(gate451inter8));
  nand2 gate1368(.a(gate451inter8), .b(gate451inter7), .O(gate451inter9));
  nand2 gate1369(.a(s_117), .b(gate451inter3), .O(gate451inter10));
  nor2  gate1370(.a(gate451inter10), .b(gate451inter9), .O(gate451inter11));
  nor2  gate1371(.a(gate451inter11), .b(gate451inter6), .O(gate451inter12));
  nand2 gate1372(.a(gate451inter12), .b(gate451inter1), .O(G1260));

  xor2  gate2381(.a(G1180), .b(G1084), .O(gate452inter0));
  nand2 gate2382(.a(gate452inter0), .b(s_262), .O(gate452inter1));
  and2  gate2383(.a(G1180), .b(G1084), .O(gate452inter2));
  inv1  gate2384(.a(s_262), .O(gate452inter3));
  inv1  gate2385(.a(s_263), .O(gate452inter4));
  nand2 gate2386(.a(gate452inter4), .b(gate452inter3), .O(gate452inter5));
  nor2  gate2387(.a(gate452inter5), .b(gate452inter2), .O(gate452inter6));
  inv1  gate2388(.a(G1084), .O(gate452inter7));
  inv1  gate2389(.a(G1180), .O(gate452inter8));
  nand2 gate2390(.a(gate452inter8), .b(gate452inter7), .O(gate452inter9));
  nand2 gate2391(.a(s_263), .b(gate452inter3), .O(gate452inter10));
  nor2  gate2392(.a(gate452inter10), .b(gate452inter9), .O(gate452inter11));
  nor2  gate2393(.a(gate452inter11), .b(gate452inter6), .O(gate452inter12));
  nand2 gate2394(.a(gate452inter12), .b(gate452inter1), .O(G1261));
nand2 gate453( .a(G18), .b(G1183), .O(G1262) );
nand2 gate454( .a(G1087), .b(G1183), .O(G1263) );
nand2 gate455( .a(G19), .b(G1186), .O(G1264) );

  xor2  gate1989(.a(G1186), .b(G1090), .O(gate456inter0));
  nand2 gate1990(.a(gate456inter0), .b(s_206), .O(gate456inter1));
  and2  gate1991(.a(G1186), .b(G1090), .O(gate456inter2));
  inv1  gate1992(.a(s_206), .O(gate456inter3));
  inv1  gate1993(.a(s_207), .O(gate456inter4));
  nand2 gate1994(.a(gate456inter4), .b(gate456inter3), .O(gate456inter5));
  nor2  gate1995(.a(gate456inter5), .b(gate456inter2), .O(gate456inter6));
  inv1  gate1996(.a(G1090), .O(gate456inter7));
  inv1  gate1997(.a(G1186), .O(gate456inter8));
  nand2 gate1998(.a(gate456inter8), .b(gate456inter7), .O(gate456inter9));
  nand2 gate1999(.a(s_207), .b(gate456inter3), .O(gate456inter10));
  nor2  gate2000(.a(gate456inter10), .b(gate456inter9), .O(gate456inter11));
  nor2  gate2001(.a(gate456inter11), .b(gate456inter6), .O(gate456inter12));
  nand2 gate2002(.a(gate456inter12), .b(gate456inter1), .O(G1265));

  xor2  gate1527(.a(G1189), .b(G20), .O(gate457inter0));
  nand2 gate1528(.a(gate457inter0), .b(s_140), .O(gate457inter1));
  and2  gate1529(.a(G1189), .b(G20), .O(gate457inter2));
  inv1  gate1530(.a(s_140), .O(gate457inter3));
  inv1  gate1531(.a(s_141), .O(gate457inter4));
  nand2 gate1532(.a(gate457inter4), .b(gate457inter3), .O(gate457inter5));
  nor2  gate1533(.a(gate457inter5), .b(gate457inter2), .O(gate457inter6));
  inv1  gate1534(.a(G20), .O(gate457inter7));
  inv1  gate1535(.a(G1189), .O(gate457inter8));
  nand2 gate1536(.a(gate457inter8), .b(gate457inter7), .O(gate457inter9));
  nand2 gate1537(.a(s_141), .b(gate457inter3), .O(gate457inter10));
  nor2  gate1538(.a(gate457inter10), .b(gate457inter9), .O(gate457inter11));
  nor2  gate1539(.a(gate457inter11), .b(gate457inter6), .O(gate457inter12));
  nand2 gate1540(.a(gate457inter12), .b(gate457inter1), .O(G1266));
nand2 gate458( .a(G1093), .b(G1189), .O(G1267) );
nand2 gate459( .a(G21), .b(G1192), .O(G1268) );

  xor2  gate1135(.a(G1192), .b(G1096), .O(gate460inter0));
  nand2 gate1136(.a(gate460inter0), .b(s_84), .O(gate460inter1));
  and2  gate1137(.a(G1192), .b(G1096), .O(gate460inter2));
  inv1  gate1138(.a(s_84), .O(gate460inter3));
  inv1  gate1139(.a(s_85), .O(gate460inter4));
  nand2 gate1140(.a(gate460inter4), .b(gate460inter3), .O(gate460inter5));
  nor2  gate1141(.a(gate460inter5), .b(gate460inter2), .O(gate460inter6));
  inv1  gate1142(.a(G1096), .O(gate460inter7));
  inv1  gate1143(.a(G1192), .O(gate460inter8));
  nand2 gate1144(.a(gate460inter8), .b(gate460inter7), .O(gate460inter9));
  nand2 gate1145(.a(s_85), .b(gate460inter3), .O(gate460inter10));
  nor2  gate1146(.a(gate460inter10), .b(gate460inter9), .O(gate460inter11));
  nor2  gate1147(.a(gate460inter11), .b(gate460inter6), .O(gate460inter12));
  nand2 gate1148(.a(gate460inter12), .b(gate460inter1), .O(G1269));

  xor2  gate925(.a(G1195), .b(G22), .O(gate461inter0));
  nand2 gate926(.a(gate461inter0), .b(s_54), .O(gate461inter1));
  and2  gate927(.a(G1195), .b(G22), .O(gate461inter2));
  inv1  gate928(.a(s_54), .O(gate461inter3));
  inv1  gate929(.a(s_55), .O(gate461inter4));
  nand2 gate930(.a(gate461inter4), .b(gate461inter3), .O(gate461inter5));
  nor2  gate931(.a(gate461inter5), .b(gate461inter2), .O(gate461inter6));
  inv1  gate932(.a(G22), .O(gate461inter7));
  inv1  gate933(.a(G1195), .O(gate461inter8));
  nand2 gate934(.a(gate461inter8), .b(gate461inter7), .O(gate461inter9));
  nand2 gate935(.a(s_55), .b(gate461inter3), .O(gate461inter10));
  nor2  gate936(.a(gate461inter10), .b(gate461inter9), .O(gate461inter11));
  nor2  gate937(.a(gate461inter11), .b(gate461inter6), .O(gate461inter12));
  nand2 gate938(.a(gate461inter12), .b(gate461inter1), .O(G1270));
nand2 gate462( .a(G1099), .b(G1195), .O(G1271) );

  xor2  gate1639(.a(G1198), .b(G23), .O(gate463inter0));
  nand2 gate1640(.a(gate463inter0), .b(s_156), .O(gate463inter1));
  and2  gate1641(.a(G1198), .b(G23), .O(gate463inter2));
  inv1  gate1642(.a(s_156), .O(gate463inter3));
  inv1  gate1643(.a(s_157), .O(gate463inter4));
  nand2 gate1644(.a(gate463inter4), .b(gate463inter3), .O(gate463inter5));
  nor2  gate1645(.a(gate463inter5), .b(gate463inter2), .O(gate463inter6));
  inv1  gate1646(.a(G23), .O(gate463inter7));
  inv1  gate1647(.a(G1198), .O(gate463inter8));
  nand2 gate1648(.a(gate463inter8), .b(gate463inter7), .O(gate463inter9));
  nand2 gate1649(.a(s_157), .b(gate463inter3), .O(gate463inter10));
  nor2  gate1650(.a(gate463inter10), .b(gate463inter9), .O(gate463inter11));
  nor2  gate1651(.a(gate463inter11), .b(gate463inter6), .O(gate463inter12));
  nand2 gate1652(.a(gate463inter12), .b(gate463inter1), .O(G1272));

  xor2  gate2535(.a(G1198), .b(G1102), .O(gate464inter0));
  nand2 gate2536(.a(gate464inter0), .b(s_284), .O(gate464inter1));
  and2  gate2537(.a(G1198), .b(G1102), .O(gate464inter2));
  inv1  gate2538(.a(s_284), .O(gate464inter3));
  inv1  gate2539(.a(s_285), .O(gate464inter4));
  nand2 gate2540(.a(gate464inter4), .b(gate464inter3), .O(gate464inter5));
  nor2  gate2541(.a(gate464inter5), .b(gate464inter2), .O(gate464inter6));
  inv1  gate2542(.a(G1102), .O(gate464inter7));
  inv1  gate2543(.a(G1198), .O(gate464inter8));
  nand2 gate2544(.a(gate464inter8), .b(gate464inter7), .O(gate464inter9));
  nand2 gate2545(.a(s_285), .b(gate464inter3), .O(gate464inter10));
  nor2  gate2546(.a(gate464inter10), .b(gate464inter9), .O(gate464inter11));
  nor2  gate2547(.a(gate464inter11), .b(gate464inter6), .O(gate464inter12));
  nand2 gate2548(.a(gate464inter12), .b(gate464inter1), .O(G1273));
nand2 gate465( .a(G24), .b(G1201), .O(G1274) );

  xor2  gate2633(.a(G1201), .b(G1105), .O(gate466inter0));
  nand2 gate2634(.a(gate466inter0), .b(s_298), .O(gate466inter1));
  and2  gate2635(.a(G1201), .b(G1105), .O(gate466inter2));
  inv1  gate2636(.a(s_298), .O(gate466inter3));
  inv1  gate2637(.a(s_299), .O(gate466inter4));
  nand2 gate2638(.a(gate466inter4), .b(gate466inter3), .O(gate466inter5));
  nor2  gate2639(.a(gate466inter5), .b(gate466inter2), .O(gate466inter6));
  inv1  gate2640(.a(G1105), .O(gate466inter7));
  inv1  gate2641(.a(G1201), .O(gate466inter8));
  nand2 gate2642(.a(gate466inter8), .b(gate466inter7), .O(gate466inter9));
  nand2 gate2643(.a(s_299), .b(gate466inter3), .O(gate466inter10));
  nor2  gate2644(.a(gate466inter10), .b(gate466inter9), .O(gate466inter11));
  nor2  gate2645(.a(gate466inter11), .b(gate466inter6), .O(gate466inter12));
  nand2 gate2646(.a(gate466inter12), .b(gate466inter1), .O(G1275));

  xor2  gate1779(.a(G1204), .b(G25), .O(gate467inter0));
  nand2 gate1780(.a(gate467inter0), .b(s_176), .O(gate467inter1));
  and2  gate1781(.a(G1204), .b(G25), .O(gate467inter2));
  inv1  gate1782(.a(s_176), .O(gate467inter3));
  inv1  gate1783(.a(s_177), .O(gate467inter4));
  nand2 gate1784(.a(gate467inter4), .b(gate467inter3), .O(gate467inter5));
  nor2  gate1785(.a(gate467inter5), .b(gate467inter2), .O(gate467inter6));
  inv1  gate1786(.a(G25), .O(gate467inter7));
  inv1  gate1787(.a(G1204), .O(gate467inter8));
  nand2 gate1788(.a(gate467inter8), .b(gate467inter7), .O(gate467inter9));
  nand2 gate1789(.a(s_177), .b(gate467inter3), .O(gate467inter10));
  nor2  gate1790(.a(gate467inter10), .b(gate467inter9), .O(gate467inter11));
  nor2  gate1791(.a(gate467inter11), .b(gate467inter6), .O(gate467inter12));
  nand2 gate1792(.a(gate467inter12), .b(gate467inter1), .O(G1276));
nand2 gate468( .a(G1108), .b(G1204), .O(G1277) );
nand2 gate469( .a(G26), .b(G1207), .O(G1278) );
nand2 gate470( .a(G1111), .b(G1207), .O(G1279) );
nand2 gate471( .a(G27), .b(G1210), .O(G1280) );

  xor2  gate2073(.a(G1210), .b(G1114), .O(gate472inter0));
  nand2 gate2074(.a(gate472inter0), .b(s_218), .O(gate472inter1));
  and2  gate2075(.a(G1210), .b(G1114), .O(gate472inter2));
  inv1  gate2076(.a(s_218), .O(gate472inter3));
  inv1  gate2077(.a(s_219), .O(gate472inter4));
  nand2 gate2078(.a(gate472inter4), .b(gate472inter3), .O(gate472inter5));
  nor2  gate2079(.a(gate472inter5), .b(gate472inter2), .O(gate472inter6));
  inv1  gate2080(.a(G1114), .O(gate472inter7));
  inv1  gate2081(.a(G1210), .O(gate472inter8));
  nand2 gate2082(.a(gate472inter8), .b(gate472inter7), .O(gate472inter9));
  nand2 gate2083(.a(s_219), .b(gate472inter3), .O(gate472inter10));
  nor2  gate2084(.a(gate472inter10), .b(gate472inter9), .O(gate472inter11));
  nor2  gate2085(.a(gate472inter11), .b(gate472inter6), .O(gate472inter12));
  nand2 gate2086(.a(gate472inter12), .b(gate472inter1), .O(G1281));

  xor2  gate2479(.a(G1213), .b(G28), .O(gate473inter0));
  nand2 gate2480(.a(gate473inter0), .b(s_276), .O(gate473inter1));
  and2  gate2481(.a(G1213), .b(G28), .O(gate473inter2));
  inv1  gate2482(.a(s_276), .O(gate473inter3));
  inv1  gate2483(.a(s_277), .O(gate473inter4));
  nand2 gate2484(.a(gate473inter4), .b(gate473inter3), .O(gate473inter5));
  nor2  gate2485(.a(gate473inter5), .b(gate473inter2), .O(gate473inter6));
  inv1  gate2486(.a(G28), .O(gate473inter7));
  inv1  gate2487(.a(G1213), .O(gate473inter8));
  nand2 gate2488(.a(gate473inter8), .b(gate473inter7), .O(gate473inter9));
  nand2 gate2489(.a(s_277), .b(gate473inter3), .O(gate473inter10));
  nor2  gate2490(.a(gate473inter10), .b(gate473inter9), .O(gate473inter11));
  nor2  gate2491(.a(gate473inter11), .b(gate473inter6), .O(gate473inter12));
  nand2 gate2492(.a(gate473inter12), .b(gate473inter1), .O(G1282));

  xor2  gate1667(.a(G1213), .b(G1117), .O(gate474inter0));
  nand2 gate1668(.a(gate474inter0), .b(s_160), .O(gate474inter1));
  and2  gate1669(.a(G1213), .b(G1117), .O(gate474inter2));
  inv1  gate1670(.a(s_160), .O(gate474inter3));
  inv1  gate1671(.a(s_161), .O(gate474inter4));
  nand2 gate1672(.a(gate474inter4), .b(gate474inter3), .O(gate474inter5));
  nor2  gate1673(.a(gate474inter5), .b(gate474inter2), .O(gate474inter6));
  inv1  gate1674(.a(G1117), .O(gate474inter7));
  inv1  gate1675(.a(G1213), .O(gate474inter8));
  nand2 gate1676(.a(gate474inter8), .b(gate474inter7), .O(gate474inter9));
  nand2 gate1677(.a(s_161), .b(gate474inter3), .O(gate474inter10));
  nor2  gate1678(.a(gate474inter10), .b(gate474inter9), .O(gate474inter11));
  nor2  gate1679(.a(gate474inter11), .b(gate474inter6), .O(gate474inter12));
  nand2 gate1680(.a(gate474inter12), .b(gate474inter1), .O(G1283));
nand2 gate475( .a(G29), .b(G1216), .O(G1284) );

  xor2  gate1555(.a(G1216), .b(G1120), .O(gate476inter0));
  nand2 gate1556(.a(gate476inter0), .b(s_144), .O(gate476inter1));
  and2  gate1557(.a(G1216), .b(G1120), .O(gate476inter2));
  inv1  gate1558(.a(s_144), .O(gate476inter3));
  inv1  gate1559(.a(s_145), .O(gate476inter4));
  nand2 gate1560(.a(gate476inter4), .b(gate476inter3), .O(gate476inter5));
  nor2  gate1561(.a(gate476inter5), .b(gate476inter2), .O(gate476inter6));
  inv1  gate1562(.a(G1120), .O(gate476inter7));
  inv1  gate1563(.a(G1216), .O(gate476inter8));
  nand2 gate1564(.a(gate476inter8), .b(gate476inter7), .O(gate476inter9));
  nand2 gate1565(.a(s_145), .b(gate476inter3), .O(gate476inter10));
  nor2  gate1566(.a(gate476inter10), .b(gate476inter9), .O(gate476inter11));
  nor2  gate1567(.a(gate476inter11), .b(gate476inter6), .O(gate476inter12));
  nand2 gate1568(.a(gate476inter12), .b(gate476inter1), .O(G1285));

  xor2  gate1611(.a(G1219), .b(G30), .O(gate477inter0));
  nand2 gate1612(.a(gate477inter0), .b(s_152), .O(gate477inter1));
  and2  gate1613(.a(G1219), .b(G30), .O(gate477inter2));
  inv1  gate1614(.a(s_152), .O(gate477inter3));
  inv1  gate1615(.a(s_153), .O(gate477inter4));
  nand2 gate1616(.a(gate477inter4), .b(gate477inter3), .O(gate477inter5));
  nor2  gate1617(.a(gate477inter5), .b(gate477inter2), .O(gate477inter6));
  inv1  gate1618(.a(G30), .O(gate477inter7));
  inv1  gate1619(.a(G1219), .O(gate477inter8));
  nand2 gate1620(.a(gate477inter8), .b(gate477inter7), .O(gate477inter9));
  nand2 gate1621(.a(s_153), .b(gate477inter3), .O(gate477inter10));
  nor2  gate1622(.a(gate477inter10), .b(gate477inter9), .O(gate477inter11));
  nor2  gate1623(.a(gate477inter11), .b(gate477inter6), .O(gate477inter12));
  nand2 gate1624(.a(gate477inter12), .b(gate477inter1), .O(G1286));

  xor2  gate911(.a(G1219), .b(G1123), .O(gate478inter0));
  nand2 gate912(.a(gate478inter0), .b(s_52), .O(gate478inter1));
  and2  gate913(.a(G1219), .b(G1123), .O(gate478inter2));
  inv1  gate914(.a(s_52), .O(gate478inter3));
  inv1  gate915(.a(s_53), .O(gate478inter4));
  nand2 gate916(.a(gate478inter4), .b(gate478inter3), .O(gate478inter5));
  nor2  gate917(.a(gate478inter5), .b(gate478inter2), .O(gate478inter6));
  inv1  gate918(.a(G1123), .O(gate478inter7));
  inv1  gate919(.a(G1219), .O(gate478inter8));
  nand2 gate920(.a(gate478inter8), .b(gate478inter7), .O(gate478inter9));
  nand2 gate921(.a(s_53), .b(gate478inter3), .O(gate478inter10));
  nor2  gate922(.a(gate478inter10), .b(gate478inter9), .O(gate478inter11));
  nor2  gate923(.a(gate478inter11), .b(gate478inter6), .O(gate478inter12));
  nand2 gate924(.a(gate478inter12), .b(gate478inter1), .O(G1287));
nand2 gate479( .a(G31), .b(G1222), .O(G1288) );

  xor2  gate1695(.a(G1222), .b(G1126), .O(gate480inter0));
  nand2 gate1696(.a(gate480inter0), .b(s_164), .O(gate480inter1));
  and2  gate1697(.a(G1222), .b(G1126), .O(gate480inter2));
  inv1  gate1698(.a(s_164), .O(gate480inter3));
  inv1  gate1699(.a(s_165), .O(gate480inter4));
  nand2 gate1700(.a(gate480inter4), .b(gate480inter3), .O(gate480inter5));
  nor2  gate1701(.a(gate480inter5), .b(gate480inter2), .O(gate480inter6));
  inv1  gate1702(.a(G1126), .O(gate480inter7));
  inv1  gate1703(.a(G1222), .O(gate480inter8));
  nand2 gate1704(.a(gate480inter8), .b(gate480inter7), .O(gate480inter9));
  nand2 gate1705(.a(s_165), .b(gate480inter3), .O(gate480inter10));
  nor2  gate1706(.a(gate480inter10), .b(gate480inter9), .O(gate480inter11));
  nor2  gate1707(.a(gate480inter11), .b(gate480inter6), .O(gate480inter12));
  nand2 gate1708(.a(gate480inter12), .b(gate480inter1), .O(G1289));
nand2 gate481( .a(G32), .b(G1225), .O(G1290) );

  xor2  gate1597(.a(G1225), .b(G1129), .O(gate482inter0));
  nand2 gate1598(.a(gate482inter0), .b(s_150), .O(gate482inter1));
  and2  gate1599(.a(G1225), .b(G1129), .O(gate482inter2));
  inv1  gate1600(.a(s_150), .O(gate482inter3));
  inv1  gate1601(.a(s_151), .O(gate482inter4));
  nand2 gate1602(.a(gate482inter4), .b(gate482inter3), .O(gate482inter5));
  nor2  gate1603(.a(gate482inter5), .b(gate482inter2), .O(gate482inter6));
  inv1  gate1604(.a(G1129), .O(gate482inter7));
  inv1  gate1605(.a(G1225), .O(gate482inter8));
  nand2 gate1606(.a(gate482inter8), .b(gate482inter7), .O(gate482inter9));
  nand2 gate1607(.a(s_151), .b(gate482inter3), .O(gate482inter10));
  nor2  gate1608(.a(gate482inter10), .b(gate482inter9), .O(gate482inter11));
  nor2  gate1609(.a(gate482inter11), .b(gate482inter6), .O(gate482inter12));
  nand2 gate1610(.a(gate482inter12), .b(gate482inter1), .O(G1291));
nand2 gate483( .a(G1228), .b(G1229), .O(G1292) );

  xor2  gate1653(.a(G1231), .b(G1230), .O(gate484inter0));
  nand2 gate1654(.a(gate484inter0), .b(s_158), .O(gate484inter1));
  and2  gate1655(.a(G1231), .b(G1230), .O(gate484inter2));
  inv1  gate1656(.a(s_158), .O(gate484inter3));
  inv1  gate1657(.a(s_159), .O(gate484inter4));
  nand2 gate1658(.a(gate484inter4), .b(gate484inter3), .O(gate484inter5));
  nor2  gate1659(.a(gate484inter5), .b(gate484inter2), .O(gate484inter6));
  inv1  gate1660(.a(G1230), .O(gate484inter7));
  inv1  gate1661(.a(G1231), .O(gate484inter8));
  nand2 gate1662(.a(gate484inter8), .b(gate484inter7), .O(gate484inter9));
  nand2 gate1663(.a(s_159), .b(gate484inter3), .O(gate484inter10));
  nor2  gate1664(.a(gate484inter10), .b(gate484inter9), .O(gate484inter11));
  nor2  gate1665(.a(gate484inter11), .b(gate484inter6), .O(gate484inter12));
  nand2 gate1666(.a(gate484inter12), .b(gate484inter1), .O(G1293));
nand2 gate485( .a(G1232), .b(G1233), .O(G1294) );

  xor2  gate2157(.a(G1235), .b(G1234), .O(gate486inter0));
  nand2 gate2158(.a(gate486inter0), .b(s_230), .O(gate486inter1));
  and2  gate2159(.a(G1235), .b(G1234), .O(gate486inter2));
  inv1  gate2160(.a(s_230), .O(gate486inter3));
  inv1  gate2161(.a(s_231), .O(gate486inter4));
  nand2 gate2162(.a(gate486inter4), .b(gate486inter3), .O(gate486inter5));
  nor2  gate2163(.a(gate486inter5), .b(gate486inter2), .O(gate486inter6));
  inv1  gate2164(.a(G1234), .O(gate486inter7));
  inv1  gate2165(.a(G1235), .O(gate486inter8));
  nand2 gate2166(.a(gate486inter8), .b(gate486inter7), .O(gate486inter9));
  nand2 gate2167(.a(s_231), .b(gate486inter3), .O(gate486inter10));
  nor2  gate2168(.a(gate486inter10), .b(gate486inter9), .O(gate486inter11));
  nor2  gate2169(.a(gate486inter11), .b(gate486inter6), .O(gate486inter12));
  nand2 gate2170(.a(gate486inter12), .b(gate486inter1), .O(G1295));
nand2 gate487( .a(G1236), .b(G1237), .O(G1296) );
nand2 gate488( .a(G1238), .b(G1239), .O(G1297) );

  xor2  gate645(.a(G1241), .b(G1240), .O(gate489inter0));
  nand2 gate646(.a(gate489inter0), .b(s_14), .O(gate489inter1));
  and2  gate647(.a(G1241), .b(G1240), .O(gate489inter2));
  inv1  gate648(.a(s_14), .O(gate489inter3));
  inv1  gate649(.a(s_15), .O(gate489inter4));
  nand2 gate650(.a(gate489inter4), .b(gate489inter3), .O(gate489inter5));
  nor2  gate651(.a(gate489inter5), .b(gate489inter2), .O(gate489inter6));
  inv1  gate652(.a(G1240), .O(gate489inter7));
  inv1  gate653(.a(G1241), .O(gate489inter8));
  nand2 gate654(.a(gate489inter8), .b(gate489inter7), .O(gate489inter9));
  nand2 gate655(.a(s_15), .b(gate489inter3), .O(gate489inter10));
  nor2  gate656(.a(gate489inter10), .b(gate489inter9), .O(gate489inter11));
  nor2  gate657(.a(gate489inter11), .b(gate489inter6), .O(gate489inter12));
  nand2 gate658(.a(gate489inter12), .b(gate489inter1), .O(G1298));
nand2 gate490( .a(G1242), .b(G1243), .O(G1299) );

  xor2  gate2325(.a(G1245), .b(G1244), .O(gate491inter0));
  nand2 gate2326(.a(gate491inter0), .b(s_254), .O(gate491inter1));
  and2  gate2327(.a(G1245), .b(G1244), .O(gate491inter2));
  inv1  gate2328(.a(s_254), .O(gate491inter3));
  inv1  gate2329(.a(s_255), .O(gate491inter4));
  nand2 gate2330(.a(gate491inter4), .b(gate491inter3), .O(gate491inter5));
  nor2  gate2331(.a(gate491inter5), .b(gate491inter2), .O(gate491inter6));
  inv1  gate2332(.a(G1244), .O(gate491inter7));
  inv1  gate2333(.a(G1245), .O(gate491inter8));
  nand2 gate2334(.a(gate491inter8), .b(gate491inter7), .O(gate491inter9));
  nand2 gate2335(.a(s_255), .b(gate491inter3), .O(gate491inter10));
  nor2  gate2336(.a(gate491inter10), .b(gate491inter9), .O(gate491inter11));
  nor2  gate2337(.a(gate491inter11), .b(gate491inter6), .O(gate491inter12));
  nand2 gate2338(.a(gate491inter12), .b(gate491inter1), .O(G1300));
nand2 gate492( .a(G1246), .b(G1247), .O(G1301) );
nand2 gate493( .a(G1248), .b(G1249), .O(G1302) );

  xor2  gate1093(.a(G1251), .b(G1250), .O(gate494inter0));
  nand2 gate1094(.a(gate494inter0), .b(s_78), .O(gate494inter1));
  and2  gate1095(.a(G1251), .b(G1250), .O(gate494inter2));
  inv1  gate1096(.a(s_78), .O(gate494inter3));
  inv1  gate1097(.a(s_79), .O(gate494inter4));
  nand2 gate1098(.a(gate494inter4), .b(gate494inter3), .O(gate494inter5));
  nor2  gate1099(.a(gate494inter5), .b(gate494inter2), .O(gate494inter6));
  inv1  gate1100(.a(G1250), .O(gate494inter7));
  inv1  gate1101(.a(G1251), .O(gate494inter8));
  nand2 gate1102(.a(gate494inter8), .b(gate494inter7), .O(gate494inter9));
  nand2 gate1103(.a(s_79), .b(gate494inter3), .O(gate494inter10));
  nor2  gate1104(.a(gate494inter10), .b(gate494inter9), .O(gate494inter11));
  nor2  gate1105(.a(gate494inter11), .b(gate494inter6), .O(gate494inter12));
  nand2 gate1106(.a(gate494inter12), .b(gate494inter1), .O(G1303));

  xor2  gate2647(.a(G1253), .b(G1252), .O(gate495inter0));
  nand2 gate2648(.a(gate495inter0), .b(s_300), .O(gate495inter1));
  and2  gate2649(.a(G1253), .b(G1252), .O(gate495inter2));
  inv1  gate2650(.a(s_300), .O(gate495inter3));
  inv1  gate2651(.a(s_301), .O(gate495inter4));
  nand2 gate2652(.a(gate495inter4), .b(gate495inter3), .O(gate495inter5));
  nor2  gate2653(.a(gate495inter5), .b(gate495inter2), .O(gate495inter6));
  inv1  gate2654(.a(G1252), .O(gate495inter7));
  inv1  gate2655(.a(G1253), .O(gate495inter8));
  nand2 gate2656(.a(gate495inter8), .b(gate495inter7), .O(gate495inter9));
  nand2 gate2657(.a(s_301), .b(gate495inter3), .O(gate495inter10));
  nor2  gate2658(.a(gate495inter10), .b(gate495inter9), .O(gate495inter11));
  nor2  gate2659(.a(gate495inter11), .b(gate495inter6), .O(gate495inter12));
  nand2 gate2660(.a(gate495inter12), .b(gate495inter1), .O(G1304));
nand2 gate496( .a(G1254), .b(G1255), .O(G1305) );
nand2 gate497( .a(G1256), .b(G1257), .O(G1306) );

  xor2  gate1205(.a(G1259), .b(G1258), .O(gate498inter0));
  nand2 gate1206(.a(gate498inter0), .b(s_94), .O(gate498inter1));
  and2  gate1207(.a(G1259), .b(G1258), .O(gate498inter2));
  inv1  gate1208(.a(s_94), .O(gate498inter3));
  inv1  gate1209(.a(s_95), .O(gate498inter4));
  nand2 gate1210(.a(gate498inter4), .b(gate498inter3), .O(gate498inter5));
  nor2  gate1211(.a(gate498inter5), .b(gate498inter2), .O(gate498inter6));
  inv1  gate1212(.a(G1258), .O(gate498inter7));
  inv1  gate1213(.a(G1259), .O(gate498inter8));
  nand2 gate1214(.a(gate498inter8), .b(gate498inter7), .O(gate498inter9));
  nand2 gate1215(.a(s_95), .b(gate498inter3), .O(gate498inter10));
  nor2  gate1216(.a(gate498inter10), .b(gate498inter9), .O(gate498inter11));
  nor2  gate1217(.a(gate498inter11), .b(gate498inter6), .O(gate498inter12));
  nand2 gate1218(.a(gate498inter12), .b(gate498inter1), .O(G1307));

  xor2  gate1331(.a(G1261), .b(G1260), .O(gate499inter0));
  nand2 gate1332(.a(gate499inter0), .b(s_112), .O(gate499inter1));
  and2  gate1333(.a(G1261), .b(G1260), .O(gate499inter2));
  inv1  gate1334(.a(s_112), .O(gate499inter3));
  inv1  gate1335(.a(s_113), .O(gate499inter4));
  nand2 gate1336(.a(gate499inter4), .b(gate499inter3), .O(gate499inter5));
  nor2  gate1337(.a(gate499inter5), .b(gate499inter2), .O(gate499inter6));
  inv1  gate1338(.a(G1260), .O(gate499inter7));
  inv1  gate1339(.a(G1261), .O(gate499inter8));
  nand2 gate1340(.a(gate499inter8), .b(gate499inter7), .O(gate499inter9));
  nand2 gate1341(.a(s_113), .b(gate499inter3), .O(gate499inter10));
  nor2  gate1342(.a(gate499inter10), .b(gate499inter9), .O(gate499inter11));
  nor2  gate1343(.a(gate499inter11), .b(gate499inter6), .O(gate499inter12));
  nand2 gate1344(.a(gate499inter12), .b(gate499inter1), .O(G1308));
nand2 gate500( .a(G1262), .b(G1263), .O(G1309) );

  xor2  gate1177(.a(G1265), .b(G1264), .O(gate501inter0));
  nand2 gate1178(.a(gate501inter0), .b(s_90), .O(gate501inter1));
  and2  gate1179(.a(G1265), .b(G1264), .O(gate501inter2));
  inv1  gate1180(.a(s_90), .O(gate501inter3));
  inv1  gate1181(.a(s_91), .O(gate501inter4));
  nand2 gate1182(.a(gate501inter4), .b(gate501inter3), .O(gate501inter5));
  nor2  gate1183(.a(gate501inter5), .b(gate501inter2), .O(gate501inter6));
  inv1  gate1184(.a(G1264), .O(gate501inter7));
  inv1  gate1185(.a(G1265), .O(gate501inter8));
  nand2 gate1186(.a(gate501inter8), .b(gate501inter7), .O(gate501inter9));
  nand2 gate1187(.a(s_91), .b(gate501inter3), .O(gate501inter10));
  nor2  gate1188(.a(gate501inter10), .b(gate501inter9), .O(gate501inter11));
  nor2  gate1189(.a(gate501inter11), .b(gate501inter6), .O(gate501inter12));
  nand2 gate1190(.a(gate501inter12), .b(gate501inter1), .O(G1310));

  xor2  gate2087(.a(G1267), .b(G1266), .O(gate502inter0));
  nand2 gate2088(.a(gate502inter0), .b(s_220), .O(gate502inter1));
  and2  gate2089(.a(G1267), .b(G1266), .O(gate502inter2));
  inv1  gate2090(.a(s_220), .O(gate502inter3));
  inv1  gate2091(.a(s_221), .O(gate502inter4));
  nand2 gate2092(.a(gate502inter4), .b(gate502inter3), .O(gate502inter5));
  nor2  gate2093(.a(gate502inter5), .b(gate502inter2), .O(gate502inter6));
  inv1  gate2094(.a(G1266), .O(gate502inter7));
  inv1  gate2095(.a(G1267), .O(gate502inter8));
  nand2 gate2096(.a(gate502inter8), .b(gate502inter7), .O(gate502inter9));
  nand2 gate2097(.a(s_221), .b(gate502inter3), .O(gate502inter10));
  nor2  gate2098(.a(gate502inter10), .b(gate502inter9), .O(gate502inter11));
  nor2  gate2099(.a(gate502inter11), .b(gate502inter6), .O(gate502inter12));
  nand2 gate2100(.a(gate502inter12), .b(gate502inter1), .O(G1311));

  xor2  gate1709(.a(G1269), .b(G1268), .O(gate503inter0));
  nand2 gate1710(.a(gate503inter0), .b(s_166), .O(gate503inter1));
  and2  gate1711(.a(G1269), .b(G1268), .O(gate503inter2));
  inv1  gate1712(.a(s_166), .O(gate503inter3));
  inv1  gate1713(.a(s_167), .O(gate503inter4));
  nand2 gate1714(.a(gate503inter4), .b(gate503inter3), .O(gate503inter5));
  nor2  gate1715(.a(gate503inter5), .b(gate503inter2), .O(gate503inter6));
  inv1  gate1716(.a(G1268), .O(gate503inter7));
  inv1  gate1717(.a(G1269), .O(gate503inter8));
  nand2 gate1718(.a(gate503inter8), .b(gate503inter7), .O(gate503inter9));
  nand2 gate1719(.a(s_167), .b(gate503inter3), .O(gate503inter10));
  nor2  gate1720(.a(gate503inter10), .b(gate503inter9), .O(gate503inter11));
  nor2  gate1721(.a(gate503inter11), .b(gate503inter6), .O(gate503inter12));
  nand2 gate1722(.a(gate503inter12), .b(gate503inter1), .O(G1312));
nand2 gate504( .a(G1270), .b(G1271), .O(G1313) );
nand2 gate505( .a(G1272), .b(G1273), .O(G1314) );
nand2 gate506( .a(G1274), .b(G1275), .O(G1315) );
nand2 gate507( .a(G1276), .b(G1277), .O(G1316) );
nand2 gate508( .a(G1278), .b(G1279), .O(G1317) );

  xor2  gate967(.a(G1281), .b(G1280), .O(gate509inter0));
  nand2 gate968(.a(gate509inter0), .b(s_60), .O(gate509inter1));
  and2  gate969(.a(G1281), .b(G1280), .O(gate509inter2));
  inv1  gate970(.a(s_60), .O(gate509inter3));
  inv1  gate971(.a(s_61), .O(gate509inter4));
  nand2 gate972(.a(gate509inter4), .b(gate509inter3), .O(gate509inter5));
  nor2  gate973(.a(gate509inter5), .b(gate509inter2), .O(gate509inter6));
  inv1  gate974(.a(G1280), .O(gate509inter7));
  inv1  gate975(.a(G1281), .O(gate509inter8));
  nand2 gate976(.a(gate509inter8), .b(gate509inter7), .O(gate509inter9));
  nand2 gate977(.a(s_61), .b(gate509inter3), .O(gate509inter10));
  nor2  gate978(.a(gate509inter10), .b(gate509inter9), .O(gate509inter11));
  nor2  gate979(.a(gate509inter11), .b(gate509inter6), .O(gate509inter12));
  nand2 gate980(.a(gate509inter12), .b(gate509inter1), .O(G1318));
nand2 gate510( .a(G1282), .b(G1283), .O(G1319) );

  xor2  gate1499(.a(G1285), .b(G1284), .O(gate511inter0));
  nand2 gate1500(.a(gate511inter0), .b(s_136), .O(gate511inter1));
  and2  gate1501(.a(G1285), .b(G1284), .O(gate511inter2));
  inv1  gate1502(.a(s_136), .O(gate511inter3));
  inv1  gate1503(.a(s_137), .O(gate511inter4));
  nand2 gate1504(.a(gate511inter4), .b(gate511inter3), .O(gate511inter5));
  nor2  gate1505(.a(gate511inter5), .b(gate511inter2), .O(gate511inter6));
  inv1  gate1506(.a(G1284), .O(gate511inter7));
  inv1  gate1507(.a(G1285), .O(gate511inter8));
  nand2 gate1508(.a(gate511inter8), .b(gate511inter7), .O(gate511inter9));
  nand2 gate1509(.a(s_137), .b(gate511inter3), .O(gate511inter10));
  nor2  gate1510(.a(gate511inter10), .b(gate511inter9), .O(gate511inter11));
  nor2  gate1511(.a(gate511inter11), .b(gate511inter6), .O(gate511inter12));
  nand2 gate1512(.a(gate511inter12), .b(gate511inter1), .O(G1320));
nand2 gate512( .a(G1286), .b(G1287), .O(G1321) );
nand2 gate513( .a(G1288), .b(G1289), .O(G1322) );
nand2 gate514( .a(G1290), .b(G1291), .O(G1323) );
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule