module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);

input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;//RE__PI;

input s_0,s_1;//RE__ALLOW(00,01,10,11);
input s_2,s_3;//RE__ALLOW(00,01,10,11);
input s_4,s_5;//RE__ALLOW(00,01,10,11);
input s_6,s_7;//RE__ALLOW(00,01,10,11);
input s_8,s_9;//RE__ALLOW(00,01,10,11);
input s_10,s_11;//RE__ALLOW(00,01,10,11);
input s_12,s_13;//RE__ALLOW(00,01,10,11);
input s_14,s_15;//RE__ALLOW(00,01,10,11);
input s_16,s_17;//RE__ALLOW(00,01,10,11);
input s_18,s_19;//RE__ALLOW(00,01,10,11);
input s_20,s_21;//RE__ALLOW(00,01,10,11);
input s_22,s_23;//RE__ALLOW(00,01,10,11);
input s_24,s_25;//RE__ALLOW(00,01,10,11);
input s_26,s_27;//RE__ALLOW(00,01,10,11);
input s_28,s_29;//RE__ALLOW(00,01,10,11);
input s_30,s_31;//RE__ALLOW(00,01,10,11);
input s_32,s_33;//RE__ALLOW(00,01,10,11);
input s_34,s_35;//RE__ALLOW(00,01,10,11);
input s_36,s_37;//RE__ALLOW(00,01,10,11);
input s_38,s_39;//RE__ALLOW(00,01,10,11);
input s_40,s_41;//RE__ALLOW(00,01,10,11);
input s_42,s_43;//RE__ALLOW(00,01,10,11);
input s_44,s_45;//RE__ALLOW(00,01,10,11);
input s_46,s_47;//RE__ALLOW(00,01,10,11);
input s_48,s_49;//RE__ALLOW(00,01,10,11);
input s_50,s_51;//RE__ALLOW(00,01,10,11);
input s_52,s_53;//RE__ALLOW(00,01,10,11);
input s_54,s_55;//RE__ALLOW(00,01,10,11);
input s_56,s_57;//RE__ALLOW(00,01,10,11);
input s_58,s_59;//RE__ALLOW(00,01,10,11);
input s_60,s_61;//RE__ALLOW(00,01,10,11);
input s_62,s_63;//RE__ALLOW(00,01,10,11);
input s_64,s_65;//RE__ALLOW(00,01,10,11);
input s_66,s_67;//RE__ALLOW(00,01,10,11);
input s_68,s_69;//RE__ALLOW(00,01,10,11);
input s_70,s_71;//RE__ALLOW(00,01,10,11);
input s_72,s_73;//RE__ALLOW(00,01,10,11);
input s_74,s_75;//RE__ALLOW(00,01,10,11);
input s_76,s_77;//RE__ALLOW(00,01,10,11);
input s_78,s_79;//RE__ALLOW(00,01,10,11);
input s_80,s_81;//RE__ALLOW(00,01,10,11);
input s_82,s_83;//RE__ALLOW(00,01,10,11);
input s_84,s_85;//RE__ALLOW(00,01,10,11);
input s_86,s_87;//RE__ALLOW(00,01,10,11);
input s_88,s_89;//RE__ALLOW(00,01,10,11);
input s_90,s_91;//RE__ALLOW(00,01,10,11);
input s_92,s_93;//RE__ALLOW(00,01,10,11);
input s_94,s_95;//RE__ALLOW(00,01,10,11);
input s_96,s_97;//RE__ALLOW(00,01,10,11);
input s_98,s_99;//RE__ALLOW(00,01,10,11);
input s_100,s_101;//RE__ALLOW(00,01,10,11);
input s_102,s_103;//RE__ALLOW(00,01,10,11);
input s_104,s_105;//RE__ALLOW(00,01,10,11);
input s_106,s_107;//RE__ALLOW(00,01,10,11);
input s_108,s_109;//RE__ALLOW(00,01,10,11);
input s_110,s_111;//RE__ALLOW(00,01,10,11);
input s_112,s_113;//RE__ALLOW(00,01,10,11);
input s_114,s_115;//RE__ALLOW(00,01,10,11);
input s_116,s_117;//RE__ALLOW(00,01,10,11);
input s_118,s_119;//RE__ALLOW(00,01,10,11);
input s_120,s_121;//RE__ALLOW(00,01,10,11);
input s_122,s_123;//RE__ALLOW(00,01,10,11);
input s_124,s_125;//RE__ALLOW(00,01,10,11);
input s_126,s_127;//RE__ALLOW(00,01,10,11);
input s_128,s_129;//RE__ALLOW(00,01,10,11);
input s_130,s_131;//RE__ALLOW(00,01,10,11);
input s_132,s_133;//RE__ALLOW(00,01,10,11);
input s_134,s_135;//RE__ALLOW(00,01,10,11);
input s_136,s_137;//RE__ALLOW(00,01,10,11);
input s_138,s_139;//RE__ALLOW(00,01,10,11);
input s_140,s_141;//RE__ALLOW(00,01,10,11);
input s_142,s_143;//RE__ALLOW(00,01,10,11);
input s_144,s_145;//RE__ALLOW(00,01,10,11);
input s_146,s_147;//RE__ALLOW(00,01,10,11);
input s_148,s_149;//RE__ALLOW(00,01,10,11);
input s_150,s_151;//RE__ALLOW(00,01,10,11);
input s_152,s_153;//RE__ALLOW(00,01,10,11);
input s_154,s_155;//RE__ALLOW(00,01,10,11);
input s_156,s_157;//RE__ALLOW(00,01,10,11);
input s_158,s_159;//RE__ALLOW(00,01,10,11);
input s_160,s_161;//RE__ALLOW(00,01,10,11);
input s_162,s_163;//RE__ALLOW(00,01,10,11);
input s_164,s_165;//RE__ALLOW(00,01,10,11);
input s_166,s_167;//RE__ALLOW(00,01,10,11);
input s_168,s_169;//RE__ALLOW(00,01,10,11);
input s_170,s_171;//RE__ALLOW(00,01,10,11);
input s_172,s_173;//RE__ALLOW(00,01,10,11);
input s_174,s_175;//RE__ALLOW(00,01,10,11);
input s_176,s_177;//RE__ALLOW(00,01,10,11);
input s_178,s_179;//RE__ALLOW(00,01,10,11);
input s_180,s_181;//RE__ALLOW(00,01,10,11);
input s_182,s_183;//RE__ALLOW(00,01,10,11);
input s_184,s_185;//RE__ALLOW(00,01,10,11);
input s_186,s_187;//RE__ALLOW(00,01,10,11);
input s_188,s_189;//RE__ALLOW(00,01,10,11);
input s_190,s_191;//RE__ALLOW(00,01,10,11);
input s_192,s_193;//RE__ALLOW(00,01,10,11);
input s_194,s_195;//RE__ALLOW(00,01,10,11);
input s_196,s_197;//RE__ALLOW(00,01,10,11);
input s_198,s_199;//RE__ALLOW(00,01,10,11);
input s_200,s_201;//RE__ALLOW(00,01,10,11);
input s_202,s_203;//RE__ALLOW(00,01,10,11);
input s_204,s_205;//RE__ALLOW(00,01,10,11);
input s_206,s_207;//RE__ALLOW(00,01,10,11);
input s_208,s_209;//RE__ALLOW(00,01,10,11);
input s_210,s_211;//RE__ALLOW(00,01,10,11);
input s_212,s_213;//RE__ALLOW(00,01,10,11);
input s_214,s_215;//RE__ALLOW(00,01,10,11);
input s_216,s_217;//RE__ALLOW(00,01,10,11);
input s_218,s_219;//RE__ALLOW(00,01,10,11);
input s_220,s_221;//RE__ALLOW(00,01,10,11);
input s_222,s_223;//RE__ALLOW(00,01,10,11);
input s_224,s_225;//RE__ALLOW(00,01,10,11);
input s_226,s_227;//RE__ALLOW(00,01,10,11);
input s_228,s_229;//RE__ALLOW(00,01,10,11);
input s_230,s_231;//RE__ALLOW(00,01,10,11);
input s_232,s_233;//RE__ALLOW(00,01,10,11);
input s_234,s_235;//RE__ALLOW(00,01,10,11);
input s_236,s_237;//RE__ALLOW(00,01,10,11);
input s_238,s_239;//RE__ALLOW(00,01,10,11);
input s_240,s_241;//RE__ALLOW(00,01,10,11);
input s_242,s_243;//RE__ALLOW(00,01,10,11);
input s_244,s_245;//RE__ALLOW(00,01,10,11);
input s_246,s_247;//RE__ALLOW(00,01,10,11);
input s_248,s_249;//RE__ALLOW(00,01,10,11);
input s_250,s_251;//RE__ALLOW(00,01,10,11);
input s_252,s_253;//RE__ALLOW(00,01,10,11);
input s_254,s_255;//RE__ALLOW(00,01,10,11);
input s_256,s_257;//RE__ALLOW(00,01,10,11);
input s_258,s_259;//RE__ALLOW(00,01,10,11);
input s_260,s_261;//RE__ALLOW(00,01,10,11);
input s_262,s_263;//RE__ALLOW(00,01,10,11);
input s_264,s_265;//RE__ALLOW(00,01,10,11);
input s_266,s_267;//RE__ALLOW(00,01,10,11);
input s_268,s_269;//RE__ALLOW(00,01,10,11);
input s_270,s_271;//RE__ALLOW(00,01,10,11);
input s_272,s_273;//RE__ALLOW(00,01,10,11);
input s_274,s_275;//RE__ALLOW(00,01,10,11);
input s_276,s_277;//RE__ALLOW(00,01,10,11);
input s_278,s_279;//RE__ALLOW(00,01,10,11);
input s_280,s_281;//RE__ALLOW(00,01,10,11);
input s_282,s_283;//RE__ALLOW(00,01,10,11);
input s_284,s_285;//RE__ALLOW(00,01,10,11);
input s_286,s_287;//RE__ALLOW(00,01,10,11);
input s_288,s_289;//RE__ALLOW(00,01,10,11);
input s_290,s_291;//RE__ALLOW(00,01,10,11);
input s_292,s_293;//RE__ALLOW(00,01,10,11);
input s_294,s_295;//RE__ALLOW(00,01,10,11);
input s_296,s_297;//RE__ALLOW(00,01,10,11);
input s_298,s_299;//RE__ALLOW(00,01,10,11);
input s_300,s_301;//RE__ALLOW(00,01,10,11);
input s_302,s_303;//RE__ALLOW(00,01,10,11);
input s_304,s_305;//RE__ALLOW(00,01,10,11);
input s_306,s_307;//RE__ALLOW(00,01,10,11);
input s_308,s_309;//RE__ALLOW(00,01,10,11);
input s_310,s_311;//RE__ALLOW(00,01,10,11);
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;

  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate209inter0, gate209inter1, gate209inter2, gate209inter3, gate209inter4, gate209inter5, gate209inter6, gate209inter7, gate209inter8, gate209inter9, gate209inter10, gate209inter11, gate209inter12, gate174inter0, gate174inter1, gate174inter2, gate174inter3, gate174inter4, gate174inter5, gate174inter6, gate174inter7, gate174inter8, gate174inter9, gate174inter10, gate174inter11, gate174inter12, gate96inter0, gate96inter1, gate96inter2, gate96inter3, gate96inter4, gate96inter5, gate96inter6, gate96inter7, gate96inter8, gate96inter9, gate96inter10, gate96inter11, gate96inter12, gate133inter0, gate133inter1, gate133inter2, gate133inter3, gate133inter4, gate133inter5, gate133inter6, gate133inter7, gate133inter8, gate133inter9, gate133inter10, gate133inter11, gate133inter12, gate76inter0, gate76inter1, gate76inter2, gate76inter3, gate76inter4, gate76inter5, gate76inter6, gate76inter7, gate76inter8, gate76inter9, gate76inter10, gate76inter11, gate76inter12, gate63inter0, gate63inter1, gate63inter2, gate63inter3, gate63inter4, gate63inter5, gate63inter6, gate63inter7, gate63inter8, gate63inter9, gate63inter10, gate63inter11, gate63inter12, gate41inter0, gate41inter1, gate41inter2, gate41inter3, gate41inter4, gate41inter5, gate41inter6, gate41inter7, gate41inter8, gate41inter9, gate41inter10, gate41inter11, gate41inter12, gate285inter0, gate285inter1, gate285inter2, gate285inter3, gate285inter4, gate285inter5, gate285inter6, gate285inter7, gate285inter8, gate285inter9, gate285inter10, gate285inter11, gate285inter12, gate36inter0, gate36inter1, gate36inter2, gate36inter3, gate36inter4, gate36inter5, gate36inter6, gate36inter7, gate36inter8, gate36inter9, gate36inter10, gate36inter11, gate36inter12, gate9inter0, gate9inter1, gate9inter2, gate9inter3, gate9inter4, gate9inter5, gate9inter6, gate9inter7, gate9inter8, gate9inter9, gate9inter10, gate9inter11, gate9inter12, gate65inter0, gate65inter1, gate65inter2, gate65inter3, gate65inter4, gate65inter5, gate65inter6, gate65inter7, gate65inter8, gate65inter9, gate65inter10, gate65inter11, gate65inter12, gate491inter0, gate491inter1, gate491inter2, gate491inter3, gate491inter4, gate491inter5, gate491inter6, gate491inter7, gate491inter8, gate491inter9, gate491inter10, gate491inter11, gate491inter12, gate47inter0, gate47inter1, gate47inter2, gate47inter3, gate47inter4, gate47inter5, gate47inter6, gate47inter7, gate47inter8, gate47inter9, gate47inter10, gate47inter11, gate47inter12, gate503inter0, gate503inter1, gate503inter2, gate503inter3, gate503inter4, gate503inter5, gate503inter6, gate503inter7, gate503inter8, gate503inter9, gate503inter10, gate503inter11, gate503inter12, gate138inter0, gate138inter1, gate138inter2, gate138inter3, gate138inter4, gate138inter5, gate138inter6, gate138inter7, gate138inter8, gate138inter9, gate138inter10, gate138inter11, gate138inter12, gate11inter0, gate11inter1, gate11inter2, gate11inter3, gate11inter4, gate11inter5, gate11inter6, gate11inter7, gate11inter8, gate11inter9, gate11inter10, gate11inter11, gate11inter12, gate249inter0, gate249inter1, gate249inter2, gate249inter3, gate249inter4, gate249inter5, gate249inter6, gate249inter7, gate249inter8, gate249inter9, gate249inter10, gate249inter11, gate249inter12, gate269inter0, gate269inter1, gate269inter2, gate269inter3, gate269inter4, gate269inter5, gate269inter6, gate269inter7, gate269inter8, gate269inter9, gate269inter10, gate269inter11, gate269inter12, gate188inter0, gate188inter1, gate188inter2, gate188inter3, gate188inter4, gate188inter5, gate188inter6, gate188inter7, gate188inter8, gate188inter9, gate188inter10, gate188inter11, gate188inter12, gate444inter0, gate444inter1, gate444inter2, gate444inter3, gate444inter4, gate444inter5, gate444inter6, gate444inter7, gate444inter8, gate444inter9, gate444inter10, gate444inter11, gate444inter12, gate493inter0, gate493inter1, gate493inter2, gate493inter3, gate493inter4, gate493inter5, gate493inter6, gate493inter7, gate493inter8, gate493inter9, gate493inter10, gate493inter11, gate493inter12, gate86inter0, gate86inter1, gate86inter2, gate86inter3, gate86inter4, gate86inter5, gate86inter6, gate86inter7, gate86inter8, gate86inter9, gate86inter10, gate86inter11, gate86inter12, gate423inter0, gate423inter1, gate423inter2, gate423inter3, gate423inter4, gate423inter5, gate423inter6, gate423inter7, gate423inter8, gate423inter9, gate423inter10, gate423inter11, gate423inter12, gate271inter0, gate271inter1, gate271inter2, gate271inter3, gate271inter4, gate271inter5, gate271inter6, gate271inter7, gate271inter8, gate271inter9, gate271inter10, gate271inter11, gate271inter12, gate225inter0, gate225inter1, gate225inter2, gate225inter3, gate225inter4, gate225inter5, gate225inter6, gate225inter7, gate225inter8, gate225inter9, gate225inter10, gate225inter11, gate225inter12, gate164inter0, gate164inter1, gate164inter2, gate164inter3, gate164inter4, gate164inter5, gate164inter6, gate164inter7, gate164inter8, gate164inter9, gate164inter10, gate164inter11, gate164inter12, gate158inter0, gate158inter1, gate158inter2, gate158inter3, gate158inter4, gate158inter5, gate158inter6, gate158inter7, gate158inter8, gate158inter9, gate158inter10, gate158inter11, gate158inter12, gate393inter0, gate393inter1, gate393inter2, gate393inter3, gate393inter4, gate393inter5, gate393inter6, gate393inter7, gate393inter8, gate393inter9, gate393inter10, gate393inter11, gate393inter12, gate187inter0, gate187inter1, gate187inter2, gate187inter3, gate187inter4, gate187inter5, gate187inter6, gate187inter7, gate187inter8, gate187inter9, gate187inter10, gate187inter11, gate187inter12, gate422inter0, gate422inter1, gate422inter2, gate422inter3, gate422inter4, gate422inter5, gate422inter6, gate422inter7, gate422inter8, gate422inter9, gate422inter10, gate422inter11, gate422inter12, gate98inter0, gate98inter1, gate98inter2, gate98inter3, gate98inter4, gate98inter5, gate98inter6, gate98inter7, gate98inter8, gate98inter9, gate98inter10, gate98inter11, gate98inter12, gate166inter0, gate166inter1, gate166inter2, gate166inter3, gate166inter4, gate166inter5, gate166inter6, gate166inter7, gate166inter8, gate166inter9, gate166inter10, gate166inter11, gate166inter12, gate279inter0, gate279inter1, gate279inter2, gate279inter3, gate279inter4, gate279inter5, gate279inter6, gate279inter7, gate279inter8, gate279inter9, gate279inter10, gate279inter11, gate279inter12, gate265inter0, gate265inter1, gate265inter2, gate265inter3, gate265inter4, gate265inter5, gate265inter6, gate265inter7, gate265inter8, gate265inter9, gate265inter10, gate265inter11, gate265inter12, gate216inter0, gate216inter1, gate216inter2, gate216inter3, gate216inter4, gate216inter5, gate216inter6, gate216inter7, gate216inter8, gate216inter9, gate216inter10, gate216inter11, gate216inter12, gate172inter0, gate172inter1, gate172inter2, gate172inter3, gate172inter4, gate172inter5, gate172inter6, gate172inter7, gate172inter8, gate172inter9, gate172inter10, gate172inter11, gate172inter12, gate449inter0, gate449inter1, gate449inter2, gate449inter3, gate449inter4, gate449inter5, gate449inter6, gate449inter7, gate449inter8, gate449inter9, gate449inter10, gate449inter11, gate449inter12, gate135inter0, gate135inter1, gate135inter2, gate135inter3, gate135inter4, gate135inter5, gate135inter6, gate135inter7, gate135inter8, gate135inter9, gate135inter10, gate135inter11, gate135inter12, gate455inter0, gate455inter1, gate455inter2, gate455inter3, gate455inter4, gate455inter5, gate455inter6, gate455inter7, gate455inter8, gate455inter9, gate455inter10, gate455inter11, gate455inter12, gate179inter0, gate179inter1, gate179inter2, gate179inter3, gate179inter4, gate179inter5, gate179inter6, gate179inter7, gate179inter8, gate179inter9, gate179inter10, gate179inter11, gate179inter12, gate155inter0, gate155inter1, gate155inter2, gate155inter3, gate155inter4, gate155inter5, gate155inter6, gate155inter7, gate155inter8, gate155inter9, gate155inter10, gate155inter11, gate155inter12, gate157inter0, gate157inter1, gate157inter2, gate157inter3, gate157inter4, gate157inter5, gate157inter6, gate157inter7, gate157inter8, gate157inter9, gate157inter10, gate157inter11, gate157inter12, gate22inter0, gate22inter1, gate22inter2, gate22inter3, gate22inter4, gate22inter5, gate22inter6, gate22inter7, gate22inter8, gate22inter9, gate22inter10, gate22inter11, gate22inter12, gate230inter0, gate230inter1, gate230inter2, gate230inter3, gate230inter4, gate230inter5, gate230inter6, gate230inter7, gate230inter8, gate230inter9, gate230inter10, gate230inter11, gate230inter12, gate59inter0, gate59inter1, gate59inter2, gate59inter3, gate59inter4, gate59inter5, gate59inter6, gate59inter7, gate59inter8, gate59inter9, gate59inter10, gate59inter11, gate59inter12, gate276inter0, gate276inter1, gate276inter2, gate276inter3, gate276inter4, gate276inter5, gate276inter6, gate276inter7, gate276inter8, gate276inter9, gate276inter10, gate276inter11, gate276inter12, gate437inter0, gate437inter1, gate437inter2, gate437inter3, gate437inter4, gate437inter5, gate437inter6, gate437inter7, gate437inter8, gate437inter9, gate437inter10, gate437inter11, gate437inter12, gate273inter0, gate273inter1, gate273inter2, gate273inter3, gate273inter4, gate273inter5, gate273inter6, gate273inter7, gate273inter8, gate273inter9, gate273inter10, gate273inter11, gate273inter12, gate507inter0, gate507inter1, gate507inter2, gate507inter3, gate507inter4, gate507inter5, gate507inter6, gate507inter7, gate507inter8, gate507inter9, gate507inter10, gate507inter11, gate507inter12, gate18inter0, gate18inter1, gate18inter2, gate18inter3, gate18inter4, gate18inter5, gate18inter6, gate18inter7, gate18inter8, gate18inter9, gate18inter10, gate18inter11, gate18inter12, gate144inter0, gate144inter1, gate144inter2, gate144inter3, gate144inter4, gate144inter5, gate144inter6, gate144inter7, gate144inter8, gate144inter9, gate144inter10, gate144inter11, gate144inter12, gate463inter0, gate463inter1, gate463inter2, gate463inter3, gate463inter4, gate463inter5, gate463inter6, gate463inter7, gate463inter8, gate463inter9, gate463inter10, gate463inter11, gate463inter12, gate73inter0, gate73inter1, gate73inter2, gate73inter3, gate73inter4, gate73inter5, gate73inter6, gate73inter7, gate73inter8, gate73inter9, gate73inter10, gate73inter11, gate73inter12, gate190inter0, gate190inter1, gate190inter2, gate190inter3, gate190inter4, gate190inter5, gate190inter6, gate190inter7, gate190inter8, gate190inter9, gate190inter10, gate190inter11, gate190inter12, gate501inter0, gate501inter1, gate501inter2, gate501inter3, gate501inter4, gate501inter5, gate501inter6, gate501inter7, gate501inter8, gate501inter9, gate501inter10, gate501inter11, gate501inter12, gate452inter0, gate452inter1, gate452inter2, gate452inter3, gate452inter4, gate452inter5, gate452inter6, gate452inter7, gate452inter8, gate452inter9, gate452inter10, gate452inter11, gate452inter12, gate134inter0, gate134inter1, gate134inter2, gate134inter3, gate134inter4, gate134inter5, gate134inter6, gate134inter7, gate134inter8, gate134inter9, gate134inter10, gate134inter11, gate134inter12, gate132inter0, gate132inter1, gate132inter2, gate132inter3, gate132inter4, gate132inter5, gate132inter6, gate132inter7, gate132inter8, gate132inter9, gate132inter10, gate132inter11, gate132inter12, gate425inter0, gate425inter1, gate425inter2, gate425inter3, gate425inter4, gate425inter5, gate425inter6, gate425inter7, gate425inter8, gate425inter9, gate425inter10, gate425inter11, gate425inter12, gate81inter0, gate81inter1, gate81inter2, gate81inter3, gate81inter4, gate81inter5, gate81inter6, gate81inter7, gate81inter8, gate81inter9, gate81inter10, gate81inter11, gate81inter12, gate514inter0, gate514inter1, gate514inter2, gate514inter3, gate514inter4, gate514inter5, gate514inter6, gate514inter7, gate514inter8, gate514inter9, gate514inter10, gate514inter11, gate514inter12, gate295inter0, gate295inter1, gate295inter2, gate295inter3, gate295inter4, gate295inter5, gate295inter6, gate295inter7, gate295inter8, gate295inter9, gate295inter10, gate295inter11, gate295inter12, gate286inter0, gate286inter1, gate286inter2, gate286inter3, gate286inter4, gate286inter5, gate286inter6, gate286inter7, gate286inter8, gate286inter9, gate286inter10, gate286inter11, gate286inter12, gate121inter0, gate121inter1, gate121inter2, gate121inter3, gate121inter4, gate121inter5, gate121inter6, gate121inter7, gate121inter8, gate121inter9, gate121inter10, gate121inter11, gate121inter12, gate147inter0, gate147inter1, gate147inter2, gate147inter3, gate147inter4, gate147inter5, gate147inter6, gate147inter7, gate147inter8, gate147inter9, gate147inter10, gate147inter11, gate147inter12, gate77inter0, gate77inter1, gate77inter2, gate77inter3, gate77inter4, gate77inter5, gate77inter6, gate77inter7, gate77inter8, gate77inter9, gate77inter10, gate77inter11, gate77inter12, gate114inter0, gate114inter1, gate114inter2, gate114inter3, gate114inter4, gate114inter5, gate114inter6, gate114inter7, gate114inter8, gate114inter9, gate114inter10, gate114inter11, gate114inter12, gate508inter0, gate508inter1, gate508inter2, gate508inter3, gate508inter4, gate508inter5, gate508inter6, gate508inter7, gate508inter8, gate508inter9, gate508inter10, gate508inter11, gate508inter12, gate54inter0, gate54inter1, gate54inter2, gate54inter3, gate54inter4, gate54inter5, gate54inter6, gate54inter7, gate54inter8, gate54inter9, gate54inter10, gate54inter11, gate54inter12, gate124inter0, gate124inter1, gate124inter2, gate124inter3, gate124inter4, gate124inter5, gate124inter6, gate124inter7, gate124inter8, gate124inter9, gate124inter10, gate124inter11, gate124inter12, gate227inter0, gate227inter1, gate227inter2, gate227inter3, gate227inter4, gate227inter5, gate227inter6, gate227inter7, gate227inter8, gate227inter9, gate227inter10, gate227inter11, gate227inter12, gate58inter0, gate58inter1, gate58inter2, gate58inter3, gate58inter4, gate58inter5, gate58inter6, gate58inter7, gate58inter8, gate58inter9, gate58inter10, gate58inter11, gate58inter12, gate60inter0, gate60inter1, gate60inter2, gate60inter3, gate60inter4, gate60inter5, gate60inter6, gate60inter7, gate60inter8, gate60inter9, gate60inter10, gate60inter11, gate60inter12, gate23inter0, gate23inter1, gate23inter2, gate23inter3, gate23inter4, gate23inter5, gate23inter6, gate23inter7, gate23inter8, gate23inter9, gate23inter10, gate23inter11, gate23inter12, gate104inter0, gate104inter1, gate104inter2, gate104inter3, gate104inter4, gate104inter5, gate104inter6, gate104inter7, gate104inter8, gate104inter9, gate104inter10, gate104inter11, gate104inter12, gate262inter0, gate262inter1, gate262inter2, gate262inter3, gate262inter4, gate262inter5, gate262inter6, gate262inter7, gate262inter8, gate262inter9, gate262inter10, gate262inter11, gate262inter12, gate152inter0, gate152inter1, gate152inter2, gate152inter3, gate152inter4, gate152inter5, gate152inter6, gate152inter7, gate152inter8, gate152inter9, gate152inter10, gate152inter11, gate152inter12, gate31inter0, gate31inter1, gate31inter2, gate31inter3, gate31inter4, gate31inter5, gate31inter6, gate31inter7, gate31inter8, gate31inter9, gate31inter10, gate31inter11, gate31inter12, gate111inter0, gate111inter1, gate111inter2, gate111inter3, gate111inter4, gate111inter5, gate111inter6, gate111inter7, gate111inter8, gate111inter9, gate111inter10, gate111inter11, gate111inter12, gate418inter0, gate418inter1, gate418inter2, gate418inter3, gate418inter4, gate418inter5, gate418inter6, gate418inter7, gate418inter8, gate418inter9, gate418inter10, gate418inter11, gate418inter12, gate413inter0, gate413inter1, gate413inter2, gate413inter3, gate413inter4, gate413inter5, gate413inter6, gate413inter7, gate413inter8, gate413inter9, gate413inter10, gate413inter11, gate413inter12, gate167inter0, gate167inter1, gate167inter2, gate167inter3, gate167inter4, gate167inter5, gate167inter6, gate167inter7, gate167inter8, gate167inter9, gate167inter10, gate167inter11, gate167inter12, gate436inter0, gate436inter1, gate436inter2, gate436inter3, gate436inter4, gate436inter5, gate436inter6, gate436inter7, gate436inter8, gate436inter9, gate436inter10, gate436inter11, gate436inter12, gate496inter0, gate496inter1, gate496inter2, gate496inter3, gate496inter4, gate496inter5, gate496inter6, gate496inter7, gate496inter8, gate496inter9, gate496inter10, gate496inter11, gate496inter12, gate92inter0, gate92inter1, gate92inter2, gate92inter3, gate92inter4, gate92inter5, gate92inter6, gate92inter7, gate92inter8, gate92inter9, gate92inter10, gate92inter11, gate92inter12, gate107inter0, gate107inter1, gate107inter2, gate107inter3, gate107inter4, gate107inter5, gate107inter6, gate107inter7, gate107inter8, gate107inter9, gate107inter10, gate107inter11, gate107inter12, gate185inter0, gate185inter1, gate185inter2, gate185inter3, gate185inter4, gate185inter5, gate185inter6, gate185inter7, gate185inter8, gate185inter9, gate185inter10, gate185inter11, gate185inter12, gate211inter0, gate211inter1, gate211inter2, gate211inter3, gate211inter4, gate211inter5, gate211inter6, gate211inter7, gate211inter8, gate211inter9, gate211inter10, gate211inter11, gate211inter12, gate474inter0, gate474inter1, gate474inter2, gate474inter3, gate474inter4, gate474inter5, gate474inter6, gate474inter7, gate474inter8, gate474inter9, gate474inter10, gate474inter11, gate474inter12, gate389inter0, gate389inter1, gate389inter2, gate389inter3, gate389inter4, gate389inter5, gate389inter6, gate389inter7, gate389inter8, gate389inter9, gate389inter10, gate389inter11, gate389inter12, gate416inter0, gate416inter1, gate416inter2, gate416inter3, gate416inter4, gate416inter5, gate416inter6, gate416inter7, gate416inter8, gate416inter9, gate416inter10, gate416inter11, gate416inter12, gate290inter0, gate290inter1, gate290inter2, gate290inter3, gate290inter4, gate290inter5, gate290inter6, gate290inter7, gate290inter8, gate290inter9, gate290inter10, gate290inter11, gate290inter12, gate223inter0, gate223inter1, gate223inter2, gate223inter3, gate223inter4, gate223inter5, gate223inter6, gate223inter7, gate223inter8, gate223inter9, gate223inter10, gate223inter11, gate223inter12, gate494inter0, gate494inter1, gate494inter2, gate494inter3, gate494inter4, gate494inter5, gate494inter6, gate494inter7, gate494inter8, gate494inter9, gate494inter10, gate494inter11, gate494inter12, gate294inter0, gate294inter1, gate294inter2, gate294inter3, gate294inter4, gate294inter5, gate294inter6, gate294inter7, gate294inter8, gate294inter9, gate294inter10, gate294inter11, gate294inter12, gate180inter0, gate180inter1, gate180inter2, gate180inter3, gate180inter4, gate180inter5, gate180inter6, gate180inter7, gate180inter8, gate180inter9, gate180inter10, gate180inter11, gate180inter12, gate287inter0, gate287inter1, gate287inter2, gate287inter3, gate287inter4, gate287inter5, gate287inter6, gate287inter7, gate287inter8, gate287inter9, gate287inter10, gate287inter11, gate287inter12, gate129inter0, gate129inter1, gate129inter2, gate129inter3, gate129inter4, gate129inter5, gate129inter6, gate129inter7, gate129inter8, gate129inter9, gate129inter10, gate129inter11, gate129inter12, gate398inter0, gate398inter1, gate398inter2, gate398inter3, gate398inter4, gate398inter5, gate398inter6, gate398inter7, gate398inter8, gate398inter9, gate398inter10, gate398inter11, gate398inter12, gate137inter0, gate137inter1, gate137inter2, gate137inter3, gate137inter4, gate137inter5, gate137inter6, gate137inter7, gate137inter8, gate137inter9, gate137inter10, gate137inter11, gate137inter12, gate128inter0, gate128inter1, gate128inter2, gate128inter3, gate128inter4, gate128inter5, gate128inter6, gate128inter7, gate128inter8, gate128inter9, gate128inter10, gate128inter11, gate128inter12, gate25inter0, gate25inter1, gate25inter2, gate25inter3, gate25inter4, gate25inter5, gate25inter6, gate25inter7, gate25inter8, gate25inter9, gate25inter10, gate25inter11, gate25inter12, gate397inter0, gate397inter1, gate397inter2, gate397inter3, gate397inter4, gate397inter5, gate397inter6, gate397inter7, gate397inter8, gate397inter9, gate397inter10, gate397inter11, gate397inter12, gate400inter0, gate400inter1, gate400inter2, gate400inter3, gate400inter4, gate400inter5, gate400inter6, gate400inter7, gate400inter8, gate400inter9, gate400inter10, gate400inter11, gate400inter12, gate102inter0, gate102inter1, gate102inter2, gate102inter3, gate102inter4, gate102inter5, gate102inter6, gate102inter7, gate102inter8, gate102inter9, gate102inter10, gate102inter11, gate102inter12, gate388inter0, gate388inter1, gate388inter2, gate388inter3, gate388inter4, gate388inter5, gate388inter6, gate388inter7, gate388inter8, gate388inter9, gate388inter10, gate388inter11, gate388inter12, gate32inter0, gate32inter1, gate32inter2, gate32inter3, gate32inter4, gate32inter5, gate32inter6, gate32inter7, gate32inter8, gate32inter9, gate32inter10, gate32inter11, gate32inter12, gate235inter0, gate235inter1, gate235inter2, gate235inter3, gate235inter4, gate235inter5, gate235inter6, gate235inter7, gate235inter8, gate235inter9, gate235inter10, gate235inter11, gate235inter12, gate473inter0, gate473inter1, gate473inter2, gate473inter3, gate473inter4, gate473inter5, gate473inter6, gate473inter7, gate473inter8, gate473inter9, gate473inter10, gate473inter11, gate473inter12, gate283inter0, gate283inter1, gate283inter2, gate283inter3, gate283inter4, gate283inter5, gate283inter6, gate283inter7, gate283inter8, gate283inter9, gate283inter10, gate283inter11, gate283inter12, gate293inter0, gate293inter1, gate293inter2, gate293inter3, gate293inter4, gate293inter5, gate293inter6, gate293inter7, gate293inter8, gate293inter9, gate293inter10, gate293inter11, gate293inter12, gate82inter0, gate82inter1, gate82inter2, gate82inter3, gate82inter4, gate82inter5, gate82inter6, gate82inter7, gate82inter8, gate82inter9, gate82inter10, gate82inter11, gate82inter12, gate261inter0, gate261inter1, gate261inter2, gate261inter3, gate261inter4, gate261inter5, gate261inter6, gate261inter7, gate261inter8, gate261inter9, gate261inter10, gate261inter11, gate261inter12, gate239inter0, gate239inter1, gate239inter2, gate239inter3, gate239inter4, gate239inter5, gate239inter6, gate239inter7, gate239inter8, gate239inter9, gate239inter10, gate239inter11, gate239inter12, gate482inter0, gate482inter1, gate482inter2, gate482inter3, gate482inter4, gate482inter5, gate482inter6, gate482inter7, gate482inter8, gate482inter9, gate482inter10, gate482inter11, gate482inter12, gate197inter0, gate197inter1, gate197inter2, gate197inter3, gate197inter4, gate197inter5, gate197inter6, gate197inter7, gate197inter8, gate197inter9, gate197inter10, gate197inter11, gate197inter12, gate21inter0, gate21inter1, gate21inter2, gate21inter3, gate21inter4, gate21inter5, gate21inter6, gate21inter7, gate21inter8, gate21inter9, gate21inter10, gate21inter11, gate21inter12, gate510inter0, gate510inter1, gate510inter2, gate510inter3, gate510inter4, gate510inter5, gate510inter6, gate510inter7, gate510inter8, gate510inter9, gate510inter10, gate510inter11, gate510inter12, gate131inter0, gate131inter1, gate131inter2, gate131inter3, gate131inter4, gate131inter5, gate131inter6, gate131inter7, gate131inter8, gate131inter9, gate131inter10, gate131inter11, gate131inter12, gate232inter0, gate232inter1, gate232inter2, gate232inter3, gate232inter4, gate232inter5, gate232inter6, gate232inter7, gate232inter8, gate232inter9, gate232inter10, gate232inter11, gate232inter12, gate215inter0, gate215inter1, gate215inter2, gate215inter3, gate215inter4, gate215inter5, gate215inter6, gate215inter7, gate215inter8, gate215inter9, gate215inter10, gate215inter11, gate215inter12, gate255inter0, gate255inter1, gate255inter2, gate255inter3, gate255inter4, gate255inter5, gate255inter6, gate255inter7, gate255inter8, gate255inter9, gate255inter10, gate255inter11, gate255inter12, gate161inter0, gate161inter1, gate161inter2, gate161inter3, gate161inter4, gate161inter5, gate161inter6, gate161inter7, gate161inter8, gate161inter9, gate161inter10, gate161inter11, gate161inter12, gate116inter0, gate116inter1, gate116inter2, gate116inter3, gate116inter4, gate116inter5, gate116inter6, gate116inter7, gate116inter8, gate116inter9, gate116inter10, gate116inter11, gate116inter12, gate201inter0, gate201inter1, gate201inter2, gate201inter3, gate201inter4, gate201inter5, gate201inter6, gate201inter7, gate201inter8, gate201inter9, gate201inter10, gate201inter11, gate201inter12, gate89inter0, gate89inter1, gate89inter2, gate89inter3, gate89inter4, gate89inter5, gate89inter6, gate89inter7, gate89inter8, gate89inter9, gate89inter10, gate89inter11, gate89inter12, gate148inter0, gate148inter1, gate148inter2, gate148inter3, gate148inter4, gate148inter5, gate148inter6, gate148inter7, gate148inter8, gate148inter9, gate148inter10, gate148inter11, gate148inter12, gate53inter0, gate53inter1, gate53inter2, gate53inter3, gate53inter4, gate53inter5, gate53inter6, gate53inter7, gate53inter8, gate53inter9, gate53inter10, gate53inter11, gate53inter12, gate193inter0, gate193inter1, gate193inter2, gate193inter3, gate193inter4, gate193inter5, gate193inter6, gate193inter7, gate193inter8, gate193inter9, gate193inter10, gate193inter11, gate193inter12, gate504inter0, gate504inter1, gate504inter2, gate504inter3, gate504inter4, gate504inter5, gate504inter6, gate504inter7, gate504inter8, gate504inter9, gate504inter10, gate504inter11, gate504inter12, gate475inter0, gate475inter1, gate475inter2, gate475inter3, gate475inter4, gate475inter5, gate475inter6, gate475inter7, gate475inter8, gate475inter9, gate475inter10, gate475inter11, gate475inter12, gate511inter0, gate511inter1, gate511inter2, gate511inter3, gate511inter4, gate511inter5, gate511inter6, gate511inter7, gate511inter8, gate511inter9, gate511inter10, gate511inter11, gate511inter12, gate221inter0, gate221inter1, gate221inter2, gate221inter3, gate221inter4, gate221inter5, gate221inter6, gate221inter7, gate221inter8, gate221inter9, gate221inter10, gate221inter11, gate221inter12, gate448inter0, gate448inter1, gate448inter2, gate448inter3, gate448inter4, gate448inter5, gate448inter6, gate448inter7, gate448inter8, gate448inter9, gate448inter10, gate448inter11, gate448inter12, gate220inter0, gate220inter1, gate220inter2, gate220inter3, gate220inter4, gate220inter5, gate220inter6, gate220inter7, gate220inter8, gate220inter9, gate220inter10, gate220inter11, gate220inter12, gate417inter0, gate417inter1, gate417inter2, gate417inter3, gate417inter4, gate417inter5, gate417inter6, gate417inter7, gate417inter8, gate417inter9, gate417inter10, gate417inter11, gate417inter12, gate87inter0, gate87inter1, gate87inter2, gate87inter3, gate87inter4, gate87inter5, gate87inter6, gate87inter7, gate87inter8, gate87inter9, gate87inter10, gate87inter11, gate87inter12, gate228inter0, gate228inter1, gate228inter2, gate228inter3, gate228inter4, gate228inter5, gate228inter6, gate228inter7, gate228inter8, gate228inter9, gate228inter10, gate228inter11, gate228inter12, gate234inter0, gate234inter1, gate234inter2, gate234inter3, gate234inter4, gate234inter5, gate234inter6, gate234inter7, gate234inter8, gate234inter9, gate234inter10, gate234inter11, gate234inter12, gate268inter0, gate268inter1, gate268inter2, gate268inter3, gate268inter4, gate268inter5, gate268inter6, gate268inter7, gate268inter8, gate268inter9, gate268inter10, gate268inter11, gate268inter12, gate192inter0, gate192inter1, gate192inter2, gate192inter3, gate192inter4, gate192inter5, gate192inter6, gate192inter7, gate192inter8, gate192inter9, gate192inter10, gate192inter11, gate192inter12, gate479inter0, gate479inter1, gate479inter2, gate479inter3, gate479inter4, gate479inter5, gate479inter6, gate479inter7, gate479inter8, gate479inter9, gate479inter10, gate479inter11, gate479inter12, gate159inter0, gate159inter1, gate159inter2, gate159inter3, gate159inter4, gate159inter5, gate159inter6, gate159inter7, gate159inter8, gate159inter9, gate159inter10, gate159inter11, gate159inter12, gate20inter0, gate20inter1, gate20inter2, gate20inter3, gate20inter4, gate20inter5, gate20inter6, gate20inter7, gate20inter8, gate20inter9, gate20inter10, gate20inter11, gate20inter12, gate257inter0, gate257inter1, gate257inter2, gate257inter3, gate257inter4, gate257inter5, gate257inter6, gate257inter7, gate257inter8, gate257inter9, gate257inter10, gate257inter11, gate257inter12, gate162inter0, gate162inter1, gate162inter2, gate162inter3, gate162inter4, gate162inter5, gate162inter6, gate162inter7, gate162inter8, gate162inter9, gate162inter10, gate162inter11, gate162inter12, gate14inter0, gate14inter1, gate14inter2, gate14inter3, gate14inter4, gate14inter5, gate14inter6, gate14inter7, gate14inter8, gate14inter9, gate14inter10, gate14inter11, gate14inter12, gate233inter0, gate233inter1, gate233inter2, gate233inter3, gate233inter4, gate233inter5, gate233inter6, gate233inter7, gate233inter8, gate233inter9, gate233inter10, gate233inter11, gate233inter12, gate431inter0, gate431inter1, gate431inter2, gate431inter3, gate431inter4, gate431inter5, gate431inter6, gate431inter7, gate431inter8, gate431inter9, gate431inter10, gate431inter11, gate431inter12, gate253inter0, gate253inter1, gate253inter2, gate253inter3, gate253inter4, gate253inter5, gate253inter6, gate253inter7, gate253inter8, gate253inter9, gate253inter10, gate253inter11, gate253inter12, gate145inter0, gate145inter1, gate145inter2, gate145inter3, gate145inter4, gate145inter5, gate145inter6, gate145inter7, gate145inter8, gate145inter9, gate145inter10, gate145inter11, gate145inter12, gate56inter0, gate56inter1, gate56inter2, gate56inter3, gate56inter4, gate56inter5, gate56inter6, gate56inter7, gate56inter8, gate56inter9, gate56inter10, gate56inter11, gate56inter12, gate229inter0, gate229inter1, gate229inter2, gate229inter3, gate229inter4, gate229inter5, gate229inter6, gate229inter7, gate229inter8, gate229inter9, gate229inter10, gate229inter11, gate229inter12, gate109inter0, gate109inter1, gate109inter2, gate109inter3, gate109inter4, gate109inter5, gate109inter6, gate109inter7, gate109inter8, gate109inter9, gate109inter10, gate109inter11, gate109inter12, gate238inter0, gate238inter1, gate238inter2, gate238inter3, gate238inter4, gate238inter5, gate238inter6, gate238inter7, gate238inter8, gate238inter9, gate238inter10, gate238inter11, gate238inter12, gate203inter0, gate203inter1, gate203inter2, gate203inter3, gate203inter4, gate203inter5, gate203inter6, gate203inter7, gate203inter8, gate203inter9, gate203inter10, gate203inter11, gate203inter12;



and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );

  xor2  gate673(.a(G2), .b(G1), .O(gate9inter0));
  nand2 gate674(.a(gate9inter0), .b(s_18), .O(gate9inter1));
  and2  gate675(.a(G2), .b(G1), .O(gate9inter2));
  inv1  gate676(.a(s_18), .O(gate9inter3));
  inv1  gate677(.a(s_19), .O(gate9inter4));
  nand2 gate678(.a(gate9inter4), .b(gate9inter3), .O(gate9inter5));
  nor2  gate679(.a(gate9inter5), .b(gate9inter2), .O(gate9inter6));
  inv1  gate680(.a(G1), .O(gate9inter7));
  inv1  gate681(.a(G2), .O(gate9inter8));
  nand2 gate682(.a(gate9inter8), .b(gate9inter7), .O(gate9inter9));
  nand2 gate683(.a(s_19), .b(gate9inter3), .O(gate9inter10));
  nor2  gate684(.a(gate9inter10), .b(gate9inter9), .O(gate9inter11));
  nor2  gate685(.a(gate9inter11), .b(gate9inter6), .O(gate9inter12));
  nand2 gate686(.a(gate9inter12), .b(gate9inter1), .O(G266));
nand2 gate10( .a(G3), .b(G4), .O(G269) );

  xor2  gate757(.a(G6), .b(G5), .O(gate11inter0));
  nand2 gate758(.a(gate11inter0), .b(s_30), .O(gate11inter1));
  and2  gate759(.a(G6), .b(G5), .O(gate11inter2));
  inv1  gate760(.a(s_30), .O(gate11inter3));
  inv1  gate761(.a(s_31), .O(gate11inter4));
  nand2 gate762(.a(gate11inter4), .b(gate11inter3), .O(gate11inter5));
  nor2  gate763(.a(gate11inter5), .b(gate11inter2), .O(gate11inter6));
  inv1  gate764(.a(G5), .O(gate11inter7));
  inv1  gate765(.a(G6), .O(gate11inter8));
  nand2 gate766(.a(gate11inter8), .b(gate11inter7), .O(gate11inter9));
  nand2 gate767(.a(s_31), .b(gate11inter3), .O(gate11inter10));
  nor2  gate768(.a(gate11inter10), .b(gate11inter9), .O(gate11inter11));
  nor2  gate769(.a(gate11inter11), .b(gate11inter6), .O(gate11inter12));
  nand2 gate770(.a(gate11inter12), .b(gate11inter1), .O(G272));
nand2 gate12( .a(G7), .b(G8), .O(G275) );
nand2 gate13( .a(G9), .b(G10), .O(G278) );

  xor2  gate2591(.a(G12), .b(G11), .O(gate14inter0));
  nand2 gate2592(.a(gate14inter0), .b(s_292), .O(gate14inter1));
  and2  gate2593(.a(G12), .b(G11), .O(gate14inter2));
  inv1  gate2594(.a(s_292), .O(gate14inter3));
  inv1  gate2595(.a(s_293), .O(gate14inter4));
  nand2 gate2596(.a(gate14inter4), .b(gate14inter3), .O(gate14inter5));
  nor2  gate2597(.a(gate14inter5), .b(gate14inter2), .O(gate14inter6));
  inv1  gate2598(.a(G11), .O(gate14inter7));
  inv1  gate2599(.a(G12), .O(gate14inter8));
  nand2 gate2600(.a(gate14inter8), .b(gate14inter7), .O(gate14inter9));
  nand2 gate2601(.a(s_293), .b(gate14inter3), .O(gate14inter10));
  nor2  gate2602(.a(gate14inter10), .b(gate14inter9), .O(gate14inter11));
  nor2  gate2603(.a(gate14inter11), .b(gate14inter6), .O(gate14inter12));
  nand2 gate2604(.a(gate14inter12), .b(gate14inter1), .O(G281));
nand2 gate15( .a(G13), .b(G14), .O(G284) );
nand2 gate16( .a(G15), .b(G16), .O(G287) );
nand2 gate17( .a(G17), .b(G18), .O(G290) );

  xor2  gate1233(.a(G20), .b(G19), .O(gate18inter0));
  nand2 gate1234(.a(gate18inter0), .b(s_98), .O(gate18inter1));
  and2  gate1235(.a(G20), .b(G19), .O(gate18inter2));
  inv1  gate1236(.a(s_98), .O(gate18inter3));
  inv1  gate1237(.a(s_99), .O(gate18inter4));
  nand2 gate1238(.a(gate18inter4), .b(gate18inter3), .O(gate18inter5));
  nor2  gate1239(.a(gate18inter5), .b(gate18inter2), .O(gate18inter6));
  inv1  gate1240(.a(G19), .O(gate18inter7));
  inv1  gate1241(.a(G20), .O(gate18inter8));
  nand2 gate1242(.a(gate18inter8), .b(gate18inter7), .O(gate18inter9));
  nand2 gate1243(.a(s_99), .b(gate18inter3), .O(gate18inter10));
  nor2  gate1244(.a(gate18inter10), .b(gate18inter9), .O(gate18inter11));
  nor2  gate1245(.a(gate18inter11), .b(gate18inter6), .O(gate18inter12));
  nand2 gate1246(.a(gate18inter12), .b(gate18inter1), .O(G293));
nand2 gate19( .a(G21), .b(G22), .O(G296) );

  xor2  gate2549(.a(G24), .b(G23), .O(gate20inter0));
  nand2 gate2550(.a(gate20inter0), .b(s_286), .O(gate20inter1));
  and2  gate2551(.a(G24), .b(G23), .O(gate20inter2));
  inv1  gate2552(.a(s_286), .O(gate20inter3));
  inv1  gate2553(.a(s_287), .O(gate20inter4));
  nand2 gate2554(.a(gate20inter4), .b(gate20inter3), .O(gate20inter5));
  nor2  gate2555(.a(gate20inter5), .b(gate20inter2), .O(gate20inter6));
  inv1  gate2556(.a(G23), .O(gate20inter7));
  inv1  gate2557(.a(G24), .O(gate20inter8));
  nand2 gate2558(.a(gate20inter8), .b(gate20inter7), .O(gate20inter9));
  nand2 gate2559(.a(s_287), .b(gate20inter3), .O(gate20inter10));
  nor2  gate2560(.a(gate20inter10), .b(gate20inter9), .O(gate20inter11));
  nor2  gate2561(.a(gate20inter11), .b(gate20inter6), .O(gate20inter12));
  nand2 gate2562(.a(gate20inter12), .b(gate20inter1), .O(G299));

  xor2  gate2171(.a(G26), .b(G25), .O(gate21inter0));
  nand2 gate2172(.a(gate21inter0), .b(s_232), .O(gate21inter1));
  and2  gate2173(.a(G26), .b(G25), .O(gate21inter2));
  inv1  gate2174(.a(s_232), .O(gate21inter3));
  inv1  gate2175(.a(s_233), .O(gate21inter4));
  nand2 gate2176(.a(gate21inter4), .b(gate21inter3), .O(gate21inter5));
  nor2  gate2177(.a(gate21inter5), .b(gate21inter2), .O(gate21inter6));
  inv1  gate2178(.a(G25), .O(gate21inter7));
  inv1  gate2179(.a(G26), .O(gate21inter8));
  nand2 gate2180(.a(gate21inter8), .b(gate21inter7), .O(gate21inter9));
  nand2 gate2181(.a(s_233), .b(gate21inter3), .O(gate21inter10));
  nor2  gate2182(.a(gate21inter10), .b(gate21inter9), .O(gate21inter11));
  nor2  gate2183(.a(gate21inter11), .b(gate21inter6), .O(gate21inter12));
  nand2 gate2184(.a(gate21inter12), .b(gate21inter1), .O(G302));

  xor2  gate1135(.a(G28), .b(G27), .O(gate22inter0));
  nand2 gate1136(.a(gate22inter0), .b(s_84), .O(gate22inter1));
  and2  gate1137(.a(G28), .b(G27), .O(gate22inter2));
  inv1  gate1138(.a(s_84), .O(gate22inter3));
  inv1  gate1139(.a(s_85), .O(gate22inter4));
  nand2 gate1140(.a(gate22inter4), .b(gate22inter3), .O(gate22inter5));
  nor2  gate1141(.a(gate22inter5), .b(gate22inter2), .O(gate22inter6));
  inv1  gate1142(.a(G27), .O(gate22inter7));
  inv1  gate1143(.a(G28), .O(gate22inter8));
  nand2 gate1144(.a(gate22inter8), .b(gate22inter7), .O(gate22inter9));
  nand2 gate1145(.a(s_85), .b(gate22inter3), .O(gate22inter10));
  nor2  gate1146(.a(gate22inter10), .b(gate22inter9), .O(gate22inter11));
  nor2  gate1147(.a(gate22inter11), .b(gate22inter6), .O(gate22inter12));
  nand2 gate1148(.a(gate22inter12), .b(gate22inter1), .O(G305));

  xor2  gate1569(.a(G30), .b(G29), .O(gate23inter0));
  nand2 gate1570(.a(gate23inter0), .b(s_146), .O(gate23inter1));
  and2  gate1571(.a(G30), .b(G29), .O(gate23inter2));
  inv1  gate1572(.a(s_146), .O(gate23inter3));
  inv1  gate1573(.a(s_147), .O(gate23inter4));
  nand2 gate1574(.a(gate23inter4), .b(gate23inter3), .O(gate23inter5));
  nor2  gate1575(.a(gate23inter5), .b(gate23inter2), .O(gate23inter6));
  inv1  gate1576(.a(G29), .O(gate23inter7));
  inv1  gate1577(.a(G30), .O(gate23inter8));
  nand2 gate1578(.a(gate23inter8), .b(gate23inter7), .O(gate23inter9));
  nand2 gate1579(.a(s_147), .b(gate23inter3), .O(gate23inter10));
  nor2  gate1580(.a(gate23inter10), .b(gate23inter9), .O(gate23inter11));
  nor2  gate1581(.a(gate23inter11), .b(gate23inter6), .O(gate23inter12));
  nand2 gate1582(.a(gate23inter12), .b(gate23inter1), .O(G308));
nand2 gate24( .a(G31), .b(G32), .O(G311) );

  xor2  gate1961(.a(G5), .b(G1), .O(gate25inter0));
  nand2 gate1962(.a(gate25inter0), .b(s_202), .O(gate25inter1));
  and2  gate1963(.a(G5), .b(G1), .O(gate25inter2));
  inv1  gate1964(.a(s_202), .O(gate25inter3));
  inv1  gate1965(.a(s_203), .O(gate25inter4));
  nand2 gate1966(.a(gate25inter4), .b(gate25inter3), .O(gate25inter5));
  nor2  gate1967(.a(gate25inter5), .b(gate25inter2), .O(gate25inter6));
  inv1  gate1968(.a(G1), .O(gate25inter7));
  inv1  gate1969(.a(G5), .O(gate25inter8));
  nand2 gate1970(.a(gate25inter8), .b(gate25inter7), .O(gate25inter9));
  nand2 gate1971(.a(s_203), .b(gate25inter3), .O(gate25inter10));
  nor2  gate1972(.a(gate25inter10), .b(gate25inter9), .O(gate25inter11));
  nor2  gate1973(.a(gate25inter11), .b(gate25inter6), .O(gate25inter12));
  nand2 gate1974(.a(gate25inter12), .b(gate25inter1), .O(G314));
nand2 gate26( .a(G9), .b(G13), .O(G317) );
nand2 gate27( .a(G2), .b(G6), .O(G320) );
nand2 gate28( .a(G10), .b(G14), .O(G323) );
nand2 gate29( .a(G3), .b(G7), .O(G326) );
nand2 gate30( .a(G11), .b(G15), .O(G329) );

  xor2  gate1625(.a(G8), .b(G4), .O(gate31inter0));
  nand2 gate1626(.a(gate31inter0), .b(s_154), .O(gate31inter1));
  and2  gate1627(.a(G8), .b(G4), .O(gate31inter2));
  inv1  gate1628(.a(s_154), .O(gate31inter3));
  inv1  gate1629(.a(s_155), .O(gate31inter4));
  nand2 gate1630(.a(gate31inter4), .b(gate31inter3), .O(gate31inter5));
  nor2  gate1631(.a(gate31inter5), .b(gate31inter2), .O(gate31inter6));
  inv1  gate1632(.a(G4), .O(gate31inter7));
  inv1  gate1633(.a(G8), .O(gate31inter8));
  nand2 gate1634(.a(gate31inter8), .b(gate31inter7), .O(gate31inter9));
  nand2 gate1635(.a(s_155), .b(gate31inter3), .O(gate31inter10));
  nor2  gate1636(.a(gate31inter10), .b(gate31inter9), .O(gate31inter11));
  nor2  gate1637(.a(gate31inter11), .b(gate31inter6), .O(gate31inter12));
  nand2 gate1638(.a(gate31inter12), .b(gate31inter1), .O(G332));

  xor2  gate2031(.a(G16), .b(G12), .O(gate32inter0));
  nand2 gate2032(.a(gate32inter0), .b(s_212), .O(gate32inter1));
  and2  gate2033(.a(G16), .b(G12), .O(gate32inter2));
  inv1  gate2034(.a(s_212), .O(gate32inter3));
  inv1  gate2035(.a(s_213), .O(gate32inter4));
  nand2 gate2036(.a(gate32inter4), .b(gate32inter3), .O(gate32inter5));
  nor2  gate2037(.a(gate32inter5), .b(gate32inter2), .O(gate32inter6));
  inv1  gate2038(.a(G12), .O(gate32inter7));
  inv1  gate2039(.a(G16), .O(gate32inter8));
  nand2 gate2040(.a(gate32inter8), .b(gate32inter7), .O(gate32inter9));
  nand2 gate2041(.a(s_213), .b(gate32inter3), .O(gate32inter10));
  nor2  gate2042(.a(gate32inter10), .b(gate32inter9), .O(gate32inter11));
  nor2  gate2043(.a(gate32inter11), .b(gate32inter6), .O(gate32inter12));
  nand2 gate2044(.a(gate32inter12), .b(gate32inter1), .O(G335));
nand2 gate33( .a(G17), .b(G21), .O(G338) );
nand2 gate34( .a(G25), .b(G29), .O(G341) );
nand2 gate35( .a(G18), .b(G22), .O(G344) );

  xor2  gate659(.a(G30), .b(G26), .O(gate36inter0));
  nand2 gate660(.a(gate36inter0), .b(s_16), .O(gate36inter1));
  and2  gate661(.a(G30), .b(G26), .O(gate36inter2));
  inv1  gate662(.a(s_16), .O(gate36inter3));
  inv1  gate663(.a(s_17), .O(gate36inter4));
  nand2 gate664(.a(gate36inter4), .b(gate36inter3), .O(gate36inter5));
  nor2  gate665(.a(gate36inter5), .b(gate36inter2), .O(gate36inter6));
  inv1  gate666(.a(G26), .O(gate36inter7));
  inv1  gate667(.a(G30), .O(gate36inter8));
  nand2 gate668(.a(gate36inter8), .b(gate36inter7), .O(gate36inter9));
  nand2 gate669(.a(s_17), .b(gate36inter3), .O(gate36inter10));
  nor2  gate670(.a(gate36inter10), .b(gate36inter9), .O(gate36inter11));
  nor2  gate671(.a(gate36inter11), .b(gate36inter6), .O(gate36inter12));
  nand2 gate672(.a(gate36inter12), .b(gate36inter1), .O(G347));
nand2 gate37( .a(G19), .b(G23), .O(G350) );
nand2 gate38( .a(G27), .b(G31), .O(G353) );
nand2 gate39( .a(G20), .b(G24), .O(G356) );
nand2 gate40( .a(G28), .b(G32), .O(G359) );

  xor2  gate631(.a(G266), .b(G1), .O(gate41inter0));
  nand2 gate632(.a(gate41inter0), .b(s_12), .O(gate41inter1));
  and2  gate633(.a(G266), .b(G1), .O(gate41inter2));
  inv1  gate634(.a(s_12), .O(gate41inter3));
  inv1  gate635(.a(s_13), .O(gate41inter4));
  nand2 gate636(.a(gate41inter4), .b(gate41inter3), .O(gate41inter5));
  nor2  gate637(.a(gate41inter5), .b(gate41inter2), .O(gate41inter6));
  inv1  gate638(.a(G1), .O(gate41inter7));
  inv1  gate639(.a(G266), .O(gate41inter8));
  nand2 gate640(.a(gate41inter8), .b(gate41inter7), .O(gate41inter9));
  nand2 gate641(.a(s_13), .b(gate41inter3), .O(gate41inter10));
  nor2  gate642(.a(gate41inter10), .b(gate41inter9), .O(gate41inter11));
  nor2  gate643(.a(gate41inter11), .b(gate41inter6), .O(gate41inter12));
  nand2 gate644(.a(gate41inter12), .b(gate41inter1), .O(G362));
nand2 gate42( .a(G2), .b(G266), .O(G363) );
nand2 gate43( .a(G3), .b(G269), .O(G364) );
nand2 gate44( .a(G4), .b(G269), .O(G365) );
nand2 gate45( .a(G5), .b(G272), .O(G366) );
nand2 gate46( .a(G6), .b(G272), .O(G367) );

  xor2  gate715(.a(G275), .b(G7), .O(gate47inter0));
  nand2 gate716(.a(gate47inter0), .b(s_24), .O(gate47inter1));
  and2  gate717(.a(G275), .b(G7), .O(gate47inter2));
  inv1  gate718(.a(s_24), .O(gate47inter3));
  inv1  gate719(.a(s_25), .O(gate47inter4));
  nand2 gate720(.a(gate47inter4), .b(gate47inter3), .O(gate47inter5));
  nor2  gate721(.a(gate47inter5), .b(gate47inter2), .O(gate47inter6));
  inv1  gate722(.a(G7), .O(gate47inter7));
  inv1  gate723(.a(G275), .O(gate47inter8));
  nand2 gate724(.a(gate47inter8), .b(gate47inter7), .O(gate47inter9));
  nand2 gate725(.a(s_25), .b(gate47inter3), .O(gate47inter10));
  nor2  gate726(.a(gate47inter10), .b(gate47inter9), .O(gate47inter11));
  nor2  gate727(.a(gate47inter11), .b(gate47inter6), .O(gate47inter12));
  nand2 gate728(.a(gate47inter12), .b(gate47inter1), .O(G368));
nand2 gate48( .a(G8), .b(G275), .O(G369) );
nand2 gate49( .a(G9), .b(G278), .O(G370) );
nand2 gate50( .a(G10), .b(G278), .O(G371) );
nand2 gate51( .a(G11), .b(G281), .O(G372) );
nand2 gate52( .a(G12), .b(G281), .O(G373) );

  xor2  gate2325(.a(G284), .b(G13), .O(gate53inter0));
  nand2 gate2326(.a(gate53inter0), .b(s_254), .O(gate53inter1));
  and2  gate2327(.a(G284), .b(G13), .O(gate53inter2));
  inv1  gate2328(.a(s_254), .O(gate53inter3));
  inv1  gate2329(.a(s_255), .O(gate53inter4));
  nand2 gate2330(.a(gate53inter4), .b(gate53inter3), .O(gate53inter5));
  nor2  gate2331(.a(gate53inter5), .b(gate53inter2), .O(gate53inter6));
  inv1  gate2332(.a(G13), .O(gate53inter7));
  inv1  gate2333(.a(G284), .O(gate53inter8));
  nand2 gate2334(.a(gate53inter8), .b(gate53inter7), .O(gate53inter9));
  nand2 gate2335(.a(s_255), .b(gate53inter3), .O(gate53inter10));
  nor2  gate2336(.a(gate53inter10), .b(gate53inter9), .O(gate53inter11));
  nor2  gate2337(.a(gate53inter11), .b(gate53inter6), .O(gate53inter12));
  nand2 gate2338(.a(gate53inter12), .b(gate53inter1), .O(G374));

  xor2  gate1499(.a(G284), .b(G14), .O(gate54inter0));
  nand2 gate1500(.a(gate54inter0), .b(s_136), .O(gate54inter1));
  and2  gate1501(.a(G284), .b(G14), .O(gate54inter2));
  inv1  gate1502(.a(s_136), .O(gate54inter3));
  inv1  gate1503(.a(s_137), .O(gate54inter4));
  nand2 gate1504(.a(gate54inter4), .b(gate54inter3), .O(gate54inter5));
  nor2  gate1505(.a(gate54inter5), .b(gate54inter2), .O(gate54inter6));
  inv1  gate1506(.a(G14), .O(gate54inter7));
  inv1  gate1507(.a(G284), .O(gate54inter8));
  nand2 gate1508(.a(gate54inter8), .b(gate54inter7), .O(gate54inter9));
  nand2 gate1509(.a(s_137), .b(gate54inter3), .O(gate54inter10));
  nor2  gate1510(.a(gate54inter10), .b(gate54inter9), .O(gate54inter11));
  nor2  gate1511(.a(gate54inter11), .b(gate54inter6), .O(gate54inter12));
  nand2 gate1512(.a(gate54inter12), .b(gate54inter1), .O(G375));
nand2 gate55( .a(G15), .b(G287), .O(G376) );

  xor2  gate2661(.a(G287), .b(G16), .O(gate56inter0));
  nand2 gate2662(.a(gate56inter0), .b(s_302), .O(gate56inter1));
  and2  gate2663(.a(G287), .b(G16), .O(gate56inter2));
  inv1  gate2664(.a(s_302), .O(gate56inter3));
  inv1  gate2665(.a(s_303), .O(gate56inter4));
  nand2 gate2666(.a(gate56inter4), .b(gate56inter3), .O(gate56inter5));
  nor2  gate2667(.a(gate56inter5), .b(gate56inter2), .O(gate56inter6));
  inv1  gate2668(.a(G16), .O(gate56inter7));
  inv1  gate2669(.a(G287), .O(gate56inter8));
  nand2 gate2670(.a(gate56inter8), .b(gate56inter7), .O(gate56inter9));
  nand2 gate2671(.a(s_303), .b(gate56inter3), .O(gate56inter10));
  nor2  gate2672(.a(gate56inter10), .b(gate56inter9), .O(gate56inter11));
  nor2  gate2673(.a(gate56inter11), .b(gate56inter6), .O(gate56inter12));
  nand2 gate2674(.a(gate56inter12), .b(gate56inter1), .O(G377));
nand2 gate57( .a(G17), .b(G290), .O(G378) );

  xor2  gate1541(.a(G290), .b(G18), .O(gate58inter0));
  nand2 gate1542(.a(gate58inter0), .b(s_142), .O(gate58inter1));
  and2  gate1543(.a(G290), .b(G18), .O(gate58inter2));
  inv1  gate1544(.a(s_142), .O(gate58inter3));
  inv1  gate1545(.a(s_143), .O(gate58inter4));
  nand2 gate1546(.a(gate58inter4), .b(gate58inter3), .O(gate58inter5));
  nor2  gate1547(.a(gate58inter5), .b(gate58inter2), .O(gate58inter6));
  inv1  gate1548(.a(G18), .O(gate58inter7));
  inv1  gate1549(.a(G290), .O(gate58inter8));
  nand2 gate1550(.a(gate58inter8), .b(gate58inter7), .O(gate58inter9));
  nand2 gate1551(.a(s_143), .b(gate58inter3), .O(gate58inter10));
  nor2  gate1552(.a(gate58inter10), .b(gate58inter9), .O(gate58inter11));
  nor2  gate1553(.a(gate58inter11), .b(gate58inter6), .O(gate58inter12));
  nand2 gate1554(.a(gate58inter12), .b(gate58inter1), .O(G379));

  xor2  gate1163(.a(G293), .b(G19), .O(gate59inter0));
  nand2 gate1164(.a(gate59inter0), .b(s_88), .O(gate59inter1));
  and2  gate1165(.a(G293), .b(G19), .O(gate59inter2));
  inv1  gate1166(.a(s_88), .O(gate59inter3));
  inv1  gate1167(.a(s_89), .O(gate59inter4));
  nand2 gate1168(.a(gate59inter4), .b(gate59inter3), .O(gate59inter5));
  nor2  gate1169(.a(gate59inter5), .b(gate59inter2), .O(gate59inter6));
  inv1  gate1170(.a(G19), .O(gate59inter7));
  inv1  gate1171(.a(G293), .O(gate59inter8));
  nand2 gate1172(.a(gate59inter8), .b(gate59inter7), .O(gate59inter9));
  nand2 gate1173(.a(s_89), .b(gate59inter3), .O(gate59inter10));
  nor2  gate1174(.a(gate59inter10), .b(gate59inter9), .O(gate59inter11));
  nor2  gate1175(.a(gate59inter11), .b(gate59inter6), .O(gate59inter12));
  nand2 gate1176(.a(gate59inter12), .b(gate59inter1), .O(G380));

  xor2  gate1555(.a(G293), .b(G20), .O(gate60inter0));
  nand2 gate1556(.a(gate60inter0), .b(s_144), .O(gate60inter1));
  and2  gate1557(.a(G293), .b(G20), .O(gate60inter2));
  inv1  gate1558(.a(s_144), .O(gate60inter3));
  inv1  gate1559(.a(s_145), .O(gate60inter4));
  nand2 gate1560(.a(gate60inter4), .b(gate60inter3), .O(gate60inter5));
  nor2  gate1561(.a(gate60inter5), .b(gate60inter2), .O(gate60inter6));
  inv1  gate1562(.a(G20), .O(gate60inter7));
  inv1  gate1563(.a(G293), .O(gate60inter8));
  nand2 gate1564(.a(gate60inter8), .b(gate60inter7), .O(gate60inter9));
  nand2 gate1565(.a(s_145), .b(gate60inter3), .O(gate60inter10));
  nor2  gate1566(.a(gate60inter10), .b(gate60inter9), .O(gate60inter11));
  nor2  gate1567(.a(gate60inter11), .b(gate60inter6), .O(gate60inter12));
  nand2 gate1568(.a(gate60inter12), .b(gate60inter1), .O(G381));
nand2 gate61( .a(G21), .b(G296), .O(G382) );
nand2 gate62( .a(G22), .b(G296), .O(G383) );

  xor2  gate617(.a(G299), .b(G23), .O(gate63inter0));
  nand2 gate618(.a(gate63inter0), .b(s_10), .O(gate63inter1));
  and2  gate619(.a(G299), .b(G23), .O(gate63inter2));
  inv1  gate620(.a(s_10), .O(gate63inter3));
  inv1  gate621(.a(s_11), .O(gate63inter4));
  nand2 gate622(.a(gate63inter4), .b(gate63inter3), .O(gate63inter5));
  nor2  gate623(.a(gate63inter5), .b(gate63inter2), .O(gate63inter6));
  inv1  gate624(.a(G23), .O(gate63inter7));
  inv1  gate625(.a(G299), .O(gate63inter8));
  nand2 gate626(.a(gate63inter8), .b(gate63inter7), .O(gate63inter9));
  nand2 gate627(.a(s_11), .b(gate63inter3), .O(gate63inter10));
  nor2  gate628(.a(gate63inter10), .b(gate63inter9), .O(gate63inter11));
  nor2  gate629(.a(gate63inter11), .b(gate63inter6), .O(gate63inter12));
  nand2 gate630(.a(gate63inter12), .b(gate63inter1), .O(G384));
nand2 gate64( .a(G24), .b(G299), .O(G385) );

  xor2  gate687(.a(G302), .b(G25), .O(gate65inter0));
  nand2 gate688(.a(gate65inter0), .b(s_20), .O(gate65inter1));
  and2  gate689(.a(G302), .b(G25), .O(gate65inter2));
  inv1  gate690(.a(s_20), .O(gate65inter3));
  inv1  gate691(.a(s_21), .O(gate65inter4));
  nand2 gate692(.a(gate65inter4), .b(gate65inter3), .O(gate65inter5));
  nor2  gate693(.a(gate65inter5), .b(gate65inter2), .O(gate65inter6));
  inv1  gate694(.a(G25), .O(gate65inter7));
  inv1  gate695(.a(G302), .O(gate65inter8));
  nand2 gate696(.a(gate65inter8), .b(gate65inter7), .O(gate65inter9));
  nand2 gate697(.a(s_21), .b(gate65inter3), .O(gate65inter10));
  nor2  gate698(.a(gate65inter10), .b(gate65inter9), .O(gate65inter11));
  nor2  gate699(.a(gate65inter11), .b(gate65inter6), .O(gate65inter12));
  nand2 gate700(.a(gate65inter12), .b(gate65inter1), .O(G386));
nand2 gate66( .a(G26), .b(G302), .O(G387) );
nand2 gate67( .a(G27), .b(G305), .O(G388) );
nand2 gate68( .a(G28), .b(G305), .O(G389) );
nand2 gate69( .a(G29), .b(G308), .O(G390) );
nand2 gate70( .a(G30), .b(G308), .O(G391) );
nand2 gate71( .a(G31), .b(G311), .O(G392) );
nand2 gate72( .a(G32), .b(G311), .O(G393) );

  xor2  gate1275(.a(G314), .b(G1), .O(gate73inter0));
  nand2 gate1276(.a(gate73inter0), .b(s_104), .O(gate73inter1));
  and2  gate1277(.a(G314), .b(G1), .O(gate73inter2));
  inv1  gate1278(.a(s_104), .O(gate73inter3));
  inv1  gate1279(.a(s_105), .O(gate73inter4));
  nand2 gate1280(.a(gate73inter4), .b(gate73inter3), .O(gate73inter5));
  nor2  gate1281(.a(gate73inter5), .b(gate73inter2), .O(gate73inter6));
  inv1  gate1282(.a(G1), .O(gate73inter7));
  inv1  gate1283(.a(G314), .O(gate73inter8));
  nand2 gate1284(.a(gate73inter8), .b(gate73inter7), .O(gate73inter9));
  nand2 gate1285(.a(s_105), .b(gate73inter3), .O(gate73inter10));
  nor2  gate1286(.a(gate73inter10), .b(gate73inter9), .O(gate73inter11));
  nor2  gate1287(.a(gate73inter11), .b(gate73inter6), .O(gate73inter12));
  nand2 gate1288(.a(gate73inter12), .b(gate73inter1), .O(G394));
nand2 gate74( .a(G5), .b(G314), .O(G395) );
nand2 gate75( .a(G9), .b(G317), .O(G396) );

  xor2  gate603(.a(G317), .b(G13), .O(gate76inter0));
  nand2 gate604(.a(gate76inter0), .b(s_8), .O(gate76inter1));
  and2  gate605(.a(G317), .b(G13), .O(gate76inter2));
  inv1  gate606(.a(s_8), .O(gate76inter3));
  inv1  gate607(.a(s_9), .O(gate76inter4));
  nand2 gate608(.a(gate76inter4), .b(gate76inter3), .O(gate76inter5));
  nor2  gate609(.a(gate76inter5), .b(gate76inter2), .O(gate76inter6));
  inv1  gate610(.a(G13), .O(gate76inter7));
  inv1  gate611(.a(G317), .O(gate76inter8));
  nand2 gate612(.a(gate76inter8), .b(gate76inter7), .O(gate76inter9));
  nand2 gate613(.a(s_9), .b(gate76inter3), .O(gate76inter10));
  nor2  gate614(.a(gate76inter10), .b(gate76inter9), .O(gate76inter11));
  nor2  gate615(.a(gate76inter11), .b(gate76inter6), .O(gate76inter12));
  nand2 gate616(.a(gate76inter12), .b(gate76inter1), .O(G397));

  xor2  gate1457(.a(G320), .b(G2), .O(gate77inter0));
  nand2 gate1458(.a(gate77inter0), .b(s_130), .O(gate77inter1));
  and2  gate1459(.a(G320), .b(G2), .O(gate77inter2));
  inv1  gate1460(.a(s_130), .O(gate77inter3));
  inv1  gate1461(.a(s_131), .O(gate77inter4));
  nand2 gate1462(.a(gate77inter4), .b(gate77inter3), .O(gate77inter5));
  nor2  gate1463(.a(gate77inter5), .b(gate77inter2), .O(gate77inter6));
  inv1  gate1464(.a(G2), .O(gate77inter7));
  inv1  gate1465(.a(G320), .O(gate77inter8));
  nand2 gate1466(.a(gate77inter8), .b(gate77inter7), .O(gate77inter9));
  nand2 gate1467(.a(s_131), .b(gate77inter3), .O(gate77inter10));
  nor2  gate1468(.a(gate77inter10), .b(gate77inter9), .O(gate77inter11));
  nor2  gate1469(.a(gate77inter11), .b(gate77inter6), .O(gate77inter12));
  nand2 gate1470(.a(gate77inter12), .b(gate77inter1), .O(G398));
nand2 gate78( .a(G6), .b(G320), .O(G399) );
nand2 gate79( .a(G10), .b(G323), .O(G400) );
nand2 gate80( .a(G14), .b(G323), .O(G401) );

  xor2  gate1373(.a(G326), .b(G3), .O(gate81inter0));
  nand2 gate1374(.a(gate81inter0), .b(s_118), .O(gate81inter1));
  and2  gate1375(.a(G326), .b(G3), .O(gate81inter2));
  inv1  gate1376(.a(s_118), .O(gate81inter3));
  inv1  gate1377(.a(s_119), .O(gate81inter4));
  nand2 gate1378(.a(gate81inter4), .b(gate81inter3), .O(gate81inter5));
  nor2  gate1379(.a(gate81inter5), .b(gate81inter2), .O(gate81inter6));
  inv1  gate1380(.a(G3), .O(gate81inter7));
  inv1  gate1381(.a(G326), .O(gate81inter8));
  nand2 gate1382(.a(gate81inter8), .b(gate81inter7), .O(gate81inter9));
  nand2 gate1383(.a(s_119), .b(gate81inter3), .O(gate81inter10));
  nor2  gate1384(.a(gate81inter10), .b(gate81inter9), .O(gate81inter11));
  nor2  gate1385(.a(gate81inter11), .b(gate81inter6), .O(gate81inter12));
  nand2 gate1386(.a(gate81inter12), .b(gate81inter1), .O(G402));

  xor2  gate2101(.a(G326), .b(G7), .O(gate82inter0));
  nand2 gate2102(.a(gate82inter0), .b(s_222), .O(gate82inter1));
  and2  gate2103(.a(G326), .b(G7), .O(gate82inter2));
  inv1  gate2104(.a(s_222), .O(gate82inter3));
  inv1  gate2105(.a(s_223), .O(gate82inter4));
  nand2 gate2106(.a(gate82inter4), .b(gate82inter3), .O(gate82inter5));
  nor2  gate2107(.a(gate82inter5), .b(gate82inter2), .O(gate82inter6));
  inv1  gate2108(.a(G7), .O(gate82inter7));
  inv1  gate2109(.a(G326), .O(gate82inter8));
  nand2 gate2110(.a(gate82inter8), .b(gate82inter7), .O(gate82inter9));
  nand2 gate2111(.a(s_223), .b(gate82inter3), .O(gate82inter10));
  nor2  gate2112(.a(gate82inter10), .b(gate82inter9), .O(gate82inter11));
  nor2  gate2113(.a(gate82inter11), .b(gate82inter6), .O(gate82inter12));
  nand2 gate2114(.a(gate82inter12), .b(gate82inter1), .O(G403));
nand2 gate83( .a(G11), .b(G329), .O(G404) );
nand2 gate84( .a(G15), .b(G329), .O(G405) );
nand2 gate85( .a(G4), .b(G332), .O(G406) );

  xor2  gate841(.a(G332), .b(G8), .O(gate86inter0));
  nand2 gate842(.a(gate86inter0), .b(s_42), .O(gate86inter1));
  and2  gate843(.a(G332), .b(G8), .O(gate86inter2));
  inv1  gate844(.a(s_42), .O(gate86inter3));
  inv1  gate845(.a(s_43), .O(gate86inter4));
  nand2 gate846(.a(gate86inter4), .b(gate86inter3), .O(gate86inter5));
  nor2  gate847(.a(gate86inter5), .b(gate86inter2), .O(gate86inter6));
  inv1  gate848(.a(G8), .O(gate86inter7));
  inv1  gate849(.a(G332), .O(gate86inter8));
  nand2 gate850(.a(gate86inter8), .b(gate86inter7), .O(gate86inter9));
  nand2 gate851(.a(s_43), .b(gate86inter3), .O(gate86inter10));
  nor2  gate852(.a(gate86inter10), .b(gate86inter9), .O(gate86inter11));
  nor2  gate853(.a(gate86inter11), .b(gate86inter6), .O(gate86inter12));
  nand2 gate854(.a(gate86inter12), .b(gate86inter1), .O(G407));

  xor2  gate2451(.a(G335), .b(G12), .O(gate87inter0));
  nand2 gate2452(.a(gate87inter0), .b(s_272), .O(gate87inter1));
  and2  gate2453(.a(G335), .b(G12), .O(gate87inter2));
  inv1  gate2454(.a(s_272), .O(gate87inter3));
  inv1  gate2455(.a(s_273), .O(gate87inter4));
  nand2 gate2456(.a(gate87inter4), .b(gate87inter3), .O(gate87inter5));
  nor2  gate2457(.a(gate87inter5), .b(gate87inter2), .O(gate87inter6));
  inv1  gate2458(.a(G12), .O(gate87inter7));
  inv1  gate2459(.a(G335), .O(gate87inter8));
  nand2 gate2460(.a(gate87inter8), .b(gate87inter7), .O(gate87inter9));
  nand2 gate2461(.a(s_273), .b(gate87inter3), .O(gate87inter10));
  nor2  gate2462(.a(gate87inter10), .b(gate87inter9), .O(gate87inter11));
  nor2  gate2463(.a(gate87inter11), .b(gate87inter6), .O(gate87inter12));
  nand2 gate2464(.a(gate87inter12), .b(gate87inter1), .O(G408));
nand2 gate88( .a(G16), .b(G335), .O(G409) );

  xor2  gate2297(.a(G338), .b(G17), .O(gate89inter0));
  nand2 gate2298(.a(gate89inter0), .b(s_250), .O(gate89inter1));
  and2  gate2299(.a(G338), .b(G17), .O(gate89inter2));
  inv1  gate2300(.a(s_250), .O(gate89inter3));
  inv1  gate2301(.a(s_251), .O(gate89inter4));
  nand2 gate2302(.a(gate89inter4), .b(gate89inter3), .O(gate89inter5));
  nor2  gate2303(.a(gate89inter5), .b(gate89inter2), .O(gate89inter6));
  inv1  gate2304(.a(G17), .O(gate89inter7));
  inv1  gate2305(.a(G338), .O(gate89inter8));
  nand2 gate2306(.a(gate89inter8), .b(gate89inter7), .O(gate89inter9));
  nand2 gate2307(.a(s_251), .b(gate89inter3), .O(gate89inter10));
  nor2  gate2308(.a(gate89inter10), .b(gate89inter9), .O(gate89inter11));
  nor2  gate2309(.a(gate89inter11), .b(gate89inter6), .O(gate89inter12));
  nand2 gate2310(.a(gate89inter12), .b(gate89inter1), .O(G410));
nand2 gate90( .a(G21), .b(G338), .O(G411) );
nand2 gate91( .a(G25), .b(G341), .O(G412) );

  xor2  gate1723(.a(G341), .b(G29), .O(gate92inter0));
  nand2 gate1724(.a(gate92inter0), .b(s_168), .O(gate92inter1));
  and2  gate1725(.a(G341), .b(G29), .O(gate92inter2));
  inv1  gate1726(.a(s_168), .O(gate92inter3));
  inv1  gate1727(.a(s_169), .O(gate92inter4));
  nand2 gate1728(.a(gate92inter4), .b(gate92inter3), .O(gate92inter5));
  nor2  gate1729(.a(gate92inter5), .b(gate92inter2), .O(gate92inter6));
  inv1  gate1730(.a(G29), .O(gate92inter7));
  inv1  gate1731(.a(G341), .O(gate92inter8));
  nand2 gate1732(.a(gate92inter8), .b(gate92inter7), .O(gate92inter9));
  nand2 gate1733(.a(s_169), .b(gate92inter3), .O(gate92inter10));
  nor2  gate1734(.a(gate92inter10), .b(gate92inter9), .O(gate92inter11));
  nor2  gate1735(.a(gate92inter11), .b(gate92inter6), .O(gate92inter12));
  nand2 gate1736(.a(gate92inter12), .b(gate92inter1), .O(G413));
nand2 gate93( .a(G18), .b(G344), .O(G414) );
nand2 gate94( .a(G22), .b(G344), .O(G415) );
nand2 gate95( .a(G26), .b(G347), .O(G416) );

  xor2  gate575(.a(G347), .b(G30), .O(gate96inter0));
  nand2 gate576(.a(gate96inter0), .b(s_4), .O(gate96inter1));
  and2  gate577(.a(G347), .b(G30), .O(gate96inter2));
  inv1  gate578(.a(s_4), .O(gate96inter3));
  inv1  gate579(.a(s_5), .O(gate96inter4));
  nand2 gate580(.a(gate96inter4), .b(gate96inter3), .O(gate96inter5));
  nor2  gate581(.a(gate96inter5), .b(gate96inter2), .O(gate96inter6));
  inv1  gate582(.a(G30), .O(gate96inter7));
  inv1  gate583(.a(G347), .O(gate96inter8));
  nand2 gate584(.a(gate96inter8), .b(gate96inter7), .O(gate96inter9));
  nand2 gate585(.a(s_5), .b(gate96inter3), .O(gate96inter10));
  nor2  gate586(.a(gate96inter10), .b(gate96inter9), .O(gate96inter11));
  nor2  gate587(.a(gate96inter11), .b(gate96inter6), .O(gate96inter12));
  nand2 gate588(.a(gate96inter12), .b(gate96inter1), .O(G417));
nand2 gate97( .a(G19), .b(G350), .O(G418) );

  xor2  gate967(.a(G350), .b(G23), .O(gate98inter0));
  nand2 gate968(.a(gate98inter0), .b(s_60), .O(gate98inter1));
  and2  gate969(.a(G350), .b(G23), .O(gate98inter2));
  inv1  gate970(.a(s_60), .O(gate98inter3));
  inv1  gate971(.a(s_61), .O(gate98inter4));
  nand2 gate972(.a(gate98inter4), .b(gate98inter3), .O(gate98inter5));
  nor2  gate973(.a(gate98inter5), .b(gate98inter2), .O(gate98inter6));
  inv1  gate974(.a(G23), .O(gate98inter7));
  inv1  gate975(.a(G350), .O(gate98inter8));
  nand2 gate976(.a(gate98inter8), .b(gate98inter7), .O(gate98inter9));
  nand2 gate977(.a(s_61), .b(gate98inter3), .O(gate98inter10));
  nor2  gate978(.a(gate98inter10), .b(gate98inter9), .O(gate98inter11));
  nor2  gate979(.a(gate98inter11), .b(gate98inter6), .O(gate98inter12));
  nand2 gate980(.a(gate98inter12), .b(gate98inter1), .O(G419));
nand2 gate99( .a(G27), .b(G353), .O(G420) );
nand2 gate100( .a(G31), .b(G353), .O(G421) );
nand2 gate101( .a(G20), .b(G356), .O(G422) );

  xor2  gate2003(.a(G356), .b(G24), .O(gate102inter0));
  nand2 gate2004(.a(gate102inter0), .b(s_208), .O(gate102inter1));
  and2  gate2005(.a(G356), .b(G24), .O(gate102inter2));
  inv1  gate2006(.a(s_208), .O(gate102inter3));
  inv1  gate2007(.a(s_209), .O(gate102inter4));
  nand2 gate2008(.a(gate102inter4), .b(gate102inter3), .O(gate102inter5));
  nor2  gate2009(.a(gate102inter5), .b(gate102inter2), .O(gate102inter6));
  inv1  gate2010(.a(G24), .O(gate102inter7));
  inv1  gate2011(.a(G356), .O(gate102inter8));
  nand2 gate2012(.a(gate102inter8), .b(gate102inter7), .O(gate102inter9));
  nand2 gate2013(.a(s_209), .b(gate102inter3), .O(gate102inter10));
  nor2  gate2014(.a(gate102inter10), .b(gate102inter9), .O(gate102inter11));
  nor2  gate2015(.a(gate102inter11), .b(gate102inter6), .O(gate102inter12));
  nand2 gate2016(.a(gate102inter12), .b(gate102inter1), .O(G423));
nand2 gate103( .a(G28), .b(G359), .O(G424) );

  xor2  gate1583(.a(G359), .b(G32), .O(gate104inter0));
  nand2 gate1584(.a(gate104inter0), .b(s_148), .O(gate104inter1));
  and2  gate1585(.a(G359), .b(G32), .O(gate104inter2));
  inv1  gate1586(.a(s_148), .O(gate104inter3));
  inv1  gate1587(.a(s_149), .O(gate104inter4));
  nand2 gate1588(.a(gate104inter4), .b(gate104inter3), .O(gate104inter5));
  nor2  gate1589(.a(gate104inter5), .b(gate104inter2), .O(gate104inter6));
  inv1  gate1590(.a(G32), .O(gate104inter7));
  inv1  gate1591(.a(G359), .O(gate104inter8));
  nand2 gate1592(.a(gate104inter8), .b(gate104inter7), .O(gate104inter9));
  nand2 gate1593(.a(s_149), .b(gate104inter3), .O(gate104inter10));
  nor2  gate1594(.a(gate104inter10), .b(gate104inter9), .O(gate104inter11));
  nor2  gate1595(.a(gate104inter11), .b(gate104inter6), .O(gate104inter12));
  nand2 gate1596(.a(gate104inter12), .b(gate104inter1), .O(G425));
nand2 gate105( .a(G362), .b(G363), .O(G426) );
nand2 gate106( .a(G364), .b(G365), .O(G429) );

  xor2  gate1737(.a(G367), .b(G366), .O(gate107inter0));
  nand2 gate1738(.a(gate107inter0), .b(s_170), .O(gate107inter1));
  and2  gate1739(.a(G367), .b(G366), .O(gate107inter2));
  inv1  gate1740(.a(s_170), .O(gate107inter3));
  inv1  gate1741(.a(s_171), .O(gate107inter4));
  nand2 gate1742(.a(gate107inter4), .b(gate107inter3), .O(gate107inter5));
  nor2  gate1743(.a(gate107inter5), .b(gate107inter2), .O(gate107inter6));
  inv1  gate1744(.a(G366), .O(gate107inter7));
  inv1  gate1745(.a(G367), .O(gate107inter8));
  nand2 gate1746(.a(gate107inter8), .b(gate107inter7), .O(gate107inter9));
  nand2 gate1747(.a(s_171), .b(gate107inter3), .O(gate107inter10));
  nor2  gate1748(.a(gate107inter10), .b(gate107inter9), .O(gate107inter11));
  nor2  gate1749(.a(gate107inter11), .b(gate107inter6), .O(gate107inter12));
  nand2 gate1750(.a(gate107inter12), .b(gate107inter1), .O(G432));
nand2 gate108( .a(G368), .b(G369), .O(G435) );

  xor2  gate2689(.a(G371), .b(G370), .O(gate109inter0));
  nand2 gate2690(.a(gate109inter0), .b(s_306), .O(gate109inter1));
  and2  gate2691(.a(G371), .b(G370), .O(gate109inter2));
  inv1  gate2692(.a(s_306), .O(gate109inter3));
  inv1  gate2693(.a(s_307), .O(gate109inter4));
  nand2 gate2694(.a(gate109inter4), .b(gate109inter3), .O(gate109inter5));
  nor2  gate2695(.a(gate109inter5), .b(gate109inter2), .O(gate109inter6));
  inv1  gate2696(.a(G370), .O(gate109inter7));
  inv1  gate2697(.a(G371), .O(gate109inter8));
  nand2 gate2698(.a(gate109inter8), .b(gate109inter7), .O(gate109inter9));
  nand2 gate2699(.a(s_307), .b(gate109inter3), .O(gate109inter10));
  nor2  gate2700(.a(gate109inter10), .b(gate109inter9), .O(gate109inter11));
  nor2  gate2701(.a(gate109inter11), .b(gate109inter6), .O(gate109inter12));
  nand2 gate2702(.a(gate109inter12), .b(gate109inter1), .O(G438));
nand2 gate110( .a(G372), .b(G373), .O(G441) );

  xor2  gate1639(.a(G375), .b(G374), .O(gate111inter0));
  nand2 gate1640(.a(gate111inter0), .b(s_156), .O(gate111inter1));
  and2  gate1641(.a(G375), .b(G374), .O(gate111inter2));
  inv1  gate1642(.a(s_156), .O(gate111inter3));
  inv1  gate1643(.a(s_157), .O(gate111inter4));
  nand2 gate1644(.a(gate111inter4), .b(gate111inter3), .O(gate111inter5));
  nor2  gate1645(.a(gate111inter5), .b(gate111inter2), .O(gate111inter6));
  inv1  gate1646(.a(G374), .O(gate111inter7));
  inv1  gate1647(.a(G375), .O(gate111inter8));
  nand2 gate1648(.a(gate111inter8), .b(gate111inter7), .O(gate111inter9));
  nand2 gate1649(.a(s_157), .b(gate111inter3), .O(gate111inter10));
  nor2  gate1650(.a(gate111inter10), .b(gate111inter9), .O(gate111inter11));
  nor2  gate1651(.a(gate111inter11), .b(gate111inter6), .O(gate111inter12));
  nand2 gate1652(.a(gate111inter12), .b(gate111inter1), .O(G444));
nand2 gate112( .a(G376), .b(G377), .O(G447) );
nand2 gate113( .a(G378), .b(G379), .O(G450) );

  xor2  gate1471(.a(G381), .b(G380), .O(gate114inter0));
  nand2 gate1472(.a(gate114inter0), .b(s_132), .O(gate114inter1));
  and2  gate1473(.a(G381), .b(G380), .O(gate114inter2));
  inv1  gate1474(.a(s_132), .O(gate114inter3));
  inv1  gate1475(.a(s_133), .O(gate114inter4));
  nand2 gate1476(.a(gate114inter4), .b(gate114inter3), .O(gate114inter5));
  nor2  gate1477(.a(gate114inter5), .b(gate114inter2), .O(gate114inter6));
  inv1  gate1478(.a(G380), .O(gate114inter7));
  inv1  gate1479(.a(G381), .O(gate114inter8));
  nand2 gate1480(.a(gate114inter8), .b(gate114inter7), .O(gate114inter9));
  nand2 gate1481(.a(s_133), .b(gate114inter3), .O(gate114inter10));
  nor2  gate1482(.a(gate114inter10), .b(gate114inter9), .O(gate114inter11));
  nor2  gate1483(.a(gate114inter11), .b(gate114inter6), .O(gate114inter12));
  nand2 gate1484(.a(gate114inter12), .b(gate114inter1), .O(G453));
nand2 gate115( .a(G382), .b(G383), .O(G456) );

  xor2  gate2269(.a(G385), .b(G384), .O(gate116inter0));
  nand2 gate2270(.a(gate116inter0), .b(s_246), .O(gate116inter1));
  and2  gate2271(.a(G385), .b(G384), .O(gate116inter2));
  inv1  gate2272(.a(s_246), .O(gate116inter3));
  inv1  gate2273(.a(s_247), .O(gate116inter4));
  nand2 gate2274(.a(gate116inter4), .b(gate116inter3), .O(gate116inter5));
  nor2  gate2275(.a(gate116inter5), .b(gate116inter2), .O(gate116inter6));
  inv1  gate2276(.a(G384), .O(gate116inter7));
  inv1  gate2277(.a(G385), .O(gate116inter8));
  nand2 gate2278(.a(gate116inter8), .b(gate116inter7), .O(gate116inter9));
  nand2 gate2279(.a(s_247), .b(gate116inter3), .O(gate116inter10));
  nor2  gate2280(.a(gate116inter10), .b(gate116inter9), .O(gate116inter11));
  nor2  gate2281(.a(gate116inter11), .b(gate116inter6), .O(gate116inter12));
  nand2 gate2282(.a(gate116inter12), .b(gate116inter1), .O(G459));
nand2 gate117( .a(G386), .b(G387), .O(G462) );
nand2 gate118( .a(G388), .b(G389), .O(G465) );
nand2 gate119( .a(G390), .b(G391), .O(G468) );
nand2 gate120( .a(G392), .b(G393), .O(G471) );

  xor2  gate1429(.a(G395), .b(G394), .O(gate121inter0));
  nand2 gate1430(.a(gate121inter0), .b(s_126), .O(gate121inter1));
  and2  gate1431(.a(G395), .b(G394), .O(gate121inter2));
  inv1  gate1432(.a(s_126), .O(gate121inter3));
  inv1  gate1433(.a(s_127), .O(gate121inter4));
  nand2 gate1434(.a(gate121inter4), .b(gate121inter3), .O(gate121inter5));
  nor2  gate1435(.a(gate121inter5), .b(gate121inter2), .O(gate121inter6));
  inv1  gate1436(.a(G394), .O(gate121inter7));
  inv1  gate1437(.a(G395), .O(gate121inter8));
  nand2 gate1438(.a(gate121inter8), .b(gate121inter7), .O(gate121inter9));
  nand2 gate1439(.a(s_127), .b(gate121inter3), .O(gate121inter10));
  nor2  gate1440(.a(gate121inter10), .b(gate121inter9), .O(gate121inter11));
  nor2  gate1441(.a(gate121inter11), .b(gate121inter6), .O(gate121inter12));
  nand2 gate1442(.a(gate121inter12), .b(gate121inter1), .O(G474));
nand2 gate122( .a(G396), .b(G397), .O(G477) );
nand2 gate123( .a(G398), .b(G399), .O(G480) );

  xor2  gate1513(.a(G401), .b(G400), .O(gate124inter0));
  nand2 gate1514(.a(gate124inter0), .b(s_138), .O(gate124inter1));
  and2  gate1515(.a(G401), .b(G400), .O(gate124inter2));
  inv1  gate1516(.a(s_138), .O(gate124inter3));
  inv1  gate1517(.a(s_139), .O(gate124inter4));
  nand2 gate1518(.a(gate124inter4), .b(gate124inter3), .O(gate124inter5));
  nor2  gate1519(.a(gate124inter5), .b(gate124inter2), .O(gate124inter6));
  inv1  gate1520(.a(G400), .O(gate124inter7));
  inv1  gate1521(.a(G401), .O(gate124inter8));
  nand2 gate1522(.a(gate124inter8), .b(gate124inter7), .O(gate124inter9));
  nand2 gate1523(.a(s_139), .b(gate124inter3), .O(gate124inter10));
  nor2  gate1524(.a(gate124inter10), .b(gate124inter9), .O(gate124inter11));
  nor2  gate1525(.a(gate124inter11), .b(gate124inter6), .O(gate124inter12));
  nand2 gate1526(.a(gate124inter12), .b(gate124inter1), .O(G483));
nand2 gate125( .a(G402), .b(G403), .O(G486) );
nand2 gate126( .a(G404), .b(G405), .O(G489) );
nand2 gate127( .a(G406), .b(G407), .O(G492) );

  xor2  gate1947(.a(G409), .b(G408), .O(gate128inter0));
  nand2 gate1948(.a(gate128inter0), .b(s_200), .O(gate128inter1));
  and2  gate1949(.a(G409), .b(G408), .O(gate128inter2));
  inv1  gate1950(.a(s_200), .O(gate128inter3));
  inv1  gate1951(.a(s_201), .O(gate128inter4));
  nand2 gate1952(.a(gate128inter4), .b(gate128inter3), .O(gate128inter5));
  nor2  gate1953(.a(gate128inter5), .b(gate128inter2), .O(gate128inter6));
  inv1  gate1954(.a(G408), .O(gate128inter7));
  inv1  gate1955(.a(G409), .O(gate128inter8));
  nand2 gate1956(.a(gate128inter8), .b(gate128inter7), .O(gate128inter9));
  nand2 gate1957(.a(s_201), .b(gate128inter3), .O(gate128inter10));
  nor2  gate1958(.a(gate128inter10), .b(gate128inter9), .O(gate128inter11));
  nor2  gate1959(.a(gate128inter11), .b(gate128inter6), .O(gate128inter12));
  nand2 gate1960(.a(gate128inter12), .b(gate128inter1), .O(G495));

  xor2  gate1905(.a(G411), .b(G410), .O(gate129inter0));
  nand2 gate1906(.a(gate129inter0), .b(s_194), .O(gate129inter1));
  and2  gate1907(.a(G411), .b(G410), .O(gate129inter2));
  inv1  gate1908(.a(s_194), .O(gate129inter3));
  inv1  gate1909(.a(s_195), .O(gate129inter4));
  nand2 gate1910(.a(gate129inter4), .b(gate129inter3), .O(gate129inter5));
  nor2  gate1911(.a(gate129inter5), .b(gate129inter2), .O(gate129inter6));
  inv1  gate1912(.a(G410), .O(gate129inter7));
  inv1  gate1913(.a(G411), .O(gate129inter8));
  nand2 gate1914(.a(gate129inter8), .b(gate129inter7), .O(gate129inter9));
  nand2 gate1915(.a(s_195), .b(gate129inter3), .O(gate129inter10));
  nor2  gate1916(.a(gate129inter10), .b(gate129inter9), .O(gate129inter11));
  nor2  gate1917(.a(gate129inter11), .b(gate129inter6), .O(gate129inter12));
  nand2 gate1918(.a(gate129inter12), .b(gate129inter1), .O(G498));
nand2 gate130( .a(G412), .b(G413), .O(G501) );

  xor2  gate2199(.a(G415), .b(G414), .O(gate131inter0));
  nand2 gate2200(.a(gate131inter0), .b(s_236), .O(gate131inter1));
  and2  gate2201(.a(G415), .b(G414), .O(gate131inter2));
  inv1  gate2202(.a(s_236), .O(gate131inter3));
  inv1  gate2203(.a(s_237), .O(gate131inter4));
  nand2 gate2204(.a(gate131inter4), .b(gate131inter3), .O(gate131inter5));
  nor2  gate2205(.a(gate131inter5), .b(gate131inter2), .O(gate131inter6));
  inv1  gate2206(.a(G414), .O(gate131inter7));
  inv1  gate2207(.a(G415), .O(gate131inter8));
  nand2 gate2208(.a(gate131inter8), .b(gate131inter7), .O(gate131inter9));
  nand2 gate2209(.a(s_237), .b(gate131inter3), .O(gate131inter10));
  nor2  gate2210(.a(gate131inter10), .b(gate131inter9), .O(gate131inter11));
  nor2  gate2211(.a(gate131inter11), .b(gate131inter6), .O(gate131inter12));
  nand2 gate2212(.a(gate131inter12), .b(gate131inter1), .O(G504));

  xor2  gate1345(.a(G417), .b(G416), .O(gate132inter0));
  nand2 gate1346(.a(gate132inter0), .b(s_114), .O(gate132inter1));
  and2  gate1347(.a(G417), .b(G416), .O(gate132inter2));
  inv1  gate1348(.a(s_114), .O(gate132inter3));
  inv1  gate1349(.a(s_115), .O(gate132inter4));
  nand2 gate1350(.a(gate132inter4), .b(gate132inter3), .O(gate132inter5));
  nor2  gate1351(.a(gate132inter5), .b(gate132inter2), .O(gate132inter6));
  inv1  gate1352(.a(G416), .O(gate132inter7));
  inv1  gate1353(.a(G417), .O(gate132inter8));
  nand2 gate1354(.a(gate132inter8), .b(gate132inter7), .O(gate132inter9));
  nand2 gate1355(.a(s_115), .b(gate132inter3), .O(gate132inter10));
  nor2  gate1356(.a(gate132inter10), .b(gate132inter9), .O(gate132inter11));
  nor2  gate1357(.a(gate132inter11), .b(gate132inter6), .O(gate132inter12));
  nand2 gate1358(.a(gate132inter12), .b(gate132inter1), .O(G507));

  xor2  gate589(.a(G419), .b(G418), .O(gate133inter0));
  nand2 gate590(.a(gate133inter0), .b(s_6), .O(gate133inter1));
  and2  gate591(.a(G419), .b(G418), .O(gate133inter2));
  inv1  gate592(.a(s_6), .O(gate133inter3));
  inv1  gate593(.a(s_7), .O(gate133inter4));
  nand2 gate594(.a(gate133inter4), .b(gate133inter3), .O(gate133inter5));
  nor2  gate595(.a(gate133inter5), .b(gate133inter2), .O(gate133inter6));
  inv1  gate596(.a(G418), .O(gate133inter7));
  inv1  gate597(.a(G419), .O(gate133inter8));
  nand2 gate598(.a(gate133inter8), .b(gate133inter7), .O(gate133inter9));
  nand2 gate599(.a(s_7), .b(gate133inter3), .O(gate133inter10));
  nor2  gate600(.a(gate133inter10), .b(gate133inter9), .O(gate133inter11));
  nor2  gate601(.a(gate133inter11), .b(gate133inter6), .O(gate133inter12));
  nand2 gate602(.a(gate133inter12), .b(gate133inter1), .O(G510));

  xor2  gate1331(.a(G421), .b(G420), .O(gate134inter0));
  nand2 gate1332(.a(gate134inter0), .b(s_112), .O(gate134inter1));
  and2  gate1333(.a(G421), .b(G420), .O(gate134inter2));
  inv1  gate1334(.a(s_112), .O(gate134inter3));
  inv1  gate1335(.a(s_113), .O(gate134inter4));
  nand2 gate1336(.a(gate134inter4), .b(gate134inter3), .O(gate134inter5));
  nor2  gate1337(.a(gate134inter5), .b(gate134inter2), .O(gate134inter6));
  inv1  gate1338(.a(G420), .O(gate134inter7));
  inv1  gate1339(.a(G421), .O(gate134inter8));
  nand2 gate1340(.a(gate134inter8), .b(gate134inter7), .O(gate134inter9));
  nand2 gate1341(.a(s_113), .b(gate134inter3), .O(gate134inter10));
  nor2  gate1342(.a(gate134inter10), .b(gate134inter9), .O(gate134inter11));
  nor2  gate1343(.a(gate134inter11), .b(gate134inter6), .O(gate134inter12));
  nand2 gate1344(.a(gate134inter12), .b(gate134inter1), .O(G513));

  xor2  gate1065(.a(G423), .b(G422), .O(gate135inter0));
  nand2 gate1066(.a(gate135inter0), .b(s_74), .O(gate135inter1));
  and2  gate1067(.a(G423), .b(G422), .O(gate135inter2));
  inv1  gate1068(.a(s_74), .O(gate135inter3));
  inv1  gate1069(.a(s_75), .O(gate135inter4));
  nand2 gate1070(.a(gate135inter4), .b(gate135inter3), .O(gate135inter5));
  nor2  gate1071(.a(gate135inter5), .b(gate135inter2), .O(gate135inter6));
  inv1  gate1072(.a(G422), .O(gate135inter7));
  inv1  gate1073(.a(G423), .O(gate135inter8));
  nand2 gate1074(.a(gate135inter8), .b(gate135inter7), .O(gate135inter9));
  nand2 gate1075(.a(s_75), .b(gate135inter3), .O(gate135inter10));
  nor2  gate1076(.a(gate135inter10), .b(gate135inter9), .O(gate135inter11));
  nor2  gate1077(.a(gate135inter11), .b(gate135inter6), .O(gate135inter12));
  nand2 gate1078(.a(gate135inter12), .b(gate135inter1), .O(G516));
nand2 gate136( .a(G424), .b(G425), .O(G519) );

  xor2  gate1933(.a(G429), .b(G426), .O(gate137inter0));
  nand2 gate1934(.a(gate137inter0), .b(s_198), .O(gate137inter1));
  and2  gate1935(.a(G429), .b(G426), .O(gate137inter2));
  inv1  gate1936(.a(s_198), .O(gate137inter3));
  inv1  gate1937(.a(s_199), .O(gate137inter4));
  nand2 gate1938(.a(gate137inter4), .b(gate137inter3), .O(gate137inter5));
  nor2  gate1939(.a(gate137inter5), .b(gate137inter2), .O(gate137inter6));
  inv1  gate1940(.a(G426), .O(gate137inter7));
  inv1  gate1941(.a(G429), .O(gate137inter8));
  nand2 gate1942(.a(gate137inter8), .b(gate137inter7), .O(gate137inter9));
  nand2 gate1943(.a(s_199), .b(gate137inter3), .O(gate137inter10));
  nor2  gate1944(.a(gate137inter10), .b(gate137inter9), .O(gate137inter11));
  nor2  gate1945(.a(gate137inter11), .b(gate137inter6), .O(gate137inter12));
  nand2 gate1946(.a(gate137inter12), .b(gate137inter1), .O(G522));

  xor2  gate743(.a(G435), .b(G432), .O(gate138inter0));
  nand2 gate744(.a(gate138inter0), .b(s_28), .O(gate138inter1));
  and2  gate745(.a(G435), .b(G432), .O(gate138inter2));
  inv1  gate746(.a(s_28), .O(gate138inter3));
  inv1  gate747(.a(s_29), .O(gate138inter4));
  nand2 gate748(.a(gate138inter4), .b(gate138inter3), .O(gate138inter5));
  nor2  gate749(.a(gate138inter5), .b(gate138inter2), .O(gate138inter6));
  inv1  gate750(.a(G432), .O(gate138inter7));
  inv1  gate751(.a(G435), .O(gate138inter8));
  nand2 gate752(.a(gate138inter8), .b(gate138inter7), .O(gate138inter9));
  nand2 gate753(.a(s_29), .b(gate138inter3), .O(gate138inter10));
  nor2  gate754(.a(gate138inter10), .b(gate138inter9), .O(gate138inter11));
  nor2  gate755(.a(gate138inter11), .b(gate138inter6), .O(gate138inter12));
  nand2 gate756(.a(gate138inter12), .b(gate138inter1), .O(G525));
nand2 gate139( .a(G438), .b(G441), .O(G528) );
nand2 gate140( .a(G444), .b(G447), .O(G531) );
nand2 gate141( .a(G450), .b(G453), .O(G534) );
nand2 gate142( .a(G456), .b(G459), .O(G537) );
nand2 gate143( .a(G462), .b(G465), .O(G540) );

  xor2  gate1247(.a(G471), .b(G468), .O(gate144inter0));
  nand2 gate1248(.a(gate144inter0), .b(s_100), .O(gate144inter1));
  and2  gate1249(.a(G471), .b(G468), .O(gate144inter2));
  inv1  gate1250(.a(s_100), .O(gate144inter3));
  inv1  gate1251(.a(s_101), .O(gate144inter4));
  nand2 gate1252(.a(gate144inter4), .b(gate144inter3), .O(gate144inter5));
  nor2  gate1253(.a(gate144inter5), .b(gate144inter2), .O(gate144inter6));
  inv1  gate1254(.a(G468), .O(gate144inter7));
  inv1  gate1255(.a(G471), .O(gate144inter8));
  nand2 gate1256(.a(gate144inter8), .b(gate144inter7), .O(gate144inter9));
  nand2 gate1257(.a(s_101), .b(gate144inter3), .O(gate144inter10));
  nor2  gate1258(.a(gate144inter10), .b(gate144inter9), .O(gate144inter11));
  nor2  gate1259(.a(gate144inter11), .b(gate144inter6), .O(gate144inter12));
  nand2 gate1260(.a(gate144inter12), .b(gate144inter1), .O(G543));

  xor2  gate2647(.a(G477), .b(G474), .O(gate145inter0));
  nand2 gate2648(.a(gate145inter0), .b(s_300), .O(gate145inter1));
  and2  gate2649(.a(G477), .b(G474), .O(gate145inter2));
  inv1  gate2650(.a(s_300), .O(gate145inter3));
  inv1  gate2651(.a(s_301), .O(gate145inter4));
  nand2 gate2652(.a(gate145inter4), .b(gate145inter3), .O(gate145inter5));
  nor2  gate2653(.a(gate145inter5), .b(gate145inter2), .O(gate145inter6));
  inv1  gate2654(.a(G474), .O(gate145inter7));
  inv1  gate2655(.a(G477), .O(gate145inter8));
  nand2 gate2656(.a(gate145inter8), .b(gate145inter7), .O(gate145inter9));
  nand2 gate2657(.a(s_301), .b(gate145inter3), .O(gate145inter10));
  nor2  gate2658(.a(gate145inter10), .b(gate145inter9), .O(gate145inter11));
  nor2  gate2659(.a(gate145inter11), .b(gate145inter6), .O(gate145inter12));
  nand2 gate2660(.a(gate145inter12), .b(gate145inter1), .O(G546));
nand2 gate146( .a(G480), .b(G483), .O(G549) );

  xor2  gate1443(.a(G489), .b(G486), .O(gate147inter0));
  nand2 gate1444(.a(gate147inter0), .b(s_128), .O(gate147inter1));
  and2  gate1445(.a(G489), .b(G486), .O(gate147inter2));
  inv1  gate1446(.a(s_128), .O(gate147inter3));
  inv1  gate1447(.a(s_129), .O(gate147inter4));
  nand2 gate1448(.a(gate147inter4), .b(gate147inter3), .O(gate147inter5));
  nor2  gate1449(.a(gate147inter5), .b(gate147inter2), .O(gate147inter6));
  inv1  gate1450(.a(G486), .O(gate147inter7));
  inv1  gate1451(.a(G489), .O(gate147inter8));
  nand2 gate1452(.a(gate147inter8), .b(gate147inter7), .O(gate147inter9));
  nand2 gate1453(.a(s_129), .b(gate147inter3), .O(gate147inter10));
  nor2  gate1454(.a(gate147inter10), .b(gate147inter9), .O(gate147inter11));
  nor2  gate1455(.a(gate147inter11), .b(gate147inter6), .O(gate147inter12));
  nand2 gate1456(.a(gate147inter12), .b(gate147inter1), .O(G552));

  xor2  gate2311(.a(G495), .b(G492), .O(gate148inter0));
  nand2 gate2312(.a(gate148inter0), .b(s_252), .O(gate148inter1));
  and2  gate2313(.a(G495), .b(G492), .O(gate148inter2));
  inv1  gate2314(.a(s_252), .O(gate148inter3));
  inv1  gate2315(.a(s_253), .O(gate148inter4));
  nand2 gate2316(.a(gate148inter4), .b(gate148inter3), .O(gate148inter5));
  nor2  gate2317(.a(gate148inter5), .b(gate148inter2), .O(gate148inter6));
  inv1  gate2318(.a(G492), .O(gate148inter7));
  inv1  gate2319(.a(G495), .O(gate148inter8));
  nand2 gate2320(.a(gate148inter8), .b(gate148inter7), .O(gate148inter9));
  nand2 gate2321(.a(s_253), .b(gate148inter3), .O(gate148inter10));
  nor2  gate2322(.a(gate148inter10), .b(gate148inter9), .O(gate148inter11));
  nor2  gate2323(.a(gate148inter11), .b(gate148inter6), .O(gate148inter12));
  nand2 gate2324(.a(gate148inter12), .b(gate148inter1), .O(G555));
nand2 gate149( .a(G498), .b(G501), .O(G558) );
nand2 gate150( .a(G504), .b(G507), .O(G561) );
nand2 gate151( .a(G510), .b(G513), .O(G564) );

  xor2  gate1611(.a(G519), .b(G516), .O(gate152inter0));
  nand2 gate1612(.a(gate152inter0), .b(s_152), .O(gate152inter1));
  and2  gate1613(.a(G519), .b(G516), .O(gate152inter2));
  inv1  gate1614(.a(s_152), .O(gate152inter3));
  inv1  gate1615(.a(s_153), .O(gate152inter4));
  nand2 gate1616(.a(gate152inter4), .b(gate152inter3), .O(gate152inter5));
  nor2  gate1617(.a(gate152inter5), .b(gate152inter2), .O(gate152inter6));
  inv1  gate1618(.a(G516), .O(gate152inter7));
  inv1  gate1619(.a(G519), .O(gate152inter8));
  nand2 gate1620(.a(gate152inter8), .b(gate152inter7), .O(gate152inter9));
  nand2 gate1621(.a(s_153), .b(gate152inter3), .O(gate152inter10));
  nor2  gate1622(.a(gate152inter10), .b(gate152inter9), .O(gate152inter11));
  nor2  gate1623(.a(gate152inter11), .b(gate152inter6), .O(gate152inter12));
  nand2 gate1624(.a(gate152inter12), .b(gate152inter1), .O(G567));
nand2 gate153( .a(G426), .b(G522), .O(G570) );
nand2 gate154( .a(G429), .b(G522), .O(G571) );

  xor2  gate1107(.a(G525), .b(G432), .O(gate155inter0));
  nand2 gate1108(.a(gate155inter0), .b(s_80), .O(gate155inter1));
  and2  gate1109(.a(G525), .b(G432), .O(gate155inter2));
  inv1  gate1110(.a(s_80), .O(gate155inter3));
  inv1  gate1111(.a(s_81), .O(gate155inter4));
  nand2 gate1112(.a(gate155inter4), .b(gate155inter3), .O(gate155inter5));
  nor2  gate1113(.a(gate155inter5), .b(gate155inter2), .O(gate155inter6));
  inv1  gate1114(.a(G432), .O(gate155inter7));
  inv1  gate1115(.a(G525), .O(gate155inter8));
  nand2 gate1116(.a(gate155inter8), .b(gate155inter7), .O(gate155inter9));
  nand2 gate1117(.a(s_81), .b(gate155inter3), .O(gate155inter10));
  nor2  gate1118(.a(gate155inter10), .b(gate155inter9), .O(gate155inter11));
  nor2  gate1119(.a(gate155inter11), .b(gate155inter6), .O(gate155inter12));
  nand2 gate1120(.a(gate155inter12), .b(gate155inter1), .O(G572));
nand2 gate156( .a(G435), .b(G525), .O(G573) );

  xor2  gate1121(.a(G528), .b(G438), .O(gate157inter0));
  nand2 gate1122(.a(gate157inter0), .b(s_82), .O(gate157inter1));
  and2  gate1123(.a(G528), .b(G438), .O(gate157inter2));
  inv1  gate1124(.a(s_82), .O(gate157inter3));
  inv1  gate1125(.a(s_83), .O(gate157inter4));
  nand2 gate1126(.a(gate157inter4), .b(gate157inter3), .O(gate157inter5));
  nor2  gate1127(.a(gate157inter5), .b(gate157inter2), .O(gate157inter6));
  inv1  gate1128(.a(G438), .O(gate157inter7));
  inv1  gate1129(.a(G528), .O(gate157inter8));
  nand2 gate1130(.a(gate157inter8), .b(gate157inter7), .O(gate157inter9));
  nand2 gate1131(.a(s_83), .b(gate157inter3), .O(gate157inter10));
  nor2  gate1132(.a(gate157inter10), .b(gate157inter9), .O(gate157inter11));
  nor2  gate1133(.a(gate157inter11), .b(gate157inter6), .O(gate157inter12));
  nand2 gate1134(.a(gate157inter12), .b(gate157inter1), .O(G574));

  xor2  gate911(.a(G528), .b(G441), .O(gate158inter0));
  nand2 gate912(.a(gate158inter0), .b(s_52), .O(gate158inter1));
  and2  gate913(.a(G528), .b(G441), .O(gate158inter2));
  inv1  gate914(.a(s_52), .O(gate158inter3));
  inv1  gate915(.a(s_53), .O(gate158inter4));
  nand2 gate916(.a(gate158inter4), .b(gate158inter3), .O(gate158inter5));
  nor2  gate917(.a(gate158inter5), .b(gate158inter2), .O(gate158inter6));
  inv1  gate918(.a(G441), .O(gate158inter7));
  inv1  gate919(.a(G528), .O(gate158inter8));
  nand2 gate920(.a(gate158inter8), .b(gate158inter7), .O(gate158inter9));
  nand2 gate921(.a(s_53), .b(gate158inter3), .O(gate158inter10));
  nor2  gate922(.a(gate158inter10), .b(gate158inter9), .O(gate158inter11));
  nor2  gate923(.a(gate158inter11), .b(gate158inter6), .O(gate158inter12));
  nand2 gate924(.a(gate158inter12), .b(gate158inter1), .O(G575));

  xor2  gate2535(.a(G531), .b(G444), .O(gate159inter0));
  nand2 gate2536(.a(gate159inter0), .b(s_284), .O(gate159inter1));
  and2  gate2537(.a(G531), .b(G444), .O(gate159inter2));
  inv1  gate2538(.a(s_284), .O(gate159inter3));
  inv1  gate2539(.a(s_285), .O(gate159inter4));
  nand2 gate2540(.a(gate159inter4), .b(gate159inter3), .O(gate159inter5));
  nor2  gate2541(.a(gate159inter5), .b(gate159inter2), .O(gate159inter6));
  inv1  gate2542(.a(G444), .O(gate159inter7));
  inv1  gate2543(.a(G531), .O(gate159inter8));
  nand2 gate2544(.a(gate159inter8), .b(gate159inter7), .O(gate159inter9));
  nand2 gate2545(.a(s_285), .b(gate159inter3), .O(gate159inter10));
  nor2  gate2546(.a(gate159inter10), .b(gate159inter9), .O(gate159inter11));
  nor2  gate2547(.a(gate159inter11), .b(gate159inter6), .O(gate159inter12));
  nand2 gate2548(.a(gate159inter12), .b(gate159inter1), .O(G576));
nand2 gate160( .a(G447), .b(G531), .O(G577) );

  xor2  gate2255(.a(G534), .b(G450), .O(gate161inter0));
  nand2 gate2256(.a(gate161inter0), .b(s_244), .O(gate161inter1));
  and2  gate2257(.a(G534), .b(G450), .O(gate161inter2));
  inv1  gate2258(.a(s_244), .O(gate161inter3));
  inv1  gate2259(.a(s_245), .O(gate161inter4));
  nand2 gate2260(.a(gate161inter4), .b(gate161inter3), .O(gate161inter5));
  nor2  gate2261(.a(gate161inter5), .b(gate161inter2), .O(gate161inter6));
  inv1  gate2262(.a(G450), .O(gate161inter7));
  inv1  gate2263(.a(G534), .O(gate161inter8));
  nand2 gate2264(.a(gate161inter8), .b(gate161inter7), .O(gate161inter9));
  nand2 gate2265(.a(s_245), .b(gate161inter3), .O(gate161inter10));
  nor2  gate2266(.a(gate161inter10), .b(gate161inter9), .O(gate161inter11));
  nor2  gate2267(.a(gate161inter11), .b(gate161inter6), .O(gate161inter12));
  nand2 gate2268(.a(gate161inter12), .b(gate161inter1), .O(G578));

  xor2  gate2577(.a(G534), .b(G453), .O(gate162inter0));
  nand2 gate2578(.a(gate162inter0), .b(s_290), .O(gate162inter1));
  and2  gate2579(.a(G534), .b(G453), .O(gate162inter2));
  inv1  gate2580(.a(s_290), .O(gate162inter3));
  inv1  gate2581(.a(s_291), .O(gate162inter4));
  nand2 gate2582(.a(gate162inter4), .b(gate162inter3), .O(gate162inter5));
  nor2  gate2583(.a(gate162inter5), .b(gate162inter2), .O(gate162inter6));
  inv1  gate2584(.a(G453), .O(gate162inter7));
  inv1  gate2585(.a(G534), .O(gate162inter8));
  nand2 gate2586(.a(gate162inter8), .b(gate162inter7), .O(gate162inter9));
  nand2 gate2587(.a(s_291), .b(gate162inter3), .O(gate162inter10));
  nor2  gate2588(.a(gate162inter10), .b(gate162inter9), .O(gate162inter11));
  nor2  gate2589(.a(gate162inter11), .b(gate162inter6), .O(gate162inter12));
  nand2 gate2590(.a(gate162inter12), .b(gate162inter1), .O(G579));
nand2 gate163( .a(G456), .b(G537), .O(G580) );

  xor2  gate897(.a(G537), .b(G459), .O(gate164inter0));
  nand2 gate898(.a(gate164inter0), .b(s_50), .O(gate164inter1));
  and2  gate899(.a(G537), .b(G459), .O(gate164inter2));
  inv1  gate900(.a(s_50), .O(gate164inter3));
  inv1  gate901(.a(s_51), .O(gate164inter4));
  nand2 gate902(.a(gate164inter4), .b(gate164inter3), .O(gate164inter5));
  nor2  gate903(.a(gate164inter5), .b(gate164inter2), .O(gate164inter6));
  inv1  gate904(.a(G459), .O(gate164inter7));
  inv1  gate905(.a(G537), .O(gate164inter8));
  nand2 gate906(.a(gate164inter8), .b(gate164inter7), .O(gate164inter9));
  nand2 gate907(.a(s_51), .b(gate164inter3), .O(gate164inter10));
  nor2  gate908(.a(gate164inter10), .b(gate164inter9), .O(gate164inter11));
  nor2  gate909(.a(gate164inter11), .b(gate164inter6), .O(gate164inter12));
  nand2 gate910(.a(gate164inter12), .b(gate164inter1), .O(G581));
nand2 gate165( .a(G462), .b(G540), .O(G582) );

  xor2  gate981(.a(G540), .b(G465), .O(gate166inter0));
  nand2 gate982(.a(gate166inter0), .b(s_62), .O(gate166inter1));
  and2  gate983(.a(G540), .b(G465), .O(gate166inter2));
  inv1  gate984(.a(s_62), .O(gate166inter3));
  inv1  gate985(.a(s_63), .O(gate166inter4));
  nand2 gate986(.a(gate166inter4), .b(gate166inter3), .O(gate166inter5));
  nor2  gate987(.a(gate166inter5), .b(gate166inter2), .O(gate166inter6));
  inv1  gate988(.a(G465), .O(gate166inter7));
  inv1  gate989(.a(G540), .O(gate166inter8));
  nand2 gate990(.a(gate166inter8), .b(gate166inter7), .O(gate166inter9));
  nand2 gate991(.a(s_63), .b(gate166inter3), .O(gate166inter10));
  nor2  gate992(.a(gate166inter10), .b(gate166inter9), .O(gate166inter11));
  nor2  gate993(.a(gate166inter11), .b(gate166inter6), .O(gate166inter12));
  nand2 gate994(.a(gate166inter12), .b(gate166inter1), .O(G583));

  xor2  gate1681(.a(G543), .b(G468), .O(gate167inter0));
  nand2 gate1682(.a(gate167inter0), .b(s_162), .O(gate167inter1));
  and2  gate1683(.a(G543), .b(G468), .O(gate167inter2));
  inv1  gate1684(.a(s_162), .O(gate167inter3));
  inv1  gate1685(.a(s_163), .O(gate167inter4));
  nand2 gate1686(.a(gate167inter4), .b(gate167inter3), .O(gate167inter5));
  nor2  gate1687(.a(gate167inter5), .b(gate167inter2), .O(gate167inter6));
  inv1  gate1688(.a(G468), .O(gate167inter7));
  inv1  gate1689(.a(G543), .O(gate167inter8));
  nand2 gate1690(.a(gate167inter8), .b(gate167inter7), .O(gate167inter9));
  nand2 gate1691(.a(s_163), .b(gate167inter3), .O(gate167inter10));
  nor2  gate1692(.a(gate167inter10), .b(gate167inter9), .O(gate167inter11));
  nor2  gate1693(.a(gate167inter11), .b(gate167inter6), .O(gate167inter12));
  nand2 gate1694(.a(gate167inter12), .b(gate167inter1), .O(G584));
nand2 gate168( .a(G471), .b(G543), .O(G585) );
nand2 gate169( .a(G474), .b(G546), .O(G586) );
nand2 gate170( .a(G477), .b(G546), .O(G587) );
nand2 gate171( .a(G480), .b(G549), .O(G588) );

  xor2  gate1037(.a(G549), .b(G483), .O(gate172inter0));
  nand2 gate1038(.a(gate172inter0), .b(s_70), .O(gate172inter1));
  and2  gate1039(.a(G549), .b(G483), .O(gate172inter2));
  inv1  gate1040(.a(s_70), .O(gate172inter3));
  inv1  gate1041(.a(s_71), .O(gate172inter4));
  nand2 gate1042(.a(gate172inter4), .b(gate172inter3), .O(gate172inter5));
  nor2  gate1043(.a(gate172inter5), .b(gate172inter2), .O(gate172inter6));
  inv1  gate1044(.a(G483), .O(gate172inter7));
  inv1  gate1045(.a(G549), .O(gate172inter8));
  nand2 gate1046(.a(gate172inter8), .b(gate172inter7), .O(gate172inter9));
  nand2 gate1047(.a(s_71), .b(gate172inter3), .O(gate172inter10));
  nor2  gate1048(.a(gate172inter10), .b(gate172inter9), .O(gate172inter11));
  nor2  gate1049(.a(gate172inter11), .b(gate172inter6), .O(gate172inter12));
  nand2 gate1050(.a(gate172inter12), .b(gate172inter1), .O(G589));
nand2 gate173( .a(G486), .b(G552), .O(G590) );

  xor2  gate561(.a(G552), .b(G489), .O(gate174inter0));
  nand2 gate562(.a(gate174inter0), .b(s_2), .O(gate174inter1));
  and2  gate563(.a(G552), .b(G489), .O(gate174inter2));
  inv1  gate564(.a(s_2), .O(gate174inter3));
  inv1  gate565(.a(s_3), .O(gate174inter4));
  nand2 gate566(.a(gate174inter4), .b(gate174inter3), .O(gate174inter5));
  nor2  gate567(.a(gate174inter5), .b(gate174inter2), .O(gate174inter6));
  inv1  gate568(.a(G489), .O(gate174inter7));
  inv1  gate569(.a(G552), .O(gate174inter8));
  nand2 gate570(.a(gate174inter8), .b(gate174inter7), .O(gate174inter9));
  nand2 gate571(.a(s_3), .b(gate174inter3), .O(gate174inter10));
  nor2  gate572(.a(gate174inter10), .b(gate174inter9), .O(gate174inter11));
  nor2  gate573(.a(gate174inter11), .b(gate174inter6), .O(gate174inter12));
  nand2 gate574(.a(gate174inter12), .b(gate174inter1), .O(G591));
nand2 gate175( .a(G492), .b(G555), .O(G592) );
nand2 gate176( .a(G495), .b(G555), .O(G593) );
nand2 gate177( .a(G498), .b(G558), .O(G594) );
nand2 gate178( .a(G501), .b(G558), .O(G595) );

  xor2  gate1093(.a(G561), .b(G504), .O(gate179inter0));
  nand2 gate1094(.a(gate179inter0), .b(s_78), .O(gate179inter1));
  and2  gate1095(.a(G561), .b(G504), .O(gate179inter2));
  inv1  gate1096(.a(s_78), .O(gate179inter3));
  inv1  gate1097(.a(s_79), .O(gate179inter4));
  nand2 gate1098(.a(gate179inter4), .b(gate179inter3), .O(gate179inter5));
  nor2  gate1099(.a(gate179inter5), .b(gate179inter2), .O(gate179inter6));
  inv1  gate1100(.a(G504), .O(gate179inter7));
  inv1  gate1101(.a(G561), .O(gate179inter8));
  nand2 gate1102(.a(gate179inter8), .b(gate179inter7), .O(gate179inter9));
  nand2 gate1103(.a(s_79), .b(gate179inter3), .O(gate179inter10));
  nor2  gate1104(.a(gate179inter10), .b(gate179inter9), .O(gate179inter11));
  nor2  gate1105(.a(gate179inter11), .b(gate179inter6), .O(gate179inter12));
  nand2 gate1106(.a(gate179inter12), .b(gate179inter1), .O(G596));

  xor2  gate1877(.a(G561), .b(G507), .O(gate180inter0));
  nand2 gate1878(.a(gate180inter0), .b(s_190), .O(gate180inter1));
  and2  gate1879(.a(G561), .b(G507), .O(gate180inter2));
  inv1  gate1880(.a(s_190), .O(gate180inter3));
  inv1  gate1881(.a(s_191), .O(gate180inter4));
  nand2 gate1882(.a(gate180inter4), .b(gate180inter3), .O(gate180inter5));
  nor2  gate1883(.a(gate180inter5), .b(gate180inter2), .O(gate180inter6));
  inv1  gate1884(.a(G507), .O(gate180inter7));
  inv1  gate1885(.a(G561), .O(gate180inter8));
  nand2 gate1886(.a(gate180inter8), .b(gate180inter7), .O(gate180inter9));
  nand2 gate1887(.a(s_191), .b(gate180inter3), .O(gate180inter10));
  nor2  gate1888(.a(gate180inter10), .b(gate180inter9), .O(gate180inter11));
  nor2  gate1889(.a(gate180inter11), .b(gate180inter6), .O(gate180inter12));
  nand2 gate1890(.a(gate180inter12), .b(gate180inter1), .O(G597));
nand2 gate181( .a(G510), .b(G564), .O(G598) );
nand2 gate182( .a(G513), .b(G564), .O(G599) );
nand2 gate183( .a(G516), .b(G567), .O(G600) );
nand2 gate184( .a(G519), .b(G567), .O(G601) );

  xor2  gate1751(.a(G571), .b(G570), .O(gate185inter0));
  nand2 gate1752(.a(gate185inter0), .b(s_172), .O(gate185inter1));
  and2  gate1753(.a(G571), .b(G570), .O(gate185inter2));
  inv1  gate1754(.a(s_172), .O(gate185inter3));
  inv1  gate1755(.a(s_173), .O(gate185inter4));
  nand2 gate1756(.a(gate185inter4), .b(gate185inter3), .O(gate185inter5));
  nor2  gate1757(.a(gate185inter5), .b(gate185inter2), .O(gate185inter6));
  inv1  gate1758(.a(G570), .O(gate185inter7));
  inv1  gate1759(.a(G571), .O(gate185inter8));
  nand2 gate1760(.a(gate185inter8), .b(gate185inter7), .O(gate185inter9));
  nand2 gate1761(.a(s_173), .b(gate185inter3), .O(gate185inter10));
  nor2  gate1762(.a(gate185inter10), .b(gate185inter9), .O(gate185inter11));
  nor2  gate1763(.a(gate185inter11), .b(gate185inter6), .O(gate185inter12));
  nand2 gate1764(.a(gate185inter12), .b(gate185inter1), .O(G602));
nand2 gate186( .a(G572), .b(G573), .O(G607) );

  xor2  gate939(.a(G575), .b(G574), .O(gate187inter0));
  nand2 gate940(.a(gate187inter0), .b(s_56), .O(gate187inter1));
  and2  gate941(.a(G575), .b(G574), .O(gate187inter2));
  inv1  gate942(.a(s_56), .O(gate187inter3));
  inv1  gate943(.a(s_57), .O(gate187inter4));
  nand2 gate944(.a(gate187inter4), .b(gate187inter3), .O(gate187inter5));
  nor2  gate945(.a(gate187inter5), .b(gate187inter2), .O(gate187inter6));
  inv1  gate946(.a(G574), .O(gate187inter7));
  inv1  gate947(.a(G575), .O(gate187inter8));
  nand2 gate948(.a(gate187inter8), .b(gate187inter7), .O(gate187inter9));
  nand2 gate949(.a(s_57), .b(gate187inter3), .O(gate187inter10));
  nor2  gate950(.a(gate187inter10), .b(gate187inter9), .O(gate187inter11));
  nor2  gate951(.a(gate187inter11), .b(gate187inter6), .O(gate187inter12));
  nand2 gate952(.a(gate187inter12), .b(gate187inter1), .O(G612));

  xor2  gate799(.a(G577), .b(G576), .O(gate188inter0));
  nand2 gate800(.a(gate188inter0), .b(s_36), .O(gate188inter1));
  and2  gate801(.a(G577), .b(G576), .O(gate188inter2));
  inv1  gate802(.a(s_36), .O(gate188inter3));
  inv1  gate803(.a(s_37), .O(gate188inter4));
  nand2 gate804(.a(gate188inter4), .b(gate188inter3), .O(gate188inter5));
  nor2  gate805(.a(gate188inter5), .b(gate188inter2), .O(gate188inter6));
  inv1  gate806(.a(G576), .O(gate188inter7));
  inv1  gate807(.a(G577), .O(gate188inter8));
  nand2 gate808(.a(gate188inter8), .b(gate188inter7), .O(gate188inter9));
  nand2 gate809(.a(s_37), .b(gate188inter3), .O(gate188inter10));
  nor2  gate810(.a(gate188inter10), .b(gate188inter9), .O(gate188inter11));
  nor2  gate811(.a(gate188inter11), .b(gate188inter6), .O(gate188inter12));
  nand2 gate812(.a(gate188inter12), .b(gate188inter1), .O(G617));
nand2 gate189( .a(G578), .b(G579), .O(G622) );

  xor2  gate1289(.a(G581), .b(G580), .O(gate190inter0));
  nand2 gate1290(.a(gate190inter0), .b(s_106), .O(gate190inter1));
  and2  gate1291(.a(G581), .b(G580), .O(gate190inter2));
  inv1  gate1292(.a(s_106), .O(gate190inter3));
  inv1  gate1293(.a(s_107), .O(gate190inter4));
  nand2 gate1294(.a(gate190inter4), .b(gate190inter3), .O(gate190inter5));
  nor2  gate1295(.a(gate190inter5), .b(gate190inter2), .O(gate190inter6));
  inv1  gate1296(.a(G580), .O(gate190inter7));
  inv1  gate1297(.a(G581), .O(gate190inter8));
  nand2 gate1298(.a(gate190inter8), .b(gate190inter7), .O(gate190inter9));
  nand2 gate1299(.a(s_107), .b(gate190inter3), .O(gate190inter10));
  nor2  gate1300(.a(gate190inter10), .b(gate190inter9), .O(gate190inter11));
  nor2  gate1301(.a(gate190inter11), .b(gate190inter6), .O(gate190inter12));
  nand2 gate1302(.a(gate190inter12), .b(gate190inter1), .O(G627));
nand2 gate191( .a(G582), .b(G583), .O(G632) );

  xor2  gate2507(.a(G585), .b(G584), .O(gate192inter0));
  nand2 gate2508(.a(gate192inter0), .b(s_280), .O(gate192inter1));
  and2  gate2509(.a(G585), .b(G584), .O(gate192inter2));
  inv1  gate2510(.a(s_280), .O(gate192inter3));
  inv1  gate2511(.a(s_281), .O(gate192inter4));
  nand2 gate2512(.a(gate192inter4), .b(gate192inter3), .O(gate192inter5));
  nor2  gate2513(.a(gate192inter5), .b(gate192inter2), .O(gate192inter6));
  inv1  gate2514(.a(G584), .O(gate192inter7));
  inv1  gate2515(.a(G585), .O(gate192inter8));
  nand2 gate2516(.a(gate192inter8), .b(gate192inter7), .O(gate192inter9));
  nand2 gate2517(.a(s_281), .b(gate192inter3), .O(gate192inter10));
  nor2  gate2518(.a(gate192inter10), .b(gate192inter9), .O(gate192inter11));
  nor2  gate2519(.a(gate192inter11), .b(gate192inter6), .O(gate192inter12));
  nand2 gate2520(.a(gate192inter12), .b(gate192inter1), .O(G637));

  xor2  gate2339(.a(G587), .b(G586), .O(gate193inter0));
  nand2 gate2340(.a(gate193inter0), .b(s_256), .O(gate193inter1));
  and2  gate2341(.a(G587), .b(G586), .O(gate193inter2));
  inv1  gate2342(.a(s_256), .O(gate193inter3));
  inv1  gate2343(.a(s_257), .O(gate193inter4));
  nand2 gate2344(.a(gate193inter4), .b(gate193inter3), .O(gate193inter5));
  nor2  gate2345(.a(gate193inter5), .b(gate193inter2), .O(gate193inter6));
  inv1  gate2346(.a(G586), .O(gate193inter7));
  inv1  gate2347(.a(G587), .O(gate193inter8));
  nand2 gate2348(.a(gate193inter8), .b(gate193inter7), .O(gate193inter9));
  nand2 gate2349(.a(s_257), .b(gate193inter3), .O(gate193inter10));
  nor2  gate2350(.a(gate193inter10), .b(gate193inter9), .O(gate193inter11));
  nor2  gate2351(.a(gate193inter11), .b(gate193inter6), .O(gate193inter12));
  nand2 gate2352(.a(gate193inter12), .b(gate193inter1), .O(G642));
nand2 gate194( .a(G588), .b(G589), .O(G645) );
nand2 gate195( .a(G590), .b(G591), .O(G648) );
nand2 gate196( .a(G592), .b(G593), .O(G651) );

  xor2  gate2157(.a(G595), .b(G594), .O(gate197inter0));
  nand2 gate2158(.a(gate197inter0), .b(s_230), .O(gate197inter1));
  and2  gate2159(.a(G595), .b(G594), .O(gate197inter2));
  inv1  gate2160(.a(s_230), .O(gate197inter3));
  inv1  gate2161(.a(s_231), .O(gate197inter4));
  nand2 gate2162(.a(gate197inter4), .b(gate197inter3), .O(gate197inter5));
  nor2  gate2163(.a(gate197inter5), .b(gate197inter2), .O(gate197inter6));
  inv1  gate2164(.a(G594), .O(gate197inter7));
  inv1  gate2165(.a(G595), .O(gate197inter8));
  nand2 gate2166(.a(gate197inter8), .b(gate197inter7), .O(gate197inter9));
  nand2 gate2167(.a(s_231), .b(gate197inter3), .O(gate197inter10));
  nor2  gate2168(.a(gate197inter10), .b(gate197inter9), .O(gate197inter11));
  nor2  gate2169(.a(gate197inter11), .b(gate197inter6), .O(gate197inter12));
  nand2 gate2170(.a(gate197inter12), .b(gate197inter1), .O(G654));
nand2 gate198( .a(G596), .b(G597), .O(G657) );
nand2 gate199( .a(G598), .b(G599), .O(G660) );
nand2 gate200( .a(G600), .b(G601), .O(G663) );

  xor2  gate2283(.a(G607), .b(G602), .O(gate201inter0));
  nand2 gate2284(.a(gate201inter0), .b(s_248), .O(gate201inter1));
  and2  gate2285(.a(G607), .b(G602), .O(gate201inter2));
  inv1  gate2286(.a(s_248), .O(gate201inter3));
  inv1  gate2287(.a(s_249), .O(gate201inter4));
  nand2 gate2288(.a(gate201inter4), .b(gate201inter3), .O(gate201inter5));
  nor2  gate2289(.a(gate201inter5), .b(gate201inter2), .O(gate201inter6));
  inv1  gate2290(.a(G602), .O(gate201inter7));
  inv1  gate2291(.a(G607), .O(gate201inter8));
  nand2 gate2292(.a(gate201inter8), .b(gate201inter7), .O(gate201inter9));
  nand2 gate2293(.a(s_249), .b(gate201inter3), .O(gate201inter10));
  nor2  gate2294(.a(gate201inter10), .b(gate201inter9), .O(gate201inter11));
  nor2  gate2295(.a(gate201inter11), .b(gate201inter6), .O(gate201inter12));
  nand2 gate2296(.a(gate201inter12), .b(gate201inter1), .O(G666));
nand2 gate202( .a(G612), .b(G617), .O(G669) );

  xor2  gate2717(.a(G612), .b(G602), .O(gate203inter0));
  nand2 gate2718(.a(gate203inter0), .b(s_310), .O(gate203inter1));
  and2  gate2719(.a(G612), .b(G602), .O(gate203inter2));
  inv1  gate2720(.a(s_310), .O(gate203inter3));
  inv1  gate2721(.a(s_311), .O(gate203inter4));
  nand2 gate2722(.a(gate203inter4), .b(gate203inter3), .O(gate203inter5));
  nor2  gate2723(.a(gate203inter5), .b(gate203inter2), .O(gate203inter6));
  inv1  gate2724(.a(G602), .O(gate203inter7));
  inv1  gate2725(.a(G612), .O(gate203inter8));
  nand2 gate2726(.a(gate203inter8), .b(gate203inter7), .O(gate203inter9));
  nand2 gate2727(.a(s_311), .b(gate203inter3), .O(gate203inter10));
  nor2  gate2728(.a(gate203inter10), .b(gate203inter9), .O(gate203inter11));
  nor2  gate2729(.a(gate203inter11), .b(gate203inter6), .O(gate203inter12));
  nand2 gate2730(.a(gate203inter12), .b(gate203inter1), .O(G672));
nand2 gate204( .a(G607), .b(G617), .O(G675) );
nand2 gate205( .a(G622), .b(G627), .O(G678) );
nand2 gate206( .a(G632), .b(G637), .O(G681) );
nand2 gate207( .a(G622), .b(G632), .O(G684) );
nand2 gate208( .a(G627), .b(G637), .O(G687) );

  xor2  gate547(.a(G666), .b(G602), .O(gate209inter0));
  nand2 gate548(.a(gate209inter0), .b(s_0), .O(gate209inter1));
  and2  gate549(.a(G666), .b(G602), .O(gate209inter2));
  inv1  gate550(.a(s_0), .O(gate209inter3));
  inv1  gate551(.a(s_1), .O(gate209inter4));
  nand2 gate552(.a(gate209inter4), .b(gate209inter3), .O(gate209inter5));
  nor2  gate553(.a(gate209inter5), .b(gate209inter2), .O(gate209inter6));
  inv1  gate554(.a(G602), .O(gate209inter7));
  inv1  gate555(.a(G666), .O(gate209inter8));
  nand2 gate556(.a(gate209inter8), .b(gate209inter7), .O(gate209inter9));
  nand2 gate557(.a(s_1), .b(gate209inter3), .O(gate209inter10));
  nor2  gate558(.a(gate209inter10), .b(gate209inter9), .O(gate209inter11));
  nor2  gate559(.a(gate209inter11), .b(gate209inter6), .O(gate209inter12));
  nand2 gate560(.a(gate209inter12), .b(gate209inter1), .O(G690));
nand2 gate210( .a(G607), .b(G666), .O(G691) );

  xor2  gate1765(.a(G669), .b(G612), .O(gate211inter0));
  nand2 gate1766(.a(gate211inter0), .b(s_174), .O(gate211inter1));
  and2  gate1767(.a(G669), .b(G612), .O(gate211inter2));
  inv1  gate1768(.a(s_174), .O(gate211inter3));
  inv1  gate1769(.a(s_175), .O(gate211inter4));
  nand2 gate1770(.a(gate211inter4), .b(gate211inter3), .O(gate211inter5));
  nor2  gate1771(.a(gate211inter5), .b(gate211inter2), .O(gate211inter6));
  inv1  gate1772(.a(G612), .O(gate211inter7));
  inv1  gate1773(.a(G669), .O(gate211inter8));
  nand2 gate1774(.a(gate211inter8), .b(gate211inter7), .O(gate211inter9));
  nand2 gate1775(.a(s_175), .b(gate211inter3), .O(gate211inter10));
  nor2  gate1776(.a(gate211inter10), .b(gate211inter9), .O(gate211inter11));
  nor2  gate1777(.a(gate211inter11), .b(gate211inter6), .O(gate211inter12));
  nand2 gate1778(.a(gate211inter12), .b(gate211inter1), .O(G692));
nand2 gate212( .a(G617), .b(G669), .O(G693) );
nand2 gate213( .a(G602), .b(G672), .O(G694) );
nand2 gate214( .a(G612), .b(G672), .O(G695) );

  xor2  gate2227(.a(G675), .b(G607), .O(gate215inter0));
  nand2 gate2228(.a(gate215inter0), .b(s_240), .O(gate215inter1));
  and2  gate2229(.a(G675), .b(G607), .O(gate215inter2));
  inv1  gate2230(.a(s_240), .O(gate215inter3));
  inv1  gate2231(.a(s_241), .O(gate215inter4));
  nand2 gate2232(.a(gate215inter4), .b(gate215inter3), .O(gate215inter5));
  nor2  gate2233(.a(gate215inter5), .b(gate215inter2), .O(gate215inter6));
  inv1  gate2234(.a(G607), .O(gate215inter7));
  inv1  gate2235(.a(G675), .O(gate215inter8));
  nand2 gate2236(.a(gate215inter8), .b(gate215inter7), .O(gate215inter9));
  nand2 gate2237(.a(s_241), .b(gate215inter3), .O(gate215inter10));
  nor2  gate2238(.a(gate215inter10), .b(gate215inter9), .O(gate215inter11));
  nor2  gate2239(.a(gate215inter11), .b(gate215inter6), .O(gate215inter12));
  nand2 gate2240(.a(gate215inter12), .b(gate215inter1), .O(G696));

  xor2  gate1023(.a(G675), .b(G617), .O(gate216inter0));
  nand2 gate1024(.a(gate216inter0), .b(s_68), .O(gate216inter1));
  and2  gate1025(.a(G675), .b(G617), .O(gate216inter2));
  inv1  gate1026(.a(s_68), .O(gate216inter3));
  inv1  gate1027(.a(s_69), .O(gate216inter4));
  nand2 gate1028(.a(gate216inter4), .b(gate216inter3), .O(gate216inter5));
  nor2  gate1029(.a(gate216inter5), .b(gate216inter2), .O(gate216inter6));
  inv1  gate1030(.a(G617), .O(gate216inter7));
  inv1  gate1031(.a(G675), .O(gate216inter8));
  nand2 gate1032(.a(gate216inter8), .b(gate216inter7), .O(gate216inter9));
  nand2 gate1033(.a(s_69), .b(gate216inter3), .O(gate216inter10));
  nor2  gate1034(.a(gate216inter10), .b(gate216inter9), .O(gate216inter11));
  nor2  gate1035(.a(gate216inter11), .b(gate216inter6), .O(gate216inter12));
  nand2 gate1036(.a(gate216inter12), .b(gate216inter1), .O(G697));
nand2 gate217( .a(G622), .b(G678), .O(G698) );
nand2 gate218( .a(G627), .b(G678), .O(G699) );
nand2 gate219( .a(G632), .b(G681), .O(G700) );

  xor2  gate2423(.a(G681), .b(G637), .O(gate220inter0));
  nand2 gate2424(.a(gate220inter0), .b(s_268), .O(gate220inter1));
  and2  gate2425(.a(G681), .b(G637), .O(gate220inter2));
  inv1  gate2426(.a(s_268), .O(gate220inter3));
  inv1  gate2427(.a(s_269), .O(gate220inter4));
  nand2 gate2428(.a(gate220inter4), .b(gate220inter3), .O(gate220inter5));
  nor2  gate2429(.a(gate220inter5), .b(gate220inter2), .O(gate220inter6));
  inv1  gate2430(.a(G637), .O(gate220inter7));
  inv1  gate2431(.a(G681), .O(gate220inter8));
  nand2 gate2432(.a(gate220inter8), .b(gate220inter7), .O(gate220inter9));
  nand2 gate2433(.a(s_269), .b(gate220inter3), .O(gate220inter10));
  nor2  gate2434(.a(gate220inter10), .b(gate220inter9), .O(gate220inter11));
  nor2  gate2435(.a(gate220inter11), .b(gate220inter6), .O(gate220inter12));
  nand2 gate2436(.a(gate220inter12), .b(gate220inter1), .O(G701));

  xor2  gate2395(.a(G684), .b(G622), .O(gate221inter0));
  nand2 gate2396(.a(gate221inter0), .b(s_264), .O(gate221inter1));
  and2  gate2397(.a(G684), .b(G622), .O(gate221inter2));
  inv1  gate2398(.a(s_264), .O(gate221inter3));
  inv1  gate2399(.a(s_265), .O(gate221inter4));
  nand2 gate2400(.a(gate221inter4), .b(gate221inter3), .O(gate221inter5));
  nor2  gate2401(.a(gate221inter5), .b(gate221inter2), .O(gate221inter6));
  inv1  gate2402(.a(G622), .O(gate221inter7));
  inv1  gate2403(.a(G684), .O(gate221inter8));
  nand2 gate2404(.a(gate221inter8), .b(gate221inter7), .O(gate221inter9));
  nand2 gate2405(.a(s_265), .b(gate221inter3), .O(gate221inter10));
  nor2  gate2406(.a(gate221inter10), .b(gate221inter9), .O(gate221inter11));
  nor2  gate2407(.a(gate221inter11), .b(gate221inter6), .O(gate221inter12));
  nand2 gate2408(.a(gate221inter12), .b(gate221inter1), .O(G702));
nand2 gate222( .a(G632), .b(G684), .O(G703) );

  xor2  gate1835(.a(G687), .b(G627), .O(gate223inter0));
  nand2 gate1836(.a(gate223inter0), .b(s_184), .O(gate223inter1));
  and2  gate1837(.a(G687), .b(G627), .O(gate223inter2));
  inv1  gate1838(.a(s_184), .O(gate223inter3));
  inv1  gate1839(.a(s_185), .O(gate223inter4));
  nand2 gate1840(.a(gate223inter4), .b(gate223inter3), .O(gate223inter5));
  nor2  gate1841(.a(gate223inter5), .b(gate223inter2), .O(gate223inter6));
  inv1  gate1842(.a(G627), .O(gate223inter7));
  inv1  gate1843(.a(G687), .O(gate223inter8));
  nand2 gate1844(.a(gate223inter8), .b(gate223inter7), .O(gate223inter9));
  nand2 gate1845(.a(s_185), .b(gate223inter3), .O(gate223inter10));
  nor2  gate1846(.a(gate223inter10), .b(gate223inter9), .O(gate223inter11));
  nor2  gate1847(.a(gate223inter11), .b(gate223inter6), .O(gate223inter12));
  nand2 gate1848(.a(gate223inter12), .b(gate223inter1), .O(G704));
nand2 gate224( .a(G637), .b(G687), .O(G705) );

  xor2  gate883(.a(G691), .b(G690), .O(gate225inter0));
  nand2 gate884(.a(gate225inter0), .b(s_48), .O(gate225inter1));
  and2  gate885(.a(G691), .b(G690), .O(gate225inter2));
  inv1  gate886(.a(s_48), .O(gate225inter3));
  inv1  gate887(.a(s_49), .O(gate225inter4));
  nand2 gate888(.a(gate225inter4), .b(gate225inter3), .O(gate225inter5));
  nor2  gate889(.a(gate225inter5), .b(gate225inter2), .O(gate225inter6));
  inv1  gate890(.a(G690), .O(gate225inter7));
  inv1  gate891(.a(G691), .O(gate225inter8));
  nand2 gate892(.a(gate225inter8), .b(gate225inter7), .O(gate225inter9));
  nand2 gate893(.a(s_49), .b(gate225inter3), .O(gate225inter10));
  nor2  gate894(.a(gate225inter10), .b(gate225inter9), .O(gate225inter11));
  nor2  gate895(.a(gate225inter11), .b(gate225inter6), .O(gate225inter12));
  nand2 gate896(.a(gate225inter12), .b(gate225inter1), .O(G706));
nand2 gate226( .a(G692), .b(G693), .O(G709) );

  xor2  gate1527(.a(G695), .b(G694), .O(gate227inter0));
  nand2 gate1528(.a(gate227inter0), .b(s_140), .O(gate227inter1));
  and2  gate1529(.a(G695), .b(G694), .O(gate227inter2));
  inv1  gate1530(.a(s_140), .O(gate227inter3));
  inv1  gate1531(.a(s_141), .O(gate227inter4));
  nand2 gate1532(.a(gate227inter4), .b(gate227inter3), .O(gate227inter5));
  nor2  gate1533(.a(gate227inter5), .b(gate227inter2), .O(gate227inter6));
  inv1  gate1534(.a(G694), .O(gate227inter7));
  inv1  gate1535(.a(G695), .O(gate227inter8));
  nand2 gate1536(.a(gate227inter8), .b(gate227inter7), .O(gate227inter9));
  nand2 gate1537(.a(s_141), .b(gate227inter3), .O(gate227inter10));
  nor2  gate1538(.a(gate227inter10), .b(gate227inter9), .O(gate227inter11));
  nor2  gate1539(.a(gate227inter11), .b(gate227inter6), .O(gate227inter12));
  nand2 gate1540(.a(gate227inter12), .b(gate227inter1), .O(G712));

  xor2  gate2465(.a(G697), .b(G696), .O(gate228inter0));
  nand2 gate2466(.a(gate228inter0), .b(s_274), .O(gate228inter1));
  and2  gate2467(.a(G697), .b(G696), .O(gate228inter2));
  inv1  gate2468(.a(s_274), .O(gate228inter3));
  inv1  gate2469(.a(s_275), .O(gate228inter4));
  nand2 gate2470(.a(gate228inter4), .b(gate228inter3), .O(gate228inter5));
  nor2  gate2471(.a(gate228inter5), .b(gate228inter2), .O(gate228inter6));
  inv1  gate2472(.a(G696), .O(gate228inter7));
  inv1  gate2473(.a(G697), .O(gate228inter8));
  nand2 gate2474(.a(gate228inter8), .b(gate228inter7), .O(gate228inter9));
  nand2 gate2475(.a(s_275), .b(gate228inter3), .O(gate228inter10));
  nor2  gate2476(.a(gate228inter10), .b(gate228inter9), .O(gate228inter11));
  nor2  gate2477(.a(gate228inter11), .b(gate228inter6), .O(gate228inter12));
  nand2 gate2478(.a(gate228inter12), .b(gate228inter1), .O(G715));

  xor2  gate2675(.a(G699), .b(G698), .O(gate229inter0));
  nand2 gate2676(.a(gate229inter0), .b(s_304), .O(gate229inter1));
  and2  gate2677(.a(G699), .b(G698), .O(gate229inter2));
  inv1  gate2678(.a(s_304), .O(gate229inter3));
  inv1  gate2679(.a(s_305), .O(gate229inter4));
  nand2 gate2680(.a(gate229inter4), .b(gate229inter3), .O(gate229inter5));
  nor2  gate2681(.a(gate229inter5), .b(gate229inter2), .O(gate229inter6));
  inv1  gate2682(.a(G698), .O(gate229inter7));
  inv1  gate2683(.a(G699), .O(gate229inter8));
  nand2 gate2684(.a(gate229inter8), .b(gate229inter7), .O(gate229inter9));
  nand2 gate2685(.a(s_305), .b(gate229inter3), .O(gate229inter10));
  nor2  gate2686(.a(gate229inter10), .b(gate229inter9), .O(gate229inter11));
  nor2  gate2687(.a(gate229inter11), .b(gate229inter6), .O(gate229inter12));
  nand2 gate2688(.a(gate229inter12), .b(gate229inter1), .O(G718));

  xor2  gate1149(.a(G701), .b(G700), .O(gate230inter0));
  nand2 gate1150(.a(gate230inter0), .b(s_86), .O(gate230inter1));
  and2  gate1151(.a(G701), .b(G700), .O(gate230inter2));
  inv1  gate1152(.a(s_86), .O(gate230inter3));
  inv1  gate1153(.a(s_87), .O(gate230inter4));
  nand2 gate1154(.a(gate230inter4), .b(gate230inter3), .O(gate230inter5));
  nor2  gate1155(.a(gate230inter5), .b(gate230inter2), .O(gate230inter6));
  inv1  gate1156(.a(G700), .O(gate230inter7));
  inv1  gate1157(.a(G701), .O(gate230inter8));
  nand2 gate1158(.a(gate230inter8), .b(gate230inter7), .O(gate230inter9));
  nand2 gate1159(.a(s_87), .b(gate230inter3), .O(gate230inter10));
  nor2  gate1160(.a(gate230inter10), .b(gate230inter9), .O(gate230inter11));
  nor2  gate1161(.a(gate230inter11), .b(gate230inter6), .O(gate230inter12));
  nand2 gate1162(.a(gate230inter12), .b(gate230inter1), .O(G721));
nand2 gate231( .a(G702), .b(G703), .O(G724) );

  xor2  gate2213(.a(G705), .b(G704), .O(gate232inter0));
  nand2 gate2214(.a(gate232inter0), .b(s_238), .O(gate232inter1));
  and2  gate2215(.a(G705), .b(G704), .O(gate232inter2));
  inv1  gate2216(.a(s_238), .O(gate232inter3));
  inv1  gate2217(.a(s_239), .O(gate232inter4));
  nand2 gate2218(.a(gate232inter4), .b(gate232inter3), .O(gate232inter5));
  nor2  gate2219(.a(gate232inter5), .b(gate232inter2), .O(gate232inter6));
  inv1  gate2220(.a(G704), .O(gate232inter7));
  inv1  gate2221(.a(G705), .O(gate232inter8));
  nand2 gate2222(.a(gate232inter8), .b(gate232inter7), .O(gate232inter9));
  nand2 gate2223(.a(s_239), .b(gate232inter3), .O(gate232inter10));
  nor2  gate2224(.a(gate232inter10), .b(gate232inter9), .O(gate232inter11));
  nor2  gate2225(.a(gate232inter11), .b(gate232inter6), .O(gate232inter12));
  nand2 gate2226(.a(gate232inter12), .b(gate232inter1), .O(G727));

  xor2  gate2605(.a(G718), .b(G242), .O(gate233inter0));
  nand2 gate2606(.a(gate233inter0), .b(s_294), .O(gate233inter1));
  and2  gate2607(.a(G718), .b(G242), .O(gate233inter2));
  inv1  gate2608(.a(s_294), .O(gate233inter3));
  inv1  gate2609(.a(s_295), .O(gate233inter4));
  nand2 gate2610(.a(gate233inter4), .b(gate233inter3), .O(gate233inter5));
  nor2  gate2611(.a(gate233inter5), .b(gate233inter2), .O(gate233inter6));
  inv1  gate2612(.a(G242), .O(gate233inter7));
  inv1  gate2613(.a(G718), .O(gate233inter8));
  nand2 gate2614(.a(gate233inter8), .b(gate233inter7), .O(gate233inter9));
  nand2 gate2615(.a(s_295), .b(gate233inter3), .O(gate233inter10));
  nor2  gate2616(.a(gate233inter10), .b(gate233inter9), .O(gate233inter11));
  nor2  gate2617(.a(gate233inter11), .b(gate233inter6), .O(gate233inter12));
  nand2 gate2618(.a(gate233inter12), .b(gate233inter1), .O(G730));

  xor2  gate2479(.a(G721), .b(G245), .O(gate234inter0));
  nand2 gate2480(.a(gate234inter0), .b(s_276), .O(gate234inter1));
  and2  gate2481(.a(G721), .b(G245), .O(gate234inter2));
  inv1  gate2482(.a(s_276), .O(gate234inter3));
  inv1  gate2483(.a(s_277), .O(gate234inter4));
  nand2 gate2484(.a(gate234inter4), .b(gate234inter3), .O(gate234inter5));
  nor2  gate2485(.a(gate234inter5), .b(gate234inter2), .O(gate234inter6));
  inv1  gate2486(.a(G245), .O(gate234inter7));
  inv1  gate2487(.a(G721), .O(gate234inter8));
  nand2 gate2488(.a(gate234inter8), .b(gate234inter7), .O(gate234inter9));
  nand2 gate2489(.a(s_277), .b(gate234inter3), .O(gate234inter10));
  nor2  gate2490(.a(gate234inter10), .b(gate234inter9), .O(gate234inter11));
  nor2  gate2491(.a(gate234inter11), .b(gate234inter6), .O(gate234inter12));
  nand2 gate2492(.a(gate234inter12), .b(gate234inter1), .O(G733));

  xor2  gate2045(.a(G724), .b(G248), .O(gate235inter0));
  nand2 gate2046(.a(gate235inter0), .b(s_214), .O(gate235inter1));
  and2  gate2047(.a(G724), .b(G248), .O(gate235inter2));
  inv1  gate2048(.a(s_214), .O(gate235inter3));
  inv1  gate2049(.a(s_215), .O(gate235inter4));
  nand2 gate2050(.a(gate235inter4), .b(gate235inter3), .O(gate235inter5));
  nor2  gate2051(.a(gate235inter5), .b(gate235inter2), .O(gate235inter6));
  inv1  gate2052(.a(G248), .O(gate235inter7));
  inv1  gate2053(.a(G724), .O(gate235inter8));
  nand2 gate2054(.a(gate235inter8), .b(gate235inter7), .O(gate235inter9));
  nand2 gate2055(.a(s_215), .b(gate235inter3), .O(gate235inter10));
  nor2  gate2056(.a(gate235inter10), .b(gate235inter9), .O(gate235inter11));
  nor2  gate2057(.a(gate235inter11), .b(gate235inter6), .O(gate235inter12));
  nand2 gate2058(.a(gate235inter12), .b(gate235inter1), .O(G736));
nand2 gate236( .a(G251), .b(G727), .O(G739) );
nand2 gate237( .a(G254), .b(G706), .O(G742) );

  xor2  gate2703(.a(G709), .b(G257), .O(gate238inter0));
  nand2 gate2704(.a(gate238inter0), .b(s_308), .O(gate238inter1));
  and2  gate2705(.a(G709), .b(G257), .O(gate238inter2));
  inv1  gate2706(.a(s_308), .O(gate238inter3));
  inv1  gate2707(.a(s_309), .O(gate238inter4));
  nand2 gate2708(.a(gate238inter4), .b(gate238inter3), .O(gate238inter5));
  nor2  gate2709(.a(gate238inter5), .b(gate238inter2), .O(gate238inter6));
  inv1  gate2710(.a(G257), .O(gate238inter7));
  inv1  gate2711(.a(G709), .O(gate238inter8));
  nand2 gate2712(.a(gate238inter8), .b(gate238inter7), .O(gate238inter9));
  nand2 gate2713(.a(s_309), .b(gate238inter3), .O(gate238inter10));
  nor2  gate2714(.a(gate238inter10), .b(gate238inter9), .O(gate238inter11));
  nor2  gate2715(.a(gate238inter11), .b(gate238inter6), .O(gate238inter12));
  nand2 gate2716(.a(gate238inter12), .b(gate238inter1), .O(G745));

  xor2  gate2129(.a(G712), .b(G260), .O(gate239inter0));
  nand2 gate2130(.a(gate239inter0), .b(s_226), .O(gate239inter1));
  and2  gate2131(.a(G712), .b(G260), .O(gate239inter2));
  inv1  gate2132(.a(s_226), .O(gate239inter3));
  inv1  gate2133(.a(s_227), .O(gate239inter4));
  nand2 gate2134(.a(gate239inter4), .b(gate239inter3), .O(gate239inter5));
  nor2  gate2135(.a(gate239inter5), .b(gate239inter2), .O(gate239inter6));
  inv1  gate2136(.a(G260), .O(gate239inter7));
  inv1  gate2137(.a(G712), .O(gate239inter8));
  nand2 gate2138(.a(gate239inter8), .b(gate239inter7), .O(gate239inter9));
  nand2 gate2139(.a(s_227), .b(gate239inter3), .O(gate239inter10));
  nor2  gate2140(.a(gate239inter10), .b(gate239inter9), .O(gate239inter11));
  nor2  gate2141(.a(gate239inter11), .b(gate239inter6), .O(gate239inter12));
  nand2 gate2142(.a(gate239inter12), .b(gate239inter1), .O(G748));
nand2 gate240( .a(G263), .b(G715), .O(G751) );
nand2 gate241( .a(G242), .b(G730), .O(G754) );
nand2 gate242( .a(G718), .b(G730), .O(G755) );
nand2 gate243( .a(G245), .b(G733), .O(G756) );
nand2 gate244( .a(G721), .b(G733), .O(G757) );
nand2 gate245( .a(G248), .b(G736), .O(G758) );
nand2 gate246( .a(G724), .b(G736), .O(G759) );
nand2 gate247( .a(G251), .b(G739), .O(G760) );
nand2 gate248( .a(G727), .b(G739), .O(G761) );

  xor2  gate771(.a(G742), .b(G254), .O(gate249inter0));
  nand2 gate772(.a(gate249inter0), .b(s_32), .O(gate249inter1));
  and2  gate773(.a(G742), .b(G254), .O(gate249inter2));
  inv1  gate774(.a(s_32), .O(gate249inter3));
  inv1  gate775(.a(s_33), .O(gate249inter4));
  nand2 gate776(.a(gate249inter4), .b(gate249inter3), .O(gate249inter5));
  nor2  gate777(.a(gate249inter5), .b(gate249inter2), .O(gate249inter6));
  inv1  gate778(.a(G254), .O(gate249inter7));
  inv1  gate779(.a(G742), .O(gate249inter8));
  nand2 gate780(.a(gate249inter8), .b(gate249inter7), .O(gate249inter9));
  nand2 gate781(.a(s_33), .b(gate249inter3), .O(gate249inter10));
  nor2  gate782(.a(gate249inter10), .b(gate249inter9), .O(gate249inter11));
  nor2  gate783(.a(gate249inter11), .b(gate249inter6), .O(gate249inter12));
  nand2 gate784(.a(gate249inter12), .b(gate249inter1), .O(G762));
nand2 gate250( .a(G706), .b(G742), .O(G763) );
nand2 gate251( .a(G257), .b(G745), .O(G764) );
nand2 gate252( .a(G709), .b(G745), .O(G765) );

  xor2  gate2633(.a(G748), .b(G260), .O(gate253inter0));
  nand2 gate2634(.a(gate253inter0), .b(s_298), .O(gate253inter1));
  and2  gate2635(.a(G748), .b(G260), .O(gate253inter2));
  inv1  gate2636(.a(s_298), .O(gate253inter3));
  inv1  gate2637(.a(s_299), .O(gate253inter4));
  nand2 gate2638(.a(gate253inter4), .b(gate253inter3), .O(gate253inter5));
  nor2  gate2639(.a(gate253inter5), .b(gate253inter2), .O(gate253inter6));
  inv1  gate2640(.a(G260), .O(gate253inter7));
  inv1  gate2641(.a(G748), .O(gate253inter8));
  nand2 gate2642(.a(gate253inter8), .b(gate253inter7), .O(gate253inter9));
  nand2 gate2643(.a(s_299), .b(gate253inter3), .O(gate253inter10));
  nor2  gate2644(.a(gate253inter10), .b(gate253inter9), .O(gate253inter11));
  nor2  gate2645(.a(gate253inter11), .b(gate253inter6), .O(gate253inter12));
  nand2 gate2646(.a(gate253inter12), .b(gate253inter1), .O(G766));
nand2 gate254( .a(G712), .b(G748), .O(G767) );

  xor2  gate2241(.a(G751), .b(G263), .O(gate255inter0));
  nand2 gate2242(.a(gate255inter0), .b(s_242), .O(gate255inter1));
  and2  gate2243(.a(G751), .b(G263), .O(gate255inter2));
  inv1  gate2244(.a(s_242), .O(gate255inter3));
  inv1  gate2245(.a(s_243), .O(gate255inter4));
  nand2 gate2246(.a(gate255inter4), .b(gate255inter3), .O(gate255inter5));
  nor2  gate2247(.a(gate255inter5), .b(gate255inter2), .O(gate255inter6));
  inv1  gate2248(.a(G263), .O(gate255inter7));
  inv1  gate2249(.a(G751), .O(gate255inter8));
  nand2 gate2250(.a(gate255inter8), .b(gate255inter7), .O(gate255inter9));
  nand2 gate2251(.a(s_243), .b(gate255inter3), .O(gate255inter10));
  nor2  gate2252(.a(gate255inter10), .b(gate255inter9), .O(gate255inter11));
  nor2  gate2253(.a(gate255inter11), .b(gate255inter6), .O(gate255inter12));
  nand2 gate2254(.a(gate255inter12), .b(gate255inter1), .O(G768));
nand2 gate256( .a(G715), .b(G751), .O(G769) );

  xor2  gate2563(.a(G755), .b(G754), .O(gate257inter0));
  nand2 gate2564(.a(gate257inter0), .b(s_288), .O(gate257inter1));
  and2  gate2565(.a(G755), .b(G754), .O(gate257inter2));
  inv1  gate2566(.a(s_288), .O(gate257inter3));
  inv1  gate2567(.a(s_289), .O(gate257inter4));
  nand2 gate2568(.a(gate257inter4), .b(gate257inter3), .O(gate257inter5));
  nor2  gate2569(.a(gate257inter5), .b(gate257inter2), .O(gate257inter6));
  inv1  gate2570(.a(G754), .O(gate257inter7));
  inv1  gate2571(.a(G755), .O(gate257inter8));
  nand2 gate2572(.a(gate257inter8), .b(gate257inter7), .O(gate257inter9));
  nand2 gate2573(.a(s_289), .b(gate257inter3), .O(gate257inter10));
  nor2  gate2574(.a(gate257inter10), .b(gate257inter9), .O(gate257inter11));
  nor2  gate2575(.a(gate257inter11), .b(gate257inter6), .O(gate257inter12));
  nand2 gate2576(.a(gate257inter12), .b(gate257inter1), .O(G770));
nand2 gate258( .a(G756), .b(G757), .O(G773) );
nand2 gate259( .a(G758), .b(G759), .O(G776) );
nand2 gate260( .a(G760), .b(G761), .O(G779) );

  xor2  gate2115(.a(G763), .b(G762), .O(gate261inter0));
  nand2 gate2116(.a(gate261inter0), .b(s_224), .O(gate261inter1));
  and2  gate2117(.a(G763), .b(G762), .O(gate261inter2));
  inv1  gate2118(.a(s_224), .O(gate261inter3));
  inv1  gate2119(.a(s_225), .O(gate261inter4));
  nand2 gate2120(.a(gate261inter4), .b(gate261inter3), .O(gate261inter5));
  nor2  gate2121(.a(gate261inter5), .b(gate261inter2), .O(gate261inter6));
  inv1  gate2122(.a(G762), .O(gate261inter7));
  inv1  gate2123(.a(G763), .O(gate261inter8));
  nand2 gate2124(.a(gate261inter8), .b(gate261inter7), .O(gate261inter9));
  nand2 gate2125(.a(s_225), .b(gate261inter3), .O(gate261inter10));
  nor2  gate2126(.a(gate261inter10), .b(gate261inter9), .O(gate261inter11));
  nor2  gate2127(.a(gate261inter11), .b(gate261inter6), .O(gate261inter12));
  nand2 gate2128(.a(gate261inter12), .b(gate261inter1), .O(G782));

  xor2  gate1597(.a(G765), .b(G764), .O(gate262inter0));
  nand2 gate1598(.a(gate262inter0), .b(s_150), .O(gate262inter1));
  and2  gate1599(.a(G765), .b(G764), .O(gate262inter2));
  inv1  gate1600(.a(s_150), .O(gate262inter3));
  inv1  gate1601(.a(s_151), .O(gate262inter4));
  nand2 gate1602(.a(gate262inter4), .b(gate262inter3), .O(gate262inter5));
  nor2  gate1603(.a(gate262inter5), .b(gate262inter2), .O(gate262inter6));
  inv1  gate1604(.a(G764), .O(gate262inter7));
  inv1  gate1605(.a(G765), .O(gate262inter8));
  nand2 gate1606(.a(gate262inter8), .b(gate262inter7), .O(gate262inter9));
  nand2 gate1607(.a(s_151), .b(gate262inter3), .O(gate262inter10));
  nor2  gate1608(.a(gate262inter10), .b(gate262inter9), .O(gate262inter11));
  nor2  gate1609(.a(gate262inter11), .b(gate262inter6), .O(gate262inter12));
  nand2 gate1610(.a(gate262inter12), .b(gate262inter1), .O(G785));
nand2 gate263( .a(G766), .b(G767), .O(G788) );
nand2 gate264( .a(G768), .b(G769), .O(G791) );

  xor2  gate1009(.a(G770), .b(G642), .O(gate265inter0));
  nand2 gate1010(.a(gate265inter0), .b(s_66), .O(gate265inter1));
  and2  gate1011(.a(G770), .b(G642), .O(gate265inter2));
  inv1  gate1012(.a(s_66), .O(gate265inter3));
  inv1  gate1013(.a(s_67), .O(gate265inter4));
  nand2 gate1014(.a(gate265inter4), .b(gate265inter3), .O(gate265inter5));
  nor2  gate1015(.a(gate265inter5), .b(gate265inter2), .O(gate265inter6));
  inv1  gate1016(.a(G642), .O(gate265inter7));
  inv1  gate1017(.a(G770), .O(gate265inter8));
  nand2 gate1018(.a(gate265inter8), .b(gate265inter7), .O(gate265inter9));
  nand2 gate1019(.a(s_67), .b(gate265inter3), .O(gate265inter10));
  nor2  gate1020(.a(gate265inter10), .b(gate265inter9), .O(gate265inter11));
  nor2  gate1021(.a(gate265inter11), .b(gate265inter6), .O(gate265inter12));
  nand2 gate1022(.a(gate265inter12), .b(gate265inter1), .O(G794));
nand2 gate266( .a(G645), .b(G773), .O(G797) );
nand2 gate267( .a(G648), .b(G776), .O(G800) );

  xor2  gate2493(.a(G779), .b(G651), .O(gate268inter0));
  nand2 gate2494(.a(gate268inter0), .b(s_278), .O(gate268inter1));
  and2  gate2495(.a(G779), .b(G651), .O(gate268inter2));
  inv1  gate2496(.a(s_278), .O(gate268inter3));
  inv1  gate2497(.a(s_279), .O(gate268inter4));
  nand2 gate2498(.a(gate268inter4), .b(gate268inter3), .O(gate268inter5));
  nor2  gate2499(.a(gate268inter5), .b(gate268inter2), .O(gate268inter6));
  inv1  gate2500(.a(G651), .O(gate268inter7));
  inv1  gate2501(.a(G779), .O(gate268inter8));
  nand2 gate2502(.a(gate268inter8), .b(gate268inter7), .O(gate268inter9));
  nand2 gate2503(.a(s_279), .b(gate268inter3), .O(gate268inter10));
  nor2  gate2504(.a(gate268inter10), .b(gate268inter9), .O(gate268inter11));
  nor2  gate2505(.a(gate268inter11), .b(gate268inter6), .O(gate268inter12));
  nand2 gate2506(.a(gate268inter12), .b(gate268inter1), .O(G803));

  xor2  gate785(.a(G782), .b(G654), .O(gate269inter0));
  nand2 gate786(.a(gate269inter0), .b(s_34), .O(gate269inter1));
  and2  gate787(.a(G782), .b(G654), .O(gate269inter2));
  inv1  gate788(.a(s_34), .O(gate269inter3));
  inv1  gate789(.a(s_35), .O(gate269inter4));
  nand2 gate790(.a(gate269inter4), .b(gate269inter3), .O(gate269inter5));
  nor2  gate791(.a(gate269inter5), .b(gate269inter2), .O(gate269inter6));
  inv1  gate792(.a(G654), .O(gate269inter7));
  inv1  gate793(.a(G782), .O(gate269inter8));
  nand2 gate794(.a(gate269inter8), .b(gate269inter7), .O(gate269inter9));
  nand2 gate795(.a(s_35), .b(gate269inter3), .O(gate269inter10));
  nor2  gate796(.a(gate269inter10), .b(gate269inter9), .O(gate269inter11));
  nor2  gate797(.a(gate269inter11), .b(gate269inter6), .O(gate269inter12));
  nand2 gate798(.a(gate269inter12), .b(gate269inter1), .O(G806));
nand2 gate270( .a(G657), .b(G785), .O(G809) );

  xor2  gate869(.a(G788), .b(G660), .O(gate271inter0));
  nand2 gate870(.a(gate271inter0), .b(s_46), .O(gate271inter1));
  and2  gate871(.a(G788), .b(G660), .O(gate271inter2));
  inv1  gate872(.a(s_46), .O(gate271inter3));
  inv1  gate873(.a(s_47), .O(gate271inter4));
  nand2 gate874(.a(gate271inter4), .b(gate271inter3), .O(gate271inter5));
  nor2  gate875(.a(gate271inter5), .b(gate271inter2), .O(gate271inter6));
  inv1  gate876(.a(G660), .O(gate271inter7));
  inv1  gate877(.a(G788), .O(gate271inter8));
  nand2 gate878(.a(gate271inter8), .b(gate271inter7), .O(gate271inter9));
  nand2 gate879(.a(s_47), .b(gate271inter3), .O(gate271inter10));
  nor2  gate880(.a(gate271inter10), .b(gate271inter9), .O(gate271inter11));
  nor2  gate881(.a(gate271inter11), .b(gate271inter6), .O(gate271inter12));
  nand2 gate882(.a(gate271inter12), .b(gate271inter1), .O(G812));
nand2 gate272( .a(G663), .b(G791), .O(G815) );

  xor2  gate1205(.a(G794), .b(G642), .O(gate273inter0));
  nand2 gate1206(.a(gate273inter0), .b(s_94), .O(gate273inter1));
  and2  gate1207(.a(G794), .b(G642), .O(gate273inter2));
  inv1  gate1208(.a(s_94), .O(gate273inter3));
  inv1  gate1209(.a(s_95), .O(gate273inter4));
  nand2 gate1210(.a(gate273inter4), .b(gate273inter3), .O(gate273inter5));
  nor2  gate1211(.a(gate273inter5), .b(gate273inter2), .O(gate273inter6));
  inv1  gate1212(.a(G642), .O(gate273inter7));
  inv1  gate1213(.a(G794), .O(gate273inter8));
  nand2 gate1214(.a(gate273inter8), .b(gate273inter7), .O(gate273inter9));
  nand2 gate1215(.a(s_95), .b(gate273inter3), .O(gate273inter10));
  nor2  gate1216(.a(gate273inter10), .b(gate273inter9), .O(gate273inter11));
  nor2  gate1217(.a(gate273inter11), .b(gate273inter6), .O(gate273inter12));
  nand2 gate1218(.a(gate273inter12), .b(gate273inter1), .O(G818));
nand2 gate274( .a(G770), .b(G794), .O(G819) );
nand2 gate275( .a(G645), .b(G797), .O(G820) );

  xor2  gate1177(.a(G797), .b(G773), .O(gate276inter0));
  nand2 gate1178(.a(gate276inter0), .b(s_90), .O(gate276inter1));
  and2  gate1179(.a(G797), .b(G773), .O(gate276inter2));
  inv1  gate1180(.a(s_90), .O(gate276inter3));
  inv1  gate1181(.a(s_91), .O(gate276inter4));
  nand2 gate1182(.a(gate276inter4), .b(gate276inter3), .O(gate276inter5));
  nor2  gate1183(.a(gate276inter5), .b(gate276inter2), .O(gate276inter6));
  inv1  gate1184(.a(G773), .O(gate276inter7));
  inv1  gate1185(.a(G797), .O(gate276inter8));
  nand2 gate1186(.a(gate276inter8), .b(gate276inter7), .O(gate276inter9));
  nand2 gate1187(.a(s_91), .b(gate276inter3), .O(gate276inter10));
  nor2  gate1188(.a(gate276inter10), .b(gate276inter9), .O(gate276inter11));
  nor2  gate1189(.a(gate276inter11), .b(gate276inter6), .O(gate276inter12));
  nand2 gate1190(.a(gate276inter12), .b(gate276inter1), .O(G821));
nand2 gate277( .a(G648), .b(G800), .O(G822) );
nand2 gate278( .a(G776), .b(G800), .O(G823) );

  xor2  gate995(.a(G803), .b(G651), .O(gate279inter0));
  nand2 gate996(.a(gate279inter0), .b(s_64), .O(gate279inter1));
  and2  gate997(.a(G803), .b(G651), .O(gate279inter2));
  inv1  gate998(.a(s_64), .O(gate279inter3));
  inv1  gate999(.a(s_65), .O(gate279inter4));
  nand2 gate1000(.a(gate279inter4), .b(gate279inter3), .O(gate279inter5));
  nor2  gate1001(.a(gate279inter5), .b(gate279inter2), .O(gate279inter6));
  inv1  gate1002(.a(G651), .O(gate279inter7));
  inv1  gate1003(.a(G803), .O(gate279inter8));
  nand2 gate1004(.a(gate279inter8), .b(gate279inter7), .O(gate279inter9));
  nand2 gate1005(.a(s_65), .b(gate279inter3), .O(gate279inter10));
  nor2  gate1006(.a(gate279inter10), .b(gate279inter9), .O(gate279inter11));
  nor2  gate1007(.a(gate279inter11), .b(gate279inter6), .O(gate279inter12));
  nand2 gate1008(.a(gate279inter12), .b(gate279inter1), .O(G824));
nand2 gate280( .a(G779), .b(G803), .O(G825) );
nand2 gate281( .a(G654), .b(G806), .O(G826) );
nand2 gate282( .a(G782), .b(G806), .O(G827) );

  xor2  gate2073(.a(G809), .b(G657), .O(gate283inter0));
  nand2 gate2074(.a(gate283inter0), .b(s_218), .O(gate283inter1));
  and2  gate2075(.a(G809), .b(G657), .O(gate283inter2));
  inv1  gate2076(.a(s_218), .O(gate283inter3));
  inv1  gate2077(.a(s_219), .O(gate283inter4));
  nand2 gate2078(.a(gate283inter4), .b(gate283inter3), .O(gate283inter5));
  nor2  gate2079(.a(gate283inter5), .b(gate283inter2), .O(gate283inter6));
  inv1  gate2080(.a(G657), .O(gate283inter7));
  inv1  gate2081(.a(G809), .O(gate283inter8));
  nand2 gate2082(.a(gate283inter8), .b(gate283inter7), .O(gate283inter9));
  nand2 gate2083(.a(s_219), .b(gate283inter3), .O(gate283inter10));
  nor2  gate2084(.a(gate283inter10), .b(gate283inter9), .O(gate283inter11));
  nor2  gate2085(.a(gate283inter11), .b(gate283inter6), .O(gate283inter12));
  nand2 gate2086(.a(gate283inter12), .b(gate283inter1), .O(G828));
nand2 gate284( .a(G785), .b(G809), .O(G829) );

  xor2  gate645(.a(G812), .b(G660), .O(gate285inter0));
  nand2 gate646(.a(gate285inter0), .b(s_14), .O(gate285inter1));
  and2  gate647(.a(G812), .b(G660), .O(gate285inter2));
  inv1  gate648(.a(s_14), .O(gate285inter3));
  inv1  gate649(.a(s_15), .O(gate285inter4));
  nand2 gate650(.a(gate285inter4), .b(gate285inter3), .O(gate285inter5));
  nor2  gate651(.a(gate285inter5), .b(gate285inter2), .O(gate285inter6));
  inv1  gate652(.a(G660), .O(gate285inter7));
  inv1  gate653(.a(G812), .O(gate285inter8));
  nand2 gate654(.a(gate285inter8), .b(gate285inter7), .O(gate285inter9));
  nand2 gate655(.a(s_15), .b(gate285inter3), .O(gate285inter10));
  nor2  gate656(.a(gate285inter10), .b(gate285inter9), .O(gate285inter11));
  nor2  gate657(.a(gate285inter11), .b(gate285inter6), .O(gate285inter12));
  nand2 gate658(.a(gate285inter12), .b(gate285inter1), .O(G830));

  xor2  gate1415(.a(G812), .b(G788), .O(gate286inter0));
  nand2 gate1416(.a(gate286inter0), .b(s_124), .O(gate286inter1));
  and2  gate1417(.a(G812), .b(G788), .O(gate286inter2));
  inv1  gate1418(.a(s_124), .O(gate286inter3));
  inv1  gate1419(.a(s_125), .O(gate286inter4));
  nand2 gate1420(.a(gate286inter4), .b(gate286inter3), .O(gate286inter5));
  nor2  gate1421(.a(gate286inter5), .b(gate286inter2), .O(gate286inter6));
  inv1  gate1422(.a(G788), .O(gate286inter7));
  inv1  gate1423(.a(G812), .O(gate286inter8));
  nand2 gate1424(.a(gate286inter8), .b(gate286inter7), .O(gate286inter9));
  nand2 gate1425(.a(s_125), .b(gate286inter3), .O(gate286inter10));
  nor2  gate1426(.a(gate286inter10), .b(gate286inter9), .O(gate286inter11));
  nor2  gate1427(.a(gate286inter11), .b(gate286inter6), .O(gate286inter12));
  nand2 gate1428(.a(gate286inter12), .b(gate286inter1), .O(G831));

  xor2  gate1891(.a(G815), .b(G663), .O(gate287inter0));
  nand2 gate1892(.a(gate287inter0), .b(s_192), .O(gate287inter1));
  and2  gate1893(.a(G815), .b(G663), .O(gate287inter2));
  inv1  gate1894(.a(s_192), .O(gate287inter3));
  inv1  gate1895(.a(s_193), .O(gate287inter4));
  nand2 gate1896(.a(gate287inter4), .b(gate287inter3), .O(gate287inter5));
  nor2  gate1897(.a(gate287inter5), .b(gate287inter2), .O(gate287inter6));
  inv1  gate1898(.a(G663), .O(gate287inter7));
  inv1  gate1899(.a(G815), .O(gate287inter8));
  nand2 gate1900(.a(gate287inter8), .b(gate287inter7), .O(gate287inter9));
  nand2 gate1901(.a(s_193), .b(gate287inter3), .O(gate287inter10));
  nor2  gate1902(.a(gate287inter10), .b(gate287inter9), .O(gate287inter11));
  nor2  gate1903(.a(gate287inter11), .b(gate287inter6), .O(gate287inter12));
  nand2 gate1904(.a(gate287inter12), .b(gate287inter1), .O(G832));
nand2 gate288( .a(G791), .b(G815), .O(G833) );
nand2 gate289( .a(G818), .b(G819), .O(G834) );

  xor2  gate1821(.a(G821), .b(G820), .O(gate290inter0));
  nand2 gate1822(.a(gate290inter0), .b(s_182), .O(gate290inter1));
  and2  gate1823(.a(G821), .b(G820), .O(gate290inter2));
  inv1  gate1824(.a(s_182), .O(gate290inter3));
  inv1  gate1825(.a(s_183), .O(gate290inter4));
  nand2 gate1826(.a(gate290inter4), .b(gate290inter3), .O(gate290inter5));
  nor2  gate1827(.a(gate290inter5), .b(gate290inter2), .O(gate290inter6));
  inv1  gate1828(.a(G820), .O(gate290inter7));
  inv1  gate1829(.a(G821), .O(gate290inter8));
  nand2 gate1830(.a(gate290inter8), .b(gate290inter7), .O(gate290inter9));
  nand2 gate1831(.a(s_183), .b(gate290inter3), .O(gate290inter10));
  nor2  gate1832(.a(gate290inter10), .b(gate290inter9), .O(gate290inter11));
  nor2  gate1833(.a(gate290inter11), .b(gate290inter6), .O(gate290inter12));
  nand2 gate1834(.a(gate290inter12), .b(gate290inter1), .O(G847));
nand2 gate291( .a(G822), .b(G823), .O(G860) );
nand2 gate292( .a(G824), .b(G825), .O(G873) );

  xor2  gate2087(.a(G829), .b(G828), .O(gate293inter0));
  nand2 gate2088(.a(gate293inter0), .b(s_220), .O(gate293inter1));
  and2  gate2089(.a(G829), .b(G828), .O(gate293inter2));
  inv1  gate2090(.a(s_220), .O(gate293inter3));
  inv1  gate2091(.a(s_221), .O(gate293inter4));
  nand2 gate2092(.a(gate293inter4), .b(gate293inter3), .O(gate293inter5));
  nor2  gate2093(.a(gate293inter5), .b(gate293inter2), .O(gate293inter6));
  inv1  gate2094(.a(G828), .O(gate293inter7));
  inv1  gate2095(.a(G829), .O(gate293inter8));
  nand2 gate2096(.a(gate293inter8), .b(gate293inter7), .O(gate293inter9));
  nand2 gate2097(.a(s_221), .b(gate293inter3), .O(gate293inter10));
  nor2  gate2098(.a(gate293inter10), .b(gate293inter9), .O(gate293inter11));
  nor2  gate2099(.a(gate293inter11), .b(gate293inter6), .O(gate293inter12));
  nand2 gate2100(.a(gate293inter12), .b(gate293inter1), .O(G886));

  xor2  gate1863(.a(G833), .b(G832), .O(gate294inter0));
  nand2 gate1864(.a(gate294inter0), .b(s_188), .O(gate294inter1));
  and2  gate1865(.a(G833), .b(G832), .O(gate294inter2));
  inv1  gate1866(.a(s_188), .O(gate294inter3));
  inv1  gate1867(.a(s_189), .O(gate294inter4));
  nand2 gate1868(.a(gate294inter4), .b(gate294inter3), .O(gate294inter5));
  nor2  gate1869(.a(gate294inter5), .b(gate294inter2), .O(gate294inter6));
  inv1  gate1870(.a(G832), .O(gate294inter7));
  inv1  gate1871(.a(G833), .O(gate294inter8));
  nand2 gate1872(.a(gate294inter8), .b(gate294inter7), .O(gate294inter9));
  nand2 gate1873(.a(s_189), .b(gate294inter3), .O(gate294inter10));
  nor2  gate1874(.a(gate294inter10), .b(gate294inter9), .O(gate294inter11));
  nor2  gate1875(.a(gate294inter11), .b(gate294inter6), .O(gate294inter12));
  nand2 gate1876(.a(gate294inter12), .b(gate294inter1), .O(G899));

  xor2  gate1401(.a(G831), .b(G830), .O(gate295inter0));
  nand2 gate1402(.a(gate295inter0), .b(s_122), .O(gate295inter1));
  and2  gate1403(.a(G831), .b(G830), .O(gate295inter2));
  inv1  gate1404(.a(s_122), .O(gate295inter3));
  inv1  gate1405(.a(s_123), .O(gate295inter4));
  nand2 gate1406(.a(gate295inter4), .b(gate295inter3), .O(gate295inter5));
  nor2  gate1407(.a(gate295inter5), .b(gate295inter2), .O(gate295inter6));
  inv1  gate1408(.a(G830), .O(gate295inter7));
  inv1  gate1409(.a(G831), .O(gate295inter8));
  nand2 gate1410(.a(gate295inter8), .b(gate295inter7), .O(gate295inter9));
  nand2 gate1411(.a(s_123), .b(gate295inter3), .O(gate295inter10));
  nor2  gate1412(.a(gate295inter10), .b(gate295inter9), .O(gate295inter11));
  nor2  gate1413(.a(gate295inter11), .b(gate295inter6), .O(gate295inter12));
  nand2 gate1414(.a(gate295inter12), .b(gate295inter1), .O(G912));
nand2 gate296( .a(G826), .b(G827), .O(G925) );
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );
nand2 gate387( .a(G1), .b(G1036), .O(G1132) );

  xor2  gate2017(.a(G1039), .b(G2), .O(gate388inter0));
  nand2 gate2018(.a(gate388inter0), .b(s_210), .O(gate388inter1));
  and2  gate2019(.a(G1039), .b(G2), .O(gate388inter2));
  inv1  gate2020(.a(s_210), .O(gate388inter3));
  inv1  gate2021(.a(s_211), .O(gate388inter4));
  nand2 gate2022(.a(gate388inter4), .b(gate388inter3), .O(gate388inter5));
  nor2  gate2023(.a(gate388inter5), .b(gate388inter2), .O(gate388inter6));
  inv1  gate2024(.a(G2), .O(gate388inter7));
  inv1  gate2025(.a(G1039), .O(gate388inter8));
  nand2 gate2026(.a(gate388inter8), .b(gate388inter7), .O(gate388inter9));
  nand2 gate2027(.a(s_211), .b(gate388inter3), .O(gate388inter10));
  nor2  gate2028(.a(gate388inter10), .b(gate388inter9), .O(gate388inter11));
  nor2  gate2029(.a(gate388inter11), .b(gate388inter6), .O(gate388inter12));
  nand2 gate2030(.a(gate388inter12), .b(gate388inter1), .O(G1135));

  xor2  gate1793(.a(G1042), .b(G3), .O(gate389inter0));
  nand2 gate1794(.a(gate389inter0), .b(s_178), .O(gate389inter1));
  and2  gate1795(.a(G1042), .b(G3), .O(gate389inter2));
  inv1  gate1796(.a(s_178), .O(gate389inter3));
  inv1  gate1797(.a(s_179), .O(gate389inter4));
  nand2 gate1798(.a(gate389inter4), .b(gate389inter3), .O(gate389inter5));
  nor2  gate1799(.a(gate389inter5), .b(gate389inter2), .O(gate389inter6));
  inv1  gate1800(.a(G3), .O(gate389inter7));
  inv1  gate1801(.a(G1042), .O(gate389inter8));
  nand2 gate1802(.a(gate389inter8), .b(gate389inter7), .O(gate389inter9));
  nand2 gate1803(.a(s_179), .b(gate389inter3), .O(gate389inter10));
  nor2  gate1804(.a(gate389inter10), .b(gate389inter9), .O(gate389inter11));
  nor2  gate1805(.a(gate389inter11), .b(gate389inter6), .O(gate389inter12));
  nand2 gate1806(.a(gate389inter12), .b(gate389inter1), .O(G1138));
nand2 gate390( .a(G4), .b(G1045), .O(G1141) );
nand2 gate391( .a(G5), .b(G1048), .O(G1144) );
nand2 gate392( .a(G6), .b(G1051), .O(G1147) );

  xor2  gate925(.a(G1054), .b(G7), .O(gate393inter0));
  nand2 gate926(.a(gate393inter0), .b(s_54), .O(gate393inter1));
  and2  gate927(.a(G1054), .b(G7), .O(gate393inter2));
  inv1  gate928(.a(s_54), .O(gate393inter3));
  inv1  gate929(.a(s_55), .O(gate393inter4));
  nand2 gate930(.a(gate393inter4), .b(gate393inter3), .O(gate393inter5));
  nor2  gate931(.a(gate393inter5), .b(gate393inter2), .O(gate393inter6));
  inv1  gate932(.a(G7), .O(gate393inter7));
  inv1  gate933(.a(G1054), .O(gate393inter8));
  nand2 gate934(.a(gate393inter8), .b(gate393inter7), .O(gate393inter9));
  nand2 gate935(.a(s_55), .b(gate393inter3), .O(gate393inter10));
  nor2  gate936(.a(gate393inter10), .b(gate393inter9), .O(gate393inter11));
  nor2  gate937(.a(gate393inter11), .b(gate393inter6), .O(gate393inter12));
  nand2 gate938(.a(gate393inter12), .b(gate393inter1), .O(G1150));
nand2 gate394( .a(G8), .b(G1057), .O(G1153) );
nand2 gate395( .a(G9), .b(G1060), .O(G1156) );
nand2 gate396( .a(G10), .b(G1063), .O(G1159) );

  xor2  gate1975(.a(G1066), .b(G11), .O(gate397inter0));
  nand2 gate1976(.a(gate397inter0), .b(s_204), .O(gate397inter1));
  and2  gate1977(.a(G1066), .b(G11), .O(gate397inter2));
  inv1  gate1978(.a(s_204), .O(gate397inter3));
  inv1  gate1979(.a(s_205), .O(gate397inter4));
  nand2 gate1980(.a(gate397inter4), .b(gate397inter3), .O(gate397inter5));
  nor2  gate1981(.a(gate397inter5), .b(gate397inter2), .O(gate397inter6));
  inv1  gate1982(.a(G11), .O(gate397inter7));
  inv1  gate1983(.a(G1066), .O(gate397inter8));
  nand2 gate1984(.a(gate397inter8), .b(gate397inter7), .O(gate397inter9));
  nand2 gate1985(.a(s_205), .b(gate397inter3), .O(gate397inter10));
  nor2  gate1986(.a(gate397inter10), .b(gate397inter9), .O(gate397inter11));
  nor2  gate1987(.a(gate397inter11), .b(gate397inter6), .O(gate397inter12));
  nand2 gate1988(.a(gate397inter12), .b(gate397inter1), .O(G1162));

  xor2  gate1919(.a(G1069), .b(G12), .O(gate398inter0));
  nand2 gate1920(.a(gate398inter0), .b(s_196), .O(gate398inter1));
  and2  gate1921(.a(G1069), .b(G12), .O(gate398inter2));
  inv1  gate1922(.a(s_196), .O(gate398inter3));
  inv1  gate1923(.a(s_197), .O(gate398inter4));
  nand2 gate1924(.a(gate398inter4), .b(gate398inter3), .O(gate398inter5));
  nor2  gate1925(.a(gate398inter5), .b(gate398inter2), .O(gate398inter6));
  inv1  gate1926(.a(G12), .O(gate398inter7));
  inv1  gate1927(.a(G1069), .O(gate398inter8));
  nand2 gate1928(.a(gate398inter8), .b(gate398inter7), .O(gate398inter9));
  nand2 gate1929(.a(s_197), .b(gate398inter3), .O(gate398inter10));
  nor2  gate1930(.a(gate398inter10), .b(gate398inter9), .O(gate398inter11));
  nor2  gate1931(.a(gate398inter11), .b(gate398inter6), .O(gate398inter12));
  nand2 gate1932(.a(gate398inter12), .b(gate398inter1), .O(G1165));
nand2 gate399( .a(G13), .b(G1072), .O(G1168) );

  xor2  gate1989(.a(G1075), .b(G14), .O(gate400inter0));
  nand2 gate1990(.a(gate400inter0), .b(s_206), .O(gate400inter1));
  and2  gate1991(.a(G1075), .b(G14), .O(gate400inter2));
  inv1  gate1992(.a(s_206), .O(gate400inter3));
  inv1  gate1993(.a(s_207), .O(gate400inter4));
  nand2 gate1994(.a(gate400inter4), .b(gate400inter3), .O(gate400inter5));
  nor2  gate1995(.a(gate400inter5), .b(gate400inter2), .O(gate400inter6));
  inv1  gate1996(.a(G14), .O(gate400inter7));
  inv1  gate1997(.a(G1075), .O(gate400inter8));
  nand2 gate1998(.a(gate400inter8), .b(gate400inter7), .O(gate400inter9));
  nand2 gate1999(.a(s_207), .b(gate400inter3), .O(gate400inter10));
  nor2  gate2000(.a(gate400inter10), .b(gate400inter9), .O(gate400inter11));
  nor2  gate2001(.a(gate400inter11), .b(gate400inter6), .O(gate400inter12));
  nand2 gate2002(.a(gate400inter12), .b(gate400inter1), .O(G1171));
nand2 gate401( .a(G15), .b(G1078), .O(G1174) );
nand2 gate402( .a(G16), .b(G1081), .O(G1177) );
nand2 gate403( .a(G17), .b(G1084), .O(G1180) );
nand2 gate404( .a(G18), .b(G1087), .O(G1183) );
nand2 gate405( .a(G19), .b(G1090), .O(G1186) );
nand2 gate406( .a(G20), .b(G1093), .O(G1189) );
nand2 gate407( .a(G21), .b(G1096), .O(G1192) );
nand2 gate408( .a(G22), .b(G1099), .O(G1195) );
nand2 gate409( .a(G23), .b(G1102), .O(G1198) );
nand2 gate410( .a(G24), .b(G1105), .O(G1201) );
nand2 gate411( .a(G25), .b(G1108), .O(G1204) );
nand2 gate412( .a(G26), .b(G1111), .O(G1207) );

  xor2  gate1667(.a(G1114), .b(G27), .O(gate413inter0));
  nand2 gate1668(.a(gate413inter0), .b(s_160), .O(gate413inter1));
  and2  gate1669(.a(G1114), .b(G27), .O(gate413inter2));
  inv1  gate1670(.a(s_160), .O(gate413inter3));
  inv1  gate1671(.a(s_161), .O(gate413inter4));
  nand2 gate1672(.a(gate413inter4), .b(gate413inter3), .O(gate413inter5));
  nor2  gate1673(.a(gate413inter5), .b(gate413inter2), .O(gate413inter6));
  inv1  gate1674(.a(G27), .O(gate413inter7));
  inv1  gate1675(.a(G1114), .O(gate413inter8));
  nand2 gate1676(.a(gate413inter8), .b(gate413inter7), .O(gate413inter9));
  nand2 gate1677(.a(s_161), .b(gate413inter3), .O(gate413inter10));
  nor2  gate1678(.a(gate413inter10), .b(gate413inter9), .O(gate413inter11));
  nor2  gate1679(.a(gate413inter11), .b(gate413inter6), .O(gate413inter12));
  nand2 gate1680(.a(gate413inter12), .b(gate413inter1), .O(G1210));
nand2 gate414( .a(G28), .b(G1117), .O(G1213) );
nand2 gate415( .a(G29), .b(G1120), .O(G1216) );

  xor2  gate1807(.a(G1123), .b(G30), .O(gate416inter0));
  nand2 gate1808(.a(gate416inter0), .b(s_180), .O(gate416inter1));
  and2  gate1809(.a(G1123), .b(G30), .O(gate416inter2));
  inv1  gate1810(.a(s_180), .O(gate416inter3));
  inv1  gate1811(.a(s_181), .O(gate416inter4));
  nand2 gate1812(.a(gate416inter4), .b(gate416inter3), .O(gate416inter5));
  nor2  gate1813(.a(gate416inter5), .b(gate416inter2), .O(gate416inter6));
  inv1  gate1814(.a(G30), .O(gate416inter7));
  inv1  gate1815(.a(G1123), .O(gate416inter8));
  nand2 gate1816(.a(gate416inter8), .b(gate416inter7), .O(gate416inter9));
  nand2 gate1817(.a(s_181), .b(gate416inter3), .O(gate416inter10));
  nor2  gate1818(.a(gate416inter10), .b(gate416inter9), .O(gate416inter11));
  nor2  gate1819(.a(gate416inter11), .b(gate416inter6), .O(gate416inter12));
  nand2 gate1820(.a(gate416inter12), .b(gate416inter1), .O(G1219));

  xor2  gate2437(.a(G1126), .b(G31), .O(gate417inter0));
  nand2 gate2438(.a(gate417inter0), .b(s_270), .O(gate417inter1));
  and2  gate2439(.a(G1126), .b(G31), .O(gate417inter2));
  inv1  gate2440(.a(s_270), .O(gate417inter3));
  inv1  gate2441(.a(s_271), .O(gate417inter4));
  nand2 gate2442(.a(gate417inter4), .b(gate417inter3), .O(gate417inter5));
  nor2  gate2443(.a(gate417inter5), .b(gate417inter2), .O(gate417inter6));
  inv1  gate2444(.a(G31), .O(gate417inter7));
  inv1  gate2445(.a(G1126), .O(gate417inter8));
  nand2 gate2446(.a(gate417inter8), .b(gate417inter7), .O(gate417inter9));
  nand2 gate2447(.a(s_271), .b(gate417inter3), .O(gate417inter10));
  nor2  gate2448(.a(gate417inter10), .b(gate417inter9), .O(gate417inter11));
  nor2  gate2449(.a(gate417inter11), .b(gate417inter6), .O(gate417inter12));
  nand2 gate2450(.a(gate417inter12), .b(gate417inter1), .O(G1222));

  xor2  gate1653(.a(G1129), .b(G32), .O(gate418inter0));
  nand2 gate1654(.a(gate418inter0), .b(s_158), .O(gate418inter1));
  and2  gate1655(.a(G1129), .b(G32), .O(gate418inter2));
  inv1  gate1656(.a(s_158), .O(gate418inter3));
  inv1  gate1657(.a(s_159), .O(gate418inter4));
  nand2 gate1658(.a(gate418inter4), .b(gate418inter3), .O(gate418inter5));
  nor2  gate1659(.a(gate418inter5), .b(gate418inter2), .O(gate418inter6));
  inv1  gate1660(.a(G32), .O(gate418inter7));
  inv1  gate1661(.a(G1129), .O(gate418inter8));
  nand2 gate1662(.a(gate418inter8), .b(gate418inter7), .O(gate418inter9));
  nand2 gate1663(.a(s_159), .b(gate418inter3), .O(gate418inter10));
  nor2  gate1664(.a(gate418inter10), .b(gate418inter9), .O(gate418inter11));
  nor2  gate1665(.a(gate418inter11), .b(gate418inter6), .O(gate418inter12));
  nand2 gate1666(.a(gate418inter12), .b(gate418inter1), .O(G1225));
nand2 gate419( .a(G1), .b(G1132), .O(G1228) );
nand2 gate420( .a(G1036), .b(G1132), .O(G1229) );
nand2 gate421( .a(G2), .b(G1135), .O(G1230) );

  xor2  gate953(.a(G1135), .b(G1039), .O(gate422inter0));
  nand2 gate954(.a(gate422inter0), .b(s_58), .O(gate422inter1));
  and2  gate955(.a(G1135), .b(G1039), .O(gate422inter2));
  inv1  gate956(.a(s_58), .O(gate422inter3));
  inv1  gate957(.a(s_59), .O(gate422inter4));
  nand2 gate958(.a(gate422inter4), .b(gate422inter3), .O(gate422inter5));
  nor2  gate959(.a(gate422inter5), .b(gate422inter2), .O(gate422inter6));
  inv1  gate960(.a(G1039), .O(gate422inter7));
  inv1  gate961(.a(G1135), .O(gate422inter8));
  nand2 gate962(.a(gate422inter8), .b(gate422inter7), .O(gate422inter9));
  nand2 gate963(.a(s_59), .b(gate422inter3), .O(gate422inter10));
  nor2  gate964(.a(gate422inter10), .b(gate422inter9), .O(gate422inter11));
  nor2  gate965(.a(gate422inter11), .b(gate422inter6), .O(gate422inter12));
  nand2 gate966(.a(gate422inter12), .b(gate422inter1), .O(G1231));

  xor2  gate855(.a(G1138), .b(G3), .O(gate423inter0));
  nand2 gate856(.a(gate423inter0), .b(s_44), .O(gate423inter1));
  and2  gate857(.a(G1138), .b(G3), .O(gate423inter2));
  inv1  gate858(.a(s_44), .O(gate423inter3));
  inv1  gate859(.a(s_45), .O(gate423inter4));
  nand2 gate860(.a(gate423inter4), .b(gate423inter3), .O(gate423inter5));
  nor2  gate861(.a(gate423inter5), .b(gate423inter2), .O(gate423inter6));
  inv1  gate862(.a(G3), .O(gate423inter7));
  inv1  gate863(.a(G1138), .O(gate423inter8));
  nand2 gate864(.a(gate423inter8), .b(gate423inter7), .O(gate423inter9));
  nand2 gate865(.a(s_45), .b(gate423inter3), .O(gate423inter10));
  nor2  gate866(.a(gate423inter10), .b(gate423inter9), .O(gate423inter11));
  nor2  gate867(.a(gate423inter11), .b(gate423inter6), .O(gate423inter12));
  nand2 gate868(.a(gate423inter12), .b(gate423inter1), .O(G1232));
nand2 gate424( .a(G1042), .b(G1138), .O(G1233) );

  xor2  gate1359(.a(G1141), .b(G4), .O(gate425inter0));
  nand2 gate1360(.a(gate425inter0), .b(s_116), .O(gate425inter1));
  and2  gate1361(.a(G1141), .b(G4), .O(gate425inter2));
  inv1  gate1362(.a(s_116), .O(gate425inter3));
  inv1  gate1363(.a(s_117), .O(gate425inter4));
  nand2 gate1364(.a(gate425inter4), .b(gate425inter3), .O(gate425inter5));
  nor2  gate1365(.a(gate425inter5), .b(gate425inter2), .O(gate425inter6));
  inv1  gate1366(.a(G4), .O(gate425inter7));
  inv1  gate1367(.a(G1141), .O(gate425inter8));
  nand2 gate1368(.a(gate425inter8), .b(gate425inter7), .O(gate425inter9));
  nand2 gate1369(.a(s_117), .b(gate425inter3), .O(gate425inter10));
  nor2  gate1370(.a(gate425inter10), .b(gate425inter9), .O(gate425inter11));
  nor2  gate1371(.a(gate425inter11), .b(gate425inter6), .O(gate425inter12));
  nand2 gate1372(.a(gate425inter12), .b(gate425inter1), .O(G1234));
nand2 gate426( .a(G1045), .b(G1141), .O(G1235) );
nand2 gate427( .a(G5), .b(G1144), .O(G1236) );
nand2 gate428( .a(G1048), .b(G1144), .O(G1237) );
nand2 gate429( .a(G6), .b(G1147), .O(G1238) );
nand2 gate430( .a(G1051), .b(G1147), .O(G1239) );

  xor2  gate2619(.a(G1150), .b(G7), .O(gate431inter0));
  nand2 gate2620(.a(gate431inter0), .b(s_296), .O(gate431inter1));
  and2  gate2621(.a(G1150), .b(G7), .O(gate431inter2));
  inv1  gate2622(.a(s_296), .O(gate431inter3));
  inv1  gate2623(.a(s_297), .O(gate431inter4));
  nand2 gate2624(.a(gate431inter4), .b(gate431inter3), .O(gate431inter5));
  nor2  gate2625(.a(gate431inter5), .b(gate431inter2), .O(gate431inter6));
  inv1  gate2626(.a(G7), .O(gate431inter7));
  inv1  gate2627(.a(G1150), .O(gate431inter8));
  nand2 gate2628(.a(gate431inter8), .b(gate431inter7), .O(gate431inter9));
  nand2 gate2629(.a(s_297), .b(gate431inter3), .O(gate431inter10));
  nor2  gate2630(.a(gate431inter10), .b(gate431inter9), .O(gate431inter11));
  nor2  gate2631(.a(gate431inter11), .b(gate431inter6), .O(gate431inter12));
  nand2 gate2632(.a(gate431inter12), .b(gate431inter1), .O(G1240));
nand2 gate432( .a(G1054), .b(G1150), .O(G1241) );
nand2 gate433( .a(G8), .b(G1153), .O(G1242) );
nand2 gate434( .a(G1057), .b(G1153), .O(G1243) );
nand2 gate435( .a(G9), .b(G1156), .O(G1244) );

  xor2  gate1695(.a(G1156), .b(G1060), .O(gate436inter0));
  nand2 gate1696(.a(gate436inter0), .b(s_164), .O(gate436inter1));
  and2  gate1697(.a(G1156), .b(G1060), .O(gate436inter2));
  inv1  gate1698(.a(s_164), .O(gate436inter3));
  inv1  gate1699(.a(s_165), .O(gate436inter4));
  nand2 gate1700(.a(gate436inter4), .b(gate436inter3), .O(gate436inter5));
  nor2  gate1701(.a(gate436inter5), .b(gate436inter2), .O(gate436inter6));
  inv1  gate1702(.a(G1060), .O(gate436inter7));
  inv1  gate1703(.a(G1156), .O(gate436inter8));
  nand2 gate1704(.a(gate436inter8), .b(gate436inter7), .O(gate436inter9));
  nand2 gate1705(.a(s_165), .b(gate436inter3), .O(gate436inter10));
  nor2  gate1706(.a(gate436inter10), .b(gate436inter9), .O(gate436inter11));
  nor2  gate1707(.a(gate436inter11), .b(gate436inter6), .O(gate436inter12));
  nand2 gate1708(.a(gate436inter12), .b(gate436inter1), .O(G1245));

  xor2  gate1191(.a(G1159), .b(G10), .O(gate437inter0));
  nand2 gate1192(.a(gate437inter0), .b(s_92), .O(gate437inter1));
  and2  gate1193(.a(G1159), .b(G10), .O(gate437inter2));
  inv1  gate1194(.a(s_92), .O(gate437inter3));
  inv1  gate1195(.a(s_93), .O(gate437inter4));
  nand2 gate1196(.a(gate437inter4), .b(gate437inter3), .O(gate437inter5));
  nor2  gate1197(.a(gate437inter5), .b(gate437inter2), .O(gate437inter6));
  inv1  gate1198(.a(G10), .O(gate437inter7));
  inv1  gate1199(.a(G1159), .O(gate437inter8));
  nand2 gate1200(.a(gate437inter8), .b(gate437inter7), .O(gate437inter9));
  nand2 gate1201(.a(s_93), .b(gate437inter3), .O(gate437inter10));
  nor2  gate1202(.a(gate437inter10), .b(gate437inter9), .O(gate437inter11));
  nor2  gate1203(.a(gate437inter11), .b(gate437inter6), .O(gate437inter12));
  nand2 gate1204(.a(gate437inter12), .b(gate437inter1), .O(G1246));
nand2 gate438( .a(G1063), .b(G1159), .O(G1247) );
nand2 gate439( .a(G11), .b(G1162), .O(G1248) );
nand2 gate440( .a(G1066), .b(G1162), .O(G1249) );
nand2 gate441( .a(G12), .b(G1165), .O(G1250) );
nand2 gate442( .a(G1069), .b(G1165), .O(G1251) );
nand2 gate443( .a(G13), .b(G1168), .O(G1252) );

  xor2  gate813(.a(G1168), .b(G1072), .O(gate444inter0));
  nand2 gate814(.a(gate444inter0), .b(s_38), .O(gate444inter1));
  and2  gate815(.a(G1168), .b(G1072), .O(gate444inter2));
  inv1  gate816(.a(s_38), .O(gate444inter3));
  inv1  gate817(.a(s_39), .O(gate444inter4));
  nand2 gate818(.a(gate444inter4), .b(gate444inter3), .O(gate444inter5));
  nor2  gate819(.a(gate444inter5), .b(gate444inter2), .O(gate444inter6));
  inv1  gate820(.a(G1072), .O(gate444inter7));
  inv1  gate821(.a(G1168), .O(gate444inter8));
  nand2 gate822(.a(gate444inter8), .b(gate444inter7), .O(gate444inter9));
  nand2 gate823(.a(s_39), .b(gate444inter3), .O(gate444inter10));
  nor2  gate824(.a(gate444inter10), .b(gate444inter9), .O(gate444inter11));
  nor2  gate825(.a(gate444inter11), .b(gate444inter6), .O(gate444inter12));
  nand2 gate826(.a(gate444inter12), .b(gate444inter1), .O(G1253));
nand2 gate445( .a(G14), .b(G1171), .O(G1254) );
nand2 gate446( .a(G1075), .b(G1171), .O(G1255) );
nand2 gate447( .a(G15), .b(G1174), .O(G1256) );

  xor2  gate2409(.a(G1174), .b(G1078), .O(gate448inter0));
  nand2 gate2410(.a(gate448inter0), .b(s_266), .O(gate448inter1));
  and2  gate2411(.a(G1174), .b(G1078), .O(gate448inter2));
  inv1  gate2412(.a(s_266), .O(gate448inter3));
  inv1  gate2413(.a(s_267), .O(gate448inter4));
  nand2 gate2414(.a(gate448inter4), .b(gate448inter3), .O(gate448inter5));
  nor2  gate2415(.a(gate448inter5), .b(gate448inter2), .O(gate448inter6));
  inv1  gate2416(.a(G1078), .O(gate448inter7));
  inv1  gate2417(.a(G1174), .O(gate448inter8));
  nand2 gate2418(.a(gate448inter8), .b(gate448inter7), .O(gate448inter9));
  nand2 gate2419(.a(s_267), .b(gate448inter3), .O(gate448inter10));
  nor2  gate2420(.a(gate448inter10), .b(gate448inter9), .O(gate448inter11));
  nor2  gate2421(.a(gate448inter11), .b(gate448inter6), .O(gate448inter12));
  nand2 gate2422(.a(gate448inter12), .b(gate448inter1), .O(G1257));

  xor2  gate1051(.a(G1177), .b(G16), .O(gate449inter0));
  nand2 gate1052(.a(gate449inter0), .b(s_72), .O(gate449inter1));
  and2  gate1053(.a(G1177), .b(G16), .O(gate449inter2));
  inv1  gate1054(.a(s_72), .O(gate449inter3));
  inv1  gate1055(.a(s_73), .O(gate449inter4));
  nand2 gate1056(.a(gate449inter4), .b(gate449inter3), .O(gate449inter5));
  nor2  gate1057(.a(gate449inter5), .b(gate449inter2), .O(gate449inter6));
  inv1  gate1058(.a(G16), .O(gate449inter7));
  inv1  gate1059(.a(G1177), .O(gate449inter8));
  nand2 gate1060(.a(gate449inter8), .b(gate449inter7), .O(gate449inter9));
  nand2 gate1061(.a(s_73), .b(gate449inter3), .O(gate449inter10));
  nor2  gate1062(.a(gate449inter10), .b(gate449inter9), .O(gate449inter11));
  nor2  gate1063(.a(gate449inter11), .b(gate449inter6), .O(gate449inter12));
  nand2 gate1064(.a(gate449inter12), .b(gate449inter1), .O(G1258));
nand2 gate450( .a(G1081), .b(G1177), .O(G1259) );
nand2 gate451( .a(G17), .b(G1180), .O(G1260) );

  xor2  gate1317(.a(G1180), .b(G1084), .O(gate452inter0));
  nand2 gate1318(.a(gate452inter0), .b(s_110), .O(gate452inter1));
  and2  gate1319(.a(G1180), .b(G1084), .O(gate452inter2));
  inv1  gate1320(.a(s_110), .O(gate452inter3));
  inv1  gate1321(.a(s_111), .O(gate452inter4));
  nand2 gate1322(.a(gate452inter4), .b(gate452inter3), .O(gate452inter5));
  nor2  gate1323(.a(gate452inter5), .b(gate452inter2), .O(gate452inter6));
  inv1  gate1324(.a(G1084), .O(gate452inter7));
  inv1  gate1325(.a(G1180), .O(gate452inter8));
  nand2 gate1326(.a(gate452inter8), .b(gate452inter7), .O(gate452inter9));
  nand2 gate1327(.a(s_111), .b(gate452inter3), .O(gate452inter10));
  nor2  gate1328(.a(gate452inter10), .b(gate452inter9), .O(gate452inter11));
  nor2  gate1329(.a(gate452inter11), .b(gate452inter6), .O(gate452inter12));
  nand2 gate1330(.a(gate452inter12), .b(gate452inter1), .O(G1261));
nand2 gate453( .a(G18), .b(G1183), .O(G1262) );
nand2 gate454( .a(G1087), .b(G1183), .O(G1263) );

  xor2  gate1079(.a(G1186), .b(G19), .O(gate455inter0));
  nand2 gate1080(.a(gate455inter0), .b(s_76), .O(gate455inter1));
  and2  gate1081(.a(G1186), .b(G19), .O(gate455inter2));
  inv1  gate1082(.a(s_76), .O(gate455inter3));
  inv1  gate1083(.a(s_77), .O(gate455inter4));
  nand2 gate1084(.a(gate455inter4), .b(gate455inter3), .O(gate455inter5));
  nor2  gate1085(.a(gate455inter5), .b(gate455inter2), .O(gate455inter6));
  inv1  gate1086(.a(G19), .O(gate455inter7));
  inv1  gate1087(.a(G1186), .O(gate455inter8));
  nand2 gate1088(.a(gate455inter8), .b(gate455inter7), .O(gate455inter9));
  nand2 gate1089(.a(s_77), .b(gate455inter3), .O(gate455inter10));
  nor2  gate1090(.a(gate455inter10), .b(gate455inter9), .O(gate455inter11));
  nor2  gate1091(.a(gate455inter11), .b(gate455inter6), .O(gate455inter12));
  nand2 gate1092(.a(gate455inter12), .b(gate455inter1), .O(G1264));
nand2 gate456( .a(G1090), .b(G1186), .O(G1265) );
nand2 gate457( .a(G20), .b(G1189), .O(G1266) );
nand2 gate458( .a(G1093), .b(G1189), .O(G1267) );
nand2 gate459( .a(G21), .b(G1192), .O(G1268) );
nand2 gate460( .a(G1096), .b(G1192), .O(G1269) );
nand2 gate461( .a(G22), .b(G1195), .O(G1270) );
nand2 gate462( .a(G1099), .b(G1195), .O(G1271) );

  xor2  gate1261(.a(G1198), .b(G23), .O(gate463inter0));
  nand2 gate1262(.a(gate463inter0), .b(s_102), .O(gate463inter1));
  and2  gate1263(.a(G1198), .b(G23), .O(gate463inter2));
  inv1  gate1264(.a(s_102), .O(gate463inter3));
  inv1  gate1265(.a(s_103), .O(gate463inter4));
  nand2 gate1266(.a(gate463inter4), .b(gate463inter3), .O(gate463inter5));
  nor2  gate1267(.a(gate463inter5), .b(gate463inter2), .O(gate463inter6));
  inv1  gate1268(.a(G23), .O(gate463inter7));
  inv1  gate1269(.a(G1198), .O(gate463inter8));
  nand2 gate1270(.a(gate463inter8), .b(gate463inter7), .O(gate463inter9));
  nand2 gate1271(.a(s_103), .b(gate463inter3), .O(gate463inter10));
  nor2  gate1272(.a(gate463inter10), .b(gate463inter9), .O(gate463inter11));
  nor2  gate1273(.a(gate463inter11), .b(gate463inter6), .O(gate463inter12));
  nand2 gate1274(.a(gate463inter12), .b(gate463inter1), .O(G1272));
nand2 gate464( .a(G1102), .b(G1198), .O(G1273) );
nand2 gate465( .a(G24), .b(G1201), .O(G1274) );
nand2 gate466( .a(G1105), .b(G1201), .O(G1275) );
nand2 gate467( .a(G25), .b(G1204), .O(G1276) );
nand2 gate468( .a(G1108), .b(G1204), .O(G1277) );
nand2 gate469( .a(G26), .b(G1207), .O(G1278) );
nand2 gate470( .a(G1111), .b(G1207), .O(G1279) );
nand2 gate471( .a(G27), .b(G1210), .O(G1280) );
nand2 gate472( .a(G1114), .b(G1210), .O(G1281) );

  xor2  gate2059(.a(G1213), .b(G28), .O(gate473inter0));
  nand2 gate2060(.a(gate473inter0), .b(s_216), .O(gate473inter1));
  and2  gate2061(.a(G1213), .b(G28), .O(gate473inter2));
  inv1  gate2062(.a(s_216), .O(gate473inter3));
  inv1  gate2063(.a(s_217), .O(gate473inter4));
  nand2 gate2064(.a(gate473inter4), .b(gate473inter3), .O(gate473inter5));
  nor2  gate2065(.a(gate473inter5), .b(gate473inter2), .O(gate473inter6));
  inv1  gate2066(.a(G28), .O(gate473inter7));
  inv1  gate2067(.a(G1213), .O(gate473inter8));
  nand2 gate2068(.a(gate473inter8), .b(gate473inter7), .O(gate473inter9));
  nand2 gate2069(.a(s_217), .b(gate473inter3), .O(gate473inter10));
  nor2  gate2070(.a(gate473inter10), .b(gate473inter9), .O(gate473inter11));
  nor2  gate2071(.a(gate473inter11), .b(gate473inter6), .O(gate473inter12));
  nand2 gate2072(.a(gate473inter12), .b(gate473inter1), .O(G1282));

  xor2  gate1779(.a(G1213), .b(G1117), .O(gate474inter0));
  nand2 gate1780(.a(gate474inter0), .b(s_176), .O(gate474inter1));
  and2  gate1781(.a(G1213), .b(G1117), .O(gate474inter2));
  inv1  gate1782(.a(s_176), .O(gate474inter3));
  inv1  gate1783(.a(s_177), .O(gate474inter4));
  nand2 gate1784(.a(gate474inter4), .b(gate474inter3), .O(gate474inter5));
  nor2  gate1785(.a(gate474inter5), .b(gate474inter2), .O(gate474inter6));
  inv1  gate1786(.a(G1117), .O(gate474inter7));
  inv1  gate1787(.a(G1213), .O(gate474inter8));
  nand2 gate1788(.a(gate474inter8), .b(gate474inter7), .O(gate474inter9));
  nand2 gate1789(.a(s_177), .b(gate474inter3), .O(gate474inter10));
  nor2  gate1790(.a(gate474inter10), .b(gate474inter9), .O(gate474inter11));
  nor2  gate1791(.a(gate474inter11), .b(gate474inter6), .O(gate474inter12));
  nand2 gate1792(.a(gate474inter12), .b(gate474inter1), .O(G1283));

  xor2  gate2367(.a(G1216), .b(G29), .O(gate475inter0));
  nand2 gate2368(.a(gate475inter0), .b(s_260), .O(gate475inter1));
  and2  gate2369(.a(G1216), .b(G29), .O(gate475inter2));
  inv1  gate2370(.a(s_260), .O(gate475inter3));
  inv1  gate2371(.a(s_261), .O(gate475inter4));
  nand2 gate2372(.a(gate475inter4), .b(gate475inter3), .O(gate475inter5));
  nor2  gate2373(.a(gate475inter5), .b(gate475inter2), .O(gate475inter6));
  inv1  gate2374(.a(G29), .O(gate475inter7));
  inv1  gate2375(.a(G1216), .O(gate475inter8));
  nand2 gate2376(.a(gate475inter8), .b(gate475inter7), .O(gate475inter9));
  nand2 gate2377(.a(s_261), .b(gate475inter3), .O(gate475inter10));
  nor2  gate2378(.a(gate475inter10), .b(gate475inter9), .O(gate475inter11));
  nor2  gate2379(.a(gate475inter11), .b(gate475inter6), .O(gate475inter12));
  nand2 gate2380(.a(gate475inter12), .b(gate475inter1), .O(G1284));
nand2 gate476( .a(G1120), .b(G1216), .O(G1285) );
nand2 gate477( .a(G30), .b(G1219), .O(G1286) );
nand2 gate478( .a(G1123), .b(G1219), .O(G1287) );

  xor2  gate2521(.a(G1222), .b(G31), .O(gate479inter0));
  nand2 gate2522(.a(gate479inter0), .b(s_282), .O(gate479inter1));
  and2  gate2523(.a(G1222), .b(G31), .O(gate479inter2));
  inv1  gate2524(.a(s_282), .O(gate479inter3));
  inv1  gate2525(.a(s_283), .O(gate479inter4));
  nand2 gate2526(.a(gate479inter4), .b(gate479inter3), .O(gate479inter5));
  nor2  gate2527(.a(gate479inter5), .b(gate479inter2), .O(gate479inter6));
  inv1  gate2528(.a(G31), .O(gate479inter7));
  inv1  gate2529(.a(G1222), .O(gate479inter8));
  nand2 gate2530(.a(gate479inter8), .b(gate479inter7), .O(gate479inter9));
  nand2 gate2531(.a(s_283), .b(gate479inter3), .O(gate479inter10));
  nor2  gate2532(.a(gate479inter10), .b(gate479inter9), .O(gate479inter11));
  nor2  gate2533(.a(gate479inter11), .b(gate479inter6), .O(gate479inter12));
  nand2 gate2534(.a(gate479inter12), .b(gate479inter1), .O(G1288));
nand2 gate480( .a(G1126), .b(G1222), .O(G1289) );
nand2 gate481( .a(G32), .b(G1225), .O(G1290) );

  xor2  gate2143(.a(G1225), .b(G1129), .O(gate482inter0));
  nand2 gate2144(.a(gate482inter0), .b(s_228), .O(gate482inter1));
  and2  gate2145(.a(G1225), .b(G1129), .O(gate482inter2));
  inv1  gate2146(.a(s_228), .O(gate482inter3));
  inv1  gate2147(.a(s_229), .O(gate482inter4));
  nand2 gate2148(.a(gate482inter4), .b(gate482inter3), .O(gate482inter5));
  nor2  gate2149(.a(gate482inter5), .b(gate482inter2), .O(gate482inter6));
  inv1  gate2150(.a(G1129), .O(gate482inter7));
  inv1  gate2151(.a(G1225), .O(gate482inter8));
  nand2 gate2152(.a(gate482inter8), .b(gate482inter7), .O(gate482inter9));
  nand2 gate2153(.a(s_229), .b(gate482inter3), .O(gate482inter10));
  nor2  gate2154(.a(gate482inter10), .b(gate482inter9), .O(gate482inter11));
  nor2  gate2155(.a(gate482inter11), .b(gate482inter6), .O(gate482inter12));
  nand2 gate2156(.a(gate482inter12), .b(gate482inter1), .O(G1291));
nand2 gate483( .a(G1228), .b(G1229), .O(G1292) );
nand2 gate484( .a(G1230), .b(G1231), .O(G1293) );
nand2 gate485( .a(G1232), .b(G1233), .O(G1294) );
nand2 gate486( .a(G1234), .b(G1235), .O(G1295) );
nand2 gate487( .a(G1236), .b(G1237), .O(G1296) );
nand2 gate488( .a(G1238), .b(G1239), .O(G1297) );
nand2 gate489( .a(G1240), .b(G1241), .O(G1298) );
nand2 gate490( .a(G1242), .b(G1243), .O(G1299) );

  xor2  gate701(.a(G1245), .b(G1244), .O(gate491inter0));
  nand2 gate702(.a(gate491inter0), .b(s_22), .O(gate491inter1));
  and2  gate703(.a(G1245), .b(G1244), .O(gate491inter2));
  inv1  gate704(.a(s_22), .O(gate491inter3));
  inv1  gate705(.a(s_23), .O(gate491inter4));
  nand2 gate706(.a(gate491inter4), .b(gate491inter3), .O(gate491inter5));
  nor2  gate707(.a(gate491inter5), .b(gate491inter2), .O(gate491inter6));
  inv1  gate708(.a(G1244), .O(gate491inter7));
  inv1  gate709(.a(G1245), .O(gate491inter8));
  nand2 gate710(.a(gate491inter8), .b(gate491inter7), .O(gate491inter9));
  nand2 gate711(.a(s_23), .b(gate491inter3), .O(gate491inter10));
  nor2  gate712(.a(gate491inter10), .b(gate491inter9), .O(gate491inter11));
  nor2  gate713(.a(gate491inter11), .b(gate491inter6), .O(gate491inter12));
  nand2 gate714(.a(gate491inter12), .b(gate491inter1), .O(G1300));
nand2 gate492( .a(G1246), .b(G1247), .O(G1301) );

  xor2  gate827(.a(G1249), .b(G1248), .O(gate493inter0));
  nand2 gate828(.a(gate493inter0), .b(s_40), .O(gate493inter1));
  and2  gate829(.a(G1249), .b(G1248), .O(gate493inter2));
  inv1  gate830(.a(s_40), .O(gate493inter3));
  inv1  gate831(.a(s_41), .O(gate493inter4));
  nand2 gate832(.a(gate493inter4), .b(gate493inter3), .O(gate493inter5));
  nor2  gate833(.a(gate493inter5), .b(gate493inter2), .O(gate493inter6));
  inv1  gate834(.a(G1248), .O(gate493inter7));
  inv1  gate835(.a(G1249), .O(gate493inter8));
  nand2 gate836(.a(gate493inter8), .b(gate493inter7), .O(gate493inter9));
  nand2 gate837(.a(s_41), .b(gate493inter3), .O(gate493inter10));
  nor2  gate838(.a(gate493inter10), .b(gate493inter9), .O(gate493inter11));
  nor2  gate839(.a(gate493inter11), .b(gate493inter6), .O(gate493inter12));
  nand2 gate840(.a(gate493inter12), .b(gate493inter1), .O(G1302));

  xor2  gate1849(.a(G1251), .b(G1250), .O(gate494inter0));
  nand2 gate1850(.a(gate494inter0), .b(s_186), .O(gate494inter1));
  and2  gate1851(.a(G1251), .b(G1250), .O(gate494inter2));
  inv1  gate1852(.a(s_186), .O(gate494inter3));
  inv1  gate1853(.a(s_187), .O(gate494inter4));
  nand2 gate1854(.a(gate494inter4), .b(gate494inter3), .O(gate494inter5));
  nor2  gate1855(.a(gate494inter5), .b(gate494inter2), .O(gate494inter6));
  inv1  gate1856(.a(G1250), .O(gate494inter7));
  inv1  gate1857(.a(G1251), .O(gate494inter8));
  nand2 gate1858(.a(gate494inter8), .b(gate494inter7), .O(gate494inter9));
  nand2 gate1859(.a(s_187), .b(gate494inter3), .O(gate494inter10));
  nor2  gate1860(.a(gate494inter10), .b(gate494inter9), .O(gate494inter11));
  nor2  gate1861(.a(gate494inter11), .b(gate494inter6), .O(gate494inter12));
  nand2 gate1862(.a(gate494inter12), .b(gate494inter1), .O(G1303));
nand2 gate495( .a(G1252), .b(G1253), .O(G1304) );

  xor2  gate1709(.a(G1255), .b(G1254), .O(gate496inter0));
  nand2 gate1710(.a(gate496inter0), .b(s_166), .O(gate496inter1));
  and2  gate1711(.a(G1255), .b(G1254), .O(gate496inter2));
  inv1  gate1712(.a(s_166), .O(gate496inter3));
  inv1  gate1713(.a(s_167), .O(gate496inter4));
  nand2 gate1714(.a(gate496inter4), .b(gate496inter3), .O(gate496inter5));
  nor2  gate1715(.a(gate496inter5), .b(gate496inter2), .O(gate496inter6));
  inv1  gate1716(.a(G1254), .O(gate496inter7));
  inv1  gate1717(.a(G1255), .O(gate496inter8));
  nand2 gate1718(.a(gate496inter8), .b(gate496inter7), .O(gate496inter9));
  nand2 gate1719(.a(s_167), .b(gate496inter3), .O(gate496inter10));
  nor2  gate1720(.a(gate496inter10), .b(gate496inter9), .O(gate496inter11));
  nor2  gate1721(.a(gate496inter11), .b(gate496inter6), .O(gate496inter12));
  nand2 gate1722(.a(gate496inter12), .b(gate496inter1), .O(G1305));
nand2 gate497( .a(G1256), .b(G1257), .O(G1306) );
nand2 gate498( .a(G1258), .b(G1259), .O(G1307) );
nand2 gate499( .a(G1260), .b(G1261), .O(G1308) );
nand2 gate500( .a(G1262), .b(G1263), .O(G1309) );

  xor2  gate1303(.a(G1265), .b(G1264), .O(gate501inter0));
  nand2 gate1304(.a(gate501inter0), .b(s_108), .O(gate501inter1));
  and2  gate1305(.a(G1265), .b(G1264), .O(gate501inter2));
  inv1  gate1306(.a(s_108), .O(gate501inter3));
  inv1  gate1307(.a(s_109), .O(gate501inter4));
  nand2 gate1308(.a(gate501inter4), .b(gate501inter3), .O(gate501inter5));
  nor2  gate1309(.a(gate501inter5), .b(gate501inter2), .O(gate501inter6));
  inv1  gate1310(.a(G1264), .O(gate501inter7));
  inv1  gate1311(.a(G1265), .O(gate501inter8));
  nand2 gate1312(.a(gate501inter8), .b(gate501inter7), .O(gate501inter9));
  nand2 gate1313(.a(s_109), .b(gate501inter3), .O(gate501inter10));
  nor2  gate1314(.a(gate501inter10), .b(gate501inter9), .O(gate501inter11));
  nor2  gate1315(.a(gate501inter11), .b(gate501inter6), .O(gate501inter12));
  nand2 gate1316(.a(gate501inter12), .b(gate501inter1), .O(G1310));
nand2 gate502( .a(G1266), .b(G1267), .O(G1311) );

  xor2  gate729(.a(G1269), .b(G1268), .O(gate503inter0));
  nand2 gate730(.a(gate503inter0), .b(s_26), .O(gate503inter1));
  and2  gate731(.a(G1269), .b(G1268), .O(gate503inter2));
  inv1  gate732(.a(s_26), .O(gate503inter3));
  inv1  gate733(.a(s_27), .O(gate503inter4));
  nand2 gate734(.a(gate503inter4), .b(gate503inter3), .O(gate503inter5));
  nor2  gate735(.a(gate503inter5), .b(gate503inter2), .O(gate503inter6));
  inv1  gate736(.a(G1268), .O(gate503inter7));
  inv1  gate737(.a(G1269), .O(gate503inter8));
  nand2 gate738(.a(gate503inter8), .b(gate503inter7), .O(gate503inter9));
  nand2 gate739(.a(s_27), .b(gate503inter3), .O(gate503inter10));
  nor2  gate740(.a(gate503inter10), .b(gate503inter9), .O(gate503inter11));
  nor2  gate741(.a(gate503inter11), .b(gate503inter6), .O(gate503inter12));
  nand2 gate742(.a(gate503inter12), .b(gate503inter1), .O(G1312));

  xor2  gate2353(.a(G1271), .b(G1270), .O(gate504inter0));
  nand2 gate2354(.a(gate504inter0), .b(s_258), .O(gate504inter1));
  and2  gate2355(.a(G1271), .b(G1270), .O(gate504inter2));
  inv1  gate2356(.a(s_258), .O(gate504inter3));
  inv1  gate2357(.a(s_259), .O(gate504inter4));
  nand2 gate2358(.a(gate504inter4), .b(gate504inter3), .O(gate504inter5));
  nor2  gate2359(.a(gate504inter5), .b(gate504inter2), .O(gate504inter6));
  inv1  gate2360(.a(G1270), .O(gate504inter7));
  inv1  gate2361(.a(G1271), .O(gate504inter8));
  nand2 gate2362(.a(gate504inter8), .b(gate504inter7), .O(gate504inter9));
  nand2 gate2363(.a(s_259), .b(gate504inter3), .O(gate504inter10));
  nor2  gate2364(.a(gate504inter10), .b(gate504inter9), .O(gate504inter11));
  nor2  gate2365(.a(gate504inter11), .b(gate504inter6), .O(gate504inter12));
  nand2 gate2366(.a(gate504inter12), .b(gate504inter1), .O(G1313));
nand2 gate505( .a(G1272), .b(G1273), .O(G1314) );
nand2 gate506( .a(G1274), .b(G1275), .O(G1315) );

  xor2  gate1219(.a(G1277), .b(G1276), .O(gate507inter0));
  nand2 gate1220(.a(gate507inter0), .b(s_96), .O(gate507inter1));
  and2  gate1221(.a(G1277), .b(G1276), .O(gate507inter2));
  inv1  gate1222(.a(s_96), .O(gate507inter3));
  inv1  gate1223(.a(s_97), .O(gate507inter4));
  nand2 gate1224(.a(gate507inter4), .b(gate507inter3), .O(gate507inter5));
  nor2  gate1225(.a(gate507inter5), .b(gate507inter2), .O(gate507inter6));
  inv1  gate1226(.a(G1276), .O(gate507inter7));
  inv1  gate1227(.a(G1277), .O(gate507inter8));
  nand2 gate1228(.a(gate507inter8), .b(gate507inter7), .O(gate507inter9));
  nand2 gate1229(.a(s_97), .b(gate507inter3), .O(gate507inter10));
  nor2  gate1230(.a(gate507inter10), .b(gate507inter9), .O(gate507inter11));
  nor2  gate1231(.a(gate507inter11), .b(gate507inter6), .O(gate507inter12));
  nand2 gate1232(.a(gate507inter12), .b(gate507inter1), .O(G1316));

  xor2  gate1485(.a(G1279), .b(G1278), .O(gate508inter0));
  nand2 gate1486(.a(gate508inter0), .b(s_134), .O(gate508inter1));
  and2  gate1487(.a(G1279), .b(G1278), .O(gate508inter2));
  inv1  gate1488(.a(s_134), .O(gate508inter3));
  inv1  gate1489(.a(s_135), .O(gate508inter4));
  nand2 gate1490(.a(gate508inter4), .b(gate508inter3), .O(gate508inter5));
  nor2  gate1491(.a(gate508inter5), .b(gate508inter2), .O(gate508inter6));
  inv1  gate1492(.a(G1278), .O(gate508inter7));
  inv1  gate1493(.a(G1279), .O(gate508inter8));
  nand2 gate1494(.a(gate508inter8), .b(gate508inter7), .O(gate508inter9));
  nand2 gate1495(.a(s_135), .b(gate508inter3), .O(gate508inter10));
  nor2  gate1496(.a(gate508inter10), .b(gate508inter9), .O(gate508inter11));
  nor2  gate1497(.a(gate508inter11), .b(gate508inter6), .O(gate508inter12));
  nand2 gate1498(.a(gate508inter12), .b(gate508inter1), .O(G1317));
nand2 gate509( .a(G1280), .b(G1281), .O(G1318) );

  xor2  gate2185(.a(G1283), .b(G1282), .O(gate510inter0));
  nand2 gate2186(.a(gate510inter0), .b(s_234), .O(gate510inter1));
  and2  gate2187(.a(G1283), .b(G1282), .O(gate510inter2));
  inv1  gate2188(.a(s_234), .O(gate510inter3));
  inv1  gate2189(.a(s_235), .O(gate510inter4));
  nand2 gate2190(.a(gate510inter4), .b(gate510inter3), .O(gate510inter5));
  nor2  gate2191(.a(gate510inter5), .b(gate510inter2), .O(gate510inter6));
  inv1  gate2192(.a(G1282), .O(gate510inter7));
  inv1  gate2193(.a(G1283), .O(gate510inter8));
  nand2 gate2194(.a(gate510inter8), .b(gate510inter7), .O(gate510inter9));
  nand2 gate2195(.a(s_235), .b(gate510inter3), .O(gate510inter10));
  nor2  gate2196(.a(gate510inter10), .b(gate510inter9), .O(gate510inter11));
  nor2  gate2197(.a(gate510inter11), .b(gate510inter6), .O(gate510inter12));
  nand2 gate2198(.a(gate510inter12), .b(gate510inter1), .O(G1319));

  xor2  gate2381(.a(G1285), .b(G1284), .O(gate511inter0));
  nand2 gate2382(.a(gate511inter0), .b(s_262), .O(gate511inter1));
  and2  gate2383(.a(G1285), .b(G1284), .O(gate511inter2));
  inv1  gate2384(.a(s_262), .O(gate511inter3));
  inv1  gate2385(.a(s_263), .O(gate511inter4));
  nand2 gate2386(.a(gate511inter4), .b(gate511inter3), .O(gate511inter5));
  nor2  gate2387(.a(gate511inter5), .b(gate511inter2), .O(gate511inter6));
  inv1  gate2388(.a(G1284), .O(gate511inter7));
  inv1  gate2389(.a(G1285), .O(gate511inter8));
  nand2 gate2390(.a(gate511inter8), .b(gate511inter7), .O(gate511inter9));
  nand2 gate2391(.a(s_263), .b(gate511inter3), .O(gate511inter10));
  nor2  gate2392(.a(gate511inter10), .b(gate511inter9), .O(gate511inter11));
  nor2  gate2393(.a(gate511inter11), .b(gate511inter6), .O(gate511inter12));
  nand2 gate2394(.a(gate511inter12), .b(gate511inter1), .O(G1320));
nand2 gate512( .a(G1286), .b(G1287), .O(G1321) );
nand2 gate513( .a(G1288), .b(G1289), .O(G1322) );

  xor2  gate1387(.a(G1291), .b(G1290), .O(gate514inter0));
  nand2 gate1388(.a(gate514inter0), .b(s_120), .O(gate514inter1));
  and2  gate1389(.a(G1291), .b(G1290), .O(gate514inter2));
  inv1  gate1390(.a(s_120), .O(gate514inter3));
  inv1  gate1391(.a(s_121), .O(gate514inter4));
  nand2 gate1392(.a(gate514inter4), .b(gate514inter3), .O(gate514inter5));
  nor2  gate1393(.a(gate514inter5), .b(gate514inter2), .O(gate514inter6));
  inv1  gate1394(.a(G1290), .O(gate514inter7));
  inv1  gate1395(.a(G1291), .O(gate514inter8));
  nand2 gate1396(.a(gate514inter8), .b(gate514inter7), .O(gate514inter9));
  nand2 gate1397(.a(s_121), .b(gate514inter3), .O(gate514inter10));
  nor2  gate1398(.a(gate514inter10), .b(gate514inter9), .O(gate514inter11));
  nor2  gate1399(.a(gate514inter11), .b(gate514inter6), .O(gate514inter12));
  nand2 gate1400(.a(gate514inter12), .b(gate514inter1), .O(G1323));
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule