module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);

input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;//RE__PI;

input s_0,s_1;//RE__ALLOW(00,01,10,11);
input s_2,s_3;//RE__ALLOW(00,01,10,11);
input s_4,s_5;//RE__ALLOW(00,01,10,11);
input s_6,s_7;//RE__ALLOW(00,01,10,11);
input s_8,s_9;//RE__ALLOW(00,01,10,11);
input s_10,s_11;//RE__ALLOW(00,01,10,11);
input s_12,s_13;//RE__ALLOW(00,01,10,11);
input s_14,s_15;//RE__ALLOW(00,01,10,11);
input s_16,s_17;//RE__ALLOW(00,01,10,11);
input s_18,s_19;//RE__ALLOW(00,01,10,11);
input s_20,s_21;//RE__ALLOW(00,01,10,11);
input s_22,s_23;//RE__ALLOW(00,01,10,11);
input s_24,s_25;//RE__ALLOW(00,01,10,11);
input s_26,s_27;//RE__ALLOW(00,01,10,11);
input s_28,s_29;//RE__ALLOW(00,01,10,11);
input s_30,s_31;//RE__ALLOW(00,01,10,11);
input s_32,s_33;//RE__ALLOW(00,01,10,11);
input s_34,s_35;//RE__ALLOW(00,01,10,11);
input s_36,s_37;//RE__ALLOW(00,01,10,11);
input s_38,s_39;//RE__ALLOW(00,01,10,11);
input s_40,s_41;//RE__ALLOW(00,01,10,11);
input s_42,s_43;//RE__ALLOW(00,01,10,11);
input s_44,s_45;//RE__ALLOW(00,01,10,11);
input s_46,s_47;//RE__ALLOW(00,01,10,11);
input s_48,s_49;//RE__ALLOW(00,01,10,11);
input s_50,s_51;//RE__ALLOW(00,01,10,11);
input s_52,s_53;//RE__ALLOW(00,01,10,11);
input s_54,s_55;//RE__ALLOW(00,01,10,11);
input s_56,s_57;//RE__ALLOW(00,01,10,11);
input s_58,s_59;//RE__ALLOW(00,01,10,11);
input s_60,s_61;//RE__ALLOW(00,01,10,11);
input s_62,s_63;//RE__ALLOW(00,01,10,11);
input s_64,s_65;//RE__ALLOW(00,01,10,11);
input s_66,s_67;//RE__ALLOW(00,01,10,11);
input s_68,s_69;//RE__ALLOW(00,01,10,11);
input s_70,s_71;//RE__ALLOW(00,01,10,11);
input s_72,s_73;//RE__ALLOW(00,01,10,11);
input s_74,s_75;//RE__ALLOW(00,01,10,11);
input s_76,s_77;//RE__ALLOW(00,01,10,11);
input s_78,s_79;//RE__ALLOW(00,01,10,11);
input s_80,s_81;//RE__ALLOW(00,01,10,11);
input s_82,s_83;//RE__ALLOW(00,01,10,11);
input s_84,s_85;//RE__ALLOW(00,01,10,11);
input s_86,s_87;//RE__ALLOW(00,01,10,11);
input s_88,s_89;//RE__ALLOW(00,01,10,11);
input s_90,s_91;//RE__ALLOW(00,01,10,11);
input s_92,s_93;//RE__ALLOW(00,01,10,11);
input s_94,s_95;//RE__ALLOW(00,01,10,11);
input s_96,s_97;//RE__ALLOW(00,01,10,11);
input s_98,s_99;//RE__ALLOW(00,01,10,11);
input s_100,s_101;//RE__ALLOW(00,01,10,11);
input s_102,s_103;//RE__ALLOW(00,01,10,11);
input s_104,s_105;//RE__ALLOW(00,01,10,11);
input s_106,s_107;//RE__ALLOW(00,01,10,11);
input s_108,s_109;//RE__ALLOW(00,01,10,11);
input s_110,s_111;//RE__ALLOW(00,01,10,11);
input s_112,s_113;//RE__ALLOW(00,01,10,11);
input s_114,s_115;//RE__ALLOW(00,01,10,11);
input s_116,s_117;//RE__ALLOW(00,01,10,11);
input s_118,s_119;//RE__ALLOW(00,01,10,11);
input s_120,s_121;//RE__ALLOW(00,01,10,11);
input s_122,s_123;//RE__ALLOW(00,01,10,11);
input s_124,s_125;//RE__ALLOW(00,01,10,11);
input s_126,s_127;//RE__ALLOW(00,01,10,11);
input s_128,s_129;//RE__ALLOW(00,01,10,11);
input s_130,s_131;//RE__ALLOW(00,01,10,11);
input s_132,s_133;//RE__ALLOW(00,01,10,11);
input s_134,s_135;//RE__ALLOW(00,01,10,11);
input s_136,s_137;//RE__ALLOW(00,01,10,11);
input s_138,s_139;//RE__ALLOW(00,01,10,11);
input s_140,s_141;//RE__ALLOW(00,01,10,11);
input s_142,s_143;//RE__ALLOW(00,01,10,11);
input s_144,s_145;//RE__ALLOW(00,01,10,11);
input s_146,s_147;//RE__ALLOW(00,01,10,11);
input s_148,s_149;//RE__ALLOW(00,01,10,11);
input s_150,s_151;//RE__ALLOW(00,01,10,11);
input s_152,s_153;//RE__ALLOW(00,01,10,11);
input s_154,s_155;//RE__ALLOW(00,01,10,11);
input s_156,s_157;//RE__ALLOW(00,01,10,11);
input s_158,s_159;//RE__ALLOW(00,01,10,11);
input s_160,s_161;//RE__ALLOW(00,01,10,11);
input s_162,s_163;//RE__ALLOW(00,01,10,11);
input s_164,s_165;//RE__ALLOW(00,01,10,11);
input s_166,s_167;//RE__ALLOW(00,01,10,11);
input s_168,s_169;//RE__ALLOW(00,01,10,11);
input s_170,s_171;//RE__ALLOW(00,01,10,11);
input s_172,s_173;//RE__ALLOW(00,01,10,11);
input s_174,s_175;//RE__ALLOW(00,01,10,11);
input s_176,s_177;//RE__ALLOW(00,01,10,11);
input s_178,s_179;//RE__ALLOW(00,01,10,11);
input s_180,s_181;//RE__ALLOW(00,01,10,11);
input s_182,s_183;//RE__ALLOW(00,01,10,11);
input s_184,s_185;//RE__ALLOW(00,01,10,11);
input s_186,s_187;//RE__ALLOW(00,01,10,11);
input s_188,s_189;//RE__ALLOW(00,01,10,11);
input s_190,s_191;//RE__ALLOW(00,01,10,11);
input s_192,s_193;//RE__ALLOW(00,01,10,11);
input s_194,s_195;//RE__ALLOW(00,01,10,11);
input s_196,s_197;//RE__ALLOW(00,01,10,11);
input s_198,s_199;//RE__ALLOW(00,01,10,11);
input s_200,s_201;//RE__ALLOW(00,01,10,11);
input s_202,s_203;//RE__ALLOW(00,01,10,11);
input s_204,s_205;//RE__ALLOW(00,01,10,11);
input s_206,s_207;//RE__ALLOW(00,01,10,11);
input s_208,s_209;//RE__ALLOW(00,01,10,11);
input s_210,s_211;//RE__ALLOW(00,01,10,11);
input s_212,s_213;//RE__ALLOW(00,01,10,11);
input s_214,s_215;//RE__ALLOW(00,01,10,11);
input s_216,s_217;//RE__ALLOW(00,01,10,11);
input s_218,s_219;//RE__ALLOW(00,01,10,11);
input s_220,s_221;//RE__ALLOW(00,01,10,11);
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;

  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate108inter0, gate108inter1, gate108inter2, gate108inter3, gate108inter4, gate108inter5, gate108inter6, gate108inter7, gate108inter8, gate108inter9, gate108inter10, gate108inter11, gate108inter12, gate92inter0, gate92inter1, gate92inter2, gate92inter3, gate92inter4, gate92inter5, gate92inter6, gate92inter7, gate92inter8, gate92inter9, gate92inter10, gate92inter11, gate92inter12, gate392inter0, gate392inter1, gate392inter2, gate392inter3, gate392inter4, gate392inter5, gate392inter6, gate392inter7, gate392inter8, gate392inter9, gate392inter10, gate392inter11, gate392inter12, gate120inter0, gate120inter1, gate120inter2, gate120inter3, gate120inter4, gate120inter5, gate120inter6, gate120inter7, gate120inter8, gate120inter9, gate120inter10, gate120inter11, gate120inter12, gate205inter0, gate205inter1, gate205inter2, gate205inter3, gate205inter4, gate205inter5, gate205inter6, gate205inter7, gate205inter8, gate205inter9, gate205inter10, gate205inter11, gate205inter12, gate186inter0, gate186inter1, gate186inter2, gate186inter3, gate186inter4, gate186inter5, gate186inter6, gate186inter7, gate186inter8, gate186inter9, gate186inter10, gate186inter11, gate186inter12, gate159inter0, gate159inter1, gate159inter2, gate159inter3, gate159inter4, gate159inter5, gate159inter6, gate159inter7, gate159inter8, gate159inter9, gate159inter10, gate159inter11, gate159inter12, gate281inter0, gate281inter1, gate281inter2, gate281inter3, gate281inter4, gate281inter5, gate281inter6, gate281inter7, gate281inter8, gate281inter9, gate281inter10, gate281inter11, gate281inter12, gate241inter0, gate241inter1, gate241inter2, gate241inter3, gate241inter4, gate241inter5, gate241inter6, gate241inter7, gate241inter8, gate241inter9, gate241inter10, gate241inter11, gate241inter12, gate426inter0, gate426inter1, gate426inter2, gate426inter3, gate426inter4, gate426inter5, gate426inter6, gate426inter7, gate426inter8, gate426inter9, gate426inter10, gate426inter11, gate426inter12, gate240inter0, gate240inter1, gate240inter2, gate240inter3, gate240inter4, gate240inter5, gate240inter6, gate240inter7, gate240inter8, gate240inter9, gate240inter10, gate240inter11, gate240inter12, gate264inter0, gate264inter1, gate264inter2, gate264inter3, gate264inter4, gate264inter5, gate264inter6, gate264inter7, gate264inter8, gate264inter9, gate264inter10, gate264inter11, gate264inter12, gate15inter0, gate15inter1, gate15inter2, gate15inter3, gate15inter4, gate15inter5, gate15inter6, gate15inter7, gate15inter8, gate15inter9, gate15inter10, gate15inter11, gate15inter12, gate164inter0, gate164inter1, gate164inter2, gate164inter3, gate164inter4, gate164inter5, gate164inter6, gate164inter7, gate164inter8, gate164inter9, gate164inter10, gate164inter11, gate164inter12, gate116inter0, gate116inter1, gate116inter2, gate116inter3, gate116inter4, gate116inter5, gate116inter6, gate116inter7, gate116inter8, gate116inter9, gate116inter10, gate116inter11, gate116inter12, gate230inter0, gate230inter1, gate230inter2, gate230inter3, gate230inter4, gate230inter5, gate230inter6, gate230inter7, gate230inter8, gate230inter9, gate230inter10, gate230inter11, gate230inter12, gate105inter0, gate105inter1, gate105inter2, gate105inter3, gate105inter4, gate105inter5, gate105inter6, gate105inter7, gate105inter8, gate105inter9, gate105inter10, gate105inter11, gate105inter12, gate282inter0, gate282inter1, gate282inter2, gate282inter3, gate282inter4, gate282inter5, gate282inter6, gate282inter7, gate282inter8, gate282inter9, gate282inter10, gate282inter11, gate282inter12, gate278inter0, gate278inter1, gate278inter2, gate278inter3, gate278inter4, gate278inter5, gate278inter6, gate278inter7, gate278inter8, gate278inter9, gate278inter10, gate278inter11, gate278inter12, gate142inter0, gate142inter1, gate142inter2, gate142inter3, gate142inter4, gate142inter5, gate142inter6, gate142inter7, gate142inter8, gate142inter9, gate142inter10, gate142inter11, gate142inter12, gate68inter0, gate68inter1, gate68inter2, gate68inter3, gate68inter4, gate68inter5, gate68inter6, gate68inter7, gate68inter8, gate68inter9, gate68inter10, gate68inter11, gate68inter12, gate63inter0, gate63inter1, gate63inter2, gate63inter3, gate63inter4, gate63inter5, gate63inter6, gate63inter7, gate63inter8, gate63inter9, gate63inter10, gate63inter11, gate63inter12, gate60inter0, gate60inter1, gate60inter2, gate60inter3, gate60inter4, gate60inter5, gate60inter6, gate60inter7, gate60inter8, gate60inter9, gate60inter10, gate60inter11, gate60inter12, gate132inter0, gate132inter1, gate132inter2, gate132inter3, gate132inter4, gate132inter5, gate132inter6, gate132inter7, gate132inter8, gate132inter9, gate132inter10, gate132inter11, gate132inter12, gate144inter0, gate144inter1, gate144inter2, gate144inter3, gate144inter4, gate144inter5, gate144inter6, gate144inter7, gate144inter8, gate144inter9, gate144inter10, gate144inter11, gate144inter12, gate466inter0, gate466inter1, gate466inter2, gate466inter3, gate466inter4, gate466inter5, gate466inter6, gate466inter7, gate466inter8, gate466inter9, gate466inter10, gate466inter11, gate466inter12, gate209inter0, gate209inter1, gate209inter2, gate209inter3, gate209inter4, gate209inter5, gate209inter6, gate209inter7, gate209inter8, gate209inter9, gate209inter10, gate209inter11, gate209inter12, gate11inter0, gate11inter1, gate11inter2, gate11inter3, gate11inter4, gate11inter5, gate11inter6, gate11inter7, gate11inter8, gate11inter9, gate11inter10, gate11inter11, gate11inter12, gate415inter0, gate415inter1, gate415inter2, gate415inter3, gate415inter4, gate415inter5, gate415inter6, gate415inter7, gate415inter8, gate415inter9, gate415inter10, gate415inter11, gate415inter12, gate412inter0, gate412inter1, gate412inter2, gate412inter3, gate412inter4, gate412inter5, gate412inter6, gate412inter7, gate412inter8, gate412inter9, gate412inter10, gate412inter11, gate412inter12, gate150inter0, gate150inter1, gate150inter2, gate150inter3, gate150inter4, gate150inter5, gate150inter6, gate150inter7, gate150inter8, gate150inter9, gate150inter10, gate150inter11, gate150inter12, gate160inter0, gate160inter1, gate160inter2, gate160inter3, gate160inter4, gate160inter5, gate160inter6, gate160inter7, gate160inter8, gate160inter9, gate160inter10, gate160inter11, gate160inter12, gate410inter0, gate410inter1, gate410inter2, gate410inter3, gate410inter4, gate410inter5, gate410inter6, gate410inter7, gate410inter8, gate410inter9, gate410inter10, gate410inter11, gate410inter12, gate212inter0, gate212inter1, gate212inter2, gate212inter3, gate212inter4, gate212inter5, gate212inter6, gate212inter7, gate212inter8, gate212inter9, gate212inter10, gate212inter11, gate212inter12, gate448inter0, gate448inter1, gate448inter2, gate448inter3, gate448inter4, gate448inter5, gate448inter6, gate448inter7, gate448inter8, gate448inter9, gate448inter10, gate448inter11, gate448inter12, gate156inter0, gate156inter1, gate156inter2, gate156inter3, gate156inter4, gate156inter5, gate156inter6, gate156inter7, gate156inter8, gate156inter9, gate156inter10, gate156inter11, gate156inter12, gate486inter0, gate486inter1, gate486inter2, gate486inter3, gate486inter4, gate486inter5, gate486inter6, gate486inter7, gate486inter8, gate486inter9, gate486inter10, gate486inter11, gate486inter12, gate404inter0, gate404inter1, gate404inter2, gate404inter3, gate404inter4, gate404inter5, gate404inter6, gate404inter7, gate404inter8, gate404inter9, gate404inter10, gate404inter11, gate404inter12, gate503inter0, gate503inter1, gate503inter2, gate503inter3, gate503inter4, gate503inter5, gate503inter6, gate503inter7, gate503inter8, gate503inter9, gate503inter10, gate503inter11, gate503inter12, gate265inter0, gate265inter1, gate265inter2, gate265inter3, gate265inter4, gate265inter5, gate265inter6, gate265inter7, gate265inter8, gate265inter9, gate265inter10, gate265inter11, gate265inter12, gate23inter0, gate23inter1, gate23inter2, gate23inter3, gate23inter4, gate23inter5, gate23inter6, gate23inter7, gate23inter8, gate23inter9, gate23inter10, gate23inter11, gate23inter12, gate501inter0, gate501inter1, gate501inter2, gate501inter3, gate501inter4, gate501inter5, gate501inter6, gate501inter7, gate501inter8, gate501inter9, gate501inter10, gate501inter11, gate501inter12, gate239inter0, gate239inter1, gate239inter2, gate239inter3, gate239inter4, gate239inter5, gate239inter6, gate239inter7, gate239inter8, gate239inter9, gate239inter10, gate239inter11, gate239inter12, gate45inter0, gate45inter1, gate45inter2, gate45inter3, gate45inter4, gate45inter5, gate45inter6, gate45inter7, gate45inter8, gate45inter9, gate45inter10, gate45inter11, gate45inter12, gate260inter0, gate260inter1, gate260inter2, gate260inter3, gate260inter4, gate260inter5, gate260inter6, gate260inter7, gate260inter8, gate260inter9, gate260inter10, gate260inter11, gate260inter12, gate31inter0, gate31inter1, gate31inter2, gate31inter3, gate31inter4, gate31inter5, gate31inter6, gate31inter7, gate31inter8, gate31inter9, gate31inter10, gate31inter11, gate31inter12, gate56inter0, gate56inter1, gate56inter2, gate56inter3, gate56inter4, gate56inter5, gate56inter6, gate56inter7, gate56inter8, gate56inter9, gate56inter10, gate56inter11, gate56inter12, gate158inter0, gate158inter1, gate158inter2, gate158inter3, gate158inter4, gate158inter5, gate158inter6, gate158inter7, gate158inter8, gate158inter9, gate158inter10, gate158inter11, gate158inter12, gate89inter0, gate89inter1, gate89inter2, gate89inter3, gate89inter4, gate89inter5, gate89inter6, gate89inter7, gate89inter8, gate89inter9, gate89inter10, gate89inter11, gate89inter12, gate179inter0, gate179inter1, gate179inter2, gate179inter3, gate179inter4, gate179inter5, gate179inter6, gate179inter7, gate179inter8, gate179inter9, gate179inter10, gate179inter11, gate179inter12, gate225inter0, gate225inter1, gate225inter2, gate225inter3, gate225inter4, gate225inter5, gate225inter6, gate225inter7, gate225inter8, gate225inter9, gate225inter10, gate225inter11, gate225inter12, gate409inter0, gate409inter1, gate409inter2, gate409inter3, gate409inter4, gate409inter5, gate409inter6, gate409inter7, gate409inter8, gate409inter9, gate409inter10, gate409inter11, gate409inter12, gate295inter0, gate295inter1, gate295inter2, gate295inter3, gate295inter4, gate295inter5, gate295inter6, gate295inter7, gate295inter8, gate295inter9, gate295inter10, gate295inter11, gate295inter12, gate485inter0, gate485inter1, gate485inter2, gate485inter3, gate485inter4, gate485inter5, gate485inter6, gate485inter7, gate485inter8, gate485inter9, gate485inter10, gate485inter11, gate485inter12, gate287inter0, gate287inter1, gate287inter2, gate287inter3, gate287inter4, gate287inter5, gate287inter6, gate287inter7, gate287inter8, gate287inter9, gate287inter10, gate287inter11, gate287inter12, gate217inter0, gate217inter1, gate217inter2, gate217inter3, gate217inter4, gate217inter5, gate217inter6, gate217inter7, gate217inter8, gate217inter9, gate217inter10, gate217inter11, gate217inter12, gate454inter0, gate454inter1, gate454inter2, gate454inter3, gate454inter4, gate454inter5, gate454inter6, gate454inter7, gate454inter8, gate454inter9, gate454inter10, gate454inter11, gate454inter12, gate274inter0, gate274inter1, gate274inter2, gate274inter3, gate274inter4, gate274inter5, gate274inter6, gate274inter7, gate274inter8, gate274inter9, gate274inter10, gate274inter11, gate274inter12, gate268inter0, gate268inter1, gate268inter2, gate268inter3, gate268inter4, gate268inter5, gate268inter6, gate268inter7, gate268inter8, gate268inter9, gate268inter10, gate268inter11, gate268inter12, gate423inter0, gate423inter1, gate423inter2, gate423inter3, gate423inter4, gate423inter5, gate423inter6, gate423inter7, gate423inter8, gate423inter9, gate423inter10, gate423inter11, gate423inter12, gate292inter0, gate292inter1, gate292inter2, gate292inter3, gate292inter4, gate292inter5, gate292inter6, gate292inter7, gate292inter8, gate292inter9, gate292inter10, gate292inter11, gate292inter12, gate223inter0, gate223inter1, gate223inter2, gate223inter3, gate223inter4, gate223inter5, gate223inter6, gate223inter7, gate223inter8, gate223inter9, gate223inter10, gate223inter11, gate223inter12, gate473inter0, gate473inter1, gate473inter2, gate473inter3, gate473inter4, gate473inter5, gate473inter6, gate473inter7, gate473inter8, gate473inter9, gate473inter10, gate473inter11, gate473inter12, gate141inter0, gate141inter1, gate141inter2, gate141inter3, gate141inter4, gate141inter5, gate141inter6, gate141inter7, gate141inter8, gate141inter9, gate141inter10, gate141inter11, gate141inter12, gate270inter0, gate270inter1, gate270inter2, gate270inter3, gate270inter4, gate270inter5, gate270inter6, gate270inter7, gate270inter8, gate270inter9, gate270inter10, gate270inter11, gate270inter12, gate471inter0, gate471inter1, gate471inter2, gate471inter3, gate471inter4, gate471inter5, gate471inter6, gate471inter7, gate471inter8, gate471inter9, gate471inter10, gate471inter11, gate471inter12, gate497inter0, gate497inter1, gate497inter2, gate497inter3, gate497inter4, gate497inter5, gate497inter6, gate497inter7, gate497inter8, gate497inter9, gate497inter10, gate497inter11, gate497inter12, gate40inter0, gate40inter1, gate40inter2, gate40inter3, gate40inter4, gate40inter5, gate40inter6, gate40inter7, gate40inter8, gate40inter9, gate40inter10, gate40inter11, gate40inter12, gate102inter0, gate102inter1, gate102inter2, gate102inter3, gate102inter4, gate102inter5, gate102inter6, gate102inter7, gate102inter8, gate102inter9, gate102inter10, gate102inter11, gate102inter12, gate509inter0, gate509inter1, gate509inter2, gate509inter3, gate509inter4, gate509inter5, gate509inter6, gate509inter7, gate509inter8, gate509inter9, gate509inter10, gate509inter11, gate509inter12, gate511inter0, gate511inter1, gate511inter2, gate511inter3, gate511inter4, gate511inter5, gate511inter6, gate511inter7, gate511inter8, gate511inter9, gate511inter10, gate511inter11, gate511inter12, gate78inter0, gate78inter1, gate78inter2, gate78inter3, gate78inter4, gate78inter5, gate78inter6, gate78inter7, gate78inter8, gate78inter9, gate78inter10, gate78inter11, gate78inter12, gate32inter0, gate32inter1, gate32inter2, gate32inter3, gate32inter4, gate32inter5, gate32inter6, gate32inter7, gate32inter8, gate32inter9, gate32inter10, gate32inter11, gate32inter12, gate489inter0, gate489inter1, gate489inter2, gate489inter3, gate489inter4, gate489inter5, gate489inter6, gate489inter7, gate489inter8, gate489inter9, gate489inter10, gate489inter11, gate489inter12, gate87inter0, gate87inter1, gate87inter2, gate87inter3, gate87inter4, gate87inter5, gate87inter6, gate87inter7, gate87inter8, gate87inter9, gate87inter10, gate87inter11, gate87inter12, gate296inter0, gate296inter1, gate296inter2, gate296inter3, gate296inter4, gate296inter5, gate296inter6, gate296inter7, gate296inter8, gate296inter9, gate296inter10, gate296inter11, gate296inter12, gate393inter0, gate393inter1, gate393inter2, gate393inter3, gate393inter4, gate393inter5, gate393inter6, gate393inter7, gate393inter8, gate393inter9, gate393inter10, gate393inter11, gate393inter12, gate111inter0, gate111inter1, gate111inter2, gate111inter3, gate111inter4, gate111inter5, gate111inter6, gate111inter7, gate111inter8, gate111inter9, gate111inter10, gate111inter11, gate111inter12, gate487inter0, gate487inter1, gate487inter2, gate487inter3, gate487inter4, gate487inter5, gate487inter6, gate487inter7, gate487inter8, gate487inter9, gate487inter10, gate487inter11, gate487inter12, gate46inter0, gate46inter1, gate46inter2, gate46inter3, gate46inter4, gate46inter5, gate46inter6, gate46inter7, gate46inter8, gate46inter9, gate46inter10, gate46inter11, gate46inter12, gate178inter0, gate178inter1, gate178inter2, gate178inter3, gate178inter4, gate178inter5, gate178inter6, gate178inter7, gate178inter8, gate178inter9, gate178inter10, gate178inter11, gate178inter12, gate491inter0, gate491inter1, gate491inter2, gate491inter3, gate491inter4, gate491inter5, gate491inter6, gate491inter7, gate491inter8, gate491inter9, gate491inter10, gate491inter11, gate491inter12, gate72inter0, gate72inter1, gate72inter2, gate72inter3, gate72inter4, gate72inter5, gate72inter6, gate72inter7, gate72inter8, gate72inter9, gate72inter10, gate72inter11, gate72inter12, gate145inter0, gate145inter1, gate145inter2, gate145inter3, gate145inter4, gate145inter5, gate145inter6, gate145inter7, gate145inter8, gate145inter9, gate145inter10, gate145inter11, gate145inter12, gate233inter0, gate233inter1, gate233inter2, gate233inter3, gate233inter4, gate233inter5, gate233inter6, gate233inter7, gate233inter8, gate233inter9, gate233inter10, gate233inter11, gate233inter12, gate514inter0, gate514inter1, gate514inter2, gate514inter3, gate514inter4, gate514inter5, gate514inter6, gate514inter7, gate514inter8, gate514inter9, gate514inter10, gate514inter11, gate514inter12, gate152inter0, gate152inter1, gate152inter2, gate152inter3, gate152inter4, gate152inter5, gate152inter6, gate152inter7, gate152inter8, gate152inter9, gate152inter10, gate152inter11, gate152inter12, gate243inter0, gate243inter1, gate243inter2, gate243inter3, gate243inter4, gate243inter5, gate243inter6, gate243inter7, gate243inter8, gate243inter9, gate243inter10, gate243inter11, gate243inter12, gate286inter0, gate286inter1, gate286inter2, gate286inter3, gate286inter4, gate286inter5, gate286inter6, gate286inter7, gate286inter8, gate286inter9, gate286inter10, gate286inter11, gate286inter12, gate417inter0, gate417inter1, gate417inter2, gate417inter3, gate417inter4, gate417inter5, gate417inter6, gate417inter7, gate417inter8, gate417inter9, gate417inter10, gate417inter11, gate417inter12, gate484inter0, gate484inter1, gate484inter2, gate484inter3, gate484inter4, gate484inter5, gate484inter6, gate484inter7, gate484inter8, gate484inter9, gate484inter10, gate484inter11, gate484inter12, gate490inter0, gate490inter1, gate490inter2, gate490inter3, gate490inter4, gate490inter5, gate490inter6, gate490inter7, gate490inter8, gate490inter9, gate490inter10, gate490inter11, gate490inter12, gate34inter0, gate34inter1, gate34inter2, gate34inter3, gate34inter4, gate34inter5, gate34inter6, gate34inter7, gate34inter8, gate34inter9, gate34inter10, gate34inter11, gate34inter12, gate199inter0, gate199inter1, gate199inter2, gate199inter3, gate199inter4, gate199inter5, gate199inter6, gate199inter7, gate199inter8, gate199inter9, gate199inter10, gate199inter11, gate199inter12, gate126inter0, gate126inter1, gate126inter2, gate126inter3, gate126inter4, gate126inter5, gate126inter6, gate126inter7, gate126inter8, gate126inter9, gate126inter10, gate126inter11, gate126inter12, gate255inter0, gate255inter1, gate255inter2, gate255inter3, gate255inter4, gate255inter5, gate255inter6, gate255inter7, gate255inter8, gate255inter9, gate255inter10, gate255inter11, gate255inter12, gate182inter0, gate182inter1, gate182inter2, gate182inter3, gate182inter4, gate182inter5, gate182inter6, gate182inter7, gate182inter8, gate182inter9, gate182inter10, gate182inter11, gate182inter12, gate508inter0, gate508inter1, gate508inter2, gate508inter3, gate508inter4, gate508inter5, gate508inter6, gate508inter7, gate508inter8, gate508inter9, gate508inter10, gate508inter11, gate508inter12, gate74inter0, gate74inter1, gate74inter2, gate74inter3, gate74inter4, gate74inter5, gate74inter6, gate74inter7, gate74inter8, gate74inter9, gate74inter10, gate74inter11, gate74inter12, gate499inter0, gate499inter1, gate499inter2, gate499inter3, gate499inter4, gate499inter5, gate499inter6, gate499inter7, gate499inter8, gate499inter9, gate499inter10, gate499inter11, gate499inter12, gate244inter0, gate244inter1, gate244inter2, gate244inter3, gate244inter4, gate244inter5, gate244inter6, gate244inter7, gate244inter8, gate244inter9, gate244inter10, gate244inter11, gate244inter12, gate19inter0, gate19inter1, gate19inter2, gate19inter3, gate19inter4, gate19inter5, gate19inter6, gate19inter7, gate19inter8, gate19inter9, gate19inter10, gate19inter11, gate19inter12, gate129inter0, gate129inter1, gate129inter2, gate129inter3, gate129inter4, gate129inter5, gate129inter6, gate129inter7, gate129inter8, gate129inter9, gate129inter10, gate129inter11, gate129inter12, gate203inter0, gate203inter1, gate203inter2, gate203inter3, gate203inter4, gate203inter5, gate203inter6, gate203inter7, gate203inter8, gate203inter9, gate203inter10, gate203inter11, gate203inter12, gate149inter0, gate149inter1, gate149inter2, gate149inter3, gate149inter4, gate149inter5, gate149inter6, gate149inter7, gate149inter8, gate149inter9, gate149inter10, gate149inter11, gate149inter12, gate437inter0, gate437inter1, gate437inter2, gate437inter3, gate437inter4, gate437inter5, gate437inter6, gate437inter7, gate437inter8, gate437inter9, gate437inter10, gate437inter11, gate437inter12, gate97inter0, gate97inter1, gate97inter2, gate97inter3, gate97inter4, gate97inter5, gate97inter6, gate97inter7, gate97inter8, gate97inter9, gate97inter10, gate97inter11, gate97inter12, gate26inter0, gate26inter1, gate26inter2, gate26inter3, gate26inter4, gate26inter5, gate26inter6, gate26inter7, gate26inter8, gate26inter9, gate26inter10, gate26inter11, gate26inter12, gate44inter0, gate44inter1, gate44inter2, gate44inter3, gate44inter4, gate44inter5, gate44inter6, gate44inter7, gate44inter8, gate44inter9, gate44inter10, gate44inter11, gate44inter12, gate211inter0, gate211inter1, gate211inter2, gate211inter3, gate211inter4, gate211inter5, gate211inter6, gate211inter7, gate211inter8, gate211inter9, gate211inter10, gate211inter11, gate211inter12, gate162inter0, gate162inter1, gate162inter2, gate162inter3, gate162inter4, gate162inter5, gate162inter6, gate162inter7, gate162inter8, gate162inter9, gate162inter10, gate162inter11, gate162inter12;



and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );
nand2 gate9( .a(G1), .b(G2), .O(G266) );
nand2 gate10( .a(G3), .b(G4), .O(G269) );

  xor2  gate925(.a(G6), .b(G5), .O(gate11inter0));
  nand2 gate926(.a(gate11inter0), .b(s_54), .O(gate11inter1));
  and2  gate927(.a(G6), .b(G5), .O(gate11inter2));
  inv1  gate928(.a(s_54), .O(gate11inter3));
  inv1  gate929(.a(s_55), .O(gate11inter4));
  nand2 gate930(.a(gate11inter4), .b(gate11inter3), .O(gate11inter5));
  nor2  gate931(.a(gate11inter5), .b(gate11inter2), .O(gate11inter6));
  inv1  gate932(.a(G5), .O(gate11inter7));
  inv1  gate933(.a(G6), .O(gate11inter8));
  nand2 gate934(.a(gate11inter8), .b(gate11inter7), .O(gate11inter9));
  nand2 gate935(.a(s_55), .b(gate11inter3), .O(gate11inter10));
  nor2  gate936(.a(gate11inter10), .b(gate11inter9), .O(gate11inter11));
  nor2  gate937(.a(gate11inter11), .b(gate11inter6), .O(gate11inter12));
  nand2 gate938(.a(gate11inter12), .b(gate11inter1), .O(G272));
nand2 gate12( .a(G7), .b(G8), .O(G275) );
nand2 gate13( .a(G9), .b(G10), .O(G278) );
nand2 gate14( .a(G11), .b(G12), .O(G281) );

  xor2  gate715(.a(G14), .b(G13), .O(gate15inter0));
  nand2 gate716(.a(gate15inter0), .b(s_24), .O(gate15inter1));
  and2  gate717(.a(G14), .b(G13), .O(gate15inter2));
  inv1  gate718(.a(s_24), .O(gate15inter3));
  inv1  gate719(.a(s_25), .O(gate15inter4));
  nand2 gate720(.a(gate15inter4), .b(gate15inter3), .O(gate15inter5));
  nor2  gate721(.a(gate15inter5), .b(gate15inter2), .O(gate15inter6));
  inv1  gate722(.a(G13), .O(gate15inter7));
  inv1  gate723(.a(G14), .O(gate15inter8));
  nand2 gate724(.a(gate15inter8), .b(gate15inter7), .O(gate15inter9));
  nand2 gate725(.a(s_25), .b(gate15inter3), .O(gate15inter10));
  nor2  gate726(.a(gate15inter10), .b(gate15inter9), .O(gate15inter11));
  nor2  gate727(.a(gate15inter11), .b(gate15inter6), .O(gate15inter12));
  nand2 gate728(.a(gate15inter12), .b(gate15inter1), .O(G284));
nand2 gate16( .a(G15), .b(G16), .O(G287) );
nand2 gate17( .a(G17), .b(G18), .O(G290) );
nand2 gate18( .a(G19), .b(G20), .O(G293) );

  xor2  gate1961(.a(G22), .b(G21), .O(gate19inter0));
  nand2 gate1962(.a(gate19inter0), .b(s_202), .O(gate19inter1));
  and2  gate1963(.a(G22), .b(G21), .O(gate19inter2));
  inv1  gate1964(.a(s_202), .O(gate19inter3));
  inv1  gate1965(.a(s_203), .O(gate19inter4));
  nand2 gate1966(.a(gate19inter4), .b(gate19inter3), .O(gate19inter5));
  nor2  gate1967(.a(gate19inter5), .b(gate19inter2), .O(gate19inter6));
  inv1  gate1968(.a(G21), .O(gate19inter7));
  inv1  gate1969(.a(G22), .O(gate19inter8));
  nand2 gate1970(.a(gate19inter8), .b(gate19inter7), .O(gate19inter9));
  nand2 gate1971(.a(s_203), .b(gate19inter3), .O(gate19inter10));
  nor2  gate1972(.a(gate19inter10), .b(gate19inter9), .O(gate19inter11));
  nor2  gate1973(.a(gate19inter11), .b(gate19inter6), .O(gate19inter12));
  nand2 gate1974(.a(gate19inter12), .b(gate19inter1), .O(G296));
nand2 gate20( .a(G23), .b(G24), .O(G299) );
nand2 gate21( .a(G25), .b(G26), .O(G302) );
nand2 gate22( .a(G27), .b(G28), .O(G305) );

  xor2  gate1107(.a(G30), .b(G29), .O(gate23inter0));
  nand2 gate1108(.a(gate23inter0), .b(s_80), .O(gate23inter1));
  and2  gate1109(.a(G30), .b(G29), .O(gate23inter2));
  inv1  gate1110(.a(s_80), .O(gate23inter3));
  inv1  gate1111(.a(s_81), .O(gate23inter4));
  nand2 gate1112(.a(gate23inter4), .b(gate23inter3), .O(gate23inter5));
  nor2  gate1113(.a(gate23inter5), .b(gate23inter2), .O(gate23inter6));
  inv1  gate1114(.a(G29), .O(gate23inter7));
  inv1  gate1115(.a(G30), .O(gate23inter8));
  nand2 gate1116(.a(gate23inter8), .b(gate23inter7), .O(gate23inter9));
  nand2 gate1117(.a(s_81), .b(gate23inter3), .O(gate23inter10));
  nor2  gate1118(.a(gate23inter10), .b(gate23inter9), .O(gate23inter11));
  nor2  gate1119(.a(gate23inter11), .b(gate23inter6), .O(gate23inter12));
  nand2 gate1120(.a(gate23inter12), .b(gate23inter1), .O(G308));
nand2 gate24( .a(G31), .b(G32), .O(G311) );
nand2 gate25( .a(G1), .b(G5), .O(G314) );

  xor2  gate2045(.a(G13), .b(G9), .O(gate26inter0));
  nand2 gate2046(.a(gate26inter0), .b(s_214), .O(gate26inter1));
  and2  gate2047(.a(G13), .b(G9), .O(gate26inter2));
  inv1  gate2048(.a(s_214), .O(gate26inter3));
  inv1  gate2049(.a(s_215), .O(gate26inter4));
  nand2 gate2050(.a(gate26inter4), .b(gate26inter3), .O(gate26inter5));
  nor2  gate2051(.a(gate26inter5), .b(gate26inter2), .O(gate26inter6));
  inv1  gate2052(.a(G9), .O(gate26inter7));
  inv1  gate2053(.a(G13), .O(gate26inter8));
  nand2 gate2054(.a(gate26inter8), .b(gate26inter7), .O(gate26inter9));
  nand2 gate2055(.a(s_215), .b(gate26inter3), .O(gate26inter10));
  nor2  gate2056(.a(gate26inter10), .b(gate26inter9), .O(gate26inter11));
  nor2  gate2057(.a(gate26inter11), .b(gate26inter6), .O(gate26inter12));
  nand2 gate2058(.a(gate26inter12), .b(gate26inter1), .O(G317));
nand2 gate27( .a(G2), .b(G6), .O(G320) );
nand2 gate28( .a(G10), .b(G14), .O(G323) );
nand2 gate29( .a(G3), .b(G7), .O(G326) );
nand2 gate30( .a(G11), .b(G15), .O(G329) );

  xor2  gate1177(.a(G8), .b(G4), .O(gate31inter0));
  nand2 gate1178(.a(gate31inter0), .b(s_90), .O(gate31inter1));
  and2  gate1179(.a(G8), .b(G4), .O(gate31inter2));
  inv1  gate1180(.a(s_90), .O(gate31inter3));
  inv1  gate1181(.a(s_91), .O(gate31inter4));
  nand2 gate1182(.a(gate31inter4), .b(gate31inter3), .O(gate31inter5));
  nor2  gate1183(.a(gate31inter5), .b(gate31inter2), .O(gate31inter6));
  inv1  gate1184(.a(G4), .O(gate31inter7));
  inv1  gate1185(.a(G8), .O(gate31inter8));
  nand2 gate1186(.a(gate31inter8), .b(gate31inter7), .O(gate31inter9));
  nand2 gate1187(.a(s_91), .b(gate31inter3), .O(gate31inter10));
  nor2  gate1188(.a(gate31inter10), .b(gate31inter9), .O(gate31inter11));
  nor2  gate1189(.a(gate31inter11), .b(gate31inter6), .O(gate31inter12));
  nand2 gate1190(.a(gate31inter12), .b(gate31inter1), .O(G332));

  xor2  gate1555(.a(G16), .b(G12), .O(gate32inter0));
  nand2 gate1556(.a(gate32inter0), .b(s_144), .O(gate32inter1));
  and2  gate1557(.a(G16), .b(G12), .O(gate32inter2));
  inv1  gate1558(.a(s_144), .O(gate32inter3));
  inv1  gate1559(.a(s_145), .O(gate32inter4));
  nand2 gate1560(.a(gate32inter4), .b(gate32inter3), .O(gate32inter5));
  nor2  gate1561(.a(gate32inter5), .b(gate32inter2), .O(gate32inter6));
  inv1  gate1562(.a(G12), .O(gate32inter7));
  inv1  gate1563(.a(G16), .O(gate32inter8));
  nand2 gate1564(.a(gate32inter8), .b(gate32inter7), .O(gate32inter9));
  nand2 gate1565(.a(s_145), .b(gate32inter3), .O(gate32inter10));
  nor2  gate1566(.a(gate32inter10), .b(gate32inter9), .O(gate32inter11));
  nor2  gate1567(.a(gate32inter11), .b(gate32inter6), .O(gate32inter12));
  nand2 gate1568(.a(gate32inter12), .b(gate32inter1), .O(G335));
nand2 gate33( .a(G17), .b(G21), .O(G338) );

  xor2  gate1835(.a(G29), .b(G25), .O(gate34inter0));
  nand2 gate1836(.a(gate34inter0), .b(s_184), .O(gate34inter1));
  and2  gate1837(.a(G29), .b(G25), .O(gate34inter2));
  inv1  gate1838(.a(s_184), .O(gate34inter3));
  inv1  gate1839(.a(s_185), .O(gate34inter4));
  nand2 gate1840(.a(gate34inter4), .b(gate34inter3), .O(gate34inter5));
  nor2  gate1841(.a(gate34inter5), .b(gate34inter2), .O(gate34inter6));
  inv1  gate1842(.a(G25), .O(gate34inter7));
  inv1  gate1843(.a(G29), .O(gate34inter8));
  nand2 gate1844(.a(gate34inter8), .b(gate34inter7), .O(gate34inter9));
  nand2 gate1845(.a(s_185), .b(gate34inter3), .O(gate34inter10));
  nor2  gate1846(.a(gate34inter10), .b(gate34inter9), .O(gate34inter11));
  nor2  gate1847(.a(gate34inter11), .b(gate34inter6), .O(gate34inter12));
  nand2 gate1848(.a(gate34inter12), .b(gate34inter1), .O(G341));
nand2 gate35( .a(G18), .b(G22), .O(G344) );
nand2 gate36( .a(G26), .b(G30), .O(G347) );
nand2 gate37( .a(G19), .b(G23), .O(G350) );
nand2 gate38( .a(G27), .b(G31), .O(G353) );
nand2 gate39( .a(G20), .b(G24), .O(G356) );

  xor2  gate1485(.a(G32), .b(G28), .O(gate40inter0));
  nand2 gate1486(.a(gate40inter0), .b(s_134), .O(gate40inter1));
  and2  gate1487(.a(G32), .b(G28), .O(gate40inter2));
  inv1  gate1488(.a(s_134), .O(gate40inter3));
  inv1  gate1489(.a(s_135), .O(gate40inter4));
  nand2 gate1490(.a(gate40inter4), .b(gate40inter3), .O(gate40inter5));
  nor2  gate1491(.a(gate40inter5), .b(gate40inter2), .O(gate40inter6));
  inv1  gate1492(.a(G28), .O(gate40inter7));
  inv1  gate1493(.a(G32), .O(gate40inter8));
  nand2 gate1494(.a(gate40inter8), .b(gate40inter7), .O(gate40inter9));
  nand2 gate1495(.a(s_135), .b(gate40inter3), .O(gate40inter10));
  nor2  gate1496(.a(gate40inter10), .b(gate40inter9), .O(gate40inter11));
  nor2  gate1497(.a(gate40inter11), .b(gate40inter6), .O(gate40inter12));
  nand2 gate1498(.a(gate40inter12), .b(gate40inter1), .O(G359));
nand2 gate41( .a(G1), .b(G266), .O(G362) );
nand2 gate42( .a(G2), .b(G266), .O(G363) );
nand2 gate43( .a(G3), .b(G269), .O(G364) );

  xor2  gate2059(.a(G269), .b(G4), .O(gate44inter0));
  nand2 gate2060(.a(gate44inter0), .b(s_216), .O(gate44inter1));
  and2  gate2061(.a(G269), .b(G4), .O(gate44inter2));
  inv1  gate2062(.a(s_216), .O(gate44inter3));
  inv1  gate2063(.a(s_217), .O(gate44inter4));
  nand2 gate2064(.a(gate44inter4), .b(gate44inter3), .O(gate44inter5));
  nor2  gate2065(.a(gate44inter5), .b(gate44inter2), .O(gate44inter6));
  inv1  gate2066(.a(G4), .O(gate44inter7));
  inv1  gate2067(.a(G269), .O(gate44inter8));
  nand2 gate2068(.a(gate44inter8), .b(gate44inter7), .O(gate44inter9));
  nand2 gate2069(.a(s_217), .b(gate44inter3), .O(gate44inter10));
  nor2  gate2070(.a(gate44inter10), .b(gate44inter9), .O(gate44inter11));
  nor2  gate2071(.a(gate44inter11), .b(gate44inter6), .O(gate44inter12));
  nand2 gate2072(.a(gate44inter12), .b(gate44inter1), .O(G365));

  xor2  gate1149(.a(G272), .b(G5), .O(gate45inter0));
  nand2 gate1150(.a(gate45inter0), .b(s_86), .O(gate45inter1));
  and2  gate1151(.a(G272), .b(G5), .O(gate45inter2));
  inv1  gate1152(.a(s_86), .O(gate45inter3));
  inv1  gate1153(.a(s_87), .O(gate45inter4));
  nand2 gate1154(.a(gate45inter4), .b(gate45inter3), .O(gate45inter5));
  nor2  gate1155(.a(gate45inter5), .b(gate45inter2), .O(gate45inter6));
  inv1  gate1156(.a(G5), .O(gate45inter7));
  inv1  gate1157(.a(G272), .O(gate45inter8));
  nand2 gate1158(.a(gate45inter8), .b(gate45inter7), .O(gate45inter9));
  nand2 gate1159(.a(s_87), .b(gate45inter3), .O(gate45inter10));
  nor2  gate1160(.a(gate45inter10), .b(gate45inter9), .O(gate45inter11));
  nor2  gate1161(.a(gate45inter11), .b(gate45inter6), .O(gate45inter12));
  nand2 gate1162(.a(gate45inter12), .b(gate45inter1), .O(G366));

  xor2  gate1653(.a(G272), .b(G6), .O(gate46inter0));
  nand2 gate1654(.a(gate46inter0), .b(s_158), .O(gate46inter1));
  and2  gate1655(.a(G272), .b(G6), .O(gate46inter2));
  inv1  gate1656(.a(s_158), .O(gate46inter3));
  inv1  gate1657(.a(s_159), .O(gate46inter4));
  nand2 gate1658(.a(gate46inter4), .b(gate46inter3), .O(gate46inter5));
  nor2  gate1659(.a(gate46inter5), .b(gate46inter2), .O(gate46inter6));
  inv1  gate1660(.a(G6), .O(gate46inter7));
  inv1  gate1661(.a(G272), .O(gate46inter8));
  nand2 gate1662(.a(gate46inter8), .b(gate46inter7), .O(gate46inter9));
  nand2 gate1663(.a(s_159), .b(gate46inter3), .O(gate46inter10));
  nor2  gate1664(.a(gate46inter10), .b(gate46inter9), .O(gate46inter11));
  nor2  gate1665(.a(gate46inter11), .b(gate46inter6), .O(gate46inter12));
  nand2 gate1666(.a(gate46inter12), .b(gate46inter1), .O(G367));
nand2 gate47( .a(G7), .b(G275), .O(G368) );
nand2 gate48( .a(G8), .b(G275), .O(G369) );
nand2 gate49( .a(G9), .b(G278), .O(G370) );
nand2 gate50( .a(G10), .b(G278), .O(G371) );
nand2 gate51( .a(G11), .b(G281), .O(G372) );
nand2 gate52( .a(G12), .b(G281), .O(G373) );
nand2 gate53( .a(G13), .b(G284), .O(G374) );
nand2 gate54( .a(G14), .b(G284), .O(G375) );
nand2 gate55( .a(G15), .b(G287), .O(G376) );

  xor2  gate1191(.a(G287), .b(G16), .O(gate56inter0));
  nand2 gate1192(.a(gate56inter0), .b(s_92), .O(gate56inter1));
  and2  gate1193(.a(G287), .b(G16), .O(gate56inter2));
  inv1  gate1194(.a(s_92), .O(gate56inter3));
  inv1  gate1195(.a(s_93), .O(gate56inter4));
  nand2 gate1196(.a(gate56inter4), .b(gate56inter3), .O(gate56inter5));
  nor2  gate1197(.a(gate56inter5), .b(gate56inter2), .O(gate56inter6));
  inv1  gate1198(.a(G16), .O(gate56inter7));
  inv1  gate1199(.a(G287), .O(gate56inter8));
  nand2 gate1200(.a(gate56inter8), .b(gate56inter7), .O(gate56inter9));
  nand2 gate1201(.a(s_93), .b(gate56inter3), .O(gate56inter10));
  nor2  gate1202(.a(gate56inter10), .b(gate56inter9), .O(gate56inter11));
  nor2  gate1203(.a(gate56inter11), .b(gate56inter6), .O(gate56inter12));
  nand2 gate1204(.a(gate56inter12), .b(gate56inter1), .O(G377));
nand2 gate57( .a(G17), .b(G290), .O(G378) );
nand2 gate58( .a(G18), .b(G290), .O(G379) );
nand2 gate59( .a(G19), .b(G293), .O(G380) );

  xor2  gate855(.a(G293), .b(G20), .O(gate60inter0));
  nand2 gate856(.a(gate60inter0), .b(s_44), .O(gate60inter1));
  and2  gate857(.a(G293), .b(G20), .O(gate60inter2));
  inv1  gate858(.a(s_44), .O(gate60inter3));
  inv1  gate859(.a(s_45), .O(gate60inter4));
  nand2 gate860(.a(gate60inter4), .b(gate60inter3), .O(gate60inter5));
  nor2  gate861(.a(gate60inter5), .b(gate60inter2), .O(gate60inter6));
  inv1  gate862(.a(G20), .O(gate60inter7));
  inv1  gate863(.a(G293), .O(gate60inter8));
  nand2 gate864(.a(gate60inter8), .b(gate60inter7), .O(gate60inter9));
  nand2 gate865(.a(s_45), .b(gate60inter3), .O(gate60inter10));
  nor2  gate866(.a(gate60inter10), .b(gate60inter9), .O(gate60inter11));
  nor2  gate867(.a(gate60inter11), .b(gate60inter6), .O(gate60inter12));
  nand2 gate868(.a(gate60inter12), .b(gate60inter1), .O(G381));
nand2 gate61( .a(G21), .b(G296), .O(G382) );
nand2 gate62( .a(G22), .b(G296), .O(G383) );

  xor2  gate841(.a(G299), .b(G23), .O(gate63inter0));
  nand2 gate842(.a(gate63inter0), .b(s_42), .O(gate63inter1));
  and2  gate843(.a(G299), .b(G23), .O(gate63inter2));
  inv1  gate844(.a(s_42), .O(gate63inter3));
  inv1  gate845(.a(s_43), .O(gate63inter4));
  nand2 gate846(.a(gate63inter4), .b(gate63inter3), .O(gate63inter5));
  nor2  gate847(.a(gate63inter5), .b(gate63inter2), .O(gate63inter6));
  inv1  gate848(.a(G23), .O(gate63inter7));
  inv1  gate849(.a(G299), .O(gate63inter8));
  nand2 gate850(.a(gate63inter8), .b(gate63inter7), .O(gate63inter9));
  nand2 gate851(.a(s_43), .b(gate63inter3), .O(gate63inter10));
  nor2  gate852(.a(gate63inter10), .b(gate63inter9), .O(gate63inter11));
  nor2  gate853(.a(gate63inter11), .b(gate63inter6), .O(gate63inter12));
  nand2 gate854(.a(gate63inter12), .b(gate63inter1), .O(G384));
nand2 gate64( .a(G24), .b(G299), .O(G385) );
nand2 gate65( .a(G25), .b(G302), .O(G386) );
nand2 gate66( .a(G26), .b(G302), .O(G387) );
nand2 gate67( .a(G27), .b(G305), .O(G388) );

  xor2  gate827(.a(G305), .b(G28), .O(gate68inter0));
  nand2 gate828(.a(gate68inter0), .b(s_40), .O(gate68inter1));
  and2  gate829(.a(G305), .b(G28), .O(gate68inter2));
  inv1  gate830(.a(s_40), .O(gate68inter3));
  inv1  gate831(.a(s_41), .O(gate68inter4));
  nand2 gate832(.a(gate68inter4), .b(gate68inter3), .O(gate68inter5));
  nor2  gate833(.a(gate68inter5), .b(gate68inter2), .O(gate68inter6));
  inv1  gate834(.a(G28), .O(gate68inter7));
  inv1  gate835(.a(G305), .O(gate68inter8));
  nand2 gate836(.a(gate68inter8), .b(gate68inter7), .O(gate68inter9));
  nand2 gate837(.a(s_41), .b(gate68inter3), .O(gate68inter10));
  nor2  gate838(.a(gate68inter10), .b(gate68inter9), .O(gate68inter11));
  nor2  gate839(.a(gate68inter11), .b(gate68inter6), .O(gate68inter12));
  nand2 gate840(.a(gate68inter12), .b(gate68inter1), .O(G389));
nand2 gate69( .a(G29), .b(G308), .O(G390) );
nand2 gate70( .a(G30), .b(G308), .O(G391) );
nand2 gate71( .a(G31), .b(G311), .O(G392) );

  xor2  gate1695(.a(G311), .b(G32), .O(gate72inter0));
  nand2 gate1696(.a(gate72inter0), .b(s_164), .O(gate72inter1));
  and2  gate1697(.a(G311), .b(G32), .O(gate72inter2));
  inv1  gate1698(.a(s_164), .O(gate72inter3));
  inv1  gate1699(.a(s_165), .O(gate72inter4));
  nand2 gate1700(.a(gate72inter4), .b(gate72inter3), .O(gate72inter5));
  nor2  gate1701(.a(gate72inter5), .b(gate72inter2), .O(gate72inter6));
  inv1  gate1702(.a(G32), .O(gate72inter7));
  inv1  gate1703(.a(G311), .O(gate72inter8));
  nand2 gate1704(.a(gate72inter8), .b(gate72inter7), .O(gate72inter9));
  nand2 gate1705(.a(s_165), .b(gate72inter3), .O(gate72inter10));
  nor2  gate1706(.a(gate72inter10), .b(gate72inter9), .O(gate72inter11));
  nor2  gate1707(.a(gate72inter11), .b(gate72inter6), .O(gate72inter12));
  nand2 gate1708(.a(gate72inter12), .b(gate72inter1), .O(G393));
nand2 gate73( .a(G1), .b(G314), .O(G394) );

  xor2  gate1919(.a(G314), .b(G5), .O(gate74inter0));
  nand2 gate1920(.a(gate74inter0), .b(s_196), .O(gate74inter1));
  and2  gate1921(.a(G314), .b(G5), .O(gate74inter2));
  inv1  gate1922(.a(s_196), .O(gate74inter3));
  inv1  gate1923(.a(s_197), .O(gate74inter4));
  nand2 gate1924(.a(gate74inter4), .b(gate74inter3), .O(gate74inter5));
  nor2  gate1925(.a(gate74inter5), .b(gate74inter2), .O(gate74inter6));
  inv1  gate1926(.a(G5), .O(gate74inter7));
  inv1  gate1927(.a(G314), .O(gate74inter8));
  nand2 gate1928(.a(gate74inter8), .b(gate74inter7), .O(gate74inter9));
  nand2 gate1929(.a(s_197), .b(gate74inter3), .O(gate74inter10));
  nor2  gate1930(.a(gate74inter10), .b(gate74inter9), .O(gate74inter11));
  nor2  gate1931(.a(gate74inter11), .b(gate74inter6), .O(gate74inter12));
  nand2 gate1932(.a(gate74inter12), .b(gate74inter1), .O(G395));
nand2 gate75( .a(G9), .b(G317), .O(G396) );
nand2 gate76( .a(G13), .b(G317), .O(G397) );
nand2 gate77( .a(G2), .b(G320), .O(G398) );

  xor2  gate1541(.a(G320), .b(G6), .O(gate78inter0));
  nand2 gate1542(.a(gate78inter0), .b(s_142), .O(gate78inter1));
  and2  gate1543(.a(G320), .b(G6), .O(gate78inter2));
  inv1  gate1544(.a(s_142), .O(gate78inter3));
  inv1  gate1545(.a(s_143), .O(gate78inter4));
  nand2 gate1546(.a(gate78inter4), .b(gate78inter3), .O(gate78inter5));
  nor2  gate1547(.a(gate78inter5), .b(gate78inter2), .O(gate78inter6));
  inv1  gate1548(.a(G6), .O(gate78inter7));
  inv1  gate1549(.a(G320), .O(gate78inter8));
  nand2 gate1550(.a(gate78inter8), .b(gate78inter7), .O(gate78inter9));
  nand2 gate1551(.a(s_143), .b(gate78inter3), .O(gate78inter10));
  nor2  gate1552(.a(gate78inter10), .b(gate78inter9), .O(gate78inter11));
  nor2  gate1553(.a(gate78inter11), .b(gate78inter6), .O(gate78inter12));
  nand2 gate1554(.a(gate78inter12), .b(gate78inter1), .O(G399));
nand2 gate79( .a(G10), .b(G323), .O(G400) );
nand2 gate80( .a(G14), .b(G323), .O(G401) );
nand2 gate81( .a(G3), .b(G326), .O(G402) );
nand2 gate82( .a(G7), .b(G326), .O(G403) );
nand2 gate83( .a(G11), .b(G329), .O(G404) );
nand2 gate84( .a(G15), .b(G329), .O(G405) );
nand2 gate85( .a(G4), .b(G332), .O(G406) );
nand2 gate86( .a(G8), .b(G332), .O(G407) );

  xor2  gate1583(.a(G335), .b(G12), .O(gate87inter0));
  nand2 gate1584(.a(gate87inter0), .b(s_148), .O(gate87inter1));
  and2  gate1585(.a(G335), .b(G12), .O(gate87inter2));
  inv1  gate1586(.a(s_148), .O(gate87inter3));
  inv1  gate1587(.a(s_149), .O(gate87inter4));
  nand2 gate1588(.a(gate87inter4), .b(gate87inter3), .O(gate87inter5));
  nor2  gate1589(.a(gate87inter5), .b(gate87inter2), .O(gate87inter6));
  inv1  gate1590(.a(G12), .O(gate87inter7));
  inv1  gate1591(.a(G335), .O(gate87inter8));
  nand2 gate1592(.a(gate87inter8), .b(gate87inter7), .O(gate87inter9));
  nand2 gate1593(.a(s_149), .b(gate87inter3), .O(gate87inter10));
  nor2  gate1594(.a(gate87inter10), .b(gate87inter9), .O(gate87inter11));
  nor2  gate1595(.a(gate87inter11), .b(gate87inter6), .O(gate87inter12));
  nand2 gate1596(.a(gate87inter12), .b(gate87inter1), .O(G408));
nand2 gate88( .a(G16), .b(G335), .O(G409) );

  xor2  gate1219(.a(G338), .b(G17), .O(gate89inter0));
  nand2 gate1220(.a(gate89inter0), .b(s_96), .O(gate89inter1));
  and2  gate1221(.a(G338), .b(G17), .O(gate89inter2));
  inv1  gate1222(.a(s_96), .O(gate89inter3));
  inv1  gate1223(.a(s_97), .O(gate89inter4));
  nand2 gate1224(.a(gate89inter4), .b(gate89inter3), .O(gate89inter5));
  nor2  gate1225(.a(gate89inter5), .b(gate89inter2), .O(gate89inter6));
  inv1  gate1226(.a(G17), .O(gate89inter7));
  inv1  gate1227(.a(G338), .O(gate89inter8));
  nand2 gate1228(.a(gate89inter8), .b(gate89inter7), .O(gate89inter9));
  nand2 gate1229(.a(s_97), .b(gate89inter3), .O(gate89inter10));
  nor2  gate1230(.a(gate89inter10), .b(gate89inter9), .O(gate89inter11));
  nor2  gate1231(.a(gate89inter11), .b(gate89inter6), .O(gate89inter12));
  nand2 gate1232(.a(gate89inter12), .b(gate89inter1), .O(G410));
nand2 gate90( .a(G21), .b(G338), .O(G411) );
nand2 gate91( .a(G25), .b(G341), .O(G412) );

  xor2  gate561(.a(G341), .b(G29), .O(gate92inter0));
  nand2 gate562(.a(gate92inter0), .b(s_2), .O(gate92inter1));
  and2  gate563(.a(G341), .b(G29), .O(gate92inter2));
  inv1  gate564(.a(s_2), .O(gate92inter3));
  inv1  gate565(.a(s_3), .O(gate92inter4));
  nand2 gate566(.a(gate92inter4), .b(gate92inter3), .O(gate92inter5));
  nor2  gate567(.a(gate92inter5), .b(gate92inter2), .O(gate92inter6));
  inv1  gate568(.a(G29), .O(gate92inter7));
  inv1  gate569(.a(G341), .O(gate92inter8));
  nand2 gate570(.a(gate92inter8), .b(gate92inter7), .O(gate92inter9));
  nand2 gate571(.a(s_3), .b(gate92inter3), .O(gate92inter10));
  nor2  gate572(.a(gate92inter10), .b(gate92inter9), .O(gate92inter11));
  nor2  gate573(.a(gate92inter11), .b(gate92inter6), .O(gate92inter12));
  nand2 gate574(.a(gate92inter12), .b(gate92inter1), .O(G413));
nand2 gate93( .a(G18), .b(G344), .O(G414) );
nand2 gate94( .a(G22), .b(G344), .O(G415) );
nand2 gate95( .a(G26), .b(G347), .O(G416) );
nand2 gate96( .a(G30), .b(G347), .O(G417) );

  xor2  gate2031(.a(G350), .b(G19), .O(gate97inter0));
  nand2 gate2032(.a(gate97inter0), .b(s_212), .O(gate97inter1));
  and2  gate2033(.a(G350), .b(G19), .O(gate97inter2));
  inv1  gate2034(.a(s_212), .O(gate97inter3));
  inv1  gate2035(.a(s_213), .O(gate97inter4));
  nand2 gate2036(.a(gate97inter4), .b(gate97inter3), .O(gate97inter5));
  nor2  gate2037(.a(gate97inter5), .b(gate97inter2), .O(gate97inter6));
  inv1  gate2038(.a(G19), .O(gate97inter7));
  inv1  gate2039(.a(G350), .O(gate97inter8));
  nand2 gate2040(.a(gate97inter8), .b(gate97inter7), .O(gate97inter9));
  nand2 gate2041(.a(s_213), .b(gate97inter3), .O(gate97inter10));
  nor2  gate2042(.a(gate97inter10), .b(gate97inter9), .O(gate97inter11));
  nor2  gate2043(.a(gate97inter11), .b(gate97inter6), .O(gate97inter12));
  nand2 gate2044(.a(gate97inter12), .b(gate97inter1), .O(G418));
nand2 gate98( .a(G23), .b(G350), .O(G419) );
nand2 gate99( .a(G27), .b(G353), .O(G420) );
nand2 gate100( .a(G31), .b(G353), .O(G421) );
nand2 gate101( .a(G20), .b(G356), .O(G422) );

  xor2  gate1499(.a(G356), .b(G24), .O(gate102inter0));
  nand2 gate1500(.a(gate102inter0), .b(s_136), .O(gate102inter1));
  and2  gate1501(.a(G356), .b(G24), .O(gate102inter2));
  inv1  gate1502(.a(s_136), .O(gate102inter3));
  inv1  gate1503(.a(s_137), .O(gate102inter4));
  nand2 gate1504(.a(gate102inter4), .b(gate102inter3), .O(gate102inter5));
  nor2  gate1505(.a(gate102inter5), .b(gate102inter2), .O(gate102inter6));
  inv1  gate1506(.a(G24), .O(gate102inter7));
  inv1  gate1507(.a(G356), .O(gate102inter8));
  nand2 gate1508(.a(gate102inter8), .b(gate102inter7), .O(gate102inter9));
  nand2 gate1509(.a(s_137), .b(gate102inter3), .O(gate102inter10));
  nor2  gate1510(.a(gate102inter10), .b(gate102inter9), .O(gate102inter11));
  nor2  gate1511(.a(gate102inter11), .b(gate102inter6), .O(gate102inter12));
  nand2 gate1512(.a(gate102inter12), .b(gate102inter1), .O(G423));
nand2 gate103( .a(G28), .b(G359), .O(G424) );
nand2 gate104( .a(G32), .b(G359), .O(G425) );

  xor2  gate771(.a(G363), .b(G362), .O(gate105inter0));
  nand2 gate772(.a(gate105inter0), .b(s_32), .O(gate105inter1));
  and2  gate773(.a(G363), .b(G362), .O(gate105inter2));
  inv1  gate774(.a(s_32), .O(gate105inter3));
  inv1  gate775(.a(s_33), .O(gate105inter4));
  nand2 gate776(.a(gate105inter4), .b(gate105inter3), .O(gate105inter5));
  nor2  gate777(.a(gate105inter5), .b(gate105inter2), .O(gate105inter6));
  inv1  gate778(.a(G362), .O(gate105inter7));
  inv1  gate779(.a(G363), .O(gate105inter8));
  nand2 gate780(.a(gate105inter8), .b(gate105inter7), .O(gate105inter9));
  nand2 gate781(.a(s_33), .b(gate105inter3), .O(gate105inter10));
  nor2  gate782(.a(gate105inter10), .b(gate105inter9), .O(gate105inter11));
  nor2  gate783(.a(gate105inter11), .b(gate105inter6), .O(gate105inter12));
  nand2 gate784(.a(gate105inter12), .b(gate105inter1), .O(G426));
nand2 gate106( .a(G364), .b(G365), .O(G429) );
nand2 gate107( .a(G366), .b(G367), .O(G432) );

  xor2  gate547(.a(G369), .b(G368), .O(gate108inter0));
  nand2 gate548(.a(gate108inter0), .b(s_0), .O(gate108inter1));
  and2  gate549(.a(G369), .b(G368), .O(gate108inter2));
  inv1  gate550(.a(s_0), .O(gate108inter3));
  inv1  gate551(.a(s_1), .O(gate108inter4));
  nand2 gate552(.a(gate108inter4), .b(gate108inter3), .O(gate108inter5));
  nor2  gate553(.a(gate108inter5), .b(gate108inter2), .O(gate108inter6));
  inv1  gate554(.a(G368), .O(gate108inter7));
  inv1  gate555(.a(G369), .O(gate108inter8));
  nand2 gate556(.a(gate108inter8), .b(gate108inter7), .O(gate108inter9));
  nand2 gate557(.a(s_1), .b(gate108inter3), .O(gate108inter10));
  nor2  gate558(.a(gate108inter10), .b(gate108inter9), .O(gate108inter11));
  nor2  gate559(.a(gate108inter11), .b(gate108inter6), .O(gate108inter12));
  nand2 gate560(.a(gate108inter12), .b(gate108inter1), .O(G435));
nand2 gate109( .a(G370), .b(G371), .O(G438) );
nand2 gate110( .a(G372), .b(G373), .O(G441) );

  xor2  gate1625(.a(G375), .b(G374), .O(gate111inter0));
  nand2 gate1626(.a(gate111inter0), .b(s_154), .O(gate111inter1));
  and2  gate1627(.a(G375), .b(G374), .O(gate111inter2));
  inv1  gate1628(.a(s_154), .O(gate111inter3));
  inv1  gate1629(.a(s_155), .O(gate111inter4));
  nand2 gate1630(.a(gate111inter4), .b(gate111inter3), .O(gate111inter5));
  nor2  gate1631(.a(gate111inter5), .b(gate111inter2), .O(gate111inter6));
  inv1  gate1632(.a(G374), .O(gate111inter7));
  inv1  gate1633(.a(G375), .O(gate111inter8));
  nand2 gate1634(.a(gate111inter8), .b(gate111inter7), .O(gate111inter9));
  nand2 gate1635(.a(s_155), .b(gate111inter3), .O(gate111inter10));
  nor2  gate1636(.a(gate111inter10), .b(gate111inter9), .O(gate111inter11));
  nor2  gate1637(.a(gate111inter11), .b(gate111inter6), .O(gate111inter12));
  nand2 gate1638(.a(gate111inter12), .b(gate111inter1), .O(G444));
nand2 gate112( .a(G376), .b(G377), .O(G447) );
nand2 gate113( .a(G378), .b(G379), .O(G450) );
nand2 gate114( .a(G380), .b(G381), .O(G453) );
nand2 gate115( .a(G382), .b(G383), .O(G456) );

  xor2  gate743(.a(G385), .b(G384), .O(gate116inter0));
  nand2 gate744(.a(gate116inter0), .b(s_28), .O(gate116inter1));
  and2  gate745(.a(G385), .b(G384), .O(gate116inter2));
  inv1  gate746(.a(s_28), .O(gate116inter3));
  inv1  gate747(.a(s_29), .O(gate116inter4));
  nand2 gate748(.a(gate116inter4), .b(gate116inter3), .O(gate116inter5));
  nor2  gate749(.a(gate116inter5), .b(gate116inter2), .O(gate116inter6));
  inv1  gate750(.a(G384), .O(gate116inter7));
  inv1  gate751(.a(G385), .O(gate116inter8));
  nand2 gate752(.a(gate116inter8), .b(gate116inter7), .O(gate116inter9));
  nand2 gate753(.a(s_29), .b(gate116inter3), .O(gate116inter10));
  nor2  gate754(.a(gate116inter10), .b(gate116inter9), .O(gate116inter11));
  nor2  gate755(.a(gate116inter11), .b(gate116inter6), .O(gate116inter12));
  nand2 gate756(.a(gate116inter12), .b(gate116inter1), .O(G459));
nand2 gate117( .a(G386), .b(G387), .O(G462) );
nand2 gate118( .a(G388), .b(G389), .O(G465) );
nand2 gate119( .a(G390), .b(G391), .O(G468) );

  xor2  gate589(.a(G393), .b(G392), .O(gate120inter0));
  nand2 gate590(.a(gate120inter0), .b(s_6), .O(gate120inter1));
  and2  gate591(.a(G393), .b(G392), .O(gate120inter2));
  inv1  gate592(.a(s_6), .O(gate120inter3));
  inv1  gate593(.a(s_7), .O(gate120inter4));
  nand2 gate594(.a(gate120inter4), .b(gate120inter3), .O(gate120inter5));
  nor2  gate595(.a(gate120inter5), .b(gate120inter2), .O(gate120inter6));
  inv1  gate596(.a(G392), .O(gate120inter7));
  inv1  gate597(.a(G393), .O(gate120inter8));
  nand2 gate598(.a(gate120inter8), .b(gate120inter7), .O(gate120inter9));
  nand2 gate599(.a(s_7), .b(gate120inter3), .O(gate120inter10));
  nor2  gate600(.a(gate120inter10), .b(gate120inter9), .O(gate120inter11));
  nor2  gate601(.a(gate120inter11), .b(gate120inter6), .O(gate120inter12));
  nand2 gate602(.a(gate120inter12), .b(gate120inter1), .O(G471));
nand2 gate121( .a(G394), .b(G395), .O(G474) );
nand2 gate122( .a(G396), .b(G397), .O(G477) );
nand2 gate123( .a(G398), .b(G399), .O(G480) );
nand2 gate124( .a(G400), .b(G401), .O(G483) );
nand2 gate125( .a(G402), .b(G403), .O(G486) );

  xor2  gate1863(.a(G405), .b(G404), .O(gate126inter0));
  nand2 gate1864(.a(gate126inter0), .b(s_188), .O(gate126inter1));
  and2  gate1865(.a(G405), .b(G404), .O(gate126inter2));
  inv1  gate1866(.a(s_188), .O(gate126inter3));
  inv1  gate1867(.a(s_189), .O(gate126inter4));
  nand2 gate1868(.a(gate126inter4), .b(gate126inter3), .O(gate126inter5));
  nor2  gate1869(.a(gate126inter5), .b(gate126inter2), .O(gate126inter6));
  inv1  gate1870(.a(G404), .O(gate126inter7));
  inv1  gate1871(.a(G405), .O(gate126inter8));
  nand2 gate1872(.a(gate126inter8), .b(gate126inter7), .O(gate126inter9));
  nand2 gate1873(.a(s_189), .b(gate126inter3), .O(gate126inter10));
  nor2  gate1874(.a(gate126inter10), .b(gate126inter9), .O(gate126inter11));
  nor2  gate1875(.a(gate126inter11), .b(gate126inter6), .O(gate126inter12));
  nand2 gate1876(.a(gate126inter12), .b(gate126inter1), .O(G489));
nand2 gate127( .a(G406), .b(G407), .O(G492) );
nand2 gate128( .a(G408), .b(G409), .O(G495) );

  xor2  gate1975(.a(G411), .b(G410), .O(gate129inter0));
  nand2 gate1976(.a(gate129inter0), .b(s_204), .O(gate129inter1));
  and2  gate1977(.a(G411), .b(G410), .O(gate129inter2));
  inv1  gate1978(.a(s_204), .O(gate129inter3));
  inv1  gate1979(.a(s_205), .O(gate129inter4));
  nand2 gate1980(.a(gate129inter4), .b(gate129inter3), .O(gate129inter5));
  nor2  gate1981(.a(gate129inter5), .b(gate129inter2), .O(gate129inter6));
  inv1  gate1982(.a(G410), .O(gate129inter7));
  inv1  gate1983(.a(G411), .O(gate129inter8));
  nand2 gate1984(.a(gate129inter8), .b(gate129inter7), .O(gate129inter9));
  nand2 gate1985(.a(s_205), .b(gate129inter3), .O(gate129inter10));
  nor2  gate1986(.a(gate129inter10), .b(gate129inter9), .O(gate129inter11));
  nor2  gate1987(.a(gate129inter11), .b(gate129inter6), .O(gate129inter12));
  nand2 gate1988(.a(gate129inter12), .b(gate129inter1), .O(G498));
nand2 gate130( .a(G412), .b(G413), .O(G501) );
nand2 gate131( .a(G414), .b(G415), .O(G504) );

  xor2  gate869(.a(G417), .b(G416), .O(gate132inter0));
  nand2 gate870(.a(gate132inter0), .b(s_46), .O(gate132inter1));
  and2  gate871(.a(G417), .b(G416), .O(gate132inter2));
  inv1  gate872(.a(s_46), .O(gate132inter3));
  inv1  gate873(.a(s_47), .O(gate132inter4));
  nand2 gate874(.a(gate132inter4), .b(gate132inter3), .O(gate132inter5));
  nor2  gate875(.a(gate132inter5), .b(gate132inter2), .O(gate132inter6));
  inv1  gate876(.a(G416), .O(gate132inter7));
  inv1  gate877(.a(G417), .O(gate132inter8));
  nand2 gate878(.a(gate132inter8), .b(gate132inter7), .O(gate132inter9));
  nand2 gate879(.a(s_47), .b(gate132inter3), .O(gate132inter10));
  nor2  gate880(.a(gate132inter10), .b(gate132inter9), .O(gate132inter11));
  nor2  gate881(.a(gate132inter11), .b(gate132inter6), .O(gate132inter12));
  nand2 gate882(.a(gate132inter12), .b(gate132inter1), .O(G507));
nand2 gate133( .a(G418), .b(G419), .O(G510) );
nand2 gate134( .a(G420), .b(G421), .O(G513) );
nand2 gate135( .a(G422), .b(G423), .O(G516) );
nand2 gate136( .a(G424), .b(G425), .O(G519) );
nand2 gate137( .a(G426), .b(G429), .O(G522) );
nand2 gate138( .a(G432), .b(G435), .O(G525) );
nand2 gate139( .a(G438), .b(G441), .O(G528) );
nand2 gate140( .a(G444), .b(G447), .O(G531) );

  xor2  gate1429(.a(G453), .b(G450), .O(gate141inter0));
  nand2 gate1430(.a(gate141inter0), .b(s_126), .O(gate141inter1));
  and2  gate1431(.a(G453), .b(G450), .O(gate141inter2));
  inv1  gate1432(.a(s_126), .O(gate141inter3));
  inv1  gate1433(.a(s_127), .O(gate141inter4));
  nand2 gate1434(.a(gate141inter4), .b(gate141inter3), .O(gate141inter5));
  nor2  gate1435(.a(gate141inter5), .b(gate141inter2), .O(gate141inter6));
  inv1  gate1436(.a(G450), .O(gate141inter7));
  inv1  gate1437(.a(G453), .O(gate141inter8));
  nand2 gate1438(.a(gate141inter8), .b(gate141inter7), .O(gate141inter9));
  nand2 gate1439(.a(s_127), .b(gate141inter3), .O(gate141inter10));
  nor2  gate1440(.a(gate141inter10), .b(gate141inter9), .O(gate141inter11));
  nor2  gate1441(.a(gate141inter11), .b(gate141inter6), .O(gate141inter12));
  nand2 gate1442(.a(gate141inter12), .b(gate141inter1), .O(G534));

  xor2  gate813(.a(G459), .b(G456), .O(gate142inter0));
  nand2 gate814(.a(gate142inter0), .b(s_38), .O(gate142inter1));
  and2  gate815(.a(G459), .b(G456), .O(gate142inter2));
  inv1  gate816(.a(s_38), .O(gate142inter3));
  inv1  gate817(.a(s_39), .O(gate142inter4));
  nand2 gate818(.a(gate142inter4), .b(gate142inter3), .O(gate142inter5));
  nor2  gate819(.a(gate142inter5), .b(gate142inter2), .O(gate142inter6));
  inv1  gate820(.a(G456), .O(gate142inter7));
  inv1  gate821(.a(G459), .O(gate142inter8));
  nand2 gate822(.a(gate142inter8), .b(gate142inter7), .O(gate142inter9));
  nand2 gate823(.a(s_39), .b(gate142inter3), .O(gate142inter10));
  nor2  gate824(.a(gate142inter10), .b(gate142inter9), .O(gate142inter11));
  nor2  gate825(.a(gate142inter11), .b(gate142inter6), .O(gate142inter12));
  nand2 gate826(.a(gate142inter12), .b(gate142inter1), .O(G537));
nand2 gate143( .a(G462), .b(G465), .O(G540) );

  xor2  gate883(.a(G471), .b(G468), .O(gate144inter0));
  nand2 gate884(.a(gate144inter0), .b(s_48), .O(gate144inter1));
  and2  gate885(.a(G471), .b(G468), .O(gate144inter2));
  inv1  gate886(.a(s_48), .O(gate144inter3));
  inv1  gate887(.a(s_49), .O(gate144inter4));
  nand2 gate888(.a(gate144inter4), .b(gate144inter3), .O(gate144inter5));
  nor2  gate889(.a(gate144inter5), .b(gate144inter2), .O(gate144inter6));
  inv1  gate890(.a(G468), .O(gate144inter7));
  inv1  gate891(.a(G471), .O(gate144inter8));
  nand2 gate892(.a(gate144inter8), .b(gate144inter7), .O(gate144inter9));
  nand2 gate893(.a(s_49), .b(gate144inter3), .O(gate144inter10));
  nor2  gate894(.a(gate144inter10), .b(gate144inter9), .O(gate144inter11));
  nor2  gate895(.a(gate144inter11), .b(gate144inter6), .O(gate144inter12));
  nand2 gate896(.a(gate144inter12), .b(gate144inter1), .O(G543));

  xor2  gate1709(.a(G477), .b(G474), .O(gate145inter0));
  nand2 gate1710(.a(gate145inter0), .b(s_166), .O(gate145inter1));
  and2  gate1711(.a(G477), .b(G474), .O(gate145inter2));
  inv1  gate1712(.a(s_166), .O(gate145inter3));
  inv1  gate1713(.a(s_167), .O(gate145inter4));
  nand2 gate1714(.a(gate145inter4), .b(gate145inter3), .O(gate145inter5));
  nor2  gate1715(.a(gate145inter5), .b(gate145inter2), .O(gate145inter6));
  inv1  gate1716(.a(G474), .O(gate145inter7));
  inv1  gate1717(.a(G477), .O(gate145inter8));
  nand2 gate1718(.a(gate145inter8), .b(gate145inter7), .O(gate145inter9));
  nand2 gate1719(.a(s_167), .b(gate145inter3), .O(gate145inter10));
  nor2  gate1720(.a(gate145inter10), .b(gate145inter9), .O(gate145inter11));
  nor2  gate1721(.a(gate145inter11), .b(gate145inter6), .O(gate145inter12));
  nand2 gate1722(.a(gate145inter12), .b(gate145inter1), .O(G546));
nand2 gate146( .a(G480), .b(G483), .O(G549) );
nand2 gate147( .a(G486), .b(G489), .O(G552) );
nand2 gate148( .a(G492), .b(G495), .O(G555) );

  xor2  gate2003(.a(G501), .b(G498), .O(gate149inter0));
  nand2 gate2004(.a(gate149inter0), .b(s_208), .O(gate149inter1));
  and2  gate2005(.a(G501), .b(G498), .O(gate149inter2));
  inv1  gate2006(.a(s_208), .O(gate149inter3));
  inv1  gate2007(.a(s_209), .O(gate149inter4));
  nand2 gate2008(.a(gate149inter4), .b(gate149inter3), .O(gate149inter5));
  nor2  gate2009(.a(gate149inter5), .b(gate149inter2), .O(gate149inter6));
  inv1  gate2010(.a(G498), .O(gate149inter7));
  inv1  gate2011(.a(G501), .O(gate149inter8));
  nand2 gate2012(.a(gate149inter8), .b(gate149inter7), .O(gate149inter9));
  nand2 gate2013(.a(s_209), .b(gate149inter3), .O(gate149inter10));
  nor2  gate2014(.a(gate149inter10), .b(gate149inter9), .O(gate149inter11));
  nor2  gate2015(.a(gate149inter11), .b(gate149inter6), .O(gate149inter12));
  nand2 gate2016(.a(gate149inter12), .b(gate149inter1), .O(G558));

  xor2  gate967(.a(G507), .b(G504), .O(gate150inter0));
  nand2 gate968(.a(gate150inter0), .b(s_60), .O(gate150inter1));
  and2  gate969(.a(G507), .b(G504), .O(gate150inter2));
  inv1  gate970(.a(s_60), .O(gate150inter3));
  inv1  gate971(.a(s_61), .O(gate150inter4));
  nand2 gate972(.a(gate150inter4), .b(gate150inter3), .O(gate150inter5));
  nor2  gate973(.a(gate150inter5), .b(gate150inter2), .O(gate150inter6));
  inv1  gate974(.a(G504), .O(gate150inter7));
  inv1  gate975(.a(G507), .O(gate150inter8));
  nand2 gate976(.a(gate150inter8), .b(gate150inter7), .O(gate150inter9));
  nand2 gate977(.a(s_61), .b(gate150inter3), .O(gate150inter10));
  nor2  gate978(.a(gate150inter10), .b(gate150inter9), .O(gate150inter11));
  nor2  gate979(.a(gate150inter11), .b(gate150inter6), .O(gate150inter12));
  nand2 gate980(.a(gate150inter12), .b(gate150inter1), .O(G561));
nand2 gate151( .a(G510), .b(G513), .O(G564) );

  xor2  gate1751(.a(G519), .b(G516), .O(gate152inter0));
  nand2 gate1752(.a(gate152inter0), .b(s_172), .O(gate152inter1));
  and2  gate1753(.a(G519), .b(G516), .O(gate152inter2));
  inv1  gate1754(.a(s_172), .O(gate152inter3));
  inv1  gate1755(.a(s_173), .O(gate152inter4));
  nand2 gate1756(.a(gate152inter4), .b(gate152inter3), .O(gate152inter5));
  nor2  gate1757(.a(gate152inter5), .b(gate152inter2), .O(gate152inter6));
  inv1  gate1758(.a(G516), .O(gate152inter7));
  inv1  gate1759(.a(G519), .O(gate152inter8));
  nand2 gate1760(.a(gate152inter8), .b(gate152inter7), .O(gate152inter9));
  nand2 gate1761(.a(s_173), .b(gate152inter3), .O(gate152inter10));
  nor2  gate1762(.a(gate152inter10), .b(gate152inter9), .O(gate152inter11));
  nor2  gate1763(.a(gate152inter11), .b(gate152inter6), .O(gate152inter12));
  nand2 gate1764(.a(gate152inter12), .b(gate152inter1), .O(G567));
nand2 gate153( .a(G426), .b(G522), .O(G570) );
nand2 gate154( .a(G429), .b(G522), .O(G571) );
nand2 gate155( .a(G432), .b(G525), .O(G572) );

  xor2  gate1037(.a(G525), .b(G435), .O(gate156inter0));
  nand2 gate1038(.a(gate156inter0), .b(s_70), .O(gate156inter1));
  and2  gate1039(.a(G525), .b(G435), .O(gate156inter2));
  inv1  gate1040(.a(s_70), .O(gate156inter3));
  inv1  gate1041(.a(s_71), .O(gate156inter4));
  nand2 gate1042(.a(gate156inter4), .b(gate156inter3), .O(gate156inter5));
  nor2  gate1043(.a(gate156inter5), .b(gate156inter2), .O(gate156inter6));
  inv1  gate1044(.a(G435), .O(gate156inter7));
  inv1  gate1045(.a(G525), .O(gate156inter8));
  nand2 gate1046(.a(gate156inter8), .b(gate156inter7), .O(gate156inter9));
  nand2 gate1047(.a(s_71), .b(gate156inter3), .O(gate156inter10));
  nor2  gate1048(.a(gate156inter10), .b(gate156inter9), .O(gate156inter11));
  nor2  gate1049(.a(gate156inter11), .b(gate156inter6), .O(gate156inter12));
  nand2 gate1050(.a(gate156inter12), .b(gate156inter1), .O(G573));
nand2 gate157( .a(G438), .b(G528), .O(G574) );

  xor2  gate1205(.a(G528), .b(G441), .O(gate158inter0));
  nand2 gate1206(.a(gate158inter0), .b(s_94), .O(gate158inter1));
  and2  gate1207(.a(G528), .b(G441), .O(gate158inter2));
  inv1  gate1208(.a(s_94), .O(gate158inter3));
  inv1  gate1209(.a(s_95), .O(gate158inter4));
  nand2 gate1210(.a(gate158inter4), .b(gate158inter3), .O(gate158inter5));
  nor2  gate1211(.a(gate158inter5), .b(gate158inter2), .O(gate158inter6));
  inv1  gate1212(.a(G441), .O(gate158inter7));
  inv1  gate1213(.a(G528), .O(gate158inter8));
  nand2 gate1214(.a(gate158inter8), .b(gate158inter7), .O(gate158inter9));
  nand2 gate1215(.a(s_95), .b(gate158inter3), .O(gate158inter10));
  nor2  gate1216(.a(gate158inter10), .b(gate158inter9), .O(gate158inter11));
  nor2  gate1217(.a(gate158inter11), .b(gate158inter6), .O(gate158inter12));
  nand2 gate1218(.a(gate158inter12), .b(gate158inter1), .O(G575));

  xor2  gate631(.a(G531), .b(G444), .O(gate159inter0));
  nand2 gate632(.a(gate159inter0), .b(s_12), .O(gate159inter1));
  and2  gate633(.a(G531), .b(G444), .O(gate159inter2));
  inv1  gate634(.a(s_12), .O(gate159inter3));
  inv1  gate635(.a(s_13), .O(gate159inter4));
  nand2 gate636(.a(gate159inter4), .b(gate159inter3), .O(gate159inter5));
  nor2  gate637(.a(gate159inter5), .b(gate159inter2), .O(gate159inter6));
  inv1  gate638(.a(G444), .O(gate159inter7));
  inv1  gate639(.a(G531), .O(gate159inter8));
  nand2 gate640(.a(gate159inter8), .b(gate159inter7), .O(gate159inter9));
  nand2 gate641(.a(s_13), .b(gate159inter3), .O(gate159inter10));
  nor2  gate642(.a(gate159inter10), .b(gate159inter9), .O(gate159inter11));
  nor2  gate643(.a(gate159inter11), .b(gate159inter6), .O(gate159inter12));
  nand2 gate644(.a(gate159inter12), .b(gate159inter1), .O(G576));

  xor2  gate981(.a(G531), .b(G447), .O(gate160inter0));
  nand2 gate982(.a(gate160inter0), .b(s_62), .O(gate160inter1));
  and2  gate983(.a(G531), .b(G447), .O(gate160inter2));
  inv1  gate984(.a(s_62), .O(gate160inter3));
  inv1  gate985(.a(s_63), .O(gate160inter4));
  nand2 gate986(.a(gate160inter4), .b(gate160inter3), .O(gate160inter5));
  nor2  gate987(.a(gate160inter5), .b(gate160inter2), .O(gate160inter6));
  inv1  gate988(.a(G447), .O(gate160inter7));
  inv1  gate989(.a(G531), .O(gate160inter8));
  nand2 gate990(.a(gate160inter8), .b(gate160inter7), .O(gate160inter9));
  nand2 gate991(.a(s_63), .b(gate160inter3), .O(gate160inter10));
  nor2  gate992(.a(gate160inter10), .b(gate160inter9), .O(gate160inter11));
  nor2  gate993(.a(gate160inter11), .b(gate160inter6), .O(gate160inter12));
  nand2 gate994(.a(gate160inter12), .b(gate160inter1), .O(G577));
nand2 gate161( .a(G450), .b(G534), .O(G578) );

  xor2  gate2087(.a(G534), .b(G453), .O(gate162inter0));
  nand2 gate2088(.a(gate162inter0), .b(s_220), .O(gate162inter1));
  and2  gate2089(.a(G534), .b(G453), .O(gate162inter2));
  inv1  gate2090(.a(s_220), .O(gate162inter3));
  inv1  gate2091(.a(s_221), .O(gate162inter4));
  nand2 gate2092(.a(gate162inter4), .b(gate162inter3), .O(gate162inter5));
  nor2  gate2093(.a(gate162inter5), .b(gate162inter2), .O(gate162inter6));
  inv1  gate2094(.a(G453), .O(gate162inter7));
  inv1  gate2095(.a(G534), .O(gate162inter8));
  nand2 gate2096(.a(gate162inter8), .b(gate162inter7), .O(gate162inter9));
  nand2 gate2097(.a(s_221), .b(gate162inter3), .O(gate162inter10));
  nor2  gate2098(.a(gate162inter10), .b(gate162inter9), .O(gate162inter11));
  nor2  gate2099(.a(gate162inter11), .b(gate162inter6), .O(gate162inter12));
  nand2 gate2100(.a(gate162inter12), .b(gate162inter1), .O(G579));
nand2 gate163( .a(G456), .b(G537), .O(G580) );

  xor2  gate729(.a(G537), .b(G459), .O(gate164inter0));
  nand2 gate730(.a(gate164inter0), .b(s_26), .O(gate164inter1));
  and2  gate731(.a(G537), .b(G459), .O(gate164inter2));
  inv1  gate732(.a(s_26), .O(gate164inter3));
  inv1  gate733(.a(s_27), .O(gate164inter4));
  nand2 gate734(.a(gate164inter4), .b(gate164inter3), .O(gate164inter5));
  nor2  gate735(.a(gate164inter5), .b(gate164inter2), .O(gate164inter6));
  inv1  gate736(.a(G459), .O(gate164inter7));
  inv1  gate737(.a(G537), .O(gate164inter8));
  nand2 gate738(.a(gate164inter8), .b(gate164inter7), .O(gate164inter9));
  nand2 gate739(.a(s_27), .b(gate164inter3), .O(gate164inter10));
  nor2  gate740(.a(gate164inter10), .b(gate164inter9), .O(gate164inter11));
  nor2  gate741(.a(gate164inter11), .b(gate164inter6), .O(gate164inter12));
  nand2 gate742(.a(gate164inter12), .b(gate164inter1), .O(G581));
nand2 gate165( .a(G462), .b(G540), .O(G582) );
nand2 gate166( .a(G465), .b(G540), .O(G583) );
nand2 gate167( .a(G468), .b(G543), .O(G584) );
nand2 gate168( .a(G471), .b(G543), .O(G585) );
nand2 gate169( .a(G474), .b(G546), .O(G586) );
nand2 gate170( .a(G477), .b(G546), .O(G587) );
nand2 gate171( .a(G480), .b(G549), .O(G588) );
nand2 gate172( .a(G483), .b(G549), .O(G589) );
nand2 gate173( .a(G486), .b(G552), .O(G590) );
nand2 gate174( .a(G489), .b(G552), .O(G591) );
nand2 gate175( .a(G492), .b(G555), .O(G592) );
nand2 gate176( .a(G495), .b(G555), .O(G593) );
nand2 gate177( .a(G498), .b(G558), .O(G594) );

  xor2  gate1667(.a(G558), .b(G501), .O(gate178inter0));
  nand2 gate1668(.a(gate178inter0), .b(s_160), .O(gate178inter1));
  and2  gate1669(.a(G558), .b(G501), .O(gate178inter2));
  inv1  gate1670(.a(s_160), .O(gate178inter3));
  inv1  gate1671(.a(s_161), .O(gate178inter4));
  nand2 gate1672(.a(gate178inter4), .b(gate178inter3), .O(gate178inter5));
  nor2  gate1673(.a(gate178inter5), .b(gate178inter2), .O(gate178inter6));
  inv1  gate1674(.a(G501), .O(gate178inter7));
  inv1  gate1675(.a(G558), .O(gate178inter8));
  nand2 gate1676(.a(gate178inter8), .b(gate178inter7), .O(gate178inter9));
  nand2 gate1677(.a(s_161), .b(gate178inter3), .O(gate178inter10));
  nor2  gate1678(.a(gate178inter10), .b(gate178inter9), .O(gate178inter11));
  nor2  gate1679(.a(gate178inter11), .b(gate178inter6), .O(gate178inter12));
  nand2 gate1680(.a(gate178inter12), .b(gate178inter1), .O(G595));

  xor2  gate1233(.a(G561), .b(G504), .O(gate179inter0));
  nand2 gate1234(.a(gate179inter0), .b(s_98), .O(gate179inter1));
  and2  gate1235(.a(G561), .b(G504), .O(gate179inter2));
  inv1  gate1236(.a(s_98), .O(gate179inter3));
  inv1  gate1237(.a(s_99), .O(gate179inter4));
  nand2 gate1238(.a(gate179inter4), .b(gate179inter3), .O(gate179inter5));
  nor2  gate1239(.a(gate179inter5), .b(gate179inter2), .O(gate179inter6));
  inv1  gate1240(.a(G504), .O(gate179inter7));
  inv1  gate1241(.a(G561), .O(gate179inter8));
  nand2 gate1242(.a(gate179inter8), .b(gate179inter7), .O(gate179inter9));
  nand2 gate1243(.a(s_99), .b(gate179inter3), .O(gate179inter10));
  nor2  gate1244(.a(gate179inter10), .b(gate179inter9), .O(gate179inter11));
  nor2  gate1245(.a(gate179inter11), .b(gate179inter6), .O(gate179inter12));
  nand2 gate1246(.a(gate179inter12), .b(gate179inter1), .O(G596));
nand2 gate180( .a(G507), .b(G561), .O(G597) );
nand2 gate181( .a(G510), .b(G564), .O(G598) );

  xor2  gate1891(.a(G564), .b(G513), .O(gate182inter0));
  nand2 gate1892(.a(gate182inter0), .b(s_192), .O(gate182inter1));
  and2  gate1893(.a(G564), .b(G513), .O(gate182inter2));
  inv1  gate1894(.a(s_192), .O(gate182inter3));
  inv1  gate1895(.a(s_193), .O(gate182inter4));
  nand2 gate1896(.a(gate182inter4), .b(gate182inter3), .O(gate182inter5));
  nor2  gate1897(.a(gate182inter5), .b(gate182inter2), .O(gate182inter6));
  inv1  gate1898(.a(G513), .O(gate182inter7));
  inv1  gate1899(.a(G564), .O(gate182inter8));
  nand2 gate1900(.a(gate182inter8), .b(gate182inter7), .O(gate182inter9));
  nand2 gate1901(.a(s_193), .b(gate182inter3), .O(gate182inter10));
  nor2  gate1902(.a(gate182inter10), .b(gate182inter9), .O(gate182inter11));
  nor2  gate1903(.a(gate182inter11), .b(gate182inter6), .O(gate182inter12));
  nand2 gate1904(.a(gate182inter12), .b(gate182inter1), .O(G599));
nand2 gate183( .a(G516), .b(G567), .O(G600) );
nand2 gate184( .a(G519), .b(G567), .O(G601) );
nand2 gate185( .a(G570), .b(G571), .O(G602) );

  xor2  gate617(.a(G573), .b(G572), .O(gate186inter0));
  nand2 gate618(.a(gate186inter0), .b(s_10), .O(gate186inter1));
  and2  gate619(.a(G573), .b(G572), .O(gate186inter2));
  inv1  gate620(.a(s_10), .O(gate186inter3));
  inv1  gate621(.a(s_11), .O(gate186inter4));
  nand2 gate622(.a(gate186inter4), .b(gate186inter3), .O(gate186inter5));
  nor2  gate623(.a(gate186inter5), .b(gate186inter2), .O(gate186inter6));
  inv1  gate624(.a(G572), .O(gate186inter7));
  inv1  gate625(.a(G573), .O(gate186inter8));
  nand2 gate626(.a(gate186inter8), .b(gate186inter7), .O(gate186inter9));
  nand2 gate627(.a(s_11), .b(gate186inter3), .O(gate186inter10));
  nor2  gate628(.a(gate186inter10), .b(gate186inter9), .O(gate186inter11));
  nor2  gate629(.a(gate186inter11), .b(gate186inter6), .O(gate186inter12));
  nand2 gate630(.a(gate186inter12), .b(gate186inter1), .O(G607));
nand2 gate187( .a(G574), .b(G575), .O(G612) );
nand2 gate188( .a(G576), .b(G577), .O(G617) );
nand2 gate189( .a(G578), .b(G579), .O(G622) );
nand2 gate190( .a(G580), .b(G581), .O(G627) );
nand2 gate191( .a(G582), .b(G583), .O(G632) );
nand2 gate192( .a(G584), .b(G585), .O(G637) );
nand2 gate193( .a(G586), .b(G587), .O(G642) );
nand2 gate194( .a(G588), .b(G589), .O(G645) );
nand2 gate195( .a(G590), .b(G591), .O(G648) );
nand2 gate196( .a(G592), .b(G593), .O(G651) );
nand2 gate197( .a(G594), .b(G595), .O(G654) );
nand2 gate198( .a(G596), .b(G597), .O(G657) );

  xor2  gate1849(.a(G599), .b(G598), .O(gate199inter0));
  nand2 gate1850(.a(gate199inter0), .b(s_186), .O(gate199inter1));
  and2  gate1851(.a(G599), .b(G598), .O(gate199inter2));
  inv1  gate1852(.a(s_186), .O(gate199inter3));
  inv1  gate1853(.a(s_187), .O(gate199inter4));
  nand2 gate1854(.a(gate199inter4), .b(gate199inter3), .O(gate199inter5));
  nor2  gate1855(.a(gate199inter5), .b(gate199inter2), .O(gate199inter6));
  inv1  gate1856(.a(G598), .O(gate199inter7));
  inv1  gate1857(.a(G599), .O(gate199inter8));
  nand2 gate1858(.a(gate199inter8), .b(gate199inter7), .O(gate199inter9));
  nand2 gate1859(.a(s_187), .b(gate199inter3), .O(gate199inter10));
  nor2  gate1860(.a(gate199inter10), .b(gate199inter9), .O(gate199inter11));
  nor2  gate1861(.a(gate199inter11), .b(gate199inter6), .O(gate199inter12));
  nand2 gate1862(.a(gate199inter12), .b(gate199inter1), .O(G660));
nand2 gate200( .a(G600), .b(G601), .O(G663) );
nand2 gate201( .a(G602), .b(G607), .O(G666) );
nand2 gate202( .a(G612), .b(G617), .O(G669) );

  xor2  gate1989(.a(G612), .b(G602), .O(gate203inter0));
  nand2 gate1990(.a(gate203inter0), .b(s_206), .O(gate203inter1));
  and2  gate1991(.a(G612), .b(G602), .O(gate203inter2));
  inv1  gate1992(.a(s_206), .O(gate203inter3));
  inv1  gate1993(.a(s_207), .O(gate203inter4));
  nand2 gate1994(.a(gate203inter4), .b(gate203inter3), .O(gate203inter5));
  nor2  gate1995(.a(gate203inter5), .b(gate203inter2), .O(gate203inter6));
  inv1  gate1996(.a(G602), .O(gate203inter7));
  inv1  gate1997(.a(G612), .O(gate203inter8));
  nand2 gate1998(.a(gate203inter8), .b(gate203inter7), .O(gate203inter9));
  nand2 gate1999(.a(s_207), .b(gate203inter3), .O(gate203inter10));
  nor2  gate2000(.a(gate203inter10), .b(gate203inter9), .O(gate203inter11));
  nor2  gate2001(.a(gate203inter11), .b(gate203inter6), .O(gate203inter12));
  nand2 gate2002(.a(gate203inter12), .b(gate203inter1), .O(G672));
nand2 gate204( .a(G607), .b(G617), .O(G675) );

  xor2  gate603(.a(G627), .b(G622), .O(gate205inter0));
  nand2 gate604(.a(gate205inter0), .b(s_8), .O(gate205inter1));
  and2  gate605(.a(G627), .b(G622), .O(gate205inter2));
  inv1  gate606(.a(s_8), .O(gate205inter3));
  inv1  gate607(.a(s_9), .O(gate205inter4));
  nand2 gate608(.a(gate205inter4), .b(gate205inter3), .O(gate205inter5));
  nor2  gate609(.a(gate205inter5), .b(gate205inter2), .O(gate205inter6));
  inv1  gate610(.a(G622), .O(gate205inter7));
  inv1  gate611(.a(G627), .O(gate205inter8));
  nand2 gate612(.a(gate205inter8), .b(gate205inter7), .O(gate205inter9));
  nand2 gate613(.a(s_9), .b(gate205inter3), .O(gate205inter10));
  nor2  gate614(.a(gate205inter10), .b(gate205inter9), .O(gate205inter11));
  nor2  gate615(.a(gate205inter11), .b(gate205inter6), .O(gate205inter12));
  nand2 gate616(.a(gate205inter12), .b(gate205inter1), .O(G678));
nand2 gate206( .a(G632), .b(G637), .O(G681) );
nand2 gate207( .a(G622), .b(G632), .O(G684) );
nand2 gate208( .a(G627), .b(G637), .O(G687) );

  xor2  gate911(.a(G666), .b(G602), .O(gate209inter0));
  nand2 gate912(.a(gate209inter0), .b(s_52), .O(gate209inter1));
  and2  gate913(.a(G666), .b(G602), .O(gate209inter2));
  inv1  gate914(.a(s_52), .O(gate209inter3));
  inv1  gate915(.a(s_53), .O(gate209inter4));
  nand2 gate916(.a(gate209inter4), .b(gate209inter3), .O(gate209inter5));
  nor2  gate917(.a(gate209inter5), .b(gate209inter2), .O(gate209inter6));
  inv1  gate918(.a(G602), .O(gate209inter7));
  inv1  gate919(.a(G666), .O(gate209inter8));
  nand2 gate920(.a(gate209inter8), .b(gate209inter7), .O(gate209inter9));
  nand2 gate921(.a(s_53), .b(gate209inter3), .O(gate209inter10));
  nor2  gate922(.a(gate209inter10), .b(gate209inter9), .O(gate209inter11));
  nor2  gate923(.a(gate209inter11), .b(gate209inter6), .O(gate209inter12));
  nand2 gate924(.a(gate209inter12), .b(gate209inter1), .O(G690));
nand2 gate210( .a(G607), .b(G666), .O(G691) );

  xor2  gate2073(.a(G669), .b(G612), .O(gate211inter0));
  nand2 gate2074(.a(gate211inter0), .b(s_218), .O(gate211inter1));
  and2  gate2075(.a(G669), .b(G612), .O(gate211inter2));
  inv1  gate2076(.a(s_218), .O(gate211inter3));
  inv1  gate2077(.a(s_219), .O(gate211inter4));
  nand2 gate2078(.a(gate211inter4), .b(gate211inter3), .O(gate211inter5));
  nor2  gate2079(.a(gate211inter5), .b(gate211inter2), .O(gate211inter6));
  inv1  gate2080(.a(G612), .O(gate211inter7));
  inv1  gate2081(.a(G669), .O(gate211inter8));
  nand2 gate2082(.a(gate211inter8), .b(gate211inter7), .O(gate211inter9));
  nand2 gate2083(.a(s_219), .b(gate211inter3), .O(gate211inter10));
  nor2  gate2084(.a(gate211inter10), .b(gate211inter9), .O(gate211inter11));
  nor2  gate2085(.a(gate211inter11), .b(gate211inter6), .O(gate211inter12));
  nand2 gate2086(.a(gate211inter12), .b(gate211inter1), .O(G692));

  xor2  gate1009(.a(G669), .b(G617), .O(gate212inter0));
  nand2 gate1010(.a(gate212inter0), .b(s_66), .O(gate212inter1));
  and2  gate1011(.a(G669), .b(G617), .O(gate212inter2));
  inv1  gate1012(.a(s_66), .O(gate212inter3));
  inv1  gate1013(.a(s_67), .O(gate212inter4));
  nand2 gate1014(.a(gate212inter4), .b(gate212inter3), .O(gate212inter5));
  nor2  gate1015(.a(gate212inter5), .b(gate212inter2), .O(gate212inter6));
  inv1  gate1016(.a(G617), .O(gate212inter7));
  inv1  gate1017(.a(G669), .O(gate212inter8));
  nand2 gate1018(.a(gate212inter8), .b(gate212inter7), .O(gate212inter9));
  nand2 gate1019(.a(s_67), .b(gate212inter3), .O(gate212inter10));
  nor2  gate1020(.a(gate212inter10), .b(gate212inter9), .O(gate212inter11));
  nor2  gate1021(.a(gate212inter11), .b(gate212inter6), .O(gate212inter12));
  nand2 gate1022(.a(gate212inter12), .b(gate212inter1), .O(G693));
nand2 gate213( .a(G602), .b(G672), .O(G694) );
nand2 gate214( .a(G612), .b(G672), .O(G695) );
nand2 gate215( .a(G607), .b(G675), .O(G696) );
nand2 gate216( .a(G617), .b(G675), .O(G697) );

  xor2  gate1317(.a(G678), .b(G622), .O(gate217inter0));
  nand2 gate1318(.a(gate217inter0), .b(s_110), .O(gate217inter1));
  and2  gate1319(.a(G678), .b(G622), .O(gate217inter2));
  inv1  gate1320(.a(s_110), .O(gate217inter3));
  inv1  gate1321(.a(s_111), .O(gate217inter4));
  nand2 gate1322(.a(gate217inter4), .b(gate217inter3), .O(gate217inter5));
  nor2  gate1323(.a(gate217inter5), .b(gate217inter2), .O(gate217inter6));
  inv1  gate1324(.a(G622), .O(gate217inter7));
  inv1  gate1325(.a(G678), .O(gate217inter8));
  nand2 gate1326(.a(gate217inter8), .b(gate217inter7), .O(gate217inter9));
  nand2 gate1327(.a(s_111), .b(gate217inter3), .O(gate217inter10));
  nor2  gate1328(.a(gate217inter10), .b(gate217inter9), .O(gate217inter11));
  nor2  gate1329(.a(gate217inter11), .b(gate217inter6), .O(gate217inter12));
  nand2 gate1330(.a(gate217inter12), .b(gate217inter1), .O(G698));
nand2 gate218( .a(G627), .b(G678), .O(G699) );
nand2 gate219( .a(G632), .b(G681), .O(G700) );
nand2 gate220( .a(G637), .b(G681), .O(G701) );
nand2 gate221( .a(G622), .b(G684), .O(G702) );
nand2 gate222( .a(G632), .b(G684), .O(G703) );

  xor2  gate1401(.a(G687), .b(G627), .O(gate223inter0));
  nand2 gate1402(.a(gate223inter0), .b(s_122), .O(gate223inter1));
  and2  gate1403(.a(G687), .b(G627), .O(gate223inter2));
  inv1  gate1404(.a(s_122), .O(gate223inter3));
  inv1  gate1405(.a(s_123), .O(gate223inter4));
  nand2 gate1406(.a(gate223inter4), .b(gate223inter3), .O(gate223inter5));
  nor2  gate1407(.a(gate223inter5), .b(gate223inter2), .O(gate223inter6));
  inv1  gate1408(.a(G627), .O(gate223inter7));
  inv1  gate1409(.a(G687), .O(gate223inter8));
  nand2 gate1410(.a(gate223inter8), .b(gate223inter7), .O(gate223inter9));
  nand2 gate1411(.a(s_123), .b(gate223inter3), .O(gate223inter10));
  nor2  gate1412(.a(gate223inter10), .b(gate223inter9), .O(gate223inter11));
  nor2  gate1413(.a(gate223inter11), .b(gate223inter6), .O(gate223inter12));
  nand2 gate1414(.a(gate223inter12), .b(gate223inter1), .O(G704));
nand2 gate224( .a(G637), .b(G687), .O(G705) );

  xor2  gate1247(.a(G691), .b(G690), .O(gate225inter0));
  nand2 gate1248(.a(gate225inter0), .b(s_100), .O(gate225inter1));
  and2  gate1249(.a(G691), .b(G690), .O(gate225inter2));
  inv1  gate1250(.a(s_100), .O(gate225inter3));
  inv1  gate1251(.a(s_101), .O(gate225inter4));
  nand2 gate1252(.a(gate225inter4), .b(gate225inter3), .O(gate225inter5));
  nor2  gate1253(.a(gate225inter5), .b(gate225inter2), .O(gate225inter6));
  inv1  gate1254(.a(G690), .O(gate225inter7));
  inv1  gate1255(.a(G691), .O(gate225inter8));
  nand2 gate1256(.a(gate225inter8), .b(gate225inter7), .O(gate225inter9));
  nand2 gate1257(.a(s_101), .b(gate225inter3), .O(gate225inter10));
  nor2  gate1258(.a(gate225inter10), .b(gate225inter9), .O(gate225inter11));
  nor2  gate1259(.a(gate225inter11), .b(gate225inter6), .O(gate225inter12));
  nand2 gate1260(.a(gate225inter12), .b(gate225inter1), .O(G706));
nand2 gate226( .a(G692), .b(G693), .O(G709) );
nand2 gate227( .a(G694), .b(G695), .O(G712) );
nand2 gate228( .a(G696), .b(G697), .O(G715) );
nand2 gate229( .a(G698), .b(G699), .O(G718) );

  xor2  gate757(.a(G701), .b(G700), .O(gate230inter0));
  nand2 gate758(.a(gate230inter0), .b(s_30), .O(gate230inter1));
  and2  gate759(.a(G701), .b(G700), .O(gate230inter2));
  inv1  gate760(.a(s_30), .O(gate230inter3));
  inv1  gate761(.a(s_31), .O(gate230inter4));
  nand2 gate762(.a(gate230inter4), .b(gate230inter3), .O(gate230inter5));
  nor2  gate763(.a(gate230inter5), .b(gate230inter2), .O(gate230inter6));
  inv1  gate764(.a(G700), .O(gate230inter7));
  inv1  gate765(.a(G701), .O(gate230inter8));
  nand2 gate766(.a(gate230inter8), .b(gate230inter7), .O(gate230inter9));
  nand2 gate767(.a(s_31), .b(gate230inter3), .O(gate230inter10));
  nor2  gate768(.a(gate230inter10), .b(gate230inter9), .O(gate230inter11));
  nor2  gate769(.a(gate230inter11), .b(gate230inter6), .O(gate230inter12));
  nand2 gate770(.a(gate230inter12), .b(gate230inter1), .O(G721));
nand2 gate231( .a(G702), .b(G703), .O(G724) );
nand2 gate232( .a(G704), .b(G705), .O(G727) );

  xor2  gate1723(.a(G718), .b(G242), .O(gate233inter0));
  nand2 gate1724(.a(gate233inter0), .b(s_168), .O(gate233inter1));
  and2  gate1725(.a(G718), .b(G242), .O(gate233inter2));
  inv1  gate1726(.a(s_168), .O(gate233inter3));
  inv1  gate1727(.a(s_169), .O(gate233inter4));
  nand2 gate1728(.a(gate233inter4), .b(gate233inter3), .O(gate233inter5));
  nor2  gate1729(.a(gate233inter5), .b(gate233inter2), .O(gate233inter6));
  inv1  gate1730(.a(G242), .O(gate233inter7));
  inv1  gate1731(.a(G718), .O(gate233inter8));
  nand2 gate1732(.a(gate233inter8), .b(gate233inter7), .O(gate233inter9));
  nand2 gate1733(.a(s_169), .b(gate233inter3), .O(gate233inter10));
  nor2  gate1734(.a(gate233inter10), .b(gate233inter9), .O(gate233inter11));
  nor2  gate1735(.a(gate233inter11), .b(gate233inter6), .O(gate233inter12));
  nand2 gate1736(.a(gate233inter12), .b(gate233inter1), .O(G730));
nand2 gate234( .a(G245), .b(G721), .O(G733) );
nand2 gate235( .a(G248), .b(G724), .O(G736) );
nand2 gate236( .a(G251), .b(G727), .O(G739) );
nand2 gate237( .a(G254), .b(G706), .O(G742) );
nand2 gate238( .a(G257), .b(G709), .O(G745) );

  xor2  gate1135(.a(G712), .b(G260), .O(gate239inter0));
  nand2 gate1136(.a(gate239inter0), .b(s_84), .O(gate239inter1));
  and2  gate1137(.a(G712), .b(G260), .O(gate239inter2));
  inv1  gate1138(.a(s_84), .O(gate239inter3));
  inv1  gate1139(.a(s_85), .O(gate239inter4));
  nand2 gate1140(.a(gate239inter4), .b(gate239inter3), .O(gate239inter5));
  nor2  gate1141(.a(gate239inter5), .b(gate239inter2), .O(gate239inter6));
  inv1  gate1142(.a(G260), .O(gate239inter7));
  inv1  gate1143(.a(G712), .O(gate239inter8));
  nand2 gate1144(.a(gate239inter8), .b(gate239inter7), .O(gate239inter9));
  nand2 gate1145(.a(s_85), .b(gate239inter3), .O(gate239inter10));
  nor2  gate1146(.a(gate239inter10), .b(gate239inter9), .O(gate239inter11));
  nor2  gate1147(.a(gate239inter11), .b(gate239inter6), .O(gate239inter12));
  nand2 gate1148(.a(gate239inter12), .b(gate239inter1), .O(G748));

  xor2  gate687(.a(G715), .b(G263), .O(gate240inter0));
  nand2 gate688(.a(gate240inter0), .b(s_20), .O(gate240inter1));
  and2  gate689(.a(G715), .b(G263), .O(gate240inter2));
  inv1  gate690(.a(s_20), .O(gate240inter3));
  inv1  gate691(.a(s_21), .O(gate240inter4));
  nand2 gate692(.a(gate240inter4), .b(gate240inter3), .O(gate240inter5));
  nor2  gate693(.a(gate240inter5), .b(gate240inter2), .O(gate240inter6));
  inv1  gate694(.a(G263), .O(gate240inter7));
  inv1  gate695(.a(G715), .O(gate240inter8));
  nand2 gate696(.a(gate240inter8), .b(gate240inter7), .O(gate240inter9));
  nand2 gate697(.a(s_21), .b(gate240inter3), .O(gate240inter10));
  nor2  gate698(.a(gate240inter10), .b(gate240inter9), .O(gate240inter11));
  nor2  gate699(.a(gate240inter11), .b(gate240inter6), .O(gate240inter12));
  nand2 gate700(.a(gate240inter12), .b(gate240inter1), .O(G751));

  xor2  gate659(.a(G730), .b(G242), .O(gate241inter0));
  nand2 gate660(.a(gate241inter0), .b(s_16), .O(gate241inter1));
  and2  gate661(.a(G730), .b(G242), .O(gate241inter2));
  inv1  gate662(.a(s_16), .O(gate241inter3));
  inv1  gate663(.a(s_17), .O(gate241inter4));
  nand2 gate664(.a(gate241inter4), .b(gate241inter3), .O(gate241inter5));
  nor2  gate665(.a(gate241inter5), .b(gate241inter2), .O(gate241inter6));
  inv1  gate666(.a(G242), .O(gate241inter7));
  inv1  gate667(.a(G730), .O(gate241inter8));
  nand2 gate668(.a(gate241inter8), .b(gate241inter7), .O(gate241inter9));
  nand2 gate669(.a(s_17), .b(gate241inter3), .O(gate241inter10));
  nor2  gate670(.a(gate241inter10), .b(gate241inter9), .O(gate241inter11));
  nor2  gate671(.a(gate241inter11), .b(gate241inter6), .O(gate241inter12));
  nand2 gate672(.a(gate241inter12), .b(gate241inter1), .O(G754));
nand2 gate242( .a(G718), .b(G730), .O(G755) );

  xor2  gate1765(.a(G733), .b(G245), .O(gate243inter0));
  nand2 gate1766(.a(gate243inter0), .b(s_174), .O(gate243inter1));
  and2  gate1767(.a(G733), .b(G245), .O(gate243inter2));
  inv1  gate1768(.a(s_174), .O(gate243inter3));
  inv1  gate1769(.a(s_175), .O(gate243inter4));
  nand2 gate1770(.a(gate243inter4), .b(gate243inter3), .O(gate243inter5));
  nor2  gate1771(.a(gate243inter5), .b(gate243inter2), .O(gate243inter6));
  inv1  gate1772(.a(G245), .O(gate243inter7));
  inv1  gate1773(.a(G733), .O(gate243inter8));
  nand2 gate1774(.a(gate243inter8), .b(gate243inter7), .O(gate243inter9));
  nand2 gate1775(.a(s_175), .b(gate243inter3), .O(gate243inter10));
  nor2  gate1776(.a(gate243inter10), .b(gate243inter9), .O(gate243inter11));
  nor2  gate1777(.a(gate243inter11), .b(gate243inter6), .O(gate243inter12));
  nand2 gate1778(.a(gate243inter12), .b(gate243inter1), .O(G756));

  xor2  gate1947(.a(G733), .b(G721), .O(gate244inter0));
  nand2 gate1948(.a(gate244inter0), .b(s_200), .O(gate244inter1));
  and2  gate1949(.a(G733), .b(G721), .O(gate244inter2));
  inv1  gate1950(.a(s_200), .O(gate244inter3));
  inv1  gate1951(.a(s_201), .O(gate244inter4));
  nand2 gate1952(.a(gate244inter4), .b(gate244inter3), .O(gate244inter5));
  nor2  gate1953(.a(gate244inter5), .b(gate244inter2), .O(gate244inter6));
  inv1  gate1954(.a(G721), .O(gate244inter7));
  inv1  gate1955(.a(G733), .O(gate244inter8));
  nand2 gate1956(.a(gate244inter8), .b(gate244inter7), .O(gate244inter9));
  nand2 gate1957(.a(s_201), .b(gate244inter3), .O(gate244inter10));
  nor2  gate1958(.a(gate244inter10), .b(gate244inter9), .O(gate244inter11));
  nor2  gate1959(.a(gate244inter11), .b(gate244inter6), .O(gate244inter12));
  nand2 gate1960(.a(gate244inter12), .b(gate244inter1), .O(G757));
nand2 gate245( .a(G248), .b(G736), .O(G758) );
nand2 gate246( .a(G724), .b(G736), .O(G759) );
nand2 gate247( .a(G251), .b(G739), .O(G760) );
nand2 gate248( .a(G727), .b(G739), .O(G761) );
nand2 gate249( .a(G254), .b(G742), .O(G762) );
nand2 gate250( .a(G706), .b(G742), .O(G763) );
nand2 gate251( .a(G257), .b(G745), .O(G764) );
nand2 gate252( .a(G709), .b(G745), .O(G765) );
nand2 gate253( .a(G260), .b(G748), .O(G766) );
nand2 gate254( .a(G712), .b(G748), .O(G767) );

  xor2  gate1877(.a(G751), .b(G263), .O(gate255inter0));
  nand2 gate1878(.a(gate255inter0), .b(s_190), .O(gate255inter1));
  and2  gate1879(.a(G751), .b(G263), .O(gate255inter2));
  inv1  gate1880(.a(s_190), .O(gate255inter3));
  inv1  gate1881(.a(s_191), .O(gate255inter4));
  nand2 gate1882(.a(gate255inter4), .b(gate255inter3), .O(gate255inter5));
  nor2  gate1883(.a(gate255inter5), .b(gate255inter2), .O(gate255inter6));
  inv1  gate1884(.a(G263), .O(gate255inter7));
  inv1  gate1885(.a(G751), .O(gate255inter8));
  nand2 gate1886(.a(gate255inter8), .b(gate255inter7), .O(gate255inter9));
  nand2 gate1887(.a(s_191), .b(gate255inter3), .O(gate255inter10));
  nor2  gate1888(.a(gate255inter10), .b(gate255inter9), .O(gate255inter11));
  nor2  gate1889(.a(gate255inter11), .b(gate255inter6), .O(gate255inter12));
  nand2 gate1890(.a(gate255inter12), .b(gate255inter1), .O(G768));
nand2 gate256( .a(G715), .b(G751), .O(G769) );
nand2 gate257( .a(G754), .b(G755), .O(G770) );
nand2 gate258( .a(G756), .b(G757), .O(G773) );
nand2 gate259( .a(G758), .b(G759), .O(G776) );

  xor2  gate1163(.a(G761), .b(G760), .O(gate260inter0));
  nand2 gate1164(.a(gate260inter0), .b(s_88), .O(gate260inter1));
  and2  gate1165(.a(G761), .b(G760), .O(gate260inter2));
  inv1  gate1166(.a(s_88), .O(gate260inter3));
  inv1  gate1167(.a(s_89), .O(gate260inter4));
  nand2 gate1168(.a(gate260inter4), .b(gate260inter3), .O(gate260inter5));
  nor2  gate1169(.a(gate260inter5), .b(gate260inter2), .O(gate260inter6));
  inv1  gate1170(.a(G760), .O(gate260inter7));
  inv1  gate1171(.a(G761), .O(gate260inter8));
  nand2 gate1172(.a(gate260inter8), .b(gate260inter7), .O(gate260inter9));
  nand2 gate1173(.a(s_89), .b(gate260inter3), .O(gate260inter10));
  nor2  gate1174(.a(gate260inter10), .b(gate260inter9), .O(gate260inter11));
  nor2  gate1175(.a(gate260inter11), .b(gate260inter6), .O(gate260inter12));
  nand2 gate1176(.a(gate260inter12), .b(gate260inter1), .O(G779));
nand2 gate261( .a(G762), .b(G763), .O(G782) );
nand2 gate262( .a(G764), .b(G765), .O(G785) );
nand2 gate263( .a(G766), .b(G767), .O(G788) );

  xor2  gate701(.a(G769), .b(G768), .O(gate264inter0));
  nand2 gate702(.a(gate264inter0), .b(s_22), .O(gate264inter1));
  and2  gate703(.a(G769), .b(G768), .O(gate264inter2));
  inv1  gate704(.a(s_22), .O(gate264inter3));
  inv1  gate705(.a(s_23), .O(gate264inter4));
  nand2 gate706(.a(gate264inter4), .b(gate264inter3), .O(gate264inter5));
  nor2  gate707(.a(gate264inter5), .b(gate264inter2), .O(gate264inter6));
  inv1  gate708(.a(G768), .O(gate264inter7));
  inv1  gate709(.a(G769), .O(gate264inter8));
  nand2 gate710(.a(gate264inter8), .b(gate264inter7), .O(gate264inter9));
  nand2 gate711(.a(s_23), .b(gate264inter3), .O(gate264inter10));
  nor2  gate712(.a(gate264inter10), .b(gate264inter9), .O(gate264inter11));
  nor2  gate713(.a(gate264inter11), .b(gate264inter6), .O(gate264inter12));
  nand2 gate714(.a(gate264inter12), .b(gate264inter1), .O(G791));

  xor2  gate1093(.a(G770), .b(G642), .O(gate265inter0));
  nand2 gate1094(.a(gate265inter0), .b(s_78), .O(gate265inter1));
  and2  gate1095(.a(G770), .b(G642), .O(gate265inter2));
  inv1  gate1096(.a(s_78), .O(gate265inter3));
  inv1  gate1097(.a(s_79), .O(gate265inter4));
  nand2 gate1098(.a(gate265inter4), .b(gate265inter3), .O(gate265inter5));
  nor2  gate1099(.a(gate265inter5), .b(gate265inter2), .O(gate265inter6));
  inv1  gate1100(.a(G642), .O(gate265inter7));
  inv1  gate1101(.a(G770), .O(gate265inter8));
  nand2 gate1102(.a(gate265inter8), .b(gate265inter7), .O(gate265inter9));
  nand2 gate1103(.a(s_79), .b(gate265inter3), .O(gate265inter10));
  nor2  gate1104(.a(gate265inter10), .b(gate265inter9), .O(gate265inter11));
  nor2  gate1105(.a(gate265inter11), .b(gate265inter6), .O(gate265inter12));
  nand2 gate1106(.a(gate265inter12), .b(gate265inter1), .O(G794));
nand2 gate266( .a(G645), .b(G773), .O(G797) );
nand2 gate267( .a(G648), .b(G776), .O(G800) );

  xor2  gate1359(.a(G779), .b(G651), .O(gate268inter0));
  nand2 gate1360(.a(gate268inter0), .b(s_116), .O(gate268inter1));
  and2  gate1361(.a(G779), .b(G651), .O(gate268inter2));
  inv1  gate1362(.a(s_116), .O(gate268inter3));
  inv1  gate1363(.a(s_117), .O(gate268inter4));
  nand2 gate1364(.a(gate268inter4), .b(gate268inter3), .O(gate268inter5));
  nor2  gate1365(.a(gate268inter5), .b(gate268inter2), .O(gate268inter6));
  inv1  gate1366(.a(G651), .O(gate268inter7));
  inv1  gate1367(.a(G779), .O(gate268inter8));
  nand2 gate1368(.a(gate268inter8), .b(gate268inter7), .O(gate268inter9));
  nand2 gate1369(.a(s_117), .b(gate268inter3), .O(gate268inter10));
  nor2  gate1370(.a(gate268inter10), .b(gate268inter9), .O(gate268inter11));
  nor2  gate1371(.a(gate268inter11), .b(gate268inter6), .O(gate268inter12));
  nand2 gate1372(.a(gate268inter12), .b(gate268inter1), .O(G803));
nand2 gate269( .a(G654), .b(G782), .O(G806) );

  xor2  gate1443(.a(G785), .b(G657), .O(gate270inter0));
  nand2 gate1444(.a(gate270inter0), .b(s_128), .O(gate270inter1));
  and2  gate1445(.a(G785), .b(G657), .O(gate270inter2));
  inv1  gate1446(.a(s_128), .O(gate270inter3));
  inv1  gate1447(.a(s_129), .O(gate270inter4));
  nand2 gate1448(.a(gate270inter4), .b(gate270inter3), .O(gate270inter5));
  nor2  gate1449(.a(gate270inter5), .b(gate270inter2), .O(gate270inter6));
  inv1  gate1450(.a(G657), .O(gate270inter7));
  inv1  gate1451(.a(G785), .O(gate270inter8));
  nand2 gate1452(.a(gate270inter8), .b(gate270inter7), .O(gate270inter9));
  nand2 gate1453(.a(s_129), .b(gate270inter3), .O(gate270inter10));
  nor2  gate1454(.a(gate270inter10), .b(gate270inter9), .O(gate270inter11));
  nor2  gate1455(.a(gate270inter11), .b(gate270inter6), .O(gate270inter12));
  nand2 gate1456(.a(gate270inter12), .b(gate270inter1), .O(G809));
nand2 gate271( .a(G660), .b(G788), .O(G812) );
nand2 gate272( .a(G663), .b(G791), .O(G815) );
nand2 gate273( .a(G642), .b(G794), .O(G818) );

  xor2  gate1345(.a(G794), .b(G770), .O(gate274inter0));
  nand2 gate1346(.a(gate274inter0), .b(s_114), .O(gate274inter1));
  and2  gate1347(.a(G794), .b(G770), .O(gate274inter2));
  inv1  gate1348(.a(s_114), .O(gate274inter3));
  inv1  gate1349(.a(s_115), .O(gate274inter4));
  nand2 gate1350(.a(gate274inter4), .b(gate274inter3), .O(gate274inter5));
  nor2  gate1351(.a(gate274inter5), .b(gate274inter2), .O(gate274inter6));
  inv1  gate1352(.a(G770), .O(gate274inter7));
  inv1  gate1353(.a(G794), .O(gate274inter8));
  nand2 gate1354(.a(gate274inter8), .b(gate274inter7), .O(gate274inter9));
  nand2 gate1355(.a(s_115), .b(gate274inter3), .O(gate274inter10));
  nor2  gate1356(.a(gate274inter10), .b(gate274inter9), .O(gate274inter11));
  nor2  gate1357(.a(gate274inter11), .b(gate274inter6), .O(gate274inter12));
  nand2 gate1358(.a(gate274inter12), .b(gate274inter1), .O(G819));
nand2 gate275( .a(G645), .b(G797), .O(G820) );
nand2 gate276( .a(G773), .b(G797), .O(G821) );
nand2 gate277( .a(G648), .b(G800), .O(G822) );

  xor2  gate799(.a(G800), .b(G776), .O(gate278inter0));
  nand2 gate800(.a(gate278inter0), .b(s_36), .O(gate278inter1));
  and2  gate801(.a(G800), .b(G776), .O(gate278inter2));
  inv1  gate802(.a(s_36), .O(gate278inter3));
  inv1  gate803(.a(s_37), .O(gate278inter4));
  nand2 gate804(.a(gate278inter4), .b(gate278inter3), .O(gate278inter5));
  nor2  gate805(.a(gate278inter5), .b(gate278inter2), .O(gate278inter6));
  inv1  gate806(.a(G776), .O(gate278inter7));
  inv1  gate807(.a(G800), .O(gate278inter8));
  nand2 gate808(.a(gate278inter8), .b(gate278inter7), .O(gate278inter9));
  nand2 gate809(.a(s_37), .b(gate278inter3), .O(gate278inter10));
  nor2  gate810(.a(gate278inter10), .b(gate278inter9), .O(gate278inter11));
  nor2  gate811(.a(gate278inter11), .b(gate278inter6), .O(gate278inter12));
  nand2 gate812(.a(gate278inter12), .b(gate278inter1), .O(G823));
nand2 gate279( .a(G651), .b(G803), .O(G824) );
nand2 gate280( .a(G779), .b(G803), .O(G825) );

  xor2  gate645(.a(G806), .b(G654), .O(gate281inter0));
  nand2 gate646(.a(gate281inter0), .b(s_14), .O(gate281inter1));
  and2  gate647(.a(G806), .b(G654), .O(gate281inter2));
  inv1  gate648(.a(s_14), .O(gate281inter3));
  inv1  gate649(.a(s_15), .O(gate281inter4));
  nand2 gate650(.a(gate281inter4), .b(gate281inter3), .O(gate281inter5));
  nor2  gate651(.a(gate281inter5), .b(gate281inter2), .O(gate281inter6));
  inv1  gate652(.a(G654), .O(gate281inter7));
  inv1  gate653(.a(G806), .O(gate281inter8));
  nand2 gate654(.a(gate281inter8), .b(gate281inter7), .O(gate281inter9));
  nand2 gate655(.a(s_15), .b(gate281inter3), .O(gate281inter10));
  nor2  gate656(.a(gate281inter10), .b(gate281inter9), .O(gate281inter11));
  nor2  gate657(.a(gate281inter11), .b(gate281inter6), .O(gate281inter12));
  nand2 gate658(.a(gate281inter12), .b(gate281inter1), .O(G826));

  xor2  gate785(.a(G806), .b(G782), .O(gate282inter0));
  nand2 gate786(.a(gate282inter0), .b(s_34), .O(gate282inter1));
  and2  gate787(.a(G806), .b(G782), .O(gate282inter2));
  inv1  gate788(.a(s_34), .O(gate282inter3));
  inv1  gate789(.a(s_35), .O(gate282inter4));
  nand2 gate790(.a(gate282inter4), .b(gate282inter3), .O(gate282inter5));
  nor2  gate791(.a(gate282inter5), .b(gate282inter2), .O(gate282inter6));
  inv1  gate792(.a(G782), .O(gate282inter7));
  inv1  gate793(.a(G806), .O(gate282inter8));
  nand2 gate794(.a(gate282inter8), .b(gate282inter7), .O(gate282inter9));
  nand2 gate795(.a(s_35), .b(gate282inter3), .O(gate282inter10));
  nor2  gate796(.a(gate282inter10), .b(gate282inter9), .O(gate282inter11));
  nor2  gate797(.a(gate282inter11), .b(gate282inter6), .O(gate282inter12));
  nand2 gate798(.a(gate282inter12), .b(gate282inter1), .O(G827));
nand2 gate283( .a(G657), .b(G809), .O(G828) );
nand2 gate284( .a(G785), .b(G809), .O(G829) );
nand2 gate285( .a(G660), .b(G812), .O(G830) );

  xor2  gate1779(.a(G812), .b(G788), .O(gate286inter0));
  nand2 gate1780(.a(gate286inter0), .b(s_176), .O(gate286inter1));
  and2  gate1781(.a(G812), .b(G788), .O(gate286inter2));
  inv1  gate1782(.a(s_176), .O(gate286inter3));
  inv1  gate1783(.a(s_177), .O(gate286inter4));
  nand2 gate1784(.a(gate286inter4), .b(gate286inter3), .O(gate286inter5));
  nor2  gate1785(.a(gate286inter5), .b(gate286inter2), .O(gate286inter6));
  inv1  gate1786(.a(G788), .O(gate286inter7));
  inv1  gate1787(.a(G812), .O(gate286inter8));
  nand2 gate1788(.a(gate286inter8), .b(gate286inter7), .O(gate286inter9));
  nand2 gate1789(.a(s_177), .b(gate286inter3), .O(gate286inter10));
  nor2  gate1790(.a(gate286inter10), .b(gate286inter9), .O(gate286inter11));
  nor2  gate1791(.a(gate286inter11), .b(gate286inter6), .O(gate286inter12));
  nand2 gate1792(.a(gate286inter12), .b(gate286inter1), .O(G831));

  xor2  gate1303(.a(G815), .b(G663), .O(gate287inter0));
  nand2 gate1304(.a(gate287inter0), .b(s_108), .O(gate287inter1));
  and2  gate1305(.a(G815), .b(G663), .O(gate287inter2));
  inv1  gate1306(.a(s_108), .O(gate287inter3));
  inv1  gate1307(.a(s_109), .O(gate287inter4));
  nand2 gate1308(.a(gate287inter4), .b(gate287inter3), .O(gate287inter5));
  nor2  gate1309(.a(gate287inter5), .b(gate287inter2), .O(gate287inter6));
  inv1  gate1310(.a(G663), .O(gate287inter7));
  inv1  gate1311(.a(G815), .O(gate287inter8));
  nand2 gate1312(.a(gate287inter8), .b(gate287inter7), .O(gate287inter9));
  nand2 gate1313(.a(s_109), .b(gate287inter3), .O(gate287inter10));
  nor2  gate1314(.a(gate287inter10), .b(gate287inter9), .O(gate287inter11));
  nor2  gate1315(.a(gate287inter11), .b(gate287inter6), .O(gate287inter12));
  nand2 gate1316(.a(gate287inter12), .b(gate287inter1), .O(G832));
nand2 gate288( .a(G791), .b(G815), .O(G833) );
nand2 gate289( .a(G818), .b(G819), .O(G834) );
nand2 gate290( .a(G820), .b(G821), .O(G847) );
nand2 gate291( .a(G822), .b(G823), .O(G860) );

  xor2  gate1387(.a(G825), .b(G824), .O(gate292inter0));
  nand2 gate1388(.a(gate292inter0), .b(s_120), .O(gate292inter1));
  and2  gate1389(.a(G825), .b(G824), .O(gate292inter2));
  inv1  gate1390(.a(s_120), .O(gate292inter3));
  inv1  gate1391(.a(s_121), .O(gate292inter4));
  nand2 gate1392(.a(gate292inter4), .b(gate292inter3), .O(gate292inter5));
  nor2  gate1393(.a(gate292inter5), .b(gate292inter2), .O(gate292inter6));
  inv1  gate1394(.a(G824), .O(gate292inter7));
  inv1  gate1395(.a(G825), .O(gate292inter8));
  nand2 gate1396(.a(gate292inter8), .b(gate292inter7), .O(gate292inter9));
  nand2 gate1397(.a(s_121), .b(gate292inter3), .O(gate292inter10));
  nor2  gate1398(.a(gate292inter10), .b(gate292inter9), .O(gate292inter11));
  nor2  gate1399(.a(gate292inter11), .b(gate292inter6), .O(gate292inter12));
  nand2 gate1400(.a(gate292inter12), .b(gate292inter1), .O(G873));
nand2 gate293( .a(G828), .b(G829), .O(G886) );
nand2 gate294( .a(G832), .b(G833), .O(G899) );

  xor2  gate1275(.a(G831), .b(G830), .O(gate295inter0));
  nand2 gate1276(.a(gate295inter0), .b(s_104), .O(gate295inter1));
  and2  gate1277(.a(G831), .b(G830), .O(gate295inter2));
  inv1  gate1278(.a(s_104), .O(gate295inter3));
  inv1  gate1279(.a(s_105), .O(gate295inter4));
  nand2 gate1280(.a(gate295inter4), .b(gate295inter3), .O(gate295inter5));
  nor2  gate1281(.a(gate295inter5), .b(gate295inter2), .O(gate295inter6));
  inv1  gate1282(.a(G830), .O(gate295inter7));
  inv1  gate1283(.a(G831), .O(gate295inter8));
  nand2 gate1284(.a(gate295inter8), .b(gate295inter7), .O(gate295inter9));
  nand2 gate1285(.a(s_105), .b(gate295inter3), .O(gate295inter10));
  nor2  gate1286(.a(gate295inter10), .b(gate295inter9), .O(gate295inter11));
  nor2  gate1287(.a(gate295inter11), .b(gate295inter6), .O(gate295inter12));
  nand2 gate1288(.a(gate295inter12), .b(gate295inter1), .O(G912));

  xor2  gate1597(.a(G827), .b(G826), .O(gate296inter0));
  nand2 gate1598(.a(gate296inter0), .b(s_150), .O(gate296inter1));
  and2  gate1599(.a(G827), .b(G826), .O(gate296inter2));
  inv1  gate1600(.a(s_150), .O(gate296inter3));
  inv1  gate1601(.a(s_151), .O(gate296inter4));
  nand2 gate1602(.a(gate296inter4), .b(gate296inter3), .O(gate296inter5));
  nor2  gate1603(.a(gate296inter5), .b(gate296inter2), .O(gate296inter6));
  inv1  gate1604(.a(G826), .O(gate296inter7));
  inv1  gate1605(.a(G827), .O(gate296inter8));
  nand2 gate1606(.a(gate296inter8), .b(gate296inter7), .O(gate296inter9));
  nand2 gate1607(.a(s_151), .b(gate296inter3), .O(gate296inter10));
  nor2  gate1608(.a(gate296inter10), .b(gate296inter9), .O(gate296inter11));
  nor2  gate1609(.a(gate296inter11), .b(gate296inter6), .O(gate296inter12));
  nand2 gate1610(.a(gate296inter12), .b(gate296inter1), .O(G925));
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );
nand2 gate387( .a(G1), .b(G1036), .O(G1132) );
nand2 gate388( .a(G2), .b(G1039), .O(G1135) );
nand2 gate389( .a(G3), .b(G1042), .O(G1138) );
nand2 gate390( .a(G4), .b(G1045), .O(G1141) );
nand2 gate391( .a(G5), .b(G1048), .O(G1144) );

  xor2  gate575(.a(G1051), .b(G6), .O(gate392inter0));
  nand2 gate576(.a(gate392inter0), .b(s_4), .O(gate392inter1));
  and2  gate577(.a(G1051), .b(G6), .O(gate392inter2));
  inv1  gate578(.a(s_4), .O(gate392inter3));
  inv1  gate579(.a(s_5), .O(gate392inter4));
  nand2 gate580(.a(gate392inter4), .b(gate392inter3), .O(gate392inter5));
  nor2  gate581(.a(gate392inter5), .b(gate392inter2), .O(gate392inter6));
  inv1  gate582(.a(G6), .O(gate392inter7));
  inv1  gate583(.a(G1051), .O(gate392inter8));
  nand2 gate584(.a(gate392inter8), .b(gate392inter7), .O(gate392inter9));
  nand2 gate585(.a(s_5), .b(gate392inter3), .O(gate392inter10));
  nor2  gate586(.a(gate392inter10), .b(gate392inter9), .O(gate392inter11));
  nor2  gate587(.a(gate392inter11), .b(gate392inter6), .O(gate392inter12));
  nand2 gate588(.a(gate392inter12), .b(gate392inter1), .O(G1147));

  xor2  gate1611(.a(G1054), .b(G7), .O(gate393inter0));
  nand2 gate1612(.a(gate393inter0), .b(s_152), .O(gate393inter1));
  and2  gate1613(.a(G1054), .b(G7), .O(gate393inter2));
  inv1  gate1614(.a(s_152), .O(gate393inter3));
  inv1  gate1615(.a(s_153), .O(gate393inter4));
  nand2 gate1616(.a(gate393inter4), .b(gate393inter3), .O(gate393inter5));
  nor2  gate1617(.a(gate393inter5), .b(gate393inter2), .O(gate393inter6));
  inv1  gate1618(.a(G7), .O(gate393inter7));
  inv1  gate1619(.a(G1054), .O(gate393inter8));
  nand2 gate1620(.a(gate393inter8), .b(gate393inter7), .O(gate393inter9));
  nand2 gate1621(.a(s_153), .b(gate393inter3), .O(gate393inter10));
  nor2  gate1622(.a(gate393inter10), .b(gate393inter9), .O(gate393inter11));
  nor2  gate1623(.a(gate393inter11), .b(gate393inter6), .O(gate393inter12));
  nand2 gate1624(.a(gate393inter12), .b(gate393inter1), .O(G1150));
nand2 gate394( .a(G8), .b(G1057), .O(G1153) );
nand2 gate395( .a(G9), .b(G1060), .O(G1156) );
nand2 gate396( .a(G10), .b(G1063), .O(G1159) );
nand2 gate397( .a(G11), .b(G1066), .O(G1162) );
nand2 gate398( .a(G12), .b(G1069), .O(G1165) );
nand2 gate399( .a(G13), .b(G1072), .O(G1168) );
nand2 gate400( .a(G14), .b(G1075), .O(G1171) );
nand2 gate401( .a(G15), .b(G1078), .O(G1174) );
nand2 gate402( .a(G16), .b(G1081), .O(G1177) );
nand2 gate403( .a(G17), .b(G1084), .O(G1180) );

  xor2  gate1065(.a(G1087), .b(G18), .O(gate404inter0));
  nand2 gate1066(.a(gate404inter0), .b(s_74), .O(gate404inter1));
  and2  gate1067(.a(G1087), .b(G18), .O(gate404inter2));
  inv1  gate1068(.a(s_74), .O(gate404inter3));
  inv1  gate1069(.a(s_75), .O(gate404inter4));
  nand2 gate1070(.a(gate404inter4), .b(gate404inter3), .O(gate404inter5));
  nor2  gate1071(.a(gate404inter5), .b(gate404inter2), .O(gate404inter6));
  inv1  gate1072(.a(G18), .O(gate404inter7));
  inv1  gate1073(.a(G1087), .O(gate404inter8));
  nand2 gate1074(.a(gate404inter8), .b(gate404inter7), .O(gate404inter9));
  nand2 gate1075(.a(s_75), .b(gate404inter3), .O(gate404inter10));
  nor2  gate1076(.a(gate404inter10), .b(gate404inter9), .O(gate404inter11));
  nor2  gate1077(.a(gate404inter11), .b(gate404inter6), .O(gate404inter12));
  nand2 gate1078(.a(gate404inter12), .b(gate404inter1), .O(G1183));
nand2 gate405( .a(G19), .b(G1090), .O(G1186) );
nand2 gate406( .a(G20), .b(G1093), .O(G1189) );
nand2 gate407( .a(G21), .b(G1096), .O(G1192) );
nand2 gate408( .a(G22), .b(G1099), .O(G1195) );

  xor2  gate1261(.a(G1102), .b(G23), .O(gate409inter0));
  nand2 gate1262(.a(gate409inter0), .b(s_102), .O(gate409inter1));
  and2  gate1263(.a(G1102), .b(G23), .O(gate409inter2));
  inv1  gate1264(.a(s_102), .O(gate409inter3));
  inv1  gate1265(.a(s_103), .O(gate409inter4));
  nand2 gate1266(.a(gate409inter4), .b(gate409inter3), .O(gate409inter5));
  nor2  gate1267(.a(gate409inter5), .b(gate409inter2), .O(gate409inter6));
  inv1  gate1268(.a(G23), .O(gate409inter7));
  inv1  gate1269(.a(G1102), .O(gate409inter8));
  nand2 gate1270(.a(gate409inter8), .b(gate409inter7), .O(gate409inter9));
  nand2 gate1271(.a(s_103), .b(gate409inter3), .O(gate409inter10));
  nor2  gate1272(.a(gate409inter10), .b(gate409inter9), .O(gate409inter11));
  nor2  gate1273(.a(gate409inter11), .b(gate409inter6), .O(gate409inter12));
  nand2 gate1274(.a(gate409inter12), .b(gate409inter1), .O(G1198));

  xor2  gate995(.a(G1105), .b(G24), .O(gate410inter0));
  nand2 gate996(.a(gate410inter0), .b(s_64), .O(gate410inter1));
  and2  gate997(.a(G1105), .b(G24), .O(gate410inter2));
  inv1  gate998(.a(s_64), .O(gate410inter3));
  inv1  gate999(.a(s_65), .O(gate410inter4));
  nand2 gate1000(.a(gate410inter4), .b(gate410inter3), .O(gate410inter5));
  nor2  gate1001(.a(gate410inter5), .b(gate410inter2), .O(gate410inter6));
  inv1  gate1002(.a(G24), .O(gate410inter7));
  inv1  gate1003(.a(G1105), .O(gate410inter8));
  nand2 gate1004(.a(gate410inter8), .b(gate410inter7), .O(gate410inter9));
  nand2 gate1005(.a(s_65), .b(gate410inter3), .O(gate410inter10));
  nor2  gate1006(.a(gate410inter10), .b(gate410inter9), .O(gate410inter11));
  nor2  gate1007(.a(gate410inter11), .b(gate410inter6), .O(gate410inter12));
  nand2 gate1008(.a(gate410inter12), .b(gate410inter1), .O(G1201));
nand2 gate411( .a(G25), .b(G1108), .O(G1204) );

  xor2  gate953(.a(G1111), .b(G26), .O(gate412inter0));
  nand2 gate954(.a(gate412inter0), .b(s_58), .O(gate412inter1));
  and2  gate955(.a(G1111), .b(G26), .O(gate412inter2));
  inv1  gate956(.a(s_58), .O(gate412inter3));
  inv1  gate957(.a(s_59), .O(gate412inter4));
  nand2 gate958(.a(gate412inter4), .b(gate412inter3), .O(gate412inter5));
  nor2  gate959(.a(gate412inter5), .b(gate412inter2), .O(gate412inter6));
  inv1  gate960(.a(G26), .O(gate412inter7));
  inv1  gate961(.a(G1111), .O(gate412inter8));
  nand2 gate962(.a(gate412inter8), .b(gate412inter7), .O(gate412inter9));
  nand2 gate963(.a(s_59), .b(gate412inter3), .O(gate412inter10));
  nor2  gate964(.a(gate412inter10), .b(gate412inter9), .O(gate412inter11));
  nor2  gate965(.a(gate412inter11), .b(gate412inter6), .O(gate412inter12));
  nand2 gate966(.a(gate412inter12), .b(gate412inter1), .O(G1207));
nand2 gate413( .a(G27), .b(G1114), .O(G1210) );
nand2 gate414( .a(G28), .b(G1117), .O(G1213) );

  xor2  gate939(.a(G1120), .b(G29), .O(gate415inter0));
  nand2 gate940(.a(gate415inter0), .b(s_56), .O(gate415inter1));
  and2  gate941(.a(G1120), .b(G29), .O(gate415inter2));
  inv1  gate942(.a(s_56), .O(gate415inter3));
  inv1  gate943(.a(s_57), .O(gate415inter4));
  nand2 gate944(.a(gate415inter4), .b(gate415inter3), .O(gate415inter5));
  nor2  gate945(.a(gate415inter5), .b(gate415inter2), .O(gate415inter6));
  inv1  gate946(.a(G29), .O(gate415inter7));
  inv1  gate947(.a(G1120), .O(gate415inter8));
  nand2 gate948(.a(gate415inter8), .b(gate415inter7), .O(gate415inter9));
  nand2 gate949(.a(s_57), .b(gate415inter3), .O(gate415inter10));
  nor2  gate950(.a(gate415inter10), .b(gate415inter9), .O(gate415inter11));
  nor2  gate951(.a(gate415inter11), .b(gate415inter6), .O(gate415inter12));
  nand2 gate952(.a(gate415inter12), .b(gate415inter1), .O(G1216));
nand2 gate416( .a(G30), .b(G1123), .O(G1219) );

  xor2  gate1793(.a(G1126), .b(G31), .O(gate417inter0));
  nand2 gate1794(.a(gate417inter0), .b(s_178), .O(gate417inter1));
  and2  gate1795(.a(G1126), .b(G31), .O(gate417inter2));
  inv1  gate1796(.a(s_178), .O(gate417inter3));
  inv1  gate1797(.a(s_179), .O(gate417inter4));
  nand2 gate1798(.a(gate417inter4), .b(gate417inter3), .O(gate417inter5));
  nor2  gate1799(.a(gate417inter5), .b(gate417inter2), .O(gate417inter6));
  inv1  gate1800(.a(G31), .O(gate417inter7));
  inv1  gate1801(.a(G1126), .O(gate417inter8));
  nand2 gate1802(.a(gate417inter8), .b(gate417inter7), .O(gate417inter9));
  nand2 gate1803(.a(s_179), .b(gate417inter3), .O(gate417inter10));
  nor2  gate1804(.a(gate417inter10), .b(gate417inter9), .O(gate417inter11));
  nor2  gate1805(.a(gate417inter11), .b(gate417inter6), .O(gate417inter12));
  nand2 gate1806(.a(gate417inter12), .b(gate417inter1), .O(G1222));
nand2 gate418( .a(G32), .b(G1129), .O(G1225) );
nand2 gate419( .a(G1), .b(G1132), .O(G1228) );
nand2 gate420( .a(G1036), .b(G1132), .O(G1229) );
nand2 gate421( .a(G2), .b(G1135), .O(G1230) );
nand2 gate422( .a(G1039), .b(G1135), .O(G1231) );

  xor2  gate1373(.a(G1138), .b(G3), .O(gate423inter0));
  nand2 gate1374(.a(gate423inter0), .b(s_118), .O(gate423inter1));
  and2  gate1375(.a(G1138), .b(G3), .O(gate423inter2));
  inv1  gate1376(.a(s_118), .O(gate423inter3));
  inv1  gate1377(.a(s_119), .O(gate423inter4));
  nand2 gate1378(.a(gate423inter4), .b(gate423inter3), .O(gate423inter5));
  nor2  gate1379(.a(gate423inter5), .b(gate423inter2), .O(gate423inter6));
  inv1  gate1380(.a(G3), .O(gate423inter7));
  inv1  gate1381(.a(G1138), .O(gate423inter8));
  nand2 gate1382(.a(gate423inter8), .b(gate423inter7), .O(gate423inter9));
  nand2 gate1383(.a(s_119), .b(gate423inter3), .O(gate423inter10));
  nor2  gate1384(.a(gate423inter10), .b(gate423inter9), .O(gate423inter11));
  nor2  gate1385(.a(gate423inter11), .b(gate423inter6), .O(gate423inter12));
  nand2 gate1386(.a(gate423inter12), .b(gate423inter1), .O(G1232));
nand2 gate424( .a(G1042), .b(G1138), .O(G1233) );
nand2 gate425( .a(G4), .b(G1141), .O(G1234) );

  xor2  gate673(.a(G1141), .b(G1045), .O(gate426inter0));
  nand2 gate674(.a(gate426inter0), .b(s_18), .O(gate426inter1));
  and2  gate675(.a(G1141), .b(G1045), .O(gate426inter2));
  inv1  gate676(.a(s_18), .O(gate426inter3));
  inv1  gate677(.a(s_19), .O(gate426inter4));
  nand2 gate678(.a(gate426inter4), .b(gate426inter3), .O(gate426inter5));
  nor2  gate679(.a(gate426inter5), .b(gate426inter2), .O(gate426inter6));
  inv1  gate680(.a(G1045), .O(gate426inter7));
  inv1  gate681(.a(G1141), .O(gate426inter8));
  nand2 gate682(.a(gate426inter8), .b(gate426inter7), .O(gate426inter9));
  nand2 gate683(.a(s_19), .b(gate426inter3), .O(gate426inter10));
  nor2  gate684(.a(gate426inter10), .b(gate426inter9), .O(gate426inter11));
  nor2  gate685(.a(gate426inter11), .b(gate426inter6), .O(gate426inter12));
  nand2 gate686(.a(gate426inter12), .b(gate426inter1), .O(G1235));
nand2 gate427( .a(G5), .b(G1144), .O(G1236) );
nand2 gate428( .a(G1048), .b(G1144), .O(G1237) );
nand2 gate429( .a(G6), .b(G1147), .O(G1238) );
nand2 gate430( .a(G1051), .b(G1147), .O(G1239) );
nand2 gate431( .a(G7), .b(G1150), .O(G1240) );
nand2 gate432( .a(G1054), .b(G1150), .O(G1241) );
nand2 gate433( .a(G8), .b(G1153), .O(G1242) );
nand2 gate434( .a(G1057), .b(G1153), .O(G1243) );
nand2 gate435( .a(G9), .b(G1156), .O(G1244) );
nand2 gate436( .a(G1060), .b(G1156), .O(G1245) );

  xor2  gate2017(.a(G1159), .b(G10), .O(gate437inter0));
  nand2 gate2018(.a(gate437inter0), .b(s_210), .O(gate437inter1));
  and2  gate2019(.a(G1159), .b(G10), .O(gate437inter2));
  inv1  gate2020(.a(s_210), .O(gate437inter3));
  inv1  gate2021(.a(s_211), .O(gate437inter4));
  nand2 gate2022(.a(gate437inter4), .b(gate437inter3), .O(gate437inter5));
  nor2  gate2023(.a(gate437inter5), .b(gate437inter2), .O(gate437inter6));
  inv1  gate2024(.a(G10), .O(gate437inter7));
  inv1  gate2025(.a(G1159), .O(gate437inter8));
  nand2 gate2026(.a(gate437inter8), .b(gate437inter7), .O(gate437inter9));
  nand2 gate2027(.a(s_211), .b(gate437inter3), .O(gate437inter10));
  nor2  gate2028(.a(gate437inter10), .b(gate437inter9), .O(gate437inter11));
  nor2  gate2029(.a(gate437inter11), .b(gate437inter6), .O(gate437inter12));
  nand2 gate2030(.a(gate437inter12), .b(gate437inter1), .O(G1246));
nand2 gate438( .a(G1063), .b(G1159), .O(G1247) );
nand2 gate439( .a(G11), .b(G1162), .O(G1248) );
nand2 gate440( .a(G1066), .b(G1162), .O(G1249) );
nand2 gate441( .a(G12), .b(G1165), .O(G1250) );
nand2 gate442( .a(G1069), .b(G1165), .O(G1251) );
nand2 gate443( .a(G13), .b(G1168), .O(G1252) );
nand2 gate444( .a(G1072), .b(G1168), .O(G1253) );
nand2 gate445( .a(G14), .b(G1171), .O(G1254) );
nand2 gate446( .a(G1075), .b(G1171), .O(G1255) );
nand2 gate447( .a(G15), .b(G1174), .O(G1256) );

  xor2  gate1023(.a(G1174), .b(G1078), .O(gate448inter0));
  nand2 gate1024(.a(gate448inter0), .b(s_68), .O(gate448inter1));
  and2  gate1025(.a(G1174), .b(G1078), .O(gate448inter2));
  inv1  gate1026(.a(s_68), .O(gate448inter3));
  inv1  gate1027(.a(s_69), .O(gate448inter4));
  nand2 gate1028(.a(gate448inter4), .b(gate448inter3), .O(gate448inter5));
  nor2  gate1029(.a(gate448inter5), .b(gate448inter2), .O(gate448inter6));
  inv1  gate1030(.a(G1078), .O(gate448inter7));
  inv1  gate1031(.a(G1174), .O(gate448inter8));
  nand2 gate1032(.a(gate448inter8), .b(gate448inter7), .O(gate448inter9));
  nand2 gate1033(.a(s_69), .b(gate448inter3), .O(gate448inter10));
  nor2  gate1034(.a(gate448inter10), .b(gate448inter9), .O(gate448inter11));
  nor2  gate1035(.a(gate448inter11), .b(gate448inter6), .O(gate448inter12));
  nand2 gate1036(.a(gate448inter12), .b(gate448inter1), .O(G1257));
nand2 gate449( .a(G16), .b(G1177), .O(G1258) );
nand2 gate450( .a(G1081), .b(G1177), .O(G1259) );
nand2 gate451( .a(G17), .b(G1180), .O(G1260) );
nand2 gate452( .a(G1084), .b(G1180), .O(G1261) );
nand2 gate453( .a(G18), .b(G1183), .O(G1262) );

  xor2  gate1331(.a(G1183), .b(G1087), .O(gate454inter0));
  nand2 gate1332(.a(gate454inter0), .b(s_112), .O(gate454inter1));
  and2  gate1333(.a(G1183), .b(G1087), .O(gate454inter2));
  inv1  gate1334(.a(s_112), .O(gate454inter3));
  inv1  gate1335(.a(s_113), .O(gate454inter4));
  nand2 gate1336(.a(gate454inter4), .b(gate454inter3), .O(gate454inter5));
  nor2  gate1337(.a(gate454inter5), .b(gate454inter2), .O(gate454inter6));
  inv1  gate1338(.a(G1087), .O(gate454inter7));
  inv1  gate1339(.a(G1183), .O(gate454inter8));
  nand2 gate1340(.a(gate454inter8), .b(gate454inter7), .O(gate454inter9));
  nand2 gate1341(.a(s_113), .b(gate454inter3), .O(gate454inter10));
  nor2  gate1342(.a(gate454inter10), .b(gate454inter9), .O(gate454inter11));
  nor2  gate1343(.a(gate454inter11), .b(gate454inter6), .O(gate454inter12));
  nand2 gate1344(.a(gate454inter12), .b(gate454inter1), .O(G1263));
nand2 gate455( .a(G19), .b(G1186), .O(G1264) );
nand2 gate456( .a(G1090), .b(G1186), .O(G1265) );
nand2 gate457( .a(G20), .b(G1189), .O(G1266) );
nand2 gate458( .a(G1093), .b(G1189), .O(G1267) );
nand2 gate459( .a(G21), .b(G1192), .O(G1268) );
nand2 gate460( .a(G1096), .b(G1192), .O(G1269) );
nand2 gate461( .a(G22), .b(G1195), .O(G1270) );
nand2 gate462( .a(G1099), .b(G1195), .O(G1271) );
nand2 gate463( .a(G23), .b(G1198), .O(G1272) );
nand2 gate464( .a(G1102), .b(G1198), .O(G1273) );
nand2 gate465( .a(G24), .b(G1201), .O(G1274) );

  xor2  gate897(.a(G1201), .b(G1105), .O(gate466inter0));
  nand2 gate898(.a(gate466inter0), .b(s_50), .O(gate466inter1));
  and2  gate899(.a(G1201), .b(G1105), .O(gate466inter2));
  inv1  gate900(.a(s_50), .O(gate466inter3));
  inv1  gate901(.a(s_51), .O(gate466inter4));
  nand2 gate902(.a(gate466inter4), .b(gate466inter3), .O(gate466inter5));
  nor2  gate903(.a(gate466inter5), .b(gate466inter2), .O(gate466inter6));
  inv1  gate904(.a(G1105), .O(gate466inter7));
  inv1  gate905(.a(G1201), .O(gate466inter8));
  nand2 gate906(.a(gate466inter8), .b(gate466inter7), .O(gate466inter9));
  nand2 gate907(.a(s_51), .b(gate466inter3), .O(gate466inter10));
  nor2  gate908(.a(gate466inter10), .b(gate466inter9), .O(gate466inter11));
  nor2  gate909(.a(gate466inter11), .b(gate466inter6), .O(gate466inter12));
  nand2 gate910(.a(gate466inter12), .b(gate466inter1), .O(G1275));
nand2 gate467( .a(G25), .b(G1204), .O(G1276) );
nand2 gate468( .a(G1108), .b(G1204), .O(G1277) );
nand2 gate469( .a(G26), .b(G1207), .O(G1278) );
nand2 gate470( .a(G1111), .b(G1207), .O(G1279) );

  xor2  gate1457(.a(G1210), .b(G27), .O(gate471inter0));
  nand2 gate1458(.a(gate471inter0), .b(s_130), .O(gate471inter1));
  and2  gate1459(.a(G1210), .b(G27), .O(gate471inter2));
  inv1  gate1460(.a(s_130), .O(gate471inter3));
  inv1  gate1461(.a(s_131), .O(gate471inter4));
  nand2 gate1462(.a(gate471inter4), .b(gate471inter3), .O(gate471inter5));
  nor2  gate1463(.a(gate471inter5), .b(gate471inter2), .O(gate471inter6));
  inv1  gate1464(.a(G27), .O(gate471inter7));
  inv1  gate1465(.a(G1210), .O(gate471inter8));
  nand2 gate1466(.a(gate471inter8), .b(gate471inter7), .O(gate471inter9));
  nand2 gate1467(.a(s_131), .b(gate471inter3), .O(gate471inter10));
  nor2  gate1468(.a(gate471inter10), .b(gate471inter9), .O(gate471inter11));
  nor2  gate1469(.a(gate471inter11), .b(gate471inter6), .O(gate471inter12));
  nand2 gate1470(.a(gate471inter12), .b(gate471inter1), .O(G1280));
nand2 gate472( .a(G1114), .b(G1210), .O(G1281) );

  xor2  gate1415(.a(G1213), .b(G28), .O(gate473inter0));
  nand2 gate1416(.a(gate473inter0), .b(s_124), .O(gate473inter1));
  and2  gate1417(.a(G1213), .b(G28), .O(gate473inter2));
  inv1  gate1418(.a(s_124), .O(gate473inter3));
  inv1  gate1419(.a(s_125), .O(gate473inter4));
  nand2 gate1420(.a(gate473inter4), .b(gate473inter3), .O(gate473inter5));
  nor2  gate1421(.a(gate473inter5), .b(gate473inter2), .O(gate473inter6));
  inv1  gate1422(.a(G28), .O(gate473inter7));
  inv1  gate1423(.a(G1213), .O(gate473inter8));
  nand2 gate1424(.a(gate473inter8), .b(gate473inter7), .O(gate473inter9));
  nand2 gate1425(.a(s_125), .b(gate473inter3), .O(gate473inter10));
  nor2  gate1426(.a(gate473inter10), .b(gate473inter9), .O(gate473inter11));
  nor2  gate1427(.a(gate473inter11), .b(gate473inter6), .O(gate473inter12));
  nand2 gate1428(.a(gate473inter12), .b(gate473inter1), .O(G1282));
nand2 gate474( .a(G1117), .b(G1213), .O(G1283) );
nand2 gate475( .a(G29), .b(G1216), .O(G1284) );
nand2 gate476( .a(G1120), .b(G1216), .O(G1285) );
nand2 gate477( .a(G30), .b(G1219), .O(G1286) );
nand2 gate478( .a(G1123), .b(G1219), .O(G1287) );
nand2 gate479( .a(G31), .b(G1222), .O(G1288) );
nand2 gate480( .a(G1126), .b(G1222), .O(G1289) );
nand2 gate481( .a(G32), .b(G1225), .O(G1290) );
nand2 gate482( .a(G1129), .b(G1225), .O(G1291) );
nand2 gate483( .a(G1228), .b(G1229), .O(G1292) );

  xor2  gate1807(.a(G1231), .b(G1230), .O(gate484inter0));
  nand2 gate1808(.a(gate484inter0), .b(s_180), .O(gate484inter1));
  and2  gate1809(.a(G1231), .b(G1230), .O(gate484inter2));
  inv1  gate1810(.a(s_180), .O(gate484inter3));
  inv1  gate1811(.a(s_181), .O(gate484inter4));
  nand2 gate1812(.a(gate484inter4), .b(gate484inter3), .O(gate484inter5));
  nor2  gate1813(.a(gate484inter5), .b(gate484inter2), .O(gate484inter6));
  inv1  gate1814(.a(G1230), .O(gate484inter7));
  inv1  gate1815(.a(G1231), .O(gate484inter8));
  nand2 gate1816(.a(gate484inter8), .b(gate484inter7), .O(gate484inter9));
  nand2 gate1817(.a(s_181), .b(gate484inter3), .O(gate484inter10));
  nor2  gate1818(.a(gate484inter10), .b(gate484inter9), .O(gate484inter11));
  nor2  gate1819(.a(gate484inter11), .b(gate484inter6), .O(gate484inter12));
  nand2 gate1820(.a(gate484inter12), .b(gate484inter1), .O(G1293));

  xor2  gate1289(.a(G1233), .b(G1232), .O(gate485inter0));
  nand2 gate1290(.a(gate485inter0), .b(s_106), .O(gate485inter1));
  and2  gate1291(.a(G1233), .b(G1232), .O(gate485inter2));
  inv1  gate1292(.a(s_106), .O(gate485inter3));
  inv1  gate1293(.a(s_107), .O(gate485inter4));
  nand2 gate1294(.a(gate485inter4), .b(gate485inter3), .O(gate485inter5));
  nor2  gate1295(.a(gate485inter5), .b(gate485inter2), .O(gate485inter6));
  inv1  gate1296(.a(G1232), .O(gate485inter7));
  inv1  gate1297(.a(G1233), .O(gate485inter8));
  nand2 gate1298(.a(gate485inter8), .b(gate485inter7), .O(gate485inter9));
  nand2 gate1299(.a(s_107), .b(gate485inter3), .O(gate485inter10));
  nor2  gate1300(.a(gate485inter10), .b(gate485inter9), .O(gate485inter11));
  nor2  gate1301(.a(gate485inter11), .b(gate485inter6), .O(gate485inter12));
  nand2 gate1302(.a(gate485inter12), .b(gate485inter1), .O(G1294));

  xor2  gate1051(.a(G1235), .b(G1234), .O(gate486inter0));
  nand2 gate1052(.a(gate486inter0), .b(s_72), .O(gate486inter1));
  and2  gate1053(.a(G1235), .b(G1234), .O(gate486inter2));
  inv1  gate1054(.a(s_72), .O(gate486inter3));
  inv1  gate1055(.a(s_73), .O(gate486inter4));
  nand2 gate1056(.a(gate486inter4), .b(gate486inter3), .O(gate486inter5));
  nor2  gate1057(.a(gate486inter5), .b(gate486inter2), .O(gate486inter6));
  inv1  gate1058(.a(G1234), .O(gate486inter7));
  inv1  gate1059(.a(G1235), .O(gate486inter8));
  nand2 gate1060(.a(gate486inter8), .b(gate486inter7), .O(gate486inter9));
  nand2 gate1061(.a(s_73), .b(gate486inter3), .O(gate486inter10));
  nor2  gate1062(.a(gate486inter10), .b(gate486inter9), .O(gate486inter11));
  nor2  gate1063(.a(gate486inter11), .b(gate486inter6), .O(gate486inter12));
  nand2 gate1064(.a(gate486inter12), .b(gate486inter1), .O(G1295));

  xor2  gate1639(.a(G1237), .b(G1236), .O(gate487inter0));
  nand2 gate1640(.a(gate487inter0), .b(s_156), .O(gate487inter1));
  and2  gate1641(.a(G1237), .b(G1236), .O(gate487inter2));
  inv1  gate1642(.a(s_156), .O(gate487inter3));
  inv1  gate1643(.a(s_157), .O(gate487inter4));
  nand2 gate1644(.a(gate487inter4), .b(gate487inter3), .O(gate487inter5));
  nor2  gate1645(.a(gate487inter5), .b(gate487inter2), .O(gate487inter6));
  inv1  gate1646(.a(G1236), .O(gate487inter7));
  inv1  gate1647(.a(G1237), .O(gate487inter8));
  nand2 gate1648(.a(gate487inter8), .b(gate487inter7), .O(gate487inter9));
  nand2 gate1649(.a(s_157), .b(gate487inter3), .O(gate487inter10));
  nor2  gate1650(.a(gate487inter10), .b(gate487inter9), .O(gate487inter11));
  nor2  gate1651(.a(gate487inter11), .b(gate487inter6), .O(gate487inter12));
  nand2 gate1652(.a(gate487inter12), .b(gate487inter1), .O(G1296));
nand2 gate488( .a(G1238), .b(G1239), .O(G1297) );

  xor2  gate1569(.a(G1241), .b(G1240), .O(gate489inter0));
  nand2 gate1570(.a(gate489inter0), .b(s_146), .O(gate489inter1));
  and2  gate1571(.a(G1241), .b(G1240), .O(gate489inter2));
  inv1  gate1572(.a(s_146), .O(gate489inter3));
  inv1  gate1573(.a(s_147), .O(gate489inter4));
  nand2 gate1574(.a(gate489inter4), .b(gate489inter3), .O(gate489inter5));
  nor2  gate1575(.a(gate489inter5), .b(gate489inter2), .O(gate489inter6));
  inv1  gate1576(.a(G1240), .O(gate489inter7));
  inv1  gate1577(.a(G1241), .O(gate489inter8));
  nand2 gate1578(.a(gate489inter8), .b(gate489inter7), .O(gate489inter9));
  nand2 gate1579(.a(s_147), .b(gate489inter3), .O(gate489inter10));
  nor2  gate1580(.a(gate489inter10), .b(gate489inter9), .O(gate489inter11));
  nor2  gate1581(.a(gate489inter11), .b(gate489inter6), .O(gate489inter12));
  nand2 gate1582(.a(gate489inter12), .b(gate489inter1), .O(G1298));

  xor2  gate1821(.a(G1243), .b(G1242), .O(gate490inter0));
  nand2 gate1822(.a(gate490inter0), .b(s_182), .O(gate490inter1));
  and2  gate1823(.a(G1243), .b(G1242), .O(gate490inter2));
  inv1  gate1824(.a(s_182), .O(gate490inter3));
  inv1  gate1825(.a(s_183), .O(gate490inter4));
  nand2 gate1826(.a(gate490inter4), .b(gate490inter3), .O(gate490inter5));
  nor2  gate1827(.a(gate490inter5), .b(gate490inter2), .O(gate490inter6));
  inv1  gate1828(.a(G1242), .O(gate490inter7));
  inv1  gate1829(.a(G1243), .O(gate490inter8));
  nand2 gate1830(.a(gate490inter8), .b(gate490inter7), .O(gate490inter9));
  nand2 gate1831(.a(s_183), .b(gate490inter3), .O(gate490inter10));
  nor2  gate1832(.a(gate490inter10), .b(gate490inter9), .O(gate490inter11));
  nor2  gate1833(.a(gate490inter11), .b(gate490inter6), .O(gate490inter12));
  nand2 gate1834(.a(gate490inter12), .b(gate490inter1), .O(G1299));

  xor2  gate1681(.a(G1245), .b(G1244), .O(gate491inter0));
  nand2 gate1682(.a(gate491inter0), .b(s_162), .O(gate491inter1));
  and2  gate1683(.a(G1245), .b(G1244), .O(gate491inter2));
  inv1  gate1684(.a(s_162), .O(gate491inter3));
  inv1  gate1685(.a(s_163), .O(gate491inter4));
  nand2 gate1686(.a(gate491inter4), .b(gate491inter3), .O(gate491inter5));
  nor2  gate1687(.a(gate491inter5), .b(gate491inter2), .O(gate491inter6));
  inv1  gate1688(.a(G1244), .O(gate491inter7));
  inv1  gate1689(.a(G1245), .O(gate491inter8));
  nand2 gate1690(.a(gate491inter8), .b(gate491inter7), .O(gate491inter9));
  nand2 gate1691(.a(s_163), .b(gate491inter3), .O(gate491inter10));
  nor2  gate1692(.a(gate491inter10), .b(gate491inter9), .O(gate491inter11));
  nor2  gate1693(.a(gate491inter11), .b(gate491inter6), .O(gate491inter12));
  nand2 gate1694(.a(gate491inter12), .b(gate491inter1), .O(G1300));
nand2 gate492( .a(G1246), .b(G1247), .O(G1301) );
nand2 gate493( .a(G1248), .b(G1249), .O(G1302) );
nand2 gate494( .a(G1250), .b(G1251), .O(G1303) );
nand2 gate495( .a(G1252), .b(G1253), .O(G1304) );
nand2 gate496( .a(G1254), .b(G1255), .O(G1305) );

  xor2  gate1471(.a(G1257), .b(G1256), .O(gate497inter0));
  nand2 gate1472(.a(gate497inter0), .b(s_132), .O(gate497inter1));
  and2  gate1473(.a(G1257), .b(G1256), .O(gate497inter2));
  inv1  gate1474(.a(s_132), .O(gate497inter3));
  inv1  gate1475(.a(s_133), .O(gate497inter4));
  nand2 gate1476(.a(gate497inter4), .b(gate497inter3), .O(gate497inter5));
  nor2  gate1477(.a(gate497inter5), .b(gate497inter2), .O(gate497inter6));
  inv1  gate1478(.a(G1256), .O(gate497inter7));
  inv1  gate1479(.a(G1257), .O(gate497inter8));
  nand2 gate1480(.a(gate497inter8), .b(gate497inter7), .O(gate497inter9));
  nand2 gate1481(.a(s_133), .b(gate497inter3), .O(gate497inter10));
  nor2  gate1482(.a(gate497inter10), .b(gate497inter9), .O(gate497inter11));
  nor2  gate1483(.a(gate497inter11), .b(gate497inter6), .O(gate497inter12));
  nand2 gate1484(.a(gate497inter12), .b(gate497inter1), .O(G1306));
nand2 gate498( .a(G1258), .b(G1259), .O(G1307) );

  xor2  gate1933(.a(G1261), .b(G1260), .O(gate499inter0));
  nand2 gate1934(.a(gate499inter0), .b(s_198), .O(gate499inter1));
  and2  gate1935(.a(G1261), .b(G1260), .O(gate499inter2));
  inv1  gate1936(.a(s_198), .O(gate499inter3));
  inv1  gate1937(.a(s_199), .O(gate499inter4));
  nand2 gate1938(.a(gate499inter4), .b(gate499inter3), .O(gate499inter5));
  nor2  gate1939(.a(gate499inter5), .b(gate499inter2), .O(gate499inter6));
  inv1  gate1940(.a(G1260), .O(gate499inter7));
  inv1  gate1941(.a(G1261), .O(gate499inter8));
  nand2 gate1942(.a(gate499inter8), .b(gate499inter7), .O(gate499inter9));
  nand2 gate1943(.a(s_199), .b(gate499inter3), .O(gate499inter10));
  nor2  gate1944(.a(gate499inter10), .b(gate499inter9), .O(gate499inter11));
  nor2  gate1945(.a(gate499inter11), .b(gate499inter6), .O(gate499inter12));
  nand2 gate1946(.a(gate499inter12), .b(gate499inter1), .O(G1308));
nand2 gate500( .a(G1262), .b(G1263), .O(G1309) );

  xor2  gate1121(.a(G1265), .b(G1264), .O(gate501inter0));
  nand2 gate1122(.a(gate501inter0), .b(s_82), .O(gate501inter1));
  and2  gate1123(.a(G1265), .b(G1264), .O(gate501inter2));
  inv1  gate1124(.a(s_82), .O(gate501inter3));
  inv1  gate1125(.a(s_83), .O(gate501inter4));
  nand2 gate1126(.a(gate501inter4), .b(gate501inter3), .O(gate501inter5));
  nor2  gate1127(.a(gate501inter5), .b(gate501inter2), .O(gate501inter6));
  inv1  gate1128(.a(G1264), .O(gate501inter7));
  inv1  gate1129(.a(G1265), .O(gate501inter8));
  nand2 gate1130(.a(gate501inter8), .b(gate501inter7), .O(gate501inter9));
  nand2 gate1131(.a(s_83), .b(gate501inter3), .O(gate501inter10));
  nor2  gate1132(.a(gate501inter10), .b(gate501inter9), .O(gate501inter11));
  nor2  gate1133(.a(gate501inter11), .b(gate501inter6), .O(gate501inter12));
  nand2 gate1134(.a(gate501inter12), .b(gate501inter1), .O(G1310));
nand2 gate502( .a(G1266), .b(G1267), .O(G1311) );

  xor2  gate1079(.a(G1269), .b(G1268), .O(gate503inter0));
  nand2 gate1080(.a(gate503inter0), .b(s_76), .O(gate503inter1));
  and2  gate1081(.a(G1269), .b(G1268), .O(gate503inter2));
  inv1  gate1082(.a(s_76), .O(gate503inter3));
  inv1  gate1083(.a(s_77), .O(gate503inter4));
  nand2 gate1084(.a(gate503inter4), .b(gate503inter3), .O(gate503inter5));
  nor2  gate1085(.a(gate503inter5), .b(gate503inter2), .O(gate503inter6));
  inv1  gate1086(.a(G1268), .O(gate503inter7));
  inv1  gate1087(.a(G1269), .O(gate503inter8));
  nand2 gate1088(.a(gate503inter8), .b(gate503inter7), .O(gate503inter9));
  nand2 gate1089(.a(s_77), .b(gate503inter3), .O(gate503inter10));
  nor2  gate1090(.a(gate503inter10), .b(gate503inter9), .O(gate503inter11));
  nor2  gate1091(.a(gate503inter11), .b(gate503inter6), .O(gate503inter12));
  nand2 gate1092(.a(gate503inter12), .b(gate503inter1), .O(G1312));
nand2 gate504( .a(G1270), .b(G1271), .O(G1313) );
nand2 gate505( .a(G1272), .b(G1273), .O(G1314) );
nand2 gate506( .a(G1274), .b(G1275), .O(G1315) );
nand2 gate507( .a(G1276), .b(G1277), .O(G1316) );

  xor2  gate1905(.a(G1279), .b(G1278), .O(gate508inter0));
  nand2 gate1906(.a(gate508inter0), .b(s_194), .O(gate508inter1));
  and2  gate1907(.a(G1279), .b(G1278), .O(gate508inter2));
  inv1  gate1908(.a(s_194), .O(gate508inter3));
  inv1  gate1909(.a(s_195), .O(gate508inter4));
  nand2 gate1910(.a(gate508inter4), .b(gate508inter3), .O(gate508inter5));
  nor2  gate1911(.a(gate508inter5), .b(gate508inter2), .O(gate508inter6));
  inv1  gate1912(.a(G1278), .O(gate508inter7));
  inv1  gate1913(.a(G1279), .O(gate508inter8));
  nand2 gate1914(.a(gate508inter8), .b(gate508inter7), .O(gate508inter9));
  nand2 gate1915(.a(s_195), .b(gate508inter3), .O(gate508inter10));
  nor2  gate1916(.a(gate508inter10), .b(gate508inter9), .O(gate508inter11));
  nor2  gate1917(.a(gate508inter11), .b(gate508inter6), .O(gate508inter12));
  nand2 gate1918(.a(gate508inter12), .b(gate508inter1), .O(G1317));

  xor2  gate1513(.a(G1281), .b(G1280), .O(gate509inter0));
  nand2 gate1514(.a(gate509inter0), .b(s_138), .O(gate509inter1));
  and2  gate1515(.a(G1281), .b(G1280), .O(gate509inter2));
  inv1  gate1516(.a(s_138), .O(gate509inter3));
  inv1  gate1517(.a(s_139), .O(gate509inter4));
  nand2 gate1518(.a(gate509inter4), .b(gate509inter3), .O(gate509inter5));
  nor2  gate1519(.a(gate509inter5), .b(gate509inter2), .O(gate509inter6));
  inv1  gate1520(.a(G1280), .O(gate509inter7));
  inv1  gate1521(.a(G1281), .O(gate509inter8));
  nand2 gate1522(.a(gate509inter8), .b(gate509inter7), .O(gate509inter9));
  nand2 gate1523(.a(s_139), .b(gate509inter3), .O(gate509inter10));
  nor2  gate1524(.a(gate509inter10), .b(gate509inter9), .O(gate509inter11));
  nor2  gate1525(.a(gate509inter11), .b(gate509inter6), .O(gate509inter12));
  nand2 gate1526(.a(gate509inter12), .b(gate509inter1), .O(G1318));
nand2 gate510( .a(G1282), .b(G1283), .O(G1319) );

  xor2  gate1527(.a(G1285), .b(G1284), .O(gate511inter0));
  nand2 gate1528(.a(gate511inter0), .b(s_140), .O(gate511inter1));
  and2  gate1529(.a(G1285), .b(G1284), .O(gate511inter2));
  inv1  gate1530(.a(s_140), .O(gate511inter3));
  inv1  gate1531(.a(s_141), .O(gate511inter4));
  nand2 gate1532(.a(gate511inter4), .b(gate511inter3), .O(gate511inter5));
  nor2  gate1533(.a(gate511inter5), .b(gate511inter2), .O(gate511inter6));
  inv1  gate1534(.a(G1284), .O(gate511inter7));
  inv1  gate1535(.a(G1285), .O(gate511inter8));
  nand2 gate1536(.a(gate511inter8), .b(gate511inter7), .O(gate511inter9));
  nand2 gate1537(.a(s_141), .b(gate511inter3), .O(gate511inter10));
  nor2  gate1538(.a(gate511inter10), .b(gate511inter9), .O(gate511inter11));
  nor2  gate1539(.a(gate511inter11), .b(gate511inter6), .O(gate511inter12));
  nand2 gate1540(.a(gate511inter12), .b(gate511inter1), .O(G1320));
nand2 gate512( .a(G1286), .b(G1287), .O(G1321) );
nand2 gate513( .a(G1288), .b(G1289), .O(G1322) );

  xor2  gate1737(.a(G1291), .b(G1290), .O(gate514inter0));
  nand2 gate1738(.a(gate514inter0), .b(s_170), .O(gate514inter1));
  and2  gate1739(.a(G1291), .b(G1290), .O(gate514inter2));
  inv1  gate1740(.a(s_170), .O(gate514inter3));
  inv1  gate1741(.a(s_171), .O(gate514inter4));
  nand2 gate1742(.a(gate514inter4), .b(gate514inter3), .O(gate514inter5));
  nor2  gate1743(.a(gate514inter5), .b(gate514inter2), .O(gate514inter6));
  inv1  gate1744(.a(G1290), .O(gate514inter7));
  inv1  gate1745(.a(G1291), .O(gate514inter8));
  nand2 gate1746(.a(gate514inter8), .b(gate514inter7), .O(gate514inter9));
  nand2 gate1747(.a(s_171), .b(gate514inter3), .O(gate514inter10));
  nor2  gate1748(.a(gate514inter10), .b(gate514inter9), .O(gate514inter11));
  nor2  gate1749(.a(gate514inter11), .b(gate514inter6), .O(gate514inter12));
  nand2 gate1750(.a(gate514inter12), .b(gate514inter1), .O(G1323));
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule