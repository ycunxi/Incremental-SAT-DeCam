module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);

input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;//RE__PI;

input s_0,s_1;//RE__ALLOW(00,01,10,11);
input s_2,s_3;//RE__ALLOW(00,01,10,11);
input s_4,s_5;//RE__ALLOW(00,01,10,11);
input s_6,s_7;//RE__ALLOW(00,01,10,11);
input s_8,s_9;//RE__ALLOW(00,01,10,11);
input s_10,s_11;//RE__ALLOW(00,01,10,11);
input s_12,s_13;//RE__ALLOW(00,01,10,11);
input s_14,s_15;//RE__ALLOW(00,01,10,11);
input s_16,s_17;//RE__ALLOW(00,01,10,11);
input s_18,s_19;//RE__ALLOW(00,01,10,11);
input s_20,s_21;//RE__ALLOW(00,01,10,11);
input s_22,s_23;//RE__ALLOW(00,01,10,11);
input s_24,s_25;//RE__ALLOW(00,01,10,11);
input s_26,s_27;//RE__ALLOW(00,01,10,11);
input s_28,s_29;//RE__ALLOW(00,01,10,11);
input s_30,s_31;//RE__ALLOW(00,01,10,11);
input s_32,s_33;//RE__ALLOW(00,01,10,11);
input s_34,s_35;//RE__ALLOW(00,01,10,11);
input s_36,s_37;//RE__ALLOW(00,01,10,11);
input s_38,s_39;//RE__ALLOW(00,01,10,11);
input s_40,s_41;//RE__ALLOW(00,01,10,11);
input s_42,s_43;//RE__ALLOW(00,01,10,11);
input s_44,s_45;//RE__ALLOW(00,01,10,11);
input s_46,s_47;//RE__ALLOW(00,01,10,11);
input s_48,s_49;//RE__ALLOW(00,01,10,11);
input s_50,s_51;//RE__ALLOW(00,01,10,11);
input s_52,s_53;//RE__ALLOW(00,01,10,11);
input s_54,s_55;//RE__ALLOW(00,01,10,11);
input s_56,s_57;//RE__ALLOW(00,01,10,11);
input s_58,s_59;//RE__ALLOW(00,01,10,11);
input s_60,s_61;//RE__ALLOW(00,01,10,11);
input s_62,s_63;//RE__ALLOW(00,01,10,11);
input s_64,s_65;//RE__ALLOW(00,01,10,11);
input s_66,s_67;//RE__ALLOW(00,01,10,11);
input s_68,s_69;//RE__ALLOW(00,01,10,11);
input s_70,s_71;//RE__ALLOW(00,01,10,11);
input s_72,s_73;//RE__ALLOW(00,01,10,11);
input s_74,s_75;//RE__ALLOW(00,01,10,11);
input s_76,s_77;//RE__ALLOW(00,01,10,11);
input s_78,s_79;//RE__ALLOW(00,01,10,11);
input s_80,s_81;//RE__ALLOW(00,01,10,11);
input s_82,s_83;//RE__ALLOW(00,01,10,11);
input s_84,s_85;//RE__ALLOW(00,01,10,11);
input s_86,s_87;//RE__ALLOW(00,01,10,11);
input s_88,s_89;//RE__ALLOW(00,01,10,11);
input s_90,s_91;//RE__ALLOW(00,01,10,11);
input s_92,s_93;//RE__ALLOW(00,01,10,11);
input s_94,s_95;//RE__ALLOW(00,01,10,11);
input s_96,s_97;//RE__ALLOW(00,01,10,11);
input s_98,s_99;//RE__ALLOW(00,01,10,11);
input s_100,s_101;//RE__ALLOW(00,01,10,11);
input s_102,s_103;//RE__ALLOW(00,01,10,11);
input s_104,s_105;//RE__ALLOW(00,01,10,11);
input s_106,s_107;//RE__ALLOW(00,01,10,11);
input s_108,s_109;//RE__ALLOW(00,01,10,11);
input s_110,s_111;//RE__ALLOW(00,01,10,11);
input s_112,s_113;//RE__ALLOW(00,01,10,11);
input s_114,s_115;//RE__ALLOW(00,01,10,11);
input s_116,s_117;//RE__ALLOW(00,01,10,11);
input s_118,s_119;//RE__ALLOW(00,01,10,11);
input s_120,s_121;//RE__ALLOW(00,01,10,11);
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;

  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate194inter0, gate194inter1, gate194inter2, gate194inter3, gate194inter4, gate194inter5, gate194inter6, gate194inter7, gate194inter8, gate194inter9, gate194inter10, gate194inter11, gate194inter12, gate468inter0, gate468inter1, gate468inter2, gate468inter3, gate468inter4, gate468inter5, gate468inter6, gate468inter7, gate468inter8, gate468inter9, gate468inter10, gate468inter11, gate468inter12, gate256inter0, gate256inter1, gate256inter2, gate256inter3, gate256inter4, gate256inter5, gate256inter6, gate256inter7, gate256inter8, gate256inter9, gate256inter10, gate256inter11, gate256inter12, gate398inter0, gate398inter1, gate398inter2, gate398inter3, gate398inter4, gate398inter5, gate398inter6, gate398inter7, gate398inter8, gate398inter9, gate398inter10, gate398inter11, gate398inter12, gate258inter0, gate258inter1, gate258inter2, gate258inter3, gate258inter4, gate258inter5, gate258inter6, gate258inter7, gate258inter8, gate258inter9, gate258inter10, gate258inter11, gate258inter12, gate244inter0, gate244inter1, gate244inter2, gate244inter3, gate244inter4, gate244inter5, gate244inter6, gate244inter7, gate244inter8, gate244inter9, gate244inter10, gate244inter11, gate244inter12, gate412inter0, gate412inter1, gate412inter2, gate412inter3, gate412inter4, gate412inter5, gate412inter6, gate412inter7, gate412inter8, gate412inter9, gate412inter10, gate412inter11, gate412inter12, gate13inter0, gate13inter1, gate13inter2, gate13inter3, gate13inter4, gate13inter5, gate13inter6, gate13inter7, gate13inter8, gate13inter9, gate13inter10, gate13inter11, gate13inter12, gate65inter0, gate65inter1, gate65inter2, gate65inter3, gate65inter4, gate65inter5, gate65inter6, gate65inter7, gate65inter8, gate65inter9, gate65inter10, gate65inter11, gate65inter12, gate128inter0, gate128inter1, gate128inter2, gate128inter3, gate128inter4, gate128inter5, gate128inter6, gate128inter7, gate128inter8, gate128inter9, gate128inter10, gate128inter11, gate128inter12, gate105inter0, gate105inter1, gate105inter2, gate105inter3, gate105inter4, gate105inter5, gate105inter6, gate105inter7, gate105inter8, gate105inter9, gate105inter10, gate105inter11, gate105inter12, gate243inter0, gate243inter1, gate243inter2, gate243inter3, gate243inter4, gate243inter5, gate243inter6, gate243inter7, gate243inter8, gate243inter9, gate243inter10, gate243inter11, gate243inter12, gate471inter0, gate471inter1, gate471inter2, gate471inter3, gate471inter4, gate471inter5, gate471inter6, gate471inter7, gate471inter8, gate471inter9, gate471inter10, gate471inter11, gate471inter12, gate176inter0, gate176inter1, gate176inter2, gate176inter3, gate176inter4, gate176inter5, gate176inter6, gate176inter7, gate176inter8, gate176inter9, gate176inter10, gate176inter11, gate176inter12, gate393inter0, gate393inter1, gate393inter2, gate393inter3, gate393inter4, gate393inter5, gate393inter6, gate393inter7, gate393inter8, gate393inter9, gate393inter10, gate393inter11, gate393inter12, gate253inter0, gate253inter1, gate253inter2, gate253inter3, gate253inter4, gate253inter5, gate253inter6, gate253inter7, gate253inter8, gate253inter9, gate253inter10, gate253inter11, gate253inter12, gate135inter0, gate135inter1, gate135inter2, gate135inter3, gate135inter4, gate135inter5, gate135inter6, gate135inter7, gate135inter8, gate135inter9, gate135inter10, gate135inter11, gate135inter12, gate481inter0, gate481inter1, gate481inter2, gate481inter3, gate481inter4, gate481inter5, gate481inter6, gate481inter7, gate481inter8, gate481inter9, gate481inter10, gate481inter11, gate481inter12, gate504inter0, gate504inter1, gate504inter2, gate504inter3, gate504inter4, gate504inter5, gate504inter6, gate504inter7, gate504inter8, gate504inter9, gate504inter10, gate504inter11, gate504inter12, gate284inter0, gate284inter1, gate284inter2, gate284inter3, gate284inter4, gate284inter5, gate284inter6, gate284inter7, gate284inter8, gate284inter9, gate284inter10, gate284inter11, gate284inter12, gate171inter0, gate171inter1, gate171inter2, gate171inter3, gate171inter4, gate171inter5, gate171inter6, gate171inter7, gate171inter8, gate171inter9, gate171inter10, gate171inter11, gate171inter12, gate53inter0, gate53inter1, gate53inter2, gate53inter3, gate53inter4, gate53inter5, gate53inter6, gate53inter7, gate53inter8, gate53inter9, gate53inter10, gate53inter11, gate53inter12, gate512inter0, gate512inter1, gate512inter2, gate512inter3, gate512inter4, gate512inter5, gate512inter6, gate512inter7, gate512inter8, gate512inter9, gate512inter10, gate512inter11, gate512inter12, gate441inter0, gate441inter1, gate441inter2, gate441inter3, gate441inter4, gate441inter5, gate441inter6, gate441inter7, gate441inter8, gate441inter9, gate441inter10, gate441inter11, gate441inter12, gate143inter0, gate143inter1, gate143inter2, gate143inter3, gate143inter4, gate143inter5, gate143inter6, gate143inter7, gate143inter8, gate143inter9, gate143inter10, gate143inter11, gate143inter12, gate19inter0, gate19inter1, gate19inter2, gate19inter3, gate19inter4, gate19inter5, gate19inter6, gate19inter7, gate19inter8, gate19inter9, gate19inter10, gate19inter11, gate19inter12, gate177inter0, gate177inter1, gate177inter2, gate177inter3, gate177inter4, gate177inter5, gate177inter6, gate177inter7, gate177inter8, gate177inter9, gate177inter10, gate177inter11, gate177inter12, gate79inter0, gate79inter1, gate79inter2, gate79inter3, gate79inter4, gate79inter5, gate79inter6, gate79inter7, gate79inter8, gate79inter9, gate79inter10, gate79inter11, gate79inter12, gate278inter0, gate278inter1, gate278inter2, gate278inter3, gate278inter4, gate278inter5, gate278inter6, gate278inter7, gate278inter8, gate278inter9, gate278inter10, gate278inter11, gate278inter12, gate275inter0, gate275inter1, gate275inter2, gate275inter3, gate275inter4, gate275inter5, gate275inter6, gate275inter7, gate275inter8, gate275inter9, gate275inter10, gate275inter11, gate275inter12, gate119inter0, gate119inter1, gate119inter2, gate119inter3, gate119inter4, gate119inter5, gate119inter6, gate119inter7, gate119inter8, gate119inter9, gate119inter10, gate119inter11, gate119inter12, gate71inter0, gate71inter1, gate71inter2, gate71inter3, gate71inter4, gate71inter5, gate71inter6, gate71inter7, gate71inter8, gate71inter9, gate71inter10, gate71inter11, gate71inter12, gate283inter0, gate283inter1, gate283inter2, gate283inter3, gate283inter4, gate283inter5, gate283inter6, gate283inter7, gate283inter8, gate283inter9, gate283inter10, gate283inter11, gate283inter12, gate26inter0, gate26inter1, gate26inter2, gate26inter3, gate26inter4, gate26inter5, gate26inter6, gate26inter7, gate26inter8, gate26inter9, gate26inter10, gate26inter11, gate26inter12, gate416inter0, gate416inter1, gate416inter2, gate416inter3, gate416inter4, gate416inter5, gate416inter6, gate416inter7, gate416inter8, gate416inter9, gate416inter10, gate416inter11, gate416inter12, gate34inter0, gate34inter1, gate34inter2, gate34inter3, gate34inter4, gate34inter5, gate34inter6, gate34inter7, gate34inter8, gate34inter9, gate34inter10, gate34inter11, gate34inter12, gate399inter0, gate399inter1, gate399inter2, gate399inter3, gate399inter4, gate399inter5, gate399inter6, gate399inter7, gate399inter8, gate399inter9, gate399inter10, gate399inter11, gate399inter12, gate9inter0, gate9inter1, gate9inter2, gate9inter3, gate9inter4, gate9inter5, gate9inter6, gate9inter7, gate9inter8, gate9inter9, gate9inter10, gate9inter11, gate9inter12, gate409inter0, gate409inter1, gate409inter2, gate409inter3, gate409inter4, gate409inter5, gate409inter6, gate409inter7, gate409inter8, gate409inter9, gate409inter10, gate409inter11, gate409inter12, gate457inter0, gate457inter1, gate457inter2, gate457inter3, gate457inter4, gate457inter5, gate457inter6, gate457inter7, gate457inter8, gate457inter9, gate457inter10, gate457inter11, gate457inter12, gate215inter0, gate215inter1, gate215inter2, gate215inter3, gate215inter4, gate215inter5, gate215inter6, gate215inter7, gate215inter8, gate215inter9, gate215inter10, gate215inter11, gate215inter12, gate201inter0, gate201inter1, gate201inter2, gate201inter3, gate201inter4, gate201inter5, gate201inter6, gate201inter7, gate201inter8, gate201inter9, gate201inter10, gate201inter11, gate201inter12, gate240inter0, gate240inter1, gate240inter2, gate240inter3, gate240inter4, gate240inter5, gate240inter6, gate240inter7, gate240inter8, gate240inter9, gate240inter10, gate240inter11, gate240inter12, gate211inter0, gate211inter1, gate211inter2, gate211inter3, gate211inter4, gate211inter5, gate211inter6, gate211inter7, gate211inter8, gate211inter9, gate211inter10, gate211inter11, gate211inter12, gate287inter0, gate287inter1, gate287inter2, gate287inter3, gate287inter4, gate287inter5, gate287inter6, gate287inter7, gate287inter8, gate287inter9, gate287inter10, gate287inter11, gate287inter12, gate224inter0, gate224inter1, gate224inter2, gate224inter3, gate224inter4, gate224inter5, gate224inter6, gate224inter7, gate224inter8, gate224inter9, gate224inter10, gate224inter11, gate224inter12, gate198inter0, gate198inter1, gate198inter2, gate198inter3, gate198inter4, gate198inter5, gate198inter6, gate198inter7, gate198inter8, gate198inter9, gate198inter10, gate198inter11, gate198inter12, gate414inter0, gate414inter1, gate414inter2, gate414inter3, gate414inter4, gate414inter5, gate414inter6, gate414inter7, gate414inter8, gate414inter9, gate414inter10, gate414inter11, gate414inter12, gate426inter0, gate426inter1, gate426inter2, gate426inter3, gate426inter4, gate426inter5, gate426inter6, gate426inter7, gate426inter8, gate426inter9, gate426inter10, gate426inter11, gate426inter12, gate236inter0, gate236inter1, gate236inter2, gate236inter3, gate236inter4, gate236inter5, gate236inter6, gate236inter7, gate236inter8, gate236inter9, gate236inter10, gate236inter11, gate236inter12, gate162inter0, gate162inter1, gate162inter2, gate162inter3, gate162inter4, gate162inter5, gate162inter6, gate162inter7, gate162inter8, gate162inter9, gate162inter10, gate162inter11, gate162inter12, gate25inter0, gate25inter1, gate25inter2, gate25inter3, gate25inter4, gate25inter5, gate25inter6, gate25inter7, gate25inter8, gate25inter9, gate25inter10, gate25inter11, gate25inter12, gate483inter0, gate483inter1, gate483inter2, gate483inter3, gate483inter4, gate483inter5, gate483inter6, gate483inter7, gate483inter8, gate483inter9, gate483inter10, gate483inter11, gate483inter12, gate212inter0, gate212inter1, gate212inter2, gate212inter3, gate212inter4, gate212inter5, gate212inter6, gate212inter7, gate212inter8, gate212inter9, gate212inter10, gate212inter11, gate212inter12, gate104inter0, gate104inter1, gate104inter2, gate104inter3, gate104inter4, gate104inter5, gate104inter6, gate104inter7, gate104inter8, gate104inter9, gate104inter10, gate104inter11, gate104inter12, gate443inter0, gate443inter1, gate443inter2, gate443inter3, gate443inter4, gate443inter5, gate443inter6, gate443inter7, gate443inter8, gate443inter9, gate443inter10, gate443inter11, gate443inter12, gate55inter0, gate55inter1, gate55inter2, gate55inter3, gate55inter4, gate55inter5, gate55inter6, gate55inter7, gate55inter8, gate55inter9, gate55inter10, gate55inter11, gate55inter12, gate142inter0, gate142inter1, gate142inter2, gate142inter3, gate142inter4, gate142inter5, gate142inter6, gate142inter7, gate142inter8, gate142inter9, gate142inter10, gate142inter11, gate142inter12, gate61inter0, gate61inter1, gate61inter2, gate61inter3, gate61inter4, gate61inter5, gate61inter6, gate61inter7, gate61inter8, gate61inter9, gate61inter10, gate61inter11, gate61inter12, gate482inter0, gate482inter1, gate482inter2, gate482inter3, gate482inter4, gate482inter5, gate482inter6, gate482inter7, gate482inter8, gate482inter9, gate482inter10, gate482inter11, gate482inter12, gate52inter0, gate52inter1, gate52inter2, gate52inter3, gate52inter4, gate52inter5, gate52inter6, gate52inter7, gate52inter8, gate52inter9, gate52inter10, gate52inter11, gate52inter12;



and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );

  xor2  gate1065(.a(G2), .b(G1), .O(gate9inter0));
  nand2 gate1066(.a(gate9inter0), .b(s_74), .O(gate9inter1));
  and2  gate1067(.a(G2), .b(G1), .O(gate9inter2));
  inv1  gate1068(.a(s_74), .O(gate9inter3));
  inv1  gate1069(.a(s_75), .O(gate9inter4));
  nand2 gate1070(.a(gate9inter4), .b(gate9inter3), .O(gate9inter5));
  nor2  gate1071(.a(gate9inter5), .b(gate9inter2), .O(gate9inter6));
  inv1  gate1072(.a(G1), .O(gate9inter7));
  inv1  gate1073(.a(G2), .O(gate9inter8));
  nand2 gate1074(.a(gate9inter8), .b(gate9inter7), .O(gate9inter9));
  nand2 gate1075(.a(s_75), .b(gate9inter3), .O(gate9inter10));
  nor2  gate1076(.a(gate9inter10), .b(gate9inter9), .O(gate9inter11));
  nor2  gate1077(.a(gate9inter11), .b(gate9inter6), .O(gate9inter12));
  nand2 gate1078(.a(gate9inter12), .b(gate9inter1), .O(G266));
nand2 gate10( .a(G3), .b(G4), .O(G269) );
nand2 gate11( .a(G5), .b(G6), .O(G272) );
nand2 gate12( .a(G7), .b(G8), .O(G275) );

  xor2  gate645(.a(G10), .b(G9), .O(gate13inter0));
  nand2 gate646(.a(gate13inter0), .b(s_14), .O(gate13inter1));
  and2  gate647(.a(G10), .b(G9), .O(gate13inter2));
  inv1  gate648(.a(s_14), .O(gate13inter3));
  inv1  gate649(.a(s_15), .O(gate13inter4));
  nand2 gate650(.a(gate13inter4), .b(gate13inter3), .O(gate13inter5));
  nor2  gate651(.a(gate13inter5), .b(gate13inter2), .O(gate13inter6));
  inv1  gate652(.a(G9), .O(gate13inter7));
  inv1  gate653(.a(G10), .O(gate13inter8));
  nand2 gate654(.a(gate13inter8), .b(gate13inter7), .O(gate13inter9));
  nand2 gate655(.a(s_15), .b(gate13inter3), .O(gate13inter10));
  nor2  gate656(.a(gate13inter10), .b(gate13inter9), .O(gate13inter11));
  nor2  gate657(.a(gate13inter11), .b(gate13inter6), .O(gate13inter12));
  nand2 gate658(.a(gate13inter12), .b(gate13inter1), .O(G278));
nand2 gate14( .a(G11), .b(G12), .O(G281) );
nand2 gate15( .a(G13), .b(G14), .O(G284) );
nand2 gate16( .a(G15), .b(G16), .O(G287) );
nand2 gate17( .a(G17), .b(G18), .O(G290) );
nand2 gate18( .a(G19), .b(G20), .O(G293) );

  xor2  gate897(.a(G22), .b(G21), .O(gate19inter0));
  nand2 gate898(.a(gate19inter0), .b(s_50), .O(gate19inter1));
  and2  gate899(.a(G22), .b(G21), .O(gate19inter2));
  inv1  gate900(.a(s_50), .O(gate19inter3));
  inv1  gate901(.a(s_51), .O(gate19inter4));
  nand2 gate902(.a(gate19inter4), .b(gate19inter3), .O(gate19inter5));
  nor2  gate903(.a(gate19inter5), .b(gate19inter2), .O(gate19inter6));
  inv1  gate904(.a(G21), .O(gate19inter7));
  inv1  gate905(.a(G22), .O(gate19inter8));
  nand2 gate906(.a(gate19inter8), .b(gate19inter7), .O(gate19inter9));
  nand2 gate907(.a(s_51), .b(gate19inter3), .O(gate19inter10));
  nor2  gate908(.a(gate19inter10), .b(gate19inter9), .O(gate19inter11));
  nor2  gate909(.a(gate19inter11), .b(gate19inter6), .O(gate19inter12));
  nand2 gate910(.a(gate19inter12), .b(gate19inter1), .O(G296));
nand2 gate20( .a(G23), .b(G24), .O(G299) );
nand2 gate21( .a(G25), .b(G26), .O(G302) );
nand2 gate22( .a(G27), .b(G28), .O(G305) );
nand2 gate23( .a(G29), .b(G30), .O(G308) );
nand2 gate24( .a(G31), .b(G32), .O(G311) );

  xor2  gate1261(.a(G5), .b(G1), .O(gate25inter0));
  nand2 gate1262(.a(gate25inter0), .b(s_102), .O(gate25inter1));
  and2  gate1263(.a(G5), .b(G1), .O(gate25inter2));
  inv1  gate1264(.a(s_102), .O(gate25inter3));
  inv1  gate1265(.a(s_103), .O(gate25inter4));
  nand2 gate1266(.a(gate25inter4), .b(gate25inter3), .O(gate25inter5));
  nor2  gate1267(.a(gate25inter5), .b(gate25inter2), .O(gate25inter6));
  inv1  gate1268(.a(G1), .O(gate25inter7));
  inv1  gate1269(.a(G5), .O(gate25inter8));
  nand2 gate1270(.a(gate25inter8), .b(gate25inter7), .O(gate25inter9));
  nand2 gate1271(.a(s_103), .b(gate25inter3), .O(gate25inter10));
  nor2  gate1272(.a(gate25inter10), .b(gate25inter9), .O(gate25inter11));
  nor2  gate1273(.a(gate25inter11), .b(gate25inter6), .O(gate25inter12));
  nand2 gate1274(.a(gate25inter12), .b(gate25inter1), .O(G314));

  xor2  gate1009(.a(G13), .b(G9), .O(gate26inter0));
  nand2 gate1010(.a(gate26inter0), .b(s_66), .O(gate26inter1));
  and2  gate1011(.a(G13), .b(G9), .O(gate26inter2));
  inv1  gate1012(.a(s_66), .O(gate26inter3));
  inv1  gate1013(.a(s_67), .O(gate26inter4));
  nand2 gate1014(.a(gate26inter4), .b(gate26inter3), .O(gate26inter5));
  nor2  gate1015(.a(gate26inter5), .b(gate26inter2), .O(gate26inter6));
  inv1  gate1016(.a(G9), .O(gate26inter7));
  inv1  gate1017(.a(G13), .O(gate26inter8));
  nand2 gate1018(.a(gate26inter8), .b(gate26inter7), .O(gate26inter9));
  nand2 gate1019(.a(s_67), .b(gate26inter3), .O(gate26inter10));
  nor2  gate1020(.a(gate26inter10), .b(gate26inter9), .O(gate26inter11));
  nor2  gate1021(.a(gate26inter11), .b(gate26inter6), .O(gate26inter12));
  nand2 gate1022(.a(gate26inter12), .b(gate26inter1), .O(G317));
nand2 gate27( .a(G2), .b(G6), .O(G320) );
nand2 gate28( .a(G10), .b(G14), .O(G323) );
nand2 gate29( .a(G3), .b(G7), .O(G326) );
nand2 gate30( .a(G11), .b(G15), .O(G329) );
nand2 gate31( .a(G4), .b(G8), .O(G332) );
nand2 gate32( .a(G12), .b(G16), .O(G335) );
nand2 gate33( .a(G17), .b(G21), .O(G338) );

  xor2  gate1037(.a(G29), .b(G25), .O(gate34inter0));
  nand2 gate1038(.a(gate34inter0), .b(s_70), .O(gate34inter1));
  and2  gate1039(.a(G29), .b(G25), .O(gate34inter2));
  inv1  gate1040(.a(s_70), .O(gate34inter3));
  inv1  gate1041(.a(s_71), .O(gate34inter4));
  nand2 gate1042(.a(gate34inter4), .b(gate34inter3), .O(gate34inter5));
  nor2  gate1043(.a(gate34inter5), .b(gate34inter2), .O(gate34inter6));
  inv1  gate1044(.a(G25), .O(gate34inter7));
  inv1  gate1045(.a(G29), .O(gate34inter8));
  nand2 gate1046(.a(gate34inter8), .b(gate34inter7), .O(gate34inter9));
  nand2 gate1047(.a(s_71), .b(gate34inter3), .O(gate34inter10));
  nor2  gate1048(.a(gate34inter10), .b(gate34inter9), .O(gate34inter11));
  nor2  gate1049(.a(gate34inter11), .b(gate34inter6), .O(gate34inter12));
  nand2 gate1050(.a(gate34inter12), .b(gate34inter1), .O(G341));
nand2 gate35( .a(G18), .b(G22), .O(G344) );
nand2 gate36( .a(G26), .b(G30), .O(G347) );
nand2 gate37( .a(G19), .b(G23), .O(G350) );
nand2 gate38( .a(G27), .b(G31), .O(G353) );
nand2 gate39( .a(G20), .b(G24), .O(G356) );
nand2 gate40( .a(G28), .b(G32), .O(G359) );
nand2 gate41( .a(G1), .b(G266), .O(G362) );
nand2 gate42( .a(G2), .b(G266), .O(G363) );
nand2 gate43( .a(G3), .b(G269), .O(G364) );
nand2 gate44( .a(G4), .b(G269), .O(G365) );
nand2 gate45( .a(G5), .b(G272), .O(G366) );
nand2 gate46( .a(G6), .b(G272), .O(G367) );
nand2 gate47( .a(G7), .b(G275), .O(G368) );
nand2 gate48( .a(G8), .b(G275), .O(G369) );
nand2 gate49( .a(G9), .b(G278), .O(G370) );
nand2 gate50( .a(G10), .b(G278), .O(G371) );
nand2 gate51( .a(G11), .b(G281), .O(G372) );

  xor2  gate1387(.a(G281), .b(G12), .O(gate52inter0));
  nand2 gate1388(.a(gate52inter0), .b(s_120), .O(gate52inter1));
  and2  gate1389(.a(G281), .b(G12), .O(gate52inter2));
  inv1  gate1390(.a(s_120), .O(gate52inter3));
  inv1  gate1391(.a(s_121), .O(gate52inter4));
  nand2 gate1392(.a(gate52inter4), .b(gate52inter3), .O(gate52inter5));
  nor2  gate1393(.a(gate52inter5), .b(gate52inter2), .O(gate52inter6));
  inv1  gate1394(.a(G12), .O(gate52inter7));
  inv1  gate1395(.a(G281), .O(gate52inter8));
  nand2 gate1396(.a(gate52inter8), .b(gate52inter7), .O(gate52inter9));
  nand2 gate1397(.a(s_121), .b(gate52inter3), .O(gate52inter10));
  nor2  gate1398(.a(gate52inter10), .b(gate52inter9), .O(gate52inter11));
  nor2  gate1399(.a(gate52inter11), .b(gate52inter6), .O(gate52inter12));
  nand2 gate1400(.a(gate52inter12), .b(gate52inter1), .O(G373));

  xor2  gate841(.a(G284), .b(G13), .O(gate53inter0));
  nand2 gate842(.a(gate53inter0), .b(s_42), .O(gate53inter1));
  and2  gate843(.a(G284), .b(G13), .O(gate53inter2));
  inv1  gate844(.a(s_42), .O(gate53inter3));
  inv1  gate845(.a(s_43), .O(gate53inter4));
  nand2 gate846(.a(gate53inter4), .b(gate53inter3), .O(gate53inter5));
  nor2  gate847(.a(gate53inter5), .b(gate53inter2), .O(gate53inter6));
  inv1  gate848(.a(G13), .O(gate53inter7));
  inv1  gate849(.a(G284), .O(gate53inter8));
  nand2 gate850(.a(gate53inter8), .b(gate53inter7), .O(gate53inter9));
  nand2 gate851(.a(s_43), .b(gate53inter3), .O(gate53inter10));
  nor2  gate852(.a(gate53inter10), .b(gate53inter9), .O(gate53inter11));
  nor2  gate853(.a(gate53inter11), .b(gate53inter6), .O(gate53inter12));
  nand2 gate854(.a(gate53inter12), .b(gate53inter1), .O(G374));
nand2 gate54( .a(G14), .b(G284), .O(G375) );

  xor2  gate1331(.a(G287), .b(G15), .O(gate55inter0));
  nand2 gate1332(.a(gate55inter0), .b(s_112), .O(gate55inter1));
  and2  gate1333(.a(G287), .b(G15), .O(gate55inter2));
  inv1  gate1334(.a(s_112), .O(gate55inter3));
  inv1  gate1335(.a(s_113), .O(gate55inter4));
  nand2 gate1336(.a(gate55inter4), .b(gate55inter3), .O(gate55inter5));
  nor2  gate1337(.a(gate55inter5), .b(gate55inter2), .O(gate55inter6));
  inv1  gate1338(.a(G15), .O(gate55inter7));
  inv1  gate1339(.a(G287), .O(gate55inter8));
  nand2 gate1340(.a(gate55inter8), .b(gate55inter7), .O(gate55inter9));
  nand2 gate1341(.a(s_113), .b(gate55inter3), .O(gate55inter10));
  nor2  gate1342(.a(gate55inter10), .b(gate55inter9), .O(gate55inter11));
  nor2  gate1343(.a(gate55inter11), .b(gate55inter6), .O(gate55inter12));
  nand2 gate1344(.a(gate55inter12), .b(gate55inter1), .O(G376));
nand2 gate56( .a(G16), .b(G287), .O(G377) );
nand2 gate57( .a(G17), .b(G290), .O(G378) );
nand2 gate58( .a(G18), .b(G290), .O(G379) );
nand2 gate59( .a(G19), .b(G293), .O(G380) );
nand2 gate60( .a(G20), .b(G293), .O(G381) );

  xor2  gate1359(.a(G296), .b(G21), .O(gate61inter0));
  nand2 gate1360(.a(gate61inter0), .b(s_116), .O(gate61inter1));
  and2  gate1361(.a(G296), .b(G21), .O(gate61inter2));
  inv1  gate1362(.a(s_116), .O(gate61inter3));
  inv1  gate1363(.a(s_117), .O(gate61inter4));
  nand2 gate1364(.a(gate61inter4), .b(gate61inter3), .O(gate61inter5));
  nor2  gate1365(.a(gate61inter5), .b(gate61inter2), .O(gate61inter6));
  inv1  gate1366(.a(G21), .O(gate61inter7));
  inv1  gate1367(.a(G296), .O(gate61inter8));
  nand2 gate1368(.a(gate61inter8), .b(gate61inter7), .O(gate61inter9));
  nand2 gate1369(.a(s_117), .b(gate61inter3), .O(gate61inter10));
  nor2  gate1370(.a(gate61inter10), .b(gate61inter9), .O(gate61inter11));
  nor2  gate1371(.a(gate61inter11), .b(gate61inter6), .O(gate61inter12));
  nand2 gate1372(.a(gate61inter12), .b(gate61inter1), .O(G382));
nand2 gate62( .a(G22), .b(G296), .O(G383) );
nand2 gate63( .a(G23), .b(G299), .O(G384) );
nand2 gate64( .a(G24), .b(G299), .O(G385) );

  xor2  gate659(.a(G302), .b(G25), .O(gate65inter0));
  nand2 gate660(.a(gate65inter0), .b(s_16), .O(gate65inter1));
  and2  gate661(.a(G302), .b(G25), .O(gate65inter2));
  inv1  gate662(.a(s_16), .O(gate65inter3));
  inv1  gate663(.a(s_17), .O(gate65inter4));
  nand2 gate664(.a(gate65inter4), .b(gate65inter3), .O(gate65inter5));
  nor2  gate665(.a(gate65inter5), .b(gate65inter2), .O(gate65inter6));
  inv1  gate666(.a(G25), .O(gate65inter7));
  inv1  gate667(.a(G302), .O(gate65inter8));
  nand2 gate668(.a(gate65inter8), .b(gate65inter7), .O(gate65inter9));
  nand2 gate669(.a(s_17), .b(gate65inter3), .O(gate65inter10));
  nor2  gate670(.a(gate65inter10), .b(gate65inter9), .O(gate65inter11));
  nor2  gate671(.a(gate65inter11), .b(gate65inter6), .O(gate65inter12));
  nand2 gate672(.a(gate65inter12), .b(gate65inter1), .O(G386));
nand2 gate66( .a(G26), .b(G302), .O(G387) );
nand2 gate67( .a(G27), .b(G305), .O(G388) );
nand2 gate68( .a(G28), .b(G305), .O(G389) );
nand2 gate69( .a(G29), .b(G308), .O(G390) );
nand2 gate70( .a(G30), .b(G308), .O(G391) );

  xor2  gate981(.a(G311), .b(G31), .O(gate71inter0));
  nand2 gate982(.a(gate71inter0), .b(s_62), .O(gate71inter1));
  and2  gate983(.a(G311), .b(G31), .O(gate71inter2));
  inv1  gate984(.a(s_62), .O(gate71inter3));
  inv1  gate985(.a(s_63), .O(gate71inter4));
  nand2 gate986(.a(gate71inter4), .b(gate71inter3), .O(gate71inter5));
  nor2  gate987(.a(gate71inter5), .b(gate71inter2), .O(gate71inter6));
  inv1  gate988(.a(G31), .O(gate71inter7));
  inv1  gate989(.a(G311), .O(gate71inter8));
  nand2 gate990(.a(gate71inter8), .b(gate71inter7), .O(gate71inter9));
  nand2 gate991(.a(s_63), .b(gate71inter3), .O(gate71inter10));
  nor2  gate992(.a(gate71inter10), .b(gate71inter9), .O(gate71inter11));
  nor2  gate993(.a(gate71inter11), .b(gate71inter6), .O(gate71inter12));
  nand2 gate994(.a(gate71inter12), .b(gate71inter1), .O(G392));
nand2 gate72( .a(G32), .b(G311), .O(G393) );
nand2 gate73( .a(G1), .b(G314), .O(G394) );
nand2 gate74( .a(G5), .b(G314), .O(G395) );
nand2 gate75( .a(G9), .b(G317), .O(G396) );
nand2 gate76( .a(G13), .b(G317), .O(G397) );
nand2 gate77( .a(G2), .b(G320), .O(G398) );
nand2 gate78( .a(G6), .b(G320), .O(G399) );

  xor2  gate925(.a(G323), .b(G10), .O(gate79inter0));
  nand2 gate926(.a(gate79inter0), .b(s_54), .O(gate79inter1));
  and2  gate927(.a(G323), .b(G10), .O(gate79inter2));
  inv1  gate928(.a(s_54), .O(gate79inter3));
  inv1  gate929(.a(s_55), .O(gate79inter4));
  nand2 gate930(.a(gate79inter4), .b(gate79inter3), .O(gate79inter5));
  nor2  gate931(.a(gate79inter5), .b(gate79inter2), .O(gate79inter6));
  inv1  gate932(.a(G10), .O(gate79inter7));
  inv1  gate933(.a(G323), .O(gate79inter8));
  nand2 gate934(.a(gate79inter8), .b(gate79inter7), .O(gate79inter9));
  nand2 gate935(.a(s_55), .b(gate79inter3), .O(gate79inter10));
  nor2  gate936(.a(gate79inter10), .b(gate79inter9), .O(gate79inter11));
  nor2  gate937(.a(gate79inter11), .b(gate79inter6), .O(gate79inter12));
  nand2 gate938(.a(gate79inter12), .b(gate79inter1), .O(G400));
nand2 gate80( .a(G14), .b(G323), .O(G401) );
nand2 gate81( .a(G3), .b(G326), .O(G402) );
nand2 gate82( .a(G7), .b(G326), .O(G403) );
nand2 gate83( .a(G11), .b(G329), .O(G404) );
nand2 gate84( .a(G15), .b(G329), .O(G405) );
nand2 gate85( .a(G4), .b(G332), .O(G406) );
nand2 gate86( .a(G8), .b(G332), .O(G407) );
nand2 gate87( .a(G12), .b(G335), .O(G408) );
nand2 gate88( .a(G16), .b(G335), .O(G409) );
nand2 gate89( .a(G17), .b(G338), .O(G410) );
nand2 gate90( .a(G21), .b(G338), .O(G411) );
nand2 gate91( .a(G25), .b(G341), .O(G412) );
nand2 gate92( .a(G29), .b(G341), .O(G413) );
nand2 gate93( .a(G18), .b(G344), .O(G414) );
nand2 gate94( .a(G22), .b(G344), .O(G415) );
nand2 gate95( .a(G26), .b(G347), .O(G416) );
nand2 gate96( .a(G30), .b(G347), .O(G417) );
nand2 gate97( .a(G19), .b(G350), .O(G418) );
nand2 gate98( .a(G23), .b(G350), .O(G419) );
nand2 gate99( .a(G27), .b(G353), .O(G420) );
nand2 gate100( .a(G31), .b(G353), .O(G421) );
nand2 gate101( .a(G20), .b(G356), .O(G422) );
nand2 gate102( .a(G24), .b(G356), .O(G423) );
nand2 gate103( .a(G28), .b(G359), .O(G424) );

  xor2  gate1303(.a(G359), .b(G32), .O(gate104inter0));
  nand2 gate1304(.a(gate104inter0), .b(s_108), .O(gate104inter1));
  and2  gate1305(.a(G359), .b(G32), .O(gate104inter2));
  inv1  gate1306(.a(s_108), .O(gate104inter3));
  inv1  gate1307(.a(s_109), .O(gate104inter4));
  nand2 gate1308(.a(gate104inter4), .b(gate104inter3), .O(gate104inter5));
  nor2  gate1309(.a(gate104inter5), .b(gate104inter2), .O(gate104inter6));
  inv1  gate1310(.a(G32), .O(gate104inter7));
  inv1  gate1311(.a(G359), .O(gate104inter8));
  nand2 gate1312(.a(gate104inter8), .b(gate104inter7), .O(gate104inter9));
  nand2 gate1313(.a(s_109), .b(gate104inter3), .O(gate104inter10));
  nor2  gate1314(.a(gate104inter10), .b(gate104inter9), .O(gate104inter11));
  nor2  gate1315(.a(gate104inter11), .b(gate104inter6), .O(gate104inter12));
  nand2 gate1316(.a(gate104inter12), .b(gate104inter1), .O(G425));

  xor2  gate687(.a(G363), .b(G362), .O(gate105inter0));
  nand2 gate688(.a(gate105inter0), .b(s_20), .O(gate105inter1));
  and2  gate689(.a(G363), .b(G362), .O(gate105inter2));
  inv1  gate690(.a(s_20), .O(gate105inter3));
  inv1  gate691(.a(s_21), .O(gate105inter4));
  nand2 gate692(.a(gate105inter4), .b(gate105inter3), .O(gate105inter5));
  nor2  gate693(.a(gate105inter5), .b(gate105inter2), .O(gate105inter6));
  inv1  gate694(.a(G362), .O(gate105inter7));
  inv1  gate695(.a(G363), .O(gate105inter8));
  nand2 gate696(.a(gate105inter8), .b(gate105inter7), .O(gate105inter9));
  nand2 gate697(.a(s_21), .b(gate105inter3), .O(gate105inter10));
  nor2  gate698(.a(gate105inter10), .b(gate105inter9), .O(gate105inter11));
  nor2  gate699(.a(gate105inter11), .b(gate105inter6), .O(gate105inter12));
  nand2 gate700(.a(gate105inter12), .b(gate105inter1), .O(G426));
nand2 gate106( .a(G364), .b(G365), .O(G429) );
nand2 gate107( .a(G366), .b(G367), .O(G432) );
nand2 gate108( .a(G368), .b(G369), .O(G435) );
nand2 gate109( .a(G370), .b(G371), .O(G438) );
nand2 gate110( .a(G372), .b(G373), .O(G441) );
nand2 gate111( .a(G374), .b(G375), .O(G444) );
nand2 gate112( .a(G376), .b(G377), .O(G447) );
nand2 gate113( .a(G378), .b(G379), .O(G450) );
nand2 gate114( .a(G380), .b(G381), .O(G453) );
nand2 gate115( .a(G382), .b(G383), .O(G456) );
nand2 gate116( .a(G384), .b(G385), .O(G459) );
nand2 gate117( .a(G386), .b(G387), .O(G462) );
nand2 gate118( .a(G388), .b(G389), .O(G465) );

  xor2  gate967(.a(G391), .b(G390), .O(gate119inter0));
  nand2 gate968(.a(gate119inter0), .b(s_60), .O(gate119inter1));
  and2  gate969(.a(G391), .b(G390), .O(gate119inter2));
  inv1  gate970(.a(s_60), .O(gate119inter3));
  inv1  gate971(.a(s_61), .O(gate119inter4));
  nand2 gate972(.a(gate119inter4), .b(gate119inter3), .O(gate119inter5));
  nor2  gate973(.a(gate119inter5), .b(gate119inter2), .O(gate119inter6));
  inv1  gate974(.a(G390), .O(gate119inter7));
  inv1  gate975(.a(G391), .O(gate119inter8));
  nand2 gate976(.a(gate119inter8), .b(gate119inter7), .O(gate119inter9));
  nand2 gate977(.a(s_61), .b(gate119inter3), .O(gate119inter10));
  nor2  gate978(.a(gate119inter10), .b(gate119inter9), .O(gate119inter11));
  nor2  gate979(.a(gate119inter11), .b(gate119inter6), .O(gate119inter12));
  nand2 gate980(.a(gate119inter12), .b(gate119inter1), .O(G468));
nand2 gate120( .a(G392), .b(G393), .O(G471) );
nand2 gate121( .a(G394), .b(G395), .O(G474) );
nand2 gate122( .a(G396), .b(G397), .O(G477) );
nand2 gate123( .a(G398), .b(G399), .O(G480) );
nand2 gate124( .a(G400), .b(G401), .O(G483) );
nand2 gate125( .a(G402), .b(G403), .O(G486) );
nand2 gate126( .a(G404), .b(G405), .O(G489) );
nand2 gate127( .a(G406), .b(G407), .O(G492) );

  xor2  gate673(.a(G409), .b(G408), .O(gate128inter0));
  nand2 gate674(.a(gate128inter0), .b(s_18), .O(gate128inter1));
  and2  gate675(.a(G409), .b(G408), .O(gate128inter2));
  inv1  gate676(.a(s_18), .O(gate128inter3));
  inv1  gate677(.a(s_19), .O(gate128inter4));
  nand2 gate678(.a(gate128inter4), .b(gate128inter3), .O(gate128inter5));
  nor2  gate679(.a(gate128inter5), .b(gate128inter2), .O(gate128inter6));
  inv1  gate680(.a(G408), .O(gate128inter7));
  inv1  gate681(.a(G409), .O(gate128inter8));
  nand2 gate682(.a(gate128inter8), .b(gate128inter7), .O(gate128inter9));
  nand2 gate683(.a(s_19), .b(gate128inter3), .O(gate128inter10));
  nor2  gate684(.a(gate128inter10), .b(gate128inter9), .O(gate128inter11));
  nor2  gate685(.a(gate128inter11), .b(gate128inter6), .O(gate128inter12));
  nand2 gate686(.a(gate128inter12), .b(gate128inter1), .O(G495));
nand2 gate129( .a(G410), .b(G411), .O(G498) );
nand2 gate130( .a(G412), .b(G413), .O(G501) );
nand2 gate131( .a(G414), .b(G415), .O(G504) );
nand2 gate132( .a(G416), .b(G417), .O(G507) );
nand2 gate133( .a(G418), .b(G419), .O(G510) );
nand2 gate134( .a(G420), .b(G421), .O(G513) );

  xor2  gate771(.a(G423), .b(G422), .O(gate135inter0));
  nand2 gate772(.a(gate135inter0), .b(s_32), .O(gate135inter1));
  and2  gate773(.a(G423), .b(G422), .O(gate135inter2));
  inv1  gate774(.a(s_32), .O(gate135inter3));
  inv1  gate775(.a(s_33), .O(gate135inter4));
  nand2 gate776(.a(gate135inter4), .b(gate135inter3), .O(gate135inter5));
  nor2  gate777(.a(gate135inter5), .b(gate135inter2), .O(gate135inter6));
  inv1  gate778(.a(G422), .O(gate135inter7));
  inv1  gate779(.a(G423), .O(gate135inter8));
  nand2 gate780(.a(gate135inter8), .b(gate135inter7), .O(gate135inter9));
  nand2 gate781(.a(s_33), .b(gate135inter3), .O(gate135inter10));
  nor2  gate782(.a(gate135inter10), .b(gate135inter9), .O(gate135inter11));
  nor2  gate783(.a(gate135inter11), .b(gate135inter6), .O(gate135inter12));
  nand2 gate784(.a(gate135inter12), .b(gate135inter1), .O(G516));
nand2 gate136( .a(G424), .b(G425), .O(G519) );
nand2 gate137( .a(G426), .b(G429), .O(G522) );
nand2 gate138( .a(G432), .b(G435), .O(G525) );
nand2 gate139( .a(G438), .b(G441), .O(G528) );
nand2 gate140( .a(G444), .b(G447), .O(G531) );
nand2 gate141( .a(G450), .b(G453), .O(G534) );

  xor2  gate1345(.a(G459), .b(G456), .O(gate142inter0));
  nand2 gate1346(.a(gate142inter0), .b(s_114), .O(gate142inter1));
  and2  gate1347(.a(G459), .b(G456), .O(gate142inter2));
  inv1  gate1348(.a(s_114), .O(gate142inter3));
  inv1  gate1349(.a(s_115), .O(gate142inter4));
  nand2 gate1350(.a(gate142inter4), .b(gate142inter3), .O(gate142inter5));
  nor2  gate1351(.a(gate142inter5), .b(gate142inter2), .O(gate142inter6));
  inv1  gate1352(.a(G456), .O(gate142inter7));
  inv1  gate1353(.a(G459), .O(gate142inter8));
  nand2 gate1354(.a(gate142inter8), .b(gate142inter7), .O(gate142inter9));
  nand2 gate1355(.a(s_115), .b(gate142inter3), .O(gate142inter10));
  nor2  gate1356(.a(gate142inter10), .b(gate142inter9), .O(gate142inter11));
  nor2  gate1357(.a(gate142inter11), .b(gate142inter6), .O(gate142inter12));
  nand2 gate1358(.a(gate142inter12), .b(gate142inter1), .O(G537));

  xor2  gate883(.a(G465), .b(G462), .O(gate143inter0));
  nand2 gate884(.a(gate143inter0), .b(s_48), .O(gate143inter1));
  and2  gate885(.a(G465), .b(G462), .O(gate143inter2));
  inv1  gate886(.a(s_48), .O(gate143inter3));
  inv1  gate887(.a(s_49), .O(gate143inter4));
  nand2 gate888(.a(gate143inter4), .b(gate143inter3), .O(gate143inter5));
  nor2  gate889(.a(gate143inter5), .b(gate143inter2), .O(gate143inter6));
  inv1  gate890(.a(G462), .O(gate143inter7));
  inv1  gate891(.a(G465), .O(gate143inter8));
  nand2 gate892(.a(gate143inter8), .b(gate143inter7), .O(gate143inter9));
  nand2 gate893(.a(s_49), .b(gate143inter3), .O(gate143inter10));
  nor2  gate894(.a(gate143inter10), .b(gate143inter9), .O(gate143inter11));
  nor2  gate895(.a(gate143inter11), .b(gate143inter6), .O(gate143inter12));
  nand2 gate896(.a(gate143inter12), .b(gate143inter1), .O(G540));
nand2 gate144( .a(G468), .b(G471), .O(G543) );
nand2 gate145( .a(G474), .b(G477), .O(G546) );
nand2 gate146( .a(G480), .b(G483), .O(G549) );
nand2 gate147( .a(G486), .b(G489), .O(G552) );
nand2 gate148( .a(G492), .b(G495), .O(G555) );
nand2 gate149( .a(G498), .b(G501), .O(G558) );
nand2 gate150( .a(G504), .b(G507), .O(G561) );
nand2 gate151( .a(G510), .b(G513), .O(G564) );
nand2 gate152( .a(G516), .b(G519), .O(G567) );
nand2 gate153( .a(G426), .b(G522), .O(G570) );
nand2 gate154( .a(G429), .b(G522), .O(G571) );
nand2 gate155( .a(G432), .b(G525), .O(G572) );
nand2 gate156( .a(G435), .b(G525), .O(G573) );
nand2 gate157( .a(G438), .b(G528), .O(G574) );
nand2 gate158( .a(G441), .b(G528), .O(G575) );
nand2 gate159( .a(G444), .b(G531), .O(G576) );
nand2 gate160( .a(G447), .b(G531), .O(G577) );
nand2 gate161( .a(G450), .b(G534), .O(G578) );

  xor2  gate1247(.a(G534), .b(G453), .O(gate162inter0));
  nand2 gate1248(.a(gate162inter0), .b(s_100), .O(gate162inter1));
  and2  gate1249(.a(G534), .b(G453), .O(gate162inter2));
  inv1  gate1250(.a(s_100), .O(gate162inter3));
  inv1  gate1251(.a(s_101), .O(gate162inter4));
  nand2 gate1252(.a(gate162inter4), .b(gate162inter3), .O(gate162inter5));
  nor2  gate1253(.a(gate162inter5), .b(gate162inter2), .O(gate162inter6));
  inv1  gate1254(.a(G453), .O(gate162inter7));
  inv1  gate1255(.a(G534), .O(gate162inter8));
  nand2 gate1256(.a(gate162inter8), .b(gate162inter7), .O(gate162inter9));
  nand2 gate1257(.a(s_101), .b(gate162inter3), .O(gate162inter10));
  nor2  gate1258(.a(gate162inter10), .b(gate162inter9), .O(gate162inter11));
  nor2  gate1259(.a(gate162inter11), .b(gate162inter6), .O(gate162inter12));
  nand2 gate1260(.a(gate162inter12), .b(gate162inter1), .O(G579));
nand2 gate163( .a(G456), .b(G537), .O(G580) );
nand2 gate164( .a(G459), .b(G537), .O(G581) );
nand2 gate165( .a(G462), .b(G540), .O(G582) );
nand2 gate166( .a(G465), .b(G540), .O(G583) );
nand2 gate167( .a(G468), .b(G543), .O(G584) );
nand2 gate168( .a(G471), .b(G543), .O(G585) );
nand2 gate169( .a(G474), .b(G546), .O(G586) );
nand2 gate170( .a(G477), .b(G546), .O(G587) );

  xor2  gate827(.a(G549), .b(G480), .O(gate171inter0));
  nand2 gate828(.a(gate171inter0), .b(s_40), .O(gate171inter1));
  and2  gate829(.a(G549), .b(G480), .O(gate171inter2));
  inv1  gate830(.a(s_40), .O(gate171inter3));
  inv1  gate831(.a(s_41), .O(gate171inter4));
  nand2 gate832(.a(gate171inter4), .b(gate171inter3), .O(gate171inter5));
  nor2  gate833(.a(gate171inter5), .b(gate171inter2), .O(gate171inter6));
  inv1  gate834(.a(G480), .O(gate171inter7));
  inv1  gate835(.a(G549), .O(gate171inter8));
  nand2 gate836(.a(gate171inter8), .b(gate171inter7), .O(gate171inter9));
  nand2 gate837(.a(s_41), .b(gate171inter3), .O(gate171inter10));
  nor2  gate838(.a(gate171inter10), .b(gate171inter9), .O(gate171inter11));
  nor2  gate839(.a(gate171inter11), .b(gate171inter6), .O(gate171inter12));
  nand2 gate840(.a(gate171inter12), .b(gate171inter1), .O(G588));
nand2 gate172( .a(G483), .b(G549), .O(G589) );
nand2 gate173( .a(G486), .b(G552), .O(G590) );
nand2 gate174( .a(G489), .b(G552), .O(G591) );
nand2 gate175( .a(G492), .b(G555), .O(G592) );

  xor2  gate729(.a(G555), .b(G495), .O(gate176inter0));
  nand2 gate730(.a(gate176inter0), .b(s_26), .O(gate176inter1));
  and2  gate731(.a(G555), .b(G495), .O(gate176inter2));
  inv1  gate732(.a(s_26), .O(gate176inter3));
  inv1  gate733(.a(s_27), .O(gate176inter4));
  nand2 gate734(.a(gate176inter4), .b(gate176inter3), .O(gate176inter5));
  nor2  gate735(.a(gate176inter5), .b(gate176inter2), .O(gate176inter6));
  inv1  gate736(.a(G495), .O(gate176inter7));
  inv1  gate737(.a(G555), .O(gate176inter8));
  nand2 gate738(.a(gate176inter8), .b(gate176inter7), .O(gate176inter9));
  nand2 gate739(.a(s_27), .b(gate176inter3), .O(gate176inter10));
  nor2  gate740(.a(gate176inter10), .b(gate176inter9), .O(gate176inter11));
  nor2  gate741(.a(gate176inter11), .b(gate176inter6), .O(gate176inter12));
  nand2 gate742(.a(gate176inter12), .b(gate176inter1), .O(G593));

  xor2  gate911(.a(G558), .b(G498), .O(gate177inter0));
  nand2 gate912(.a(gate177inter0), .b(s_52), .O(gate177inter1));
  and2  gate913(.a(G558), .b(G498), .O(gate177inter2));
  inv1  gate914(.a(s_52), .O(gate177inter3));
  inv1  gate915(.a(s_53), .O(gate177inter4));
  nand2 gate916(.a(gate177inter4), .b(gate177inter3), .O(gate177inter5));
  nor2  gate917(.a(gate177inter5), .b(gate177inter2), .O(gate177inter6));
  inv1  gate918(.a(G498), .O(gate177inter7));
  inv1  gate919(.a(G558), .O(gate177inter8));
  nand2 gate920(.a(gate177inter8), .b(gate177inter7), .O(gate177inter9));
  nand2 gate921(.a(s_53), .b(gate177inter3), .O(gate177inter10));
  nor2  gate922(.a(gate177inter10), .b(gate177inter9), .O(gate177inter11));
  nor2  gate923(.a(gate177inter11), .b(gate177inter6), .O(gate177inter12));
  nand2 gate924(.a(gate177inter12), .b(gate177inter1), .O(G594));
nand2 gate178( .a(G501), .b(G558), .O(G595) );
nand2 gate179( .a(G504), .b(G561), .O(G596) );
nand2 gate180( .a(G507), .b(G561), .O(G597) );
nand2 gate181( .a(G510), .b(G564), .O(G598) );
nand2 gate182( .a(G513), .b(G564), .O(G599) );
nand2 gate183( .a(G516), .b(G567), .O(G600) );
nand2 gate184( .a(G519), .b(G567), .O(G601) );
nand2 gate185( .a(G570), .b(G571), .O(G602) );
nand2 gate186( .a(G572), .b(G573), .O(G607) );
nand2 gate187( .a(G574), .b(G575), .O(G612) );
nand2 gate188( .a(G576), .b(G577), .O(G617) );
nand2 gate189( .a(G578), .b(G579), .O(G622) );
nand2 gate190( .a(G580), .b(G581), .O(G627) );
nand2 gate191( .a(G582), .b(G583), .O(G632) );
nand2 gate192( .a(G584), .b(G585), .O(G637) );
nand2 gate193( .a(G586), .b(G587), .O(G642) );

  xor2  gate547(.a(G589), .b(G588), .O(gate194inter0));
  nand2 gate548(.a(gate194inter0), .b(s_0), .O(gate194inter1));
  and2  gate549(.a(G589), .b(G588), .O(gate194inter2));
  inv1  gate550(.a(s_0), .O(gate194inter3));
  inv1  gate551(.a(s_1), .O(gate194inter4));
  nand2 gate552(.a(gate194inter4), .b(gate194inter3), .O(gate194inter5));
  nor2  gate553(.a(gate194inter5), .b(gate194inter2), .O(gate194inter6));
  inv1  gate554(.a(G588), .O(gate194inter7));
  inv1  gate555(.a(G589), .O(gate194inter8));
  nand2 gate556(.a(gate194inter8), .b(gate194inter7), .O(gate194inter9));
  nand2 gate557(.a(s_1), .b(gate194inter3), .O(gate194inter10));
  nor2  gate558(.a(gate194inter10), .b(gate194inter9), .O(gate194inter11));
  nor2  gate559(.a(gate194inter11), .b(gate194inter6), .O(gate194inter12));
  nand2 gate560(.a(gate194inter12), .b(gate194inter1), .O(G645));
nand2 gate195( .a(G590), .b(G591), .O(G648) );
nand2 gate196( .a(G592), .b(G593), .O(G651) );
nand2 gate197( .a(G594), .b(G595), .O(G654) );

  xor2  gate1191(.a(G597), .b(G596), .O(gate198inter0));
  nand2 gate1192(.a(gate198inter0), .b(s_92), .O(gate198inter1));
  and2  gate1193(.a(G597), .b(G596), .O(gate198inter2));
  inv1  gate1194(.a(s_92), .O(gate198inter3));
  inv1  gate1195(.a(s_93), .O(gate198inter4));
  nand2 gate1196(.a(gate198inter4), .b(gate198inter3), .O(gate198inter5));
  nor2  gate1197(.a(gate198inter5), .b(gate198inter2), .O(gate198inter6));
  inv1  gate1198(.a(G596), .O(gate198inter7));
  inv1  gate1199(.a(G597), .O(gate198inter8));
  nand2 gate1200(.a(gate198inter8), .b(gate198inter7), .O(gate198inter9));
  nand2 gate1201(.a(s_93), .b(gate198inter3), .O(gate198inter10));
  nor2  gate1202(.a(gate198inter10), .b(gate198inter9), .O(gate198inter11));
  nor2  gate1203(.a(gate198inter11), .b(gate198inter6), .O(gate198inter12));
  nand2 gate1204(.a(gate198inter12), .b(gate198inter1), .O(G657));
nand2 gate199( .a(G598), .b(G599), .O(G660) );
nand2 gate200( .a(G600), .b(G601), .O(G663) );

  xor2  gate1121(.a(G607), .b(G602), .O(gate201inter0));
  nand2 gate1122(.a(gate201inter0), .b(s_82), .O(gate201inter1));
  and2  gate1123(.a(G607), .b(G602), .O(gate201inter2));
  inv1  gate1124(.a(s_82), .O(gate201inter3));
  inv1  gate1125(.a(s_83), .O(gate201inter4));
  nand2 gate1126(.a(gate201inter4), .b(gate201inter3), .O(gate201inter5));
  nor2  gate1127(.a(gate201inter5), .b(gate201inter2), .O(gate201inter6));
  inv1  gate1128(.a(G602), .O(gate201inter7));
  inv1  gate1129(.a(G607), .O(gate201inter8));
  nand2 gate1130(.a(gate201inter8), .b(gate201inter7), .O(gate201inter9));
  nand2 gate1131(.a(s_83), .b(gate201inter3), .O(gate201inter10));
  nor2  gate1132(.a(gate201inter10), .b(gate201inter9), .O(gate201inter11));
  nor2  gate1133(.a(gate201inter11), .b(gate201inter6), .O(gate201inter12));
  nand2 gate1134(.a(gate201inter12), .b(gate201inter1), .O(G666));
nand2 gate202( .a(G612), .b(G617), .O(G669) );
nand2 gate203( .a(G602), .b(G612), .O(G672) );
nand2 gate204( .a(G607), .b(G617), .O(G675) );
nand2 gate205( .a(G622), .b(G627), .O(G678) );
nand2 gate206( .a(G632), .b(G637), .O(G681) );
nand2 gate207( .a(G622), .b(G632), .O(G684) );
nand2 gate208( .a(G627), .b(G637), .O(G687) );
nand2 gate209( .a(G602), .b(G666), .O(G690) );
nand2 gate210( .a(G607), .b(G666), .O(G691) );

  xor2  gate1149(.a(G669), .b(G612), .O(gate211inter0));
  nand2 gate1150(.a(gate211inter0), .b(s_86), .O(gate211inter1));
  and2  gate1151(.a(G669), .b(G612), .O(gate211inter2));
  inv1  gate1152(.a(s_86), .O(gate211inter3));
  inv1  gate1153(.a(s_87), .O(gate211inter4));
  nand2 gate1154(.a(gate211inter4), .b(gate211inter3), .O(gate211inter5));
  nor2  gate1155(.a(gate211inter5), .b(gate211inter2), .O(gate211inter6));
  inv1  gate1156(.a(G612), .O(gate211inter7));
  inv1  gate1157(.a(G669), .O(gate211inter8));
  nand2 gate1158(.a(gate211inter8), .b(gate211inter7), .O(gate211inter9));
  nand2 gate1159(.a(s_87), .b(gate211inter3), .O(gate211inter10));
  nor2  gate1160(.a(gate211inter10), .b(gate211inter9), .O(gate211inter11));
  nor2  gate1161(.a(gate211inter11), .b(gate211inter6), .O(gate211inter12));
  nand2 gate1162(.a(gate211inter12), .b(gate211inter1), .O(G692));

  xor2  gate1289(.a(G669), .b(G617), .O(gate212inter0));
  nand2 gate1290(.a(gate212inter0), .b(s_106), .O(gate212inter1));
  and2  gate1291(.a(G669), .b(G617), .O(gate212inter2));
  inv1  gate1292(.a(s_106), .O(gate212inter3));
  inv1  gate1293(.a(s_107), .O(gate212inter4));
  nand2 gate1294(.a(gate212inter4), .b(gate212inter3), .O(gate212inter5));
  nor2  gate1295(.a(gate212inter5), .b(gate212inter2), .O(gate212inter6));
  inv1  gate1296(.a(G617), .O(gate212inter7));
  inv1  gate1297(.a(G669), .O(gate212inter8));
  nand2 gate1298(.a(gate212inter8), .b(gate212inter7), .O(gate212inter9));
  nand2 gate1299(.a(s_107), .b(gate212inter3), .O(gate212inter10));
  nor2  gate1300(.a(gate212inter10), .b(gate212inter9), .O(gate212inter11));
  nor2  gate1301(.a(gate212inter11), .b(gate212inter6), .O(gate212inter12));
  nand2 gate1302(.a(gate212inter12), .b(gate212inter1), .O(G693));
nand2 gate213( .a(G602), .b(G672), .O(G694) );
nand2 gate214( .a(G612), .b(G672), .O(G695) );

  xor2  gate1107(.a(G675), .b(G607), .O(gate215inter0));
  nand2 gate1108(.a(gate215inter0), .b(s_80), .O(gate215inter1));
  and2  gate1109(.a(G675), .b(G607), .O(gate215inter2));
  inv1  gate1110(.a(s_80), .O(gate215inter3));
  inv1  gate1111(.a(s_81), .O(gate215inter4));
  nand2 gate1112(.a(gate215inter4), .b(gate215inter3), .O(gate215inter5));
  nor2  gate1113(.a(gate215inter5), .b(gate215inter2), .O(gate215inter6));
  inv1  gate1114(.a(G607), .O(gate215inter7));
  inv1  gate1115(.a(G675), .O(gate215inter8));
  nand2 gate1116(.a(gate215inter8), .b(gate215inter7), .O(gate215inter9));
  nand2 gate1117(.a(s_81), .b(gate215inter3), .O(gate215inter10));
  nor2  gate1118(.a(gate215inter10), .b(gate215inter9), .O(gate215inter11));
  nor2  gate1119(.a(gate215inter11), .b(gate215inter6), .O(gate215inter12));
  nand2 gate1120(.a(gate215inter12), .b(gate215inter1), .O(G696));
nand2 gate216( .a(G617), .b(G675), .O(G697) );
nand2 gate217( .a(G622), .b(G678), .O(G698) );
nand2 gate218( .a(G627), .b(G678), .O(G699) );
nand2 gate219( .a(G632), .b(G681), .O(G700) );
nand2 gate220( .a(G637), .b(G681), .O(G701) );
nand2 gate221( .a(G622), .b(G684), .O(G702) );
nand2 gate222( .a(G632), .b(G684), .O(G703) );
nand2 gate223( .a(G627), .b(G687), .O(G704) );

  xor2  gate1177(.a(G687), .b(G637), .O(gate224inter0));
  nand2 gate1178(.a(gate224inter0), .b(s_90), .O(gate224inter1));
  and2  gate1179(.a(G687), .b(G637), .O(gate224inter2));
  inv1  gate1180(.a(s_90), .O(gate224inter3));
  inv1  gate1181(.a(s_91), .O(gate224inter4));
  nand2 gate1182(.a(gate224inter4), .b(gate224inter3), .O(gate224inter5));
  nor2  gate1183(.a(gate224inter5), .b(gate224inter2), .O(gate224inter6));
  inv1  gate1184(.a(G637), .O(gate224inter7));
  inv1  gate1185(.a(G687), .O(gate224inter8));
  nand2 gate1186(.a(gate224inter8), .b(gate224inter7), .O(gate224inter9));
  nand2 gate1187(.a(s_91), .b(gate224inter3), .O(gate224inter10));
  nor2  gate1188(.a(gate224inter10), .b(gate224inter9), .O(gate224inter11));
  nor2  gate1189(.a(gate224inter11), .b(gate224inter6), .O(gate224inter12));
  nand2 gate1190(.a(gate224inter12), .b(gate224inter1), .O(G705));
nand2 gate225( .a(G690), .b(G691), .O(G706) );
nand2 gate226( .a(G692), .b(G693), .O(G709) );
nand2 gate227( .a(G694), .b(G695), .O(G712) );
nand2 gate228( .a(G696), .b(G697), .O(G715) );
nand2 gate229( .a(G698), .b(G699), .O(G718) );
nand2 gate230( .a(G700), .b(G701), .O(G721) );
nand2 gate231( .a(G702), .b(G703), .O(G724) );
nand2 gate232( .a(G704), .b(G705), .O(G727) );
nand2 gate233( .a(G242), .b(G718), .O(G730) );
nand2 gate234( .a(G245), .b(G721), .O(G733) );
nand2 gate235( .a(G248), .b(G724), .O(G736) );

  xor2  gate1233(.a(G727), .b(G251), .O(gate236inter0));
  nand2 gate1234(.a(gate236inter0), .b(s_98), .O(gate236inter1));
  and2  gate1235(.a(G727), .b(G251), .O(gate236inter2));
  inv1  gate1236(.a(s_98), .O(gate236inter3));
  inv1  gate1237(.a(s_99), .O(gate236inter4));
  nand2 gate1238(.a(gate236inter4), .b(gate236inter3), .O(gate236inter5));
  nor2  gate1239(.a(gate236inter5), .b(gate236inter2), .O(gate236inter6));
  inv1  gate1240(.a(G251), .O(gate236inter7));
  inv1  gate1241(.a(G727), .O(gate236inter8));
  nand2 gate1242(.a(gate236inter8), .b(gate236inter7), .O(gate236inter9));
  nand2 gate1243(.a(s_99), .b(gate236inter3), .O(gate236inter10));
  nor2  gate1244(.a(gate236inter10), .b(gate236inter9), .O(gate236inter11));
  nor2  gate1245(.a(gate236inter11), .b(gate236inter6), .O(gate236inter12));
  nand2 gate1246(.a(gate236inter12), .b(gate236inter1), .O(G739));
nand2 gate237( .a(G254), .b(G706), .O(G742) );
nand2 gate238( .a(G257), .b(G709), .O(G745) );
nand2 gate239( .a(G260), .b(G712), .O(G748) );

  xor2  gate1135(.a(G715), .b(G263), .O(gate240inter0));
  nand2 gate1136(.a(gate240inter0), .b(s_84), .O(gate240inter1));
  and2  gate1137(.a(G715), .b(G263), .O(gate240inter2));
  inv1  gate1138(.a(s_84), .O(gate240inter3));
  inv1  gate1139(.a(s_85), .O(gate240inter4));
  nand2 gate1140(.a(gate240inter4), .b(gate240inter3), .O(gate240inter5));
  nor2  gate1141(.a(gate240inter5), .b(gate240inter2), .O(gate240inter6));
  inv1  gate1142(.a(G263), .O(gate240inter7));
  inv1  gate1143(.a(G715), .O(gate240inter8));
  nand2 gate1144(.a(gate240inter8), .b(gate240inter7), .O(gate240inter9));
  nand2 gate1145(.a(s_85), .b(gate240inter3), .O(gate240inter10));
  nor2  gate1146(.a(gate240inter10), .b(gate240inter9), .O(gate240inter11));
  nor2  gate1147(.a(gate240inter11), .b(gate240inter6), .O(gate240inter12));
  nand2 gate1148(.a(gate240inter12), .b(gate240inter1), .O(G751));
nand2 gate241( .a(G242), .b(G730), .O(G754) );
nand2 gate242( .a(G718), .b(G730), .O(G755) );

  xor2  gate701(.a(G733), .b(G245), .O(gate243inter0));
  nand2 gate702(.a(gate243inter0), .b(s_22), .O(gate243inter1));
  and2  gate703(.a(G733), .b(G245), .O(gate243inter2));
  inv1  gate704(.a(s_22), .O(gate243inter3));
  inv1  gate705(.a(s_23), .O(gate243inter4));
  nand2 gate706(.a(gate243inter4), .b(gate243inter3), .O(gate243inter5));
  nor2  gate707(.a(gate243inter5), .b(gate243inter2), .O(gate243inter6));
  inv1  gate708(.a(G245), .O(gate243inter7));
  inv1  gate709(.a(G733), .O(gate243inter8));
  nand2 gate710(.a(gate243inter8), .b(gate243inter7), .O(gate243inter9));
  nand2 gate711(.a(s_23), .b(gate243inter3), .O(gate243inter10));
  nor2  gate712(.a(gate243inter10), .b(gate243inter9), .O(gate243inter11));
  nor2  gate713(.a(gate243inter11), .b(gate243inter6), .O(gate243inter12));
  nand2 gate714(.a(gate243inter12), .b(gate243inter1), .O(G756));

  xor2  gate617(.a(G733), .b(G721), .O(gate244inter0));
  nand2 gate618(.a(gate244inter0), .b(s_10), .O(gate244inter1));
  and2  gate619(.a(G733), .b(G721), .O(gate244inter2));
  inv1  gate620(.a(s_10), .O(gate244inter3));
  inv1  gate621(.a(s_11), .O(gate244inter4));
  nand2 gate622(.a(gate244inter4), .b(gate244inter3), .O(gate244inter5));
  nor2  gate623(.a(gate244inter5), .b(gate244inter2), .O(gate244inter6));
  inv1  gate624(.a(G721), .O(gate244inter7));
  inv1  gate625(.a(G733), .O(gate244inter8));
  nand2 gate626(.a(gate244inter8), .b(gate244inter7), .O(gate244inter9));
  nand2 gate627(.a(s_11), .b(gate244inter3), .O(gate244inter10));
  nor2  gate628(.a(gate244inter10), .b(gate244inter9), .O(gate244inter11));
  nor2  gate629(.a(gate244inter11), .b(gate244inter6), .O(gate244inter12));
  nand2 gate630(.a(gate244inter12), .b(gate244inter1), .O(G757));
nand2 gate245( .a(G248), .b(G736), .O(G758) );
nand2 gate246( .a(G724), .b(G736), .O(G759) );
nand2 gate247( .a(G251), .b(G739), .O(G760) );
nand2 gate248( .a(G727), .b(G739), .O(G761) );
nand2 gate249( .a(G254), .b(G742), .O(G762) );
nand2 gate250( .a(G706), .b(G742), .O(G763) );
nand2 gate251( .a(G257), .b(G745), .O(G764) );
nand2 gate252( .a(G709), .b(G745), .O(G765) );

  xor2  gate757(.a(G748), .b(G260), .O(gate253inter0));
  nand2 gate758(.a(gate253inter0), .b(s_30), .O(gate253inter1));
  and2  gate759(.a(G748), .b(G260), .O(gate253inter2));
  inv1  gate760(.a(s_30), .O(gate253inter3));
  inv1  gate761(.a(s_31), .O(gate253inter4));
  nand2 gate762(.a(gate253inter4), .b(gate253inter3), .O(gate253inter5));
  nor2  gate763(.a(gate253inter5), .b(gate253inter2), .O(gate253inter6));
  inv1  gate764(.a(G260), .O(gate253inter7));
  inv1  gate765(.a(G748), .O(gate253inter8));
  nand2 gate766(.a(gate253inter8), .b(gate253inter7), .O(gate253inter9));
  nand2 gate767(.a(s_31), .b(gate253inter3), .O(gate253inter10));
  nor2  gate768(.a(gate253inter10), .b(gate253inter9), .O(gate253inter11));
  nor2  gate769(.a(gate253inter11), .b(gate253inter6), .O(gate253inter12));
  nand2 gate770(.a(gate253inter12), .b(gate253inter1), .O(G766));
nand2 gate254( .a(G712), .b(G748), .O(G767) );
nand2 gate255( .a(G263), .b(G751), .O(G768) );

  xor2  gate575(.a(G751), .b(G715), .O(gate256inter0));
  nand2 gate576(.a(gate256inter0), .b(s_4), .O(gate256inter1));
  and2  gate577(.a(G751), .b(G715), .O(gate256inter2));
  inv1  gate578(.a(s_4), .O(gate256inter3));
  inv1  gate579(.a(s_5), .O(gate256inter4));
  nand2 gate580(.a(gate256inter4), .b(gate256inter3), .O(gate256inter5));
  nor2  gate581(.a(gate256inter5), .b(gate256inter2), .O(gate256inter6));
  inv1  gate582(.a(G715), .O(gate256inter7));
  inv1  gate583(.a(G751), .O(gate256inter8));
  nand2 gate584(.a(gate256inter8), .b(gate256inter7), .O(gate256inter9));
  nand2 gate585(.a(s_5), .b(gate256inter3), .O(gate256inter10));
  nor2  gate586(.a(gate256inter10), .b(gate256inter9), .O(gate256inter11));
  nor2  gate587(.a(gate256inter11), .b(gate256inter6), .O(gate256inter12));
  nand2 gate588(.a(gate256inter12), .b(gate256inter1), .O(G769));
nand2 gate257( .a(G754), .b(G755), .O(G770) );

  xor2  gate603(.a(G757), .b(G756), .O(gate258inter0));
  nand2 gate604(.a(gate258inter0), .b(s_8), .O(gate258inter1));
  and2  gate605(.a(G757), .b(G756), .O(gate258inter2));
  inv1  gate606(.a(s_8), .O(gate258inter3));
  inv1  gate607(.a(s_9), .O(gate258inter4));
  nand2 gate608(.a(gate258inter4), .b(gate258inter3), .O(gate258inter5));
  nor2  gate609(.a(gate258inter5), .b(gate258inter2), .O(gate258inter6));
  inv1  gate610(.a(G756), .O(gate258inter7));
  inv1  gate611(.a(G757), .O(gate258inter8));
  nand2 gate612(.a(gate258inter8), .b(gate258inter7), .O(gate258inter9));
  nand2 gate613(.a(s_9), .b(gate258inter3), .O(gate258inter10));
  nor2  gate614(.a(gate258inter10), .b(gate258inter9), .O(gate258inter11));
  nor2  gate615(.a(gate258inter11), .b(gate258inter6), .O(gate258inter12));
  nand2 gate616(.a(gate258inter12), .b(gate258inter1), .O(G773));
nand2 gate259( .a(G758), .b(G759), .O(G776) );
nand2 gate260( .a(G760), .b(G761), .O(G779) );
nand2 gate261( .a(G762), .b(G763), .O(G782) );
nand2 gate262( .a(G764), .b(G765), .O(G785) );
nand2 gate263( .a(G766), .b(G767), .O(G788) );
nand2 gate264( .a(G768), .b(G769), .O(G791) );
nand2 gate265( .a(G642), .b(G770), .O(G794) );
nand2 gate266( .a(G645), .b(G773), .O(G797) );
nand2 gate267( .a(G648), .b(G776), .O(G800) );
nand2 gate268( .a(G651), .b(G779), .O(G803) );
nand2 gate269( .a(G654), .b(G782), .O(G806) );
nand2 gate270( .a(G657), .b(G785), .O(G809) );
nand2 gate271( .a(G660), .b(G788), .O(G812) );
nand2 gate272( .a(G663), .b(G791), .O(G815) );
nand2 gate273( .a(G642), .b(G794), .O(G818) );
nand2 gate274( .a(G770), .b(G794), .O(G819) );

  xor2  gate953(.a(G797), .b(G645), .O(gate275inter0));
  nand2 gate954(.a(gate275inter0), .b(s_58), .O(gate275inter1));
  and2  gate955(.a(G797), .b(G645), .O(gate275inter2));
  inv1  gate956(.a(s_58), .O(gate275inter3));
  inv1  gate957(.a(s_59), .O(gate275inter4));
  nand2 gate958(.a(gate275inter4), .b(gate275inter3), .O(gate275inter5));
  nor2  gate959(.a(gate275inter5), .b(gate275inter2), .O(gate275inter6));
  inv1  gate960(.a(G645), .O(gate275inter7));
  inv1  gate961(.a(G797), .O(gate275inter8));
  nand2 gate962(.a(gate275inter8), .b(gate275inter7), .O(gate275inter9));
  nand2 gate963(.a(s_59), .b(gate275inter3), .O(gate275inter10));
  nor2  gate964(.a(gate275inter10), .b(gate275inter9), .O(gate275inter11));
  nor2  gate965(.a(gate275inter11), .b(gate275inter6), .O(gate275inter12));
  nand2 gate966(.a(gate275inter12), .b(gate275inter1), .O(G820));
nand2 gate276( .a(G773), .b(G797), .O(G821) );
nand2 gate277( .a(G648), .b(G800), .O(G822) );

  xor2  gate939(.a(G800), .b(G776), .O(gate278inter0));
  nand2 gate940(.a(gate278inter0), .b(s_56), .O(gate278inter1));
  and2  gate941(.a(G800), .b(G776), .O(gate278inter2));
  inv1  gate942(.a(s_56), .O(gate278inter3));
  inv1  gate943(.a(s_57), .O(gate278inter4));
  nand2 gate944(.a(gate278inter4), .b(gate278inter3), .O(gate278inter5));
  nor2  gate945(.a(gate278inter5), .b(gate278inter2), .O(gate278inter6));
  inv1  gate946(.a(G776), .O(gate278inter7));
  inv1  gate947(.a(G800), .O(gate278inter8));
  nand2 gate948(.a(gate278inter8), .b(gate278inter7), .O(gate278inter9));
  nand2 gate949(.a(s_57), .b(gate278inter3), .O(gate278inter10));
  nor2  gate950(.a(gate278inter10), .b(gate278inter9), .O(gate278inter11));
  nor2  gate951(.a(gate278inter11), .b(gate278inter6), .O(gate278inter12));
  nand2 gate952(.a(gate278inter12), .b(gate278inter1), .O(G823));
nand2 gate279( .a(G651), .b(G803), .O(G824) );
nand2 gate280( .a(G779), .b(G803), .O(G825) );
nand2 gate281( .a(G654), .b(G806), .O(G826) );
nand2 gate282( .a(G782), .b(G806), .O(G827) );

  xor2  gate995(.a(G809), .b(G657), .O(gate283inter0));
  nand2 gate996(.a(gate283inter0), .b(s_64), .O(gate283inter1));
  and2  gate997(.a(G809), .b(G657), .O(gate283inter2));
  inv1  gate998(.a(s_64), .O(gate283inter3));
  inv1  gate999(.a(s_65), .O(gate283inter4));
  nand2 gate1000(.a(gate283inter4), .b(gate283inter3), .O(gate283inter5));
  nor2  gate1001(.a(gate283inter5), .b(gate283inter2), .O(gate283inter6));
  inv1  gate1002(.a(G657), .O(gate283inter7));
  inv1  gate1003(.a(G809), .O(gate283inter8));
  nand2 gate1004(.a(gate283inter8), .b(gate283inter7), .O(gate283inter9));
  nand2 gate1005(.a(s_65), .b(gate283inter3), .O(gate283inter10));
  nor2  gate1006(.a(gate283inter10), .b(gate283inter9), .O(gate283inter11));
  nor2  gate1007(.a(gate283inter11), .b(gate283inter6), .O(gate283inter12));
  nand2 gate1008(.a(gate283inter12), .b(gate283inter1), .O(G828));

  xor2  gate813(.a(G809), .b(G785), .O(gate284inter0));
  nand2 gate814(.a(gate284inter0), .b(s_38), .O(gate284inter1));
  and2  gate815(.a(G809), .b(G785), .O(gate284inter2));
  inv1  gate816(.a(s_38), .O(gate284inter3));
  inv1  gate817(.a(s_39), .O(gate284inter4));
  nand2 gate818(.a(gate284inter4), .b(gate284inter3), .O(gate284inter5));
  nor2  gate819(.a(gate284inter5), .b(gate284inter2), .O(gate284inter6));
  inv1  gate820(.a(G785), .O(gate284inter7));
  inv1  gate821(.a(G809), .O(gate284inter8));
  nand2 gate822(.a(gate284inter8), .b(gate284inter7), .O(gate284inter9));
  nand2 gate823(.a(s_39), .b(gate284inter3), .O(gate284inter10));
  nor2  gate824(.a(gate284inter10), .b(gate284inter9), .O(gate284inter11));
  nor2  gate825(.a(gate284inter11), .b(gate284inter6), .O(gate284inter12));
  nand2 gate826(.a(gate284inter12), .b(gate284inter1), .O(G829));
nand2 gate285( .a(G660), .b(G812), .O(G830) );
nand2 gate286( .a(G788), .b(G812), .O(G831) );

  xor2  gate1163(.a(G815), .b(G663), .O(gate287inter0));
  nand2 gate1164(.a(gate287inter0), .b(s_88), .O(gate287inter1));
  and2  gate1165(.a(G815), .b(G663), .O(gate287inter2));
  inv1  gate1166(.a(s_88), .O(gate287inter3));
  inv1  gate1167(.a(s_89), .O(gate287inter4));
  nand2 gate1168(.a(gate287inter4), .b(gate287inter3), .O(gate287inter5));
  nor2  gate1169(.a(gate287inter5), .b(gate287inter2), .O(gate287inter6));
  inv1  gate1170(.a(G663), .O(gate287inter7));
  inv1  gate1171(.a(G815), .O(gate287inter8));
  nand2 gate1172(.a(gate287inter8), .b(gate287inter7), .O(gate287inter9));
  nand2 gate1173(.a(s_89), .b(gate287inter3), .O(gate287inter10));
  nor2  gate1174(.a(gate287inter10), .b(gate287inter9), .O(gate287inter11));
  nor2  gate1175(.a(gate287inter11), .b(gate287inter6), .O(gate287inter12));
  nand2 gate1176(.a(gate287inter12), .b(gate287inter1), .O(G832));
nand2 gate288( .a(G791), .b(G815), .O(G833) );
nand2 gate289( .a(G818), .b(G819), .O(G834) );
nand2 gate290( .a(G820), .b(G821), .O(G847) );
nand2 gate291( .a(G822), .b(G823), .O(G860) );
nand2 gate292( .a(G824), .b(G825), .O(G873) );
nand2 gate293( .a(G828), .b(G829), .O(G886) );
nand2 gate294( .a(G832), .b(G833), .O(G899) );
nand2 gate295( .a(G830), .b(G831), .O(G912) );
nand2 gate296( .a(G826), .b(G827), .O(G925) );
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );
nand2 gate387( .a(G1), .b(G1036), .O(G1132) );
nand2 gate388( .a(G2), .b(G1039), .O(G1135) );
nand2 gate389( .a(G3), .b(G1042), .O(G1138) );
nand2 gate390( .a(G4), .b(G1045), .O(G1141) );
nand2 gate391( .a(G5), .b(G1048), .O(G1144) );
nand2 gate392( .a(G6), .b(G1051), .O(G1147) );

  xor2  gate743(.a(G1054), .b(G7), .O(gate393inter0));
  nand2 gate744(.a(gate393inter0), .b(s_28), .O(gate393inter1));
  and2  gate745(.a(G1054), .b(G7), .O(gate393inter2));
  inv1  gate746(.a(s_28), .O(gate393inter3));
  inv1  gate747(.a(s_29), .O(gate393inter4));
  nand2 gate748(.a(gate393inter4), .b(gate393inter3), .O(gate393inter5));
  nor2  gate749(.a(gate393inter5), .b(gate393inter2), .O(gate393inter6));
  inv1  gate750(.a(G7), .O(gate393inter7));
  inv1  gate751(.a(G1054), .O(gate393inter8));
  nand2 gate752(.a(gate393inter8), .b(gate393inter7), .O(gate393inter9));
  nand2 gate753(.a(s_29), .b(gate393inter3), .O(gate393inter10));
  nor2  gate754(.a(gate393inter10), .b(gate393inter9), .O(gate393inter11));
  nor2  gate755(.a(gate393inter11), .b(gate393inter6), .O(gate393inter12));
  nand2 gate756(.a(gate393inter12), .b(gate393inter1), .O(G1150));
nand2 gate394( .a(G8), .b(G1057), .O(G1153) );
nand2 gate395( .a(G9), .b(G1060), .O(G1156) );
nand2 gate396( .a(G10), .b(G1063), .O(G1159) );
nand2 gate397( .a(G11), .b(G1066), .O(G1162) );

  xor2  gate589(.a(G1069), .b(G12), .O(gate398inter0));
  nand2 gate590(.a(gate398inter0), .b(s_6), .O(gate398inter1));
  and2  gate591(.a(G1069), .b(G12), .O(gate398inter2));
  inv1  gate592(.a(s_6), .O(gate398inter3));
  inv1  gate593(.a(s_7), .O(gate398inter4));
  nand2 gate594(.a(gate398inter4), .b(gate398inter3), .O(gate398inter5));
  nor2  gate595(.a(gate398inter5), .b(gate398inter2), .O(gate398inter6));
  inv1  gate596(.a(G12), .O(gate398inter7));
  inv1  gate597(.a(G1069), .O(gate398inter8));
  nand2 gate598(.a(gate398inter8), .b(gate398inter7), .O(gate398inter9));
  nand2 gate599(.a(s_7), .b(gate398inter3), .O(gate398inter10));
  nor2  gate600(.a(gate398inter10), .b(gate398inter9), .O(gate398inter11));
  nor2  gate601(.a(gate398inter11), .b(gate398inter6), .O(gate398inter12));
  nand2 gate602(.a(gate398inter12), .b(gate398inter1), .O(G1165));

  xor2  gate1051(.a(G1072), .b(G13), .O(gate399inter0));
  nand2 gate1052(.a(gate399inter0), .b(s_72), .O(gate399inter1));
  and2  gate1053(.a(G1072), .b(G13), .O(gate399inter2));
  inv1  gate1054(.a(s_72), .O(gate399inter3));
  inv1  gate1055(.a(s_73), .O(gate399inter4));
  nand2 gate1056(.a(gate399inter4), .b(gate399inter3), .O(gate399inter5));
  nor2  gate1057(.a(gate399inter5), .b(gate399inter2), .O(gate399inter6));
  inv1  gate1058(.a(G13), .O(gate399inter7));
  inv1  gate1059(.a(G1072), .O(gate399inter8));
  nand2 gate1060(.a(gate399inter8), .b(gate399inter7), .O(gate399inter9));
  nand2 gate1061(.a(s_73), .b(gate399inter3), .O(gate399inter10));
  nor2  gate1062(.a(gate399inter10), .b(gate399inter9), .O(gate399inter11));
  nor2  gate1063(.a(gate399inter11), .b(gate399inter6), .O(gate399inter12));
  nand2 gate1064(.a(gate399inter12), .b(gate399inter1), .O(G1168));
nand2 gate400( .a(G14), .b(G1075), .O(G1171) );
nand2 gate401( .a(G15), .b(G1078), .O(G1174) );
nand2 gate402( .a(G16), .b(G1081), .O(G1177) );
nand2 gate403( .a(G17), .b(G1084), .O(G1180) );
nand2 gate404( .a(G18), .b(G1087), .O(G1183) );
nand2 gate405( .a(G19), .b(G1090), .O(G1186) );
nand2 gate406( .a(G20), .b(G1093), .O(G1189) );
nand2 gate407( .a(G21), .b(G1096), .O(G1192) );
nand2 gate408( .a(G22), .b(G1099), .O(G1195) );

  xor2  gate1079(.a(G1102), .b(G23), .O(gate409inter0));
  nand2 gate1080(.a(gate409inter0), .b(s_76), .O(gate409inter1));
  and2  gate1081(.a(G1102), .b(G23), .O(gate409inter2));
  inv1  gate1082(.a(s_76), .O(gate409inter3));
  inv1  gate1083(.a(s_77), .O(gate409inter4));
  nand2 gate1084(.a(gate409inter4), .b(gate409inter3), .O(gate409inter5));
  nor2  gate1085(.a(gate409inter5), .b(gate409inter2), .O(gate409inter6));
  inv1  gate1086(.a(G23), .O(gate409inter7));
  inv1  gate1087(.a(G1102), .O(gate409inter8));
  nand2 gate1088(.a(gate409inter8), .b(gate409inter7), .O(gate409inter9));
  nand2 gate1089(.a(s_77), .b(gate409inter3), .O(gate409inter10));
  nor2  gate1090(.a(gate409inter10), .b(gate409inter9), .O(gate409inter11));
  nor2  gate1091(.a(gate409inter11), .b(gate409inter6), .O(gate409inter12));
  nand2 gate1092(.a(gate409inter12), .b(gate409inter1), .O(G1198));
nand2 gate410( .a(G24), .b(G1105), .O(G1201) );
nand2 gate411( .a(G25), .b(G1108), .O(G1204) );

  xor2  gate631(.a(G1111), .b(G26), .O(gate412inter0));
  nand2 gate632(.a(gate412inter0), .b(s_12), .O(gate412inter1));
  and2  gate633(.a(G1111), .b(G26), .O(gate412inter2));
  inv1  gate634(.a(s_12), .O(gate412inter3));
  inv1  gate635(.a(s_13), .O(gate412inter4));
  nand2 gate636(.a(gate412inter4), .b(gate412inter3), .O(gate412inter5));
  nor2  gate637(.a(gate412inter5), .b(gate412inter2), .O(gate412inter6));
  inv1  gate638(.a(G26), .O(gate412inter7));
  inv1  gate639(.a(G1111), .O(gate412inter8));
  nand2 gate640(.a(gate412inter8), .b(gate412inter7), .O(gate412inter9));
  nand2 gate641(.a(s_13), .b(gate412inter3), .O(gate412inter10));
  nor2  gate642(.a(gate412inter10), .b(gate412inter9), .O(gate412inter11));
  nor2  gate643(.a(gate412inter11), .b(gate412inter6), .O(gate412inter12));
  nand2 gate644(.a(gate412inter12), .b(gate412inter1), .O(G1207));
nand2 gate413( .a(G27), .b(G1114), .O(G1210) );

  xor2  gate1205(.a(G1117), .b(G28), .O(gate414inter0));
  nand2 gate1206(.a(gate414inter0), .b(s_94), .O(gate414inter1));
  and2  gate1207(.a(G1117), .b(G28), .O(gate414inter2));
  inv1  gate1208(.a(s_94), .O(gate414inter3));
  inv1  gate1209(.a(s_95), .O(gate414inter4));
  nand2 gate1210(.a(gate414inter4), .b(gate414inter3), .O(gate414inter5));
  nor2  gate1211(.a(gate414inter5), .b(gate414inter2), .O(gate414inter6));
  inv1  gate1212(.a(G28), .O(gate414inter7));
  inv1  gate1213(.a(G1117), .O(gate414inter8));
  nand2 gate1214(.a(gate414inter8), .b(gate414inter7), .O(gate414inter9));
  nand2 gate1215(.a(s_95), .b(gate414inter3), .O(gate414inter10));
  nor2  gate1216(.a(gate414inter10), .b(gate414inter9), .O(gate414inter11));
  nor2  gate1217(.a(gate414inter11), .b(gate414inter6), .O(gate414inter12));
  nand2 gate1218(.a(gate414inter12), .b(gate414inter1), .O(G1213));
nand2 gate415( .a(G29), .b(G1120), .O(G1216) );

  xor2  gate1023(.a(G1123), .b(G30), .O(gate416inter0));
  nand2 gate1024(.a(gate416inter0), .b(s_68), .O(gate416inter1));
  and2  gate1025(.a(G1123), .b(G30), .O(gate416inter2));
  inv1  gate1026(.a(s_68), .O(gate416inter3));
  inv1  gate1027(.a(s_69), .O(gate416inter4));
  nand2 gate1028(.a(gate416inter4), .b(gate416inter3), .O(gate416inter5));
  nor2  gate1029(.a(gate416inter5), .b(gate416inter2), .O(gate416inter6));
  inv1  gate1030(.a(G30), .O(gate416inter7));
  inv1  gate1031(.a(G1123), .O(gate416inter8));
  nand2 gate1032(.a(gate416inter8), .b(gate416inter7), .O(gate416inter9));
  nand2 gate1033(.a(s_69), .b(gate416inter3), .O(gate416inter10));
  nor2  gate1034(.a(gate416inter10), .b(gate416inter9), .O(gate416inter11));
  nor2  gate1035(.a(gate416inter11), .b(gate416inter6), .O(gate416inter12));
  nand2 gate1036(.a(gate416inter12), .b(gate416inter1), .O(G1219));
nand2 gate417( .a(G31), .b(G1126), .O(G1222) );
nand2 gate418( .a(G32), .b(G1129), .O(G1225) );
nand2 gate419( .a(G1), .b(G1132), .O(G1228) );
nand2 gate420( .a(G1036), .b(G1132), .O(G1229) );
nand2 gate421( .a(G2), .b(G1135), .O(G1230) );
nand2 gate422( .a(G1039), .b(G1135), .O(G1231) );
nand2 gate423( .a(G3), .b(G1138), .O(G1232) );
nand2 gate424( .a(G1042), .b(G1138), .O(G1233) );
nand2 gate425( .a(G4), .b(G1141), .O(G1234) );

  xor2  gate1219(.a(G1141), .b(G1045), .O(gate426inter0));
  nand2 gate1220(.a(gate426inter0), .b(s_96), .O(gate426inter1));
  and2  gate1221(.a(G1141), .b(G1045), .O(gate426inter2));
  inv1  gate1222(.a(s_96), .O(gate426inter3));
  inv1  gate1223(.a(s_97), .O(gate426inter4));
  nand2 gate1224(.a(gate426inter4), .b(gate426inter3), .O(gate426inter5));
  nor2  gate1225(.a(gate426inter5), .b(gate426inter2), .O(gate426inter6));
  inv1  gate1226(.a(G1045), .O(gate426inter7));
  inv1  gate1227(.a(G1141), .O(gate426inter8));
  nand2 gate1228(.a(gate426inter8), .b(gate426inter7), .O(gate426inter9));
  nand2 gate1229(.a(s_97), .b(gate426inter3), .O(gate426inter10));
  nor2  gate1230(.a(gate426inter10), .b(gate426inter9), .O(gate426inter11));
  nor2  gate1231(.a(gate426inter11), .b(gate426inter6), .O(gate426inter12));
  nand2 gate1232(.a(gate426inter12), .b(gate426inter1), .O(G1235));
nand2 gate427( .a(G5), .b(G1144), .O(G1236) );
nand2 gate428( .a(G1048), .b(G1144), .O(G1237) );
nand2 gate429( .a(G6), .b(G1147), .O(G1238) );
nand2 gate430( .a(G1051), .b(G1147), .O(G1239) );
nand2 gate431( .a(G7), .b(G1150), .O(G1240) );
nand2 gate432( .a(G1054), .b(G1150), .O(G1241) );
nand2 gate433( .a(G8), .b(G1153), .O(G1242) );
nand2 gate434( .a(G1057), .b(G1153), .O(G1243) );
nand2 gate435( .a(G9), .b(G1156), .O(G1244) );
nand2 gate436( .a(G1060), .b(G1156), .O(G1245) );
nand2 gate437( .a(G10), .b(G1159), .O(G1246) );
nand2 gate438( .a(G1063), .b(G1159), .O(G1247) );
nand2 gate439( .a(G11), .b(G1162), .O(G1248) );
nand2 gate440( .a(G1066), .b(G1162), .O(G1249) );

  xor2  gate869(.a(G1165), .b(G12), .O(gate441inter0));
  nand2 gate870(.a(gate441inter0), .b(s_46), .O(gate441inter1));
  and2  gate871(.a(G1165), .b(G12), .O(gate441inter2));
  inv1  gate872(.a(s_46), .O(gate441inter3));
  inv1  gate873(.a(s_47), .O(gate441inter4));
  nand2 gate874(.a(gate441inter4), .b(gate441inter3), .O(gate441inter5));
  nor2  gate875(.a(gate441inter5), .b(gate441inter2), .O(gate441inter6));
  inv1  gate876(.a(G12), .O(gate441inter7));
  inv1  gate877(.a(G1165), .O(gate441inter8));
  nand2 gate878(.a(gate441inter8), .b(gate441inter7), .O(gate441inter9));
  nand2 gate879(.a(s_47), .b(gate441inter3), .O(gate441inter10));
  nor2  gate880(.a(gate441inter10), .b(gate441inter9), .O(gate441inter11));
  nor2  gate881(.a(gate441inter11), .b(gate441inter6), .O(gate441inter12));
  nand2 gate882(.a(gate441inter12), .b(gate441inter1), .O(G1250));
nand2 gate442( .a(G1069), .b(G1165), .O(G1251) );

  xor2  gate1317(.a(G1168), .b(G13), .O(gate443inter0));
  nand2 gate1318(.a(gate443inter0), .b(s_110), .O(gate443inter1));
  and2  gate1319(.a(G1168), .b(G13), .O(gate443inter2));
  inv1  gate1320(.a(s_110), .O(gate443inter3));
  inv1  gate1321(.a(s_111), .O(gate443inter4));
  nand2 gate1322(.a(gate443inter4), .b(gate443inter3), .O(gate443inter5));
  nor2  gate1323(.a(gate443inter5), .b(gate443inter2), .O(gate443inter6));
  inv1  gate1324(.a(G13), .O(gate443inter7));
  inv1  gate1325(.a(G1168), .O(gate443inter8));
  nand2 gate1326(.a(gate443inter8), .b(gate443inter7), .O(gate443inter9));
  nand2 gate1327(.a(s_111), .b(gate443inter3), .O(gate443inter10));
  nor2  gate1328(.a(gate443inter10), .b(gate443inter9), .O(gate443inter11));
  nor2  gate1329(.a(gate443inter11), .b(gate443inter6), .O(gate443inter12));
  nand2 gate1330(.a(gate443inter12), .b(gate443inter1), .O(G1252));
nand2 gate444( .a(G1072), .b(G1168), .O(G1253) );
nand2 gate445( .a(G14), .b(G1171), .O(G1254) );
nand2 gate446( .a(G1075), .b(G1171), .O(G1255) );
nand2 gate447( .a(G15), .b(G1174), .O(G1256) );
nand2 gate448( .a(G1078), .b(G1174), .O(G1257) );
nand2 gate449( .a(G16), .b(G1177), .O(G1258) );
nand2 gate450( .a(G1081), .b(G1177), .O(G1259) );
nand2 gate451( .a(G17), .b(G1180), .O(G1260) );
nand2 gate452( .a(G1084), .b(G1180), .O(G1261) );
nand2 gate453( .a(G18), .b(G1183), .O(G1262) );
nand2 gate454( .a(G1087), .b(G1183), .O(G1263) );
nand2 gate455( .a(G19), .b(G1186), .O(G1264) );
nand2 gate456( .a(G1090), .b(G1186), .O(G1265) );

  xor2  gate1093(.a(G1189), .b(G20), .O(gate457inter0));
  nand2 gate1094(.a(gate457inter0), .b(s_78), .O(gate457inter1));
  and2  gate1095(.a(G1189), .b(G20), .O(gate457inter2));
  inv1  gate1096(.a(s_78), .O(gate457inter3));
  inv1  gate1097(.a(s_79), .O(gate457inter4));
  nand2 gate1098(.a(gate457inter4), .b(gate457inter3), .O(gate457inter5));
  nor2  gate1099(.a(gate457inter5), .b(gate457inter2), .O(gate457inter6));
  inv1  gate1100(.a(G20), .O(gate457inter7));
  inv1  gate1101(.a(G1189), .O(gate457inter8));
  nand2 gate1102(.a(gate457inter8), .b(gate457inter7), .O(gate457inter9));
  nand2 gate1103(.a(s_79), .b(gate457inter3), .O(gate457inter10));
  nor2  gate1104(.a(gate457inter10), .b(gate457inter9), .O(gate457inter11));
  nor2  gate1105(.a(gate457inter11), .b(gate457inter6), .O(gate457inter12));
  nand2 gate1106(.a(gate457inter12), .b(gate457inter1), .O(G1266));
nand2 gate458( .a(G1093), .b(G1189), .O(G1267) );
nand2 gate459( .a(G21), .b(G1192), .O(G1268) );
nand2 gate460( .a(G1096), .b(G1192), .O(G1269) );
nand2 gate461( .a(G22), .b(G1195), .O(G1270) );
nand2 gate462( .a(G1099), .b(G1195), .O(G1271) );
nand2 gate463( .a(G23), .b(G1198), .O(G1272) );
nand2 gate464( .a(G1102), .b(G1198), .O(G1273) );
nand2 gate465( .a(G24), .b(G1201), .O(G1274) );
nand2 gate466( .a(G1105), .b(G1201), .O(G1275) );
nand2 gate467( .a(G25), .b(G1204), .O(G1276) );

  xor2  gate561(.a(G1204), .b(G1108), .O(gate468inter0));
  nand2 gate562(.a(gate468inter0), .b(s_2), .O(gate468inter1));
  and2  gate563(.a(G1204), .b(G1108), .O(gate468inter2));
  inv1  gate564(.a(s_2), .O(gate468inter3));
  inv1  gate565(.a(s_3), .O(gate468inter4));
  nand2 gate566(.a(gate468inter4), .b(gate468inter3), .O(gate468inter5));
  nor2  gate567(.a(gate468inter5), .b(gate468inter2), .O(gate468inter6));
  inv1  gate568(.a(G1108), .O(gate468inter7));
  inv1  gate569(.a(G1204), .O(gate468inter8));
  nand2 gate570(.a(gate468inter8), .b(gate468inter7), .O(gate468inter9));
  nand2 gate571(.a(s_3), .b(gate468inter3), .O(gate468inter10));
  nor2  gate572(.a(gate468inter10), .b(gate468inter9), .O(gate468inter11));
  nor2  gate573(.a(gate468inter11), .b(gate468inter6), .O(gate468inter12));
  nand2 gate574(.a(gate468inter12), .b(gate468inter1), .O(G1277));
nand2 gate469( .a(G26), .b(G1207), .O(G1278) );
nand2 gate470( .a(G1111), .b(G1207), .O(G1279) );

  xor2  gate715(.a(G1210), .b(G27), .O(gate471inter0));
  nand2 gate716(.a(gate471inter0), .b(s_24), .O(gate471inter1));
  and2  gate717(.a(G1210), .b(G27), .O(gate471inter2));
  inv1  gate718(.a(s_24), .O(gate471inter3));
  inv1  gate719(.a(s_25), .O(gate471inter4));
  nand2 gate720(.a(gate471inter4), .b(gate471inter3), .O(gate471inter5));
  nor2  gate721(.a(gate471inter5), .b(gate471inter2), .O(gate471inter6));
  inv1  gate722(.a(G27), .O(gate471inter7));
  inv1  gate723(.a(G1210), .O(gate471inter8));
  nand2 gate724(.a(gate471inter8), .b(gate471inter7), .O(gate471inter9));
  nand2 gate725(.a(s_25), .b(gate471inter3), .O(gate471inter10));
  nor2  gate726(.a(gate471inter10), .b(gate471inter9), .O(gate471inter11));
  nor2  gate727(.a(gate471inter11), .b(gate471inter6), .O(gate471inter12));
  nand2 gate728(.a(gate471inter12), .b(gate471inter1), .O(G1280));
nand2 gate472( .a(G1114), .b(G1210), .O(G1281) );
nand2 gate473( .a(G28), .b(G1213), .O(G1282) );
nand2 gate474( .a(G1117), .b(G1213), .O(G1283) );
nand2 gate475( .a(G29), .b(G1216), .O(G1284) );
nand2 gate476( .a(G1120), .b(G1216), .O(G1285) );
nand2 gate477( .a(G30), .b(G1219), .O(G1286) );
nand2 gate478( .a(G1123), .b(G1219), .O(G1287) );
nand2 gate479( .a(G31), .b(G1222), .O(G1288) );
nand2 gate480( .a(G1126), .b(G1222), .O(G1289) );

  xor2  gate785(.a(G1225), .b(G32), .O(gate481inter0));
  nand2 gate786(.a(gate481inter0), .b(s_34), .O(gate481inter1));
  and2  gate787(.a(G1225), .b(G32), .O(gate481inter2));
  inv1  gate788(.a(s_34), .O(gate481inter3));
  inv1  gate789(.a(s_35), .O(gate481inter4));
  nand2 gate790(.a(gate481inter4), .b(gate481inter3), .O(gate481inter5));
  nor2  gate791(.a(gate481inter5), .b(gate481inter2), .O(gate481inter6));
  inv1  gate792(.a(G32), .O(gate481inter7));
  inv1  gate793(.a(G1225), .O(gate481inter8));
  nand2 gate794(.a(gate481inter8), .b(gate481inter7), .O(gate481inter9));
  nand2 gate795(.a(s_35), .b(gate481inter3), .O(gate481inter10));
  nor2  gate796(.a(gate481inter10), .b(gate481inter9), .O(gate481inter11));
  nor2  gate797(.a(gate481inter11), .b(gate481inter6), .O(gate481inter12));
  nand2 gate798(.a(gate481inter12), .b(gate481inter1), .O(G1290));

  xor2  gate1373(.a(G1225), .b(G1129), .O(gate482inter0));
  nand2 gate1374(.a(gate482inter0), .b(s_118), .O(gate482inter1));
  and2  gate1375(.a(G1225), .b(G1129), .O(gate482inter2));
  inv1  gate1376(.a(s_118), .O(gate482inter3));
  inv1  gate1377(.a(s_119), .O(gate482inter4));
  nand2 gate1378(.a(gate482inter4), .b(gate482inter3), .O(gate482inter5));
  nor2  gate1379(.a(gate482inter5), .b(gate482inter2), .O(gate482inter6));
  inv1  gate1380(.a(G1129), .O(gate482inter7));
  inv1  gate1381(.a(G1225), .O(gate482inter8));
  nand2 gate1382(.a(gate482inter8), .b(gate482inter7), .O(gate482inter9));
  nand2 gate1383(.a(s_119), .b(gate482inter3), .O(gate482inter10));
  nor2  gate1384(.a(gate482inter10), .b(gate482inter9), .O(gate482inter11));
  nor2  gate1385(.a(gate482inter11), .b(gate482inter6), .O(gate482inter12));
  nand2 gate1386(.a(gate482inter12), .b(gate482inter1), .O(G1291));

  xor2  gate1275(.a(G1229), .b(G1228), .O(gate483inter0));
  nand2 gate1276(.a(gate483inter0), .b(s_104), .O(gate483inter1));
  and2  gate1277(.a(G1229), .b(G1228), .O(gate483inter2));
  inv1  gate1278(.a(s_104), .O(gate483inter3));
  inv1  gate1279(.a(s_105), .O(gate483inter4));
  nand2 gate1280(.a(gate483inter4), .b(gate483inter3), .O(gate483inter5));
  nor2  gate1281(.a(gate483inter5), .b(gate483inter2), .O(gate483inter6));
  inv1  gate1282(.a(G1228), .O(gate483inter7));
  inv1  gate1283(.a(G1229), .O(gate483inter8));
  nand2 gate1284(.a(gate483inter8), .b(gate483inter7), .O(gate483inter9));
  nand2 gate1285(.a(s_105), .b(gate483inter3), .O(gate483inter10));
  nor2  gate1286(.a(gate483inter10), .b(gate483inter9), .O(gate483inter11));
  nor2  gate1287(.a(gate483inter11), .b(gate483inter6), .O(gate483inter12));
  nand2 gate1288(.a(gate483inter12), .b(gate483inter1), .O(G1292));
nand2 gate484( .a(G1230), .b(G1231), .O(G1293) );
nand2 gate485( .a(G1232), .b(G1233), .O(G1294) );
nand2 gate486( .a(G1234), .b(G1235), .O(G1295) );
nand2 gate487( .a(G1236), .b(G1237), .O(G1296) );
nand2 gate488( .a(G1238), .b(G1239), .O(G1297) );
nand2 gate489( .a(G1240), .b(G1241), .O(G1298) );
nand2 gate490( .a(G1242), .b(G1243), .O(G1299) );
nand2 gate491( .a(G1244), .b(G1245), .O(G1300) );
nand2 gate492( .a(G1246), .b(G1247), .O(G1301) );
nand2 gate493( .a(G1248), .b(G1249), .O(G1302) );
nand2 gate494( .a(G1250), .b(G1251), .O(G1303) );
nand2 gate495( .a(G1252), .b(G1253), .O(G1304) );
nand2 gate496( .a(G1254), .b(G1255), .O(G1305) );
nand2 gate497( .a(G1256), .b(G1257), .O(G1306) );
nand2 gate498( .a(G1258), .b(G1259), .O(G1307) );
nand2 gate499( .a(G1260), .b(G1261), .O(G1308) );
nand2 gate500( .a(G1262), .b(G1263), .O(G1309) );
nand2 gate501( .a(G1264), .b(G1265), .O(G1310) );
nand2 gate502( .a(G1266), .b(G1267), .O(G1311) );
nand2 gate503( .a(G1268), .b(G1269), .O(G1312) );

  xor2  gate799(.a(G1271), .b(G1270), .O(gate504inter0));
  nand2 gate800(.a(gate504inter0), .b(s_36), .O(gate504inter1));
  and2  gate801(.a(G1271), .b(G1270), .O(gate504inter2));
  inv1  gate802(.a(s_36), .O(gate504inter3));
  inv1  gate803(.a(s_37), .O(gate504inter4));
  nand2 gate804(.a(gate504inter4), .b(gate504inter3), .O(gate504inter5));
  nor2  gate805(.a(gate504inter5), .b(gate504inter2), .O(gate504inter6));
  inv1  gate806(.a(G1270), .O(gate504inter7));
  inv1  gate807(.a(G1271), .O(gate504inter8));
  nand2 gate808(.a(gate504inter8), .b(gate504inter7), .O(gate504inter9));
  nand2 gate809(.a(s_37), .b(gate504inter3), .O(gate504inter10));
  nor2  gate810(.a(gate504inter10), .b(gate504inter9), .O(gate504inter11));
  nor2  gate811(.a(gate504inter11), .b(gate504inter6), .O(gate504inter12));
  nand2 gate812(.a(gate504inter12), .b(gate504inter1), .O(G1313));
nand2 gate505( .a(G1272), .b(G1273), .O(G1314) );
nand2 gate506( .a(G1274), .b(G1275), .O(G1315) );
nand2 gate507( .a(G1276), .b(G1277), .O(G1316) );
nand2 gate508( .a(G1278), .b(G1279), .O(G1317) );
nand2 gate509( .a(G1280), .b(G1281), .O(G1318) );
nand2 gate510( .a(G1282), .b(G1283), .O(G1319) );
nand2 gate511( .a(G1284), .b(G1285), .O(G1320) );

  xor2  gate855(.a(G1287), .b(G1286), .O(gate512inter0));
  nand2 gate856(.a(gate512inter0), .b(s_44), .O(gate512inter1));
  and2  gate857(.a(G1287), .b(G1286), .O(gate512inter2));
  inv1  gate858(.a(s_44), .O(gate512inter3));
  inv1  gate859(.a(s_45), .O(gate512inter4));
  nand2 gate860(.a(gate512inter4), .b(gate512inter3), .O(gate512inter5));
  nor2  gate861(.a(gate512inter5), .b(gate512inter2), .O(gate512inter6));
  inv1  gate862(.a(G1286), .O(gate512inter7));
  inv1  gate863(.a(G1287), .O(gate512inter8));
  nand2 gate864(.a(gate512inter8), .b(gate512inter7), .O(gate512inter9));
  nand2 gate865(.a(s_45), .b(gate512inter3), .O(gate512inter10));
  nor2  gate866(.a(gate512inter10), .b(gate512inter9), .O(gate512inter11));
  nor2  gate867(.a(gate512inter11), .b(gate512inter6), .O(gate512inter12));
  nand2 gate868(.a(gate512inter12), .b(gate512inter1), .O(G1321));
nand2 gate513( .a(G1288), .b(G1289), .O(G1322) );
nand2 gate514( .a(G1290), .b(G1291), .O(G1323) );
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule