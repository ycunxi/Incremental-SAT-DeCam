module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);

input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;//RE__PI;

input s_0,s_1;//RE__ALLOW(00,01,10,11);
input s_2,s_3;//RE__ALLOW(00,01,10,11);
input s_4,s_5;//RE__ALLOW(00,01,10,11);
input s_6,s_7;//RE__ALLOW(00,01,10,11);
input s_8,s_9;//RE__ALLOW(00,01,10,11);
input s_10,s_11;//RE__ALLOW(00,01,10,11);
input s_12,s_13;//RE__ALLOW(00,01,10,11);
input s_14,s_15;//RE__ALLOW(00,01,10,11);
input s_16,s_17;//RE__ALLOW(00,01,10,11);
input s_18,s_19;//RE__ALLOW(00,01,10,11);
input s_20,s_21;//RE__ALLOW(00,01,10,11);
input s_22,s_23;//RE__ALLOW(00,01,10,11);
input s_24,s_25;//RE__ALLOW(00,01,10,11);
input s_26,s_27;//RE__ALLOW(00,01,10,11);
input s_28,s_29;//RE__ALLOW(00,01,10,11);
input s_30,s_31;//RE__ALLOW(00,01,10,11);
input s_32,s_33;//RE__ALLOW(00,01,10,11);
input s_34,s_35;//RE__ALLOW(00,01,10,11);
input s_36,s_37;//RE__ALLOW(00,01,10,11);
input s_38,s_39;//RE__ALLOW(00,01,10,11);
input s_40,s_41;//RE__ALLOW(00,01,10,11);
input s_42,s_43;//RE__ALLOW(00,01,10,11);
input s_44,s_45;//RE__ALLOW(00,01,10,11);
input s_46,s_47;//RE__ALLOW(00,01,10,11);
input s_48,s_49;//RE__ALLOW(00,01,10,11);
input s_50,s_51;//RE__ALLOW(00,01,10,11);
input s_52,s_53;//RE__ALLOW(00,01,10,11);
input s_54,s_55;//RE__ALLOW(00,01,10,11);
input s_56,s_57;//RE__ALLOW(00,01,10,11);
input s_58,s_59;//RE__ALLOW(00,01,10,11);
input s_60,s_61;//RE__ALLOW(00,01,10,11);
input s_62,s_63;//RE__ALLOW(00,01,10,11);
input s_64,s_65;//RE__ALLOW(00,01,10,11);
input s_66,s_67;//RE__ALLOW(00,01,10,11);
input s_68,s_69;//RE__ALLOW(00,01,10,11);
input s_70,s_71;//RE__ALLOW(00,01,10,11);
input s_72,s_73;//RE__ALLOW(00,01,10,11);
input s_74,s_75;//RE__ALLOW(00,01,10,11);
input s_76,s_77;//RE__ALLOW(00,01,10,11);
input s_78,s_79;//RE__ALLOW(00,01,10,11);
input s_80,s_81;//RE__ALLOW(00,01,10,11);
input s_82,s_83;//RE__ALLOW(00,01,10,11);
input s_84,s_85;//RE__ALLOW(00,01,10,11);
input s_86,s_87;//RE__ALLOW(00,01,10,11);
input s_88,s_89;//RE__ALLOW(00,01,10,11);
input s_90,s_91;//RE__ALLOW(00,01,10,11);
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;

  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate221inter0, gate221inter1, gate221inter2, gate221inter3, gate221inter4, gate221inter5, gate221inter6, gate221inter7, gate221inter8, gate221inter9, gate221inter10, gate221inter11, gate221inter12, gate137inter0, gate137inter1, gate137inter2, gate137inter3, gate137inter4, gate137inter5, gate137inter6, gate137inter7, gate137inter8, gate137inter9, gate137inter10, gate137inter11, gate137inter12, gate68inter0, gate68inter1, gate68inter2, gate68inter3, gate68inter4, gate68inter5, gate68inter6, gate68inter7, gate68inter8, gate68inter9, gate68inter10, gate68inter11, gate68inter12, gate135inter0, gate135inter1, gate135inter2, gate135inter3, gate135inter4, gate135inter5, gate135inter6, gate135inter7, gate135inter8, gate135inter9, gate135inter10, gate135inter11, gate135inter12, gate21inter0, gate21inter1, gate21inter2, gate21inter3, gate21inter4, gate21inter5, gate21inter6, gate21inter7, gate21inter8, gate21inter9, gate21inter10, gate21inter11, gate21inter12, gate15inter0, gate15inter1, gate15inter2, gate15inter3, gate15inter4, gate15inter5, gate15inter6, gate15inter7, gate15inter8, gate15inter9, gate15inter10, gate15inter11, gate15inter12, gate231inter0, gate231inter1, gate231inter2, gate231inter3, gate231inter4, gate231inter5, gate231inter6, gate231inter7, gate231inter8, gate231inter9, gate231inter10, gate231inter11, gate231inter12, gate200inter0, gate200inter1, gate200inter2, gate200inter3, gate200inter4, gate200inter5, gate200inter6, gate200inter7, gate200inter8, gate200inter9, gate200inter10, gate200inter11, gate200inter12, gate485inter0, gate485inter1, gate485inter2, gate485inter3, gate485inter4, gate485inter5, gate485inter6, gate485inter7, gate485inter8, gate485inter9, gate485inter10, gate485inter11, gate485inter12, gate134inter0, gate134inter1, gate134inter2, gate134inter3, gate134inter4, gate134inter5, gate134inter6, gate134inter7, gate134inter8, gate134inter9, gate134inter10, gate134inter11, gate134inter12, gate400inter0, gate400inter1, gate400inter2, gate400inter3, gate400inter4, gate400inter5, gate400inter6, gate400inter7, gate400inter8, gate400inter9, gate400inter10, gate400inter11, gate400inter12, gate250inter0, gate250inter1, gate250inter2, gate250inter3, gate250inter4, gate250inter5, gate250inter6, gate250inter7, gate250inter8, gate250inter9, gate250inter10, gate250inter11, gate250inter12, gate161inter0, gate161inter1, gate161inter2, gate161inter3, gate161inter4, gate161inter5, gate161inter6, gate161inter7, gate161inter8, gate161inter9, gate161inter10, gate161inter11, gate161inter12, gate471inter0, gate471inter1, gate471inter2, gate471inter3, gate471inter4, gate471inter5, gate471inter6, gate471inter7, gate471inter8, gate471inter9, gate471inter10, gate471inter11, gate471inter12, gate486inter0, gate486inter1, gate486inter2, gate486inter3, gate486inter4, gate486inter5, gate486inter6, gate486inter7, gate486inter8, gate486inter9, gate486inter10, gate486inter11, gate486inter12, gate194inter0, gate194inter1, gate194inter2, gate194inter3, gate194inter4, gate194inter5, gate194inter6, gate194inter7, gate194inter8, gate194inter9, gate194inter10, gate194inter11, gate194inter12, gate443inter0, gate443inter1, gate443inter2, gate443inter3, gate443inter4, gate443inter5, gate443inter6, gate443inter7, gate443inter8, gate443inter9, gate443inter10, gate443inter11, gate443inter12, gate503inter0, gate503inter1, gate503inter2, gate503inter3, gate503inter4, gate503inter5, gate503inter6, gate503inter7, gate503inter8, gate503inter9, gate503inter10, gate503inter11, gate503inter12, gate463inter0, gate463inter1, gate463inter2, gate463inter3, gate463inter4, gate463inter5, gate463inter6, gate463inter7, gate463inter8, gate463inter9, gate463inter10, gate463inter11, gate463inter12, gate234inter0, gate234inter1, gate234inter2, gate234inter3, gate234inter4, gate234inter5, gate234inter6, gate234inter7, gate234inter8, gate234inter9, gate234inter10, gate234inter11, gate234inter12, gate225inter0, gate225inter1, gate225inter2, gate225inter3, gate225inter4, gate225inter5, gate225inter6, gate225inter7, gate225inter8, gate225inter9, gate225inter10, gate225inter11, gate225inter12, gate91inter0, gate91inter1, gate91inter2, gate91inter3, gate91inter4, gate91inter5, gate91inter6, gate91inter7, gate91inter8, gate91inter9, gate91inter10, gate91inter11, gate91inter12, gate494inter0, gate494inter1, gate494inter2, gate494inter3, gate494inter4, gate494inter5, gate494inter6, gate494inter7, gate494inter8, gate494inter9, gate494inter10, gate494inter11, gate494inter12, gate207inter0, gate207inter1, gate207inter2, gate207inter3, gate207inter4, gate207inter5, gate207inter6, gate207inter7, gate207inter8, gate207inter9, gate207inter10, gate207inter11, gate207inter12, gate398inter0, gate398inter1, gate398inter2, gate398inter3, gate398inter4, gate398inter5, gate398inter6, gate398inter7, gate398inter8, gate398inter9, gate398inter10, gate398inter11, gate398inter12, gate255inter0, gate255inter1, gate255inter2, gate255inter3, gate255inter4, gate255inter5, gate255inter6, gate255inter7, gate255inter8, gate255inter9, gate255inter10, gate255inter11, gate255inter12, gate37inter0, gate37inter1, gate37inter2, gate37inter3, gate37inter4, gate37inter5, gate37inter6, gate37inter7, gate37inter8, gate37inter9, gate37inter10, gate37inter11, gate37inter12, gate417inter0, gate417inter1, gate417inter2, gate417inter3, gate417inter4, gate417inter5, gate417inter6, gate417inter7, gate417inter8, gate417inter9, gate417inter10, gate417inter11, gate417inter12, gate25inter0, gate25inter1, gate25inter2, gate25inter3, gate25inter4, gate25inter5, gate25inter6, gate25inter7, gate25inter8, gate25inter9, gate25inter10, gate25inter11, gate25inter12, gate423inter0, gate423inter1, gate423inter2, gate423inter3, gate423inter4, gate423inter5, gate423inter6, gate423inter7, gate423inter8, gate423inter9, gate423inter10, gate423inter11, gate423inter12, gate45inter0, gate45inter1, gate45inter2, gate45inter3, gate45inter4, gate45inter5, gate45inter6, gate45inter7, gate45inter8, gate45inter9, gate45inter10, gate45inter11, gate45inter12, gate86inter0, gate86inter1, gate86inter2, gate86inter3, gate86inter4, gate86inter5, gate86inter6, gate86inter7, gate86inter8, gate86inter9, gate86inter10, gate86inter11, gate86inter12, gate394inter0, gate394inter1, gate394inter2, gate394inter3, gate394inter4, gate394inter5, gate394inter6, gate394inter7, gate394inter8, gate394inter9, gate394inter10, gate394inter11, gate394inter12, gate23inter0, gate23inter1, gate23inter2, gate23inter3, gate23inter4, gate23inter5, gate23inter6, gate23inter7, gate23inter8, gate23inter9, gate23inter10, gate23inter11, gate23inter12, gate257inter0, gate257inter1, gate257inter2, gate257inter3, gate257inter4, gate257inter5, gate257inter6, gate257inter7, gate257inter8, gate257inter9, gate257inter10, gate257inter11, gate257inter12, gate273inter0, gate273inter1, gate273inter2, gate273inter3, gate273inter4, gate273inter5, gate273inter6, gate273inter7, gate273inter8, gate273inter9, gate273inter10, gate273inter11, gate273inter12, gate145inter0, gate145inter1, gate145inter2, gate145inter3, gate145inter4, gate145inter5, gate145inter6, gate145inter7, gate145inter8, gate145inter9, gate145inter10, gate145inter11, gate145inter12, gate89inter0, gate89inter1, gate89inter2, gate89inter3, gate89inter4, gate89inter5, gate89inter6, gate89inter7, gate89inter8, gate89inter9, gate89inter10, gate89inter11, gate89inter12, gate510inter0, gate510inter1, gate510inter2, gate510inter3, gate510inter4, gate510inter5, gate510inter6, gate510inter7, gate510inter8, gate510inter9, gate510inter10, gate510inter11, gate510inter12, gate191inter0, gate191inter1, gate191inter2, gate191inter3, gate191inter4, gate191inter5, gate191inter6, gate191inter7, gate191inter8, gate191inter9, gate191inter10, gate191inter11, gate191inter12, gate95inter0, gate95inter1, gate95inter2, gate95inter3, gate95inter4, gate95inter5, gate95inter6, gate95inter7, gate95inter8, gate95inter9, gate95inter10, gate95inter11, gate95inter12, gate12inter0, gate12inter1, gate12inter2, gate12inter3, gate12inter4, gate12inter5, gate12inter6, gate12inter7, gate12inter8, gate12inter9, gate12inter10, gate12inter11, gate12inter12, gate422inter0, gate422inter1, gate422inter2, gate422inter3, gate422inter4, gate422inter5, gate422inter6, gate422inter7, gate422inter8, gate422inter9, gate422inter10, gate422inter11, gate422inter12, gate93inter0, gate93inter1, gate93inter2, gate93inter3, gate93inter4, gate93inter5, gate93inter6, gate93inter7, gate93inter8, gate93inter9, gate93inter10, gate93inter11, gate93inter12, gate124inter0, gate124inter1, gate124inter2, gate124inter3, gate124inter4, gate124inter5, gate124inter6, gate124inter7, gate124inter8, gate124inter9, gate124inter10, gate124inter11, gate124inter12, gate261inter0, gate261inter1, gate261inter2, gate261inter3, gate261inter4, gate261inter5, gate261inter6, gate261inter7, gate261inter8, gate261inter9, gate261inter10, gate261inter11, gate261inter12;



and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );
nand2 gate9( .a(G1), .b(G2), .O(G266) );
nand2 gate10( .a(G3), .b(G4), .O(G269) );
nand2 gate11( .a(G5), .b(G6), .O(G272) );

  xor2  gate1121(.a(G8), .b(G7), .O(gate12inter0));
  nand2 gate1122(.a(gate12inter0), .b(s_82), .O(gate12inter1));
  and2  gate1123(.a(G8), .b(G7), .O(gate12inter2));
  inv1  gate1124(.a(s_82), .O(gate12inter3));
  inv1  gate1125(.a(s_83), .O(gate12inter4));
  nand2 gate1126(.a(gate12inter4), .b(gate12inter3), .O(gate12inter5));
  nor2  gate1127(.a(gate12inter5), .b(gate12inter2), .O(gate12inter6));
  inv1  gate1128(.a(G7), .O(gate12inter7));
  inv1  gate1129(.a(G8), .O(gate12inter8));
  nand2 gate1130(.a(gate12inter8), .b(gate12inter7), .O(gate12inter9));
  nand2 gate1131(.a(s_83), .b(gate12inter3), .O(gate12inter10));
  nor2  gate1132(.a(gate12inter10), .b(gate12inter9), .O(gate12inter11));
  nor2  gate1133(.a(gate12inter11), .b(gate12inter6), .O(gate12inter12));
  nand2 gate1134(.a(gate12inter12), .b(gate12inter1), .O(G275));
nand2 gate13( .a(G9), .b(G10), .O(G278) );
nand2 gate14( .a(G11), .b(G12), .O(G281) );

  xor2  gate617(.a(G14), .b(G13), .O(gate15inter0));
  nand2 gate618(.a(gate15inter0), .b(s_10), .O(gate15inter1));
  and2  gate619(.a(G14), .b(G13), .O(gate15inter2));
  inv1  gate620(.a(s_10), .O(gate15inter3));
  inv1  gate621(.a(s_11), .O(gate15inter4));
  nand2 gate622(.a(gate15inter4), .b(gate15inter3), .O(gate15inter5));
  nor2  gate623(.a(gate15inter5), .b(gate15inter2), .O(gate15inter6));
  inv1  gate624(.a(G13), .O(gate15inter7));
  inv1  gate625(.a(G14), .O(gate15inter8));
  nand2 gate626(.a(gate15inter8), .b(gate15inter7), .O(gate15inter9));
  nand2 gate627(.a(s_11), .b(gate15inter3), .O(gate15inter10));
  nor2  gate628(.a(gate15inter10), .b(gate15inter9), .O(gate15inter11));
  nor2  gate629(.a(gate15inter11), .b(gate15inter6), .O(gate15inter12));
  nand2 gate630(.a(gate15inter12), .b(gate15inter1), .O(G284));
nand2 gate16( .a(G15), .b(G16), .O(G287) );
nand2 gate17( .a(G17), .b(G18), .O(G290) );
nand2 gate18( .a(G19), .b(G20), .O(G293) );
nand2 gate19( .a(G21), .b(G22), .O(G296) );
nand2 gate20( .a(G23), .b(G24), .O(G299) );

  xor2  gate603(.a(G26), .b(G25), .O(gate21inter0));
  nand2 gate604(.a(gate21inter0), .b(s_8), .O(gate21inter1));
  and2  gate605(.a(G26), .b(G25), .O(gate21inter2));
  inv1  gate606(.a(s_8), .O(gate21inter3));
  inv1  gate607(.a(s_9), .O(gate21inter4));
  nand2 gate608(.a(gate21inter4), .b(gate21inter3), .O(gate21inter5));
  nor2  gate609(.a(gate21inter5), .b(gate21inter2), .O(gate21inter6));
  inv1  gate610(.a(G25), .O(gate21inter7));
  inv1  gate611(.a(G26), .O(gate21inter8));
  nand2 gate612(.a(gate21inter8), .b(gate21inter7), .O(gate21inter9));
  nand2 gate613(.a(s_9), .b(gate21inter3), .O(gate21inter10));
  nor2  gate614(.a(gate21inter10), .b(gate21inter9), .O(gate21inter11));
  nor2  gate615(.a(gate21inter11), .b(gate21inter6), .O(gate21inter12));
  nand2 gate616(.a(gate21inter12), .b(gate21inter1), .O(G302));
nand2 gate22( .a(G27), .b(G28), .O(G305) );

  xor2  gate1009(.a(G30), .b(G29), .O(gate23inter0));
  nand2 gate1010(.a(gate23inter0), .b(s_66), .O(gate23inter1));
  and2  gate1011(.a(G30), .b(G29), .O(gate23inter2));
  inv1  gate1012(.a(s_66), .O(gate23inter3));
  inv1  gate1013(.a(s_67), .O(gate23inter4));
  nand2 gate1014(.a(gate23inter4), .b(gate23inter3), .O(gate23inter5));
  nor2  gate1015(.a(gate23inter5), .b(gate23inter2), .O(gate23inter6));
  inv1  gate1016(.a(G29), .O(gate23inter7));
  inv1  gate1017(.a(G30), .O(gate23inter8));
  nand2 gate1018(.a(gate23inter8), .b(gate23inter7), .O(gate23inter9));
  nand2 gate1019(.a(s_67), .b(gate23inter3), .O(gate23inter10));
  nor2  gate1020(.a(gate23inter10), .b(gate23inter9), .O(gate23inter11));
  nor2  gate1021(.a(gate23inter11), .b(gate23inter6), .O(gate23inter12));
  nand2 gate1022(.a(gate23inter12), .b(gate23inter1), .O(G308));
nand2 gate24( .a(G31), .b(G32), .O(G311) );

  xor2  gate939(.a(G5), .b(G1), .O(gate25inter0));
  nand2 gate940(.a(gate25inter0), .b(s_56), .O(gate25inter1));
  and2  gate941(.a(G5), .b(G1), .O(gate25inter2));
  inv1  gate942(.a(s_56), .O(gate25inter3));
  inv1  gate943(.a(s_57), .O(gate25inter4));
  nand2 gate944(.a(gate25inter4), .b(gate25inter3), .O(gate25inter5));
  nor2  gate945(.a(gate25inter5), .b(gate25inter2), .O(gate25inter6));
  inv1  gate946(.a(G1), .O(gate25inter7));
  inv1  gate947(.a(G5), .O(gate25inter8));
  nand2 gate948(.a(gate25inter8), .b(gate25inter7), .O(gate25inter9));
  nand2 gate949(.a(s_57), .b(gate25inter3), .O(gate25inter10));
  nor2  gate950(.a(gate25inter10), .b(gate25inter9), .O(gate25inter11));
  nor2  gate951(.a(gate25inter11), .b(gate25inter6), .O(gate25inter12));
  nand2 gate952(.a(gate25inter12), .b(gate25inter1), .O(G314));
nand2 gate26( .a(G9), .b(G13), .O(G317) );
nand2 gate27( .a(G2), .b(G6), .O(G320) );
nand2 gate28( .a(G10), .b(G14), .O(G323) );
nand2 gate29( .a(G3), .b(G7), .O(G326) );
nand2 gate30( .a(G11), .b(G15), .O(G329) );
nand2 gate31( .a(G4), .b(G8), .O(G332) );
nand2 gate32( .a(G12), .b(G16), .O(G335) );
nand2 gate33( .a(G17), .b(G21), .O(G338) );
nand2 gate34( .a(G25), .b(G29), .O(G341) );
nand2 gate35( .a(G18), .b(G22), .O(G344) );
nand2 gate36( .a(G26), .b(G30), .O(G347) );

  xor2  gate911(.a(G23), .b(G19), .O(gate37inter0));
  nand2 gate912(.a(gate37inter0), .b(s_52), .O(gate37inter1));
  and2  gate913(.a(G23), .b(G19), .O(gate37inter2));
  inv1  gate914(.a(s_52), .O(gate37inter3));
  inv1  gate915(.a(s_53), .O(gate37inter4));
  nand2 gate916(.a(gate37inter4), .b(gate37inter3), .O(gate37inter5));
  nor2  gate917(.a(gate37inter5), .b(gate37inter2), .O(gate37inter6));
  inv1  gate918(.a(G19), .O(gate37inter7));
  inv1  gate919(.a(G23), .O(gate37inter8));
  nand2 gate920(.a(gate37inter8), .b(gate37inter7), .O(gate37inter9));
  nand2 gate921(.a(s_53), .b(gate37inter3), .O(gate37inter10));
  nor2  gate922(.a(gate37inter10), .b(gate37inter9), .O(gate37inter11));
  nor2  gate923(.a(gate37inter11), .b(gate37inter6), .O(gate37inter12));
  nand2 gate924(.a(gate37inter12), .b(gate37inter1), .O(G350));
nand2 gate38( .a(G27), .b(G31), .O(G353) );
nand2 gate39( .a(G20), .b(G24), .O(G356) );
nand2 gate40( .a(G28), .b(G32), .O(G359) );
nand2 gate41( .a(G1), .b(G266), .O(G362) );
nand2 gate42( .a(G2), .b(G266), .O(G363) );
nand2 gate43( .a(G3), .b(G269), .O(G364) );
nand2 gate44( .a(G4), .b(G269), .O(G365) );

  xor2  gate967(.a(G272), .b(G5), .O(gate45inter0));
  nand2 gate968(.a(gate45inter0), .b(s_60), .O(gate45inter1));
  and2  gate969(.a(G272), .b(G5), .O(gate45inter2));
  inv1  gate970(.a(s_60), .O(gate45inter3));
  inv1  gate971(.a(s_61), .O(gate45inter4));
  nand2 gate972(.a(gate45inter4), .b(gate45inter3), .O(gate45inter5));
  nor2  gate973(.a(gate45inter5), .b(gate45inter2), .O(gate45inter6));
  inv1  gate974(.a(G5), .O(gate45inter7));
  inv1  gate975(.a(G272), .O(gate45inter8));
  nand2 gate976(.a(gate45inter8), .b(gate45inter7), .O(gate45inter9));
  nand2 gate977(.a(s_61), .b(gate45inter3), .O(gate45inter10));
  nor2  gate978(.a(gate45inter10), .b(gate45inter9), .O(gate45inter11));
  nor2  gate979(.a(gate45inter11), .b(gate45inter6), .O(gate45inter12));
  nand2 gate980(.a(gate45inter12), .b(gate45inter1), .O(G366));
nand2 gate46( .a(G6), .b(G272), .O(G367) );
nand2 gate47( .a(G7), .b(G275), .O(G368) );
nand2 gate48( .a(G8), .b(G275), .O(G369) );
nand2 gate49( .a(G9), .b(G278), .O(G370) );
nand2 gate50( .a(G10), .b(G278), .O(G371) );
nand2 gate51( .a(G11), .b(G281), .O(G372) );
nand2 gate52( .a(G12), .b(G281), .O(G373) );
nand2 gate53( .a(G13), .b(G284), .O(G374) );
nand2 gate54( .a(G14), .b(G284), .O(G375) );
nand2 gate55( .a(G15), .b(G287), .O(G376) );
nand2 gate56( .a(G16), .b(G287), .O(G377) );
nand2 gate57( .a(G17), .b(G290), .O(G378) );
nand2 gate58( .a(G18), .b(G290), .O(G379) );
nand2 gate59( .a(G19), .b(G293), .O(G380) );
nand2 gate60( .a(G20), .b(G293), .O(G381) );
nand2 gate61( .a(G21), .b(G296), .O(G382) );
nand2 gate62( .a(G22), .b(G296), .O(G383) );
nand2 gate63( .a(G23), .b(G299), .O(G384) );
nand2 gate64( .a(G24), .b(G299), .O(G385) );
nand2 gate65( .a(G25), .b(G302), .O(G386) );
nand2 gate66( .a(G26), .b(G302), .O(G387) );
nand2 gate67( .a(G27), .b(G305), .O(G388) );

  xor2  gate575(.a(G305), .b(G28), .O(gate68inter0));
  nand2 gate576(.a(gate68inter0), .b(s_4), .O(gate68inter1));
  and2  gate577(.a(G305), .b(G28), .O(gate68inter2));
  inv1  gate578(.a(s_4), .O(gate68inter3));
  inv1  gate579(.a(s_5), .O(gate68inter4));
  nand2 gate580(.a(gate68inter4), .b(gate68inter3), .O(gate68inter5));
  nor2  gate581(.a(gate68inter5), .b(gate68inter2), .O(gate68inter6));
  inv1  gate582(.a(G28), .O(gate68inter7));
  inv1  gate583(.a(G305), .O(gate68inter8));
  nand2 gate584(.a(gate68inter8), .b(gate68inter7), .O(gate68inter9));
  nand2 gate585(.a(s_5), .b(gate68inter3), .O(gate68inter10));
  nor2  gate586(.a(gate68inter10), .b(gate68inter9), .O(gate68inter11));
  nor2  gate587(.a(gate68inter11), .b(gate68inter6), .O(gate68inter12));
  nand2 gate588(.a(gate68inter12), .b(gate68inter1), .O(G389));
nand2 gate69( .a(G29), .b(G308), .O(G390) );
nand2 gate70( .a(G30), .b(G308), .O(G391) );
nand2 gate71( .a(G31), .b(G311), .O(G392) );
nand2 gate72( .a(G32), .b(G311), .O(G393) );
nand2 gate73( .a(G1), .b(G314), .O(G394) );
nand2 gate74( .a(G5), .b(G314), .O(G395) );
nand2 gate75( .a(G9), .b(G317), .O(G396) );
nand2 gate76( .a(G13), .b(G317), .O(G397) );
nand2 gate77( .a(G2), .b(G320), .O(G398) );
nand2 gate78( .a(G6), .b(G320), .O(G399) );
nand2 gate79( .a(G10), .b(G323), .O(G400) );
nand2 gate80( .a(G14), .b(G323), .O(G401) );
nand2 gate81( .a(G3), .b(G326), .O(G402) );
nand2 gate82( .a(G7), .b(G326), .O(G403) );
nand2 gate83( .a(G11), .b(G329), .O(G404) );
nand2 gate84( .a(G15), .b(G329), .O(G405) );
nand2 gate85( .a(G4), .b(G332), .O(G406) );

  xor2  gate981(.a(G332), .b(G8), .O(gate86inter0));
  nand2 gate982(.a(gate86inter0), .b(s_62), .O(gate86inter1));
  and2  gate983(.a(G332), .b(G8), .O(gate86inter2));
  inv1  gate984(.a(s_62), .O(gate86inter3));
  inv1  gate985(.a(s_63), .O(gate86inter4));
  nand2 gate986(.a(gate86inter4), .b(gate86inter3), .O(gate86inter5));
  nor2  gate987(.a(gate86inter5), .b(gate86inter2), .O(gate86inter6));
  inv1  gate988(.a(G8), .O(gate86inter7));
  inv1  gate989(.a(G332), .O(gate86inter8));
  nand2 gate990(.a(gate86inter8), .b(gate86inter7), .O(gate86inter9));
  nand2 gate991(.a(s_63), .b(gate86inter3), .O(gate86inter10));
  nor2  gate992(.a(gate86inter10), .b(gate86inter9), .O(gate86inter11));
  nor2  gate993(.a(gate86inter11), .b(gate86inter6), .O(gate86inter12));
  nand2 gate994(.a(gate86inter12), .b(gate86inter1), .O(G407));
nand2 gate87( .a(G12), .b(G335), .O(G408) );
nand2 gate88( .a(G16), .b(G335), .O(G409) );

  xor2  gate1065(.a(G338), .b(G17), .O(gate89inter0));
  nand2 gate1066(.a(gate89inter0), .b(s_74), .O(gate89inter1));
  and2  gate1067(.a(G338), .b(G17), .O(gate89inter2));
  inv1  gate1068(.a(s_74), .O(gate89inter3));
  inv1  gate1069(.a(s_75), .O(gate89inter4));
  nand2 gate1070(.a(gate89inter4), .b(gate89inter3), .O(gate89inter5));
  nor2  gate1071(.a(gate89inter5), .b(gate89inter2), .O(gate89inter6));
  inv1  gate1072(.a(G17), .O(gate89inter7));
  inv1  gate1073(.a(G338), .O(gate89inter8));
  nand2 gate1074(.a(gate89inter8), .b(gate89inter7), .O(gate89inter9));
  nand2 gate1075(.a(s_75), .b(gate89inter3), .O(gate89inter10));
  nor2  gate1076(.a(gate89inter10), .b(gate89inter9), .O(gate89inter11));
  nor2  gate1077(.a(gate89inter11), .b(gate89inter6), .O(gate89inter12));
  nand2 gate1078(.a(gate89inter12), .b(gate89inter1), .O(G410));
nand2 gate90( .a(G21), .b(G338), .O(G411) );

  xor2  gate841(.a(G341), .b(G25), .O(gate91inter0));
  nand2 gate842(.a(gate91inter0), .b(s_42), .O(gate91inter1));
  and2  gate843(.a(G341), .b(G25), .O(gate91inter2));
  inv1  gate844(.a(s_42), .O(gate91inter3));
  inv1  gate845(.a(s_43), .O(gate91inter4));
  nand2 gate846(.a(gate91inter4), .b(gate91inter3), .O(gate91inter5));
  nor2  gate847(.a(gate91inter5), .b(gate91inter2), .O(gate91inter6));
  inv1  gate848(.a(G25), .O(gate91inter7));
  inv1  gate849(.a(G341), .O(gate91inter8));
  nand2 gate850(.a(gate91inter8), .b(gate91inter7), .O(gate91inter9));
  nand2 gate851(.a(s_43), .b(gate91inter3), .O(gate91inter10));
  nor2  gate852(.a(gate91inter10), .b(gate91inter9), .O(gate91inter11));
  nor2  gate853(.a(gate91inter11), .b(gate91inter6), .O(gate91inter12));
  nand2 gate854(.a(gate91inter12), .b(gate91inter1), .O(G412));
nand2 gate92( .a(G29), .b(G341), .O(G413) );

  xor2  gate1149(.a(G344), .b(G18), .O(gate93inter0));
  nand2 gate1150(.a(gate93inter0), .b(s_86), .O(gate93inter1));
  and2  gate1151(.a(G344), .b(G18), .O(gate93inter2));
  inv1  gate1152(.a(s_86), .O(gate93inter3));
  inv1  gate1153(.a(s_87), .O(gate93inter4));
  nand2 gate1154(.a(gate93inter4), .b(gate93inter3), .O(gate93inter5));
  nor2  gate1155(.a(gate93inter5), .b(gate93inter2), .O(gate93inter6));
  inv1  gate1156(.a(G18), .O(gate93inter7));
  inv1  gate1157(.a(G344), .O(gate93inter8));
  nand2 gate1158(.a(gate93inter8), .b(gate93inter7), .O(gate93inter9));
  nand2 gate1159(.a(s_87), .b(gate93inter3), .O(gate93inter10));
  nor2  gate1160(.a(gate93inter10), .b(gate93inter9), .O(gate93inter11));
  nor2  gate1161(.a(gate93inter11), .b(gate93inter6), .O(gate93inter12));
  nand2 gate1162(.a(gate93inter12), .b(gate93inter1), .O(G414));
nand2 gate94( .a(G22), .b(G344), .O(G415) );

  xor2  gate1107(.a(G347), .b(G26), .O(gate95inter0));
  nand2 gate1108(.a(gate95inter0), .b(s_80), .O(gate95inter1));
  and2  gate1109(.a(G347), .b(G26), .O(gate95inter2));
  inv1  gate1110(.a(s_80), .O(gate95inter3));
  inv1  gate1111(.a(s_81), .O(gate95inter4));
  nand2 gate1112(.a(gate95inter4), .b(gate95inter3), .O(gate95inter5));
  nor2  gate1113(.a(gate95inter5), .b(gate95inter2), .O(gate95inter6));
  inv1  gate1114(.a(G26), .O(gate95inter7));
  inv1  gate1115(.a(G347), .O(gate95inter8));
  nand2 gate1116(.a(gate95inter8), .b(gate95inter7), .O(gate95inter9));
  nand2 gate1117(.a(s_81), .b(gate95inter3), .O(gate95inter10));
  nor2  gate1118(.a(gate95inter10), .b(gate95inter9), .O(gate95inter11));
  nor2  gate1119(.a(gate95inter11), .b(gate95inter6), .O(gate95inter12));
  nand2 gate1120(.a(gate95inter12), .b(gate95inter1), .O(G416));
nand2 gate96( .a(G30), .b(G347), .O(G417) );
nand2 gate97( .a(G19), .b(G350), .O(G418) );
nand2 gate98( .a(G23), .b(G350), .O(G419) );
nand2 gate99( .a(G27), .b(G353), .O(G420) );
nand2 gate100( .a(G31), .b(G353), .O(G421) );
nand2 gate101( .a(G20), .b(G356), .O(G422) );
nand2 gate102( .a(G24), .b(G356), .O(G423) );
nand2 gate103( .a(G28), .b(G359), .O(G424) );
nand2 gate104( .a(G32), .b(G359), .O(G425) );
nand2 gate105( .a(G362), .b(G363), .O(G426) );
nand2 gate106( .a(G364), .b(G365), .O(G429) );
nand2 gate107( .a(G366), .b(G367), .O(G432) );
nand2 gate108( .a(G368), .b(G369), .O(G435) );
nand2 gate109( .a(G370), .b(G371), .O(G438) );
nand2 gate110( .a(G372), .b(G373), .O(G441) );
nand2 gate111( .a(G374), .b(G375), .O(G444) );
nand2 gate112( .a(G376), .b(G377), .O(G447) );
nand2 gate113( .a(G378), .b(G379), .O(G450) );
nand2 gate114( .a(G380), .b(G381), .O(G453) );
nand2 gate115( .a(G382), .b(G383), .O(G456) );
nand2 gate116( .a(G384), .b(G385), .O(G459) );
nand2 gate117( .a(G386), .b(G387), .O(G462) );
nand2 gate118( .a(G388), .b(G389), .O(G465) );
nand2 gate119( .a(G390), .b(G391), .O(G468) );
nand2 gate120( .a(G392), .b(G393), .O(G471) );
nand2 gate121( .a(G394), .b(G395), .O(G474) );
nand2 gate122( .a(G396), .b(G397), .O(G477) );
nand2 gate123( .a(G398), .b(G399), .O(G480) );

  xor2  gate1163(.a(G401), .b(G400), .O(gate124inter0));
  nand2 gate1164(.a(gate124inter0), .b(s_88), .O(gate124inter1));
  and2  gate1165(.a(G401), .b(G400), .O(gate124inter2));
  inv1  gate1166(.a(s_88), .O(gate124inter3));
  inv1  gate1167(.a(s_89), .O(gate124inter4));
  nand2 gate1168(.a(gate124inter4), .b(gate124inter3), .O(gate124inter5));
  nor2  gate1169(.a(gate124inter5), .b(gate124inter2), .O(gate124inter6));
  inv1  gate1170(.a(G400), .O(gate124inter7));
  inv1  gate1171(.a(G401), .O(gate124inter8));
  nand2 gate1172(.a(gate124inter8), .b(gate124inter7), .O(gate124inter9));
  nand2 gate1173(.a(s_89), .b(gate124inter3), .O(gate124inter10));
  nor2  gate1174(.a(gate124inter10), .b(gate124inter9), .O(gate124inter11));
  nor2  gate1175(.a(gate124inter11), .b(gate124inter6), .O(gate124inter12));
  nand2 gate1176(.a(gate124inter12), .b(gate124inter1), .O(G483));
nand2 gate125( .a(G402), .b(G403), .O(G486) );
nand2 gate126( .a(G404), .b(G405), .O(G489) );
nand2 gate127( .a(G406), .b(G407), .O(G492) );
nand2 gate128( .a(G408), .b(G409), .O(G495) );
nand2 gate129( .a(G410), .b(G411), .O(G498) );
nand2 gate130( .a(G412), .b(G413), .O(G501) );
nand2 gate131( .a(G414), .b(G415), .O(G504) );
nand2 gate132( .a(G416), .b(G417), .O(G507) );
nand2 gate133( .a(G418), .b(G419), .O(G510) );

  xor2  gate673(.a(G421), .b(G420), .O(gate134inter0));
  nand2 gate674(.a(gate134inter0), .b(s_18), .O(gate134inter1));
  and2  gate675(.a(G421), .b(G420), .O(gate134inter2));
  inv1  gate676(.a(s_18), .O(gate134inter3));
  inv1  gate677(.a(s_19), .O(gate134inter4));
  nand2 gate678(.a(gate134inter4), .b(gate134inter3), .O(gate134inter5));
  nor2  gate679(.a(gate134inter5), .b(gate134inter2), .O(gate134inter6));
  inv1  gate680(.a(G420), .O(gate134inter7));
  inv1  gate681(.a(G421), .O(gate134inter8));
  nand2 gate682(.a(gate134inter8), .b(gate134inter7), .O(gate134inter9));
  nand2 gate683(.a(s_19), .b(gate134inter3), .O(gate134inter10));
  nor2  gate684(.a(gate134inter10), .b(gate134inter9), .O(gate134inter11));
  nor2  gate685(.a(gate134inter11), .b(gate134inter6), .O(gate134inter12));
  nand2 gate686(.a(gate134inter12), .b(gate134inter1), .O(G513));

  xor2  gate589(.a(G423), .b(G422), .O(gate135inter0));
  nand2 gate590(.a(gate135inter0), .b(s_6), .O(gate135inter1));
  and2  gate591(.a(G423), .b(G422), .O(gate135inter2));
  inv1  gate592(.a(s_6), .O(gate135inter3));
  inv1  gate593(.a(s_7), .O(gate135inter4));
  nand2 gate594(.a(gate135inter4), .b(gate135inter3), .O(gate135inter5));
  nor2  gate595(.a(gate135inter5), .b(gate135inter2), .O(gate135inter6));
  inv1  gate596(.a(G422), .O(gate135inter7));
  inv1  gate597(.a(G423), .O(gate135inter8));
  nand2 gate598(.a(gate135inter8), .b(gate135inter7), .O(gate135inter9));
  nand2 gate599(.a(s_7), .b(gate135inter3), .O(gate135inter10));
  nor2  gate600(.a(gate135inter10), .b(gate135inter9), .O(gate135inter11));
  nor2  gate601(.a(gate135inter11), .b(gate135inter6), .O(gate135inter12));
  nand2 gate602(.a(gate135inter12), .b(gate135inter1), .O(G516));
nand2 gate136( .a(G424), .b(G425), .O(G519) );

  xor2  gate561(.a(G429), .b(G426), .O(gate137inter0));
  nand2 gate562(.a(gate137inter0), .b(s_2), .O(gate137inter1));
  and2  gate563(.a(G429), .b(G426), .O(gate137inter2));
  inv1  gate564(.a(s_2), .O(gate137inter3));
  inv1  gate565(.a(s_3), .O(gate137inter4));
  nand2 gate566(.a(gate137inter4), .b(gate137inter3), .O(gate137inter5));
  nor2  gate567(.a(gate137inter5), .b(gate137inter2), .O(gate137inter6));
  inv1  gate568(.a(G426), .O(gate137inter7));
  inv1  gate569(.a(G429), .O(gate137inter8));
  nand2 gate570(.a(gate137inter8), .b(gate137inter7), .O(gate137inter9));
  nand2 gate571(.a(s_3), .b(gate137inter3), .O(gate137inter10));
  nor2  gate572(.a(gate137inter10), .b(gate137inter9), .O(gate137inter11));
  nor2  gate573(.a(gate137inter11), .b(gate137inter6), .O(gate137inter12));
  nand2 gate574(.a(gate137inter12), .b(gate137inter1), .O(G522));
nand2 gate138( .a(G432), .b(G435), .O(G525) );
nand2 gate139( .a(G438), .b(G441), .O(G528) );
nand2 gate140( .a(G444), .b(G447), .O(G531) );
nand2 gate141( .a(G450), .b(G453), .O(G534) );
nand2 gate142( .a(G456), .b(G459), .O(G537) );
nand2 gate143( .a(G462), .b(G465), .O(G540) );
nand2 gate144( .a(G468), .b(G471), .O(G543) );

  xor2  gate1051(.a(G477), .b(G474), .O(gate145inter0));
  nand2 gate1052(.a(gate145inter0), .b(s_72), .O(gate145inter1));
  and2  gate1053(.a(G477), .b(G474), .O(gate145inter2));
  inv1  gate1054(.a(s_72), .O(gate145inter3));
  inv1  gate1055(.a(s_73), .O(gate145inter4));
  nand2 gate1056(.a(gate145inter4), .b(gate145inter3), .O(gate145inter5));
  nor2  gate1057(.a(gate145inter5), .b(gate145inter2), .O(gate145inter6));
  inv1  gate1058(.a(G474), .O(gate145inter7));
  inv1  gate1059(.a(G477), .O(gate145inter8));
  nand2 gate1060(.a(gate145inter8), .b(gate145inter7), .O(gate145inter9));
  nand2 gate1061(.a(s_73), .b(gate145inter3), .O(gate145inter10));
  nor2  gate1062(.a(gate145inter10), .b(gate145inter9), .O(gate145inter11));
  nor2  gate1063(.a(gate145inter11), .b(gate145inter6), .O(gate145inter12));
  nand2 gate1064(.a(gate145inter12), .b(gate145inter1), .O(G546));
nand2 gate146( .a(G480), .b(G483), .O(G549) );
nand2 gate147( .a(G486), .b(G489), .O(G552) );
nand2 gate148( .a(G492), .b(G495), .O(G555) );
nand2 gate149( .a(G498), .b(G501), .O(G558) );
nand2 gate150( .a(G504), .b(G507), .O(G561) );
nand2 gate151( .a(G510), .b(G513), .O(G564) );
nand2 gate152( .a(G516), .b(G519), .O(G567) );
nand2 gate153( .a(G426), .b(G522), .O(G570) );
nand2 gate154( .a(G429), .b(G522), .O(G571) );
nand2 gate155( .a(G432), .b(G525), .O(G572) );
nand2 gate156( .a(G435), .b(G525), .O(G573) );
nand2 gate157( .a(G438), .b(G528), .O(G574) );
nand2 gate158( .a(G441), .b(G528), .O(G575) );
nand2 gate159( .a(G444), .b(G531), .O(G576) );
nand2 gate160( .a(G447), .b(G531), .O(G577) );

  xor2  gate715(.a(G534), .b(G450), .O(gate161inter0));
  nand2 gate716(.a(gate161inter0), .b(s_24), .O(gate161inter1));
  and2  gate717(.a(G534), .b(G450), .O(gate161inter2));
  inv1  gate718(.a(s_24), .O(gate161inter3));
  inv1  gate719(.a(s_25), .O(gate161inter4));
  nand2 gate720(.a(gate161inter4), .b(gate161inter3), .O(gate161inter5));
  nor2  gate721(.a(gate161inter5), .b(gate161inter2), .O(gate161inter6));
  inv1  gate722(.a(G450), .O(gate161inter7));
  inv1  gate723(.a(G534), .O(gate161inter8));
  nand2 gate724(.a(gate161inter8), .b(gate161inter7), .O(gate161inter9));
  nand2 gate725(.a(s_25), .b(gate161inter3), .O(gate161inter10));
  nor2  gate726(.a(gate161inter10), .b(gate161inter9), .O(gate161inter11));
  nor2  gate727(.a(gate161inter11), .b(gate161inter6), .O(gate161inter12));
  nand2 gate728(.a(gate161inter12), .b(gate161inter1), .O(G578));
nand2 gate162( .a(G453), .b(G534), .O(G579) );
nand2 gate163( .a(G456), .b(G537), .O(G580) );
nand2 gate164( .a(G459), .b(G537), .O(G581) );
nand2 gate165( .a(G462), .b(G540), .O(G582) );
nand2 gate166( .a(G465), .b(G540), .O(G583) );
nand2 gate167( .a(G468), .b(G543), .O(G584) );
nand2 gate168( .a(G471), .b(G543), .O(G585) );
nand2 gate169( .a(G474), .b(G546), .O(G586) );
nand2 gate170( .a(G477), .b(G546), .O(G587) );
nand2 gate171( .a(G480), .b(G549), .O(G588) );
nand2 gate172( .a(G483), .b(G549), .O(G589) );
nand2 gate173( .a(G486), .b(G552), .O(G590) );
nand2 gate174( .a(G489), .b(G552), .O(G591) );
nand2 gate175( .a(G492), .b(G555), .O(G592) );
nand2 gate176( .a(G495), .b(G555), .O(G593) );
nand2 gate177( .a(G498), .b(G558), .O(G594) );
nand2 gate178( .a(G501), .b(G558), .O(G595) );
nand2 gate179( .a(G504), .b(G561), .O(G596) );
nand2 gate180( .a(G507), .b(G561), .O(G597) );
nand2 gate181( .a(G510), .b(G564), .O(G598) );
nand2 gate182( .a(G513), .b(G564), .O(G599) );
nand2 gate183( .a(G516), .b(G567), .O(G600) );
nand2 gate184( .a(G519), .b(G567), .O(G601) );
nand2 gate185( .a(G570), .b(G571), .O(G602) );
nand2 gate186( .a(G572), .b(G573), .O(G607) );
nand2 gate187( .a(G574), .b(G575), .O(G612) );
nand2 gate188( .a(G576), .b(G577), .O(G617) );
nand2 gate189( .a(G578), .b(G579), .O(G622) );
nand2 gate190( .a(G580), .b(G581), .O(G627) );

  xor2  gate1093(.a(G583), .b(G582), .O(gate191inter0));
  nand2 gate1094(.a(gate191inter0), .b(s_78), .O(gate191inter1));
  and2  gate1095(.a(G583), .b(G582), .O(gate191inter2));
  inv1  gate1096(.a(s_78), .O(gate191inter3));
  inv1  gate1097(.a(s_79), .O(gate191inter4));
  nand2 gate1098(.a(gate191inter4), .b(gate191inter3), .O(gate191inter5));
  nor2  gate1099(.a(gate191inter5), .b(gate191inter2), .O(gate191inter6));
  inv1  gate1100(.a(G582), .O(gate191inter7));
  inv1  gate1101(.a(G583), .O(gate191inter8));
  nand2 gate1102(.a(gate191inter8), .b(gate191inter7), .O(gate191inter9));
  nand2 gate1103(.a(s_79), .b(gate191inter3), .O(gate191inter10));
  nor2  gate1104(.a(gate191inter10), .b(gate191inter9), .O(gate191inter11));
  nor2  gate1105(.a(gate191inter11), .b(gate191inter6), .O(gate191inter12));
  nand2 gate1106(.a(gate191inter12), .b(gate191inter1), .O(G632));
nand2 gate192( .a(G584), .b(G585), .O(G637) );
nand2 gate193( .a(G586), .b(G587), .O(G642) );

  xor2  gate757(.a(G589), .b(G588), .O(gate194inter0));
  nand2 gate758(.a(gate194inter0), .b(s_30), .O(gate194inter1));
  and2  gate759(.a(G589), .b(G588), .O(gate194inter2));
  inv1  gate760(.a(s_30), .O(gate194inter3));
  inv1  gate761(.a(s_31), .O(gate194inter4));
  nand2 gate762(.a(gate194inter4), .b(gate194inter3), .O(gate194inter5));
  nor2  gate763(.a(gate194inter5), .b(gate194inter2), .O(gate194inter6));
  inv1  gate764(.a(G588), .O(gate194inter7));
  inv1  gate765(.a(G589), .O(gate194inter8));
  nand2 gate766(.a(gate194inter8), .b(gate194inter7), .O(gate194inter9));
  nand2 gate767(.a(s_31), .b(gate194inter3), .O(gate194inter10));
  nor2  gate768(.a(gate194inter10), .b(gate194inter9), .O(gate194inter11));
  nor2  gate769(.a(gate194inter11), .b(gate194inter6), .O(gate194inter12));
  nand2 gate770(.a(gate194inter12), .b(gate194inter1), .O(G645));
nand2 gate195( .a(G590), .b(G591), .O(G648) );
nand2 gate196( .a(G592), .b(G593), .O(G651) );
nand2 gate197( .a(G594), .b(G595), .O(G654) );
nand2 gate198( .a(G596), .b(G597), .O(G657) );
nand2 gate199( .a(G598), .b(G599), .O(G660) );

  xor2  gate645(.a(G601), .b(G600), .O(gate200inter0));
  nand2 gate646(.a(gate200inter0), .b(s_14), .O(gate200inter1));
  and2  gate647(.a(G601), .b(G600), .O(gate200inter2));
  inv1  gate648(.a(s_14), .O(gate200inter3));
  inv1  gate649(.a(s_15), .O(gate200inter4));
  nand2 gate650(.a(gate200inter4), .b(gate200inter3), .O(gate200inter5));
  nor2  gate651(.a(gate200inter5), .b(gate200inter2), .O(gate200inter6));
  inv1  gate652(.a(G600), .O(gate200inter7));
  inv1  gate653(.a(G601), .O(gate200inter8));
  nand2 gate654(.a(gate200inter8), .b(gate200inter7), .O(gate200inter9));
  nand2 gate655(.a(s_15), .b(gate200inter3), .O(gate200inter10));
  nor2  gate656(.a(gate200inter10), .b(gate200inter9), .O(gate200inter11));
  nor2  gate657(.a(gate200inter11), .b(gate200inter6), .O(gate200inter12));
  nand2 gate658(.a(gate200inter12), .b(gate200inter1), .O(G663));
nand2 gate201( .a(G602), .b(G607), .O(G666) );
nand2 gate202( .a(G612), .b(G617), .O(G669) );
nand2 gate203( .a(G602), .b(G612), .O(G672) );
nand2 gate204( .a(G607), .b(G617), .O(G675) );
nand2 gate205( .a(G622), .b(G627), .O(G678) );
nand2 gate206( .a(G632), .b(G637), .O(G681) );

  xor2  gate869(.a(G632), .b(G622), .O(gate207inter0));
  nand2 gate870(.a(gate207inter0), .b(s_46), .O(gate207inter1));
  and2  gate871(.a(G632), .b(G622), .O(gate207inter2));
  inv1  gate872(.a(s_46), .O(gate207inter3));
  inv1  gate873(.a(s_47), .O(gate207inter4));
  nand2 gate874(.a(gate207inter4), .b(gate207inter3), .O(gate207inter5));
  nor2  gate875(.a(gate207inter5), .b(gate207inter2), .O(gate207inter6));
  inv1  gate876(.a(G622), .O(gate207inter7));
  inv1  gate877(.a(G632), .O(gate207inter8));
  nand2 gate878(.a(gate207inter8), .b(gate207inter7), .O(gate207inter9));
  nand2 gate879(.a(s_47), .b(gate207inter3), .O(gate207inter10));
  nor2  gate880(.a(gate207inter10), .b(gate207inter9), .O(gate207inter11));
  nor2  gate881(.a(gate207inter11), .b(gate207inter6), .O(gate207inter12));
  nand2 gate882(.a(gate207inter12), .b(gate207inter1), .O(G684));
nand2 gate208( .a(G627), .b(G637), .O(G687) );
nand2 gate209( .a(G602), .b(G666), .O(G690) );
nand2 gate210( .a(G607), .b(G666), .O(G691) );
nand2 gate211( .a(G612), .b(G669), .O(G692) );
nand2 gate212( .a(G617), .b(G669), .O(G693) );
nand2 gate213( .a(G602), .b(G672), .O(G694) );
nand2 gate214( .a(G612), .b(G672), .O(G695) );
nand2 gate215( .a(G607), .b(G675), .O(G696) );
nand2 gate216( .a(G617), .b(G675), .O(G697) );
nand2 gate217( .a(G622), .b(G678), .O(G698) );
nand2 gate218( .a(G627), .b(G678), .O(G699) );
nand2 gate219( .a(G632), .b(G681), .O(G700) );
nand2 gate220( .a(G637), .b(G681), .O(G701) );

  xor2  gate547(.a(G684), .b(G622), .O(gate221inter0));
  nand2 gate548(.a(gate221inter0), .b(s_0), .O(gate221inter1));
  and2  gate549(.a(G684), .b(G622), .O(gate221inter2));
  inv1  gate550(.a(s_0), .O(gate221inter3));
  inv1  gate551(.a(s_1), .O(gate221inter4));
  nand2 gate552(.a(gate221inter4), .b(gate221inter3), .O(gate221inter5));
  nor2  gate553(.a(gate221inter5), .b(gate221inter2), .O(gate221inter6));
  inv1  gate554(.a(G622), .O(gate221inter7));
  inv1  gate555(.a(G684), .O(gate221inter8));
  nand2 gate556(.a(gate221inter8), .b(gate221inter7), .O(gate221inter9));
  nand2 gate557(.a(s_1), .b(gate221inter3), .O(gate221inter10));
  nor2  gate558(.a(gate221inter10), .b(gate221inter9), .O(gate221inter11));
  nor2  gate559(.a(gate221inter11), .b(gate221inter6), .O(gate221inter12));
  nand2 gate560(.a(gate221inter12), .b(gate221inter1), .O(G702));
nand2 gate222( .a(G632), .b(G684), .O(G703) );
nand2 gate223( .a(G627), .b(G687), .O(G704) );
nand2 gate224( .a(G637), .b(G687), .O(G705) );

  xor2  gate827(.a(G691), .b(G690), .O(gate225inter0));
  nand2 gate828(.a(gate225inter0), .b(s_40), .O(gate225inter1));
  and2  gate829(.a(G691), .b(G690), .O(gate225inter2));
  inv1  gate830(.a(s_40), .O(gate225inter3));
  inv1  gate831(.a(s_41), .O(gate225inter4));
  nand2 gate832(.a(gate225inter4), .b(gate225inter3), .O(gate225inter5));
  nor2  gate833(.a(gate225inter5), .b(gate225inter2), .O(gate225inter6));
  inv1  gate834(.a(G690), .O(gate225inter7));
  inv1  gate835(.a(G691), .O(gate225inter8));
  nand2 gate836(.a(gate225inter8), .b(gate225inter7), .O(gate225inter9));
  nand2 gate837(.a(s_41), .b(gate225inter3), .O(gate225inter10));
  nor2  gate838(.a(gate225inter10), .b(gate225inter9), .O(gate225inter11));
  nor2  gate839(.a(gate225inter11), .b(gate225inter6), .O(gate225inter12));
  nand2 gate840(.a(gate225inter12), .b(gate225inter1), .O(G706));
nand2 gate226( .a(G692), .b(G693), .O(G709) );
nand2 gate227( .a(G694), .b(G695), .O(G712) );
nand2 gate228( .a(G696), .b(G697), .O(G715) );
nand2 gate229( .a(G698), .b(G699), .O(G718) );
nand2 gate230( .a(G700), .b(G701), .O(G721) );

  xor2  gate631(.a(G703), .b(G702), .O(gate231inter0));
  nand2 gate632(.a(gate231inter0), .b(s_12), .O(gate231inter1));
  and2  gate633(.a(G703), .b(G702), .O(gate231inter2));
  inv1  gate634(.a(s_12), .O(gate231inter3));
  inv1  gate635(.a(s_13), .O(gate231inter4));
  nand2 gate636(.a(gate231inter4), .b(gate231inter3), .O(gate231inter5));
  nor2  gate637(.a(gate231inter5), .b(gate231inter2), .O(gate231inter6));
  inv1  gate638(.a(G702), .O(gate231inter7));
  inv1  gate639(.a(G703), .O(gate231inter8));
  nand2 gate640(.a(gate231inter8), .b(gate231inter7), .O(gate231inter9));
  nand2 gate641(.a(s_13), .b(gate231inter3), .O(gate231inter10));
  nor2  gate642(.a(gate231inter10), .b(gate231inter9), .O(gate231inter11));
  nor2  gate643(.a(gate231inter11), .b(gate231inter6), .O(gate231inter12));
  nand2 gate644(.a(gate231inter12), .b(gate231inter1), .O(G724));
nand2 gate232( .a(G704), .b(G705), .O(G727) );
nand2 gate233( .a(G242), .b(G718), .O(G730) );

  xor2  gate813(.a(G721), .b(G245), .O(gate234inter0));
  nand2 gate814(.a(gate234inter0), .b(s_38), .O(gate234inter1));
  and2  gate815(.a(G721), .b(G245), .O(gate234inter2));
  inv1  gate816(.a(s_38), .O(gate234inter3));
  inv1  gate817(.a(s_39), .O(gate234inter4));
  nand2 gate818(.a(gate234inter4), .b(gate234inter3), .O(gate234inter5));
  nor2  gate819(.a(gate234inter5), .b(gate234inter2), .O(gate234inter6));
  inv1  gate820(.a(G245), .O(gate234inter7));
  inv1  gate821(.a(G721), .O(gate234inter8));
  nand2 gate822(.a(gate234inter8), .b(gate234inter7), .O(gate234inter9));
  nand2 gate823(.a(s_39), .b(gate234inter3), .O(gate234inter10));
  nor2  gate824(.a(gate234inter10), .b(gate234inter9), .O(gate234inter11));
  nor2  gate825(.a(gate234inter11), .b(gate234inter6), .O(gate234inter12));
  nand2 gate826(.a(gate234inter12), .b(gate234inter1), .O(G733));
nand2 gate235( .a(G248), .b(G724), .O(G736) );
nand2 gate236( .a(G251), .b(G727), .O(G739) );
nand2 gate237( .a(G254), .b(G706), .O(G742) );
nand2 gate238( .a(G257), .b(G709), .O(G745) );
nand2 gate239( .a(G260), .b(G712), .O(G748) );
nand2 gate240( .a(G263), .b(G715), .O(G751) );
nand2 gate241( .a(G242), .b(G730), .O(G754) );
nand2 gate242( .a(G718), .b(G730), .O(G755) );
nand2 gate243( .a(G245), .b(G733), .O(G756) );
nand2 gate244( .a(G721), .b(G733), .O(G757) );
nand2 gate245( .a(G248), .b(G736), .O(G758) );
nand2 gate246( .a(G724), .b(G736), .O(G759) );
nand2 gate247( .a(G251), .b(G739), .O(G760) );
nand2 gate248( .a(G727), .b(G739), .O(G761) );
nand2 gate249( .a(G254), .b(G742), .O(G762) );

  xor2  gate701(.a(G742), .b(G706), .O(gate250inter0));
  nand2 gate702(.a(gate250inter0), .b(s_22), .O(gate250inter1));
  and2  gate703(.a(G742), .b(G706), .O(gate250inter2));
  inv1  gate704(.a(s_22), .O(gate250inter3));
  inv1  gate705(.a(s_23), .O(gate250inter4));
  nand2 gate706(.a(gate250inter4), .b(gate250inter3), .O(gate250inter5));
  nor2  gate707(.a(gate250inter5), .b(gate250inter2), .O(gate250inter6));
  inv1  gate708(.a(G706), .O(gate250inter7));
  inv1  gate709(.a(G742), .O(gate250inter8));
  nand2 gate710(.a(gate250inter8), .b(gate250inter7), .O(gate250inter9));
  nand2 gate711(.a(s_23), .b(gate250inter3), .O(gate250inter10));
  nor2  gate712(.a(gate250inter10), .b(gate250inter9), .O(gate250inter11));
  nor2  gate713(.a(gate250inter11), .b(gate250inter6), .O(gate250inter12));
  nand2 gate714(.a(gate250inter12), .b(gate250inter1), .O(G763));
nand2 gate251( .a(G257), .b(G745), .O(G764) );
nand2 gate252( .a(G709), .b(G745), .O(G765) );
nand2 gate253( .a(G260), .b(G748), .O(G766) );
nand2 gate254( .a(G712), .b(G748), .O(G767) );

  xor2  gate897(.a(G751), .b(G263), .O(gate255inter0));
  nand2 gate898(.a(gate255inter0), .b(s_50), .O(gate255inter1));
  and2  gate899(.a(G751), .b(G263), .O(gate255inter2));
  inv1  gate900(.a(s_50), .O(gate255inter3));
  inv1  gate901(.a(s_51), .O(gate255inter4));
  nand2 gate902(.a(gate255inter4), .b(gate255inter3), .O(gate255inter5));
  nor2  gate903(.a(gate255inter5), .b(gate255inter2), .O(gate255inter6));
  inv1  gate904(.a(G263), .O(gate255inter7));
  inv1  gate905(.a(G751), .O(gate255inter8));
  nand2 gate906(.a(gate255inter8), .b(gate255inter7), .O(gate255inter9));
  nand2 gate907(.a(s_51), .b(gate255inter3), .O(gate255inter10));
  nor2  gate908(.a(gate255inter10), .b(gate255inter9), .O(gate255inter11));
  nor2  gate909(.a(gate255inter11), .b(gate255inter6), .O(gate255inter12));
  nand2 gate910(.a(gate255inter12), .b(gate255inter1), .O(G768));
nand2 gate256( .a(G715), .b(G751), .O(G769) );

  xor2  gate1023(.a(G755), .b(G754), .O(gate257inter0));
  nand2 gate1024(.a(gate257inter0), .b(s_68), .O(gate257inter1));
  and2  gate1025(.a(G755), .b(G754), .O(gate257inter2));
  inv1  gate1026(.a(s_68), .O(gate257inter3));
  inv1  gate1027(.a(s_69), .O(gate257inter4));
  nand2 gate1028(.a(gate257inter4), .b(gate257inter3), .O(gate257inter5));
  nor2  gate1029(.a(gate257inter5), .b(gate257inter2), .O(gate257inter6));
  inv1  gate1030(.a(G754), .O(gate257inter7));
  inv1  gate1031(.a(G755), .O(gate257inter8));
  nand2 gate1032(.a(gate257inter8), .b(gate257inter7), .O(gate257inter9));
  nand2 gate1033(.a(s_69), .b(gate257inter3), .O(gate257inter10));
  nor2  gate1034(.a(gate257inter10), .b(gate257inter9), .O(gate257inter11));
  nor2  gate1035(.a(gate257inter11), .b(gate257inter6), .O(gate257inter12));
  nand2 gate1036(.a(gate257inter12), .b(gate257inter1), .O(G770));
nand2 gate258( .a(G756), .b(G757), .O(G773) );
nand2 gate259( .a(G758), .b(G759), .O(G776) );
nand2 gate260( .a(G760), .b(G761), .O(G779) );

  xor2  gate1177(.a(G763), .b(G762), .O(gate261inter0));
  nand2 gate1178(.a(gate261inter0), .b(s_90), .O(gate261inter1));
  and2  gate1179(.a(G763), .b(G762), .O(gate261inter2));
  inv1  gate1180(.a(s_90), .O(gate261inter3));
  inv1  gate1181(.a(s_91), .O(gate261inter4));
  nand2 gate1182(.a(gate261inter4), .b(gate261inter3), .O(gate261inter5));
  nor2  gate1183(.a(gate261inter5), .b(gate261inter2), .O(gate261inter6));
  inv1  gate1184(.a(G762), .O(gate261inter7));
  inv1  gate1185(.a(G763), .O(gate261inter8));
  nand2 gate1186(.a(gate261inter8), .b(gate261inter7), .O(gate261inter9));
  nand2 gate1187(.a(s_91), .b(gate261inter3), .O(gate261inter10));
  nor2  gate1188(.a(gate261inter10), .b(gate261inter9), .O(gate261inter11));
  nor2  gate1189(.a(gate261inter11), .b(gate261inter6), .O(gate261inter12));
  nand2 gate1190(.a(gate261inter12), .b(gate261inter1), .O(G782));
nand2 gate262( .a(G764), .b(G765), .O(G785) );
nand2 gate263( .a(G766), .b(G767), .O(G788) );
nand2 gate264( .a(G768), .b(G769), .O(G791) );
nand2 gate265( .a(G642), .b(G770), .O(G794) );
nand2 gate266( .a(G645), .b(G773), .O(G797) );
nand2 gate267( .a(G648), .b(G776), .O(G800) );
nand2 gate268( .a(G651), .b(G779), .O(G803) );
nand2 gate269( .a(G654), .b(G782), .O(G806) );
nand2 gate270( .a(G657), .b(G785), .O(G809) );
nand2 gate271( .a(G660), .b(G788), .O(G812) );
nand2 gate272( .a(G663), .b(G791), .O(G815) );

  xor2  gate1037(.a(G794), .b(G642), .O(gate273inter0));
  nand2 gate1038(.a(gate273inter0), .b(s_70), .O(gate273inter1));
  and2  gate1039(.a(G794), .b(G642), .O(gate273inter2));
  inv1  gate1040(.a(s_70), .O(gate273inter3));
  inv1  gate1041(.a(s_71), .O(gate273inter4));
  nand2 gate1042(.a(gate273inter4), .b(gate273inter3), .O(gate273inter5));
  nor2  gate1043(.a(gate273inter5), .b(gate273inter2), .O(gate273inter6));
  inv1  gate1044(.a(G642), .O(gate273inter7));
  inv1  gate1045(.a(G794), .O(gate273inter8));
  nand2 gate1046(.a(gate273inter8), .b(gate273inter7), .O(gate273inter9));
  nand2 gate1047(.a(s_71), .b(gate273inter3), .O(gate273inter10));
  nor2  gate1048(.a(gate273inter10), .b(gate273inter9), .O(gate273inter11));
  nor2  gate1049(.a(gate273inter11), .b(gate273inter6), .O(gate273inter12));
  nand2 gate1050(.a(gate273inter12), .b(gate273inter1), .O(G818));
nand2 gate274( .a(G770), .b(G794), .O(G819) );
nand2 gate275( .a(G645), .b(G797), .O(G820) );
nand2 gate276( .a(G773), .b(G797), .O(G821) );
nand2 gate277( .a(G648), .b(G800), .O(G822) );
nand2 gate278( .a(G776), .b(G800), .O(G823) );
nand2 gate279( .a(G651), .b(G803), .O(G824) );
nand2 gate280( .a(G779), .b(G803), .O(G825) );
nand2 gate281( .a(G654), .b(G806), .O(G826) );
nand2 gate282( .a(G782), .b(G806), .O(G827) );
nand2 gate283( .a(G657), .b(G809), .O(G828) );
nand2 gate284( .a(G785), .b(G809), .O(G829) );
nand2 gate285( .a(G660), .b(G812), .O(G830) );
nand2 gate286( .a(G788), .b(G812), .O(G831) );
nand2 gate287( .a(G663), .b(G815), .O(G832) );
nand2 gate288( .a(G791), .b(G815), .O(G833) );
nand2 gate289( .a(G818), .b(G819), .O(G834) );
nand2 gate290( .a(G820), .b(G821), .O(G847) );
nand2 gate291( .a(G822), .b(G823), .O(G860) );
nand2 gate292( .a(G824), .b(G825), .O(G873) );
nand2 gate293( .a(G828), .b(G829), .O(G886) );
nand2 gate294( .a(G832), .b(G833), .O(G899) );
nand2 gate295( .a(G830), .b(G831), .O(G912) );
nand2 gate296( .a(G826), .b(G827), .O(G925) );
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );
nand2 gate387( .a(G1), .b(G1036), .O(G1132) );
nand2 gate388( .a(G2), .b(G1039), .O(G1135) );
nand2 gate389( .a(G3), .b(G1042), .O(G1138) );
nand2 gate390( .a(G4), .b(G1045), .O(G1141) );
nand2 gate391( .a(G5), .b(G1048), .O(G1144) );
nand2 gate392( .a(G6), .b(G1051), .O(G1147) );
nand2 gate393( .a(G7), .b(G1054), .O(G1150) );

  xor2  gate995(.a(G1057), .b(G8), .O(gate394inter0));
  nand2 gate996(.a(gate394inter0), .b(s_64), .O(gate394inter1));
  and2  gate997(.a(G1057), .b(G8), .O(gate394inter2));
  inv1  gate998(.a(s_64), .O(gate394inter3));
  inv1  gate999(.a(s_65), .O(gate394inter4));
  nand2 gate1000(.a(gate394inter4), .b(gate394inter3), .O(gate394inter5));
  nor2  gate1001(.a(gate394inter5), .b(gate394inter2), .O(gate394inter6));
  inv1  gate1002(.a(G8), .O(gate394inter7));
  inv1  gate1003(.a(G1057), .O(gate394inter8));
  nand2 gate1004(.a(gate394inter8), .b(gate394inter7), .O(gate394inter9));
  nand2 gate1005(.a(s_65), .b(gate394inter3), .O(gate394inter10));
  nor2  gate1006(.a(gate394inter10), .b(gate394inter9), .O(gate394inter11));
  nor2  gate1007(.a(gate394inter11), .b(gate394inter6), .O(gate394inter12));
  nand2 gate1008(.a(gate394inter12), .b(gate394inter1), .O(G1153));
nand2 gate395( .a(G9), .b(G1060), .O(G1156) );
nand2 gate396( .a(G10), .b(G1063), .O(G1159) );
nand2 gate397( .a(G11), .b(G1066), .O(G1162) );

  xor2  gate883(.a(G1069), .b(G12), .O(gate398inter0));
  nand2 gate884(.a(gate398inter0), .b(s_48), .O(gate398inter1));
  and2  gate885(.a(G1069), .b(G12), .O(gate398inter2));
  inv1  gate886(.a(s_48), .O(gate398inter3));
  inv1  gate887(.a(s_49), .O(gate398inter4));
  nand2 gate888(.a(gate398inter4), .b(gate398inter3), .O(gate398inter5));
  nor2  gate889(.a(gate398inter5), .b(gate398inter2), .O(gate398inter6));
  inv1  gate890(.a(G12), .O(gate398inter7));
  inv1  gate891(.a(G1069), .O(gate398inter8));
  nand2 gate892(.a(gate398inter8), .b(gate398inter7), .O(gate398inter9));
  nand2 gate893(.a(s_49), .b(gate398inter3), .O(gate398inter10));
  nor2  gate894(.a(gate398inter10), .b(gate398inter9), .O(gate398inter11));
  nor2  gate895(.a(gate398inter11), .b(gate398inter6), .O(gate398inter12));
  nand2 gate896(.a(gate398inter12), .b(gate398inter1), .O(G1165));
nand2 gate399( .a(G13), .b(G1072), .O(G1168) );

  xor2  gate687(.a(G1075), .b(G14), .O(gate400inter0));
  nand2 gate688(.a(gate400inter0), .b(s_20), .O(gate400inter1));
  and2  gate689(.a(G1075), .b(G14), .O(gate400inter2));
  inv1  gate690(.a(s_20), .O(gate400inter3));
  inv1  gate691(.a(s_21), .O(gate400inter4));
  nand2 gate692(.a(gate400inter4), .b(gate400inter3), .O(gate400inter5));
  nor2  gate693(.a(gate400inter5), .b(gate400inter2), .O(gate400inter6));
  inv1  gate694(.a(G14), .O(gate400inter7));
  inv1  gate695(.a(G1075), .O(gate400inter8));
  nand2 gate696(.a(gate400inter8), .b(gate400inter7), .O(gate400inter9));
  nand2 gate697(.a(s_21), .b(gate400inter3), .O(gate400inter10));
  nor2  gate698(.a(gate400inter10), .b(gate400inter9), .O(gate400inter11));
  nor2  gate699(.a(gate400inter11), .b(gate400inter6), .O(gate400inter12));
  nand2 gate700(.a(gate400inter12), .b(gate400inter1), .O(G1171));
nand2 gate401( .a(G15), .b(G1078), .O(G1174) );
nand2 gate402( .a(G16), .b(G1081), .O(G1177) );
nand2 gate403( .a(G17), .b(G1084), .O(G1180) );
nand2 gate404( .a(G18), .b(G1087), .O(G1183) );
nand2 gate405( .a(G19), .b(G1090), .O(G1186) );
nand2 gate406( .a(G20), .b(G1093), .O(G1189) );
nand2 gate407( .a(G21), .b(G1096), .O(G1192) );
nand2 gate408( .a(G22), .b(G1099), .O(G1195) );
nand2 gate409( .a(G23), .b(G1102), .O(G1198) );
nand2 gate410( .a(G24), .b(G1105), .O(G1201) );
nand2 gate411( .a(G25), .b(G1108), .O(G1204) );
nand2 gate412( .a(G26), .b(G1111), .O(G1207) );
nand2 gate413( .a(G27), .b(G1114), .O(G1210) );
nand2 gate414( .a(G28), .b(G1117), .O(G1213) );
nand2 gate415( .a(G29), .b(G1120), .O(G1216) );
nand2 gate416( .a(G30), .b(G1123), .O(G1219) );

  xor2  gate925(.a(G1126), .b(G31), .O(gate417inter0));
  nand2 gate926(.a(gate417inter0), .b(s_54), .O(gate417inter1));
  and2  gate927(.a(G1126), .b(G31), .O(gate417inter2));
  inv1  gate928(.a(s_54), .O(gate417inter3));
  inv1  gate929(.a(s_55), .O(gate417inter4));
  nand2 gate930(.a(gate417inter4), .b(gate417inter3), .O(gate417inter5));
  nor2  gate931(.a(gate417inter5), .b(gate417inter2), .O(gate417inter6));
  inv1  gate932(.a(G31), .O(gate417inter7));
  inv1  gate933(.a(G1126), .O(gate417inter8));
  nand2 gate934(.a(gate417inter8), .b(gate417inter7), .O(gate417inter9));
  nand2 gate935(.a(s_55), .b(gate417inter3), .O(gate417inter10));
  nor2  gate936(.a(gate417inter10), .b(gate417inter9), .O(gate417inter11));
  nor2  gate937(.a(gate417inter11), .b(gate417inter6), .O(gate417inter12));
  nand2 gate938(.a(gate417inter12), .b(gate417inter1), .O(G1222));
nand2 gate418( .a(G32), .b(G1129), .O(G1225) );
nand2 gate419( .a(G1), .b(G1132), .O(G1228) );
nand2 gate420( .a(G1036), .b(G1132), .O(G1229) );
nand2 gate421( .a(G2), .b(G1135), .O(G1230) );

  xor2  gate1135(.a(G1135), .b(G1039), .O(gate422inter0));
  nand2 gate1136(.a(gate422inter0), .b(s_84), .O(gate422inter1));
  and2  gate1137(.a(G1135), .b(G1039), .O(gate422inter2));
  inv1  gate1138(.a(s_84), .O(gate422inter3));
  inv1  gate1139(.a(s_85), .O(gate422inter4));
  nand2 gate1140(.a(gate422inter4), .b(gate422inter3), .O(gate422inter5));
  nor2  gate1141(.a(gate422inter5), .b(gate422inter2), .O(gate422inter6));
  inv1  gate1142(.a(G1039), .O(gate422inter7));
  inv1  gate1143(.a(G1135), .O(gate422inter8));
  nand2 gate1144(.a(gate422inter8), .b(gate422inter7), .O(gate422inter9));
  nand2 gate1145(.a(s_85), .b(gate422inter3), .O(gate422inter10));
  nor2  gate1146(.a(gate422inter10), .b(gate422inter9), .O(gate422inter11));
  nor2  gate1147(.a(gate422inter11), .b(gate422inter6), .O(gate422inter12));
  nand2 gate1148(.a(gate422inter12), .b(gate422inter1), .O(G1231));

  xor2  gate953(.a(G1138), .b(G3), .O(gate423inter0));
  nand2 gate954(.a(gate423inter0), .b(s_58), .O(gate423inter1));
  and2  gate955(.a(G1138), .b(G3), .O(gate423inter2));
  inv1  gate956(.a(s_58), .O(gate423inter3));
  inv1  gate957(.a(s_59), .O(gate423inter4));
  nand2 gate958(.a(gate423inter4), .b(gate423inter3), .O(gate423inter5));
  nor2  gate959(.a(gate423inter5), .b(gate423inter2), .O(gate423inter6));
  inv1  gate960(.a(G3), .O(gate423inter7));
  inv1  gate961(.a(G1138), .O(gate423inter8));
  nand2 gate962(.a(gate423inter8), .b(gate423inter7), .O(gate423inter9));
  nand2 gate963(.a(s_59), .b(gate423inter3), .O(gate423inter10));
  nor2  gate964(.a(gate423inter10), .b(gate423inter9), .O(gate423inter11));
  nor2  gate965(.a(gate423inter11), .b(gate423inter6), .O(gate423inter12));
  nand2 gate966(.a(gate423inter12), .b(gate423inter1), .O(G1232));
nand2 gate424( .a(G1042), .b(G1138), .O(G1233) );
nand2 gate425( .a(G4), .b(G1141), .O(G1234) );
nand2 gate426( .a(G1045), .b(G1141), .O(G1235) );
nand2 gate427( .a(G5), .b(G1144), .O(G1236) );
nand2 gate428( .a(G1048), .b(G1144), .O(G1237) );
nand2 gate429( .a(G6), .b(G1147), .O(G1238) );
nand2 gate430( .a(G1051), .b(G1147), .O(G1239) );
nand2 gate431( .a(G7), .b(G1150), .O(G1240) );
nand2 gate432( .a(G1054), .b(G1150), .O(G1241) );
nand2 gate433( .a(G8), .b(G1153), .O(G1242) );
nand2 gate434( .a(G1057), .b(G1153), .O(G1243) );
nand2 gate435( .a(G9), .b(G1156), .O(G1244) );
nand2 gate436( .a(G1060), .b(G1156), .O(G1245) );
nand2 gate437( .a(G10), .b(G1159), .O(G1246) );
nand2 gate438( .a(G1063), .b(G1159), .O(G1247) );
nand2 gate439( .a(G11), .b(G1162), .O(G1248) );
nand2 gate440( .a(G1066), .b(G1162), .O(G1249) );
nand2 gate441( .a(G12), .b(G1165), .O(G1250) );
nand2 gate442( .a(G1069), .b(G1165), .O(G1251) );

  xor2  gate771(.a(G1168), .b(G13), .O(gate443inter0));
  nand2 gate772(.a(gate443inter0), .b(s_32), .O(gate443inter1));
  and2  gate773(.a(G1168), .b(G13), .O(gate443inter2));
  inv1  gate774(.a(s_32), .O(gate443inter3));
  inv1  gate775(.a(s_33), .O(gate443inter4));
  nand2 gate776(.a(gate443inter4), .b(gate443inter3), .O(gate443inter5));
  nor2  gate777(.a(gate443inter5), .b(gate443inter2), .O(gate443inter6));
  inv1  gate778(.a(G13), .O(gate443inter7));
  inv1  gate779(.a(G1168), .O(gate443inter8));
  nand2 gate780(.a(gate443inter8), .b(gate443inter7), .O(gate443inter9));
  nand2 gate781(.a(s_33), .b(gate443inter3), .O(gate443inter10));
  nor2  gate782(.a(gate443inter10), .b(gate443inter9), .O(gate443inter11));
  nor2  gate783(.a(gate443inter11), .b(gate443inter6), .O(gate443inter12));
  nand2 gate784(.a(gate443inter12), .b(gate443inter1), .O(G1252));
nand2 gate444( .a(G1072), .b(G1168), .O(G1253) );
nand2 gate445( .a(G14), .b(G1171), .O(G1254) );
nand2 gate446( .a(G1075), .b(G1171), .O(G1255) );
nand2 gate447( .a(G15), .b(G1174), .O(G1256) );
nand2 gate448( .a(G1078), .b(G1174), .O(G1257) );
nand2 gate449( .a(G16), .b(G1177), .O(G1258) );
nand2 gate450( .a(G1081), .b(G1177), .O(G1259) );
nand2 gate451( .a(G17), .b(G1180), .O(G1260) );
nand2 gate452( .a(G1084), .b(G1180), .O(G1261) );
nand2 gate453( .a(G18), .b(G1183), .O(G1262) );
nand2 gate454( .a(G1087), .b(G1183), .O(G1263) );
nand2 gate455( .a(G19), .b(G1186), .O(G1264) );
nand2 gate456( .a(G1090), .b(G1186), .O(G1265) );
nand2 gate457( .a(G20), .b(G1189), .O(G1266) );
nand2 gate458( .a(G1093), .b(G1189), .O(G1267) );
nand2 gate459( .a(G21), .b(G1192), .O(G1268) );
nand2 gate460( .a(G1096), .b(G1192), .O(G1269) );
nand2 gate461( .a(G22), .b(G1195), .O(G1270) );
nand2 gate462( .a(G1099), .b(G1195), .O(G1271) );

  xor2  gate799(.a(G1198), .b(G23), .O(gate463inter0));
  nand2 gate800(.a(gate463inter0), .b(s_36), .O(gate463inter1));
  and2  gate801(.a(G1198), .b(G23), .O(gate463inter2));
  inv1  gate802(.a(s_36), .O(gate463inter3));
  inv1  gate803(.a(s_37), .O(gate463inter4));
  nand2 gate804(.a(gate463inter4), .b(gate463inter3), .O(gate463inter5));
  nor2  gate805(.a(gate463inter5), .b(gate463inter2), .O(gate463inter6));
  inv1  gate806(.a(G23), .O(gate463inter7));
  inv1  gate807(.a(G1198), .O(gate463inter8));
  nand2 gate808(.a(gate463inter8), .b(gate463inter7), .O(gate463inter9));
  nand2 gate809(.a(s_37), .b(gate463inter3), .O(gate463inter10));
  nor2  gate810(.a(gate463inter10), .b(gate463inter9), .O(gate463inter11));
  nor2  gate811(.a(gate463inter11), .b(gate463inter6), .O(gate463inter12));
  nand2 gate812(.a(gate463inter12), .b(gate463inter1), .O(G1272));
nand2 gate464( .a(G1102), .b(G1198), .O(G1273) );
nand2 gate465( .a(G24), .b(G1201), .O(G1274) );
nand2 gate466( .a(G1105), .b(G1201), .O(G1275) );
nand2 gate467( .a(G25), .b(G1204), .O(G1276) );
nand2 gate468( .a(G1108), .b(G1204), .O(G1277) );
nand2 gate469( .a(G26), .b(G1207), .O(G1278) );
nand2 gate470( .a(G1111), .b(G1207), .O(G1279) );

  xor2  gate729(.a(G1210), .b(G27), .O(gate471inter0));
  nand2 gate730(.a(gate471inter0), .b(s_26), .O(gate471inter1));
  and2  gate731(.a(G1210), .b(G27), .O(gate471inter2));
  inv1  gate732(.a(s_26), .O(gate471inter3));
  inv1  gate733(.a(s_27), .O(gate471inter4));
  nand2 gate734(.a(gate471inter4), .b(gate471inter3), .O(gate471inter5));
  nor2  gate735(.a(gate471inter5), .b(gate471inter2), .O(gate471inter6));
  inv1  gate736(.a(G27), .O(gate471inter7));
  inv1  gate737(.a(G1210), .O(gate471inter8));
  nand2 gate738(.a(gate471inter8), .b(gate471inter7), .O(gate471inter9));
  nand2 gate739(.a(s_27), .b(gate471inter3), .O(gate471inter10));
  nor2  gate740(.a(gate471inter10), .b(gate471inter9), .O(gate471inter11));
  nor2  gate741(.a(gate471inter11), .b(gate471inter6), .O(gate471inter12));
  nand2 gate742(.a(gate471inter12), .b(gate471inter1), .O(G1280));
nand2 gate472( .a(G1114), .b(G1210), .O(G1281) );
nand2 gate473( .a(G28), .b(G1213), .O(G1282) );
nand2 gate474( .a(G1117), .b(G1213), .O(G1283) );
nand2 gate475( .a(G29), .b(G1216), .O(G1284) );
nand2 gate476( .a(G1120), .b(G1216), .O(G1285) );
nand2 gate477( .a(G30), .b(G1219), .O(G1286) );
nand2 gate478( .a(G1123), .b(G1219), .O(G1287) );
nand2 gate479( .a(G31), .b(G1222), .O(G1288) );
nand2 gate480( .a(G1126), .b(G1222), .O(G1289) );
nand2 gate481( .a(G32), .b(G1225), .O(G1290) );
nand2 gate482( .a(G1129), .b(G1225), .O(G1291) );
nand2 gate483( .a(G1228), .b(G1229), .O(G1292) );
nand2 gate484( .a(G1230), .b(G1231), .O(G1293) );

  xor2  gate659(.a(G1233), .b(G1232), .O(gate485inter0));
  nand2 gate660(.a(gate485inter0), .b(s_16), .O(gate485inter1));
  and2  gate661(.a(G1233), .b(G1232), .O(gate485inter2));
  inv1  gate662(.a(s_16), .O(gate485inter3));
  inv1  gate663(.a(s_17), .O(gate485inter4));
  nand2 gate664(.a(gate485inter4), .b(gate485inter3), .O(gate485inter5));
  nor2  gate665(.a(gate485inter5), .b(gate485inter2), .O(gate485inter6));
  inv1  gate666(.a(G1232), .O(gate485inter7));
  inv1  gate667(.a(G1233), .O(gate485inter8));
  nand2 gate668(.a(gate485inter8), .b(gate485inter7), .O(gate485inter9));
  nand2 gate669(.a(s_17), .b(gate485inter3), .O(gate485inter10));
  nor2  gate670(.a(gate485inter10), .b(gate485inter9), .O(gate485inter11));
  nor2  gate671(.a(gate485inter11), .b(gate485inter6), .O(gate485inter12));
  nand2 gate672(.a(gate485inter12), .b(gate485inter1), .O(G1294));

  xor2  gate743(.a(G1235), .b(G1234), .O(gate486inter0));
  nand2 gate744(.a(gate486inter0), .b(s_28), .O(gate486inter1));
  and2  gate745(.a(G1235), .b(G1234), .O(gate486inter2));
  inv1  gate746(.a(s_28), .O(gate486inter3));
  inv1  gate747(.a(s_29), .O(gate486inter4));
  nand2 gate748(.a(gate486inter4), .b(gate486inter3), .O(gate486inter5));
  nor2  gate749(.a(gate486inter5), .b(gate486inter2), .O(gate486inter6));
  inv1  gate750(.a(G1234), .O(gate486inter7));
  inv1  gate751(.a(G1235), .O(gate486inter8));
  nand2 gate752(.a(gate486inter8), .b(gate486inter7), .O(gate486inter9));
  nand2 gate753(.a(s_29), .b(gate486inter3), .O(gate486inter10));
  nor2  gate754(.a(gate486inter10), .b(gate486inter9), .O(gate486inter11));
  nor2  gate755(.a(gate486inter11), .b(gate486inter6), .O(gate486inter12));
  nand2 gate756(.a(gate486inter12), .b(gate486inter1), .O(G1295));
nand2 gate487( .a(G1236), .b(G1237), .O(G1296) );
nand2 gate488( .a(G1238), .b(G1239), .O(G1297) );
nand2 gate489( .a(G1240), .b(G1241), .O(G1298) );
nand2 gate490( .a(G1242), .b(G1243), .O(G1299) );
nand2 gate491( .a(G1244), .b(G1245), .O(G1300) );
nand2 gate492( .a(G1246), .b(G1247), .O(G1301) );
nand2 gate493( .a(G1248), .b(G1249), .O(G1302) );

  xor2  gate855(.a(G1251), .b(G1250), .O(gate494inter0));
  nand2 gate856(.a(gate494inter0), .b(s_44), .O(gate494inter1));
  and2  gate857(.a(G1251), .b(G1250), .O(gate494inter2));
  inv1  gate858(.a(s_44), .O(gate494inter3));
  inv1  gate859(.a(s_45), .O(gate494inter4));
  nand2 gate860(.a(gate494inter4), .b(gate494inter3), .O(gate494inter5));
  nor2  gate861(.a(gate494inter5), .b(gate494inter2), .O(gate494inter6));
  inv1  gate862(.a(G1250), .O(gate494inter7));
  inv1  gate863(.a(G1251), .O(gate494inter8));
  nand2 gate864(.a(gate494inter8), .b(gate494inter7), .O(gate494inter9));
  nand2 gate865(.a(s_45), .b(gate494inter3), .O(gate494inter10));
  nor2  gate866(.a(gate494inter10), .b(gate494inter9), .O(gate494inter11));
  nor2  gate867(.a(gate494inter11), .b(gate494inter6), .O(gate494inter12));
  nand2 gate868(.a(gate494inter12), .b(gate494inter1), .O(G1303));
nand2 gate495( .a(G1252), .b(G1253), .O(G1304) );
nand2 gate496( .a(G1254), .b(G1255), .O(G1305) );
nand2 gate497( .a(G1256), .b(G1257), .O(G1306) );
nand2 gate498( .a(G1258), .b(G1259), .O(G1307) );
nand2 gate499( .a(G1260), .b(G1261), .O(G1308) );
nand2 gate500( .a(G1262), .b(G1263), .O(G1309) );
nand2 gate501( .a(G1264), .b(G1265), .O(G1310) );
nand2 gate502( .a(G1266), .b(G1267), .O(G1311) );

  xor2  gate785(.a(G1269), .b(G1268), .O(gate503inter0));
  nand2 gate786(.a(gate503inter0), .b(s_34), .O(gate503inter1));
  and2  gate787(.a(G1269), .b(G1268), .O(gate503inter2));
  inv1  gate788(.a(s_34), .O(gate503inter3));
  inv1  gate789(.a(s_35), .O(gate503inter4));
  nand2 gate790(.a(gate503inter4), .b(gate503inter3), .O(gate503inter5));
  nor2  gate791(.a(gate503inter5), .b(gate503inter2), .O(gate503inter6));
  inv1  gate792(.a(G1268), .O(gate503inter7));
  inv1  gate793(.a(G1269), .O(gate503inter8));
  nand2 gate794(.a(gate503inter8), .b(gate503inter7), .O(gate503inter9));
  nand2 gate795(.a(s_35), .b(gate503inter3), .O(gate503inter10));
  nor2  gate796(.a(gate503inter10), .b(gate503inter9), .O(gate503inter11));
  nor2  gate797(.a(gate503inter11), .b(gate503inter6), .O(gate503inter12));
  nand2 gate798(.a(gate503inter12), .b(gate503inter1), .O(G1312));
nand2 gate504( .a(G1270), .b(G1271), .O(G1313) );
nand2 gate505( .a(G1272), .b(G1273), .O(G1314) );
nand2 gate506( .a(G1274), .b(G1275), .O(G1315) );
nand2 gate507( .a(G1276), .b(G1277), .O(G1316) );
nand2 gate508( .a(G1278), .b(G1279), .O(G1317) );
nand2 gate509( .a(G1280), .b(G1281), .O(G1318) );

  xor2  gate1079(.a(G1283), .b(G1282), .O(gate510inter0));
  nand2 gate1080(.a(gate510inter0), .b(s_76), .O(gate510inter1));
  and2  gate1081(.a(G1283), .b(G1282), .O(gate510inter2));
  inv1  gate1082(.a(s_76), .O(gate510inter3));
  inv1  gate1083(.a(s_77), .O(gate510inter4));
  nand2 gate1084(.a(gate510inter4), .b(gate510inter3), .O(gate510inter5));
  nor2  gate1085(.a(gate510inter5), .b(gate510inter2), .O(gate510inter6));
  inv1  gate1086(.a(G1282), .O(gate510inter7));
  inv1  gate1087(.a(G1283), .O(gate510inter8));
  nand2 gate1088(.a(gate510inter8), .b(gate510inter7), .O(gate510inter9));
  nand2 gate1089(.a(s_77), .b(gate510inter3), .O(gate510inter10));
  nor2  gate1090(.a(gate510inter10), .b(gate510inter9), .O(gate510inter11));
  nor2  gate1091(.a(gate510inter11), .b(gate510inter6), .O(gate510inter12));
  nand2 gate1092(.a(gate510inter12), .b(gate510inter1), .O(G1319));
nand2 gate511( .a(G1284), .b(G1285), .O(G1320) );
nand2 gate512( .a(G1286), .b(G1287), .O(G1321) );
nand2 gate513( .a(G1288), .b(G1289), .O(G1322) );
nand2 gate514( .a(G1290), .b(G1291), .O(G1323) );
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule