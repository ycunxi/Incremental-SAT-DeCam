module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);

input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;//RE__PI;

input s_0,s_1;//RE__ALLOW(00,01,10,11);
input s_2,s_3;//RE__ALLOW(00,01,10,11);
input s_4,s_5;//RE__ALLOW(00,01,10,11);
input s_6,s_7;//RE__ALLOW(00,01,10,11);
input s_8,s_9;//RE__ALLOW(00,01,10,11);
input s_10,s_11;//RE__ALLOW(00,01,10,11);
input s_12,s_13;//RE__ALLOW(00,01,10,11);
input s_14,s_15;//RE__ALLOW(00,01,10,11);
input s_16,s_17;//RE__ALLOW(00,01,10,11);
input s_18,s_19;//RE__ALLOW(00,01,10,11);
input s_20,s_21;//RE__ALLOW(00,01,10,11);
input s_22,s_23;//RE__ALLOW(00,01,10,11);
input s_24,s_25;//RE__ALLOW(00,01,10,11);
input s_26,s_27;//RE__ALLOW(00,01,10,11);
input s_28,s_29;//RE__ALLOW(00,01,10,11);
input s_30,s_31;//RE__ALLOW(00,01,10,11);
input s_32,s_33;//RE__ALLOW(00,01,10,11);
input s_34,s_35;//RE__ALLOW(00,01,10,11);
input s_36,s_37;//RE__ALLOW(00,01,10,11);
input s_38,s_39;//RE__ALLOW(00,01,10,11);
input s_40,s_41;//RE__ALLOW(00,01,10,11);
input s_42,s_43;//RE__ALLOW(00,01,10,11);
input s_44,s_45;//RE__ALLOW(00,01,10,11);
input s_46,s_47;//RE__ALLOW(00,01,10,11);
input s_48,s_49;//RE__ALLOW(00,01,10,11);
input s_50,s_51;//RE__ALLOW(00,01,10,11);
input s_52,s_53;//RE__ALLOW(00,01,10,11);
input s_54,s_55;//RE__ALLOW(00,01,10,11);
input s_56,s_57;//RE__ALLOW(00,01,10,11);
input s_58,s_59;//RE__ALLOW(00,01,10,11);
input s_60,s_61;//RE__ALLOW(00,01,10,11);
input s_62,s_63;//RE__ALLOW(00,01,10,11);
input s_64,s_65;//RE__ALLOW(00,01,10,11);
input s_66,s_67;//RE__ALLOW(00,01,10,11);
input s_68,s_69;//RE__ALLOW(00,01,10,11);
input s_70,s_71;//RE__ALLOW(00,01,10,11);
input s_72,s_73;//RE__ALLOW(00,01,10,11);
input s_74,s_75;//RE__ALLOW(00,01,10,11);
input s_76,s_77;//RE__ALLOW(00,01,10,11);
input s_78,s_79;//RE__ALLOW(00,01,10,11);
input s_80,s_81;//RE__ALLOW(00,01,10,11);
input s_82,s_83;//RE__ALLOW(00,01,10,11);
input s_84,s_85;//RE__ALLOW(00,01,10,11);
input s_86,s_87;//RE__ALLOW(00,01,10,11);
input s_88,s_89;//RE__ALLOW(00,01,10,11);
input s_90,s_91;//RE__ALLOW(00,01,10,11);
input s_92,s_93;//RE__ALLOW(00,01,10,11);
input s_94,s_95;//RE__ALLOW(00,01,10,11);
input s_96,s_97;//RE__ALLOW(00,01,10,11);
input s_98,s_99;//RE__ALLOW(00,01,10,11);
input s_100,s_101;//RE__ALLOW(00,01,10,11);
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;

  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate198inter0, gate198inter1, gate198inter2, gate198inter3, gate198inter4, gate198inter5, gate198inter6, gate198inter7, gate198inter8, gate198inter9, gate198inter10, gate198inter11, gate198inter12, gate463inter0, gate463inter1, gate463inter2, gate463inter3, gate463inter4, gate463inter5, gate463inter6, gate463inter7, gate463inter8, gate463inter9, gate463inter10, gate463inter11, gate463inter12, gate398inter0, gate398inter1, gate398inter2, gate398inter3, gate398inter4, gate398inter5, gate398inter6, gate398inter7, gate398inter8, gate398inter9, gate398inter10, gate398inter11, gate398inter12, gate53inter0, gate53inter1, gate53inter2, gate53inter3, gate53inter4, gate53inter5, gate53inter6, gate53inter7, gate53inter8, gate53inter9, gate53inter10, gate53inter11, gate53inter12, gate407inter0, gate407inter1, gate407inter2, gate407inter3, gate407inter4, gate407inter5, gate407inter6, gate407inter7, gate407inter8, gate407inter9, gate407inter10, gate407inter11, gate407inter12, gate21inter0, gate21inter1, gate21inter2, gate21inter3, gate21inter4, gate21inter5, gate21inter6, gate21inter7, gate21inter8, gate21inter9, gate21inter10, gate21inter11, gate21inter12, gate137inter0, gate137inter1, gate137inter2, gate137inter3, gate137inter4, gate137inter5, gate137inter6, gate137inter7, gate137inter8, gate137inter9, gate137inter10, gate137inter11, gate137inter12, gate278inter0, gate278inter1, gate278inter2, gate278inter3, gate278inter4, gate278inter5, gate278inter6, gate278inter7, gate278inter8, gate278inter9, gate278inter10, gate278inter11, gate278inter12, gate449inter0, gate449inter1, gate449inter2, gate449inter3, gate449inter4, gate449inter5, gate449inter6, gate449inter7, gate449inter8, gate449inter9, gate449inter10, gate449inter11, gate449inter12, gate109inter0, gate109inter1, gate109inter2, gate109inter3, gate109inter4, gate109inter5, gate109inter6, gate109inter7, gate109inter8, gate109inter9, gate109inter10, gate109inter11, gate109inter12, gate258inter0, gate258inter1, gate258inter2, gate258inter3, gate258inter4, gate258inter5, gate258inter6, gate258inter7, gate258inter8, gate258inter9, gate258inter10, gate258inter11, gate258inter12, gate205inter0, gate205inter1, gate205inter2, gate205inter3, gate205inter4, gate205inter5, gate205inter6, gate205inter7, gate205inter8, gate205inter9, gate205inter10, gate205inter11, gate205inter12, gate86inter0, gate86inter1, gate86inter2, gate86inter3, gate86inter4, gate86inter5, gate86inter6, gate86inter7, gate86inter8, gate86inter9, gate86inter10, gate86inter11, gate86inter12, gate132inter0, gate132inter1, gate132inter2, gate132inter3, gate132inter4, gate132inter5, gate132inter6, gate132inter7, gate132inter8, gate132inter9, gate132inter10, gate132inter11, gate132inter12, gate421inter0, gate421inter1, gate421inter2, gate421inter3, gate421inter4, gate421inter5, gate421inter6, gate421inter7, gate421inter8, gate421inter9, gate421inter10, gate421inter11, gate421inter12, gate36inter0, gate36inter1, gate36inter2, gate36inter3, gate36inter4, gate36inter5, gate36inter6, gate36inter7, gate36inter8, gate36inter9, gate36inter10, gate36inter11, gate36inter12, gate152inter0, gate152inter1, gate152inter2, gate152inter3, gate152inter4, gate152inter5, gate152inter6, gate152inter7, gate152inter8, gate152inter9, gate152inter10, gate152inter11, gate152inter12, gate247inter0, gate247inter1, gate247inter2, gate247inter3, gate247inter4, gate247inter5, gate247inter6, gate247inter7, gate247inter8, gate247inter9, gate247inter10, gate247inter11, gate247inter12, gate438inter0, gate438inter1, gate438inter2, gate438inter3, gate438inter4, gate438inter5, gate438inter6, gate438inter7, gate438inter8, gate438inter9, gate438inter10, gate438inter11, gate438inter12, gate236inter0, gate236inter1, gate236inter2, gate236inter3, gate236inter4, gate236inter5, gate236inter6, gate236inter7, gate236inter8, gate236inter9, gate236inter10, gate236inter11, gate236inter12, gate501inter0, gate501inter1, gate501inter2, gate501inter3, gate501inter4, gate501inter5, gate501inter6, gate501inter7, gate501inter8, gate501inter9, gate501inter10, gate501inter11, gate501inter12, gate171inter0, gate171inter1, gate171inter2, gate171inter3, gate171inter4, gate171inter5, gate171inter6, gate171inter7, gate171inter8, gate171inter9, gate171inter10, gate171inter11, gate171inter12, gate18inter0, gate18inter1, gate18inter2, gate18inter3, gate18inter4, gate18inter5, gate18inter6, gate18inter7, gate18inter8, gate18inter9, gate18inter10, gate18inter11, gate18inter12, gate125inter0, gate125inter1, gate125inter2, gate125inter3, gate125inter4, gate125inter5, gate125inter6, gate125inter7, gate125inter8, gate125inter9, gate125inter10, gate125inter11, gate125inter12, gate142inter0, gate142inter1, gate142inter2, gate142inter3, gate142inter4, gate142inter5, gate142inter6, gate142inter7, gate142inter8, gate142inter9, gate142inter10, gate142inter11, gate142inter12, gate70inter0, gate70inter1, gate70inter2, gate70inter3, gate70inter4, gate70inter5, gate70inter6, gate70inter7, gate70inter8, gate70inter9, gate70inter10, gate70inter11, gate70inter12, gate255inter0, gate255inter1, gate255inter2, gate255inter3, gate255inter4, gate255inter5, gate255inter6, gate255inter7, gate255inter8, gate255inter9, gate255inter10, gate255inter11, gate255inter12, gate146inter0, gate146inter1, gate146inter2, gate146inter3, gate146inter4, gate146inter5, gate146inter6, gate146inter7, gate146inter8, gate146inter9, gate146inter10, gate146inter11, gate146inter12, gate424inter0, gate424inter1, gate424inter2, gate424inter3, gate424inter4, gate424inter5, gate424inter6, gate424inter7, gate424inter8, gate424inter9, gate424inter10, gate424inter11, gate424inter12, gate461inter0, gate461inter1, gate461inter2, gate461inter3, gate461inter4, gate461inter5, gate461inter6, gate461inter7, gate461inter8, gate461inter9, gate461inter10, gate461inter11, gate461inter12, gate47inter0, gate47inter1, gate47inter2, gate47inter3, gate47inter4, gate47inter5, gate47inter6, gate47inter7, gate47inter8, gate47inter9, gate47inter10, gate47inter11, gate47inter12, gate245inter0, gate245inter1, gate245inter2, gate245inter3, gate245inter4, gate245inter5, gate245inter6, gate245inter7, gate245inter8, gate245inter9, gate245inter10, gate245inter11, gate245inter12, gate294inter0, gate294inter1, gate294inter2, gate294inter3, gate294inter4, gate294inter5, gate294inter6, gate294inter7, gate294inter8, gate294inter9, gate294inter10, gate294inter11, gate294inter12, gate32inter0, gate32inter1, gate32inter2, gate32inter3, gate32inter4, gate32inter5, gate32inter6, gate32inter7, gate32inter8, gate32inter9, gate32inter10, gate32inter11, gate32inter12, gate181inter0, gate181inter1, gate181inter2, gate181inter3, gate181inter4, gate181inter5, gate181inter6, gate181inter7, gate181inter8, gate181inter9, gate181inter10, gate181inter11, gate181inter12, gate148inter0, gate148inter1, gate148inter2, gate148inter3, gate148inter4, gate148inter5, gate148inter6, gate148inter7, gate148inter8, gate148inter9, gate148inter10, gate148inter11, gate148inter12, gate504inter0, gate504inter1, gate504inter2, gate504inter3, gate504inter4, gate504inter5, gate504inter6, gate504inter7, gate504inter8, gate504inter9, gate504inter10, gate504inter11, gate504inter12, gate131inter0, gate131inter1, gate131inter2, gate131inter3, gate131inter4, gate131inter5, gate131inter6, gate131inter7, gate131inter8, gate131inter9, gate131inter10, gate131inter11, gate131inter12, gate200inter0, gate200inter1, gate200inter2, gate200inter3, gate200inter4, gate200inter5, gate200inter6, gate200inter7, gate200inter8, gate200inter9, gate200inter10, gate200inter11, gate200inter12, gate31inter0, gate31inter1, gate31inter2, gate31inter3, gate31inter4, gate31inter5, gate31inter6, gate31inter7, gate31inter8, gate31inter9, gate31inter10, gate31inter11, gate31inter12, gate456inter0, gate456inter1, gate456inter2, gate456inter3, gate456inter4, gate456inter5, gate456inter6, gate456inter7, gate456inter8, gate456inter9, gate456inter10, gate456inter11, gate456inter12, gate257inter0, gate257inter1, gate257inter2, gate257inter3, gate257inter4, gate257inter5, gate257inter6, gate257inter7, gate257inter8, gate257inter9, gate257inter10, gate257inter11, gate257inter12, gate503inter0, gate503inter1, gate503inter2, gate503inter3, gate503inter4, gate503inter5, gate503inter6, gate503inter7, gate503inter8, gate503inter9, gate503inter10, gate503inter11, gate503inter12, gate50inter0, gate50inter1, gate50inter2, gate50inter3, gate50inter4, gate50inter5, gate50inter6, gate50inter7, gate50inter8, gate50inter9, gate50inter10, gate50inter11, gate50inter12, gate473inter0, gate473inter1, gate473inter2, gate473inter3, gate473inter4, gate473inter5, gate473inter6, gate473inter7, gate473inter8, gate473inter9, gate473inter10, gate473inter11, gate473inter12, gate296inter0, gate296inter1, gate296inter2, gate296inter3, gate296inter4, gate296inter5, gate296inter6, gate296inter7, gate296inter8, gate296inter9, gate296inter10, gate296inter11, gate296inter12, gate87inter0, gate87inter1, gate87inter2, gate87inter3, gate87inter4, gate87inter5, gate87inter6, gate87inter7, gate87inter8, gate87inter9, gate87inter10, gate87inter11, gate87inter12, gate62inter0, gate62inter1, gate62inter2, gate62inter3, gate62inter4, gate62inter5, gate62inter6, gate62inter7, gate62inter8, gate62inter9, gate62inter10, gate62inter11, gate62inter12, gate42inter0, gate42inter1, gate42inter2, gate42inter3, gate42inter4, gate42inter5, gate42inter6, gate42inter7, gate42inter8, gate42inter9, gate42inter10, gate42inter11, gate42inter12, gate208inter0, gate208inter1, gate208inter2, gate208inter3, gate208inter4, gate208inter5, gate208inter6, gate208inter7, gate208inter8, gate208inter9, gate208inter10, gate208inter11, gate208inter12, gate510inter0, gate510inter1, gate510inter2, gate510inter3, gate510inter4, gate510inter5, gate510inter6, gate510inter7, gate510inter8, gate510inter9, gate510inter10, gate510inter11, gate510inter12;



and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );
nand2 gate9( .a(G1), .b(G2), .O(G266) );
nand2 gate10( .a(G3), .b(G4), .O(G269) );
nand2 gate11( .a(G5), .b(G6), .O(G272) );
nand2 gate12( .a(G7), .b(G8), .O(G275) );
nand2 gate13( .a(G9), .b(G10), .O(G278) );
nand2 gate14( .a(G11), .b(G12), .O(G281) );
nand2 gate15( .a(G13), .b(G14), .O(G284) );
nand2 gate16( .a(G15), .b(G16), .O(G287) );
nand2 gate17( .a(G17), .b(G18), .O(G290) );

  xor2  gate855(.a(G20), .b(G19), .O(gate18inter0));
  nand2 gate856(.a(gate18inter0), .b(s_44), .O(gate18inter1));
  and2  gate857(.a(G20), .b(G19), .O(gate18inter2));
  inv1  gate858(.a(s_44), .O(gate18inter3));
  inv1  gate859(.a(s_45), .O(gate18inter4));
  nand2 gate860(.a(gate18inter4), .b(gate18inter3), .O(gate18inter5));
  nor2  gate861(.a(gate18inter5), .b(gate18inter2), .O(gate18inter6));
  inv1  gate862(.a(G19), .O(gate18inter7));
  inv1  gate863(.a(G20), .O(gate18inter8));
  nand2 gate864(.a(gate18inter8), .b(gate18inter7), .O(gate18inter9));
  nand2 gate865(.a(s_45), .b(gate18inter3), .O(gate18inter10));
  nor2  gate866(.a(gate18inter10), .b(gate18inter9), .O(gate18inter11));
  nor2  gate867(.a(gate18inter11), .b(gate18inter6), .O(gate18inter12));
  nand2 gate868(.a(gate18inter12), .b(gate18inter1), .O(G293));
nand2 gate19( .a(G21), .b(G22), .O(G296) );
nand2 gate20( .a(G23), .b(G24), .O(G299) );

  xor2  gate617(.a(G26), .b(G25), .O(gate21inter0));
  nand2 gate618(.a(gate21inter0), .b(s_10), .O(gate21inter1));
  and2  gate619(.a(G26), .b(G25), .O(gate21inter2));
  inv1  gate620(.a(s_10), .O(gate21inter3));
  inv1  gate621(.a(s_11), .O(gate21inter4));
  nand2 gate622(.a(gate21inter4), .b(gate21inter3), .O(gate21inter5));
  nor2  gate623(.a(gate21inter5), .b(gate21inter2), .O(gate21inter6));
  inv1  gate624(.a(G25), .O(gate21inter7));
  inv1  gate625(.a(G26), .O(gate21inter8));
  nand2 gate626(.a(gate21inter8), .b(gate21inter7), .O(gate21inter9));
  nand2 gate627(.a(s_11), .b(gate21inter3), .O(gate21inter10));
  nor2  gate628(.a(gate21inter10), .b(gate21inter9), .O(gate21inter11));
  nor2  gate629(.a(gate21inter11), .b(gate21inter6), .O(gate21inter12));
  nand2 gate630(.a(gate21inter12), .b(gate21inter1), .O(G302));
nand2 gate22( .a(G27), .b(G28), .O(G305) );
nand2 gate23( .a(G29), .b(G30), .O(G308) );
nand2 gate24( .a(G31), .b(G32), .O(G311) );
nand2 gate25( .a(G1), .b(G5), .O(G314) );
nand2 gate26( .a(G9), .b(G13), .O(G317) );
nand2 gate27( .a(G2), .b(G6), .O(G320) );
nand2 gate28( .a(G10), .b(G14), .O(G323) );
nand2 gate29( .a(G3), .b(G7), .O(G326) );
nand2 gate30( .a(G11), .b(G15), .O(G329) );

  xor2  gate1093(.a(G8), .b(G4), .O(gate31inter0));
  nand2 gate1094(.a(gate31inter0), .b(s_78), .O(gate31inter1));
  and2  gate1095(.a(G8), .b(G4), .O(gate31inter2));
  inv1  gate1096(.a(s_78), .O(gate31inter3));
  inv1  gate1097(.a(s_79), .O(gate31inter4));
  nand2 gate1098(.a(gate31inter4), .b(gate31inter3), .O(gate31inter5));
  nor2  gate1099(.a(gate31inter5), .b(gate31inter2), .O(gate31inter6));
  inv1  gate1100(.a(G4), .O(gate31inter7));
  inv1  gate1101(.a(G8), .O(gate31inter8));
  nand2 gate1102(.a(gate31inter8), .b(gate31inter7), .O(gate31inter9));
  nand2 gate1103(.a(s_79), .b(gate31inter3), .O(gate31inter10));
  nor2  gate1104(.a(gate31inter10), .b(gate31inter9), .O(gate31inter11));
  nor2  gate1105(.a(gate31inter11), .b(gate31inter6), .O(gate31inter12));
  nand2 gate1106(.a(gate31inter12), .b(gate31inter1), .O(G332));

  xor2  gate1009(.a(G16), .b(G12), .O(gate32inter0));
  nand2 gate1010(.a(gate32inter0), .b(s_66), .O(gate32inter1));
  and2  gate1011(.a(G16), .b(G12), .O(gate32inter2));
  inv1  gate1012(.a(s_66), .O(gate32inter3));
  inv1  gate1013(.a(s_67), .O(gate32inter4));
  nand2 gate1014(.a(gate32inter4), .b(gate32inter3), .O(gate32inter5));
  nor2  gate1015(.a(gate32inter5), .b(gate32inter2), .O(gate32inter6));
  inv1  gate1016(.a(G12), .O(gate32inter7));
  inv1  gate1017(.a(G16), .O(gate32inter8));
  nand2 gate1018(.a(gate32inter8), .b(gate32inter7), .O(gate32inter9));
  nand2 gate1019(.a(s_67), .b(gate32inter3), .O(gate32inter10));
  nor2  gate1020(.a(gate32inter10), .b(gate32inter9), .O(gate32inter11));
  nor2  gate1021(.a(gate32inter11), .b(gate32inter6), .O(gate32inter12));
  nand2 gate1022(.a(gate32inter12), .b(gate32inter1), .O(G335));
nand2 gate33( .a(G17), .b(G21), .O(G338) );
nand2 gate34( .a(G25), .b(G29), .O(G341) );
nand2 gate35( .a(G18), .b(G22), .O(G344) );

  xor2  gate757(.a(G30), .b(G26), .O(gate36inter0));
  nand2 gate758(.a(gate36inter0), .b(s_30), .O(gate36inter1));
  and2  gate759(.a(G30), .b(G26), .O(gate36inter2));
  inv1  gate760(.a(s_30), .O(gate36inter3));
  inv1  gate761(.a(s_31), .O(gate36inter4));
  nand2 gate762(.a(gate36inter4), .b(gate36inter3), .O(gate36inter5));
  nor2  gate763(.a(gate36inter5), .b(gate36inter2), .O(gate36inter6));
  inv1  gate764(.a(G26), .O(gate36inter7));
  inv1  gate765(.a(G30), .O(gate36inter8));
  nand2 gate766(.a(gate36inter8), .b(gate36inter7), .O(gate36inter9));
  nand2 gate767(.a(s_31), .b(gate36inter3), .O(gate36inter10));
  nor2  gate768(.a(gate36inter10), .b(gate36inter9), .O(gate36inter11));
  nor2  gate769(.a(gate36inter11), .b(gate36inter6), .O(gate36inter12));
  nand2 gate770(.a(gate36inter12), .b(gate36inter1), .O(G347));
nand2 gate37( .a(G19), .b(G23), .O(G350) );
nand2 gate38( .a(G27), .b(G31), .O(G353) );
nand2 gate39( .a(G20), .b(G24), .O(G356) );
nand2 gate40( .a(G28), .b(G32), .O(G359) );
nand2 gate41( .a(G1), .b(G266), .O(G362) );

  xor2  gate1219(.a(G266), .b(G2), .O(gate42inter0));
  nand2 gate1220(.a(gate42inter0), .b(s_96), .O(gate42inter1));
  and2  gate1221(.a(G266), .b(G2), .O(gate42inter2));
  inv1  gate1222(.a(s_96), .O(gate42inter3));
  inv1  gate1223(.a(s_97), .O(gate42inter4));
  nand2 gate1224(.a(gate42inter4), .b(gate42inter3), .O(gate42inter5));
  nor2  gate1225(.a(gate42inter5), .b(gate42inter2), .O(gate42inter6));
  inv1  gate1226(.a(G2), .O(gate42inter7));
  inv1  gate1227(.a(G266), .O(gate42inter8));
  nand2 gate1228(.a(gate42inter8), .b(gate42inter7), .O(gate42inter9));
  nand2 gate1229(.a(s_97), .b(gate42inter3), .O(gate42inter10));
  nor2  gate1230(.a(gate42inter10), .b(gate42inter9), .O(gate42inter11));
  nor2  gate1231(.a(gate42inter11), .b(gate42inter6), .O(gate42inter12));
  nand2 gate1232(.a(gate42inter12), .b(gate42inter1), .O(G363));
nand2 gate43( .a(G3), .b(G269), .O(G364) );
nand2 gate44( .a(G4), .b(G269), .O(G365) );
nand2 gate45( .a(G5), .b(G272), .O(G366) );
nand2 gate46( .a(G6), .b(G272), .O(G367) );

  xor2  gate967(.a(G275), .b(G7), .O(gate47inter0));
  nand2 gate968(.a(gate47inter0), .b(s_60), .O(gate47inter1));
  and2  gate969(.a(G275), .b(G7), .O(gate47inter2));
  inv1  gate970(.a(s_60), .O(gate47inter3));
  inv1  gate971(.a(s_61), .O(gate47inter4));
  nand2 gate972(.a(gate47inter4), .b(gate47inter3), .O(gate47inter5));
  nor2  gate973(.a(gate47inter5), .b(gate47inter2), .O(gate47inter6));
  inv1  gate974(.a(G7), .O(gate47inter7));
  inv1  gate975(.a(G275), .O(gate47inter8));
  nand2 gate976(.a(gate47inter8), .b(gate47inter7), .O(gate47inter9));
  nand2 gate977(.a(s_61), .b(gate47inter3), .O(gate47inter10));
  nor2  gate978(.a(gate47inter10), .b(gate47inter9), .O(gate47inter11));
  nor2  gate979(.a(gate47inter11), .b(gate47inter6), .O(gate47inter12));
  nand2 gate980(.a(gate47inter12), .b(gate47inter1), .O(G368));
nand2 gate48( .a(G8), .b(G275), .O(G369) );
nand2 gate49( .a(G9), .b(G278), .O(G370) );

  xor2  gate1149(.a(G278), .b(G10), .O(gate50inter0));
  nand2 gate1150(.a(gate50inter0), .b(s_86), .O(gate50inter1));
  and2  gate1151(.a(G278), .b(G10), .O(gate50inter2));
  inv1  gate1152(.a(s_86), .O(gate50inter3));
  inv1  gate1153(.a(s_87), .O(gate50inter4));
  nand2 gate1154(.a(gate50inter4), .b(gate50inter3), .O(gate50inter5));
  nor2  gate1155(.a(gate50inter5), .b(gate50inter2), .O(gate50inter6));
  inv1  gate1156(.a(G10), .O(gate50inter7));
  inv1  gate1157(.a(G278), .O(gate50inter8));
  nand2 gate1158(.a(gate50inter8), .b(gate50inter7), .O(gate50inter9));
  nand2 gate1159(.a(s_87), .b(gate50inter3), .O(gate50inter10));
  nor2  gate1160(.a(gate50inter10), .b(gate50inter9), .O(gate50inter11));
  nor2  gate1161(.a(gate50inter11), .b(gate50inter6), .O(gate50inter12));
  nand2 gate1162(.a(gate50inter12), .b(gate50inter1), .O(G371));
nand2 gate51( .a(G11), .b(G281), .O(G372) );
nand2 gate52( .a(G12), .b(G281), .O(G373) );

  xor2  gate589(.a(G284), .b(G13), .O(gate53inter0));
  nand2 gate590(.a(gate53inter0), .b(s_6), .O(gate53inter1));
  and2  gate591(.a(G284), .b(G13), .O(gate53inter2));
  inv1  gate592(.a(s_6), .O(gate53inter3));
  inv1  gate593(.a(s_7), .O(gate53inter4));
  nand2 gate594(.a(gate53inter4), .b(gate53inter3), .O(gate53inter5));
  nor2  gate595(.a(gate53inter5), .b(gate53inter2), .O(gate53inter6));
  inv1  gate596(.a(G13), .O(gate53inter7));
  inv1  gate597(.a(G284), .O(gate53inter8));
  nand2 gate598(.a(gate53inter8), .b(gate53inter7), .O(gate53inter9));
  nand2 gate599(.a(s_7), .b(gate53inter3), .O(gate53inter10));
  nor2  gate600(.a(gate53inter10), .b(gate53inter9), .O(gate53inter11));
  nor2  gate601(.a(gate53inter11), .b(gate53inter6), .O(gate53inter12));
  nand2 gate602(.a(gate53inter12), .b(gate53inter1), .O(G374));
nand2 gate54( .a(G14), .b(G284), .O(G375) );
nand2 gate55( .a(G15), .b(G287), .O(G376) );
nand2 gate56( .a(G16), .b(G287), .O(G377) );
nand2 gate57( .a(G17), .b(G290), .O(G378) );
nand2 gate58( .a(G18), .b(G290), .O(G379) );
nand2 gate59( .a(G19), .b(G293), .O(G380) );
nand2 gate60( .a(G20), .b(G293), .O(G381) );
nand2 gate61( .a(G21), .b(G296), .O(G382) );

  xor2  gate1205(.a(G296), .b(G22), .O(gate62inter0));
  nand2 gate1206(.a(gate62inter0), .b(s_94), .O(gate62inter1));
  and2  gate1207(.a(G296), .b(G22), .O(gate62inter2));
  inv1  gate1208(.a(s_94), .O(gate62inter3));
  inv1  gate1209(.a(s_95), .O(gate62inter4));
  nand2 gate1210(.a(gate62inter4), .b(gate62inter3), .O(gate62inter5));
  nor2  gate1211(.a(gate62inter5), .b(gate62inter2), .O(gate62inter6));
  inv1  gate1212(.a(G22), .O(gate62inter7));
  inv1  gate1213(.a(G296), .O(gate62inter8));
  nand2 gate1214(.a(gate62inter8), .b(gate62inter7), .O(gate62inter9));
  nand2 gate1215(.a(s_95), .b(gate62inter3), .O(gate62inter10));
  nor2  gate1216(.a(gate62inter10), .b(gate62inter9), .O(gate62inter11));
  nor2  gate1217(.a(gate62inter11), .b(gate62inter6), .O(gate62inter12));
  nand2 gate1218(.a(gate62inter12), .b(gate62inter1), .O(G383));
nand2 gate63( .a(G23), .b(G299), .O(G384) );
nand2 gate64( .a(G24), .b(G299), .O(G385) );
nand2 gate65( .a(G25), .b(G302), .O(G386) );
nand2 gate66( .a(G26), .b(G302), .O(G387) );
nand2 gate67( .a(G27), .b(G305), .O(G388) );
nand2 gate68( .a(G28), .b(G305), .O(G389) );
nand2 gate69( .a(G29), .b(G308), .O(G390) );

  xor2  gate897(.a(G308), .b(G30), .O(gate70inter0));
  nand2 gate898(.a(gate70inter0), .b(s_50), .O(gate70inter1));
  and2  gate899(.a(G308), .b(G30), .O(gate70inter2));
  inv1  gate900(.a(s_50), .O(gate70inter3));
  inv1  gate901(.a(s_51), .O(gate70inter4));
  nand2 gate902(.a(gate70inter4), .b(gate70inter3), .O(gate70inter5));
  nor2  gate903(.a(gate70inter5), .b(gate70inter2), .O(gate70inter6));
  inv1  gate904(.a(G30), .O(gate70inter7));
  inv1  gate905(.a(G308), .O(gate70inter8));
  nand2 gate906(.a(gate70inter8), .b(gate70inter7), .O(gate70inter9));
  nand2 gate907(.a(s_51), .b(gate70inter3), .O(gate70inter10));
  nor2  gate908(.a(gate70inter10), .b(gate70inter9), .O(gate70inter11));
  nor2  gate909(.a(gate70inter11), .b(gate70inter6), .O(gate70inter12));
  nand2 gate910(.a(gate70inter12), .b(gate70inter1), .O(G391));
nand2 gate71( .a(G31), .b(G311), .O(G392) );
nand2 gate72( .a(G32), .b(G311), .O(G393) );
nand2 gate73( .a(G1), .b(G314), .O(G394) );
nand2 gate74( .a(G5), .b(G314), .O(G395) );
nand2 gate75( .a(G9), .b(G317), .O(G396) );
nand2 gate76( .a(G13), .b(G317), .O(G397) );
nand2 gate77( .a(G2), .b(G320), .O(G398) );
nand2 gate78( .a(G6), .b(G320), .O(G399) );
nand2 gate79( .a(G10), .b(G323), .O(G400) );
nand2 gate80( .a(G14), .b(G323), .O(G401) );
nand2 gate81( .a(G3), .b(G326), .O(G402) );
nand2 gate82( .a(G7), .b(G326), .O(G403) );
nand2 gate83( .a(G11), .b(G329), .O(G404) );
nand2 gate84( .a(G15), .b(G329), .O(G405) );
nand2 gate85( .a(G4), .b(G332), .O(G406) );

  xor2  gate715(.a(G332), .b(G8), .O(gate86inter0));
  nand2 gate716(.a(gate86inter0), .b(s_24), .O(gate86inter1));
  and2  gate717(.a(G332), .b(G8), .O(gate86inter2));
  inv1  gate718(.a(s_24), .O(gate86inter3));
  inv1  gate719(.a(s_25), .O(gate86inter4));
  nand2 gate720(.a(gate86inter4), .b(gate86inter3), .O(gate86inter5));
  nor2  gate721(.a(gate86inter5), .b(gate86inter2), .O(gate86inter6));
  inv1  gate722(.a(G8), .O(gate86inter7));
  inv1  gate723(.a(G332), .O(gate86inter8));
  nand2 gate724(.a(gate86inter8), .b(gate86inter7), .O(gate86inter9));
  nand2 gate725(.a(s_25), .b(gate86inter3), .O(gate86inter10));
  nor2  gate726(.a(gate86inter10), .b(gate86inter9), .O(gate86inter11));
  nor2  gate727(.a(gate86inter11), .b(gate86inter6), .O(gate86inter12));
  nand2 gate728(.a(gate86inter12), .b(gate86inter1), .O(G407));

  xor2  gate1191(.a(G335), .b(G12), .O(gate87inter0));
  nand2 gate1192(.a(gate87inter0), .b(s_92), .O(gate87inter1));
  and2  gate1193(.a(G335), .b(G12), .O(gate87inter2));
  inv1  gate1194(.a(s_92), .O(gate87inter3));
  inv1  gate1195(.a(s_93), .O(gate87inter4));
  nand2 gate1196(.a(gate87inter4), .b(gate87inter3), .O(gate87inter5));
  nor2  gate1197(.a(gate87inter5), .b(gate87inter2), .O(gate87inter6));
  inv1  gate1198(.a(G12), .O(gate87inter7));
  inv1  gate1199(.a(G335), .O(gate87inter8));
  nand2 gate1200(.a(gate87inter8), .b(gate87inter7), .O(gate87inter9));
  nand2 gate1201(.a(s_93), .b(gate87inter3), .O(gate87inter10));
  nor2  gate1202(.a(gate87inter10), .b(gate87inter9), .O(gate87inter11));
  nor2  gate1203(.a(gate87inter11), .b(gate87inter6), .O(gate87inter12));
  nand2 gate1204(.a(gate87inter12), .b(gate87inter1), .O(G408));
nand2 gate88( .a(G16), .b(G335), .O(G409) );
nand2 gate89( .a(G17), .b(G338), .O(G410) );
nand2 gate90( .a(G21), .b(G338), .O(G411) );
nand2 gate91( .a(G25), .b(G341), .O(G412) );
nand2 gate92( .a(G29), .b(G341), .O(G413) );
nand2 gate93( .a(G18), .b(G344), .O(G414) );
nand2 gate94( .a(G22), .b(G344), .O(G415) );
nand2 gate95( .a(G26), .b(G347), .O(G416) );
nand2 gate96( .a(G30), .b(G347), .O(G417) );
nand2 gate97( .a(G19), .b(G350), .O(G418) );
nand2 gate98( .a(G23), .b(G350), .O(G419) );
nand2 gate99( .a(G27), .b(G353), .O(G420) );
nand2 gate100( .a(G31), .b(G353), .O(G421) );
nand2 gate101( .a(G20), .b(G356), .O(G422) );
nand2 gate102( .a(G24), .b(G356), .O(G423) );
nand2 gate103( .a(G28), .b(G359), .O(G424) );
nand2 gate104( .a(G32), .b(G359), .O(G425) );
nand2 gate105( .a(G362), .b(G363), .O(G426) );
nand2 gate106( .a(G364), .b(G365), .O(G429) );
nand2 gate107( .a(G366), .b(G367), .O(G432) );
nand2 gate108( .a(G368), .b(G369), .O(G435) );

  xor2  gate673(.a(G371), .b(G370), .O(gate109inter0));
  nand2 gate674(.a(gate109inter0), .b(s_18), .O(gate109inter1));
  and2  gate675(.a(G371), .b(G370), .O(gate109inter2));
  inv1  gate676(.a(s_18), .O(gate109inter3));
  inv1  gate677(.a(s_19), .O(gate109inter4));
  nand2 gate678(.a(gate109inter4), .b(gate109inter3), .O(gate109inter5));
  nor2  gate679(.a(gate109inter5), .b(gate109inter2), .O(gate109inter6));
  inv1  gate680(.a(G370), .O(gate109inter7));
  inv1  gate681(.a(G371), .O(gate109inter8));
  nand2 gate682(.a(gate109inter8), .b(gate109inter7), .O(gate109inter9));
  nand2 gate683(.a(s_19), .b(gate109inter3), .O(gate109inter10));
  nor2  gate684(.a(gate109inter10), .b(gate109inter9), .O(gate109inter11));
  nor2  gate685(.a(gate109inter11), .b(gate109inter6), .O(gate109inter12));
  nand2 gate686(.a(gate109inter12), .b(gate109inter1), .O(G438));
nand2 gate110( .a(G372), .b(G373), .O(G441) );
nand2 gate111( .a(G374), .b(G375), .O(G444) );
nand2 gate112( .a(G376), .b(G377), .O(G447) );
nand2 gate113( .a(G378), .b(G379), .O(G450) );
nand2 gate114( .a(G380), .b(G381), .O(G453) );
nand2 gate115( .a(G382), .b(G383), .O(G456) );
nand2 gate116( .a(G384), .b(G385), .O(G459) );
nand2 gate117( .a(G386), .b(G387), .O(G462) );
nand2 gate118( .a(G388), .b(G389), .O(G465) );
nand2 gate119( .a(G390), .b(G391), .O(G468) );
nand2 gate120( .a(G392), .b(G393), .O(G471) );
nand2 gate121( .a(G394), .b(G395), .O(G474) );
nand2 gate122( .a(G396), .b(G397), .O(G477) );
nand2 gate123( .a(G398), .b(G399), .O(G480) );
nand2 gate124( .a(G400), .b(G401), .O(G483) );

  xor2  gate869(.a(G403), .b(G402), .O(gate125inter0));
  nand2 gate870(.a(gate125inter0), .b(s_46), .O(gate125inter1));
  and2  gate871(.a(G403), .b(G402), .O(gate125inter2));
  inv1  gate872(.a(s_46), .O(gate125inter3));
  inv1  gate873(.a(s_47), .O(gate125inter4));
  nand2 gate874(.a(gate125inter4), .b(gate125inter3), .O(gate125inter5));
  nor2  gate875(.a(gate125inter5), .b(gate125inter2), .O(gate125inter6));
  inv1  gate876(.a(G402), .O(gate125inter7));
  inv1  gate877(.a(G403), .O(gate125inter8));
  nand2 gate878(.a(gate125inter8), .b(gate125inter7), .O(gate125inter9));
  nand2 gate879(.a(s_47), .b(gate125inter3), .O(gate125inter10));
  nor2  gate880(.a(gate125inter10), .b(gate125inter9), .O(gate125inter11));
  nor2  gate881(.a(gate125inter11), .b(gate125inter6), .O(gate125inter12));
  nand2 gate882(.a(gate125inter12), .b(gate125inter1), .O(G486));
nand2 gate126( .a(G404), .b(G405), .O(G489) );
nand2 gate127( .a(G406), .b(G407), .O(G492) );
nand2 gate128( .a(G408), .b(G409), .O(G495) );
nand2 gate129( .a(G410), .b(G411), .O(G498) );
nand2 gate130( .a(G412), .b(G413), .O(G501) );

  xor2  gate1065(.a(G415), .b(G414), .O(gate131inter0));
  nand2 gate1066(.a(gate131inter0), .b(s_74), .O(gate131inter1));
  and2  gate1067(.a(G415), .b(G414), .O(gate131inter2));
  inv1  gate1068(.a(s_74), .O(gate131inter3));
  inv1  gate1069(.a(s_75), .O(gate131inter4));
  nand2 gate1070(.a(gate131inter4), .b(gate131inter3), .O(gate131inter5));
  nor2  gate1071(.a(gate131inter5), .b(gate131inter2), .O(gate131inter6));
  inv1  gate1072(.a(G414), .O(gate131inter7));
  inv1  gate1073(.a(G415), .O(gate131inter8));
  nand2 gate1074(.a(gate131inter8), .b(gate131inter7), .O(gate131inter9));
  nand2 gate1075(.a(s_75), .b(gate131inter3), .O(gate131inter10));
  nor2  gate1076(.a(gate131inter10), .b(gate131inter9), .O(gate131inter11));
  nor2  gate1077(.a(gate131inter11), .b(gate131inter6), .O(gate131inter12));
  nand2 gate1078(.a(gate131inter12), .b(gate131inter1), .O(G504));

  xor2  gate729(.a(G417), .b(G416), .O(gate132inter0));
  nand2 gate730(.a(gate132inter0), .b(s_26), .O(gate132inter1));
  and2  gate731(.a(G417), .b(G416), .O(gate132inter2));
  inv1  gate732(.a(s_26), .O(gate132inter3));
  inv1  gate733(.a(s_27), .O(gate132inter4));
  nand2 gate734(.a(gate132inter4), .b(gate132inter3), .O(gate132inter5));
  nor2  gate735(.a(gate132inter5), .b(gate132inter2), .O(gate132inter6));
  inv1  gate736(.a(G416), .O(gate132inter7));
  inv1  gate737(.a(G417), .O(gate132inter8));
  nand2 gate738(.a(gate132inter8), .b(gate132inter7), .O(gate132inter9));
  nand2 gate739(.a(s_27), .b(gate132inter3), .O(gate132inter10));
  nor2  gate740(.a(gate132inter10), .b(gate132inter9), .O(gate132inter11));
  nor2  gate741(.a(gate132inter11), .b(gate132inter6), .O(gate132inter12));
  nand2 gate742(.a(gate132inter12), .b(gate132inter1), .O(G507));
nand2 gate133( .a(G418), .b(G419), .O(G510) );
nand2 gate134( .a(G420), .b(G421), .O(G513) );
nand2 gate135( .a(G422), .b(G423), .O(G516) );
nand2 gate136( .a(G424), .b(G425), .O(G519) );

  xor2  gate631(.a(G429), .b(G426), .O(gate137inter0));
  nand2 gate632(.a(gate137inter0), .b(s_12), .O(gate137inter1));
  and2  gate633(.a(G429), .b(G426), .O(gate137inter2));
  inv1  gate634(.a(s_12), .O(gate137inter3));
  inv1  gate635(.a(s_13), .O(gate137inter4));
  nand2 gate636(.a(gate137inter4), .b(gate137inter3), .O(gate137inter5));
  nor2  gate637(.a(gate137inter5), .b(gate137inter2), .O(gate137inter6));
  inv1  gate638(.a(G426), .O(gate137inter7));
  inv1  gate639(.a(G429), .O(gate137inter8));
  nand2 gate640(.a(gate137inter8), .b(gate137inter7), .O(gate137inter9));
  nand2 gate641(.a(s_13), .b(gate137inter3), .O(gate137inter10));
  nor2  gate642(.a(gate137inter10), .b(gate137inter9), .O(gate137inter11));
  nor2  gate643(.a(gate137inter11), .b(gate137inter6), .O(gate137inter12));
  nand2 gate644(.a(gate137inter12), .b(gate137inter1), .O(G522));
nand2 gate138( .a(G432), .b(G435), .O(G525) );
nand2 gate139( .a(G438), .b(G441), .O(G528) );
nand2 gate140( .a(G444), .b(G447), .O(G531) );
nand2 gate141( .a(G450), .b(G453), .O(G534) );

  xor2  gate883(.a(G459), .b(G456), .O(gate142inter0));
  nand2 gate884(.a(gate142inter0), .b(s_48), .O(gate142inter1));
  and2  gate885(.a(G459), .b(G456), .O(gate142inter2));
  inv1  gate886(.a(s_48), .O(gate142inter3));
  inv1  gate887(.a(s_49), .O(gate142inter4));
  nand2 gate888(.a(gate142inter4), .b(gate142inter3), .O(gate142inter5));
  nor2  gate889(.a(gate142inter5), .b(gate142inter2), .O(gate142inter6));
  inv1  gate890(.a(G456), .O(gate142inter7));
  inv1  gate891(.a(G459), .O(gate142inter8));
  nand2 gate892(.a(gate142inter8), .b(gate142inter7), .O(gate142inter9));
  nand2 gate893(.a(s_49), .b(gate142inter3), .O(gate142inter10));
  nor2  gate894(.a(gate142inter10), .b(gate142inter9), .O(gate142inter11));
  nor2  gate895(.a(gate142inter11), .b(gate142inter6), .O(gate142inter12));
  nand2 gate896(.a(gate142inter12), .b(gate142inter1), .O(G537));
nand2 gate143( .a(G462), .b(G465), .O(G540) );
nand2 gate144( .a(G468), .b(G471), .O(G543) );
nand2 gate145( .a(G474), .b(G477), .O(G546) );

  xor2  gate925(.a(G483), .b(G480), .O(gate146inter0));
  nand2 gate926(.a(gate146inter0), .b(s_54), .O(gate146inter1));
  and2  gate927(.a(G483), .b(G480), .O(gate146inter2));
  inv1  gate928(.a(s_54), .O(gate146inter3));
  inv1  gate929(.a(s_55), .O(gate146inter4));
  nand2 gate930(.a(gate146inter4), .b(gate146inter3), .O(gate146inter5));
  nor2  gate931(.a(gate146inter5), .b(gate146inter2), .O(gate146inter6));
  inv1  gate932(.a(G480), .O(gate146inter7));
  inv1  gate933(.a(G483), .O(gate146inter8));
  nand2 gate934(.a(gate146inter8), .b(gate146inter7), .O(gate146inter9));
  nand2 gate935(.a(s_55), .b(gate146inter3), .O(gate146inter10));
  nor2  gate936(.a(gate146inter10), .b(gate146inter9), .O(gate146inter11));
  nor2  gate937(.a(gate146inter11), .b(gate146inter6), .O(gate146inter12));
  nand2 gate938(.a(gate146inter12), .b(gate146inter1), .O(G549));
nand2 gate147( .a(G486), .b(G489), .O(G552) );

  xor2  gate1037(.a(G495), .b(G492), .O(gate148inter0));
  nand2 gate1038(.a(gate148inter0), .b(s_70), .O(gate148inter1));
  and2  gate1039(.a(G495), .b(G492), .O(gate148inter2));
  inv1  gate1040(.a(s_70), .O(gate148inter3));
  inv1  gate1041(.a(s_71), .O(gate148inter4));
  nand2 gate1042(.a(gate148inter4), .b(gate148inter3), .O(gate148inter5));
  nor2  gate1043(.a(gate148inter5), .b(gate148inter2), .O(gate148inter6));
  inv1  gate1044(.a(G492), .O(gate148inter7));
  inv1  gate1045(.a(G495), .O(gate148inter8));
  nand2 gate1046(.a(gate148inter8), .b(gate148inter7), .O(gate148inter9));
  nand2 gate1047(.a(s_71), .b(gate148inter3), .O(gate148inter10));
  nor2  gate1048(.a(gate148inter10), .b(gate148inter9), .O(gate148inter11));
  nor2  gate1049(.a(gate148inter11), .b(gate148inter6), .O(gate148inter12));
  nand2 gate1050(.a(gate148inter12), .b(gate148inter1), .O(G555));
nand2 gate149( .a(G498), .b(G501), .O(G558) );
nand2 gate150( .a(G504), .b(G507), .O(G561) );
nand2 gate151( .a(G510), .b(G513), .O(G564) );

  xor2  gate771(.a(G519), .b(G516), .O(gate152inter0));
  nand2 gate772(.a(gate152inter0), .b(s_32), .O(gate152inter1));
  and2  gate773(.a(G519), .b(G516), .O(gate152inter2));
  inv1  gate774(.a(s_32), .O(gate152inter3));
  inv1  gate775(.a(s_33), .O(gate152inter4));
  nand2 gate776(.a(gate152inter4), .b(gate152inter3), .O(gate152inter5));
  nor2  gate777(.a(gate152inter5), .b(gate152inter2), .O(gate152inter6));
  inv1  gate778(.a(G516), .O(gate152inter7));
  inv1  gate779(.a(G519), .O(gate152inter8));
  nand2 gate780(.a(gate152inter8), .b(gate152inter7), .O(gate152inter9));
  nand2 gate781(.a(s_33), .b(gate152inter3), .O(gate152inter10));
  nor2  gate782(.a(gate152inter10), .b(gate152inter9), .O(gate152inter11));
  nor2  gate783(.a(gate152inter11), .b(gate152inter6), .O(gate152inter12));
  nand2 gate784(.a(gate152inter12), .b(gate152inter1), .O(G567));
nand2 gate153( .a(G426), .b(G522), .O(G570) );
nand2 gate154( .a(G429), .b(G522), .O(G571) );
nand2 gate155( .a(G432), .b(G525), .O(G572) );
nand2 gate156( .a(G435), .b(G525), .O(G573) );
nand2 gate157( .a(G438), .b(G528), .O(G574) );
nand2 gate158( .a(G441), .b(G528), .O(G575) );
nand2 gate159( .a(G444), .b(G531), .O(G576) );
nand2 gate160( .a(G447), .b(G531), .O(G577) );
nand2 gate161( .a(G450), .b(G534), .O(G578) );
nand2 gate162( .a(G453), .b(G534), .O(G579) );
nand2 gate163( .a(G456), .b(G537), .O(G580) );
nand2 gate164( .a(G459), .b(G537), .O(G581) );
nand2 gate165( .a(G462), .b(G540), .O(G582) );
nand2 gate166( .a(G465), .b(G540), .O(G583) );
nand2 gate167( .a(G468), .b(G543), .O(G584) );
nand2 gate168( .a(G471), .b(G543), .O(G585) );
nand2 gate169( .a(G474), .b(G546), .O(G586) );
nand2 gate170( .a(G477), .b(G546), .O(G587) );

  xor2  gate841(.a(G549), .b(G480), .O(gate171inter0));
  nand2 gate842(.a(gate171inter0), .b(s_42), .O(gate171inter1));
  and2  gate843(.a(G549), .b(G480), .O(gate171inter2));
  inv1  gate844(.a(s_42), .O(gate171inter3));
  inv1  gate845(.a(s_43), .O(gate171inter4));
  nand2 gate846(.a(gate171inter4), .b(gate171inter3), .O(gate171inter5));
  nor2  gate847(.a(gate171inter5), .b(gate171inter2), .O(gate171inter6));
  inv1  gate848(.a(G480), .O(gate171inter7));
  inv1  gate849(.a(G549), .O(gate171inter8));
  nand2 gate850(.a(gate171inter8), .b(gate171inter7), .O(gate171inter9));
  nand2 gate851(.a(s_43), .b(gate171inter3), .O(gate171inter10));
  nor2  gate852(.a(gate171inter10), .b(gate171inter9), .O(gate171inter11));
  nor2  gate853(.a(gate171inter11), .b(gate171inter6), .O(gate171inter12));
  nand2 gate854(.a(gate171inter12), .b(gate171inter1), .O(G588));
nand2 gate172( .a(G483), .b(G549), .O(G589) );
nand2 gate173( .a(G486), .b(G552), .O(G590) );
nand2 gate174( .a(G489), .b(G552), .O(G591) );
nand2 gate175( .a(G492), .b(G555), .O(G592) );
nand2 gate176( .a(G495), .b(G555), .O(G593) );
nand2 gate177( .a(G498), .b(G558), .O(G594) );
nand2 gate178( .a(G501), .b(G558), .O(G595) );
nand2 gate179( .a(G504), .b(G561), .O(G596) );
nand2 gate180( .a(G507), .b(G561), .O(G597) );

  xor2  gate1023(.a(G564), .b(G510), .O(gate181inter0));
  nand2 gate1024(.a(gate181inter0), .b(s_68), .O(gate181inter1));
  and2  gate1025(.a(G564), .b(G510), .O(gate181inter2));
  inv1  gate1026(.a(s_68), .O(gate181inter3));
  inv1  gate1027(.a(s_69), .O(gate181inter4));
  nand2 gate1028(.a(gate181inter4), .b(gate181inter3), .O(gate181inter5));
  nor2  gate1029(.a(gate181inter5), .b(gate181inter2), .O(gate181inter6));
  inv1  gate1030(.a(G510), .O(gate181inter7));
  inv1  gate1031(.a(G564), .O(gate181inter8));
  nand2 gate1032(.a(gate181inter8), .b(gate181inter7), .O(gate181inter9));
  nand2 gate1033(.a(s_69), .b(gate181inter3), .O(gate181inter10));
  nor2  gate1034(.a(gate181inter10), .b(gate181inter9), .O(gate181inter11));
  nor2  gate1035(.a(gate181inter11), .b(gate181inter6), .O(gate181inter12));
  nand2 gate1036(.a(gate181inter12), .b(gate181inter1), .O(G598));
nand2 gate182( .a(G513), .b(G564), .O(G599) );
nand2 gate183( .a(G516), .b(G567), .O(G600) );
nand2 gate184( .a(G519), .b(G567), .O(G601) );
nand2 gate185( .a(G570), .b(G571), .O(G602) );
nand2 gate186( .a(G572), .b(G573), .O(G607) );
nand2 gate187( .a(G574), .b(G575), .O(G612) );
nand2 gate188( .a(G576), .b(G577), .O(G617) );
nand2 gate189( .a(G578), .b(G579), .O(G622) );
nand2 gate190( .a(G580), .b(G581), .O(G627) );
nand2 gate191( .a(G582), .b(G583), .O(G632) );
nand2 gate192( .a(G584), .b(G585), .O(G637) );
nand2 gate193( .a(G586), .b(G587), .O(G642) );
nand2 gate194( .a(G588), .b(G589), .O(G645) );
nand2 gate195( .a(G590), .b(G591), .O(G648) );
nand2 gate196( .a(G592), .b(G593), .O(G651) );
nand2 gate197( .a(G594), .b(G595), .O(G654) );

  xor2  gate547(.a(G597), .b(G596), .O(gate198inter0));
  nand2 gate548(.a(gate198inter0), .b(s_0), .O(gate198inter1));
  and2  gate549(.a(G597), .b(G596), .O(gate198inter2));
  inv1  gate550(.a(s_0), .O(gate198inter3));
  inv1  gate551(.a(s_1), .O(gate198inter4));
  nand2 gate552(.a(gate198inter4), .b(gate198inter3), .O(gate198inter5));
  nor2  gate553(.a(gate198inter5), .b(gate198inter2), .O(gate198inter6));
  inv1  gate554(.a(G596), .O(gate198inter7));
  inv1  gate555(.a(G597), .O(gate198inter8));
  nand2 gate556(.a(gate198inter8), .b(gate198inter7), .O(gate198inter9));
  nand2 gate557(.a(s_1), .b(gate198inter3), .O(gate198inter10));
  nor2  gate558(.a(gate198inter10), .b(gate198inter9), .O(gate198inter11));
  nor2  gate559(.a(gate198inter11), .b(gate198inter6), .O(gate198inter12));
  nand2 gate560(.a(gate198inter12), .b(gate198inter1), .O(G657));
nand2 gate199( .a(G598), .b(G599), .O(G660) );

  xor2  gate1079(.a(G601), .b(G600), .O(gate200inter0));
  nand2 gate1080(.a(gate200inter0), .b(s_76), .O(gate200inter1));
  and2  gate1081(.a(G601), .b(G600), .O(gate200inter2));
  inv1  gate1082(.a(s_76), .O(gate200inter3));
  inv1  gate1083(.a(s_77), .O(gate200inter4));
  nand2 gate1084(.a(gate200inter4), .b(gate200inter3), .O(gate200inter5));
  nor2  gate1085(.a(gate200inter5), .b(gate200inter2), .O(gate200inter6));
  inv1  gate1086(.a(G600), .O(gate200inter7));
  inv1  gate1087(.a(G601), .O(gate200inter8));
  nand2 gate1088(.a(gate200inter8), .b(gate200inter7), .O(gate200inter9));
  nand2 gate1089(.a(s_77), .b(gate200inter3), .O(gate200inter10));
  nor2  gate1090(.a(gate200inter10), .b(gate200inter9), .O(gate200inter11));
  nor2  gate1091(.a(gate200inter11), .b(gate200inter6), .O(gate200inter12));
  nand2 gate1092(.a(gate200inter12), .b(gate200inter1), .O(G663));
nand2 gate201( .a(G602), .b(G607), .O(G666) );
nand2 gate202( .a(G612), .b(G617), .O(G669) );
nand2 gate203( .a(G602), .b(G612), .O(G672) );
nand2 gate204( .a(G607), .b(G617), .O(G675) );

  xor2  gate701(.a(G627), .b(G622), .O(gate205inter0));
  nand2 gate702(.a(gate205inter0), .b(s_22), .O(gate205inter1));
  and2  gate703(.a(G627), .b(G622), .O(gate205inter2));
  inv1  gate704(.a(s_22), .O(gate205inter3));
  inv1  gate705(.a(s_23), .O(gate205inter4));
  nand2 gate706(.a(gate205inter4), .b(gate205inter3), .O(gate205inter5));
  nor2  gate707(.a(gate205inter5), .b(gate205inter2), .O(gate205inter6));
  inv1  gate708(.a(G622), .O(gate205inter7));
  inv1  gate709(.a(G627), .O(gate205inter8));
  nand2 gate710(.a(gate205inter8), .b(gate205inter7), .O(gate205inter9));
  nand2 gate711(.a(s_23), .b(gate205inter3), .O(gate205inter10));
  nor2  gate712(.a(gate205inter10), .b(gate205inter9), .O(gate205inter11));
  nor2  gate713(.a(gate205inter11), .b(gate205inter6), .O(gate205inter12));
  nand2 gate714(.a(gate205inter12), .b(gate205inter1), .O(G678));
nand2 gate206( .a(G632), .b(G637), .O(G681) );
nand2 gate207( .a(G622), .b(G632), .O(G684) );

  xor2  gate1233(.a(G637), .b(G627), .O(gate208inter0));
  nand2 gate1234(.a(gate208inter0), .b(s_98), .O(gate208inter1));
  and2  gate1235(.a(G637), .b(G627), .O(gate208inter2));
  inv1  gate1236(.a(s_98), .O(gate208inter3));
  inv1  gate1237(.a(s_99), .O(gate208inter4));
  nand2 gate1238(.a(gate208inter4), .b(gate208inter3), .O(gate208inter5));
  nor2  gate1239(.a(gate208inter5), .b(gate208inter2), .O(gate208inter6));
  inv1  gate1240(.a(G627), .O(gate208inter7));
  inv1  gate1241(.a(G637), .O(gate208inter8));
  nand2 gate1242(.a(gate208inter8), .b(gate208inter7), .O(gate208inter9));
  nand2 gate1243(.a(s_99), .b(gate208inter3), .O(gate208inter10));
  nor2  gate1244(.a(gate208inter10), .b(gate208inter9), .O(gate208inter11));
  nor2  gate1245(.a(gate208inter11), .b(gate208inter6), .O(gate208inter12));
  nand2 gate1246(.a(gate208inter12), .b(gate208inter1), .O(G687));
nand2 gate209( .a(G602), .b(G666), .O(G690) );
nand2 gate210( .a(G607), .b(G666), .O(G691) );
nand2 gate211( .a(G612), .b(G669), .O(G692) );
nand2 gate212( .a(G617), .b(G669), .O(G693) );
nand2 gate213( .a(G602), .b(G672), .O(G694) );
nand2 gate214( .a(G612), .b(G672), .O(G695) );
nand2 gate215( .a(G607), .b(G675), .O(G696) );
nand2 gate216( .a(G617), .b(G675), .O(G697) );
nand2 gate217( .a(G622), .b(G678), .O(G698) );
nand2 gate218( .a(G627), .b(G678), .O(G699) );
nand2 gate219( .a(G632), .b(G681), .O(G700) );
nand2 gate220( .a(G637), .b(G681), .O(G701) );
nand2 gate221( .a(G622), .b(G684), .O(G702) );
nand2 gate222( .a(G632), .b(G684), .O(G703) );
nand2 gate223( .a(G627), .b(G687), .O(G704) );
nand2 gate224( .a(G637), .b(G687), .O(G705) );
nand2 gate225( .a(G690), .b(G691), .O(G706) );
nand2 gate226( .a(G692), .b(G693), .O(G709) );
nand2 gate227( .a(G694), .b(G695), .O(G712) );
nand2 gate228( .a(G696), .b(G697), .O(G715) );
nand2 gate229( .a(G698), .b(G699), .O(G718) );
nand2 gate230( .a(G700), .b(G701), .O(G721) );
nand2 gate231( .a(G702), .b(G703), .O(G724) );
nand2 gate232( .a(G704), .b(G705), .O(G727) );
nand2 gate233( .a(G242), .b(G718), .O(G730) );
nand2 gate234( .a(G245), .b(G721), .O(G733) );
nand2 gate235( .a(G248), .b(G724), .O(G736) );

  xor2  gate813(.a(G727), .b(G251), .O(gate236inter0));
  nand2 gate814(.a(gate236inter0), .b(s_38), .O(gate236inter1));
  and2  gate815(.a(G727), .b(G251), .O(gate236inter2));
  inv1  gate816(.a(s_38), .O(gate236inter3));
  inv1  gate817(.a(s_39), .O(gate236inter4));
  nand2 gate818(.a(gate236inter4), .b(gate236inter3), .O(gate236inter5));
  nor2  gate819(.a(gate236inter5), .b(gate236inter2), .O(gate236inter6));
  inv1  gate820(.a(G251), .O(gate236inter7));
  inv1  gate821(.a(G727), .O(gate236inter8));
  nand2 gate822(.a(gate236inter8), .b(gate236inter7), .O(gate236inter9));
  nand2 gate823(.a(s_39), .b(gate236inter3), .O(gate236inter10));
  nor2  gate824(.a(gate236inter10), .b(gate236inter9), .O(gate236inter11));
  nor2  gate825(.a(gate236inter11), .b(gate236inter6), .O(gate236inter12));
  nand2 gate826(.a(gate236inter12), .b(gate236inter1), .O(G739));
nand2 gate237( .a(G254), .b(G706), .O(G742) );
nand2 gate238( .a(G257), .b(G709), .O(G745) );
nand2 gate239( .a(G260), .b(G712), .O(G748) );
nand2 gate240( .a(G263), .b(G715), .O(G751) );
nand2 gate241( .a(G242), .b(G730), .O(G754) );
nand2 gate242( .a(G718), .b(G730), .O(G755) );
nand2 gate243( .a(G245), .b(G733), .O(G756) );
nand2 gate244( .a(G721), .b(G733), .O(G757) );

  xor2  gate981(.a(G736), .b(G248), .O(gate245inter0));
  nand2 gate982(.a(gate245inter0), .b(s_62), .O(gate245inter1));
  and2  gate983(.a(G736), .b(G248), .O(gate245inter2));
  inv1  gate984(.a(s_62), .O(gate245inter3));
  inv1  gate985(.a(s_63), .O(gate245inter4));
  nand2 gate986(.a(gate245inter4), .b(gate245inter3), .O(gate245inter5));
  nor2  gate987(.a(gate245inter5), .b(gate245inter2), .O(gate245inter6));
  inv1  gate988(.a(G248), .O(gate245inter7));
  inv1  gate989(.a(G736), .O(gate245inter8));
  nand2 gate990(.a(gate245inter8), .b(gate245inter7), .O(gate245inter9));
  nand2 gate991(.a(s_63), .b(gate245inter3), .O(gate245inter10));
  nor2  gate992(.a(gate245inter10), .b(gate245inter9), .O(gate245inter11));
  nor2  gate993(.a(gate245inter11), .b(gate245inter6), .O(gate245inter12));
  nand2 gate994(.a(gate245inter12), .b(gate245inter1), .O(G758));
nand2 gate246( .a(G724), .b(G736), .O(G759) );

  xor2  gate785(.a(G739), .b(G251), .O(gate247inter0));
  nand2 gate786(.a(gate247inter0), .b(s_34), .O(gate247inter1));
  and2  gate787(.a(G739), .b(G251), .O(gate247inter2));
  inv1  gate788(.a(s_34), .O(gate247inter3));
  inv1  gate789(.a(s_35), .O(gate247inter4));
  nand2 gate790(.a(gate247inter4), .b(gate247inter3), .O(gate247inter5));
  nor2  gate791(.a(gate247inter5), .b(gate247inter2), .O(gate247inter6));
  inv1  gate792(.a(G251), .O(gate247inter7));
  inv1  gate793(.a(G739), .O(gate247inter8));
  nand2 gate794(.a(gate247inter8), .b(gate247inter7), .O(gate247inter9));
  nand2 gate795(.a(s_35), .b(gate247inter3), .O(gate247inter10));
  nor2  gate796(.a(gate247inter10), .b(gate247inter9), .O(gate247inter11));
  nor2  gate797(.a(gate247inter11), .b(gate247inter6), .O(gate247inter12));
  nand2 gate798(.a(gate247inter12), .b(gate247inter1), .O(G760));
nand2 gate248( .a(G727), .b(G739), .O(G761) );
nand2 gate249( .a(G254), .b(G742), .O(G762) );
nand2 gate250( .a(G706), .b(G742), .O(G763) );
nand2 gate251( .a(G257), .b(G745), .O(G764) );
nand2 gate252( .a(G709), .b(G745), .O(G765) );
nand2 gate253( .a(G260), .b(G748), .O(G766) );
nand2 gate254( .a(G712), .b(G748), .O(G767) );

  xor2  gate911(.a(G751), .b(G263), .O(gate255inter0));
  nand2 gate912(.a(gate255inter0), .b(s_52), .O(gate255inter1));
  and2  gate913(.a(G751), .b(G263), .O(gate255inter2));
  inv1  gate914(.a(s_52), .O(gate255inter3));
  inv1  gate915(.a(s_53), .O(gate255inter4));
  nand2 gate916(.a(gate255inter4), .b(gate255inter3), .O(gate255inter5));
  nor2  gate917(.a(gate255inter5), .b(gate255inter2), .O(gate255inter6));
  inv1  gate918(.a(G263), .O(gate255inter7));
  inv1  gate919(.a(G751), .O(gate255inter8));
  nand2 gate920(.a(gate255inter8), .b(gate255inter7), .O(gate255inter9));
  nand2 gate921(.a(s_53), .b(gate255inter3), .O(gate255inter10));
  nor2  gate922(.a(gate255inter10), .b(gate255inter9), .O(gate255inter11));
  nor2  gate923(.a(gate255inter11), .b(gate255inter6), .O(gate255inter12));
  nand2 gate924(.a(gate255inter12), .b(gate255inter1), .O(G768));
nand2 gate256( .a(G715), .b(G751), .O(G769) );

  xor2  gate1121(.a(G755), .b(G754), .O(gate257inter0));
  nand2 gate1122(.a(gate257inter0), .b(s_82), .O(gate257inter1));
  and2  gate1123(.a(G755), .b(G754), .O(gate257inter2));
  inv1  gate1124(.a(s_82), .O(gate257inter3));
  inv1  gate1125(.a(s_83), .O(gate257inter4));
  nand2 gate1126(.a(gate257inter4), .b(gate257inter3), .O(gate257inter5));
  nor2  gate1127(.a(gate257inter5), .b(gate257inter2), .O(gate257inter6));
  inv1  gate1128(.a(G754), .O(gate257inter7));
  inv1  gate1129(.a(G755), .O(gate257inter8));
  nand2 gate1130(.a(gate257inter8), .b(gate257inter7), .O(gate257inter9));
  nand2 gate1131(.a(s_83), .b(gate257inter3), .O(gate257inter10));
  nor2  gate1132(.a(gate257inter10), .b(gate257inter9), .O(gate257inter11));
  nor2  gate1133(.a(gate257inter11), .b(gate257inter6), .O(gate257inter12));
  nand2 gate1134(.a(gate257inter12), .b(gate257inter1), .O(G770));

  xor2  gate687(.a(G757), .b(G756), .O(gate258inter0));
  nand2 gate688(.a(gate258inter0), .b(s_20), .O(gate258inter1));
  and2  gate689(.a(G757), .b(G756), .O(gate258inter2));
  inv1  gate690(.a(s_20), .O(gate258inter3));
  inv1  gate691(.a(s_21), .O(gate258inter4));
  nand2 gate692(.a(gate258inter4), .b(gate258inter3), .O(gate258inter5));
  nor2  gate693(.a(gate258inter5), .b(gate258inter2), .O(gate258inter6));
  inv1  gate694(.a(G756), .O(gate258inter7));
  inv1  gate695(.a(G757), .O(gate258inter8));
  nand2 gate696(.a(gate258inter8), .b(gate258inter7), .O(gate258inter9));
  nand2 gate697(.a(s_21), .b(gate258inter3), .O(gate258inter10));
  nor2  gate698(.a(gate258inter10), .b(gate258inter9), .O(gate258inter11));
  nor2  gate699(.a(gate258inter11), .b(gate258inter6), .O(gate258inter12));
  nand2 gate700(.a(gate258inter12), .b(gate258inter1), .O(G773));
nand2 gate259( .a(G758), .b(G759), .O(G776) );
nand2 gate260( .a(G760), .b(G761), .O(G779) );
nand2 gate261( .a(G762), .b(G763), .O(G782) );
nand2 gate262( .a(G764), .b(G765), .O(G785) );
nand2 gate263( .a(G766), .b(G767), .O(G788) );
nand2 gate264( .a(G768), .b(G769), .O(G791) );
nand2 gate265( .a(G642), .b(G770), .O(G794) );
nand2 gate266( .a(G645), .b(G773), .O(G797) );
nand2 gate267( .a(G648), .b(G776), .O(G800) );
nand2 gate268( .a(G651), .b(G779), .O(G803) );
nand2 gate269( .a(G654), .b(G782), .O(G806) );
nand2 gate270( .a(G657), .b(G785), .O(G809) );
nand2 gate271( .a(G660), .b(G788), .O(G812) );
nand2 gate272( .a(G663), .b(G791), .O(G815) );
nand2 gate273( .a(G642), .b(G794), .O(G818) );
nand2 gate274( .a(G770), .b(G794), .O(G819) );
nand2 gate275( .a(G645), .b(G797), .O(G820) );
nand2 gate276( .a(G773), .b(G797), .O(G821) );
nand2 gate277( .a(G648), .b(G800), .O(G822) );

  xor2  gate645(.a(G800), .b(G776), .O(gate278inter0));
  nand2 gate646(.a(gate278inter0), .b(s_14), .O(gate278inter1));
  and2  gate647(.a(G800), .b(G776), .O(gate278inter2));
  inv1  gate648(.a(s_14), .O(gate278inter3));
  inv1  gate649(.a(s_15), .O(gate278inter4));
  nand2 gate650(.a(gate278inter4), .b(gate278inter3), .O(gate278inter5));
  nor2  gate651(.a(gate278inter5), .b(gate278inter2), .O(gate278inter6));
  inv1  gate652(.a(G776), .O(gate278inter7));
  inv1  gate653(.a(G800), .O(gate278inter8));
  nand2 gate654(.a(gate278inter8), .b(gate278inter7), .O(gate278inter9));
  nand2 gate655(.a(s_15), .b(gate278inter3), .O(gate278inter10));
  nor2  gate656(.a(gate278inter10), .b(gate278inter9), .O(gate278inter11));
  nor2  gate657(.a(gate278inter11), .b(gate278inter6), .O(gate278inter12));
  nand2 gate658(.a(gate278inter12), .b(gate278inter1), .O(G823));
nand2 gate279( .a(G651), .b(G803), .O(G824) );
nand2 gate280( .a(G779), .b(G803), .O(G825) );
nand2 gate281( .a(G654), .b(G806), .O(G826) );
nand2 gate282( .a(G782), .b(G806), .O(G827) );
nand2 gate283( .a(G657), .b(G809), .O(G828) );
nand2 gate284( .a(G785), .b(G809), .O(G829) );
nand2 gate285( .a(G660), .b(G812), .O(G830) );
nand2 gate286( .a(G788), .b(G812), .O(G831) );
nand2 gate287( .a(G663), .b(G815), .O(G832) );
nand2 gate288( .a(G791), .b(G815), .O(G833) );
nand2 gate289( .a(G818), .b(G819), .O(G834) );
nand2 gate290( .a(G820), .b(G821), .O(G847) );
nand2 gate291( .a(G822), .b(G823), .O(G860) );
nand2 gate292( .a(G824), .b(G825), .O(G873) );
nand2 gate293( .a(G828), .b(G829), .O(G886) );

  xor2  gate995(.a(G833), .b(G832), .O(gate294inter0));
  nand2 gate996(.a(gate294inter0), .b(s_64), .O(gate294inter1));
  and2  gate997(.a(G833), .b(G832), .O(gate294inter2));
  inv1  gate998(.a(s_64), .O(gate294inter3));
  inv1  gate999(.a(s_65), .O(gate294inter4));
  nand2 gate1000(.a(gate294inter4), .b(gate294inter3), .O(gate294inter5));
  nor2  gate1001(.a(gate294inter5), .b(gate294inter2), .O(gate294inter6));
  inv1  gate1002(.a(G832), .O(gate294inter7));
  inv1  gate1003(.a(G833), .O(gate294inter8));
  nand2 gate1004(.a(gate294inter8), .b(gate294inter7), .O(gate294inter9));
  nand2 gate1005(.a(s_65), .b(gate294inter3), .O(gate294inter10));
  nor2  gate1006(.a(gate294inter10), .b(gate294inter9), .O(gate294inter11));
  nor2  gate1007(.a(gate294inter11), .b(gate294inter6), .O(gate294inter12));
  nand2 gate1008(.a(gate294inter12), .b(gate294inter1), .O(G899));
nand2 gate295( .a(G830), .b(G831), .O(G912) );

  xor2  gate1177(.a(G827), .b(G826), .O(gate296inter0));
  nand2 gate1178(.a(gate296inter0), .b(s_90), .O(gate296inter1));
  and2  gate1179(.a(G827), .b(G826), .O(gate296inter2));
  inv1  gate1180(.a(s_90), .O(gate296inter3));
  inv1  gate1181(.a(s_91), .O(gate296inter4));
  nand2 gate1182(.a(gate296inter4), .b(gate296inter3), .O(gate296inter5));
  nor2  gate1183(.a(gate296inter5), .b(gate296inter2), .O(gate296inter6));
  inv1  gate1184(.a(G826), .O(gate296inter7));
  inv1  gate1185(.a(G827), .O(gate296inter8));
  nand2 gate1186(.a(gate296inter8), .b(gate296inter7), .O(gate296inter9));
  nand2 gate1187(.a(s_91), .b(gate296inter3), .O(gate296inter10));
  nor2  gate1188(.a(gate296inter10), .b(gate296inter9), .O(gate296inter11));
  nor2  gate1189(.a(gate296inter11), .b(gate296inter6), .O(gate296inter12));
  nand2 gate1190(.a(gate296inter12), .b(gate296inter1), .O(G925));
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );
nand2 gate387( .a(G1), .b(G1036), .O(G1132) );
nand2 gate388( .a(G2), .b(G1039), .O(G1135) );
nand2 gate389( .a(G3), .b(G1042), .O(G1138) );
nand2 gate390( .a(G4), .b(G1045), .O(G1141) );
nand2 gate391( .a(G5), .b(G1048), .O(G1144) );
nand2 gate392( .a(G6), .b(G1051), .O(G1147) );
nand2 gate393( .a(G7), .b(G1054), .O(G1150) );
nand2 gate394( .a(G8), .b(G1057), .O(G1153) );
nand2 gate395( .a(G9), .b(G1060), .O(G1156) );
nand2 gate396( .a(G10), .b(G1063), .O(G1159) );
nand2 gate397( .a(G11), .b(G1066), .O(G1162) );

  xor2  gate575(.a(G1069), .b(G12), .O(gate398inter0));
  nand2 gate576(.a(gate398inter0), .b(s_4), .O(gate398inter1));
  and2  gate577(.a(G1069), .b(G12), .O(gate398inter2));
  inv1  gate578(.a(s_4), .O(gate398inter3));
  inv1  gate579(.a(s_5), .O(gate398inter4));
  nand2 gate580(.a(gate398inter4), .b(gate398inter3), .O(gate398inter5));
  nor2  gate581(.a(gate398inter5), .b(gate398inter2), .O(gate398inter6));
  inv1  gate582(.a(G12), .O(gate398inter7));
  inv1  gate583(.a(G1069), .O(gate398inter8));
  nand2 gate584(.a(gate398inter8), .b(gate398inter7), .O(gate398inter9));
  nand2 gate585(.a(s_5), .b(gate398inter3), .O(gate398inter10));
  nor2  gate586(.a(gate398inter10), .b(gate398inter9), .O(gate398inter11));
  nor2  gate587(.a(gate398inter11), .b(gate398inter6), .O(gate398inter12));
  nand2 gate588(.a(gate398inter12), .b(gate398inter1), .O(G1165));
nand2 gate399( .a(G13), .b(G1072), .O(G1168) );
nand2 gate400( .a(G14), .b(G1075), .O(G1171) );
nand2 gate401( .a(G15), .b(G1078), .O(G1174) );
nand2 gate402( .a(G16), .b(G1081), .O(G1177) );
nand2 gate403( .a(G17), .b(G1084), .O(G1180) );
nand2 gate404( .a(G18), .b(G1087), .O(G1183) );
nand2 gate405( .a(G19), .b(G1090), .O(G1186) );
nand2 gate406( .a(G20), .b(G1093), .O(G1189) );

  xor2  gate603(.a(G1096), .b(G21), .O(gate407inter0));
  nand2 gate604(.a(gate407inter0), .b(s_8), .O(gate407inter1));
  and2  gate605(.a(G1096), .b(G21), .O(gate407inter2));
  inv1  gate606(.a(s_8), .O(gate407inter3));
  inv1  gate607(.a(s_9), .O(gate407inter4));
  nand2 gate608(.a(gate407inter4), .b(gate407inter3), .O(gate407inter5));
  nor2  gate609(.a(gate407inter5), .b(gate407inter2), .O(gate407inter6));
  inv1  gate610(.a(G21), .O(gate407inter7));
  inv1  gate611(.a(G1096), .O(gate407inter8));
  nand2 gate612(.a(gate407inter8), .b(gate407inter7), .O(gate407inter9));
  nand2 gate613(.a(s_9), .b(gate407inter3), .O(gate407inter10));
  nor2  gate614(.a(gate407inter10), .b(gate407inter9), .O(gate407inter11));
  nor2  gate615(.a(gate407inter11), .b(gate407inter6), .O(gate407inter12));
  nand2 gate616(.a(gate407inter12), .b(gate407inter1), .O(G1192));
nand2 gate408( .a(G22), .b(G1099), .O(G1195) );
nand2 gate409( .a(G23), .b(G1102), .O(G1198) );
nand2 gate410( .a(G24), .b(G1105), .O(G1201) );
nand2 gate411( .a(G25), .b(G1108), .O(G1204) );
nand2 gate412( .a(G26), .b(G1111), .O(G1207) );
nand2 gate413( .a(G27), .b(G1114), .O(G1210) );
nand2 gate414( .a(G28), .b(G1117), .O(G1213) );
nand2 gate415( .a(G29), .b(G1120), .O(G1216) );
nand2 gate416( .a(G30), .b(G1123), .O(G1219) );
nand2 gate417( .a(G31), .b(G1126), .O(G1222) );
nand2 gate418( .a(G32), .b(G1129), .O(G1225) );
nand2 gate419( .a(G1), .b(G1132), .O(G1228) );
nand2 gate420( .a(G1036), .b(G1132), .O(G1229) );

  xor2  gate743(.a(G1135), .b(G2), .O(gate421inter0));
  nand2 gate744(.a(gate421inter0), .b(s_28), .O(gate421inter1));
  and2  gate745(.a(G1135), .b(G2), .O(gate421inter2));
  inv1  gate746(.a(s_28), .O(gate421inter3));
  inv1  gate747(.a(s_29), .O(gate421inter4));
  nand2 gate748(.a(gate421inter4), .b(gate421inter3), .O(gate421inter5));
  nor2  gate749(.a(gate421inter5), .b(gate421inter2), .O(gate421inter6));
  inv1  gate750(.a(G2), .O(gate421inter7));
  inv1  gate751(.a(G1135), .O(gate421inter8));
  nand2 gate752(.a(gate421inter8), .b(gate421inter7), .O(gate421inter9));
  nand2 gate753(.a(s_29), .b(gate421inter3), .O(gate421inter10));
  nor2  gate754(.a(gate421inter10), .b(gate421inter9), .O(gate421inter11));
  nor2  gate755(.a(gate421inter11), .b(gate421inter6), .O(gate421inter12));
  nand2 gate756(.a(gate421inter12), .b(gate421inter1), .O(G1230));
nand2 gate422( .a(G1039), .b(G1135), .O(G1231) );
nand2 gate423( .a(G3), .b(G1138), .O(G1232) );

  xor2  gate939(.a(G1138), .b(G1042), .O(gate424inter0));
  nand2 gate940(.a(gate424inter0), .b(s_56), .O(gate424inter1));
  and2  gate941(.a(G1138), .b(G1042), .O(gate424inter2));
  inv1  gate942(.a(s_56), .O(gate424inter3));
  inv1  gate943(.a(s_57), .O(gate424inter4));
  nand2 gate944(.a(gate424inter4), .b(gate424inter3), .O(gate424inter5));
  nor2  gate945(.a(gate424inter5), .b(gate424inter2), .O(gate424inter6));
  inv1  gate946(.a(G1042), .O(gate424inter7));
  inv1  gate947(.a(G1138), .O(gate424inter8));
  nand2 gate948(.a(gate424inter8), .b(gate424inter7), .O(gate424inter9));
  nand2 gate949(.a(s_57), .b(gate424inter3), .O(gate424inter10));
  nor2  gate950(.a(gate424inter10), .b(gate424inter9), .O(gate424inter11));
  nor2  gate951(.a(gate424inter11), .b(gate424inter6), .O(gate424inter12));
  nand2 gate952(.a(gate424inter12), .b(gate424inter1), .O(G1233));
nand2 gate425( .a(G4), .b(G1141), .O(G1234) );
nand2 gate426( .a(G1045), .b(G1141), .O(G1235) );
nand2 gate427( .a(G5), .b(G1144), .O(G1236) );
nand2 gate428( .a(G1048), .b(G1144), .O(G1237) );
nand2 gate429( .a(G6), .b(G1147), .O(G1238) );
nand2 gate430( .a(G1051), .b(G1147), .O(G1239) );
nand2 gate431( .a(G7), .b(G1150), .O(G1240) );
nand2 gate432( .a(G1054), .b(G1150), .O(G1241) );
nand2 gate433( .a(G8), .b(G1153), .O(G1242) );
nand2 gate434( .a(G1057), .b(G1153), .O(G1243) );
nand2 gate435( .a(G9), .b(G1156), .O(G1244) );
nand2 gate436( .a(G1060), .b(G1156), .O(G1245) );
nand2 gate437( .a(G10), .b(G1159), .O(G1246) );

  xor2  gate799(.a(G1159), .b(G1063), .O(gate438inter0));
  nand2 gate800(.a(gate438inter0), .b(s_36), .O(gate438inter1));
  and2  gate801(.a(G1159), .b(G1063), .O(gate438inter2));
  inv1  gate802(.a(s_36), .O(gate438inter3));
  inv1  gate803(.a(s_37), .O(gate438inter4));
  nand2 gate804(.a(gate438inter4), .b(gate438inter3), .O(gate438inter5));
  nor2  gate805(.a(gate438inter5), .b(gate438inter2), .O(gate438inter6));
  inv1  gate806(.a(G1063), .O(gate438inter7));
  inv1  gate807(.a(G1159), .O(gate438inter8));
  nand2 gate808(.a(gate438inter8), .b(gate438inter7), .O(gate438inter9));
  nand2 gate809(.a(s_37), .b(gate438inter3), .O(gate438inter10));
  nor2  gate810(.a(gate438inter10), .b(gate438inter9), .O(gate438inter11));
  nor2  gate811(.a(gate438inter11), .b(gate438inter6), .O(gate438inter12));
  nand2 gate812(.a(gate438inter12), .b(gate438inter1), .O(G1247));
nand2 gate439( .a(G11), .b(G1162), .O(G1248) );
nand2 gate440( .a(G1066), .b(G1162), .O(G1249) );
nand2 gate441( .a(G12), .b(G1165), .O(G1250) );
nand2 gate442( .a(G1069), .b(G1165), .O(G1251) );
nand2 gate443( .a(G13), .b(G1168), .O(G1252) );
nand2 gate444( .a(G1072), .b(G1168), .O(G1253) );
nand2 gate445( .a(G14), .b(G1171), .O(G1254) );
nand2 gate446( .a(G1075), .b(G1171), .O(G1255) );
nand2 gate447( .a(G15), .b(G1174), .O(G1256) );
nand2 gate448( .a(G1078), .b(G1174), .O(G1257) );

  xor2  gate659(.a(G1177), .b(G16), .O(gate449inter0));
  nand2 gate660(.a(gate449inter0), .b(s_16), .O(gate449inter1));
  and2  gate661(.a(G1177), .b(G16), .O(gate449inter2));
  inv1  gate662(.a(s_16), .O(gate449inter3));
  inv1  gate663(.a(s_17), .O(gate449inter4));
  nand2 gate664(.a(gate449inter4), .b(gate449inter3), .O(gate449inter5));
  nor2  gate665(.a(gate449inter5), .b(gate449inter2), .O(gate449inter6));
  inv1  gate666(.a(G16), .O(gate449inter7));
  inv1  gate667(.a(G1177), .O(gate449inter8));
  nand2 gate668(.a(gate449inter8), .b(gate449inter7), .O(gate449inter9));
  nand2 gate669(.a(s_17), .b(gate449inter3), .O(gate449inter10));
  nor2  gate670(.a(gate449inter10), .b(gate449inter9), .O(gate449inter11));
  nor2  gate671(.a(gate449inter11), .b(gate449inter6), .O(gate449inter12));
  nand2 gate672(.a(gate449inter12), .b(gate449inter1), .O(G1258));
nand2 gate450( .a(G1081), .b(G1177), .O(G1259) );
nand2 gate451( .a(G17), .b(G1180), .O(G1260) );
nand2 gate452( .a(G1084), .b(G1180), .O(G1261) );
nand2 gate453( .a(G18), .b(G1183), .O(G1262) );
nand2 gate454( .a(G1087), .b(G1183), .O(G1263) );
nand2 gate455( .a(G19), .b(G1186), .O(G1264) );

  xor2  gate1107(.a(G1186), .b(G1090), .O(gate456inter0));
  nand2 gate1108(.a(gate456inter0), .b(s_80), .O(gate456inter1));
  and2  gate1109(.a(G1186), .b(G1090), .O(gate456inter2));
  inv1  gate1110(.a(s_80), .O(gate456inter3));
  inv1  gate1111(.a(s_81), .O(gate456inter4));
  nand2 gate1112(.a(gate456inter4), .b(gate456inter3), .O(gate456inter5));
  nor2  gate1113(.a(gate456inter5), .b(gate456inter2), .O(gate456inter6));
  inv1  gate1114(.a(G1090), .O(gate456inter7));
  inv1  gate1115(.a(G1186), .O(gate456inter8));
  nand2 gate1116(.a(gate456inter8), .b(gate456inter7), .O(gate456inter9));
  nand2 gate1117(.a(s_81), .b(gate456inter3), .O(gate456inter10));
  nor2  gate1118(.a(gate456inter10), .b(gate456inter9), .O(gate456inter11));
  nor2  gate1119(.a(gate456inter11), .b(gate456inter6), .O(gate456inter12));
  nand2 gate1120(.a(gate456inter12), .b(gate456inter1), .O(G1265));
nand2 gate457( .a(G20), .b(G1189), .O(G1266) );
nand2 gate458( .a(G1093), .b(G1189), .O(G1267) );
nand2 gate459( .a(G21), .b(G1192), .O(G1268) );
nand2 gate460( .a(G1096), .b(G1192), .O(G1269) );

  xor2  gate953(.a(G1195), .b(G22), .O(gate461inter0));
  nand2 gate954(.a(gate461inter0), .b(s_58), .O(gate461inter1));
  and2  gate955(.a(G1195), .b(G22), .O(gate461inter2));
  inv1  gate956(.a(s_58), .O(gate461inter3));
  inv1  gate957(.a(s_59), .O(gate461inter4));
  nand2 gate958(.a(gate461inter4), .b(gate461inter3), .O(gate461inter5));
  nor2  gate959(.a(gate461inter5), .b(gate461inter2), .O(gate461inter6));
  inv1  gate960(.a(G22), .O(gate461inter7));
  inv1  gate961(.a(G1195), .O(gate461inter8));
  nand2 gate962(.a(gate461inter8), .b(gate461inter7), .O(gate461inter9));
  nand2 gate963(.a(s_59), .b(gate461inter3), .O(gate461inter10));
  nor2  gate964(.a(gate461inter10), .b(gate461inter9), .O(gate461inter11));
  nor2  gate965(.a(gate461inter11), .b(gate461inter6), .O(gate461inter12));
  nand2 gate966(.a(gate461inter12), .b(gate461inter1), .O(G1270));
nand2 gate462( .a(G1099), .b(G1195), .O(G1271) );

  xor2  gate561(.a(G1198), .b(G23), .O(gate463inter0));
  nand2 gate562(.a(gate463inter0), .b(s_2), .O(gate463inter1));
  and2  gate563(.a(G1198), .b(G23), .O(gate463inter2));
  inv1  gate564(.a(s_2), .O(gate463inter3));
  inv1  gate565(.a(s_3), .O(gate463inter4));
  nand2 gate566(.a(gate463inter4), .b(gate463inter3), .O(gate463inter5));
  nor2  gate567(.a(gate463inter5), .b(gate463inter2), .O(gate463inter6));
  inv1  gate568(.a(G23), .O(gate463inter7));
  inv1  gate569(.a(G1198), .O(gate463inter8));
  nand2 gate570(.a(gate463inter8), .b(gate463inter7), .O(gate463inter9));
  nand2 gate571(.a(s_3), .b(gate463inter3), .O(gate463inter10));
  nor2  gate572(.a(gate463inter10), .b(gate463inter9), .O(gate463inter11));
  nor2  gate573(.a(gate463inter11), .b(gate463inter6), .O(gate463inter12));
  nand2 gate574(.a(gate463inter12), .b(gate463inter1), .O(G1272));
nand2 gate464( .a(G1102), .b(G1198), .O(G1273) );
nand2 gate465( .a(G24), .b(G1201), .O(G1274) );
nand2 gate466( .a(G1105), .b(G1201), .O(G1275) );
nand2 gate467( .a(G25), .b(G1204), .O(G1276) );
nand2 gate468( .a(G1108), .b(G1204), .O(G1277) );
nand2 gate469( .a(G26), .b(G1207), .O(G1278) );
nand2 gate470( .a(G1111), .b(G1207), .O(G1279) );
nand2 gate471( .a(G27), .b(G1210), .O(G1280) );
nand2 gate472( .a(G1114), .b(G1210), .O(G1281) );

  xor2  gate1163(.a(G1213), .b(G28), .O(gate473inter0));
  nand2 gate1164(.a(gate473inter0), .b(s_88), .O(gate473inter1));
  and2  gate1165(.a(G1213), .b(G28), .O(gate473inter2));
  inv1  gate1166(.a(s_88), .O(gate473inter3));
  inv1  gate1167(.a(s_89), .O(gate473inter4));
  nand2 gate1168(.a(gate473inter4), .b(gate473inter3), .O(gate473inter5));
  nor2  gate1169(.a(gate473inter5), .b(gate473inter2), .O(gate473inter6));
  inv1  gate1170(.a(G28), .O(gate473inter7));
  inv1  gate1171(.a(G1213), .O(gate473inter8));
  nand2 gate1172(.a(gate473inter8), .b(gate473inter7), .O(gate473inter9));
  nand2 gate1173(.a(s_89), .b(gate473inter3), .O(gate473inter10));
  nor2  gate1174(.a(gate473inter10), .b(gate473inter9), .O(gate473inter11));
  nor2  gate1175(.a(gate473inter11), .b(gate473inter6), .O(gate473inter12));
  nand2 gate1176(.a(gate473inter12), .b(gate473inter1), .O(G1282));
nand2 gate474( .a(G1117), .b(G1213), .O(G1283) );
nand2 gate475( .a(G29), .b(G1216), .O(G1284) );
nand2 gate476( .a(G1120), .b(G1216), .O(G1285) );
nand2 gate477( .a(G30), .b(G1219), .O(G1286) );
nand2 gate478( .a(G1123), .b(G1219), .O(G1287) );
nand2 gate479( .a(G31), .b(G1222), .O(G1288) );
nand2 gate480( .a(G1126), .b(G1222), .O(G1289) );
nand2 gate481( .a(G32), .b(G1225), .O(G1290) );
nand2 gate482( .a(G1129), .b(G1225), .O(G1291) );
nand2 gate483( .a(G1228), .b(G1229), .O(G1292) );
nand2 gate484( .a(G1230), .b(G1231), .O(G1293) );
nand2 gate485( .a(G1232), .b(G1233), .O(G1294) );
nand2 gate486( .a(G1234), .b(G1235), .O(G1295) );
nand2 gate487( .a(G1236), .b(G1237), .O(G1296) );
nand2 gate488( .a(G1238), .b(G1239), .O(G1297) );
nand2 gate489( .a(G1240), .b(G1241), .O(G1298) );
nand2 gate490( .a(G1242), .b(G1243), .O(G1299) );
nand2 gate491( .a(G1244), .b(G1245), .O(G1300) );
nand2 gate492( .a(G1246), .b(G1247), .O(G1301) );
nand2 gate493( .a(G1248), .b(G1249), .O(G1302) );
nand2 gate494( .a(G1250), .b(G1251), .O(G1303) );
nand2 gate495( .a(G1252), .b(G1253), .O(G1304) );
nand2 gate496( .a(G1254), .b(G1255), .O(G1305) );
nand2 gate497( .a(G1256), .b(G1257), .O(G1306) );
nand2 gate498( .a(G1258), .b(G1259), .O(G1307) );
nand2 gate499( .a(G1260), .b(G1261), .O(G1308) );
nand2 gate500( .a(G1262), .b(G1263), .O(G1309) );

  xor2  gate827(.a(G1265), .b(G1264), .O(gate501inter0));
  nand2 gate828(.a(gate501inter0), .b(s_40), .O(gate501inter1));
  and2  gate829(.a(G1265), .b(G1264), .O(gate501inter2));
  inv1  gate830(.a(s_40), .O(gate501inter3));
  inv1  gate831(.a(s_41), .O(gate501inter4));
  nand2 gate832(.a(gate501inter4), .b(gate501inter3), .O(gate501inter5));
  nor2  gate833(.a(gate501inter5), .b(gate501inter2), .O(gate501inter6));
  inv1  gate834(.a(G1264), .O(gate501inter7));
  inv1  gate835(.a(G1265), .O(gate501inter8));
  nand2 gate836(.a(gate501inter8), .b(gate501inter7), .O(gate501inter9));
  nand2 gate837(.a(s_41), .b(gate501inter3), .O(gate501inter10));
  nor2  gate838(.a(gate501inter10), .b(gate501inter9), .O(gate501inter11));
  nor2  gate839(.a(gate501inter11), .b(gate501inter6), .O(gate501inter12));
  nand2 gate840(.a(gate501inter12), .b(gate501inter1), .O(G1310));
nand2 gate502( .a(G1266), .b(G1267), .O(G1311) );

  xor2  gate1135(.a(G1269), .b(G1268), .O(gate503inter0));
  nand2 gate1136(.a(gate503inter0), .b(s_84), .O(gate503inter1));
  and2  gate1137(.a(G1269), .b(G1268), .O(gate503inter2));
  inv1  gate1138(.a(s_84), .O(gate503inter3));
  inv1  gate1139(.a(s_85), .O(gate503inter4));
  nand2 gate1140(.a(gate503inter4), .b(gate503inter3), .O(gate503inter5));
  nor2  gate1141(.a(gate503inter5), .b(gate503inter2), .O(gate503inter6));
  inv1  gate1142(.a(G1268), .O(gate503inter7));
  inv1  gate1143(.a(G1269), .O(gate503inter8));
  nand2 gate1144(.a(gate503inter8), .b(gate503inter7), .O(gate503inter9));
  nand2 gate1145(.a(s_85), .b(gate503inter3), .O(gate503inter10));
  nor2  gate1146(.a(gate503inter10), .b(gate503inter9), .O(gate503inter11));
  nor2  gate1147(.a(gate503inter11), .b(gate503inter6), .O(gate503inter12));
  nand2 gate1148(.a(gate503inter12), .b(gate503inter1), .O(G1312));

  xor2  gate1051(.a(G1271), .b(G1270), .O(gate504inter0));
  nand2 gate1052(.a(gate504inter0), .b(s_72), .O(gate504inter1));
  and2  gate1053(.a(G1271), .b(G1270), .O(gate504inter2));
  inv1  gate1054(.a(s_72), .O(gate504inter3));
  inv1  gate1055(.a(s_73), .O(gate504inter4));
  nand2 gate1056(.a(gate504inter4), .b(gate504inter3), .O(gate504inter5));
  nor2  gate1057(.a(gate504inter5), .b(gate504inter2), .O(gate504inter6));
  inv1  gate1058(.a(G1270), .O(gate504inter7));
  inv1  gate1059(.a(G1271), .O(gate504inter8));
  nand2 gate1060(.a(gate504inter8), .b(gate504inter7), .O(gate504inter9));
  nand2 gate1061(.a(s_73), .b(gate504inter3), .O(gate504inter10));
  nor2  gate1062(.a(gate504inter10), .b(gate504inter9), .O(gate504inter11));
  nor2  gate1063(.a(gate504inter11), .b(gate504inter6), .O(gate504inter12));
  nand2 gate1064(.a(gate504inter12), .b(gate504inter1), .O(G1313));
nand2 gate505( .a(G1272), .b(G1273), .O(G1314) );
nand2 gate506( .a(G1274), .b(G1275), .O(G1315) );
nand2 gate507( .a(G1276), .b(G1277), .O(G1316) );
nand2 gate508( .a(G1278), .b(G1279), .O(G1317) );
nand2 gate509( .a(G1280), .b(G1281), .O(G1318) );

  xor2  gate1247(.a(G1283), .b(G1282), .O(gate510inter0));
  nand2 gate1248(.a(gate510inter0), .b(s_100), .O(gate510inter1));
  and2  gate1249(.a(G1283), .b(G1282), .O(gate510inter2));
  inv1  gate1250(.a(s_100), .O(gate510inter3));
  inv1  gate1251(.a(s_101), .O(gate510inter4));
  nand2 gate1252(.a(gate510inter4), .b(gate510inter3), .O(gate510inter5));
  nor2  gate1253(.a(gate510inter5), .b(gate510inter2), .O(gate510inter6));
  inv1  gate1254(.a(G1282), .O(gate510inter7));
  inv1  gate1255(.a(G1283), .O(gate510inter8));
  nand2 gate1256(.a(gate510inter8), .b(gate510inter7), .O(gate510inter9));
  nand2 gate1257(.a(s_101), .b(gate510inter3), .O(gate510inter10));
  nor2  gate1258(.a(gate510inter10), .b(gate510inter9), .O(gate510inter11));
  nor2  gate1259(.a(gate510inter11), .b(gate510inter6), .O(gate510inter12));
  nand2 gate1260(.a(gate510inter12), .b(gate510inter1), .O(G1319));
nand2 gate511( .a(G1284), .b(G1285), .O(G1320) );
nand2 gate512( .a(G1286), .b(G1287), .O(G1321) );
nand2 gate513( .a(G1288), .b(G1289), .O(G1322) );
nand2 gate514( .a(G1290), .b(G1291), .O(G1323) );
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule