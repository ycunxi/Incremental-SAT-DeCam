module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);

input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;//RE__PI;

input s_0,s_1;//RE__ALLOW(00,01,10,11);
input s_2,s_3;//RE__ALLOW(00,01,10,11);
input s_4,s_5;//RE__ALLOW(00,01,10,11);
input s_6,s_7;//RE__ALLOW(00,01,10,11);
input s_8,s_9;//RE__ALLOW(00,01,10,11);
input s_10,s_11;//RE__ALLOW(00,01,10,11);
input s_12,s_13;//RE__ALLOW(00,01,10,11);
input s_14,s_15;//RE__ALLOW(00,01,10,11);
input s_16,s_17;//RE__ALLOW(00,01,10,11);
input s_18,s_19;//RE__ALLOW(00,01,10,11);
input s_20,s_21;//RE__ALLOW(00,01,10,11);
input s_22,s_23;//RE__ALLOW(00,01,10,11);
input s_24,s_25;//RE__ALLOW(00,01,10,11);
input s_26,s_27;//RE__ALLOW(00,01,10,11);
input s_28,s_29;//RE__ALLOW(00,01,10,11);
input s_30,s_31;//RE__ALLOW(00,01,10,11);
input s_32,s_33;//RE__ALLOW(00,01,10,11);
input s_34,s_35;//RE__ALLOW(00,01,10,11);
input s_36,s_37;//RE__ALLOW(00,01,10,11);
input s_38,s_39;//RE__ALLOW(00,01,10,11);
input s_40,s_41;//RE__ALLOW(00,01,10,11);
input s_42,s_43;//RE__ALLOW(00,01,10,11);
input s_44,s_45;//RE__ALLOW(00,01,10,11);
input s_46,s_47;//RE__ALLOW(00,01,10,11);
input s_48,s_49;//RE__ALLOW(00,01,10,11);
input s_50,s_51;//RE__ALLOW(00,01,10,11);
input s_52,s_53;//RE__ALLOW(00,01,10,11);
input s_54,s_55;//RE__ALLOW(00,01,10,11);
input s_56,s_57;//RE__ALLOW(00,01,10,11);
input s_58,s_59;//RE__ALLOW(00,01,10,11);
input s_60,s_61;//RE__ALLOW(00,01,10,11);
input s_62,s_63;//RE__ALLOW(00,01,10,11);
input s_64,s_65;//RE__ALLOW(00,01,10,11);
input s_66,s_67;//RE__ALLOW(00,01,10,11);
input s_68,s_69;//RE__ALLOW(00,01,10,11);
input s_70,s_71;//RE__ALLOW(00,01,10,11);
input s_72,s_73;//RE__ALLOW(00,01,10,11);
input s_74,s_75;//RE__ALLOW(00,01,10,11);
input s_76,s_77;//RE__ALLOW(00,01,10,11);
input s_78,s_79;//RE__ALLOW(00,01,10,11);
input s_80,s_81;//RE__ALLOW(00,01,10,11);
input s_82,s_83;//RE__ALLOW(00,01,10,11);
input s_84,s_85;//RE__ALLOW(00,01,10,11);
input s_86,s_87;//RE__ALLOW(00,01,10,11);
input s_88,s_89;//RE__ALLOW(00,01,10,11);
input s_90,s_91;//RE__ALLOW(00,01,10,11);
input s_92,s_93;//RE__ALLOW(00,01,10,11);
input s_94,s_95;//RE__ALLOW(00,01,10,11);
input s_96,s_97;//RE__ALLOW(00,01,10,11);
input s_98,s_99;//RE__ALLOW(00,01,10,11);
input s_100,s_101;//RE__ALLOW(00,01,10,11);
input s_102,s_103;//RE__ALLOW(00,01,10,11);
input s_104,s_105;//RE__ALLOW(00,01,10,11);
input s_106,s_107;//RE__ALLOW(00,01,10,11);
input s_108,s_109;//RE__ALLOW(00,01,10,11);
input s_110,s_111;//RE__ALLOW(00,01,10,11);
input s_112,s_113;//RE__ALLOW(00,01,10,11);
input s_114,s_115;//RE__ALLOW(00,01,10,11);
input s_116,s_117;//RE__ALLOW(00,01,10,11);
input s_118,s_119;//RE__ALLOW(00,01,10,11);
input s_120,s_121;//RE__ALLOW(00,01,10,11);
input s_122,s_123;//RE__ALLOW(00,01,10,11);
input s_124,s_125;//RE__ALLOW(00,01,10,11);
input s_126,s_127;//RE__ALLOW(00,01,10,11);
input s_128,s_129;//RE__ALLOW(00,01,10,11);
input s_130,s_131;//RE__ALLOW(00,01,10,11);
input s_132,s_133;//RE__ALLOW(00,01,10,11);
input s_134,s_135;//RE__ALLOW(00,01,10,11);
input s_136,s_137;//RE__ALLOW(00,01,10,11);
input s_138,s_139;//RE__ALLOW(00,01,10,11);
input s_140,s_141;//RE__ALLOW(00,01,10,11);
input s_142,s_143;//RE__ALLOW(00,01,10,11);
input s_144,s_145;//RE__ALLOW(00,01,10,11);
input s_146,s_147;//RE__ALLOW(00,01,10,11);
input s_148,s_149;//RE__ALLOW(00,01,10,11);
input s_150,s_151;//RE__ALLOW(00,01,10,11);
input s_152,s_153;//RE__ALLOW(00,01,10,11);
input s_154,s_155;//RE__ALLOW(00,01,10,11);
input s_156,s_157;//RE__ALLOW(00,01,10,11);
input s_158,s_159;//RE__ALLOW(00,01,10,11);
input s_160,s_161;//RE__ALLOW(00,01,10,11);
input s_162,s_163;//RE__ALLOW(00,01,10,11);
input s_164,s_165;//RE__ALLOW(00,01,10,11);
input s_166,s_167;//RE__ALLOW(00,01,10,11);
input s_168,s_169;//RE__ALLOW(00,01,10,11);
input s_170,s_171;//RE__ALLOW(00,01,10,11);
input s_172,s_173;//RE__ALLOW(00,01,10,11);
input s_174,s_175;//RE__ALLOW(00,01,10,11);
input s_176,s_177;//RE__ALLOW(00,01,10,11);
input s_178,s_179;//RE__ALLOW(00,01,10,11);
input s_180,s_181;//RE__ALLOW(00,01,10,11);
input s_182,s_183;//RE__ALLOW(00,01,10,11);
input s_184,s_185;//RE__ALLOW(00,01,10,11);
input s_186,s_187;//RE__ALLOW(00,01,10,11);
input s_188,s_189;//RE__ALLOW(00,01,10,11);
input s_190,s_191;//RE__ALLOW(00,01,10,11);
input s_192,s_193;//RE__ALLOW(00,01,10,11);
input s_194,s_195;//RE__ALLOW(00,01,10,11);
input s_196,s_197;//RE__ALLOW(00,01,10,11);
input s_198,s_199;//RE__ALLOW(00,01,10,11);
input s_200,s_201;//RE__ALLOW(00,01,10,11);
input s_202,s_203;//RE__ALLOW(00,01,10,11);
input s_204,s_205;//RE__ALLOW(00,01,10,11);
input s_206,s_207;//RE__ALLOW(00,01,10,11);
input s_208,s_209;//RE__ALLOW(00,01,10,11);
input s_210,s_211;//RE__ALLOW(00,01,10,11);
input s_212,s_213;//RE__ALLOW(00,01,10,11);
input s_214,s_215;//RE__ALLOW(00,01,10,11);
input s_216,s_217;//RE__ALLOW(00,01,10,11);
input s_218,s_219;//RE__ALLOW(00,01,10,11);
input s_220,s_221;//RE__ALLOW(00,01,10,11);
input s_222,s_223;//RE__ALLOW(00,01,10,11);
input s_224,s_225;//RE__ALLOW(00,01,10,11);
input s_226,s_227;//RE__ALLOW(00,01,10,11);
input s_228,s_229;//RE__ALLOW(00,01,10,11);
input s_230,s_231;//RE__ALLOW(00,01,10,11);
input s_232,s_233;//RE__ALLOW(00,01,10,11);
input s_234,s_235;//RE__ALLOW(00,01,10,11);
input s_236,s_237;//RE__ALLOW(00,01,10,11);
input s_238,s_239;//RE__ALLOW(00,01,10,11);
input s_240,s_241;//RE__ALLOW(00,01,10,11);
input s_242,s_243;//RE__ALLOW(00,01,10,11);
input s_244,s_245;//RE__ALLOW(00,01,10,11);
input s_246,s_247;//RE__ALLOW(00,01,10,11);
input s_248,s_249;//RE__ALLOW(00,01,10,11);
input s_250,s_251;//RE__ALLOW(00,01,10,11);
input s_252,s_253;//RE__ALLOW(00,01,10,11);
input s_254,s_255;//RE__ALLOW(00,01,10,11);
input s_256,s_257;//RE__ALLOW(00,01,10,11);
input s_258,s_259;//RE__ALLOW(00,01,10,11);
input s_260,s_261;//RE__ALLOW(00,01,10,11);
input s_262,s_263;//RE__ALLOW(00,01,10,11);
input s_264,s_265;//RE__ALLOW(00,01,10,11);
input s_266,s_267;//RE__ALLOW(00,01,10,11);
input s_268,s_269;//RE__ALLOW(00,01,10,11);
input s_270,s_271;//RE__ALLOW(00,01,10,11);
input s_272,s_273;//RE__ALLOW(00,01,10,11);
input s_274,s_275;//RE__ALLOW(00,01,10,11);
input s_276,s_277;//RE__ALLOW(00,01,10,11);
input s_278,s_279;//RE__ALLOW(00,01,10,11);
input s_280,s_281;//RE__ALLOW(00,01,10,11);
input s_282,s_283;//RE__ALLOW(00,01,10,11);
input s_284,s_285;//RE__ALLOW(00,01,10,11);
input s_286,s_287;//RE__ALLOW(00,01,10,11);
input s_288,s_289;//RE__ALLOW(00,01,10,11);
input s_290,s_291;//RE__ALLOW(00,01,10,11);
input s_292,s_293;//RE__ALLOW(00,01,10,11);
input s_294,s_295;//RE__ALLOW(00,01,10,11);
input s_296,s_297;//RE__ALLOW(00,01,10,11);
input s_298,s_299;//RE__ALLOW(00,01,10,11);
input s_300,s_301;//RE__ALLOW(00,01,10,11);
input s_302,s_303;//RE__ALLOW(00,01,10,11);
input s_304,s_305;//RE__ALLOW(00,01,10,11);
input s_306,s_307;//RE__ALLOW(00,01,10,11);
input s_308,s_309;//RE__ALLOW(00,01,10,11);
input s_310,s_311;//RE__ALLOW(00,01,10,11);
input s_312,s_313;//RE__ALLOW(00,01,10,11);
input s_314,s_315;//RE__ALLOW(00,01,10,11);
input s_316,s_317;//RE__ALLOW(00,01,10,11);
input s_318,s_319;//RE__ALLOW(00,01,10,11);
input s_320,s_321;//RE__ALLOW(00,01,10,11);
input s_322,s_323;//RE__ALLOW(00,01,10,11);
input s_324,s_325;//RE__ALLOW(00,01,10,11);
input s_326,s_327;//RE__ALLOW(00,01,10,11);
input s_328,s_329;//RE__ALLOW(00,01,10,11);
input s_330,s_331;//RE__ALLOW(00,01,10,11);
input s_332,s_333;//RE__ALLOW(00,01,10,11);
input s_334,s_335;//RE__ALLOW(00,01,10,11);
input s_336,s_337;//RE__ALLOW(00,01,10,11);
input s_338,s_339;//RE__ALLOW(00,01,10,11);
input s_340,s_341;//RE__ALLOW(00,01,10,11);
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;

  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate196inter0, gate196inter1, gate196inter2, gate196inter3, gate196inter4, gate196inter5, gate196inter6, gate196inter7, gate196inter8, gate196inter9, gate196inter10, gate196inter11, gate196inter12, gate459inter0, gate459inter1, gate459inter2, gate459inter3, gate459inter4, gate459inter5, gate459inter6, gate459inter7, gate459inter8, gate459inter9, gate459inter10, gate459inter11, gate459inter12, gate489inter0, gate489inter1, gate489inter2, gate489inter3, gate489inter4, gate489inter5, gate489inter6, gate489inter7, gate489inter8, gate489inter9, gate489inter10, gate489inter11, gate489inter12, gate508inter0, gate508inter1, gate508inter2, gate508inter3, gate508inter4, gate508inter5, gate508inter6, gate508inter7, gate508inter8, gate508inter9, gate508inter10, gate508inter11, gate508inter12, gate234inter0, gate234inter1, gate234inter2, gate234inter3, gate234inter4, gate234inter5, gate234inter6, gate234inter7, gate234inter8, gate234inter9, gate234inter10, gate234inter11, gate234inter12, gate22inter0, gate22inter1, gate22inter2, gate22inter3, gate22inter4, gate22inter5, gate22inter6, gate22inter7, gate22inter8, gate22inter9, gate22inter10, gate22inter11, gate22inter12, gate510inter0, gate510inter1, gate510inter2, gate510inter3, gate510inter4, gate510inter5, gate510inter6, gate510inter7, gate510inter8, gate510inter9, gate510inter10, gate510inter11, gate510inter12, gate50inter0, gate50inter1, gate50inter2, gate50inter3, gate50inter4, gate50inter5, gate50inter6, gate50inter7, gate50inter8, gate50inter9, gate50inter10, gate50inter11, gate50inter12, gate486inter0, gate486inter1, gate486inter2, gate486inter3, gate486inter4, gate486inter5, gate486inter6, gate486inter7, gate486inter8, gate486inter9, gate486inter10, gate486inter11, gate486inter12, gate187inter0, gate187inter1, gate187inter2, gate187inter3, gate187inter4, gate187inter5, gate187inter6, gate187inter7, gate187inter8, gate187inter9, gate187inter10, gate187inter11, gate187inter12, gate266inter0, gate266inter1, gate266inter2, gate266inter3, gate266inter4, gate266inter5, gate266inter6, gate266inter7, gate266inter8, gate266inter9, gate266inter10, gate266inter11, gate266inter12, gate13inter0, gate13inter1, gate13inter2, gate13inter3, gate13inter4, gate13inter5, gate13inter6, gate13inter7, gate13inter8, gate13inter9, gate13inter10, gate13inter11, gate13inter12, gate282inter0, gate282inter1, gate282inter2, gate282inter3, gate282inter4, gate282inter5, gate282inter6, gate282inter7, gate282inter8, gate282inter9, gate282inter10, gate282inter11, gate282inter12, gate33inter0, gate33inter1, gate33inter2, gate33inter3, gate33inter4, gate33inter5, gate33inter6, gate33inter7, gate33inter8, gate33inter9, gate33inter10, gate33inter11, gate33inter12, gate506inter0, gate506inter1, gate506inter2, gate506inter3, gate506inter4, gate506inter5, gate506inter6, gate506inter7, gate506inter8, gate506inter9, gate506inter10, gate506inter11, gate506inter12, gate208inter0, gate208inter1, gate208inter2, gate208inter3, gate208inter4, gate208inter5, gate208inter6, gate208inter7, gate208inter8, gate208inter9, gate208inter10, gate208inter11, gate208inter12, gate290inter0, gate290inter1, gate290inter2, gate290inter3, gate290inter4, gate290inter5, gate290inter6, gate290inter7, gate290inter8, gate290inter9, gate290inter10, gate290inter11, gate290inter12, gate205inter0, gate205inter1, gate205inter2, gate205inter3, gate205inter4, gate205inter5, gate205inter6, gate205inter7, gate205inter8, gate205inter9, gate205inter10, gate205inter11, gate205inter12, gate285inter0, gate285inter1, gate285inter2, gate285inter3, gate285inter4, gate285inter5, gate285inter6, gate285inter7, gate285inter8, gate285inter9, gate285inter10, gate285inter11, gate285inter12, gate228inter0, gate228inter1, gate228inter2, gate228inter3, gate228inter4, gate228inter5, gate228inter6, gate228inter7, gate228inter8, gate228inter9, gate228inter10, gate228inter11, gate228inter12, gate243inter0, gate243inter1, gate243inter2, gate243inter3, gate243inter4, gate243inter5, gate243inter6, gate243inter7, gate243inter8, gate243inter9, gate243inter10, gate243inter11, gate243inter12, gate51inter0, gate51inter1, gate51inter2, gate51inter3, gate51inter4, gate51inter5, gate51inter6, gate51inter7, gate51inter8, gate51inter9, gate51inter10, gate51inter11, gate51inter12, gate477inter0, gate477inter1, gate477inter2, gate477inter3, gate477inter4, gate477inter5, gate477inter6, gate477inter7, gate477inter8, gate477inter9, gate477inter10, gate477inter11, gate477inter12, gate262inter0, gate262inter1, gate262inter2, gate262inter3, gate262inter4, gate262inter5, gate262inter6, gate262inter7, gate262inter8, gate262inter9, gate262inter10, gate262inter11, gate262inter12, gate256inter0, gate256inter1, gate256inter2, gate256inter3, gate256inter4, gate256inter5, gate256inter6, gate256inter7, gate256inter8, gate256inter9, gate256inter10, gate256inter11, gate256inter12, gate391inter0, gate391inter1, gate391inter2, gate391inter3, gate391inter4, gate391inter5, gate391inter6, gate391inter7, gate391inter8, gate391inter9, gate391inter10, gate391inter11, gate391inter12, gate431inter0, gate431inter1, gate431inter2, gate431inter3, gate431inter4, gate431inter5, gate431inter6, gate431inter7, gate431inter8, gate431inter9, gate431inter10, gate431inter11, gate431inter12, gate483inter0, gate483inter1, gate483inter2, gate483inter3, gate483inter4, gate483inter5, gate483inter6, gate483inter7, gate483inter8, gate483inter9, gate483inter10, gate483inter11, gate483inter12, gate21inter0, gate21inter1, gate21inter2, gate21inter3, gate21inter4, gate21inter5, gate21inter6, gate21inter7, gate21inter8, gate21inter9, gate21inter10, gate21inter11, gate21inter12, gate429inter0, gate429inter1, gate429inter2, gate429inter3, gate429inter4, gate429inter5, gate429inter6, gate429inter7, gate429inter8, gate429inter9, gate429inter10, gate429inter11, gate429inter12, gate191inter0, gate191inter1, gate191inter2, gate191inter3, gate191inter4, gate191inter5, gate191inter6, gate191inter7, gate191inter8, gate191inter9, gate191inter10, gate191inter11, gate191inter12, gate60inter0, gate60inter1, gate60inter2, gate60inter3, gate60inter4, gate60inter5, gate60inter6, gate60inter7, gate60inter8, gate60inter9, gate60inter10, gate60inter11, gate60inter12, gate455inter0, gate455inter1, gate455inter2, gate455inter3, gate455inter4, gate455inter5, gate455inter6, gate455inter7, gate455inter8, gate455inter9, gate455inter10, gate455inter11, gate455inter12, gate231inter0, gate231inter1, gate231inter2, gate231inter3, gate231inter4, gate231inter5, gate231inter6, gate231inter7, gate231inter8, gate231inter9, gate231inter10, gate231inter11, gate231inter12, gate35inter0, gate35inter1, gate35inter2, gate35inter3, gate35inter4, gate35inter5, gate35inter6, gate35inter7, gate35inter8, gate35inter9, gate35inter10, gate35inter11, gate35inter12, gate467inter0, gate467inter1, gate467inter2, gate467inter3, gate467inter4, gate467inter5, gate467inter6, gate467inter7, gate467inter8, gate467inter9, gate467inter10, gate467inter11, gate467inter12, gate47inter0, gate47inter1, gate47inter2, gate47inter3, gate47inter4, gate47inter5, gate47inter6, gate47inter7, gate47inter8, gate47inter9, gate47inter10, gate47inter11, gate47inter12, gate87inter0, gate87inter1, gate87inter2, gate87inter3, gate87inter4, gate87inter5, gate87inter6, gate87inter7, gate87inter8, gate87inter9, gate87inter10, gate87inter11, gate87inter12, gate250inter0, gate250inter1, gate250inter2, gate250inter3, gate250inter4, gate250inter5, gate250inter6, gate250inter7, gate250inter8, gate250inter9, gate250inter10, gate250inter11, gate250inter12, gate147inter0, gate147inter1, gate147inter2, gate147inter3, gate147inter4, gate147inter5, gate147inter6, gate147inter7, gate147inter8, gate147inter9, gate147inter10, gate147inter11, gate147inter12, gate203inter0, gate203inter1, gate203inter2, gate203inter3, gate203inter4, gate203inter5, gate203inter6, gate203inter7, gate203inter8, gate203inter9, gate203inter10, gate203inter11, gate203inter12, gate245inter0, gate245inter1, gate245inter2, gate245inter3, gate245inter4, gate245inter5, gate245inter6, gate245inter7, gate245inter8, gate245inter9, gate245inter10, gate245inter11, gate245inter12, gate103inter0, gate103inter1, gate103inter2, gate103inter3, gate103inter4, gate103inter5, gate103inter6, gate103inter7, gate103inter8, gate103inter9, gate103inter10, gate103inter11, gate103inter12, gate283inter0, gate283inter1, gate283inter2, gate283inter3, gate283inter4, gate283inter5, gate283inter6, gate283inter7, gate283inter8, gate283inter9, gate283inter10, gate283inter11, gate283inter12, gate140inter0, gate140inter1, gate140inter2, gate140inter3, gate140inter4, gate140inter5, gate140inter6, gate140inter7, gate140inter8, gate140inter9, gate140inter10, gate140inter11, gate140inter12, gate421inter0, gate421inter1, gate421inter2, gate421inter3, gate421inter4, gate421inter5, gate421inter6, gate421inter7, gate421inter8, gate421inter9, gate421inter10, gate421inter11, gate421inter12, gate148inter0, gate148inter1, gate148inter2, gate148inter3, gate148inter4, gate148inter5, gate148inter6, gate148inter7, gate148inter8, gate148inter9, gate148inter10, gate148inter11, gate148inter12, gate288inter0, gate288inter1, gate288inter2, gate288inter3, gate288inter4, gate288inter5, gate288inter6, gate288inter7, gate288inter8, gate288inter9, gate288inter10, gate288inter11, gate288inter12, gate452inter0, gate452inter1, gate452inter2, gate452inter3, gate452inter4, gate452inter5, gate452inter6, gate452inter7, gate452inter8, gate452inter9, gate452inter10, gate452inter11, gate452inter12, gate10inter0, gate10inter1, gate10inter2, gate10inter3, gate10inter4, gate10inter5, gate10inter6, gate10inter7, gate10inter8, gate10inter9, gate10inter10, gate10inter11, gate10inter12, gate418inter0, gate418inter1, gate418inter2, gate418inter3, gate418inter4, gate418inter5, gate418inter6, gate418inter7, gate418inter8, gate418inter9, gate418inter10, gate418inter11, gate418inter12, gate159inter0, gate159inter1, gate159inter2, gate159inter3, gate159inter4, gate159inter5, gate159inter6, gate159inter7, gate159inter8, gate159inter9, gate159inter10, gate159inter11, gate159inter12, gate441inter0, gate441inter1, gate441inter2, gate441inter3, gate441inter4, gate441inter5, gate441inter6, gate441inter7, gate441inter8, gate441inter9, gate441inter10, gate441inter11, gate441inter12, gate169inter0, gate169inter1, gate169inter2, gate169inter3, gate169inter4, gate169inter5, gate169inter6, gate169inter7, gate169inter8, gate169inter9, gate169inter10, gate169inter11, gate169inter12, gate168inter0, gate168inter1, gate168inter2, gate168inter3, gate168inter4, gate168inter5, gate168inter6, gate168inter7, gate168inter8, gate168inter9, gate168inter10, gate168inter11, gate168inter12, gate163inter0, gate163inter1, gate163inter2, gate163inter3, gate163inter4, gate163inter5, gate163inter6, gate163inter7, gate163inter8, gate163inter9, gate163inter10, gate163inter11, gate163inter12, gate487inter0, gate487inter1, gate487inter2, gate487inter3, gate487inter4, gate487inter5, gate487inter6, gate487inter7, gate487inter8, gate487inter9, gate487inter10, gate487inter11, gate487inter12, gate458inter0, gate458inter1, gate458inter2, gate458inter3, gate458inter4, gate458inter5, gate458inter6, gate458inter7, gate458inter8, gate458inter9, gate458inter10, gate458inter11, gate458inter12, gate197inter0, gate197inter1, gate197inter2, gate197inter3, gate197inter4, gate197inter5, gate197inter6, gate197inter7, gate197inter8, gate197inter9, gate197inter10, gate197inter11, gate197inter12, gate198inter0, gate198inter1, gate198inter2, gate198inter3, gate198inter4, gate198inter5, gate198inter6, gate198inter7, gate198inter8, gate198inter9, gate198inter10, gate198inter11, gate198inter12, gate117inter0, gate117inter1, gate117inter2, gate117inter3, gate117inter4, gate117inter5, gate117inter6, gate117inter7, gate117inter8, gate117inter9, gate117inter10, gate117inter11, gate117inter12, gate265inter0, gate265inter1, gate265inter2, gate265inter3, gate265inter4, gate265inter5, gate265inter6, gate265inter7, gate265inter8, gate265inter9, gate265inter10, gate265inter11, gate265inter12, gate223inter0, gate223inter1, gate223inter2, gate223inter3, gate223inter4, gate223inter5, gate223inter6, gate223inter7, gate223inter8, gate223inter9, gate223inter10, gate223inter11, gate223inter12, gate460inter0, gate460inter1, gate460inter2, gate460inter3, gate460inter4, gate460inter5, gate460inter6, gate460inter7, gate460inter8, gate460inter9, gate460inter10, gate460inter11, gate460inter12, gate174inter0, gate174inter1, gate174inter2, gate174inter3, gate174inter4, gate174inter5, gate174inter6, gate174inter7, gate174inter8, gate174inter9, gate174inter10, gate174inter11, gate174inter12, gate58inter0, gate58inter1, gate58inter2, gate58inter3, gate58inter4, gate58inter5, gate58inter6, gate58inter7, gate58inter8, gate58inter9, gate58inter10, gate58inter11, gate58inter12, gate456inter0, gate456inter1, gate456inter2, gate456inter3, gate456inter4, gate456inter5, gate456inter6, gate456inter7, gate456inter8, gate456inter9, gate456inter10, gate456inter11, gate456inter12, gate402inter0, gate402inter1, gate402inter2, gate402inter3, gate402inter4, gate402inter5, gate402inter6, gate402inter7, gate402inter8, gate402inter9, gate402inter10, gate402inter11, gate402inter12, gate408inter0, gate408inter1, gate408inter2, gate408inter3, gate408inter4, gate408inter5, gate408inter6, gate408inter7, gate408inter8, gate408inter9, gate408inter10, gate408inter11, gate408inter12, gate31inter0, gate31inter1, gate31inter2, gate31inter3, gate31inter4, gate31inter5, gate31inter6, gate31inter7, gate31inter8, gate31inter9, gate31inter10, gate31inter11, gate31inter12, gate188inter0, gate188inter1, gate188inter2, gate188inter3, gate188inter4, gate188inter5, gate188inter6, gate188inter7, gate188inter8, gate188inter9, gate188inter10, gate188inter11, gate188inter12, gate412inter0, gate412inter1, gate412inter2, gate412inter3, gate412inter4, gate412inter5, gate412inter6, gate412inter7, gate412inter8, gate412inter9, gate412inter10, gate412inter11, gate412inter12, gate445inter0, gate445inter1, gate445inter2, gate445inter3, gate445inter4, gate445inter5, gate445inter6, gate445inter7, gate445inter8, gate445inter9, gate445inter10, gate445inter11, gate445inter12, gate118inter0, gate118inter1, gate118inter2, gate118inter3, gate118inter4, gate118inter5, gate118inter6, gate118inter7, gate118inter8, gate118inter9, gate118inter10, gate118inter11, gate118inter12, gate430inter0, gate430inter1, gate430inter2, gate430inter3, gate430inter4, gate430inter5, gate430inter6, gate430inter7, gate430inter8, gate430inter9, gate430inter10, gate430inter11, gate430inter12, gate48inter0, gate48inter1, gate48inter2, gate48inter3, gate48inter4, gate48inter5, gate48inter6, gate48inter7, gate48inter8, gate48inter9, gate48inter10, gate48inter11, gate48inter12, gate137inter0, gate137inter1, gate137inter2, gate137inter3, gate137inter4, gate137inter5, gate137inter6, gate137inter7, gate137inter8, gate137inter9, gate137inter10, gate137inter11, gate137inter12, gate417inter0, gate417inter1, gate417inter2, gate417inter3, gate417inter4, gate417inter5, gate417inter6, gate417inter7, gate417inter8, gate417inter9, gate417inter10, gate417inter11, gate417inter12, gate183inter0, gate183inter1, gate183inter2, gate183inter3, gate183inter4, gate183inter5, gate183inter6, gate183inter7, gate183inter8, gate183inter9, gate183inter10, gate183inter11, gate183inter12, gate400inter0, gate400inter1, gate400inter2, gate400inter3, gate400inter4, gate400inter5, gate400inter6, gate400inter7, gate400inter8, gate400inter9, gate400inter10, gate400inter11, gate400inter12, gate143inter0, gate143inter1, gate143inter2, gate143inter3, gate143inter4, gate143inter5, gate143inter6, gate143inter7, gate143inter8, gate143inter9, gate143inter10, gate143inter11, gate143inter12, gate406inter0, gate406inter1, gate406inter2, gate406inter3, gate406inter4, gate406inter5, gate406inter6, gate406inter7, gate406inter8, gate406inter9, gate406inter10, gate406inter11, gate406inter12, gate185inter0, gate185inter1, gate185inter2, gate185inter3, gate185inter4, gate185inter5, gate185inter6, gate185inter7, gate185inter8, gate185inter9, gate185inter10, gate185inter11, gate185inter12, gate99inter0, gate99inter1, gate99inter2, gate99inter3, gate99inter4, gate99inter5, gate99inter6, gate99inter7, gate99inter8, gate99inter9, gate99inter10, gate99inter11, gate99inter12, gate128inter0, gate128inter1, gate128inter2, gate128inter3, gate128inter4, gate128inter5, gate128inter6, gate128inter7, gate128inter8, gate128inter9, gate128inter10, gate128inter11, gate128inter12, gate113inter0, gate113inter1, gate113inter2, gate113inter3, gate113inter4, gate113inter5, gate113inter6, gate113inter7, gate113inter8, gate113inter9, gate113inter10, gate113inter11, gate113inter12, gate162inter0, gate162inter1, gate162inter2, gate162inter3, gate162inter4, gate162inter5, gate162inter6, gate162inter7, gate162inter8, gate162inter9, gate162inter10, gate162inter11, gate162inter12, gate270inter0, gate270inter1, gate270inter2, gate270inter3, gate270inter4, gate270inter5, gate270inter6, gate270inter7, gate270inter8, gate270inter9, gate270inter10, gate270inter11, gate270inter12, gate182inter0, gate182inter1, gate182inter2, gate182inter3, gate182inter4, gate182inter5, gate182inter6, gate182inter7, gate182inter8, gate182inter9, gate182inter10, gate182inter11, gate182inter12, gate201inter0, gate201inter1, gate201inter2, gate201inter3, gate201inter4, gate201inter5, gate201inter6, gate201inter7, gate201inter8, gate201inter9, gate201inter10, gate201inter11, gate201inter12, gate286inter0, gate286inter1, gate286inter2, gate286inter3, gate286inter4, gate286inter5, gate286inter6, gate286inter7, gate286inter8, gate286inter9, gate286inter10, gate286inter11, gate286inter12, gate123inter0, gate123inter1, gate123inter2, gate123inter3, gate123inter4, gate123inter5, gate123inter6, gate123inter7, gate123inter8, gate123inter9, gate123inter10, gate123inter11, gate123inter12, gate279inter0, gate279inter1, gate279inter2, gate279inter3, gate279inter4, gate279inter5, gate279inter6, gate279inter7, gate279inter8, gate279inter9, gate279inter10, gate279inter11, gate279inter12, gate504inter0, gate504inter1, gate504inter2, gate504inter3, gate504inter4, gate504inter5, gate504inter6, gate504inter7, gate504inter8, gate504inter9, gate504inter10, gate504inter11, gate504inter12, gate253inter0, gate253inter1, gate253inter2, gate253inter3, gate253inter4, gate253inter5, gate253inter6, gate253inter7, gate253inter8, gate253inter9, gate253inter10, gate253inter11, gate253inter12, gate155inter0, gate155inter1, gate155inter2, gate155inter3, gate155inter4, gate155inter5, gate155inter6, gate155inter7, gate155inter8, gate155inter9, gate155inter10, gate155inter11, gate155inter12, gate259inter0, gate259inter1, gate259inter2, gate259inter3, gate259inter4, gate259inter5, gate259inter6, gate259inter7, gate259inter8, gate259inter9, gate259inter10, gate259inter11, gate259inter12, gate134inter0, gate134inter1, gate134inter2, gate134inter3, gate134inter4, gate134inter5, gate134inter6, gate134inter7, gate134inter8, gate134inter9, gate134inter10, gate134inter11, gate134inter12, gate263inter0, gate263inter1, gate263inter2, gate263inter3, gate263inter4, gate263inter5, gate263inter6, gate263inter7, gate263inter8, gate263inter9, gate263inter10, gate263inter11, gate263inter12, gate65inter0, gate65inter1, gate65inter2, gate65inter3, gate65inter4, gate65inter5, gate65inter6, gate65inter7, gate65inter8, gate65inter9, gate65inter10, gate65inter11, gate65inter12, gate77inter0, gate77inter1, gate77inter2, gate77inter3, gate77inter4, gate77inter5, gate77inter6, gate77inter7, gate77inter8, gate77inter9, gate77inter10, gate77inter11, gate77inter12, gate42inter0, gate42inter1, gate42inter2, gate42inter3, gate42inter4, gate42inter5, gate42inter6, gate42inter7, gate42inter8, gate42inter9, gate42inter10, gate42inter11, gate42inter12, gate23inter0, gate23inter1, gate23inter2, gate23inter3, gate23inter4, gate23inter5, gate23inter6, gate23inter7, gate23inter8, gate23inter9, gate23inter10, gate23inter11, gate23inter12, gate229inter0, gate229inter1, gate229inter2, gate229inter3, gate229inter4, gate229inter5, gate229inter6, gate229inter7, gate229inter8, gate229inter9, gate229inter10, gate229inter11, gate229inter12, gate254inter0, gate254inter1, gate254inter2, gate254inter3, gate254inter4, gate254inter5, gate254inter6, gate254inter7, gate254inter8, gate254inter9, gate254inter10, gate254inter11, gate254inter12, gate179inter0, gate179inter1, gate179inter2, gate179inter3, gate179inter4, gate179inter5, gate179inter6, gate179inter7, gate179inter8, gate179inter9, gate179inter10, gate179inter11, gate179inter12, gate449inter0, gate449inter1, gate449inter2, gate449inter3, gate449inter4, gate449inter5, gate449inter6, gate449inter7, gate449inter8, gate449inter9, gate449inter10, gate449inter11, gate449inter12, gate443inter0, gate443inter1, gate443inter2, gate443inter3, gate443inter4, gate443inter5, gate443inter6, gate443inter7, gate443inter8, gate443inter9, gate443inter10, gate443inter11, gate443inter12, gate45inter0, gate45inter1, gate45inter2, gate45inter3, gate45inter4, gate45inter5, gate45inter6, gate45inter7, gate45inter8, gate45inter9, gate45inter10, gate45inter11, gate45inter12, gate20inter0, gate20inter1, gate20inter2, gate20inter3, gate20inter4, gate20inter5, gate20inter6, gate20inter7, gate20inter8, gate20inter9, gate20inter10, gate20inter11, gate20inter12, gate247inter0, gate247inter1, gate247inter2, gate247inter3, gate247inter4, gate247inter5, gate247inter6, gate247inter7, gate247inter8, gate247inter9, gate247inter10, gate247inter11, gate247inter12, gate175inter0, gate175inter1, gate175inter2, gate175inter3, gate175inter4, gate175inter5, gate175inter6, gate175inter7, gate175inter8, gate175inter9, gate175inter10, gate175inter11, gate175inter12, gate255inter0, gate255inter1, gate255inter2, gate255inter3, gate255inter4, gate255inter5, gate255inter6, gate255inter7, gate255inter8, gate255inter9, gate255inter10, gate255inter11, gate255inter12, gate171inter0, gate171inter1, gate171inter2, gate171inter3, gate171inter4, gate171inter5, gate171inter6, gate171inter7, gate171inter8, gate171inter9, gate171inter10, gate171inter11, gate171inter12, gate9inter0, gate9inter1, gate9inter2, gate9inter3, gate9inter4, gate9inter5, gate9inter6, gate9inter7, gate9inter8, gate9inter9, gate9inter10, gate9inter11, gate9inter12, gate496inter0, gate496inter1, gate496inter2, gate496inter3, gate496inter4, gate496inter5, gate496inter6, gate496inter7, gate496inter8, gate496inter9, gate496inter10, gate496inter11, gate496inter12, gate132inter0, gate132inter1, gate132inter2, gate132inter3, gate132inter4, gate132inter5, gate132inter6, gate132inter7, gate132inter8, gate132inter9, gate132inter10, gate132inter11, gate132inter12, gate446inter0, gate446inter1, gate446inter2, gate446inter3, gate446inter4, gate446inter5, gate446inter6, gate446inter7, gate446inter8, gate446inter9, gate446inter10, gate446inter11, gate446inter12, gate435inter0, gate435inter1, gate435inter2, gate435inter3, gate435inter4, gate435inter5, gate435inter6, gate435inter7, gate435inter8, gate435inter9, gate435inter10, gate435inter11, gate435inter12, gate151inter0, gate151inter1, gate151inter2, gate151inter3, gate151inter4, gate151inter5, gate151inter6, gate151inter7, gate151inter8, gate151inter9, gate151inter10, gate151inter11, gate151inter12, gate86inter0, gate86inter1, gate86inter2, gate86inter3, gate86inter4, gate86inter5, gate86inter6, gate86inter7, gate86inter8, gate86inter9, gate86inter10, gate86inter11, gate86inter12, gate27inter0, gate27inter1, gate27inter2, gate27inter3, gate27inter4, gate27inter5, gate27inter6, gate27inter7, gate27inter8, gate27inter9, gate27inter10, gate27inter11, gate27inter12, gate36inter0, gate36inter1, gate36inter2, gate36inter3, gate36inter4, gate36inter5, gate36inter6, gate36inter7, gate36inter8, gate36inter9, gate36inter10, gate36inter11, gate36inter12, gate160inter0, gate160inter1, gate160inter2, gate160inter3, gate160inter4, gate160inter5, gate160inter6, gate160inter7, gate160inter8, gate160inter9, gate160inter10, gate160inter11, gate160inter12, gate136inter0, gate136inter1, gate136inter2, gate136inter3, gate136inter4, gate136inter5, gate136inter6, gate136inter7, gate136inter8, gate136inter9, gate136inter10, gate136inter11, gate136inter12, gate14inter0, gate14inter1, gate14inter2, gate14inter3, gate14inter4, gate14inter5, gate14inter6, gate14inter7, gate14inter8, gate14inter9, gate14inter10, gate14inter11, gate14inter12, gate261inter0, gate261inter1, gate261inter2, gate261inter3, gate261inter4, gate261inter5, gate261inter6, gate261inter7, gate261inter8, gate261inter9, gate261inter10, gate261inter11, gate261inter12, gate44inter0, gate44inter1, gate44inter2, gate44inter3, gate44inter4, gate44inter5, gate44inter6, gate44inter7, gate44inter8, gate44inter9, gate44inter10, gate44inter11, gate44inter12, gate112inter0, gate112inter1, gate112inter2, gate112inter3, gate112inter4, gate112inter5, gate112inter6, gate112inter7, gate112inter8, gate112inter9, gate112inter10, gate112inter11, gate112inter12, gate436inter0, gate436inter1, gate436inter2, gate436inter3, gate436inter4, gate436inter5, gate436inter6, gate436inter7, gate436inter8, gate436inter9, gate436inter10, gate436inter11, gate436inter12, gate17inter0, gate17inter1, gate17inter2, gate17inter3, gate17inter4, gate17inter5, gate17inter6, gate17inter7, gate17inter8, gate17inter9, gate17inter10, gate17inter11, gate17inter12, gate478inter0, gate478inter1, gate478inter2, gate478inter3, gate478inter4, gate478inter5, gate478inter6, gate478inter7, gate478inter8, gate478inter9, gate478inter10, gate478inter11, gate478inter12, gate104inter0, gate104inter1, gate104inter2, gate104inter3, gate104inter4, gate104inter5, gate104inter6, gate104inter7, gate104inter8, gate104inter9, gate104inter10, gate104inter11, gate104inter12, gate173inter0, gate173inter1, gate173inter2, gate173inter3, gate173inter4, gate173inter5, gate173inter6, gate173inter7, gate173inter8, gate173inter9, gate173inter10, gate173inter11, gate173inter12, gate502inter0, gate502inter1, gate502inter2, gate502inter3, gate502inter4, gate502inter5, gate502inter6, gate502inter7, gate502inter8, gate502inter9, gate502inter10, gate502inter11, gate502inter12, gate281inter0, gate281inter1, gate281inter2, gate281inter3, gate281inter4, gate281inter5, gate281inter6, gate281inter7, gate281inter8, gate281inter9, gate281inter10, gate281inter11, gate281inter12, gate235inter0, gate235inter1, gate235inter2, gate235inter3, gate235inter4, gate235inter5, gate235inter6, gate235inter7, gate235inter8, gate235inter9, gate235inter10, gate235inter11, gate235inter12, gate248inter0, gate248inter1, gate248inter2, gate248inter3, gate248inter4, gate248inter5, gate248inter6, gate248inter7, gate248inter8, gate248inter9, gate248inter10, gate248inter11, gate248inter12, gate108inter0, gate108inter1, gate108inter2, gate108inter3, gate108inter4, gate108inter5, gate108inter6, gate108inter7, gate108inter8, gate108inter9, gate108inter10, gate108inter11, gate108inter12, gate457inter0, gate457inter1, gate457inter2, gate457inter3, gate457inter4, gate457inter5, gate457inter6, gate457inter7, gate457inter8, gate457inter9, gate457inter10, gate457inter11, gate457inter12, gate399inter0, gate399inter1, gate399inter2, gate399inter3, gate399inter4, gate399inter5, gate399inter6, gate399inter7, gate399inter8, gate399inter9, gate399inter10, gate399inter11, gate399inter12, gate206inter0, gate206inter1, gate206inter2, gate206inter3, gate206inter4, gate206inter5, gate206inter6, gate206inter7, gate206inter8, gate206inter9, gate206inter10, gate206inter11, gate206inter12, gate41inter0, gate41inter1, gate41inter2, gate41inter3, gate41inter4, gate41inter5, gate41inter6, gate41inter7, gate41inter8, gate41inter9, gate41inter10, gate41inter11, gate41inter12, gate410inter0, gate410inter1, gate410inter2, gate410inter3, gate410inter4, gate410inter5, gate410inter6, gate410inter7, gate410inter8, gate410inter9, gate410inter10, gate410inter11, gate410inter12, gate167inter0, gate167inter1, gate167inter2, gate167inter3, gate167inter4, gate167inter5, gate167inter6, gate167inter7, gate167inter8, gate167inter9, gate167inter10, gate167inter11, gate167inter12, gate387inter0, gate387inter1, gate387inter2, gate387inter3, gate387inter4, gate387inter5, gate387inter6, gate387inter7, gate387inter8, gate387inter9, gate387inter10, gate387inter11, gate387inter12, gate120inter0, gate120inter1, gate120inter2, gate120inter3, gate120inter4, gate120inter5, gate120inter6, gate120inter7, gate120inter8, gate120inter9, gate120inter10, gate120inter11, gate120inter12, gate291inter0, gate291inter1, gate291inter2, gate291inter3, gate291inter4, gate291inter5, gate291inter6, gate291inter7, gate291inter8, gate291inter9, gate291inter10, gate291inter11, gate291inter12, gate122inter0, gate122inter1, gate122inter2, gate122inter3, gate122inter4, gate122inter5, gate122inter6, gate122inter7, gate122inter8, gate122inter9, gate122inter10, gate122inter11, gate122inter12, gate438inter0, gate438inter1, gate438inter2, gate438inter3, gate438inter4, gate438inter5, gate438inter6, gate438inter7, gate438inter8, gate438inter9, gate438inter10, gate438inter11, gate438inter12, gate18inter0, gate18inter1, gate18inter2, gate18inter3, gate18inter4, gate18inter5, gate18inter6, gate18inter7, gate18inter8, gate18inter9, gate18inter10, gate18inter11, gate18inter12, gate209inter0, gate209inter1, gate209inter2, gate209inter3, gate209inter4, gate209inter5, gate209inter6, gate209inter7, gate209inter8, gate209inter9, gate209inter10, gate209inter11, gate209inter12, gate442inter0, gate442inter1, gate442inter2, gate442inter3, gate442inter4, gate442inter5, gate442inter6, gate442inter7, gate442inter8, gate442inter9, gate442inter10, gate442inter11, gate442inter12, gate512inter0, gate512inter1, gate512inter2, gate512inter3, gate512inter4, gate512inter5, gate512inter6, gate512inter7, gate512inter8, gate512inter9, gate512inter10, gate512inter11, gate512inter12, gate125inter0, gate125inter1, gate125inter2, gate125inter3, gate125inter4, gate125inter5, gate125inter6, gate125inter7, gate125inter8, gate125inter9, gate125inter10, gate125inter11, gate125inter12, gate271inter0, gate271inter1, gate271inter2, gate271inter3, gate271inter4, gate271inter5, gate271inter6, gate271inter7, gate271inter8, gate271inter9, gate271inter10, gate271inter11, gate271inter12, gate85inter0, gate85inter1, gate85inter2, gate85inter3, gate85inter4, gate85inter5, gate85inter6, gate85inter7, gate85inter8, gate85inter9, gate85inter10, gate85inter11, gate85inter12, gate415inter0, gate415inter1, gate415inter2, gate415inter3, gate415inter4, gate415inter5, gate415inter6, gate415inter7, gate415inter8, gate415inter9, gate415inter10, gate415inter11, gate415inter12, gate210inter0, gate210inter1, gate210inter2, gate210inter3, gate210inter4, gate210inter5, gate210inter6, gate210inter7, gate210inter8, gate210inter9, gate210inter10, gate210inter11, gate210inter12, gate199inter0, gate199inter1, gate199inter2, gate199inter3, gate199inter4, gate199inter5, gate199inter6, gate199inter7, gate199inter8, gate199inter9, gate199inter10, gate199inter11, gate199inter12, gate32inter0, gate32inter1, gate32inter2, gate32inter3, gate32inter4, gate32inter5, gate32inter6, gate32inter7, gate32inter8, gate32inter9, gate32inter10, gate32inter11, gate32inter12, gate479inter0, gate479inter1, gate479inter2, gate479inter3, gate479inter4, gate479inter5, gate479inter6, gate479inter7, gate479inter8, gate479inter9, gate479inter10, gate479inter11, gate479inter12, gate394inter0, gate394inter1, gate394inter2, gate394inter3, gate394inter4, gate394inter5, gate394inter6, gate394inter7, gate394inter8, gate394inter9, gate394inter10, gate394inter11, gate394inter12, gate181inter0, gate181inter1, gate181inter2, gate181inter3, gate181inter4, gate181inter5, gate181inter6, gate181inter7, gate181inter8, gate181inter9, gate181inter10, gate181inter11, gate181inter12, gate403inter0, gate403inter1, gate403inter2, gate403inter3, gate403inter4, gate403inter5, gate403inter6, gate403inter7, gate403inter8, gate403inter9, gate403inter10, gate403inter11, gate403inter12, gate177inter0, gate177inter1, gate177inter2, gate177inter3, gate177inter4, gate177inter5, gate177inter6, gate177inter7, gate177inter8, gate177inter9, gate177inter10, gate177inter11, gate177inter12, gate434inter0, gate434inter1, gate434inter2, gate434inter3, gate434inter4, gate434inter5, gate434inter6, gate434inter7, gate434inter8, gate434inter9, gate434inter10, gate434inter11, gate434inter12, gate276inter0, gate276inter1, gate276inter2, gate276inter3, gate276inter4, gate276inter5, gate276inter6, gate276inter7, gate276inter8, gate276inter9, gate276inter10, gate276inter11, gate276inter12, gate12inter0, gate12inter1, gate12inter2, gate12inter3, gate12inter4, gate12inter5, gate12inter6, gate12inter7, gate12inter8, gate12inter9, gate12inter10, gate12inter11, gate12inter12, gate268inter0, gate268inter1, gate268inter2, gate268inter3, gate268inter4, gate268inter5, gate268inter6, gate268inter7, gate268inter8, gate268inter9, gate268inter10, gate268inter11, gate268inter12, gate222inter0, gate222inter1, gate222inter2, gate222inter3, gate222inter4, gate222inter5, gate222inter6, gate222inter7, gate222inter8, gate222inter9, gate222inter10, gate222inter11, gate222inter12;



and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );

  xor2  gate2143(.a(G2), .b(G1), .O(gate9inter0));
  nand2 gate2144(.a(gate9inter0), .b(s_228), .O(gate9inter1));
  and2  gate2145(.a(G2), .b(G1), .O(gate9inter2));
  inv1  gate2146(.a(s_228), .O(gate9inter3));
  inv1  gate2147(.a(s_229), .O(gate9inter4));
  nand2 gate2148(.a(gate9inter4), .b(gate9inter3), .O(gate9inter5));
  nor2  gate2149(.a(gate9inter5), .b(gate9inter2), .O(gate9inter6));
  inv1  gate2150(.a(G1), .O(gate9inter7));
  inv1  gate2151(.a(G2), .O(gate9inter8));
  nand2 gate2152(.a(gate9inter8), .b(gate9inter7), .O(gate9inter9));
  nand2 gate2153(.a(s_229), .b(gate9inter3), .O(gate9inter10));
  nor2  gate2154(.a(gate9inter10), .b(gate9inter9), .O(gate9inter11));
  nor2  gate2155(.a(gate9inter11), .b(gate9inter6), .O(gate9inter12));
  nand2 gate2156(.a(gate9inter12), .b(gate9inter1), .O(G266));

  xor2  gate1233(.a(G4), .b(G3), .O(gate10inter0));
  nand2 gate1234(.a(gate10inter0), .b(s_98), .O(gate10inter1));
  and2  gate1235(.a(G4), .b(G3), .O(gate10inter2));
  inv1  gate1236(.a(s_98), .O(gate10inter3));
  inv1  gate1237(.a(s_99), .O(gate10inter4));
  nand2 gate1238(.a(gate10inter4), .b(gate10inter3), .O(gate10inter5));
  nor2  gate1239(.a(gate10inter5), .b(gate10inter2), .O(gate10inter6));
  inv1  gate1240(.a(G3), .O(gate10inter7));
  inv1  gate1241(.a(G4), .O(gate10inter8));
  nand2 gate1242(.a(gate10inter8), .b(gate10inter7), .O(gate10inter9));
  nand2 gate1243(.a(s_99), .b(gate10inter3), .O(gate10inter10));
  nor2  gate1244(.a(gate10inter10), .b(gate10inter9), .O(gate10inter11));
  nor2  gate1245(.a(gate10inter11), .b(gate10inter6), .O(gate10inter12));
  nand2 gate1246(.a(gate10inter12), .b(gate10inter1), .O(G269));
nand2 gate11( .a(G5), .b(G6), .O(G272) );

  xor2  gate2899(.a(G8), .b(G7), .O(gate12inter0));
  nand2 gate2900(.a(gate12inter0), .b(s_336), .O(gate12inter1));
  and2  gate2901(.a(G8), .b(G7), .O(gate12inter2));
  inv1  gate2902(.a(s_336), .O(gate12inter3));
  inv1  gate2903(.a(s_337), .O(gate12inter4));
  nand2 gate2904(.a(gate12inter4), .b(gate12inter3), .O(gate12inter5));
  nor2  gate2905(.a(gate12inter5), .b(gate12inter2), .O(gate12inter6));
  inv1  gate2906(.a(G7), .O(gate12inter7));
  inv1  gate2907(.a(G8), .O(gate12inter8));
  nand2 gate2908(.a(gate12inter8), .b(gate12inter7), .O(gate12inter9));
  nand2 gate2909(.a(s_337), .b(gate12inter3), .O(gate12inter10));
  nor2  gate2910(.a(gate12inter10), .b(gate12inter9), .O(gate12inter11));
  nor2  gate2911(.a(gate12inter11), .b(gate12inter6), .O(gate12inter12));
  nand2 gate2912(.a(gate12inter12), .b(gate12inter1), .O(G275));

  xor2  gate701(.a(G10), .b(G9), .O(gate13inter0));
  nand2 gate702(.a(gate13inter0), .b(s_22), .O(gate13inter1));
  and2  gate703(.a(G10), .b(G9), .O(gate13inter2));
  inv1  gate704(.a(s_22), .O(gate13inter3));
  inv1  gate705(.a(s_23), .O(gate13inter4));
  nand2 gate706(.a(gate13inter4), .b(gate13inter3), .O(gate13inter5));
  nor2  gate707(.a(gate13inter5), .b(gate13inter2), .O(gate13inter6));
  inv1  gate708(.a(G9), .O(gate13inter7));
  inv1  gate709(.a(G10), .O(gate13inter8));
  nand2 gate710(.a(gate13inter8), .b(gate13inter7), .O(gate13inter9));
  nand2 gate711(.a(s_23), .b(gate13inter3), .O(gate13inter10));
  nor2  gate712(.a(gate13inter10), .b(gate13inter9), .O(gate13inter11));
  nor2  gate713(.a(gate13inter11), .b(gate13inter6), .O(gate13inter12));
  nand2 gate714(.a(gate13inter12), .b(gate13inter1), .O(G278));

  xor2  gate2297(.a(G12), .b(G11), .O(gate14inter0));
  nand2 gate2298(.a(gate14inter0), .b(s_250), .O(gate14inter1));
  and2  gate2299(.a(G12), .b(G11), .O(gate14inter2));
  inv1  gate2300(.a(s_250), .O(gate14inter3));
  inv1  gate2301(.a(s_251), .O(gate14inter4));
  nand2 gate2302(.a(gate14inter4), .b(gate14inter3), .O(gate14inter5));
  nor2  gate2303(.a(gate14inter5), .b(gate14inter2), .O(gate14inter6));
  inv1  gate2304(.a(G11), .O(gate14inter7));
  inv1  gate2305(.a(G12), .O(gate14inter8));
  nand2 gate2306(.a(gate14inter8), .b(gate14inter7), .O(gate14inter9));
  nand2 gate2307(.a(s_251), .b(gate14inter3), .O(gate14inter10));
  nor2  gate2308(.a(gate14inter10), .b(gate14inter9), .O(gate14inter11));
  nor2  gate2309(.a(gate14inter11), .b(gate14inter6), .O(gate14inter12));
  nand2 gate2310(.a(gate14inter12), .b(gate14inter1), .O(G281));
nand2 gate15( .a(G13), .b(G14), .O(G284) );
nand2 gate16( .a(G15), .b(G16), .O(G287) );

  xor2  gate2367(.a(G18), .b(G17), .O(gate17inter0));
  nand2 gate2368(.a(gate17inter0), .b(s_260), .O(gate17inter1));
  and2  gate2369(.a(G18), .b(G17), .O(gate17inter2));
  inv1  gate2370(.a(s_260), .O(gate17inter3));
  inv1  gate2371(.a(s_261), .O(gate17inter4));
  nand2 gate2372(.a(gate17inter4), .b(gate17inter3), .O(gate17inter5));
  nor2  gate2373(.a(gate17inter5), .b(gate17inter2), .O(gate17inter6));
  inv1  gate2374(.a(G17), .O(gate17inter7));
  inv1  gate2375(.a(G18), .O(gate17inter8));
  nand2 gate2376(.a(gate17inter8), .b(gate17inter7), .O(gate17inter9));
  nand2 gate2377(.a(s_261), .b(gate17inter3), .O(gate17inter10));
  nor2  gate2378(.a(gate17inter10), .b(gate17inter9), .O(gate17inter11));
  nor2  gate2379(.a(gate17inter11), .b(gate17inter6), .O(gate17inter12));
  nand2 gate2380(.a(gate17inter12), .b(gate17inter1), .O(G290));

  xor2  gate2647(.a(G20), .b(G19), .O(gate18inter0));
  nand2 gate2648(.a(gate18inter0), .b(s_300), .O(gate18inter1));
  and2  gate2649(.a(G20), .b(G19), .O(gate18inter2));
  inv1  gate2650(.a(s_300), .O(gate18inter3));
  inv1  gate2651(.a(s_301), .O(gate18inter4));
  nand2 gate2652(.a(gate18inter4), .b(gate18inter3), .O(gate18inter5));
  nor2  gate2653(.a(gate18inter5), .b(gate18inter2), .O(gate18inter6));
  inv1  gate2654(.a(G19), .O(gate18inter7));
  inv1  gate2655(.a(G20), .O(gate18inter8));
  nand2 gate2656(.a(gate18inter8), .b(gate18inter7), .O(gate18inter9));
  nand2 gate2657(.a(s_301), .b(gate18inter3), .O(gate18inter10));
  nor2  gate2658(.a(gate18inter10), .b(gate18inter9), .O(gate18inter11));
  nor2  gate2659(.a(gate18inter11), .b(gate18inter6), .O(gate18inter12));
  nand2 gate2660(.a(gate18inter12), .b(gate18inter1), .O(G293));
nand2 gate19( .a(G21), .b(G22), .O(G296) );

  xor2  gate2073(.a(G24), .b(G23), .O(gate20inter0));
  nand2 gate2074(.a(gate20inter0), .b(s_218), .O(gate20inter1));
  and2  gate2075(.a(G24), .b(G23), .O(gate20inter2));
  inv1  gate2076(.a(s_218), .O(gate20inter3));
  inv1  gate2077(.a(s_219), .O(gate20inter4));
  nand2 gate2078(.a(gate20inter4), .b(gate20inter3), .O(gate20inter5));
  nor2  gate2079(.a(gate20inter5), .b(gate20inter2), .O(gate20inter6));
  inv1  gate2080(.a(G23), .O(gate20inter7));
  inv1  gate2081(.a(G24), .O(gate20inter8));
  nand2 gate2082(.a(gate20inter8), .b(gate20inter7), .O(gate20inter9));
  nand2 gate2083(.a(s_219), .b(gate20inter3), .O(gate20inter10));
  nor2  gate2084(.a(gate20inter10), .b(gate20inter9), .O(gate20inter11));
  nor2  gate2085(.a(gate20inter11), .b(gate20inter6), .O(gate20inter12));
  nand2 gate2086(.a(gate20inter12), .b(gate20inter1), .O(G299));

  xor2  gate939(.a(G26), .b(G25), .O(gate21inter0));
  nand2 gate940(.a(gate21inter0), .b(s_56), .O(gate21inter1));
  and2  gate941(.a(G26), .b(G25), .O(gate21inter2));
  inv1  gate942(.a(s_56), .O(gate21inter3));
  inv1  gate943(.a(s_57), .O(gate21inter4));
  nand2 gate944(.a(gate21inter4), .b(gate21inter3), .O(gate21inter5));
  nor2  gate945(.a(gate21inter5), .b(gate21inter2), .O(gate21inter6));
  inv1  gate946(.a(G25), .O(gate21inter7));
  inv1  gate947(.a(G26), .O(gate21inter8));
  nand2 gate948(.a(gate21inter8), .b(gate21inter7), .O(gate21inter9));
  nand2 gate949(.a(s_57), .b(gate21inter3), .O(gate21inter10));
  nor2  gate950(.a(gate21inter10), .b(gate21inter9), .O(gate21inter11));
  nor2  gate951(.a(gate21inter11), .b(gate21inter6), .O(gate21inter12));
  nand2 gate952(.a(gate21inter12), .b(gate21inter1), .O(G302));

  xor2  gate617(.a(G28), .b(G27), .O(gate22inter0));
  nand2 gate618(.a(gate22inter0), .b(s_10), .O(gate22inter1));
  and2  gate619(.a(G28), .b(G27), .O(gate22inter2));
  inv1  gate620(.a(s_10), .O(gate22inter3));
  inv1  gate621(.a(s_11), .O(gate22inter4));
  nand2 gate622(.a(gate22inter4), .b(gate22inter3), .O(gate22inter5));
  nor2  gate623(.a(gate22inter5), .b(gate22inter2), .O(gate22inter6));
  inv1  gate624(.a(G27), .O(gate22inter7));
  inv1  gate625(.a(G28), .O(gate22inter8));
  nand2 gate626(.a(gate22inter8), .b(gate22inter7), .O(gate22inter9));
  nand2 gate627(.a(s_11), .b(gate22inter3), .O(gate22inter10));
  nor2  gate628(.a(gate22inter10), .b(gate22inter9), .O(gate22inter11));
  nor2  gate629(.a(gate22inter11), .b(gate22inter6), .O(gate22inter12));
  nand2 gate630(.a(gate22inter12), .b(gate22inter1), .O(G305));

  xor2  gate1975(.a(G30), .b(G29), .O(gate23inter0));
  nand2 gate1976(.a(gate23inter0), .b(s_204), .O(gate23inter1));
  and2  gate1977(.a(G30), .b(G29), .O(gate23inter2));
  inv1  gate1978(.a(s_204), .O(gate23inter3));
  inv1  gate1979(.a(s_205), .O(gate23inter4));
  nand2 gate1980(.a(gate23inter4), .b(gate23inter3), .O(gate23inter5));
  nor2  gate1981(.a(gate23inter5), .b(gate23inter2), .O(gate23inter6));
  inv1  gate1982(.a(G29), .O(gate23inter7));
  inv1  gate1983(.a(G30), .O(gate23inter8));
  nand2 gate1984(.a(gate23inter8), .b(gate23inter7), .O(gate23inter9));
  nand2 gate1985(.a(s_205), .b(gate23inter3), .O(gate23inter10));
  nor2  gate1986(.a(gate23inter10), .b(gate23inter9), .O(gate23inter11));
  nor2  gate1987(.a(gate23inter11), .b(gate23inter6), .O(gate23inter12));
  nand2 gate1988(.a(gate23inter12), .b(gate23inter1), .O(G308));
nand2 gate24( .a(G31), .b(G32), .O(G311) );
nand2 gate25( .a(G1), .b(G5), .O(G314) );
nand2 gate26( .a(G9), .b(G13), .O(G317) );

  xor2  gate2241(.a(G6), .b(G2), .O(gate27inter0));
  nand2 gate2242(.a(gate27inter0), .b(s_242), .O(gate27inter1));
  and2  gate2243(.a(G6), .b(G2), .O(gate27inter2));
  inv1  gate2244(.a(s_242), .O(gate27inter3));
  inv1  gate2245(.a(s_243), .O(gate27inter4));
  nand2 gate2246(.a(gate27inter4), .b(gate27inter3), .O(gate27inter5));
  nor2  gate2247(.a(gate27inter5), .b(gate27inter2), .O(gate27inter6));
  inv1  gate2248(.a(G2), .O(gate27inter7));
  inv1  gate2249(.a(G6), .O(gate27inter8));
  nand2 gate2250(.a(gate27inter8), .b(gate27inter7), .O(gate27inter9));
  nand2 gate2251(.a(s_243), .b(gate27inter3), .O(gate27inter10));
  nor2  gate2252(.a(gate27inter10), .b(gate27inter9), .O(gate27inter11));
  nor2  gate2253(.a(gate27inter11), .b(gate27inter6), .O(gate27inter12));
  nand2 gate2254(.a(gate27inter12), .b(gate27inter1), .O(G320));
nand2 gate28( .a(G10), .b(G14), .O(G323) );
nand2 gate29( .a(G3), .b(G7), .O(G326) );
nand2 gate30( .a(G11), .b(G15), .O(G329) );

  xor2  gate1513(.a(G8), .b(G4), .O(gate31inter0));
  nand2 gate1514(.a(gate31inter0), .b(s_138), .O(gate31inter1));
  and2  gate1515(.a(G8), .b(G4), .O(gate31inter2));
  inv1  gate1516(.a(s_138), .O(gate31inter3));
  inv1  gate1517(.a(s_139), .O(gate31inter4));
  nand2 gate1518(.a(gate31inter4), .b(gate31inter3), .O(gate31inter5));
  nor2  gate1519(.a(gate31inter5), .b(gate31inter2), .O(gate31inter6));
  inv1  gate1520(.a(G4), .O(gate31inter7));
  inv1  gate1521(.a(G8), .O(gate31inter8));
  nand2 gate1522(.a(gate31inter8), .b(gate31inter7), .O(gate31inter9));
  nand2 gate1523(.a(s_139), .b(gate31inter3), .O(gate31inter10));
  nor2  gate1524(.a(gate31inter10), .b(gate31inter9), .O(gate31inter11));
  nor2  gate1525(.a(gate31inter11), .b(gate31inter6), .O(gate31inter12));
  nand2 gate1526(.a(gate31inter12), .b(gate31inter1), .O(G332));

  xor2  gate2787(.a(G16), .b(G12), .O(gate32inter0));
  nand2 gate2788(.a(gate32inter0), .b(s_320), .O(gate32inter1));
  and2  gate2789(.a(G16), .b(G12), .O(gate32inter2));
  inv1  gate2790(.a(s_320), .O(gate32inter3));
  inv1  gate2791(.a(s_321), .O(gate32inter4));
  nand2 gate2792(.a(gate32inter4), .b(gate32inter3), .O(gate32inter5));
  nor2  gate2793(.a(gate32inter5), .b(gate32inter2), .O(gate32inter6));
  inv1  gate2794(.a(G12), .O(gate32inter7));
  inv1  gate2795(.a(G16), .O(gate32inter8));
  nand2 gate2796(.a(gate32inter8), .b(gate32inter7), .O(gate32inter9));
  nand2 gate2797(.a(s_321), .b(gate32inter3), .O(gate32inter10));
  nor2  gate2798(.a(gate32inter10), .b(gate32inter9), .O(gate32inter11));
  nor2  gate2799(.a(gate32inter11), .b(gate32inter6), .O(gate32inter12));
  nand2 gate2800(.a(gate32inter12), .b(gate32inter1), .O(G335));

  xor2  gate729(.a(G21), .b(G17), .O(gate33inter0));
  nand2 gate730(.a(gate33inter0), .b(s_26), .O(gate33inter1));
  and2  gate731(.a(G21), .b(G17), .O(gate33inter2));
  inv1  gate732(.a(s_26), .O(gate33inter3));
  inv1  gate733(.a(s_27), .O(gate33inter4));
  nand2 gate734(.a(gate33inter4), .b(gate33inter3), .O(gate33inter5));
  nor2  gate735(.a(gate33inter5), .b(gate33inter2), .O(gate33inter6));
  inv1  gate736(.a(G17), .O(gate33inter7));
  inv1  gate737(.a(G21), .O(gate33inter8));
  nand2 gate738(.a(gate33inter8), .b(gate33inter7), .O(gate33inter9));
  nand2 gate739(.a(s_27), .b(gate33inter3), .O(gate33inter10));
  nor2  gate740(.a(gate33inter10), .b(gate33inter9), .O(gate33inter11));
  nor2  gate741(.a(gate33inter11), .b(gate33inter6), .O(gate33inter12));
  nand2 gate742(.a(gate33inter12), .b(gate33inter1), .O(G338));
nand2 gate34( .a(G25), .b(G29), .O(G341) );

  xor2  gate1023(.a(G22), .b(G18), .O(gate35inter0));
  nand2 gate1024(.a(gate35inter0), .b(s_68), .O(gate35inter1));
  and2  gate1025(.a(G22), .b(G18), .O(gate35inter2));
  inv1  gate1026(.a(s_68), .O(gate35inter3));
  inv1  gate1027(.a(s_69), .O(gate35inter4));
  nand2 gate1028(.a(gate35inter4), .b(gate35inter3), .O(gate35inter5));
  nor2  gate1029(.a(gate35inter5), .b(gate35inter2), .O(gate35inter6));
  inv1  gate1030(.a(G18), .O(gate35inter7));
  inv1  gate1031(.a(G22), .O(gate35inter8));
  nand2 gate1032(.a(gate35inter8), .b(gate35inter7), .O(gate35inter9));
  nand2 gate1033(.a(s_69), .b(gate35inter3), .O(gate35inter10));
  nor2  gate1034(.a(gate35inter10), .b(gate35inter9), .O(gate35inter11));
  nor2  gate1035(.a(gate35inter11), .b(gate35inter6), .O(gate35inter12));
  nand2 gate1036(.a(gate35inter12), .b(gate35inter1), .O(G344));

  xor2  gate2255(.a(G30), .b(G26), .O(gate36inter0));
  nand2 gate2256(.a(gate36inter0), .b(s_244), .O(gate36inter1));
  and2  gate2257(.a(G30), .b(G26), .O(gate36inter2));
  inv1  gate2258(.a(s_244), .O(gate36inter3));
  inv1  gate2259(.a(s_245), .O(gate36inter4));
  nand2 gate2260(.a(gate36inter4), .b(gate36inter3), .O(gate36inter5));
  nor2  gate2261(.a(gate36inter5), .b(gate36inter2), .O(gate36inter6));
  inv1  gate2262(.a(G26), .O(gate36inter7));
  inv1  gate2263(.a(G30), .O(gate36inter8));
  nand2 gate2264(.a(gate36inter8), .b(gate36inter7), .O(gate36inter9));
  nand2 gate2265(.a(s_245), .b(gate36inter3), .O(gate36inter10));
  nor2  gate2266(.a(gate36inter10), .b(gate36inter9), .O(gate36inter11));
  nor2  gate2267(.a(gate36inter11), .b(gate36inter6), .O(gate36inter12));
  nand2 gate2268(.a(gate36inter12), .b(gate36inter1), .O(G347));
nand2 gate37( .a(G19), .b(G23), .O(G350) );
nand2 gate38( .a(G27), .b(G31), .O(G353) );
nand2 gate39( .a(G20), .b(G24), .O(G356) );
nand2 gate40( .a(G28), .b(G32), .O(G359) );

  xor2  gate2535(.a(G266), .b(G1), .O(gate41inter0));
  nand2 gate2536(.a(gate41inter0), .b(s_284), .O(gate41inter1));
  and2  gate2537(.a(G266), .b(G1), .O(gate41inter2));
  inv1  gate2538(.a(s_284), .O(gate41inter3));
  inv1  gate2539(.a(s_285), .O(gate41inter4));
  nand2 gate2540(.a(gate41inter4), .b(gate41inter3), .O(gate41inter5));
  nor2  gate2541(.a(gate41inter5), .b(gate41inter2), .O(gate41inter6));
  inv1  gate2542(.a(G1), .O(gate41inter7));
  inv1  gate2543(.a(G266), .O(gate41inter8));
  nand2 gate2544(.a(gate41inter8), .b(gate41inter7), .O(gate41inter9));
  nand2 gate2545(.a(s_285), .b(gate41inter3), .O(gate41inter10));
  nor2  gate2546(.a(gate41inter10), .b(gate41inter9), .O(gate41inter11));
  nor2  gate2547(.a(gate41inter11), .b(gate41inter6), .O(gate41inter12));
  nand2 gate2548(.a(gate41inter12), .b(gate41inter1), .O(G362));

  xor2  gate1961(.a(G266), .b(G2), .O(gate42inter0));
  nand2 gate1962(.a(gate42inter0), .b(s_202), .O(gate42inter1));
  and2  gate1963(.a(G266), .b(G2), .O(gate42inter2));
  inv1  gate1964(.a(s_202), .O(gate42inter3));
  inv1  gate1965(.a(s_203), .O(gate42inter4));
  nand2 gate1966(.a(gate42inter4), .b(gate42inter3), .O(gate42inter5));
  nor2  gate1967(.a(gate42inter5), .b(gate42inter2), .O(gate42inter6));
  inv1  gate1968(.a(G2), .O(gate42inter7));
  inv1  gate1969(.a(G266), .O(gate42inter8));
  nand2 gate1970(.a(gate42inter8), .b(gate42inter7), .O(gate42inter9));
  nand2 gate1971(.a(s_203), .b(gate42inter3), .O(gate42inter10));
  nor2  gate1972(.a(gate42inter10), .b(gate42inter9), .O(gate42inter11));
  nor2  gate1973(.a(gate42inter11), .b(gate42inter6), .O(gate42inter12));
  nand2 gate1974(.a(gate42inter12), .b(gate42inter1), .O(G363));
nand2 gate43( .a(G3), .b(G269), .O(G364) );

  xor2  gate2325(.a(G269), .b(G4), .O(gate44inter0));
  nand2 gate2326(.a(gate44inter0), .b(s_254), .O(gate44inter1));
  and2  gate2327(.a(G269), .b(G4), .O(gate44inter2));
  inv1  gate2328(.a(s_254), .O(gate44inter3));
  inv1  gate2329(.a(s_255), .O(gate44inter4));
  nand2 gate2330(.a(gate44inter4), .b(gate44inter3), .O(gate44inter5));
  nor2  gate2331(.a(gate44inter5), .b(gate44inter2), .O(gate44inter6));
  inv1  gate2332(.a(G4), .O(gate44inter7));
  inv1  gate2333(.a(G269), .O(gate44inter8));
  nand2 gate2334(.a(gate44inter8), .b(gate44inter7), .O(gate44inter9));
  nand2 gate2335(.a(s_255), .b(gate44inter3), .O(gate44inter10));
  nor2  gate2336(.a(gate44inter10), .b(gate44inter9), .O(gate44inter11));
  nor2  gate2337(.a(gate44inter11), .b(gate44inter6), .O(gate44inter12));
  nand2 gate2338(.a(gate44inter12), .b(gate44inter1), .O(G365));

  xor2  gate2059(.a(G272), .b(G5), .O(gate45inter0));
  nand2 gate2060(.a(gate45inter0), .b(s_216), .O(gate45inter1));
  and2  gate2061(.a(G272), .b(G5), .O(gate45inter2));
  inv1  gate2062(.a(s_216), .O(gate45inter3));
  inv1  gate2063(.a(s_217), .O(gate45inter4));
  nand2 gate2064(.a(gate45inter4), .b(gate45inter3), .O(gate45inter5));
  nor2  gate2065(.a(gate45inter5), .b(gate45inter2), .O(gate45inter6));
  inv1  gate2066(.a(G5), .O(gate45inter7));
  inv1  gate2067(.a(G272), .O(gate45inter8));
  nand2 gate2068(.a(gate45inter8), .b(gate45inter7), .O(gate45inter9));
  nand2 gate2069(.a(s_217), .b(gate45inter3), .O(gate45inter10));
  nor2  gate2070(.a(gate45inter10), .b(gate45inter9), .O(gate45inter11));
  nor2  gate2071(.a(gate45inter11), .b(gate45inter6), .O(gate45inter12));
  nand2 gate2072(.a(gate45inter12), .b(gate45inter1), .O(G366));
nand2 gate46( .a(G6), .b(G272), .O(G367) );

  xor2  gate1051(.a(G275), .b(G7), .O(gate47inter0));
  nand2 gate1052(.a(gate47inter0), .b(s_72), .O(gate47inter1));
  and2  gate1053(.a(G275), .b(G7), .O(gate47inter2));
  inv1  gate1054(.a(s_72), .O(gate47inter3));
  inv1  gate1055(.a(s_73), .O(gate47inter4));
  nand2 gate1056(.a(gate47inter4), .b(gate47inter3), .O(gate47inter5));
  nor2  gate1057(.a(gate47inter5), .b(gate47inter2), .O(gate47inter6));
  inv1  gate1058(.a(G7), .O(gate47inter7));
  inv1  gate1059(.a(G275), .O(gate47inter8));
  nand2 gate1060(.a(gate47inter8), .b(gate47inter7), .O(gate47inter9));
  nand2 gate1061(.a(s_73), .b(gate47inter3), .O(gate47inter10));
  nor2  gate1062(.a(gate47inter10), .b(gate47inter9), .O(gate47inter11));
  nor2  gate1063(.a(gate47inter11), .b(gate47inter6), .O(gate47inter12));
  nand2 gate1064(.a(gate47inter12), .b(gate47inter1), .O(G368));

  xor2  gate1597(.a(G275), .b(G8), .O(gate48inter0));
  nand2 gate1598(.a(gate48inter0), .b(s_150), .O(gate48inter1));
  and2  gate1599(.a(G275), .b(G8), .O(gate48inter2));
  inv1  gate1600(.a(s_150), .O(gate48inter3));
  inv1  gate1601(.a(s_151), .O(gate48inter4));
  nand2 gate1602(.a(gate48inter4), .b(gate48inter3), .O(gate48inter5));
  nor2  gate1603(.a(gate48inter5), .b(gate48inter2), .O(gate48inter6));
  inv1  gate1604(.a(G8), .O(gate48inter7));
  inv1  gate1605(.a(G275), .O(gate48inter8));
  nand2 gate1606(.a(gate48inter8), .b(gate48inter7), .O(gate48inter9));
  nand2 gate1607(.a(s_151), .b(gate48inter3), .O(gate48inter10));
  nor2  gate1608(.a(gate48inter10), .b(gate48inter9), .O(gate48inter11));
  nor2  gate1609(.a(gate48inter11), .b(gate48inter6), .O(gate48inter12));
  nand2 gate1610(.a(gate48inter12), .b(gate48inter1), .O(G369));
nand2 gate49( .a(G9), .b(G278), .O(G370) );

  xor2  gate645(.a(G278), .b(G10), .O(gate50inter0));
  nand2 gate646(.a(gate50inter0), .b(s_14), .O(gate50inter1));
  and2  gate647(.a(G278), .b(G10), .O(gate50inter2));
  inv1  gate648(.a(s_14), .O(gate50inter3));
  inv1  gate649(.a(s_15), .O(gate50inter4));
  nand2 gate650(.a(gate50inter4), .b(gate50inter3), .O(gate50inter5));
  nor2  gate651(.a(gate50inter5), .b(gate50inter2), .O(gate50inter6));
  inv1  gate652(.a(G10), .O(gate50inter7));
  inv1  gate653(.a(G278), .O(gate50inter8));
  nand2 gate654(.a(gate50inter8), .b(gate50inter7), .O(gate50inter9));
  nand2 gate655(.a(s_15), .b(gate50inter3), .O(gate50inter10));
  nor2  gate656(.a(gate50inter10), .b(gate50inter9), .O(gate50inter11));
  nor2  gate657(.a(gate50inter11), .b(gate50inter6), .O(gate50inter12));
  nand2 gate658(.a(gate50inter12), .b(gate50inter1), .O(G371));

  xor2  gate841(.a(G281), .b(G11), .O(gate51inter0));
  nand2 gate842(.a(gate51inter0), .b(s_42), .O(gate51inter1));
  and2  gate843(.a(G281), .b(G11), .O(gate51inter2));
  inv1  gate844(.a(s_42), .O(gate51inter3));
  inv1  gate845(.a(s_43), .O(gate51inter4));
  nand2 gate846(.a(gate51inter4), .b(gate51inter3), .O(gate51inter5));
  nor2  gate847(.a(gate51inter5), .b(gate51inter2), .O(gate51inter6));
  inv1  gate848(.a(G11), .O(gate51inter7));
  inv1  gate849(.a(G281), .O(gate51inter8));
  nand2 gate850(.a(gate51inter8), .b(gate51inter7), .O(gate51inter9));
  nand2 gate851(.a(s_43), .b(gate51inter3), .O(gate51inter10));
  nor2  gate852(.a(gate51inter10), .b(gate51inter9), .O(gate51inter11));
  nor2  gate853(.a(gate51inter11), .b(gate51inter6), .O(gate51inter12));
  nand2 gate854(.a(gate51inter12), .b(gate51inter1), .O(G372));
nand2 gate52( .a(G12), .b(G281), .O(G373) );
nand2 gate53( .a(G13), .b(G284), .O(G374) );
nand2 gate54( .a(G14), .b(G284), .O(G375) );
nand2 gate55( .a(G15), .b(G287), .O(G376) );
nand2 gate56( .a(G16), .b(G287), .O(G377) );
nand2 gate57( .a(G17), .b(G290), .O(G378) );

  xor2  gate1457(.a(G290), .b(G18), .O(gate58inter0));
  nand2 gate1458(.a(gate58inter0), .b(s_130), .O(gate58inter1));
  and2  gate1459(.a(G290), .b(G18), .O(gate58inter2));
  inv1  gate1460(.a(s_130), .O(gate58inter3));
  inv1  gate1461(.a(s_131), .O(gate58inter4));
  nand2 gate1462(.a(gate58inter4), .b(gate58inter3), .O(gate58inter5));
  nor2  gate1463(.a(gate58inter5), .b(gate58inter2), .O(gate58inter6));
  inv1  gate1464(.a(G18), .O(gate58inter7));
  inv1  gate1465(.a(G290), .O(gate58inter8));
  nand2 gate1466(.a(gate58inter8), .b(gate58inter7), .O(gate58inter9));
  nand2 gate1467(.a(s_131), .b(gate58inter3), .O(gate58inter10));
  nor2  gate1468(.a(gate58inter10), .b(gate58inter9), .O(gate58inter11));
  nor2  gate1469(.a(gate58inter11), .b(gate58inter6), .O(gate58inter12));
  nand2 gate1470(.a(gate58inter12), .b(gate58inter1), .O(G379));
nand2 gate59( .a(G19), .b(G293), .O(G380) );

  xor2  gate981(.a(G293), .b(G20), .O(gate60inter0));
  nand2 gate982(.a(gate60inter0), .b(s_62), .O(gate60inter1));
  and2  gate983(.a(G293), .b(G20), .O(gate60inter2));
  inv1  gate984(.a(s_62), .O(gate60inter3));
  inv1  gate985(.a(s_63), .O(gate60inter4));
  nand2 gate986(.a(gate60inter4), .b(gate60inter3), .O(gate60inter5));
  nor2  gate987(.a(gate60inter5), .b(gate60inter2), .O(gate60inter6));
  inv1  gate988(.a(G20), .O(gate60inter7));
  inv1  gate989(.a(G293), .O(gate60inter8));
  nand2 gate990(.a(gate60inter8), .b(gate60inter7), .O(gate60inter9));
  nand2 gate991(.a(s_63), .b(gate60inter3), .O(gate60inter10));
  nor2  gate992(.a(gate60inter10), .b(gate60inter9), .O(gate60inter11));
  nor2  gate993(.a(gate60inter11), .b(gate60inter6), .O(gate60inter12));
  nand2 gate994(.a(gate60inter12), .b(gate60inter1), .O(G381));
nand2 gate61( .a(G21), .b(G296), .O(G382) );
nand2 gate62( .a(G22), .b(G296), .O(G383) );
nand2 gate63( .a(G23), .b(G299), .O(G384) );
nand2 gate64( .a(G24), .b(G299), .O(G385) );

  xor2  gate1933(.a(G302), .b(G25), .O(gate65inter0));
  nand2 gate1934(.a(gate65inter0), .b(s_198), .O(gate65inter1));
  and2  gate1935(.a(G302), .b(G25), .O(gate65inter2));
  inv1  gate1936(.a(s_198), .O(gate65inter3));
  inv1  gate1937(.a(s_199), .O(gate65inter4));
  nand2 gate1938(.a(gate65inter4), .b(gate65inter3), .O(gate65inter5));
  nor2  gate1939(.a(gate65inter5), .b(gate65inter2), .O(gate65inter6));
  inv1  gate1940(.a(G25), .O(gate65inter7));
  inv1  gate1941(.a(G302), .O(gate65inter8));
  nand2 gate1942(.a(gate65inter8), .b(gate65inter7), .O(gate65inter9));
  nand2 gate1943(.a(s_199), .b(gate65inter3), .O(gate65inter10));
  nor2  gate1944(.a(gate65inter10), .b(gate65inter9), .O(gate65inter11));
  nor2  gate1945(.a(gate65inter11), .b(gate65inter6), .O(gate65inter12));
  nand2 gate1946(.a(gate65inter12), .b(gate65inter1), .O(G386));
nand2 gate66( .a(G26), .b(G302), .O(G387) );
nand2 gate67( .a(G27), .b(G305), .O(G388) );
nand2 gate68( .a(G28), .b(G305), .O(G389) );
nand2 gate69( .a(G29), .b(G308), .O(G390) );
nand2 gate70( .a(G30), .b(G308), .O(G391) );
nand2 gate71( .a(G31), .b(G311), .O(G392) );
nand2 gate72( .a(G32), .b(G311), .O(G393) );
nand2 gate73( .a(G1), .b(G314), .O(G394) );
nand2 gate74( .a(G5), .b(G314), .O(G395) );
nand2 gate75( .a(G9), .b(G317), .O(G396) );
nand2 gate76( .a(G13), .b(G317), .O(G397) );

  xor2  gate1947(.a(G320), .b(G2), .O(gate77inter0));
  nand2 gate1948(.a(gate77inter0), .b(s_200), .O(gate77inter1));
  and2  gate1949(.a(G320), .b(G2), .O(gate77inter2));
  inv1  gate1950(.a(s_200), .O(gate77inter3));
  inv1  gate1951(.a(s_201), .O(gate77inter4));
  nand2 gate1952(.a(gate77inter4), .b(gate77inter3), .O(gate77inter5));
  nor2  gate1953(.a(gate77inter5), .b(gate77inter2), .O(gate77inter6));
  inv1  gate1954(.a(G2), .O(gate77inter7));
  inv1  gate1955(.a(G320), .O(gate77inter8));
  nand2 gate1956(.a(gate77inter8), .b(gate77inter7), .O(gate77inter9));
  nand2 gate1957(.a(s_201), .b(gate77inter3), .O(gate77inter10));
  nor2  gate1958(.a(gate77inter10), .b(gate77inter9), .O(gate77inter11));
  nor2  gate1959(.a(gate77inter11), .b(gate77inter6), .O(gate77inter12));
  nand2 gate1960(.a(gate77inter12), .b(gate77inter1), .O(G398));
nand2 gate78( .a(G6), .b(G320), .O(G399) );
nand2 gate79( .a(G10), .b(G323), .O(G400) );
nand2 gate80( .a(G14), .b(G323), .O(G401) );
nand2 gate81( .a(G3), .b(G326), .O(G402) );
nand2 gate82( .a(G7), .b(G326), .O(G403) );
nand2 gate83( .a(G11), .b(G329), .O(G404) );
nand2 gate84( .a(G15), .b(G329), .O(G405) );

  xor2  gate2731(.a(G332), .b(G4), .O(gate85inter0));
  nand2 gate2732(.a(gate85inter0), .b(s_312), .O(gate85inter1));
  and2  gate2733(.a(G332), .b(G4), .O(gate85inter2));
  inv1  gate2734(.a(s_312), .O(gate85inter3));
  inv1  gate2735(.a(s_313), .O(gate85inter4));
  nand2 gate2736(.a(gate85inter4), .b(gate85inter3), .O(gate85inter5));
  nor2  gate2737(.a(gate85inter5), .b(gate85inter2), .O(gate85inter6));
  inv1  gate2738(.a(G4), .O(gate85inter7));
  inv1  gate2739(.a(G332), .O(gate85inter8));
  nand2 gate2740(.a(gate85inter8), .b(gate85inter7), .O(gate85inter9));
  nand2 gate2741(.a(s_313), .b(gate85inter3), .O(gate85inter10));
  nor2  gate2742(.a(gate85inter10), .b(gate85inter9), .O(gate85inter11));
  nor2  gate2743(.a(gate85inter11), .b(gate85inter6), .O(gate85inter12));
  nand2 gate2744(.a(gate85inter12), .b(gate85inter1), .O(G406));

  xor2  gate2227(.a(G332), .b(G8), .O(gate86inter0));
  nand2 gate2228(.a(gate86inter0), .b(s_240), .O(gate86inter1));
  and2  gate2229(.a(G332), .b(G8), .O(gate86inter2));
  inv1  gate2230(.a(s_240), .O(gate86inter3));
  inv1  gate2231(.a(s_241), .O(gate86inter4));
  nand2 gate2232(.a(gate86inter4), .b(gate86inter3), .O(gate86inter5));
  nor2  gate2233(.a(gate86inter5), .b(gate86inter2), .O(gate86inter6));
  inv1  gate2234(.a(G8), .O(gate86inter7));
  inv1  gate2235(.a(G332), .O(gate86inter8));
  nand2 gate2236(.a(gate86inter8), .b(gate86inter7), .O(gate86inter9));
  nand2 gate2237(.a(s_241), .b(gate86inter3), .O(gate86inter10));
  nor2  gate2238(.a(gate86inter10), .b(gate86inter9), .O(gate86inter11));
  nor2  gate2239(.a(gate86inter11), .b(gate86inter6), .O(gate86inter12));
  nand2 gate2240(.a(gate86inter12), .b(gate86inter1), .O(G407));

  xor2  gate1065(.a(G335), .b(G12), .O(gate87inter0));
  nand2 gate1066(.a(gate87inter0), .b(s_74), .O(gate87inter1));
  and2  gate1067(.a(G335), .b(G12), .O(gate87inter2));
  inv1  gate1068(.a(s_74), .O(gate87inter3));
  inv1  gate1069(.a(s_75), .O(gate87inter4));
  nand2 gate1070(.a(gate87inter4), .b(gate87inter3), .O(gate87inter5));
  nor2  gate1071(.a(gate87inter5), .b(gate87inter2), .O(gate87inter6));
  inv1  gate1072(.a(G12), .O(gate87inter7));
  inv1  gate1073(.a(G335), .O(gate87inter8));
  nand2 gate1074(.a(gate87inter8), .b(gate87inter7), .O(gate87inter9));
  nand2 gate1075(.a(s_75), .b(gate87inter3), .O(gate87inter10));
  nor2  gate1076(.a(gate87inter10), .b(gate87inter9), .O(gate87inter11));
  nor2  gate1077(.a(gate87inter11), .b(gate87inter6), .O(gate87inter12));
  nand2 gate1078(.a(gate87inter12), .b(gate87inter1), .O(G408));
nand2 gate88( .a(G16), .b(G335), .O(G409) );
nand2 gate89( .a(G17), .b(G338), .O(G410) );
nand2 gate90( .a(G21), .b(G338), .O(G411) );
nand2 gate91( .a(G25), .b(G341), .O(G412) );
nand2 gate92( .a(G29), .b(G341), .O(G413) );
nand2 gate93( .a(G18), .b(G344), .O(G414) );
nand2 gate94( .a(G22), .b(G344), .O(G415) );
nand2 gate95( .a(G26), .b(G347), .O(G416) );
nand2 gate96( .a(G30), .b(G347), .O(G417) );
nand2 gate97( .a(G19), .b(G350), .O(G418) );
nand2 gate98( .a(G23), .b(G350), .O(G419) );

  xor2  gate1709(.a(G353), .b(G27), .O(gate99inter0));
  nand2 gate1710(.a(gate99inter0), .b(s_166), .O(gate99inter1));
  and2  gate1711(.a(G353), .b(G27), .O(gate99inter2));
  inv1  gate1712(.a(s_166), .O(gate99inter3));
  inv1  gate1713(.a(s_167), .O(gate99inter4));
  nand2 gate1714(.a(gate99inter4), .b(gate99inter3), .O(gate99inter5));
  nor2  gate1715(.a(gate99inter5), .b(gate99inter2), .O(gate99inter6));
  inv1  gate1716(.a(G27), .O(gate99inter7));
  inv1  gate1717(.a(G353), .O(gate99inter8));
  nand2 gate1718(.a(gate99inter8), .b(gate99inter7), .O(gate99inter9));
  nand2 gate1719(.a(s_167), .b(gate99inter3), .O(gate99inter10));
  nor2  gate1720(.a(gate99inter10), .b(gate99inter9), .O(gate99inter11));
  nor2  gate1721(.a(gate99inter11), .b(gate99inter6), .O(gate99inter12));
  nand2 gate1722(.a(gate99inter12), .b(gate99inter1), .O(G420));
nand2 gate100( .a(G31), .b(G353), .O(G421) );
nand2 gate101( .a(G20), .b(G356), .O(G422) );
nand2 gate102( .a(G24), .b(G356), .O(G423) );

  xor2  gate1135(.a(G359), .b(G28), .O(gate103inter0));
  nand2 gate1136(.a(gate103inter0), .b(s_84), .O(gate103inter1));
  and2  gate1137(.a(G359), .b(G28), .O(gate103inter2));
  inv1  gate1138(.a(s_84), .O(gate103inter3));
  inv1  gate1139(.a(s_85), .O(gate103inter4));
  nand2 gate1140(.a(gate103inter4), .b(gate103inter3), .O(gate103inter5));
  nor2  gate1141(.a(gate103inter5), .b(gate103inter2), .O(gate103inter6));
  inv1  gate1142(.a(G28), .O(gate103inter7));
  inv1  gate1143(.a(G359), .O(gate103inter8));
  nand2 gate1144(.a(gate103inter8), .b(gate103inter7), .O(gate103inter9));
  nand2 gate1145(.a(s_85), .b(gate103inter3), .O(gate103inter10));
  nor2  gate1146(.a(gate103inter10), .b(gate103inter9), .O(gate103inter11));
  nor2  gate1147(.a(gate103inter11), .b(gate103inter6), .O(gate103inter12));
  nand2 gate1148(.a(gate103inter12), .b(gate103inter1), .O(G424));

  xor2  gate2395(.a(G359), .b(G32), .O(gate104inter0));
  nand2 gate2396(.a(gate104inter0), .b(s_264), .O(gate104inter1));
  and2  gate2397(.a(G359), .b(G32), .O(gate104inter2));
  inv1  gate2398(.a(s_264), .O(gate104inter3));
  inv1  gate2399(.a(s_265), .O(gate104inter4));
  nand2 gate2400(.a(gate104inter4), .b(gate104inter3), .O(gate104inter5));
  nor2  gate2401(.a(gate104inter5), .b(gate104inter2), .O(gate104inter6));
  inv1  gate2402(.a(G32), .O(gate104inter7));
  inv1  gate2403(.a(G359), .O(gate104inter8));
  nand2 gate2404(.a(gate104inter8), .b(gate104inter7), .O(gate104inter9));
  nand2 gate2405(.a(s_265), .b(gate104inter3), .O(gate104inter10));
  nor2  gate2406(.a(gate104inter10), .b(gate104inter9), .O(gate104inter11));
  nor2  gate2407(.a(gate104inter11), .b(gate104inter6), .O(gate104inter12));
  nand2 gate2408(.a(gate104inter12), .b(gate104inter1), .O(G425));
nand2 gate105( .a(G362), .b(G363), .O(G426) );
nand2 gate106( .a(G364), .b(G365), .O(G429) );
nand2 gate107( .a(G366), .b(G367), .O(G432) );

  xor2  gate2479(.a(G369), .b(G368), .O(gate108inter0));
  nand2 gate2480(.a(gate108inter0), .b(s_276), .O(gate108inter1));
  and2  gate2481(.a(G369), .b(G368), .O(gate108inter2));
  inv1  gate2482(.a(s_276), .O(gate108inter3));
  inv1  gate2483(.a(s_277), .O(gate108inter4));
  nand2 gate2484(.a(gate108inter4), .b(gate108inter3), .O(gate108inter5));
  nor2  gate2485(.a(gate108inter5), .b(gate108inter2), .O(gate108inter6));
  inv1  gate2486(.a(G368), .O(gate108inter7));
  inv1  gate2487(.a(G369), .O(gate108inter8));
  nand2 gate2488(.a(gate108inter8), .b(gate108inter7), .O(gate108inter9));
  nand2 gate2489(.a(s_277), .b(gate108inter3), .O(gate108inter10));
  nor2  gate2490(.a(gate108inter10), .b(gate108inter9), .O(gate108inter11));
  nor2  gate2491(.a(gate108inter11), .b(gate108inter6), .O(gate108inter12));
  nand2 gate2492(.a(gate108inter12), .b(gate108inter1), .O(G435));
nand2 gate109( .a(G370), .b(G371), .O(G438) );
nand2 gate110( .a(G372), .b(G373), .O(G441) );
nand2 gate111( .a(G374), .b(G375), .O(G444) );

  xor2  gate2339(.a(G377), .b(G376), .O(gate112inter0));
  nand2 gate2340(.a(gate112inter0), .b(s_256), .O(gate112inter1));
  and2  gate2341(.a(G377), .b(G376), .O(gate112inter2));
  inv1  gate2342(.a(s_256), .O(gate112inter3));
  inv1  gate2343(.a(s_257), .O(gate112inter4));
  nand2 gate2344(.a(gate112inter4), .b(gate112inter3), .O(gate112inter5));
  nor2  gate2345(.a(gate112inter5), .b(gate112inter2), .O(gate112inter6));
  inv1  gate2346(.a(G376), .O(gate112inter7));
  inv1  gate2347(.a(G377), .O(gate112inter8));
  nand2 gate2348(.a(gate112inter8), .b(gate112inter7), .O(gate112inter9));
  nand2 gate2349(.a(s_257), .b(gate112inter3), .O(gate112inter10));
  nor2  gate2350(.a(gate112inter10), .b(gate112inter9), .O(gate112inter11));
  nor2  gate2351(.a(gate112inter11), .b(gate112inter6), .O(gate112inter12));
  nand2 gate2352(.a(gate112inter12), .b(gate112inter1), .O(G447));

  xor2  gate1737(.a(G379), .b(G378), .O(gate113inter0));
  nand2 gate1738(.a(gate113inter0), .b(s_170), .O(gate113inter1));
  and2  gate1739(.a(G379), .b(G378), .O(gate113inter2));
  inv1  gate1740(.a(s_170), .O(gate113inter3));
  inv1  gate1741(.a(s_171), .O(gate113inter4));
  nand2 gate1742(.a(gate113inter4), .b(gate113inter3), .O(gate113inter5));
  nor2  gate1743(.a(gate113inter5), .b(gate113inter2), .O(gate113inter6));
  inv1  gate1744(.a(G378), .O(gate113inter7));
  inv1  gate1745(.a(G379), .O(gate113inter8));
  nand2 gate1746(.a(gate113inter8), .b(gate113inter7), .O(gate113inter9));
  nand2 gate1747(.a(s_171), .b(gate113inter3), .O(gate113inter10));
  nor2  gate1748(.a(gate113inter10), .b(gate113inter9), .O(gate113inter11));
  nor2  gate1749(.a(gate113inter11), .b(gate113inter6), .O(gate113inter12));
  nand2 gate1750(.a(gate113inter12), .b(gate113inter1), .O(G450));
nand2 gate114( .a(G380), .b(G381), .O(G453) );
nand2 gate115( .a(G382), .b(G383), .O(G456) );
nand2 gate116( .a(G384), .b(G385), .O(G459) );

  xor2  gate1387(.a(G387), .b(G386), .O(gate117inter0));
  nand2 gate1388(.a(gate117inter0), .b(s_120), .O(gate117inter1));
  and2  gate1389(.a(G387), .b(G386), .O(gate117inter2));
  inv1  gate1390(.a(s_120), .O(gate117inter3));
  inv1  gate1391(.a(s_121), .O(gate117inter4));
  nand2 gate1392(.a(gate117inter4), .b(gate117inter3), .O(gate117inter5));
  nor2  gate1393(.a(gate117inter5), .b(gate117inter2), .O(gate117inter6));
  inv1  gate1394(.a(G386), .O(gate117inter7));
  inv1  gate1395(.a(G387), .O(gate117inter8));
  nand2 gate1396(.a(gate117inter8), .b(gate117inter7), .O(gate117inter9));
  nand2 gate1397(.a(s_121), .b(gate117inter3), .O(gate117inter10));
  nor2  gate1398(.a(gate117inter10), .b(gate117inter9), .O(gate117inter11));
  nor2  gate1399(.a(gate117inter11), .b(gate117inter6), .O(gate117inter12));
  nand2 gate1400(.a(gate117inter12), .b(gate117inter1), .O(G462));

  xor2  gate1569(.a(G389), .b(G388), .O(gate118inter0));
  nand2 gate1570(.a(gate118inter0), .b(s_146), .O(gate118inter1));
  and2  gate1571(.a(G389), .b(G388), .O(gate118inter2));
  inv1  gate1572(.a(s_146), .O(gate118inter3));
  inv1  gate1573(.a(s_147), .O(gate118inter4));
  nand2 gate1574(.a(gate118inter4), .b(gate118inter3), .O(gate118inter5));
  nor2  gate1575(.a(gate118inter5), .b(gate118inter2), .O(gate118inter6));
  inv1  gate1576(.a(G388), .O(gate118inter7));
  inv1  gate1577(.a(G389), .O(gate118inter8));
  nand2 gate1578(.a(gate118inter8), .b(gate118inter7), .O(gate118inter9));
  nand2 gate1579(.a(s_147), .b(gate118inter3), .O(gate118inter10));
  nor2  gate1580(.a(gate118inter10), .b(gate118inter9), .O(gate118inter11));
  nor2  gate1581(.a(gate118inter11), .b(gate118inter6), .O(gate118inter12));
  nand2 gate1582(.a(gate118inter12), .b(gate118inter1), .O(G465));
nand2 gate119( .a(G390), .b(G391), .O(G468) );

  xor2  gate2591(.a(G393), .b(G392), .O(gate120inter0));
  nand2 gate2592(.a(gate120inter0), .b(s_292), .O(gate120inter1));
  and2  gate2593(.a(G393), .b(G392), .O(gate120inter2));
  inv1  gate2594(.a(s_292), .O(gate120inter3));
  inv1  gate2595(.a(s_293), .O(gate120inter4));
  nand2 gate2596(.a(gate120inter4), .b(gate120inter3), .O(gate120inter5));
  nor2  gate2597(.a(gate120inter5), .b(gate120inter2), .O(gate120inter6));
  inv1  gate2598(.a(G392), .O(gate120inter7));
  inv1  gate2599(.a(G393), .O(gate120inter8));
  nand2 gate2600(.a(gate120inter8), .b(gate120inter7), .O(gate120inter9));
  nand2 gate2601(.a(s_293), .b(gate120inter3), .O(gate120inter10));
  nor2  gate2602(.a(gate120inter10), .b(gate120inter9), .O(gate120inter11));
  nor2  gate2603(.a(gate120inter11), .b(gate120inter6), .O(gate120inter12));
  nand2 gate2604(.a(gate120inter12), .b(gate120inter1), .O(G471));
nand2 gate121( .a(G394), .b(G395), .O(G474) );

  xor2  gate2619(.a(G397), .b(G396), .O(gate122inter0));
  nand2 gate2620(.a(gate122inter0), .b(s_296), .O(gate122inter1));
  and2  gate2621(.a(G397), .b(G396), .O(gate122inter2));
  inv1  gate2622(.a(s_296), .O(gate122inter3));
  inv1  gate2623(.a(s_297), .O(gate122inter4));
  nand2 gate2624(.a(gate122inter4), .b(gate122inter3), .O(gate122inter5));
  nor2  gate2625(.a(gate122inter5), .b(gate122inter2), .O(gate122inter6));
  inv1  gate2626(.a(G396), .O(gate122inter7));
  inv1  gate2627(.a(G397), .O(gate122inter8));
  nand2 gate2628(.a(gate122inter8), .b(gate122inter7), .O(gate122inter9));
  nand2 gate2629(.a(s_297), .b(gate122inter3), .O(gate122inter10));
  nor2  gate2630(.a(gate122inter10), .b(gate122inter9), .O(gate122inter11));
  nor2  gate2631(.a(gate122inter11), .b(gate122inter6), .O(gate122inter12));
  nand2 gate2632(.a(gate122inter12), .b(gate122inter1), .O(G477));

  xor2  gate1821(.a(G399), .b(G398), .O(gate123inter0));
  nand2 gate1822(.a(gate123inter0), .b(s_182), .O(gate123inter1));
  and2  gate1823(.a(G399), .b(G398), .O(gate123inter2));
  inv1  gate1824(.a(s_182), .O(gate123inter3));
  inv1  gate1825(.a(s_183), .O(gate123inter4));
  nand2 gate1826(.a(gate123inter4), .b(gate123inter3), .O(gate123inter5));
  nor2  gate1827(.a(gate123inter5), .b(gate123inter2), .O(gate123inter6));
  inv1  gate1828(.a(G398), .O(gate123inter7));
  inv1  gate1829(.a(G399), .O(gate123inter8));
  nand2 gate1830(.a(gate123inter8), .b(gate123inter7), .O(gate123inter9));
  nand2 gate1831(.a(s_183), .b(gate123inter3), .O(gate123inter10));
  nor2  gate1832(.a(gate123inter10), .b(gate123inter9), .O(gate123inter11));
  nor2  gate1833(.a(gate123inter11), .b(gate123inter6), .O(gate123inter12));
  nand2 gate1834(.a(gate123inter12), .b(gate123inter1), .O(G480));
nand2 gate124( .a(G400), .b(G401), .O(G483) );

  xor2  gate2703(.a(G403), .b(G402), .O(gate125inter0));
  nand2 gate2704(.a(gate125inter0), .b(s_308), .O(gate125inter1));
  and2  gate2705(.a(G403), .b(G402), .O(gate125inter2));
  inv1  gate2706(.a(s_308), .O(gate125inter3));
  inv1  gate2707(.a(s_309), .O(gate125inter4));
  nand2 gate2708(.a(gate125inter4), .b(gate125inter3), .O(gate125inter5));
  nor2  gate2709(.a(gate125inter5), .b(gate125inter2), .O(gate125inter6));
  inv1  gate2710(.a(G402), .O(gate125inter7));
  inv1  gate2711(.a(G403), .O(gate125inter8));
  nand2 gate2712(.a(gate125inter8), .b(gate125inter7), .O(gate125inter9));
  nand2 gate2713(.a(s_309), .b(gate125inter3), .O(gate125inter10));
  nor2  gate2714(.a(gate125inter10), .b(gate125inter9), .O(gate125inter11));
  nor2  gate2715(.a(gate125inter11), .b(gate125inter6), .O(gate125inter12));
  nand2 gate2716(.a(gate125inter12), .b(gate125inter1), .O(G486));
nand2 gate126( .a(G404), .b(G405), .O(G489) );
nand2 gate127( .a(G406), .b(G407), .O(G492) );

  xor2  gate1723(.a(G409), .b(G408), .O(gate128inter0));
  nand2 gate1724(.a(gate128inter0), .b(s_168), .O(gate128inter1));
  and2  gate1725(.a(G409), .b(G408), .O(gate128inter2));
  inv1  gate1726(.a(s_168), .O(gate128inter3));
  inv1  gate1727(.a(s_169), .O(gate128inter4));
  nand2 gate1728(.a(gate128inter4), .b(gate128inter3), .O(gate128inter5));
  nor2  gate1729(.a(gate128inter5), .b(gate128inter2), .O(gate128inter6));
  inv1  gate1730(.a(G408), .O(gate128inter7));
  inv1  gate1731(.a(G409), .O(gate128inter8));
  nand2 gate1732(.a(gate128inter8), .b(gate128inter7), .O(gate128inter9));
  nand2 gate1733(.a(s_169), .b(gate128inter3), .O(gate128inter10));
  nor2  gate1734(.a(gate128inter10), .b(gate128inter9), .O(gate128inter11));
  nor2  gate1735(.a(gate128inter11), .b(gate128inter6), .O(gate128inter12));
  nand2 gate1736(.a(gate128inter12), .b(gate128inter1), .O(G495));
nand2 gate129( .a(G410), .b(G411), .O(G498) );
nand2 gate130( .a(G412), .b(G413), .O(G501) );
nand2 gate131( .a(G414), .b(G415), .O(G504) );

  xor2  gate2171(.a(G417), .b(G416), .O(gate132inter0));
  nand2 gate2172(.a(gate132inter0), .b(s_232), .O(gate132inter1));
  and2  gate2173(.a(G417), .b(G416), .O(gate132inter2));
  inv1  gate2174(.a(s_232), .O(gate132inter3));
  inv1  gate2175(.a(s_233), .O(gate132inter4));
  nand2 gate2176(.a(gate132inter4), .b(gate132inter3), .O(gate132inter5));
  nor2  gate2177(.a(gate132inter5), .b(gate132inter2), .O(gate132inter6));
  inv1  gate2178(.a(G416), .O(gate132inter7));
  inv1  gate2179(.a(G417), .O(gate132inter8));
  nand2 gate2180(.a(gate132inter8), .b(gate132inter7), .O(gate132inter9));
  nand2 gate2181(.a(s_233), .b(gate132inter3), .O(gate132inter10));
  nor2  gate2182(.a(gate132inter10), .b(gate132inter9), .O(gate132inter11));
  nor2  gate2183(.a(gate132inter11), .b(gate132inter6), .O(gate132inter12));
  nand2 gate2184(.a(gate132inter12), .b(gate132inter1), .O(G507));
nand2 gate133( .a(G418), .b(G419), .O(G510) );

  xor2  gate1905(.a(G421), .b(G420), .O(gate134inter0));
  nand2 gate1906(.a(gate134inter0), .b(s_194), .O(gate134inter1));
  and2  gate1907(.a(G421), .b(G420), .O(gate134inter2));
  inv1  gate1908(.a(s_194), .O(gate134inter3));
  inv1  gate1909(.a(s_195), .O(gate134inter4));
  nand2 gate1910(.a(gate134inter4), .b(gate134inter3), .O(gate134inter5));
  nor2  gate1911(.a(gate134inter5), .b(gate134inter2), .O(gate134inter6));
  inv1  gate1912(.a(G420), .O(gate134inter7));
  inv1  gate1913(.a(G421), .O(gate134inter8));
  nand2 gate1914(.a(gate134inter8), .b(gate134inter7), .O(gate134inter9));
  nand2 gate1915(.a(s_195), .b(gate134inter3), .O(gate134inter10));
  nor2  gate1916(.a(gate134inter10), .b(gate134inter9), .O(gate134inter11));
  nor2  gate1917(.a(gate134inter11), .b(gate134inter6), .O(gate134inter12));
  nand2 gate1918(.a(gate134inter12), .b(gate134inter1), .O(G513));
nand2 gate135( .a(G422), .b(G423), .O(G516) );

  xor2  gate2283(.a(G425), .b(G424), .O(gate136inter0));
  nand2 gate2284(.a(gate136inter0), .b(s_248), .O(gate136inter1));
  and2  gate2285(.a(G425), .b(G424), .O(gate136inter2));
  inv1  gate2286(.a(s_248), .O(gate136inter3));
  inv1  gate2287(.a(s_249), .O(gate136inter4));
  nand2 gate2288(.a(gate136inter4), .b(gate136inter3), .O(gate136inter5));
  nor2  gate2289(.a(gate136inter5), .b(gate136inter2), .O(gate136inter6));
  inv1  gate2290(.a(G424), .O(gate136inter7));
  inv1  gate2291(.a(G425), .O(gate136inter8));
  nand2 gate2292(.a(gate136inter8), .b(gate136inter7), .O(gate136inter9));
  nand2 gate2293(.a(s_249), .b(gate136inter3), .O(gate136inter10));
  nor2  gate2294(.a(gate136inter10), .b(gate136inter9), .O(gate136inter11));
  nor2  gate2295(.a(gate136inter11), .b(gate136inter6), .O(gate136inter12));
  nand2 gate2296(.a(gate136inter12), .b(gate136inter1), .O(G519));

  xor2  gate1611(.a(G429), .b(G426), .O(gate137inter0));
  nand2 gate1612(.a(gate137inter0), .b(s_152), .O(gate137inter1));
  and2  gate1613(.a(G429), .b(G426), .O(gate137inter2));
  inv1  gate1614(.a(s_152), .O(gate137inter3));
  inv1  gate1615(.a(s_153), .O(gate137inter4));
  nand2 gate1616(.a(gate137inter4), .b(gate137inter3), .O(gate137inter5));
  nor2  gate1617(.a(gate137inter5), .b(gate137inter2), .O(gate137inter6));
  inv1  gate1618(.a(G426), .O(gate137inter7));
  inv1  gate1619(.a(G429), .O(gate137inter8));
  nand2 gate1620(.a(gate137inter8), .b(gate137inter7), .O(gate137inter9));
  nand2 gate1621(.a(s_153), .b(gate137inter3), .O(gate137inter10));
  nor2  gate1622(.a(gate137inter10), .b(gate137inter9), .O(gate137inter11));
  nor2  gate1623(.a(gate137inter11), .b(gate137inter6), .O(gate137inter12));
  nand2 gate1624(.a(gate137inter12), .b(gate137inter1), .O(G522));
nand2 gate138( .a(G432), .b(G435), .O(G525) );
nand2 gate139( .a(G438), .b(G441), .O(G528) );

  xor2  gate1163(.a(G447), .b(G444), .O(gate140inter0));
  nand2 gate1164(.a(gate140inter0), .b(s_88), .O(gate140inter1));
  and2  gate1165(.a(G447), .b(G444), .O(gate140inter2));
  inv1  gate1166(.a(s_88), .O(gate140inter3));
  inv1  gate1167(.a(s_89), .O(gate140inter4));
  nand2 gate1168(.a(gate140inter4), .b(gate140inter3), .O(gate140inter5));
  nor2  gate1169(.a(gate140inter5), .b(gate140inter2), .O(gate140inter6));
  inv1  gate1170(.a(G444), .O(gate140inter7));
  inv1  gate1171(.a(G447), .O(gate140inter8));
  nand2 gate1172(.a(gate140inter8), .b(gate140inter7), .O(gate140inter9));
  nand2 gate1173(.a(s_89), .b(gate140inter3), .O(gate140inter10));
  nor2  gate1174(.a(gate140inter10), .b(gate140inter9), .O(gate140inter11));
  nor2  gate1175(.a(gate140inter11), .b(gate140inter6), .O(gate140inter12));
  nand2 gate1176(.a(gate140inter12), .b(gate140inter1), .O(G531));
nand2 gate141( .a(G450), .b(G453), .O(G534) );
nand2 gate142( .a(G456), .b(G459), .O(G537) );

  xor2  gate1667(.a(G465), .b(G462), .O(gate143inter0));
  nand2 gate1668(.a(gate143inter0), .b(s_160), .O(gate143inter1));
  and2  gate1669(.a(G465), .b(G462), .O(gate143inter2));
  inv1  gate1670(.a(s_160), .O(gate143inter3));
  inv1  gate1671(.a(s_161), .O(gate143inter4));
  nand2 gate1672(.a(gate143inter4), .b(gate143inter3), .O(gate143inter5));
  nor2  gate1673(.a(gate143inter5), .b(gate143inter2), .O(gate143inter6));
  inv1  gate1674(.a(G462), .O(gate143inter7));
  inv1  gate1675(.a(G465), .O(gate143inter8));
  nand2 gate1676(.a(gate143inter8), .b(gate143inter7), .O(gate143inter9));
  nand2 gate1677(.a(s_161), .b(gate143inter3), .O(gate143inter10));
  nor2  gate1678(.a(gate143inter10), .b(gate143inter9), .O(gate143inter11));
  nor2  gate1679(.a(gate143inter11), .b(gate143inter6), .O(gate143inter12));
  nand2 gate1680(.a(gate143inter12), .b(gate143inter1), .O(G540));
nand2 gate144( .a(G468), .b(G471), .O(G543) );
nand2 gate145( .a(G474), .b(G477), .O(G546) );
nand2 gate146( .a(G480), .b(G483), .O(G549) );

  xor2  gate1093(.a(G489), .b(G486), .O(gate147inter0));
  nand2 gate1094(.a(gate147inter0), .b(s_78), .O(gate147inter1));
  and2  gate1095(.a(G489), .b(G486), .O(gate147inter2));
  inv1  gate1096(.a(s_78), .O(gate147inter3));
  inv1  gate1097(.a(s_79), .O(gate147inter4));
  nand2 gate1098(.a(gate147inter4), .b(gate147inter3), .O(gate147inter5));
  nor2  gate1099(.a(gate147inter5), .b(gate147inter2), .O(gate147inter6));
  inv1  gate1100(.a(G486), .O(gate147inter7));
  inv1  gate1101(.a(G489), .O(gate147inter8));
  nand2 gate1102(.a(gate147inter8), .b(gate147inter7), .O(gate147inter9));
  nand2 gate1103(.a(s_79), .b(gate147inter3), .O(gate147inter10));
  nor2  gate1104(.a(gate147inter10), .b(gate147inter9), .O(gate147inter11));
  nor2  gate1105(.a(gate147inter11), .b(gate147inter6), .O(gate147inter12));
  nand2 gate1106(.a(gate147inter12), .b(gate147inter1), .O(G552));

  xor2  gate1191(.a(G495), .b(G492), .O(gate148inter0));
  nand2 gate1192(.a(gate148inter0), .b(s_92), .O(gate148inter1));
  and2  gate1193(.a(G495), .b(G492), .O(gate148inter2));
  inv1  gate1194(.a(s_92), .O(gate148inter3));
  inv1  gate1195(.a(s_93), .O(gate148inter4));
  nand2 gate1196(.a(gate148inter4), .b(gate148inter3), .O(gate148inter5));
  nor2  gate1197(.a(gate148inter5), .b(gate148inter2), .O(gate148inter6));
  inv1  gate1198(.a(G492), .O(gate148inter7));
  inv1  gate1199(.a(G495), .O(gate148inter8));
  nand2 gate1200(.a(gate148inter8), .b(gate148inter7), .O(gate148inter9));
  nand2 gate1201(.a(s_93), .b(gate148inter3), .O(gate148inter10));
  nor2  gate1202(.a(gate148inter10), .b(gate148inter9), .O(gate148inter11));
  nor2  gate1203(.a(gate148inter11), .b(gate148inter6), .O(gate148inter12));
  nand2 gate1204(.a(gate148inter12), .b(gate148inter1), .O(G555));
nand2 gate149( .a(G498), .b(G501), .O(G558) );
nand2 gate150( .a(G504), .b(G507), .O(G561) );

  xor2  gate2213(.a(G513), .b(G510), .O(gate151inter0));
  nand2 gate2214(.a(gate151inter0), .b(s_238), .O(gate151inter1));
  and2  gate2215(.a(G513), .b(G510), .O(gate151inter2));
  inv1  gate2216(.a(s_238), .O(gate151inter3));
  inv1  gate2217(.a(s_239), .O(gate151inter4));
  nand2 gate2218(.a(gate151inter4), .b(gate151inter3), .O(gate151inter5));
  nor2  gate2219(.a(gate151inter5), .b(gate151inter2), .O(gate151inter6));
  inv1  gate2220(.a(G510), .O(gate151inter7));
  inv1  gate2221(.a(G513), .O(gate151inter8));
  nand2 gate2222(.a(gate151inter8), .b(gate151inter7), .O(gate151inter9));
  nand2 gate2223(.a(s_239), .b(gate151inter3), .O(gate151inter10));
  nor2  gate2224(.a(gate151inter10), .b(gate151inter9), .O(gate151inter11));
  nor2  gate2225(.a(gate151inter11), .b(gate151inter6), .O(gate151inter12));
  nand2 gate2226(.a(gate151inter12), .b(gate151inter1), .O(G564));
nand2 gate152( .a(G516), .b(G519), .O(G567) );
nand2 gate153( .a(G426), .b(G522), .O(G570) );
nand2 gate154( .a(G429), .b(G522), .O(G571) );

  xor2  gate1877(.a(G525), .b(G432), .O(gate155inter0));
  nand2 gate1878(.a(gate155inter0), .b(s_190), .O(gate155inter1));
  and2  gate1879(.a(G525), .b(G432), .O(gate155inter2));
  inv1  gate1880(.a(s_190), .O(gate155inter3));
  inv1  gate1881(.a(s_191), .O(gate155inter4));
  nand2 gate1882(.a(gate155inter4), .b(gate155inter3), .O(gate155inter5));
  nor2  gate1883(.a(gate155inter5), .b(gate155inter2), .O(gate155inter6));
  inv1  gate1884(.a(G432), .O(gate155inter7));
  inv1  gate1885(.a(G525), .O(gate155inter8));
  nand2 gate1886(.a(gate155inter8), .b(gate155inter7), .O(gate155inter9));
  nand2 gate1887(.a(s_191), .b(gate155inter3), .O(gate155inter10));
  nor2  gate1888(.a(gate155inter10), .b(gate155inter9), .O(gate155inter11));
  nor2  gate1889(.a(gate155inter11), .b(gate155inter6), .O(gate155inter12));
  nand2 gate1890(.a(gate155inter12), .b(gate155inter1), .O(G572));
nand2 gate156( .a(G435), .b(G525), .O(G573) );
nand2 gate157( .a(G438), .b(G528), .O(G574) );
nand2 gate158( .a(G441), .b(G528), .O(G575) );

  xor2  gate1261(.a(G531), .b(G444), .O(gate159inter0));
  nand2 gate1262(.a(gate159inter0), .b(s_102), .O(gate159inter1));
  and2  gate1263(.a(G531), .b(G444), .O(gate159inter2));
  inv1  gate1264(.a(s_102), .O(gate159inter3));
  inv1  gate1265(.a(s_103), .O(gate159inter4));
  nand2 gate1266(.a(gate159inter4), .b(gate159inter3), .O(gate159inter5));
  nor2  gate1267(.a(gate159inter5), .b(gate159inter2), .O(gate159inter6));
  inv1  gate1268(.a(G444), .O(gate159inter7));
  inv1  gate1269(.a(G531), .O(gate159inter8));
  nand2 gate1270(.a(gate159inter8), .b(gate159inter7), .O(gate159inter9));
  nand2 gate1271(.a(s_103), .b(gate159inter3), .O(gate159inter10));
  nor2  gate1272(.a(gate159inter10), .b(gate159inter9), .O(gate159inter11));
  nor2  gate1273(.a(gate159inter11), .b(gate159inter6), .O(gate159inter12));
  nand2 gate1274(.a(gate159inter12), .b(gate159inter1), .O(G576));

  xor2  gate2269(.a(G531), .b(G447), .O(gate160inter0));
  nand2 gate2270(.a(gate160inter0), .b(s_246), .O(gate160inter1));
  and2  gate2271(.a(G531), .b(G447), .O(gate160inter2));
  inv1  gate2272(.a(s_246), .O(gate160inter3));
  inv1  gate2273(.a(s_247), .O(gate160inter4));
  nand2 gate2274(.a(gate160inter4), .b(gate160inter3), .O(gate160inter5));
  nor2  gate2275(.a(gate160inter5), .b(gate160inter2), .O(gate160inter6));
  inv1  gate2276(.a(G447), .O(gate160inter7));
  inv1  gate2277(.a(G531), .O(gate160inter8));
  nand2 gate2278(.a(gate160inter8), .b(gate160inter7), .O(gate160inter9));
  nand2 gate2279(.a(s_247), .b(gate160inter3), .O(gate160inter10));
  nor2  gate2280(.a(gate160inter10), .b(gate160inter9), .O(gate160inter11));
  nor2  gate2281(.a(gate160inter11), .b(gate160inter6), .O(gate160inter12));
  nand2 gate2282(.a(gate160inter12), .b(gate160inter1), .O(G577));
nand2 gate161( .a(G450), .b(G534), .O(G578) );

  xor2  gate1751(.a(G534), .b(G453), .O(gate162inter0));
  nand2 gate1752(.a(gate162inter0), .b(s_172), .O(gate162inter1));
  and2  gate1753(.a(G534), .b(G453), .O(gate162inter2));
  inv1  gate1754(.a(s_172), .O(gate162inter3));
  inv1  gate1755(.a(s_173), .O(gate162inter4));
  nand2 gate1756(.a(gate162inter4), .b(gate162inter3), .O(gate162inter5));
  nor2  gate1757(.a(gate162inter5), .b(gate162inter2), .O(gate162inter6));
  inv1  gate1758(.a(G453), .O(gate162inter7));
  inv1  gate1759(.a(G534), .O(gate162inter8));
  nand2 gate1760(.a(gate162inter8), .b(gate162inter7), .O(gate162inter9));
  nand2 gate1761(.a(s_173), .b(gate162inter3), .O(gate162inter10));
  nor2  gate1762(.a(gate162inter10), .b(gate162inter9), .O(gate162inter11));
  nor2  gate1763(.a(gate162inter11), .b(gate162inter6), .O(gate162inter12));
  nand2 gate1764(.a(gate162inter12), .b(gate162inter1), .O(G579));

  xor2  gate1317(.a(G537), .b(G456), .O(gate163inter0));
  nand2 gate1318(.a(gate163inter0), .b(s_110), .O(gate163inter1));
  and2  gate1319(.a(G537), .b(G456), .O(gate163inter2));
  inv1  gate1320(.a(s_110), .O(gate163inter3));
  inv1  gate1321(.a(s_111), .O(gate163inter4));
  nand2 gate1322(.a(gate163inter4), .b(gate163inter3), .O(gate163inter5));
  nor2  gate1323(.a(gate163inter5), .b(gate163inter2), .O(gate163inter6));
  inv1  gate1324(.a(G456), .O(gate163inter7));
  inv1  gate1325(.a(G537), .O(gate163inter8));
  nand2 gate1326(.a(gate163inter8), .b(gate163inter7), .O(gate163inter9));
  nand2 gate1327(.a(s_111), .b(gate163inter3), .O(gate163inter10));
  nor2  gate1328(.a(gate163inter10), .b(gate163inter9), .O(gate163inter11));
  nor2  gate1329(.a(gate163inter11), .b(gate163inter6), .O(gate163inter12));
  nand2 gate1330(.a(gate163inter12), .b(gate163inter1), .O(G580));
nand2 gate164( .a(G459), .b(G537), .O(G581) );
nand2 gate165( .a(G462), .b(G540), .O(G582) );
nand2 gate166( .a(G465), .b(G540), .O(G583) );

  xor2  gate2563(.a(G543), .b(G468), .O(gate167inter0));
  nand2 gate2564(.a(gate167inter0), .b(s_288), .O(gate167inter1));
  and2  gate2565(.a(G543), .b(G468), .O(gate167inter2));
  inv1  gate2566(.a(s_288), .O(gate167inter3));
  inv1  gate2567(.a(s_289), .O(gate167inter4));
  nand2 gate2568(.a(gate167inter4), .b(gate167inter3), .O(gate167inter5));
  nor2  gate2569(.a(gate167inter5), .b(gate167inter2), .O(gate167inter6));
  inv1  gate2570(.a(G468), .O(gate167inter7));
  inv1  gate2571(.a(G543), .O(gate167inter8));
  nand2 gate2572(.a(gate167inter8), .b(gate167inter7), .O(gate167inter9));
  nand2 gate2573(.a(s_289), .b(gate167inter3), .O(gate167inter10));
  nor2  gate2574(.a(gate167inter10), .b(gate167inter9), .O(gate167inter11));
  nor2  gate2575(.a(gate167inter11), .b(gate167inter6), .O(gate167inter12));
  nand2 gate2576(.a(gate167inter12), .b(gate167inter1), .O(G584));

  xor2  gate1303(.a(G543), .b(G471), .O(gate168inter0));
  nand2 gate1304(.a(gate168inter0), .b(s_108), .O(gate168inter1));
  and2  gate1305(.a(G543), .b(G471), .O(gate168inter2));
  inv1  gate1306(.a(s_108), .O(gate168inter3));
  inv1  gate1307(.a(s_109), .O(gate168inter4));
  nand2 gate1308(.a(gate168inter4), .b(gate168inter3), .O(gate168inter5));
  nor2  gate1309(.a(gate168inter5), .b(gate168inter2), .O(gate168inter6));
  inv1  gate1310(.a(G471), .O(gate168inter7));
  inv1  gate1311(.a(G543), .O(gate168inter8));
  nand2 gate1312(.a(gate168inter8), .b(gate168inter7), .O(gate168inter9));
  nand2 gate1313(.a(s_109), .b(gate168inter3), .O(gate168inter10));
  nor2  gate1314(.a(gate168inter10), .b(gate168inter9), .O(gate168inter11));
  nor2  gate1315(.a(gate168inter11), .b(gate168inter6), .O(gate168inter12));
  nand2 gate1316(.a(gate168inter12), .b(gate168inter1), .O(G585));

  xor2  gate1289(.a(G546), .b(G474), .O(gate169inter0));
  nand2 gate1290(.a(gate169inter0), .b(s_106), .O(gate169inter1));
  and2  gate1291(.a(G546), .b(G474), .O(gate169inter2));
  inv1  gate1292(.a(s_106), .O(gate169inter3));
  inv1  gate1293(.a(s_107), .O(gate169inter4));
  nand2 gate1294(.a(gate169inter4), .b(gate169inter3), .O(gate169inter5));
  nor2  gate1295(.a(gate169inter5), .b(gate169inter2), .O(gate169inter6));
  inv1  gate1296(.a(G474), .O(gate169inter7));
  inv1  gate1297(.a(G546), .O(gate169inter8));
  nand2 gate1298(.a(gate169inter8), .b(gate169inter7), .O(gate169inter9));
  nand2 gate1299(.a(s_107), .b(gate169inter3), .O(gate169inter10));
  nor2  gate1300(.a(gate169inter10), .b(gate169inter9), .O(gate169inter11));
  nor2  gate1301(.a(gate169inter11), .b(gate169inter6), .O(gate169inter12));
  nand2 gate1302(.a(gate169inter12), .b(gate169inter1), .O(G586));
nand2 gate170( .a(G477), .b(G546), .O(G587) );

  xor2  gate2129(.a(G549), .b(G480), .O(gate171inter0));
  nand2 gate2130(.a(gate171inter0), .b(s_226), .O(gate171inter1));
  and2  gate2131(.a(G549), .b(G480), .O(gate171inter2));
  inv1  gate2132(.a(s_226), .O(gate171inter3));
  inv1  gate2133(.a(s_227), .O(gate171inter4));
  nand2 gate2134(.a(gate171inter4), .b(gate171inter3), .O(gate171inter5));
  nor2  gate2135(.a(gate171inter5), .b(gate171inter2), .O(gate171inter6));
  inv1  gate2136(.a(G480), .O(gate171inter7));
  inv1  gate2137(.a(G549), .O(gate171inter8));
  nand2 gate2138(.a(gate171inter8), .b(gate171inter7), .O(gate171inter9));
  nand2 gate2139(.a(s_227), .b(gate171inter3), .O(gate171inter10));
  nor2  gate2140(.a(gate171inter10), .b(gate171inter9), .O(gate171inter11));
  nor2  gate2141(.a(gate171inter11), .b(gate171inter6), .O(gate171inter12));
  nand2 gate2142(.a(gate171inter12), .b(gate171inter1), .O(G588));
nand2 gate172( .a(G483), .b(G549), .O(G589) );

  xor2  gate2409(.a(G552), .b(G486), .O(gate173inter0));
  nand2 gate2410(.a(gate173inter0), .b(s_266), .O(gate173inter1));
  and2  gate2411(.a(G552), .b(G486), .O(gate173inter2));
  inv1  gate2412(.a(s_266), .O(gate173inter3));
  inv1  gate2413(.a(s_267), .O(gate173inter4));
  nand2 gate2414(.a(gate173inter4), .b(gate173inter3), .O(gate173inter5));
  nor2  gate2415(.a(gate173inter5), .b(gate173inter2), .O(gate173inter6));
  inv1  gate2416(.a(G486), .O(gate173inter7));
  inv1  gate2417(.a(G552), .O(gate173inter8));
  nand2 gate2418(.a(gate173inter8), .b(gate173inter7), .O(gate173inter9));
  nand2 gate2419(.a(s_267), .b(gate173inter3), .O(gate173inter10));
  nor2  gate2420(.a(gate173inter10), .b(gate173inter9), .O(gate173inter11));
  nor2  gate2421(.a(gate173inter11), .b(gate173inter6), .O(gate173inter12));
  nand2 gate2422(.a(gate173inter12), .b(gate173inter1), .O(G590));

  xor2  gate1443(.a(G552), .b(G489), .O(gate174inter0));
  nand2 gate1444(.a(gate174inter0), .b(s_128), .O(gate174inter1));
  and2  gate1445(.a(G552), .b(G489), .O(gate174inter2));
  inv1  gate1446(.a(s_128), .O(gate174inter3));
  inv1  gate1447(.a(s_129), .O(gate174inter4));
  nand2 gate1448(.a(gate174inter4), .b(gate174inter3), .O(gate174inter5));
  nor2  gate1449(.a(gate174inter5), .b(gate174inter2), .O(gate174inter6));
  inv1  gate1450(.a(G489), .O(gate174inter7));
  inv1  gate1451(.a(G552), .O(gate174inter8));
  nand2 gate1452(.a(gate174inter8), .b(gate174inter7), .O(gate174inter9));
  nand2 gate1453(.a(s_129), .b(gate174inter3), .O(gate174inter10));
  nor2  gate1454(.a(gate174inter10), .b(gate174inter9), .O(gate174inter11));
  nor2  gate1455(.a(gate174inter11), .b(gate174inter6), .O(gate174inter12));
  nand2 gate1456(.a(gate174inter12), .b(gate174inter1), .O(G591));

  xor2  gate2101(.a(G555), .b(G492), .O(gate175inter0));
  nand2 gate2102(.a(gate175inter0), .b(s_222), .O(gate175inter1));
  and2  gate2103(.a(G555), .b(G492), .O(gate175inter2));
  inv1  gate2104(.a(s_222), .O(gate175inter3));
  inv1  gate2105(.a(s_223), .O(gate175inter4));
  nand2 gate2106(.a(gate175inter4), .b(gate175inter3), .O(gate175inter5));
  nor2  gate2107(.a(gate175inter5), .b(gate175inter2), .O(gate175inter6));
  inv1  gate2108(.a(G492), .O(gate175inter7));
  inv1  gate2109(.a(G555), .O(gate175inter8));
  nand2 gate2110(.a(gate175inter8), .b(gate175inter7), .O(gate175inter9));
  nand2 gate2111(.a(s_223), .b(gate175inter3), .O(gate175inter10));
  nor2  gate2112(.a(gate175inter10), .b(gate175inter9), .O(gate175inter11));
  nor2  gate2113(.a(gate175inter11), .b(gate175inter6), .O(gate175inter12));
  nand2 gate2114(.a(gate175inter12), .b(gate175inter1), .O(G592));
nand2 gate176( .a(G495), .b(G555), .O(G593) );

  xor2  gate2857(.a(G558), .b(G498), .O(gate177inter0));
  nand2 gate2858(.a(gate177inter0), .b(s_330), .O(gate177inter1));
  and2  gate2859(.a(G558), .b(G498), .O(gate177inter2));
  inv1  gate2860(.a(s_330), .O(gate177inter3));
  inv1  gate2861(.a(s_331), .O(gate177inter4));
  nand2 gate2862(.a(gate177inter4), .b(gate177inter3), .O(gate177inter5));
  nor2  gate2863(.a(gate177inter5), .b(gate177inter2), .O(gate177inter6));
  inv1  gate2864(.a(G498), .O(gate177inter7));
  inv1  gate2865(.a(G558), .O(gate177inter8));
  nand2 gate2866(.a(gate177inter8), .b(gate177inter7), .O(gate177inter9));
  nand2 gate2867(.a(s_331), .b(gate177inter3), .O(gate177inter10));
  nor2  gate2868(.a(gate177inter10), .b(gate177inter9), .O(gate177inter11));
  nor2  gate2869(.a(gate177inter11), .b(gate177inter6), .O(gate177inter12));
  nand2 gate2870(.a(gate177inter12), .b(gate177inter1), .O(G594));
nand2 gate178( .a(G501), .b(G558), .O(G595) );

  xor2  gate2017(.a(G561), .b(G504), .O(gate179inter0));
  nand2 gate2018(.a(gate179inter0), .b(s_210), .O(gate179inter1));
  and2  gate2019(.a(G561), .b(G504), .O(gate179inter2));
  inv1  gate2020(.a(s_210), .O(gate179inter3));
  inv1  gate2021(.a(s_211), .O(gate179inter4));
  nand2 gate2022(.a(gate179inter4), .b(gate179inter3), .O(gate179inter5));
  nor2  gate2023(.a(gate179inter5), .b(gate179inter2), .O(gate179inter6));
  inv1  gate2024(.a(G504), .O(gate179inter7));
  inv1  gate2025(.a(G561), .O(gate179inter8));
  nand2 gate2026(.a(gate179inter8), .b(gate179inter7), .O(gate179inter9));
  nand2 gate2027(.a(s_211), .b(gate179inter3), .O(gate179inter10));
  nor2  gate2028(.a(gate179inter10), .b(gate179inter9), .O(gate179inter11));
  nor2  gate2029(.a(gate179inter11), .b(gate179inter6), .O(gate179inter12));
  nand2 gate2030(.a(gate179inter12), .b(gate179inter1), .O(G596));
nand2 gate180( .a(G507), .b(G561), .O(G597) );

  xor2  gate2829(.a(G564), .b(G510), .O(gate181inter0));
  nand2 gate2830(.a(gate181inter0), .b(s_326), .O(gate181inter1));
  and2  gate2831(.a(G564), .b(G510), .O(gate181inter2));
  inv1  gate2832(.a(s_326), .O(gate181inter3));
  inv1  gate2833(.a(s_327), .O(gate181inter4));
  nand2 gate2834(.a(gate181inter4), .b(gate181inter3), .O(gate181inter5));
  nor2  gate2835(.a(gate181inter5), .b(gate181inter2), .O(gate181inter6));
  inv1  gate2836(.a(G510), .O(gate181inter7));
  inv1  gate2837(.a(G564), .O(gate181inter8));
  nand2 gate2838(.a(gate181inter8), .b(gate181inter7), .O(gate181inter9));
  nand2 gate2839(.a(s_327), .b(gate181inter3), .O(gate181inter10));
  nor2  gate2840(.a(gate181inter10), .b(gate181inter9), .O(gate181inter11));
  nor2  gate2841(.a(gate181inter11), .b(gate181inter6), .O(gate181inter12));
  nand2 gate2842(.a(gate181inter12), .b(gate181inter1), .O(G598));

  xor2  gate1779(.a(G564), .b(G513), .O(gate182inter0));
  nand2 gate1780(.a(gate182inter0), .b(s_176), .O(gate182inter1));
  and2  gate1781(.a(G564), .b(G513), .O(gate182inter2));
  inv1  gate1782(.a(s_176), .O(gate182inter3));
  inv1  gate1783(.a(s_177), .O(gate182inter4));
  nand2 gate1784(.a(gate182inter4), .b(gate182inter3), .O(gate182inter5));
  nor2  gate1785(.a(gate182inter5), .b(gate182inter2), .O(gate182inter6));
  inv1  gate1786(.a(G513), .O(gate182inter7));
  inv1  gate1787(.a(G564), .O(gate182inter8));
  nand2 gate1788(.a(gate182inter8), .b(gate182inter7), .O(gate182inter9));
  nand2 gate1789(.a(s_177), .b(gate182inter3), .O(gate182inter10));
  nor2  gate1790(.a(gate182inter10), .b(gate182inter9), .O(gate182inter11));
  nor2  gate1791(.a(gate182inter11), .b(gate182inter6), .O(gate182inter12));
  nand2 gate1792(.a(gate182inter12), .b(gate182inter1), .O(G599));

  xor2  gate1639(.a(G567), .b(G516), .O(gate183inter0));
  nand2 gate1640(.a(gate183inter0), .b(s_156), .O(gate183inter1));
  and2  gate1641(.a(G567), .b(G516), .O(gate183inter2));
  inv1  gate1642(.a(s_156), .O(gate183inter3));
  inv1  gate1643(.a(s_157), .O(gate183inter4));
  nand2 gate1644(.a(gate183inter4), .b(gate183inter3), .O(gate183inter5));
  nor2  gate1645(.a(gate183inter5), .b(gate183inter2), .O(gate183inter6));
  inv1  gate1646(.a(G516), .O(gate183inter7));
  inv1  gate1647(.a(G567), .O(gate183inter8));
  nand2 gate1648(.a(gate183inter8), .b(gate183inter7), .O(gate183inter9));
  nand2 gate1649(.a(s_157), .b(gate183inter3), .O(gate183inter10));
  nor2  gate1650(.a(gate183inter10), .b(gate183inter9), .O(gate183inter11));
  nor2  gate1651(.a(gate183inter11), .b(gate183inter6), .O(gate183inter12));
  nand2 gate1652(.a(gate183inter12), .b(gate183inter1), .O(G600));
nand2 gate184( .a(G519), .b(G567), .O(G601) );

  xor2  gate1695(.a(G571), .b(G570), .O(gate185inter0));
  nand2 gate1696(.a(gate185inter0), .b(s_164), .O(gate185inter1));
  and2  gate1697(.a(G571), .b(G570), .O(gate185inter2));
  inv1  gate1698(.a(s_164), .O(gate185inter3));
  inv1  gate1699(.a(s_165), .O(gate185inter4));
  nand2 gate1700(.a(gate185inter4), .b(gate185inter3), .O(gate185inter5));
  nor2  gate1701(.a(gate185inter5), .b(gate185inter2), .O(gate185inter6));
  inv1  gate1702(.a(G570), .O(gate185inter7));
  inv1  gate1703(.a(G571), .O(gate185inter8));
  nand2 gate1704(.a(gate185inter8), .b(gate185inter7), .O(gate185inter9));
  nand2 gate1705(.a(s_165), .b(gate185inter3), .O(gate185inter10));
  nor2  gate1706(.a(gate185inter10), .b(gate185inter9), .O(gate185inter11));
  nor2  gate1707(.a(gate185inter11), .b(gate185inter6), .O(gate185inter12));
  nand2 gate1708(.a(gate185inter12), .b(gate185inter1), .O(G602));
nand2 gate186( .a(G572), .b(G573), .O(G607) );

  xor2  gate673(.a(G575), .b(G574), .O(gate187inter0));
  nand2 gate674(.a(gate187inter0), .b(s_18), .O(gate187inter1));
  and2  gate675(.a(G575), .b(G574), .O(gate187inter2));
  inv1  gate676(.a(s_18), .O(gate187inter3));
  inv1  gate677(.a(s_19), .O(gate187inter4));
  nand2 gate678(.a(gate187inter4), .b(gate187inter3), .O(gate187inter5));
  nor2  gate679(.a(gate187inter5), .b(gate187inter2), .O(gate187inter6));
  inv1  gate680(.a(G574), .O(gate187inter7));
  inv1  gate681(.a(G575), .O(gate187inter8));
  nand2 gate682(.a(gate187inter8), .b(gate187inter7), .O(gate187inter9));
  nand2 gate683(.a(s_19), .b(gate187inter3), .O(gate187inter10));
  nor2  gate684(.a(gate187inter10), .b(gate187inter9), .O(gate187inter11));
  nor2  gate685(.a(gate187inter11), .b(gate187inter6), .O(gate187inter12));
  nand2 gate686(.a(gate187inter12), .b(gate187inter1), .O(G612));

  xor2  gate1527(.a(G577), .b(G576), .O(gate188inter0));
  nand2 gate1528(.a(gate188inter0), .b(s_140), .O(gate188inter1));
  and2  gate1529(.a(G577), .b(G576), .O(gate188inter2));
  inv1  gate1530(.a(s_140), .O(gate188inter3));
  inv1  gate1531(.a(s_141), .O(gate188inter4));
  nand2 gate1532(.a(gate188inter4), .b(gate188inter3), .O(gate188inter5));
  nor2  gate1533(.a(gate188inter5), .b(gate188inter2), .O(gate188inter6));
  inv1  gate1534(.a(G576), .O(gate188inter7));
  inv1  gate1535(.a(G577), .O(gate188inter8));
  nand2 gate1536(.a(gate188inter8), .b(gate188inter7), .O(gate188inter9));
  nand2 gate1537(.a(s_141), .b(gate188inter3), .O(gate188inter10));
  nor2  gate1538(.a(gate188inter10), .b(gate188inter9), .O(gate188inter11));
  nor2  gate1539(.a(gate188inter11), .b(gate188inter6), .O(gate188inter12));
  nand2 gate1540(.a(gate188inter12), .b(gate188inter1), .O(G617));
nand2 gate189( .a(G578), .b(G579), .O(G622) );
nand2 gate190( .a(G580), .b(G581), .O(G627) );

  xor2  gate967(.a(G583), .b(G582), .O(gate191inter0));
  nand2 gate968(.a(gate191inter0), .b(s_60), .O(gate191inter1));
  and2  gate969(.a(G583), .b(G582), .O(gate191inter2));
  inv1  gate970(.a(s_60), .O(gate191inter3));
  inv1  gate971(.a(s_61), .O(gate191inter4));
  nand2 gate972(.a(gate191inter4), .b(gate191inter3), .O(gate191inter5));
  nor2  gate973(.a(gate191inter5), .b(gate191inter2), .O(gate191inter6));
  inv1  gate974(.a(G582), .O(gate191inter7));
  inv1  gate975(.a(G583), .O(gate191inter8));
  nand2 gate976(.a(gate191inter8), .b(gate191inter7), .O(gate191inter9));
  nand2 gate977(.a(s_61), .b(gate191inter3), .O(gate191inter10));
  nor2  gate978(.a(gate191inter10), .b(gate191inter9), .O(gate191inter11));
  nor2  gate979(.a(gate191inter11), .b(gate191inter6), .O(gate191inter12));
  nand2 gate980(.a(gate191inter12), .b(gate191inter1), .O(G632));
nand2 gate192( .a(G584), .b(G585), .O(G637) );
nand2 gate193( .a(G586), .b(G587), .O(G642) );
nand2 gate194( .a(G588), .b(G589), .O(G645) );
nand2 gate195( .a(G590), .b(G591), .O(G648) );

  xor2  gate547(.a(G593), .b(G592), .O(gate196inter0));
  nand2 gate548(.a(gate196inter0), .b(s_0), .O(gate196inter1));
  and2  gate549(.a(G593), .b(G592), .O(gate196inter2));
  inv1  gate550(.a(s_0), .O(gate196inter3));
  inv1  gate551(.a(s_1), .O(gate196inter4));
  nand2 gate552(.a(gate196inter4), .b(gate196inter3), .O(gate196inter5));
  nor2  gate553(.a(gate196inter5), .b(gate196inter2), .O(gate196inter6));
  inv1  gate554(.a(G592), .O(gate196inter7));
  inv1  gate555(.a(G593), .O(gate196inter8));
  nand2 gate556(.a(gate196inter8), .b(gate196inter7), .O(gate196inter9));
  nand2 gate557(.a(s_1), .b(gate196inter3), .O(gate196inter10));
  nor2  gate558(.a(gate196inter10), .b(gate196inter9), .O(gate196inter11));
  nor2  gate559(.a(gate196inter11), .b(gate196inter6), .O(gate196inter12));
  nand2 gate560(.a(gate196inter12), .b(gate196inter1), .O(G651));

  xor2  gate1359(.a(G595), .b(G594), .O(gate197inter0));
  nand2 gate1360(.a(gate197inter0), .b(s_116), .O(gate197inter1));
  and2  gate1361(.a(G595), .b(G594), .O(gate197inter2));
  inv1  gate1362(.a(s_116), .O(gate197inter3));
  inv1  gate1363(.a(s_117), .O(gate197inter4));
  nand2 gate1364(.a(gate197inter4), .b(gate197inter3), .O(gate197inter5));
  nor2  gate1365(.a(gate197inter5), .b(gate197inter2), .O(gate197inter6));
  inv1  gate1366(.a(G594), .O(gate197inter7));
  inv1  gate1367(.a(G595), .O(gate197inter8));
  nand2 gate1368(.a(gate197inter8), .b(gate197inter7), .O(gate197inter9));
  nand2 gate1369(.a(s_117), .b(gate197inter3), .O(gate197inter10));
  nor2  gate1370(.a(gate197inter10), .b(gate197inter9), .O(gate197inter11));
  nor2  gate1371(.a(gate197inter11), .b(gate197inter6), .O(gate197inter12));
  nand2 gate1372(.a(gate197inter12), .b(gate197inter1), .O(G654));

  xor2  gate1373(.a(G597), .b(G596), .O(gate198inter0));
  nand2 gate1374(.a(gate198inter0), .b(s_118), .O(gate198inter1));
  and2  gate1375(.a(G597), .b(G596), .O(gate198inter2));
  inv1  gate1376(.a(s_118), .O(gate198inter3));
  inv1  gate1377(.a(s_119), .O(gate198inter4));
  nand2 gate1378(.a(gate198inter4), .b(gate198inter3), .O(gate198inter5));
  nor2  gate1379(.a(gate198inter5), .b(gate198inter2), .O(gate198inter6));
  inv1  gate1380(.a(G596), .O(gate198inter7));
  inv1  gate1381(.a(G597), .O(gate198inter8));
  nand2 gate1382(.a(gate198inter8), .b(gate198inter7), .O(gate198inter9));
  nand2 gate1383(.a(s_119), .b(gate198inter3), .O(gate198inter10));
  nor2  gate1384(.a(gate198inter10), .b(gate198inter9), .O(gate198inter11));
  nor2  gate1385(.a(gate198inter11), .b(gate198inter6), .O(gate198inter12));
  nand2 gate1386(.a(gate198inter12), .b(gate198inter1), .O(G657));

  xor2  gate2773(.a(G599), .b(G598), .O(gate199inter0));
  nand2 gate2774(.a(gate199inter0), .b(s_318), .O(gate199inter1));
  and2  gate2775(.a(G599), .b(G598), .O(gate199inter2));
  inv1  gate2776(.a(s_318), .O(gate199inter3));
  inv1  gate2777(.a(s_319), .O(gate199inter4));
  nand2 gate2778(.a(gate199inter4), .b(gate199inter3), .O(gate199inter5));
  nor2  gate2779(.a(gate199inter5), .b(gate199inter2), .O(gate199inter6));
  inv1  gate2780(.a(G598), .O(gate199inter7));
  inv1  gate2781(.a(G599), .O(gate199inter8));
  nand2 gate2782(.a(gate199inter8), .b(gate199inter7), .O(gate199inter9));
  nand2 gate2783(.a(s_319), .b(gate199inter3), .O(gate199inter10));
  nor2  gate2784(.a(gate199inter10), .b(gate199inter9), .O(gate199inter11));
  nor2  gate2785(.a(gate199inter11), .b(gate199inter6), .O(gate199inter12));
  nand2 gate2786(.a(gate199inter12), .b(gate199inter1), .O(G660));
nand2 gate200( .a(G600), .b(G601), .O(G663) );

  xor2  gate1793(.a(G607), .b(G602), .O(gate201inter0));
  nand2 gate1794(.a(gate201inter0), .b(s_178), .O(gate201inter1));
  and2  gate1795(.a(G607), .b(G602), .O(gate201inter2));
  inv1  gate1796(.a(s_178), .O(gate201inter3));
  inv1  gate1797(.a(s_179), .O(gate201inter4));
  nand2 gate1798(.a(gate201inter4), .b(gate201inter3), .O(gate201inter5));
  nor2  gate1799(.a(gate201inter5), .b(gate201inter2), .O(gate201inter6));
  inv1  gate1800(.a(G602), .O(gate201inter7));
  inv1  gate1801(.a(G607), .O(gate201inter8));
  nand2 gate1802(.a(gate201inter8), .b(gate201inter7), .O(gate201inter9));
  nand2 gate1803(.a(s_179), .b(gate201inter3), .O(gate201inter10));
  nor2  gate1804(.a(gate201inter10), .b(gate201inter9), .O(gate201inter11));
  nor2  gate1805(.a(gate201inter11), .b(gate201inter6), .O(gate201inter12));
  nand2 gate1806(.a(gate201inter12), .b(gate201inter1), .O(G666));
nand2 gate202( .a(G612), .b(G617), .O(G669) );

  xor2  gate1107(.a(G612), .b(G602), .O(gate203inter0));
  nand2 gate1108(.a(gate203inter0), .b(s_80), .O(gate203inter1));
  and2  gate1109(.a(G612), .b(G602), .O(gate203inter2));
  inv1  gate1110(.a(s_80), .O(gate203inter3));
  inv1  gate1111(.a(s_81), .O(gate203inter4));
  nand2 gate1112(.a(gate203inter4), .b(gate203inter3), .O(gate203inter5));
  nor2  gate1113(.a(gate203inter5), .b(gate203inter2), .O(gate203inter6));
  inv1  gate1114(.a(G602), .O(gate203inter7));
  inv1  gate1115(.a(G612), .O(gate203inter8));
  nand2 gate1116(.a(gate203inter8), .b(gate203inter7), .O(gate203inter9));
  nand2 gate1117(.a(s_81), .b(gate203inter3), .O(gate203inter10));
  nor2  gate1118(.a(gate203inter10), .b(gate203inter9), .O(gate203inter11));
  nor2  gate1119(.a(gate203inter11), .b(gate203inter6), .O(gate203inter12));
  nand2 gate1120(.a(gate203inter12), .b(gate203inter1), .O(G672));
nand2 gate204( .a(G607), .b(G617), .O(G675) );

  xor2  gate785(.a(G627), .b(G622), .O(gate205inter0));
  nand2 gate786(.a(gate205inter0), .b(s_34), .O(gate205inter1));
  and2  gate787(.a(G627), .b(G622), .O(gate205inter2));
  inv1  gate788(.a(s_34), .O(gate205inter3));
  inv1  gate789(.a(s_35), .O(gate205inter4));
  nand2 gate790(.a(gate205inter4), .b(gate205inter3), .O(gate205inter5));
  nor2  gate791(.a(gate205inter5), .b(gate205inter2), .O(gate205inter6));
  inv1  gate792(.a(G622), .O(gate205inter7));
  inv1  gate793(.a(G627), .O(gate205inter8));
  nand2 gate794(.a(gate205inter8), .b(gate205inter7), .O(gate205inter9));
  nand2 gate795(.a(s_35), .b(gate205inter3), .O(gate205inter10));
  nor2  gate796(.a(gate205inter10), .b(gate205inter9), .O(gate205inter11));
  nor2  gate797(.a(gate205inter11), .b(gate205inter6), .O(gate205inter12));
  nand2 gate798(.a(gate205inter12), .b(gate205inter1), .O(G678));

  xor2  gate2521(.a(G637), .b(G632), .O(gate206inter0));
  nand2 gate2522(.a(gate206inter0), .b(s_282), .O(gate206inter1));
  and2  gate2523(.a(G637), .b(G632), .O(gate206inter2));
  inv1  gate2524(.a(s_282), .O(gate206inter3));
  inv1  gate2525(.a(s_283), .O(gate206inter4));
  nand2 gate2526(.a(gate206inter4), .b(gate206inter3), .O(gate206inter5));
  nor2  gate2527(.a(gate206inter5), .b(gate206inter2), .O(gate206inter6));
  inv1  gate2528(.a(G632), .O(gate206inter7));
  inv1  gate2529(.a(G637), .O(gate206inter8));
  nand2 gate2530(.a(gate206inter8), .b(gate206inter7), .O(gate206inter9));
  nand2 gate2531(.a(s_283), .b(gate206inter3), .O(gate206inter10));
  nor2  gate2532(.a(gate206inter10), .b(gate206inter9), .O(gate206inter11));
  nor2  gate2533(.a(gate206inter11), .b(gate206inter6), .O(gate206inter12));
  nand2 gate2534(.a(gate206inter12), .b(gate206inter1), .O(G681));
nand2 gate207( .a(G622), .b(G632), .O(G684) );

  xor2  gate757(.a(G637), .b(G627), .O(gate208inter0));
  nand2 gate758(.a(gate208inter0), .b(s_30), .O(gate208inter1));
  and2  gate759(.a(G637), .b(G627), .O(gate208inter2));
  inv1  gate760(.a(s_30), .O(gate208inter3));
  inv1  gate761(.a(s_31), .O(gate208inter4));
  nand2 gate762(.a(gate208inter4), .b(gate208inter3), .O(gate208inter5));
  nor2  gate763(.a(gate208inter5), .b(gate208inter2), .O(gate208inter6));
  inv1  gate764(.a(G627), .O(gate208inter7));
  inv1  gate765(.a(G637), .O(gate208inter8));
  nand2 gate766(.a(gate208inter8), .b(gate208inter7), .O(gate208inter9));
  nand2 gate767(.a(s_31), .b(gate208inter3), .O(gate208inter10));
  nor2  gate768(.a(gate208inter10), .b(gate208inter9), .O(gate208inter11));
  nor2  gate769(.a(gate208inter11), .b(gate208inter6), .O(gate208inter12));
  nand2 gate770(.a(gate208inter12), .b(gate208inter1), .O(G687));

  xor2  gate2661(.a(G666), .b(G602), .O(gate209inter0));
  nand2 gate2662(.a(gate209inter0), .b(s_302), .O(gate209inter1));
  and2  gate2663(.a(G666), .b(G602), .O(gate209inter2));
  inv1  gate2664(.a(s_302), .O(gate209inter3));
  inv1  gate2665(.a(s_303), .O(gate209inter4));
  nand2 gate2666(.a(gate209inter4), .b(gate209inter3), .O(gate209inter5));
  nor2  gate2667(.a(gate209inter5), .b(gate209inter2), .O(gate209inter6));
  inv1  gate2668(.a(G602), .O(gate209inter7));
  inv1  gate2669(.a(G666), .O(gate209inter8));
  nand2 gate2670(.a(gate209inter8), .b(gate209inter7), .O(gate209inter9));
  nand2 gate2671(.a(s_303), .b(gate209inter3), .O(gate209inter10));
  nor2  gate2672(.a(gate209inter10), .b(gate209inter9), .O(gate209inter11));
  nor2  gate2673(.a(gate209inter11), .b(gate209inter6), .O(gate209inter12));
  nand2 gate2674(.a(gate209inter12), .b(gate209inter1), .O(G690));

  xor2  gate2759(.a(G666), .b(G607), .O(gate210inter0));
  nand2 gate2760(.a(gate210inter0), .b(s_316), .O(gate210inter1));
  and2  gate2761(.a(G666), .b(G607), .O(gate210inter2));
  inv1  gate2762(.a(s_316), .O(gate210inter3));
  inv1  gate2763(.a(s_317), .O(gate210inter4));
  nand2 gate2764(.a(gate210inter4), .b(gate210inter3), .O(gate210inter5));
  nor2  gate2765(.a(gate210inter5), .b(gate210inter2), .O(gate210inter6));
  inv1  gate2766(.a(G607), .O(gate210inter7));
  inv1  gate2767(.a(G666), .O(gate210inter8));
  nand2 gate2768(.a(gate210inter8), .b(gate210inter7), .O(gate210inter9));
  nand2 gate2769(.a(s_317), .b(gate210inter3), .O(gate210inter10));
  nor2  gate2770(.a(gate210inter10), .b(gate210inter9), .O(gate210inter11));
  nor2  gate2771(.a(gate210inter11), .b(gate210inter6), .O(gate210inter12));
  nand2 gate2772(.a(gate210inter12), .b(gate210inter1), .O(G691));
nand2 gate211( .a(G612), .b(G669), .O(G692) );
nand2 gate212( .a(G617), .b(G669), .O(G693) );
nand2 gate213( .a(G602), .b(G672), .O(G694) );
nand2 gate214( .a(G612), .b(G672), .O(G695) );
nand2 gate215( .a(G607), .b(G675), .O(G696) );
nand2 gate216( .a(G617), .b(G675), .O(G697) );
nand2 gate217( .a(G622), .b(G678), .O(G698) );
nand2 gate218( .a(G627), .b(G678), .O(G699) );
nand2 gate219( .a(G632), .b(G681), .O(G700) );
nand2 gate220( .a(G637), .b(G681), .O(G701) );
nand2 gate221( .a(G622), .b(G684), .O(G702) );

  xor2  gate2927(.a(G684), .b(G632), .O(gate222inter0));
  nand2 gate2928(.a(gate222inter0), .b(s_340), .O(gate222inter1));
  and2  gate2929(.a(G684), .b(G632), .O(gate222inter2));
  inv1  gate2930(.a(s_340), .O(gate222inter3));
  inv1  gate2931(.a(s_341), .O(gate222inter4));
  nand2 gate2932(.a(gate222inter4), .b(gate222inter3), .O(gate222inter5));
  nor2  gate2933(.a(gate222inter5), .b(gate222inter2), .O(gate222inter6));
  inv1  gate2934(.a(G632), .O(gate222inter7));
  inv1  gate2935(.a(G684), .O(gate222inter8));
  nand2 gate2936(.a(gate222inter8), .b(gate222inter7), .O(gate222inter9));
  nand2 gate2937(.a(s_341), .b(gate222inter3), .O(gate222inter10));
  nor2  gate2938(.a(gate222inter10), .b(gate222inter9), .O(gate222inter11));
  nor2  gate2939(.a(gate222inter11), .b(gate222inter6), .O(gate222inter12));
  nand2 gate2940(.a(gate222inter12), .b(gate222inter1), .O(G703));

  xor2  gate1415(.a(G687), .b(G627), .O(gate223inter0));
  nand2 gate1416(.a(gate223inter0), .b(s_124), .O(gate223inter1));
  and2  gate1417(.a(G687), .b(G627), .O(gate223inter2));
  inv1  gate1418(.a(s_124), .O(gate223inter3));
  inv1  gate1419(.a(s_125), .O(gate223inter4));
  nand2 gate1420(.a(gate223inter4), .b(gate223inter3), .O(gate223inter5));
  nor2  gate1421(.a(gate223inter5), .b(gate223inter2), .O(gate223inter6));
  inv1  gate1422(.a(G627), .O(gate223inter7));
  inv1  gate1423(.a(G687), .O(gate223inter8));
  nand2 gate1424(.a(gate223inter8), .b(gate223inter7), .O(gate223inter9));
  nand2 gate1425(.a(s_125), .b(gate223inter3), .O(gate223inter10));
  nor2  gate1426(.a(gate223inter10), .b(gate223inter9), .O(gate223inter11));
  nor2  gate1427(.a(gate223inter11), .b(gate223inter6), .O(gate223inter12));
  nand2 gate1428(.a(gate223inter12), .b(gate223inter1), .O(G704));
nand2 gate224( .a(G637), .b(G687), .O(G705) );
nand2 gate225( .a(G690), .b(G691), .O(G706) );
nand2 gate226( .a(G692), .b(G693), .O(G709) );
nand2 gate227( .a(G694), .b(G695), .O(G712) );

  xor2  gate813(.a(G697), .b(G696), .O(gate228inter0));
  nand2 gate814(.a(gate228inter0), .b(s_38), .O(gate228inter1));
  and2  gate815(.a(G697), .b(G696), .O(gate228inter2));
  inv1  gate816(.a(s_38), .O(gate228inter3));
  inv1  gate817(.a(s_39), .O(gate228inter4));
  nand2 gate818(.a(gate228inter4), .b(gate228inter3), .O(gate228inter5));
  nor2  gate819(.a(gate228inter5), .b(gate228inter2), .O(gate228inter6));
  inv1  gate820(.a(G696), .O(gate228inter7));
  inv1  gate821(.a(G697), .O(gate228inter8));
  nand2 gate822(.a(gate228inter8), .b(gate228inter7), .O(gate228inter9));
  nand2 gate823(.a(s_39), .b(gate228inter3), .O(gate228inter10));
  nor2  gate824(.a(gate228inter10), .b(gate228inter9), .O(gate228inter11));
  nor2  gate825(.a(gate228inter11), .b(gate228inter6), .O(gate228inter12));
  nand2 gate826(.a(gate228inter12), .b(gate228inter1), .O(G715));

  xor2  gate1989(.a(G699), .b(G698), .O(gate229inter0));
  nand2 gate1990(.a(gate229inter0), .b(s_206), .O(gate229inter1));
  and2  gate1991(.a(G699), .b(G698), .O(gate229inter2));
  inv1  gate1992(.a(s_206), .O(gate229inter3));
  inv1  gate1993(.a(s_207), .O(gate229inter4));
  nand2 gate1994(.a(gate229inter4), .b(gate229inter3), .O(gate229inter5));
  nor2  gate1995(.a(gate229inter5), .b(gate229inter2), .O(gate229inter6));
  inv1  gate1996(.a(G698), .O(gate229inter7));
  inv1  gate1997(.a(G699), .O(gate229inter8));
  nand2 gate1998(.a(gate229inter8), .b(gate229inter7), .O(gate229inter9));
  nand2 gate1999(.a(s_207), .b(gate229inter3), .O(gate229inter10));
  nor2  gate2000(.a(gate229inter10), .b(gate229inter9), .O(gate229inter11));
  nor2  gate2001(.a(gate229inter11), .b(gate229inter6), .O(gate229inter12));
  nand2 gate2002(.a(gate229inter12), .b(gate229inter1), .O(G718));
nand2 gate230( .a(G700), .b(G701), .O(G721) );

  xor2  gate1009(.a(G703), .b(G702), .O(gate231inter0));
  nand2 gate1010(.a(gate231inter0), .b(s_66), .O(gate231inter1));
  and2  gate1011(.a(G703), .b(G702), .O(gate231inter2));
  inv1  gate1012(.a(s_66), .O(gate231inter3));
  inv1  gate1013(.a(s_67), .O(gate231inter4));
  nand2 gate1014(.a(gate231inter4), .b(gate231inter3), .O(gate231inter5));
  nor2  gate1015(.a(gate231inter5), .b(gate231inter2), .O(gate231inter6));
  inv1  gate1016(.a(G702), .O(gate231inter7));
  inv1  gate1017(.a(G703), .O(gate231inter8));
  nand2 gate1018(.a(gate231inter8), .b(gate231inter7), .O(gate231inter9));
  nand2 gate1019(.a(s_67), .b(gate231inter3), .O(gate231inter10));
  nor2  gate1020(.a(gate231inter10), .b(gate231inter9), .O(gate231inter11));
  nor2  gate1021(.a(gate231inter11), .b(gate231inter6), .O(gate231inter12));
  nand2 gate1022(.a(gate231inter12), .b(gate231inter1), .O(G724));
nand2 gate232( .a(G704), .b(G705), .O(G727) );
nand2 gate233( .a(G242), .b(G718), .O(G730) );

  xor2  gate603(.a(G721), .b(G245), .O(gate234inter0));
  nand2 gate604(.a(gate234inter0), .b(s_8), .O(gate234inter1));
  and2  gate605(.a(G721), .b(G245), .O(gate234inter2));
  inv1  gate606(.a(s_8), .O(gate234inter3));
  inv1  gate607(.a(s_9), .O(gate234inter4));
  nand2 gate608(.a(gate234inter4), .b(gate234inter3), .O(gate234inter5));
  nor2  gate609(.a(gate234inter5), .b(gate234inter2), .O(gate234inter6));
  inv1  gate610(.a(G245), .O(gate234inter7));
  inv1  gate611(.a(G721), .O(gate234inter8));
  nand2 gate612(.a(gate234inter8), .b(gate234inter7), .O(gate234inter9));
  nand2 gate613(.a(s_9), .b(gate234inter3), .O(gate234inter10));
  nor2  gate614(.a(gate234inter10), .b(gate234inter9), .O(gate234inter11));
  nor2  gate615(.a(gate234inter11), .b(gate234inter6), .O(gate234inter12));
  nand2 gate616(.a(gate234inter12), .b(gate234inter1), .O(G733));

  xor2  gate2451(.a(G724), .b(G248), .O(gate235inter0));
  nand2 gate2452(.a(gate235inter0), .b(s_272), .O(gate235inter1));
  and2  gate2453(.a(G724), .b(G248), .O(gate235inter2));
  inv1  gate2454(.a(s_272), .O(gate235inter3));
  inv1  gate2455(.a(s_273), .O(gate235inter4));
  nand2 gate2456(.a(gate235inter4), .b(gate235inter3), .O(gate235inter5));
  nor2  gate2457(.a(gate235inter5), .b(gate235inter2), .O(gate235inter6));
  inv1  gate2458(.a(G248), .O(gate235inter7));
  inv1  gate2459(.a(G724), .O(gate235inter8));
  nand2 gate2460(.a(gate235inter8), .b(gate235inter7), .O(gate235inter9));
  nand2 gate2461(.a(s_273), .b(gate235inter3), .O(gate235inter10));
  nor2  gate2462(.a(gate235inter10), .b(gate235inter9), .O(gate235inter11));
  nor2  gate2463(.a(gate235inter11), .b(gate235inter6), .O(gate235inter12));
  nand2 gate2464(.a(gate235inter12), .b(gate235inter1), .O(G736));
nand2 gate236( .a(G251), .b(G727), .O(G739) );
nand2 gate237( .a(G254), .b(G706), .O(G742) );
nand2 gate238( .a(G257), .b(G709), .O(G745) );
nand2 gate239( .a(G260), .b(G712), .O(G748) );
nand2 gate240( .a(G263), .b(G715), .O(G751) );
nand2 gate241( .a(G242), .b(G730), .O(G754) );
nand2 gate242( .a(G718), .b(G730), .O(G755) );

  xor2  gate827(.a(G733), .b(G245), .O(gate243inter0));
  nand2 gate828(.a(gate243inter0), .b(s_40), .O(gate243inter1));
  and2  gate829(.a(G733), .b(G245), .O(gate243inter2));
  inv1  gate830(.a(s_40), .O(gate243inter3));
  inv1  gate831(.a(s_41), .O(gate243inter4));
  nand2 gate832(.a(gate243inter4), .b(gate243inter3), .O(gate243inter5));
  nor2  gate833(.a(gate243inter5), .b(gate243inter2), .O(gate243inter6));
  inv1  gate834(.a(G245), .O(gate243inter7));
  inv1  gate835(.a(G733), .O(gate243inter8));
  nand2 gate836(.a(gate243inter8), .b(gate243inter7), .O(gate243inter9));
  nand2 gate837(.a(s_41), .b(gate243inter3), .O(gate243inter10));
  nor2  gate838(.a(gate243inter10), .b(gate243inter9), .O(gate243inter11));
  nor2  gate839(.a(gate243inter11), .b(gate243inter6), .O(gate243inter12));
  nand2 gate840(.a(gate243inter12), .b(gate243inter1), .O(G756));
nand2 gate244( .a(G721), .b(G733), .O(G757) );

  xor2  gate1121(.a(G736), .b(G248), .O(gate245inter0));
  nand2 gate1122(.a(gate245inter0), .b(s_82), .O(gate245inter1));
  and2  gate1123(.a(G736), .b(G248), .O(gate245inter2));
  inv1  gate1124(.a(s_82), .O(gate245inter3));
  inv1  gate1125(.a(s_83), .O(gate245inter4));
  nand2 gate1126(.a(gate245inter4), .b(gate245inter3), .O(gate245inter5));
  nor2  gate1127(.a(gate245inter5), .b(gate245inter2), .O(gate245inter6));
  inv1  gate1128(.a(G248), .O(gate245inter7));
  inv1  gate1129(.a(G736), .O(gate245inter8));
  nand2 gate1130(.a(gate245inter8), .b(gate245inter7), .O(gate245inter9));
  nand2 gate1131(.a(s_83), .b(gate245inter3), .O(gate245inter10));
  nor2  gate1132(.a(gate245inter10), .b(gate245inter9), .O(gate245inter11));
  nor2  gate1133(.a(gate245inter11), .b(gate245inter6), .O(gate245inter12));
  nand2 gate1134(.a(gate245inter12), .b(gate245inter1), .O(G758));
nand2 gate246( .a(G724), .b(G736), .O(G759) );

  xor2  gate2087(.a(G739), .b(G251), .O(gate247inter0));
  nand2 gate2088(.a(gate247inter0), .b(s_220), .O(gate247inter1));
  and2  gate2089(.a(G739), .b(G251), .O(gate247inter2));
  inv1  gate2090(.a(s_220), .O(gate247inter3));
  inv1  gate2091(.a(s_221), .O(gate247inter4));
  nand2 gate2092(.a(gate247inter4), .b(gate247inter3), .O(gate247inter5));
  nor2  gate2093(.a(gate247inter5), .b(gate247inter2), .O(gate247inter6));
  inv1  gate2094(.a(G251), .O(gate247inter7));
  inv1  gate2095(.a(G739), .O(gate247inter8));
  nand2 gate2096(.a(gate247inter8), .b(gate247inter7), .O(gate247inter9));
  nand2 gate2097(.a(s_221), .b(gate247inter3), .O(gate247inter10));
  nor2  gate2098(.a(gate247inter10), .b(gate247inter9), .O(gate247inter11));
  nor2  gate2099(.a(gate247inter11), .b(gate247inter6), .O(gate247inter12));
  nand2 gate2100(.a(gate247inter12), .b(gate247inter1), .O(G760));

  xor2  gate2465(.a(G739), .b(G727), .O(gate248inter0));
  nand2 gate2466(.a(gate248inter0), .b(s_274), .O(gate248inter1));
  and2  gate2467(.a(G739), .b(G727), .O(gate248inter2));
  inv1  gate2468(.a(s_274), .O(gate248inter3));
  inv1  gate2469(.a(s_275), .O(gate248inter4));
  nand2 gate2470(.a(gate248inter4), .b(gate248inter3), .O(gate248inter5));
  nor2  gate2471(.a(gate248inter5), .b(gate248inter2), .O(gate248inter6));
  inv1  gate2472(.a(G727), .O(gate248inter7));
  inv1  gate2473(.a(G739), .O(gate248inter8));
  nand2 gate2474(.a(gate248inter8), .b(gate248inter7), .O(gate248inter9));
  nand2 gate2475(.a(s_275), .b(gate248inter3), .O(gate248inter10));
  nor2  gate2476(.a(gate248inter10), .b(gate248inter9), .O(gate248inter11));
  nor2  gate2477(.a(gate248inter11), .b(gate248inter6), .O(gate248inter12));
  nand2 gate2478(.a(gate248inter12), .b(gate248inter1), .O(G761));
nand2 gate249( .a(G254), .b(G742), .O(G762) );

  xor2  gate1079(.a(G742), .b(G706), .O(gate250inter0));
  nand2 gate1080(.a(gate250inter0), .b(s_76), .O(gate250inter1));
  and2  gate1081(.a(G742), .b(G706), .O(gate250inter2));
  inv1  gate1082(.a(s_76), .O(gate250inter3));
  inv1  gate1083(.a(s_77), .O(gate250inter4));
  nand2 gate1084(.a(gate250inter4), .b(gate250inter3), .O(gate250inter5));
  nor2  gate1085(.a(gate250inter5), .b(gate250inter2), .O(gate250inter6));
  inv1  gate1086(.a(G706), .O(gate250inter7));
  inv1  gate1087(.a(G742), .O(gate250inter8));
  nand2 gate1088(.a(gate250inter8), .b(gate250inter7), .O(gate250inter9));
  nand2 gate1089(.a(s_77), .b(gate250inter3), .O(gate250inter10));
  nor2  gate1090(.a(gate250inter10), .b(gate250inter9), .O(gate250inter11));
  nor2  gate1091(.a(gate250inter11), .b(gate250inter6), .O(gate250inter12));
  nand2 gate1092(.a(gate250inter12), .b(gate250inter1), .O(G763));
nand2 gate251( .a(G257), .b(G745), .O(G764) );
nand2 gate252( .a(G709), .b(G745), .O(G765) );

  xor2  gate1863(.a(G748), .b(G260), .O(gate253inter0));
  nand2 gate1864(.a(gate253inter0), .b(s_188), .O(gate253inter1));
  and2  gate1865(.a(G748), .b(G260), .O(gate253inter2));
  inv1  gate1866(.a(s_188), .O(gate253inter3));
  inv1  gate1867(.a(s_189), .O(gate253inter4));
  nand2 gate1868(.a(gate253inter4), .b(gate253inter3), .O(gate253inter5));
  nor2  gate1869(.a(gate253inter5), .b(gate253inter2), .O(gate253inter6));
  inv1  gate1870(.a(G260), .O(gate253inter7));
  inv1  gate1871(.a(G748), .O(gate253inter8));
  nand2 gate1872(.a(gate253inter8), .b(gate253inter7), .O(gate253inter9));
  nand2 gate1873(.a(s_189), .b(gate253inter3), .O(gate253inter10));
  nor2  gate1874(.a(gate253inter10), .b(gate253inter9), .O(gate253inter11));
  nor2  gate1875(.a(gate253inter11), .b(gate253inter6), .O(gate253inter12));
  nand2 gate1876(.a(gate253inter12), .b(gate253inter1), .O(G766));

  xor2  gate2003(.a(G748), .b(G712), .O(gate254inter0));
  nand2 gate2004(.a(gate254inter0), .b(s_208), .O(gate254inter1));
  and2  gate2005(.a(G748), .b(G712), .O(gate254inter2));
  inv1  gate2006(.a(s_208), .O(gate254inter3));
  inv1  gate2007(.a(s_209), .O(gate254inter4));
  nand2 gate2008(.a(gate254inter4), .b(gate254inter3), .O(gate254inter5));
  nor2  gate2009(.a(gate254inter5), .b(gate254inter2), .O(gate254inter6));
  inv1  gate2010(.a(G712), .O(gate254inter7));
  inv1  gate2011(.a(G748), .O(gate254inter8));
  nand2 gate2012(.a(gate254inter8), .b(gate254inter7), .O(gate254inter9));
  nand2 gate2013(.a(s_209), .b(gate254inter3), .O(gate254inter10));
  nor2  gate2014(.a(gate254inter10), .b(gate254inter9), .O(gate254inter11));
  nor2  gate2015(.a(gate254inter11), .b(gate254inter6), .O(gate254inter12));
  nand2 gate2016(.a(gate254inter12), .b(gate254inter1), .O(G767));

  xor2  gate2115(.a(G751), .b(G263), .O(gate255inter0));
  nand2 gate2116(.a(gate255inter0), .b(s_224), .O(gate255inter1));
  and2  gate2117(.a(G751), .b(G263), .O(gate255inter2));
  inv1  gate2118(.a(s_224), .O(gate255inter3));
  inv1  gate2119(.a(s_225), .O(gate255inter4));
  nand2 gate2120(.a(gate255inter4), .b(gate255inter3), .O(gate255inter5));
  nor2  gate2121(.a(gate255inter5), .b(gate255inter2), .O(gate255inter6));
  inv1  gate2122(.a(G263), .O(gate255inter7));
  inv1  gate2123(.a(G751), .O(gate255inter8));
  nand2 gate2124(.a(gate255inter8), .b(gate255inter7), .O(gate255inter9));
  nand2 gate2125(.a(s_225), .b(gate255inter3), .O(gate255inter10));
  nor2  gate2126(.a(gate255inter10), .b(gate255inter9), .O(gate255inter11));
  nor2  gate2127(.a(gate255inter11), .b(gate255inter6), .O(gate255inter12));
  nand2 gate2128(.a(gate255inter12), .b(gate255inter1), .O(G768));

  xor2  gate883(.a(G751), .b(G715), .O(gate256inter0));
  nand2 gate884(.a(gate256inter0), .b(s_48), .O(gate256inter1));
  and2  gate885(.a(G751), .b(G715), .O(gate256inter2));
  inv1  gate886(.a(s_48), .O(gate256inter3));
  inv1  gate887(.a(s_49), .O(gate256inter4));
  nand2 gate888(.a(gate256inter4), .b(gate256inter3), .O(gate256inter5));
  nor2  gate889(.a(gate256inter5), .b(gate256inter2), .O(gate256inter6));
  inv1  gate890(.a(G715), .O(gate256inter7));
  inv1  gate891(.a(G751), .O(gate256inter8));
  nand2 gate892(.a(gate256inter8), .b(gate256inter7), .O(gate256inter9));
  nand2 gate893(.a(s_49), .b(gate256inter3), .O(gate256inter10));
  nor2  gate894(.a(gate256inter10), .b(gate256inter9), .O(gate256inter11));
  nor2  gate895(.a(gate256inter11), .b(gate256inter6), .O(gate256inter12));
  nand2 gate896(.a(gate256inter12), .b(gate256inter1), .O(G769));
nand2 gate257( .a(G754), .b(G755), .O(G770) );
nand2 gate258( .a(G756), .b(G757), .O(G773) );

  xor2  gate1891(.a(G759), .b(G758), .O(gate259inter0));
  nand2 gate1892(.a(gate259inter0), .b(s_192), .O(gate259inter1));
  and2  gate1893(.a(G759), .b(G758), .O(gate259inter2));
  inv1  gate1894(.a(s_192), .O(gate259inter3));
  inv1  gate1895(.a(s_193), .O(gate259inter4));
  nand2 gate1896(.a(gate259inter4), .b(gate259inter3), .O(gate259inter5));
  nor2  gate1897(.a(gate259inter5), .b(gate259inter2), .O(gate259inter6));
  inv1  gate1898(.a(G758), .O(gate259inter7));
  inv1  gate1899(.a(G759), .O(gate259inter8));
  nand2 gate1900(.a(gate259inter8), .b(gate259inter7), .O(gate259inter9));
  nand2 gate1901(.a(s_193), .b(gate259inter3), .O(gate259inter10));
  nor2  gate1902(.a(gate259inter10), .b(gate259inter9), .O(gate259inter11));
  nor2  gate1903(.a(gate259inter11), .b(gate259inter6), .O(gate259inter12));
  nand2 gate1904(.a(gate259inter12), .b(gate259inter1), .O(G776));
nand2 gate260( .a(G760), .b(G761), .O(G779) );

  xor2  gate2311(.a(G763), .b(G762), .O(gate261inter0));
  nand2 gate2312(.a(gate261inter0), .b(s_252), .O(gate261inter1));
  and2  gate2313(.a(G763), .b(G762), .O(gate261inter2));
  inv1  gate2314(.a(s_252), .O(gate261inter3));
  inv1  gate2315(.a(s_253), .O(gate261inter4));
  nand2 gate2316(.a(gate261inter4), .b(gate261inter3), .O(gate261inter5));
  nor2  gate2317(.a(gate261inter5), .b(gate261inter2), .O(gate261inter6));
  inv1  gate2318(.a(G762), .O(gate261inter7));
  inv1  gate2319(.a(G763), .O(gate261inter8));
  nand2 gate2320(.a(gate261inter8), .b(gate261inter7), .O(gate261inter9));
  nand2 gate2321(.a(s_253), .b(gate261inter3), .O(gate261inter10));
  nor2  gate2322(.a(gate261inter10), .b(gate261inter9), .O(gate261inter11));
  nor2  gate2323(.a(gate261inter11), .b(gate261inter6), .O(gate261inter12));
  nand2 gate2324(.a(gate261inter12), .b(gate261inter1), .O(G782));

  xor2  gate869(.a(G765), .b(G764), .O(gate262inter0));
  nand2 gate870(.a(gate262inter0), .b(s_46), .O(gate262inter1));
  and2  gate871(.a(G765), .b(G764), .O(gate262inter2));
  inv1  gate872(.a(s_46), .O(gate262inter3));
  inv1  gate873(.a(s_47), .O(gate262inter4));
  nand2 gate874(.a(gate262inter4), .b(gate262inter3), .O(gate262inter5));
  nor2  gate875(.a(gate262inter5), .b(gate262inter2), .O(gate262inter6));
  inv1  gate876(.a(G764), .O(gate262inter7));
  inv1  gate877(.a(G765), .O(gate262inter8));
  nand2 gate878(.a(gate262inter8), .b(gate262inter7), .O(gate262inter9));
  nand2 gate879(.a(s_47), .b(gate262inter3), .O(gate262inter10));
  nor2  gate880(.a(gate262inter10), .b(gate262inter9), .O(gate262inter11));
  nor2  gate881(.a(gate262inter11), .b(gate262inter6), .O(gate262inter12));
  nand2 gate882(.a(gate262inter12), .b(gate262inter1), .O(G785));

  xor2  gate1919(.a(G767), .b(G766), .O(gate263inter0));
  nand2 gate1920(.a(gate263inter0), .b(s_196), .O(gate263inter1));
  and2  gate1921(.a(G767), .b(G766), .O(gate263inter2));
  inv1  gate1922(.a(s_196), .O(gate263inter3));
  inv1  gate1923(.a(s_197), .O(gate263inter4));
  nand2 gate1924(.a(gate263inter4), .b(gate263inter3), .O(gate263inter5));
  nor2  gate1925(.a(gate263inter5), .b(gate263inter2), .O(gate263inter6));
  inv1  gate1926(.a(G766), .O(gate263inter7));
  inv1  gate1927(.a(G767), .O(gate263inter8));
  nand2 gate1928(.a(gate263inter8), .b(gate263inter7), .O(gate263inter9));
  nand2 gate1929(.a(s_197), .b(gate263inter3), .O(gate263inter10));
  nor2  gate1930(.a(gate263inter10), .b(gate263inter9), .O(gate263inter11));
  nor2  gate1931(.a(gate263inter11), .b(gate263inter6), .O(gate263inter12));
  nand2 gate1932(.a(gate263inter12), .b(gate263inter1), .O(G788));
nand2 gate264( .a(G768), .b(G769), .O(G791) );

  xor2  gate1401(.a(G770), .b(G642), .O(gate265inter0));
  nand2 gate1402(.a(gate265inter0), .b(s_122), .O(gate265inter1));
  and2  gate1403(.a(G770), .b(G642), .O(gate265inter2));
  inv1  gate1404(.a(s_122), .O(gate265inter3));
  inv1  gate1405(.a(s_123), .O(gate265inter4));
  nand2 gate1406(.a(gate265inter4), .b(gate265inter3), .O(gate265inter5));
  nor2  gate1407(.a(gate265inter5), .b(gate265inter2), .O(gate265inter6));
  inv1  gate1408(.a(G642), .O(gate265inter7));
  inv1  gate1409(.a(G770), .O(gate265inter8));
  nand2 gate1410(.a(gate265inter8), .b(gate265inter7), .O(gate265inter9));
  nand2 gate1411(.a(s_123), .b(gate265inter3), .O(gate265inter10));
  nor2  gate1412(.a(gate265inter10), .b(gate265inter9), .O(gate265inter11));
  nor2  gate1413(.a(gate265inter11), .b(gate265inter6), .O(gate265inter12));
  nand2 gate1414(.a(gate265inter12), .b(gate265inter1), .O(G794));

  xor2  gate687(.a(G773), .b(G645), .O(gate266inter0));
  nand2 gate688(.a(gate266inter0), .b(s_20), .O(gate266inter1));
  and2  gate689(.a(G773), .b(G645), .O(gate266inter2));
  inv1  gate690(.a(s_20), .O(gate266inter3));
  inv1  gate691(.a(s_21), .O(gate266inter4));
  nand2 gate692(.a(gate266inter4), .b(gate266inter3), .O(gate266inter5));
  nor2  gate693(.a(gate266inter5), .b(gate266inter2), .O(gate266inter6));
  inv1  gate694(.a(G645), .O(gate266inter7));
  inv1  gate695(.a(G773), .O(gate266inter8));
  nand2 gate696(.a(gate266inter8), .b(gate266inter7), .O(gate266inter9));
  nand2 gate697(.a(s_21), .b(gate266inter3), .O(gate266inter10));
  nor2  gate698(.a(gate266inter10), .b(gate266inter9), .O(gate266inter11));
  nor2  gate699(.a(gate266inter11), .b(gate266inter6), .O(gate266inter12));
  nand2 gate700(.a(gate266inter12), .b(gate266inter1), .O(G797));
nand2 gate267( .a(G648), .b(G776), .O(G800) );

  xor2  gate2913(.a(G779), .b(G651), .O(gate268inter0));
  nand2 gate2914(.a(gate268inter0), .b(s_338), .O(gate268inter1));
  and2  gate2915(.a(G779), .b(G651), .O(gate268inter2));
  inv1  gate2916(.a(s_338), .O(gate268inter3));
  inv1  gate2917(.a(s_339), .O(gate268inter4));
  nand2 gate2918(.a(gate268inter4), .b(gate268inter3), .O(gate268inter5));
  nor2  gate2919(.a(gate268inter5), .b(gate268inter2), .O(gate268inter6));
  inv1  gate2920(.a(G651), .O(gate268inter7));
  inv1  gate2921(.a(G779), .O(gate268inter8));
  nand2 gate2922(.a(gate268inter8), .b(gate268inter7), .O(gate268inter9));
  nand2 gate2923(.a(s_339), .b(gate268inter3), .O(gate268inter10));
  nor2  gate2924(.a(gate268inter10), .b(gate268inter9), .O(gate268inter11));
  nor2  gate2925(.a(gate268inter11), .b(gate268inter6), .O(gate268inter12));
  nand2 gate2926(.a(gate268inter12), .b(gate268inter1), .O(G803));
nand2 gate269( .a(G654), .b(G782), .O(G806) );

  xor2  gate1765(.a(G785), .b(G657), .O(gate270inter0));
  nand2 gate1766(.a(gate270inter0), .b(s_174), .O(gate270inter1));
  and2  gate1767(.a(G785), .b(G657), .O(gate270inter2));
  inv1  gate1768(.a(s_174), .O(gate270inter3));
  inv1  gate1769(.a(s_175), .O(gate270inter4));
  nand2 gate1770(.a(gate270inter4), .b(gate270inter3), .O(gate270inter5));
  nor2  gate1771(.a(gate270inter5), .b(gate270inter2), .O(gate270inter6));
  inv1  gate1772(.a(G657), .O(gate270inter7));
  inv1  gate1773(.a(G785), .O(gate270inter8));
  nand2 gate1774(.a(gate270inter8), .b(gate270inter7), .O(gate270inter9));
  nand2 gate1775(.a(s_175), .b(gate270inter3), .O(gate270inter10));
  nor2  gate1776(.a(gate270inter10), .b(gate270inter9), .O(gate270inter11));
  nor2  gate1777(.a(gate270inter11), .b(gate270inter6), .O(gate270inter12));
  nand2 gate1778(.a(gate270inter12), .b(gate270inter1), .O(G809));

  xor2  gate2717(.a(G788), .b(G660), .O(gate271inter0));
  nand2 gate2718(.a(gate271inter0), .b(s_310), .O(gate271inter1));
  and2  gate2719(.a(G788), .b(G660), .O(gate271inter2));
  inv1  gate2720(.a(s_310), .O(gate271inter3));
  inv1  gate2721(.a(s_311), .O(gate271inter4));
  nand2 gate2722(.a(gate271inter4), .b(gate271inter3), .O(gate271inter5));
  nor2  gate2723(.a(gate271inter5), .b(gate271inter2), .O(gate271inter6));
  inv1  gate2724(.a(G660), .O(gate271inter7));
  inv1  gate2725(.a(G788), .O(gate271inter8));
  nand2 gate2726(.a(gate271inter8), .b(gate271inter7), .O(gate271inter9));
  nand2 gate2727(.a(s_311), .b(gate271inter3), .O(gate271inter10));
  nor2  gate2728(.a(gate271inter10), .b(gate271inter9), .O(gate271inter11));
  nor2  gate2729(.a(gate271inter11), .b(gate271inter6), .O(gate271inter12));
  nand2 gate2730(.a(gate271inter12), .b(gate271inter1), .O(G812));
nand2 gate272( .a(G663), .b(G791), .O(G815) );
nand2 gate273( .a(G642), .b(G794), .O(G818) );
nand2 gate274( .a(G770), .b(G794), .O(G819) );
nand2 gate275( .a(G645), .b(G797), .O(G820) );

  xor2  gate2885(.a(G797), .b(G773), .O(gate276inter0));
  nand2 gate2886(.a(gate276inter0), .b(s_334), .O(gate276inter1));
  and2  gate2887(.a(G797), .b(G773), .O(gate276inter2));
  inv1  gate2888(.a(s_334), .O(gate276inter3));
  inv1  gate2889(.a(s_335), .O(gate276inter4));
  nand2 gate2890(.a(gate276inter4), .b(gate276inter3), .O(gate276inter5));
  nor2  gate2891(.a(gate276inter5), .b(gate276inter2), .O(gate276inter6));
  inv1  gate2892(.a(G773), .O(gate276inter7));
  inv1  gate2893(.a(G797), .O(gate276inter8));
  nand2 gate2894(.a(gate276inter8), .b(gate276inter7), .O(gate276inter9));
  nand2 gate2895(.a(s_335), .b(gate276inter3), .O(gate276inter10));
  nor2  gate2896(.a(gate276inter10), .b(gate276inter9), .O(gate276inter11));
  nor2  gate2897(.a(gate276inter11), .b(gate276inter6), .O(gate276inter12));
  nand2 gate2898(.a(gate276inter12), .b(gate276inter1), .O(G821));
nand2 gate277( .a(G648), .b(G800), .O(G822) );
nand2 gate278( .a(G776), .b(G800), .O(G823) );

  xor2  gate1835(.a(G803), .b(G651), .O(gate279inter0));
  nand2 gate1836(.a(gate279inter0), .b(s_184), .O(gate279inter1));
  and2  gate1837(.a(G803), .b(G651), .O(gate279inter2));
  inv1  gate1838(.a(s_184), .O(gate279inter3));
  inv1  gate1839(.a(s_185), .O(gate279inter4));
  nand2 gate1840(.a(gate279inter4), .b(gate279inter3), .O(gate279inter5));
  nor2  gate1841(.a(gate279inter5), .b(gate279inter2), .O(gate279inter6));
  inv1  gate1842(.a(G651), .O(gate279inter7));
  inv1  gate1843(.a(G803), .O(gate279inter8));
  nand2 gate1844(.a(gate279inter8), .b(gate279inter7), .O(gate279inter9));
  nand2 gate1845(.a(s_185), .b(gate279inter3), .O(gate279inter10));
  nor2  gate1846(.a(gate279inter10), .b(gate279inter9), .O(gate279inter11));
  nor2  gate1847(.a(gate279inter11), .b(gate279inter6), .O(gate279inter12));
  nand2 gate1848(.a(gate279inter12), .b(gate279inter1), .O(G824));
nand2 gate280( .a(G779), .b(G803), .O(G825) );

  xor2  gate2437(.a(G806), .b(G654), .O(gate281inter0));
  nand2 gate2438(.a(gate281inter0), .b(s_270), .O(gate281inter1));
  and2  gate2439(.a(G806), .b(G654), .O(gate281inter2));
  inv1  gate2440(.a(s_270), .O(gate281inter3));
  inv1  gate2441(.a(s_271), .O(gate281inter4));
  nand2 gate2442(.a(gate281inter4), .b(gate281inter3), .O(gate281inter5));
  nor2  gate2443(.a(gate281inter5), .b(gate281inter2), .O(gate281inter6));
  inv1  gate2444(.a(G654), .O(gate281inter7));
  inv1  gate2445(.a(G806), .O(gate281inter8));
  nand2 gate2446(.a(gate281inter8), .b(gate281inter7), .O(gate281inter9));
  nand2 gate2447(.a(s_271), .b(gate281inter3), .O(gate281inter10));
  nor2  gate2448(.a(gate281inter10), .b(gate281inter9), .O(gate281inter11));
  nor2  gate2449(.a(gate281inter11), .b(gate281inter6), .O(gate281inter12));
  nand2 gate2450(.a(gate281inter12), .b(gate281inter1), .O(G826));

  xor2  gate715(.a(G806), .b(G782), .O(gate282inter0));
  nand2 gate716(.a(gate282inter0), .b(s_24), .O(gate282inter1));
  and2  gate717(.a(G806), .b(G782), .O(gate282inter2));
  inv1  gate718(.a(s_24), .O(gate282inter3));
  inv1  gate719(.a(s_25), .O(gate282inter4));
  nand2 gate720(.a(gate282inter4), .b(gate282inter3), .O(gate282inter5));
  nor2  gate721(.a(gate282inter5), .b(gate282inter2), .O(gate282inter6));
  inv1  gate722(.a(G782), .O(gate282inter7));
  inv1  gate723(.a(G806), .O(gate282inter8));
  nand2 gate724(.a(gate282inter8), .b(gate282inter7), .O(gate282inter9));
  nand2 gate725(.a(s_25), .b(gate282inter3), .O(gate282inter10));
  nor2  gate726(.a(gate282inter10), .b(gate282inter9), .O(gate282inter11));
  nor2  gate727(.a(gate282inter11), .b(gate282inter6), .O(gate282inter12));
  nand2 gate728(.a(gate282inter12), .b(gate282inter1), .O(G827));

  xor2  gate1149(.a(G809), .b(G657), .O(gate283inter0));
  nand2 gate1150(.a(gate283inter0), .b(s_86), .O(gate283inter1));
  and2  gate1151(.a(G809), .b(G657), .O(gate283inter2));
  inv1  gate1152(.a(s_86), .O(gate283inter3));
  inv1  gate1153(.a(s_87), .O(gate283inter4));
  nand2 gate1154(.a(gate283inter4), .b(gate283inter3), .O(gate283inter5));
  nor2  gate1155(.a(gate283inter5), .b(gate283inter2), .O(gate283inter6));
  inv1  gate1156(.a(G657), .O(gate283inter7));
  inv1  gate1157(.a(G809), .O(gate283inter8));
  nand2 gate1158(.a(gate283inter8), .b(gate283inter7), .O(gate283inter9));
  nand2 gate1159(.a(s_87), .b(gate283inter3), .O(gate283inter10));
  nor2  gate1160(.a(gate283inter10), .b(gate283inter9), .O(gate283inter11));
  nor2  gate1161(.a(gate283inter11), .b(gate283inter6), .O(gate283inter12));
  nand2 gate1162(.a(gate283inter12), .b(gate283inter1), .O(G828));
nand2 gate284( .a(G785), .b(G809), .O(G829) );

  xor2  gate799(.a(G812), .b(G660), .O(gate285inter0));
  nand2 gate800(.a(gate285inter0), .b(s_36), .O(gate285inter1));
  and2  gate801(.a(G812), .b(G660), .O(gate285inter2));
  inv1  gate802(.a(s_36), .O(gate285inter3));
  inv1  gate803(.a(s_37), .O(gate285inter4));
  nand2 gate804(.a(gate285inter4), .b(gate285inter3), .O(gate285inter5));
  nor2  gate805(.a(gate285inter5), .b(gate285inter2), .O(gate285inter6));
  inv1  gate806(.a(G660), .O(gate285inter7));
  inv1  gate807(.a(G812), .O(gate285inter8));
  nand2 gate808(.a(gate285inter8), .b(gate285inter7), .O(gate285inter9));
  nand2 gate809(.a(s_37), .b(gate285inter3), .O(gate285inter10));
  nor2  gate810(.a(gate285inter10), .b(gate285inter9), .O(gate285inter11));
  nor2  gate811(.a(gate285inter11), .b(gate285inter6), .O(gate285inter12));
  nand2 gate812(.a(gate285inter12), .b(gate285inter1), .O(G830));

  xor2  gate1807(.a(G812), .b(G788), .O(gate286inter0));
  nand2 gate1808(.a(gate286inter0), .b(s_180), .O(gate286inter1));
  and2  gate1809(.a(G812), .b(G788), .O(gate286inter2));
  inv1  gate1810(.a(s_180), .O(gate286inter3));
  inv1  gate1811(.a(s_181), .O(gate286inter4));
  nand2 gate1812(.a(gate286inter4), .b(gate286inter3), .O(gate286inter5));
  nor2  gate1813(.a(gate286inter5), .b(gate286inter2), .O(gate286inter6));
  inv1  gate1814(.a(G788), .O(gate286inter7));
  inv1  gate1815(.a(G812), .O(gate286inter8));
  nand2 gate1816(.a(gate286inter8), .b(gate286inter7), .O(gate286inter9));
  nand2 gate1817(.a(s_181), .b(gate286inter3), .O(gate286inter10));
  nor2  gate1818(.a(gate286inter10), .b(gate286inter9), .O(gate286inter11));
  nor2  gate1819(.a(gate286inter11), .b(gate286inter6), .O(gate286inter12));
  nand2 gate1820(.a(gate286inter12), .b(gate286inter1), .O(G831));
nand2 gate287( .a(G663), .b(G815), .O(G832) );

  xor2  gate1205(.a(G815), .b(G791), .O(gate288inter0));
  nand2 gate1206(.a(gate288inter0), .b(s_94), .O(gate288inter1));
  and2  gate1207(.a(G815), .b(G791), .O(gate288inter2));
  inv1  gate1208(.a(s_94), .O(gate288inter3));
  inv1  gate1209(.a(s_95), .O(gate288inter4));
  nand2 gate1210(.a(gate288inter4), .b(gate288inter3), .O(gate288inter5));
  nor2  gate1211(.a(gate288inter5), .b(gate288inter2), .O(gate288inter6));
  inv1  gate1212(.a(G791), .O(gate288inter7));
  inv1  gate1213(.a(G815), .O(gate288inter8));
  nand2 gate1214(.a(gate288inter8), .b(gate288inter7), .O(gate288inter9));
  nand2 gate1215(.a(s_95), .b(gate288inter3), .O(gate288inter10));
  nor2  gate1216(.a(gate288inter10), .b(gate288inter9), .O(gate288inter11));
  nor2  gate1217(.a(gate288inter11), .b(gate288inter6), .O(gate288inter12));
  nand2 gate1218(.a(gate288inter12), .b(gate288inter1), .O(G833));
nand2 gate289( .a(G818), .b(G819), .O(G834) );

  xor2  gate771(.a(G821), .b(G820), .O(gate290inter0));
  nand2 gate772(.a(gate290inter0), .b(s_32), .O(gate290inter1));
  and2  gate773(.a(G821), .b(G820), .O(gate290inter2));
  inv1  gate774(.a(s_32), .O(gate290inter3));
  inv1  gate775(.a(s_33), .O(gate290inter4));
  nand2 gate776(.a(gate290inter4), .b(gate290inter3), .O(gate290inter5));
  nor2  gate777(.a(gate290inter5), .b(gate290inter2), .O(gate290inter6));
  inv1  gate778(.a(G820), .O(gate290inter7));
  inv1  gate779(.a(G821), .O(gate290inter8));
  nand2 gate780(.a(gate290inter8), .b(gate290inter7), .O(gate290inter9));
  nand2 gate781(.a(s_33), .b(gate290inter3), .O(gate290inter10));
  nor2  gate782(.a(gate290inter10), .b(gate290inter9), .O(gate290inter11));
  nor2  gate783(.a(gate290inter11), .b(gate290inter6), .O(gate290inter12));
  nand2 gate784(.a(gate290inter12), .b(gate290inter1), .O(G847));

  xor2  gate2605(.a(G823), .b(G822), .O(gate291inter0));
  nand2 gate2606(.a(gate291inter0), .b(s_294), .O(gate291inter1));
  and2  gate2607(.a(G823), .b(G822), .O(gate291inter2));
  inv1  gate2608(.a(s_294), .O(gate291inter3));
  inv1  gate2609(.a(s_295), .O(gate291inter4));
  nand2 gate2610(.a(gate291inter4), .b(gate291inter3), .O(gate291inter5));
  nor2  gate2611(.a(gate291inter5), .b(gate291inter2), .O(gate291inter6));
  inv1  gate2612(.a(G822), .O(gate291inter7));
  inv1  gate2613(.a(G823), .O(gate291inter8));
  nand2 gate2614(.a(gate291inter8), .b(gate291inter7), .O(gate291inter9));
  nand2 gate2615(.a(s_295), .b(gate291inter3), .O(gate291inter10));
  nor2  gate2616(.a(gate291inter10), .b(gate291inter9), .O(gate291inter11));
  nor2  gate2617(.a(gate291inter11), .b(gate291inter6), .O(gate291inter12));
  nand2 gate2618(.a(gate291inter12), .b(gate291inter1), .O(G860));
nand2 gate292( .a(G824), .b(G825), .O(G873) );
nand2 gate293( .a(G828), .b(G829), .O(G886) );
nand2 gate294( .a(G832), .b(G833), .O(G899) );
nand2 gate295( .a(G830), .b(G831), .O(G912) );
nand2 gate296( .a(G826), .b(G827), .O(G925) );
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );

  xor2  gate2577(.a(G1036), .b(G1), .O(gate387inter0));
  nand2 gate2578(.a(gate387inter0), .b(s_290), .O(gate387inter1));
  and2  gate2579(.a(G1036), .b(G1), .O(gate387inter2));
  inv1  gate2580(.a(s_290), .O(gate387inter3));
  inv1  gate2581(.a(s_291), .O(gate387inter4));
  nand2 gate2582(.a(gate387inter4), .b(gate387inter3), .O(gate387inter5));
  nor2  gate2583(.a(gate387inter5), .b(gate387inter2), .O(gate387inter6));
  inv1  gate2584(.a(G1), .O(gate387inter7));
  inv1  gate2585(.a(G1036), .O(gate387inter8));
  nand2 gate2586(.a(gate387inter8), .b(gate387inter7), .O(gate387inter9));
  nand2 gate2587(.a(s_291), .b(gate387inter3), .O(gate387inter10));
  nor2  gate2588(.a(gate387inter10), .b(gate387inter9), .O(gate387inter11));
  nor2  gate2589(.a(gate387inter11), .b(gate387inter6), .O(gate387inter12));
  nand2 gate2590(.a(gate387inter12), .b(gate387inter1), .O(G1132));
nand2 gate388( .a(G2), .b(G1039), .O(G1135) );
nand2 gate389( .a(G3), .b(G1042), .O(G1138) );
nand2 gate390( .a(G4), .b(G1045), .O(G1141) );

  xor2  gate897(.a(G1048), .b(G5), .O(gate391inter0));
  nand2 gate898(.a(gate391inter0), .b(s_50), .O(gate391inter1));
  and2  gate899(.a(G1048), .b(G5), .O(gate391inter2));
  inv1  gate900(.a(s_50), .O(gate391inter3));
  inv1  gate901(.a(s_51), .O(gate391inter4));
  nand2 gate902(.a(gate391inter4), .b(gate391inter3), .O(gate391inter5));
  nor2  gate903(.a(gate391inter5), .b(gate391inter2), .O(gate391inter6));
  inv1  gate904(.a(G5), .O(gate391inter7));
  inv1  gate905(.a(G1048), .O(gate391inter8));
  nand2 gate906(.a(gate391inter8), .b(gate391inter7), .O(gate391inter9));
  nand2 gate907(.a(s_51), .b(gate391inter3), .O(gate391inter10));
  nor2  gate908(.a(gate391inter10), .b(gate391inter9), .O(gate391inter11));
  nor2  gate909(.a(gate391inter11), .b(gate391inter6), .O(gate391inter12));
  nand2 gate910(.a(gate391inter12), .b(gate391inter1), .O(G1144));
nand2 gate392( .a(G6), .b(G1051), .O(G1147) );
nand2 gate393( .a(G7), .b(G1054), .O(G1150) );

  xor2  gate2815(.a(G1057), .b(G8), .O(gate394inter0));
  nand2 gate2816(.a(gate394inter0), .b(s_324), .O(gate394inter1));
  and2  gate2817(.a(G1057), .b(G8), .O(gate394inter2));
  inv1  gate2818(.a(s_324), .O(gate394inter3));
  inv1  gate2819(.a(s_325), .O(gate394inter4));
  nand2 gate2820(.a(gate394inter4), .b(gate394inter3), .O(gate394inter5));
  nor2  gate2821(.a(gate394inter5), .b(gate394inter2), .O(gate394inter6));
  inv1  gate2822(.a(G8), .O(gate394inter7));
  inv1  gate2823(.a(G1057), .O(gate394inter8));
  nand2 gate2824(.a(gate394inter8), .b(gate394inter7), .O(gate394inter9));
  nand2 gate2825(.a(s_325), .b(gate394inter3), .O(gate394inter10));
  nor2  gate2826(.a(gate394inter10), .b(gate394inter9), .O(gate394inter11));
  nor2  gate2827(.a(gate394inter11), .b(gate394inter6), .O(gate394inter12));
  nand2 gate2828(.a(gate394inter12), .b(gate394inter1), .O(G1153));
nand2 gate395( .a(G9), .b(G1060), .O(G1156) );
nand2 gate396( .a(G10), .b(G1063), .O(G1159) );
nand2 gate397( .a(G11), .b(G1066), .O(G1162) );
nand2 gate398( .a(G12), .b(G1069), .O(G1165) );

  xor2  gate2507(.a(G1072), .b(G13), .O(gate399inter0));
  nand2 gate2508(.a(gate399inter0), .b(s_280), .O(gate399inter1));
  and2  gate2509(.a(G1072), .b(G13), .O(gate399inter2));
  inv1  gate2510(.a(s_280), .O(gate399inter3));
  inv1  gate2511(.a(s_281), .O(gate399inter4));
  nand2 gate2512(.a(gate399inter4), .b(gate399inter3), .O(gate399inter5));
  nor2  gate2513(.a(gate399inter5), .b(gate399inter2), .O(gate399inter6));
  inv1  gate2514(.a(G13), .O(gate399inter7));
  inv1  gate2515(.a(G1072), .O(gate399inter8));
  nand2 gate2516(.a(gate399inter8), .b(gate399inter7), .O(gate399inter9));
  nand2 gate2517(.a(s_281), .b(gate399inter3), .O(gate399inter10));
  nor2  gate2518(.a(gate399inter10), .b(gate399inter9), .O(gate399inter11));
  nor2  gate2519(.a(gate399inter11), .b(gate399inter6), .O(gate399inter12));
  nand2 gate2520(.a(gate399inter12), .b(gate399inter1), .O(G1168));

  xor2  gate1653(.a(G1075), .b(G14), .O(gate400inter0));
  nand2 gate1654(.a(gate400inter0), .b(s_158), .O(gate400inter1));
  and2  gate1655(.a(G1075), .b(G14), .O(gate400inter2));
  inv1  gate1656(.a(s_158), .O(gate400inter3));
  inv1  gate1657(.a(s_159), .O(gate400inter4));
  nand2 gate1658(.a(gate400inter4), .b(gate400inter3), .O(gate400inter5));
  nor2  gate1659(.a(gate400inter5), .b(gate400inter2), .O(gate400inter6));
  inv1  gate1660(.a(G14), .O(gate400inter7));
  inv1  gate1661(.a(G1075), .O(gate400inter8));
  nand2 gate1662(.a(gate400inter8), .b(gate400inter7), .O(gate400inter9));
  nand2 gate1663(.a(s_159), .b(gate400inter3), .O(gate400inter10));
  nor2  gate1664(.a(gate400inter10), .b(gate400inter9), .O(gate400inter11));
  nor2  gate1665(.a(gate400inter11), .b(gate400inter6), .O(gate400inter12));
  nand2 gate1666(.a(gate400inter12), .b(gate400inter1), .O(G1171));
nand2 gate401( .a(G15), .b(G1078), .O(G1174) );

  xor2  gate1485(.a(G1081), .b(G16), .O(gate402inter0));
  nand2 gate1486(.a(gate402inter0), .b(s_134), .O(gate402inter1));
  and2  gate1487(.a(G1081), .b(G16), .O(gate402inter2));
  inv1  gate1488(.a(s_134), .O(gate402inter3));
  inv1  gate1489(.a(s_135), .O(gate402inter4));
  nand2 gate1490(.a(gate402inter4), .b(gate402inter3), .O(gate402inter5));
  nor2  gate1491(.a(gate402inter5), .b(gate402inter2), .O(gate402inter6));
  inv1  gate1492(.a(G16), .O(gate402inter7));
  inv1  gate1493(.a(G1081), .O(gate402inter8));
  nand2 gate1494(.a(gate402inter8), .b(gate402inter7), .O(gate402inter9));
  nand2 gate1495(.a(s_135), .b(gate402inter3), .O(gate402inter10));
  nor2  gate1496(.a(gate402inter10), .b(gate402inter9), .O(gate402inter11));
  nor2  gate1497(.a(gate402inter11), .b(gate402inter6), .O(gate402inter12));
  nand2 gate1498(.a(gate402inter12), .b(gate402inter1), .O(G1177));

  xor2  gate2843(.a(G1084), .b(G17), .O(gate403inter0));
  nand2 gate2844(.a(gate403inter0), .b(s_328), .O(gate403inter1));
  and2  gate2845(.a(G1084), .b(G17), .O(gate403inter2));
  inv1  gate2846(.a(s_328), .O(gate403inter3));
  inv1  gate2847(.a(s_329), .O(gate403inter4));
  nand2 gate2848(.a(gate403inter4), .b(gate403inter3), .O(gate403inter5));
  nor2  gate2849(.a(gate403inter5), .b(gate403inter2), .O(gate403inter6));
  inv1  gate2850(.a(G17), .O(gate403inter7));
  inv1  gate2851(.a(G1084), .O(gate403inter8));
  nand2 gate2852(.a(gate403inter8), .b(gate403inter7), .O(gate403inter9));
  nand2 gate2853(.a(s_329), .b(gate403inter3), .O(gate403inter10));
  nor2  gate2854(.a(gate403inter10), .b(gate403inter9), .O(gate403inter11));
  nor2  gate2855(.a(gate403inter11), .b(gate403inter6), .O(gate403inter12));
  nand2 gate2856(.a(gate403inter12), .b(gate403inter1), .O(G1180));
nand2 gate404( .a(G18), .b(G1087), .O(G1183) );
nand2 gate405( .a(G19), .b(G1090), .O(G1186) );

  xor2  gate1681(.a(G1093), .b(G20), .O(gate406inter0));
  nand2 gate1682(.a(gate406inter0), .b(s_162), .O(gate406inter1));
  and2  gate1683(.a(G1093), .b(G20), .O(gate406inter2));
  inv1  gate1684(.a(s_162), .O(gate406inter3));
  inv1  gate1685(.a(s_163), .O(gate406inter4));
  nand2 gate1686(.a(gate406inter4), .b(gate406inter3), .O(gate406inter5));
  nor2  gate1687(.a(gate406inter5), .b(gate406inter2), .O(gate406inter6));
  inv1  gate1688(.a(G20), .O(gate406inter7));
  inv1  gate1689(.a(G1093), .O(gate406inter8));
  nand2 gate1690(.a(gate406inter8), .b(gate406inter7), .O(gate406inter9));
  nand2 gate1691(.a(s_163), .b(gate406inter3), .O(gate406inter10));
  nor2  gate1692(.a(gate406inter10), .b(gate406inter9), .O(gate406inter11));
  nor2  gate1693(.a(gate406inter11), .b(gate406inter6), .O(gate406inter12));
  nand2 gate1694(.a(gate406inter12), .b(gate406inter1), .O(G1189));
nand2 gate407( .a(G21), .b(G1096), .O(G1192) );

  xor2  gate1499(.a(G1099), .b(G22), .O(gate408inter0));
  nand2 gate1500(.a(gate408inter0), .b(s_136), .O(gate408inter1));
  and2  gate1501(.a(G1099), .b(G22), .O(gate408inter2));
  inv1  gate1502(.a(s_136), .O(gate408inter3));
  inv1  gate1503(.a(s_137), .O(gate408inter4));
  nand2 gate1504(.a(gate408inter4), .b(gate408inter3), .O(gate408inter5));
  nor2  gate1505(.a(gate408inter5), .b(gate408inter2), .O(gate408inter6));
  inv1  gate1506(.a(G22), .O(gate408inter7));
  inv1  gate1507(.a(G1099), .O(gate408inter8));
  nand2 gate1508(.a(gate408inter8), .b(gate408inter7), .O(gate408inter9));
  nand2 gate1509(.a(s_137), .b(gate408inter3), .O(gate408inter10));
  nor2  gate1510(.a(gate408inter10), .b(gate408inter9), .O(gate408inter11));
  nor2  gate1511(.a(gate408inter11), .b(gate408inter6), .O(gate408inter12));
  nand2 gate1512(.a(gate408inter12), .b(gate408inter1), .O(G1195));
nand2 gate409( .a(G23), .b(G1102), .O(G1198) );

  xor2  gate2549(.a(G1105), .b(G24), .O(gate410inter0));
  nand2 gate2550(.a(gate410inter0), .b(s_286), .O(gate410inter1));
  and2  gate2551(.a(G1105), .b(G24), .O(gate410inter2));
  inv1  gate2552(.a(s_286), .O(gate410inter3));
  inv1  gate2553(.a(s_287), .O(gate410inter4));
  nand2 gate2554(.a(gate410inter4), .b(gate410inter3), .O(gate410inter5));
  nor2  gate2555(.a(gate410inter5), .b(gate410inter2), .O(gate410inter6));
  inv1  gate2556(.a(G24), .O(gate410inter7));
  inv1  gate2557(.a(G1105), .O(gate410inter8));
  nand2 gate2558(.a(gate410inter8), .b(gate410inter7), .O(gate410inter9));
  nand2 gate2559(.a(s_287), .b(gate410inter3), .O(gate410inter10));
  nor2  gate2560(.a(gate410inter10), .b(gate410inter9), .O(gate410inter11));
  nor2  gate2561(.a(gate410inter11), .b(gate410inter6), .O(gate410inter12));
  nand2 gate2562(.a(gate410inter12), .b(gate410inter1), .O(G1201));
nand2 gate411( .a(G25), .b(G1108), .O(G1204) );

  xor2  gate1541(.a(G1111), .b(G26), .O(gate412inter0));
  nand2 gate1542(.a(gate412inter0), .b(s_142), .O(gate412inter1));
  and2  gate1543(.a(G1111), .b(G26), .O(gate412inter2));
  inv1  gate1544(.a(s_142), .O(gate412inter3));
  inv1  gate1545(.a(s_143), .O(gate412inter4));
  nand2 gate1546(.a(gate412inter4), .b(gate412inter3), .O(gate412inter5));
  nor2  gate1547(.a(gate412inter5), .b(gate412inter2), .O(gate412inter6));
  inv1  gate1548(.a(G26), .O(gate412inter7));
  inv1  gate1549(.a(G1111), .O(gate412inter8));
  nand2 gate1550(.a(gate412inter8), .b(gate412inter7), .O(gate412inter9));
  nand2 gate1551(.a(s_143), .b(gate412inter3), .O(gate412inter10));
  nor2  gate1552(.a(gate412inter10), .b(gate412inter9), .O(gate412inter11));
  nor2  gate1553(.a(gate412inter11), .b(gate412inter6), .O(gate412inter12));
  nand2 gate1554(.a(gate412inter12), .b(gate412inter1), .O(G1207));
nand2 gate413( .a(G27), .b(G1114), .O(G1210) );
nand2 gate414( .a(G28), .b(G1117), .O(G1213) );

  xor2  gate2745(.a(G1120), .b(G29), .O(gate415inter0));
  nand2 gate2746(.a(gate415inter0), .b(s_314), .O(gate415inter1));
  and2  gate2747(.a(G1120), .b(G29), .O(gate415inter2));
  inv1  gate2748(.a(s_314), .O(gate415inter3));
  inv1  gate2749(.a(s_315), .O(gate415inter4));
  nand2 gate2750(.a(gate415inter4), .b(gate415inter3), .O(gate415inter5));
  nor2  gate2751(.a(gate415inter5), .b(gate415inter2), .O(gate415inter6));
  inv1  gate2752(.a(G29), .O(gate415inter7));
  inv1  gate2753(.a(G1120), .O(gate415inter8));
  nand2 gate2754(.a(gate415inter8), .b(gate415inter7), .O(gate415inter9));
  nand2 gate2755(.a(s_315), .b(gate415inter3), .O(gate415inter10));
  nor2  gate2756(.a(gate415inter10), .b(gate415inter9), .O(gate415inter11));
  nor2  gate2757(.a(gate415inter11), .b(gate415inter6), .O(gate415inter12));
  nand2 gate2758(.a(gate415inter12), .b(gate415inter1), .O(G1216));
nand2 gate416( .a(G30), .b(G1123), .O(G1219) );

  xor2  gate1625(.a(G1126), .b(G31), .O(gate417inter0));
  nand2 gate1626(.a(gate417inter0), .b(s_154), .O(gate417inter1));
  and2  gate1627(.a(G1126), .b(G31), .O(gate417inter2));
  inv1  gate1628(.a(s_154), .O(gate417inter3));
  inv1  gate1629(.a(s_155), .O(gate417inter4));
  nand2 gate1630(.a(gate417inter4), .b(gate417inter3), .O(gate417inter5));
  nor2  gate1631(.a(gate417inter5), .b(gate417inter2), .O(gate417inter6));
  inv1  gate1632(.a(G31), .O(gate417inter7));
  inv1  gate1633(.a(G1126), .O(gate417inter8));
  nand2 gate1634(.a(gate417inter8), .b(gate417inter7), .O(gate417inter9));
  nand2 gate1635(.a(s_155), .b(gate417inter3), .O(gate417inter10));
  nor2  gate1636(.a(gate417inter10), .b(gate417inter9), .O(gate417inter11));
  nor2  gate1637(.a(gate417inter11), .b(gate417inter6), .O(gate417inter12));
  nand2 gate1638(.a(gate417inter12), .b(gate417inter1), .O(G1222));

  xor2  gate1247(.a(G1129), .b(G32), .O(gate418inter0));
  nand2 gate1248(.a(gate418inter0), .b(s_100), .O(gate418inter1));
  and2  gate1249(.a(G1129), .b(G32), .O(gate418inter2));
  inv1  gate1250(.a(s_100), .O(gate418inter3));
  inv1  gate1251(.a(s_101), .O(gate418inter4));
  nand2 gate1252(.a(gate418inter4), .b(gate418inter3), .O(gate418inter5));
  nor2  gate1253(.a(gate418inter5), .b(gate418inter2), .O(gate418inter6));
  inv1  gate1254(.a(G32), .O(gate418inter7));
  inv1  gate1255(.a(G1129), .O(gate418inter8));
  nand2 gate1256(.a(gate418inter8), .b(gate418inter7), .O(gate418inter9));
  nand2 gate1257(.a(s_101), .b(gate418inter3), .O(gate418inter10));
  nor2  gate1258(.a(gate418inter10), .b(gate418inter9), .O(gate418inter11));
  nor2  gate1259(.a(gate418inter11), .b(gate418inter6), .O(gate418inter12));
  nand2 gate1260(.a(gate418inter12), .b(gate418inter1), .O(G1225));
nand2 gate419( .a(G1), .b(G1132), .O(G1228) );
nand2 gate420( .a(G1036), .b(G1132), .O(G1229) );

  xor2  gate1177(.a(G1135), .b(G2), .O(gate421inter0));
  nand2 gate1178(.a(gate421inter0), .b(s_90), .O(gate421inter1));
  and2  gate1179(.a(G1135), .b(G2), .O(gate421inter2));
  inv1  gate1180(.a(s_90), .O(gate421inter3));
  inv1  gate1181(.a(s_91), .O(gate421inter4));
  nand2 gate1182(.a(gate421inter4), .b(gate421inter3), .O(gate421inter5));
  nor2  gate1183(.a(gate421inter5), .b(gate421inter2), .O(gate421inter6));
  inv1  gate1184(.a(G2), .O(gate421inter7));
  inv1  gate1185(.a(G1135), .O(gate421inter8));
  nand2 gate1186(.a(gate421inter8), .b(gate421inter7), .O(gate421inter9));
  nand2 gate1187(.a(s_91), .b(gate421inter3), .O(gate421inter10));
  nor2  gate1188(.a(gate421inter10), .b(gate421inter9), .O(gate421inter11));
  nor2  gate1189(.a(gate421inter11), .b(gate421inter6), .O(gate421inter12));
  nand2 gate1190(.a(gate421inter12), .b(gate421inter1), .O(G1230));
nand2 gate422( .a(G1039), .b(G1135), .O(G1231) );
nand2 gate423( .a(G3), .b(G1138), .O(G1232) );
nand2 gate424( .a(G1042), .b(G1138), .O(G1233) );
nand2 gate425( .a(G4), .b(G1141), .O(G1234) );
nand2 gate426( .a(G1045), .b(G1141), .O(G1235) );
nand2 gate427( .a(G5), .b(G1144), .O(G1236) );
nand2 gate428( .a(G1048), .b(G1144), .O(G1237) );

  xor2  gate953(.a(G1147), .b(G6), .O(gate429inter0));
  nand2 gate954(.a(gate429inter0), .b(s_58), .O(gate429inter1));
  and2  gate955(.a(G1147), .b(G6), .O(gate429inter2));
  inv1  gate956(.a(s_58), .O(gate429inter3));
  inv1  gate957(.a(s_59), .O(gate429inter4));
  nand2 gate958(.a(gate429inter4), .b(gate429inter3), .O(gate429inter5));
  nor2  gate959(.a(gate429inter5), .b(gate429inter2), .O(gate429inter6));
  inv1  gate960(.a(G6), .O(gate429inter7));
  inv1  gate961(.a(G1147), .O(gate429inter8));
  nand2 gate962(.a(gate429inter8), .b(gate429inter7), .O(gate429inter9));
  nand2 gate963(.a(s_59), .b(gate429inter3), .O(gate429inter10));
  nor2  gate964(.a(gate429inter10), .b(gate429inter9), .O(gate429inter11));
  nor2  gate965(.a(gate429inter11), .b(gate429inter6), .O(gate429inter12));
  nand2 gate966(.a(gate429inter12), .b(gate429inter1), .O(G1238));

  xor2  gate1583(.a(G1147), .b(G1051), .O(gate430inter0));
  nand2 gate1584(.a(gate430inter0), .b(s_148), .O(gate430inter1));
  and2  gate1585(.a(G1147), .b(G1051), .O(gate430inter2));
  inv1  gate1586(.a(s_148), .O(gate430inter3));
  inv1  gate1587(.a(s_149), .O(gate430inter4));
  nand2 gate1588(.a(gate430inter4), .b(gate430inter3), .O(gate430inter5));
  nor2  gate1589(.a(gate430inter5), .b(gate430inter2), .O(gate430inter6));
  inv1  gate1590(.a(G1051), .O(gate430inter7));
  inv1  gate1591(.a(G1147), .O(gate430inter8));
  nand2 gate1592(.a(gate430inter8), .b(gate430inter7), .O(gate430inter9));
  nand2 gate1593(.a(s_149), .b(gate430inter3), .O(gate430inter10));
  nor2  gate1594(.a(gate430inter10), .b(gate430inter9), .O(gate430inter11));
  nor2  gate1595(.a(gate430inter11), .b(gate430inter6), .O(gate430inter12));
  nand2 gate1596(.a(gate430inter12), .b(gate430inter1), .O(G1239));

  xor2  gate911(.a(G1150), .b(G7), .O(gate431inter0));
  nand2 gate912(.a(gate431inter0), .b(s_52), .O(gate431inter1));
  and2  gate913(.a(G1150), .b(G7), .O(gate431inter2));
  inv1  gate914(.a(s_52), .O(gate431inter3));
  inv1  gate915(.a(s_53), .O(gate431inter4));
  nand2 gate916(.a(gate431inter4), .b(gate431inter3), .O(gate431inter5));
  nor2  gate917(.a(gate431inter5), .b(gate431inter2), .O(gate431inter6));
  inv1  gate918(.a(G7), .O(gate431inter7));
  inv1  gate919(.a(G1150), .O(gate431inter8));
  nand2 gate920(.a(gate431inter8), .b(gate431inter7), .O(gate431inter9));
  nand2 gate921(.a(s_53), .b(gate431inter3), .O(gate431inter10));
  nor2  gate922(.a(gate431inter10), .b(gate431inter9), .O(gate431inter11));
  nor2  gate923(.a(gate431inter11), .b(gate431inter6), .O(gate431inter12));
  nand2 gate924(.a(gate431inter12), .b(gate431inter1), .O(G1240));
nand2 gate432( .a(G1054), .b(G1150), .O(G1241) );
nand2 gate433( .a(G8), .b(G1153), .O(G1242) );

  xor2  gate2871(.a(G1153), .b(G1057), .O(gate434inter0));
  nand2 gate2872(.a(gate434inter0), .b(s_332), .O(gate434inter1));
  and2  gate2873(.a(G1153), .b(G1057), .O(gate434inter2));
  inv1  gate2874(.a(s_332), .O(gate434inter3));
  inv1  gate2875(.a(s_333), .O(gate434inter4));
  nand2 gate2876(.a(gate434inter4), .b(gate434inter3), .O(gate434inter5));
  nor2  gate2877(.a(gate434inter5), .b(gate434inter2), .O(gate434inter6));
  inv1  gate2878(.a(G1057), .O(gate434inter7));
  inv1  gate2879(.a(G1153), .O(gate434inter8));
  nand2 gate2880(.a(gate434inter8), .b(gate434inter7), .O(gate434inter9));
  nand2 gate2881(.a(s_333), .b(gate434inter3), .O(gate434inter10));
  nor2  gate2882(.a(gate434inter10), .b(gate434inter9), .O(gate434inter11));
  nor2  gate2883(.a(gate434inter11), .b(gate434inter6), .O(gate434inter12));
  nand2 gate2884(.a(gate434inter12), .b(gate434inter1), .O(G1243));

  xor2  gate2199(.a(G1156), .b(G9), .O(gate435inter0));
  nand2 gate2200(.a(gate435inter0), .b(s_236), .O(gate435inter1));
  and2  gate2201(.a(G1156), .b(G9), .O(gate435inter2));
  inv1  gate2202(.a(s_236), .O(gate435inter3));
  inv1  gate2203(.a(s_237), .O(gate435inter4));
  nand2 gate2204(.a(gate435inter4), .b(gate435inter3), .O(gate435inter5));
  nor2  gate2205(.a(gate435inter5), .b(gate435inter2), .O(gate435inter6));
  inv1  gate2206(.a(G9), .O(gate435inter7));
  inv1  gate2207(.a(G1156), .O(gate435inter8));
  nand2 gate2208(.a(gate435inter8), .b(gate435inter7), .O(gate435inter9));
  nand2 gate2209(.a(s_237), .b(gate435inter3), .O(gate435inter10));
  nor2  gate2210(.a(gate435inter10), .b(gate435inter9), .O(gate435inter11));
  nor2  gate2211(.a(gate435inter11), .b(gate435inter6), .O(gate435inter12));
  nand2 gate2212(.a(gate435inter12), .b(gate435inter1), .O(G1244));

  xor2  gate2353(.a(G1156), .b(G1060), .O(gate436inter0));
  nand2 gate2354(.a(gate436inter0), .b(s_258), .O(gate436inter1));
  and2  gate2355(.a(G1156), .b(G1060), .O(gate436inter2));
  inv1  gate2356(.a(s_258), .O(gate436inter3));
  inv1  gate2357(.a(s_259), .O(gate436inter4));
  nand2 gate2358(.a(gate436inter4), .b(gate436inter3), .O(gate436inter5));
  nor2  gate2359(.a(gate436inter5), .b(gate436inter2), .O(gate436inter6));
  inv1  gate2360(.a(G1060), .O(gate436inter7));
  inv1  gate2361(.a(G1156), .O(gate436inter8));
  nand2 gate2362(.a(gate436inter8), .b(gate436inter7), .O(gate436inter9));
  nand2 gate2363(.a(s_259), .b(gate436inter3), .O(gate436inter10));
  nor2  gate2364(.a(gate436inter10), .b(gate436inter9), .O(gate436inter11));
  nor2  gate2365(.a(gate436inter11), .b(gate436inter6), .O(gate436inter12));
  nand2 gate2366(.a(gate436inter12), .b(gate436inter1), .O(G1245));
nand2 gate437( .a(G10), .b(G1159), .O(G1246) );

  xor2  gate2633(.a(G1159), .b(G1063), .O(gate438inter0));
  nand2 gate2634(.a(gate438inter0), .b(s_298), .O(gate438inter1));
  and2  gate2635(.a(G1159), .b(G1063), .O(gate438inter2));
  inv1  gate2636(.a(s_298), .O(gate438inter3));
  inv1  gate2637(.a(s_299), .O(gate438inter4));
  nand2 gate2638(.a(gate438inter4), .b(gate438inter3), .O(gate438inter5));
  nor2  gate2639(.a(gate438inter5), .b(gate438inter2), .O(gate438inter6));
  inv1  gate2640(.a(G1063), .O(gate438inter7));
  inv1  gate2641(.a(G1159), .O(gate438inter8));
  nand2 gate2642(.a(gate438inter8), .b(gate438inter7), .O(gate438inter9));
  nand2 gate2643(.a(s_299), .b(gate438inter3), .O(gate438inter10));
  nor2  gate2644(.a(gate438inter10), .b(gate438inter9), .O(gate438inter11));
  nor2  gate2645(.a(gate438inter11), .b(gate438inter6), .O(gate438inter12));
  nand2 gate2646(.a(gate438inter12), .b(gate438inter1), .O(G1247));
nand2 gate439( .a(G11), .b(G1162), .O(G1248) );
nand2 gate440( .a(G1066), .b(G1162), .O(G1249) );

  xor2  gate1275(.a(G1165), .b(G12), .O(gate441inter0));
  nand2 gate1276(.a(gate441inter0), .b(s_104), .O(gate441inter1));
  and2  gate1277(.a(G1165), .b(G12), .O(gate441inter2));
  inv1  gate1278(.a(s_104), .O(gate441inter3));
  inv1  gate1279(.a(s_105), .O(gate441inter4));
  nand2 gate1280(.a(gate441inter4), .b(gate441inter3), .O(gate441inter5));
  nor2  gate1281(.a(gate441inter5), .b(gate441inter2), .O(gate441inter6));
  inv1  gate1282(.a(G12), .O(gate441inter7));
  inv1  gate1283(.a(G1165), .O(gate441inter8));
  nand2 gate1284(.a(gate441inter8), .b(gate441inter7), .O(gate441inter9));
  nand2 gate1285(.a(s_105), .b(gate441inter3), .O(gate441inter10));
  nor2  gate1286(.a(gate441inter10), .b(gate441inter9), .O(gate441inter11));
  nor2  gate1287(.a(gate441inter11), .b(gate441inter6), .O(gate441inter12));
  nand2 gate1288(.a(gate441inter12), .b(gate441inter1), .O(G1250));

  xor2  gate2675(.a(G1165), .b(G1069), .O(gate442inter0));
  nand2 gate2676(.a(gate442inter0), .b(s_304), .O(gate442inter1));
  and2  gate2677(.a(G1165), .b(G1069), .O(gate442inter2));
  inv1  gate2678(.a(s_304), .O(gate442inter3));
  inv1  gate2679(.a(s_305), .O(gate442inter4));
  nand2 gate2680(.a(gate442inter4), .b(gate442inter3), .O(gate442inter5));
  nor2  gate2681(.a(gate442inter5), .b(gate442inter2), .O(gate442inter6));
  inv1  gate2682(.a(G1069), .O(gate442inter7));
  inv1  gate2683(.a(G1165), .O(gate442inter8));
  nand2 gate2684(.a(gate442inter8), .b(gate442inter7), .O(gate442inter9));
  nand2 gate2685(.a(s_305), .b(gate442inter3), .O(gate442inter10));
  nor2  gate2686(.a(gate442inter10), .b(gate442inter9), .O(gate442inter11));
  nor2  gate2687(.a(gate442inter11), .b(gate442inter6), .O(gate442inter12));
  nand2 gate2688(.a(gate442inter12), .b(gate442inter1), .O(G1251));

  xor2  gate2045(.a(G1168), .b(G13), .O(gate443inter0));
  nand2 gate2046(.a(gate443inter0), .b(s_214), .O(gate443inter1));
  and2  gate2047(.a(G1168), .b(G13), .O(gate443inter2));
  inv1  gate2048(.a(s_214), .O(gate443inter3));
  inv1  gate2049(.a(s_215), .O(gate443inter4));
  nand2 gate2050(.a(gate443inter4), .b(gate443inter3), .O(gate443inter5));
  nor2  gate2051(.a(gate443inter5), .b(gate443inter2), .O(gate443inter6));
  inv1  gate2052(.a(G13), .O(gate443inter7));
  inv1  gate2053(.a(G1168), .O(gate443inter8));
  nand2 gate2054(.a(gate443inter8), .b(gate443inter7), .O(gate443inter9));
  nand2 gate2055(.a(s_215), .b(gate443inter3), .O(gate443inter10));
  nor2  gate2056(.a(gate443inter10), .b(gate443inter9), .O(gate443inter11));
  nor2  gate2057(.a(gate443inter11), .b(gate443inter6), .O(gate443inter12));
  nand2 gate2058(.a(gate443inter12), .b(gate443inter1), .O(G1252));
nand2 gate444( .a(G1072), .b(G1168), .O(G1253) );

  xor2  gate1555(.a(G1171), .b(G14), .O(gate445inter0));
  nand2 gate1556(.a(gate445inter0), .b(s_144), .O(gate445inter1));
  and2  gate1557(.a(G1171), .b(G14), .O(gate445inter2));
  inv1  gate1558(.a(s_144), .O(gate445inter3));
  inv1  gate1559(.a(s_145), .O(gate445inter4));
  nand2 gate1560(.a(gate445inter4), .b(gate445inter3), .O(gate445inter5));
  nor2  gate1561(.a(gate445inter5), .b(gate445inter2), .O(gate445inter6));
  inv1  gate1562(.a(G14), .O(gate445inter7));
  inv1  gate1563(.a(G1171), .O(gate445inter8));
  nand2 gate1564(.a(gate445inter8), .b(gate445inter7), .O(gate445inter9));
  nand2 gate1565(.a(s_145), .b(gate445inter3), .O(gate445inter10));
  nor2  gate1566(.a(gate445inter10), .b(gate445inter9), .O(gate445inter11));
  nor2  gate1567(.a(gate445inter11), .b(gate445inter6), .O(gate445inter12));
  nand2 gate1568(.a(gate445inter12), .b(gate445inter1), .O(G1254));

  xor2  gate2185(.a(G1171), .b(G1075), .O(gate446inter0));
  nand2 gate2186(.a(gate446inter0), .b(s_234), .O(gate446inter1));
  and2  gate2187(.a(G1171), .b(G1075), .O(gate446inter2));
  inv1  gate2188(.a(s_234), .O(gate446inter3));
  inv1  gate2189(.a(s_235), .O(gate446inter4));
  nand2 gate2190(.a(gate446inter4), .b(gate446inter3), .O(gate446inter5));
  nor2  gate2191(.a(gate446inter5), .b(gate446inter2), .O(gate446inter6));
  inv1  gate2192(.a(G1075), .O(gate446inter7));
  inv1  gate2193(.a(G1171), .O(gate446inter8));
  nand2 gate2194(.a(gate446inter8), .b(gate446inter7), .O(gate446inter9));
  nand2 gate2195(.a(s_235), .b(gate446inter3), .O(gate446inter10));
  nor2  gate2196(.a(gate446inter10), .b(gate446inter9), .O(gate446inter11));
  nor2  gate2197(.a(gate446inter11), .b(gate446inter6), .O(gate446inter12));
  nand2 gate2198(.a(gate446inter12), .b(gate446inter1), .O(G1255));
nand2 gate447( .a(G15), .b(G1174), .O(G1256) );
nand2 gate448( .a(G1078), .b(G1174), .O(G1257) );

  xor2  gate2031(.a(G1177), .b(G16), .O(gate449inter0));
  nand2 gate2032(.a(gate449inter0), .b(s_212), .O(gate449inter1));
  and2  gate2033(.a(G1177), .b(G16), .O(gate449inter2));
  inv1  gate2034(.a(s_212), .O(gate449inter3));
  inv1  gate2035(.a(s_213), .O(gate449inter4));
  nand2 gate2036(.a(gate449inter4), .b(gate449inter3), .O(gate449inter5));
  nor2  gate2037(.a(gate449inter5), .b(gate449inter2), .O(gate449inter6));
  inv1  gate2038(.a(G16), .O(gate449inter7));
  inv1  gate2039(.a(G1177), .O(gate449inter8));
  nand2 gate2040(.a(gate449inter8), .b(gate449inter7), .O(gate449inter9));
  nand2 gate2041(.a(s_213), .b(gate449inter3), .O(gate449inter10));
  nor2  gate2042(.a(gate449inter10), .b(gate449inter9), .O(gate449inter11));
  nor2  gate2043(.a(gate449inter11), .b(gate449inter6), .O(gate449inter12));
  nand2 gate2044(.a(gate449inter12), .b(gate449inter1), .O(G1258));
nand2 gate450( .a(G1081), .b(G1177), .O(G1259) );
nand2 gate451( .a(G17), .b(G1180), .O(G1260) );

  xor2  gate1219(.a(G1180), .b(G1084), .O(gate452inter0));
  nand2 gate1220(.a(gate452inter0), .b(s_96), .O(gate452inter1));
  and2  gate1221(.a(G1180), .b(G1084), .O(gate452inter2));
  inv1  gate1222(.a(s_96), .O(gate452inter3));
  inv1  gate1223(.a(s_97), .O(gate452inter4));
  nand2 gate1224(.a(gate452inter4), .b(gate452inter3), .O(gate452inter5));
  nor2  gate1225(.a(gate452inter5), .b(gate452inter2), .O(gate452inter6));
  inv1  gate1226(.a(G1084), .O(gate452inter7));
  inv1  gate1227(.a(G1180), .O(gate452inter8));
  nand2 gate1228(.a(gate452inter8), .b(gate452inter7), .O(gate452inter9));
  nand2 gate1229(.a(s_97), .b(gate452inter3), .O(gate452inter10));
  nor2  gate1230(.a(gate452inter10), .b(gate452inter9), .O(gate452inter11));
  nor2  gate1231(.a(gate452inter11), .b(gate452inter6), .O(gate452inter12));
  nand2 gate1232(.a(gate452inter12), .b(gate452inter1), .O(G1261));
nand2 gate453( .a(G18), .b(G1183), .O(G1262) );
nand2 gate454( .a(G1087), .b(G1183), .O(G1263) );

  xor2  gate995(.a(G1186), .b(G19), .O(gate455inter0));
  nand2 gate996(.a(gate455inter0), .b(s_64), .O(gate455inter1));
  and2  gate997(.a(G1186), .b(G19), .O(gate455inter2));
  inv1  gate998(.a(s_64), .O(gate455inter3));
  inv1  gate999(.a(s_65), .O(gate455inter4));
  nand2 gate1000(.a(gate455inter4), .b(gate455inter3), .O(gate455inter5));
  nor2  gate1001(.a(gate455inter5), .b(gate455inter2), .O(gate455inter6));
  inv1  gate1002(.a(G19), .O(gate455inter7));
  inv1  gate1003(.a(G1186), .O(gate455inter8));
  nand2 gate1004(.a(gate455inter8), .b(gate455inter7), .O(gate455inter9));
  nand2 gate1005(.a(s_65), .b(gate455inter3), .O(gate455inter10));
  nor2  gate1006(.a(gate455inter10), .b(gate455inter9), .O(gate455inter11));
  nor2  gate1007(.a(gate455inter11), .b(gate455inter6), .O(gate455inter12));
  nand2 gate1008(.a(gate455inter12), .b(gate455inter1), .O(G1264));

  xor2  gate1471(.a(G1186), .b(G1090), .O(gate456inter0));
  nand2 gate1472(.a(gate456inter0), .b(s_132), .O(gate456inter1));
  and2  gate1473(.a(G1186), .b(G1090), .O(gate456inter2));
  inv1  gate1474(.a(s_132), .O(gate456inter3));
  inv1  gate1475(.a(s_133), .O(gate456inter4));
  nand2 gate1476(.a(gate456inter4), .b(gate456inter3), .O(gate456inter5));
  nor2  gate1477(.a(gate456inter5), .b(gate456inter2), .O(gate456inter6));
  inv1  gate1478(.a(G1090), .O(gate456inter7));
  inv1  gate1479(.a(G1186), .O(gate456inter8));
  nand2 gate1480(.a(gate456inter8), .b(gate456inter7), .O(gate456inter9));
  nand2 gate1481(.a(s_133), .b(gate456inter3), .O(gate456inter10));
  nor2  gate1482(.a(gate456inter10), .b(gate456inter9), .O(gate456inter11));
  nor2  gate1483(.a(gate456inter11), .b(gate456inter6), .O(gate456inter12));
  nand2 gate1484(.a(gate456inter12), .b(gate456inter1), .O(G1265));

  xor2  gate2493(.a(G1189), .b(G20), .O(gate457inter0));
  nand2 gate2494(.a(gate457inter0), .b(s_278), .O(gate457inter1));
  and2  gate2495(.a(G1189), .b(G20), .O(gate457inter2));
  inv1  gate2496(.a(s_278), .O(gate457inter3));
  inv1  gate2497(.a(s_279), .O(gate457inter4));
  nand2 gate2498(.a(gate457inter4), .b(gate457inter3), .O(gate457inter5));
  nor2  gate2499(.a(gate457inter5), .b(gate457inter2), .O(gate457inter6));
  inv1  gate2500(.a(G20), .O(gate457inter7));
  inv1  gate2501(.a(G1189), .O(gate457inter8));
  nand2 gate2502(.a(gate457inter8), .b(gate457inter7), .O(gate457inter9));
  nand2 gate2503(.a(s_279), .b(gate457inter3), .O(gate457inter10));
  nor2  gate2504(.a(gate457inter10), .b(gate457inter9), .O(gate457inter11));
  nor2  gate2505(.a(gate457inter11), .b(gate457inter6), .O(gate457inter12));
  nand2 gate2506(.a(gate457inter12), .b(gate457inter1), .O(G1266));

  xor2  gate1345(.a(G1189), .b(G1093), .O(gate458inter0));
  nand2 gate1346(.a(gate458inter0), .b(s_114), .O(gate458inter1));
  and2  gate1347(.a(G1189), .b(G1093), .O(gate458inter2));
  inv1  gate1348(.a(s_114), .O(gate458inter3));
  inv1  gate1349(.a(s_115), .O(gate458inter4));
  nand2 gate1350(.a(gate458inter4), .b(gate458inter3), .O(gate458inter5));
  nor2  gate1351(.a(gate458inter5), .b(gate458inter2), .O(gate458inter6));
  inv1  gate1352(.a(G1093), .O(gate458inter7));
  inv1  gate1353(.a(G1189), .O(gate458inter8));
  nand2 gate1354(.a(gate458inter8), .b(gate458inter7), .O(gate458inter9));
  nand2 gate1355(.a(s_115), .b(gate458inter3), .O(gate458inter10));
  nor2  gate1356(.a(gate458inter10), .b(gate458inter9), .O(gate458inter11));
  nor2  gate1357(.a(gate458inter11), .b(gate458inter6), .O(gate458inter12));
  nand2 gate1358(.a(gate458inter12), .b(gate458inter1), .O(G1267));

  xor2  gate561(.a(G1192), .b(G21), .O(gate459inter0));
  nand2 gate562(.a(gate459inter0), .b(s_2), .O(gate459inter1));
  and2  gate563(.a(G1192), .b(G21), .O(gate459inter2));
  inv1  gate564(.a(s_2), .O(gate459inter3));
  inv1  gate565(.a(s_3), .O(gate459inter4));
  nand2 gate566(.a(gate459inter4), .b(gate459inter3), .O(gate459inter5));
  nor2  gate567(.a(gate459inter5), .b(gate459inter2), .O(gate459inter6));
  inv1  gate568(.a(G21), .O(gate459inter7));
  inv1  gate569(.a(G1192), .O(gate459inter8));
  nand2 gate570(.a(gate459inter8), .b(gate459inter7), .O(gate459inter9));
  nand2 gate571(.a(s_3), .b(gate459inter3), .O(gate459inter10));
  nor2  gate572(.a(gate459inter10), .b(gate459inter9), .O(gate459inter11));
  nor2  gate573(.a(gate459inter11), .b(gate459inter6), .O(gate459inter12));
  nand2 gate574(.a(gate459inter12), .b(gate459inter1), .O(G1268));

  xor2  gate1429(.a(G1192), .b(G1096), .O(gate460inter0));
  nand2 gate1430(.a(gate460inter0), .b(s_126), .O(gate460inter1));
  and2  gate1431(.a(G1192), .b(G1096), .O(gate460inter2));
  inv1  gate1432(.a(s_126), .O(gate460inter3));
  inv1  gate1433(.a(s_127), .O(gate460inter4));
  nand2 gate1434(.a(gate460inter4), .b(gate460inter3), .O(gate460inter5));
  nor2  gate1435(.a(gate460inter5), .b(gate460inter2), .O(gate460inter6));
  inv1  gate1436(.a(G1096), .O(gate460inter7));
  inv1  gate1437(.a(G1192), .O(gate460inter8));
  nand2 gate1438(.a(gate460inter8), .b(gate460inter7), .O(gate460inter9));
  nand2 gate1439(.a(s_127), .b(gate460inter3), .O(gate460inter10));
  nor2  gate1440(.a(gate460inter10), .b(gate460inter9), .O(gate460inter11));
  nor2  gate1441(.a(gate460inter11), .b(gate460inter6), .O(gate460inter12));
  nand2 gate1442(.a(gate460inter12), .b(gate460inter1), .O(G1269));
nand2 gate461( .a(G22), .b(G1195), .O(G1270) );
nand2 gate462( .a(G1099), .b(G1195), .O(G1271) );
nand2 gate463( .a(G23), .b(G1198), .O(G1272) );
nand2 gate464( .a(G1102), .b(G1198), .O(G1273) );
nand2 gate465( .a(G24), .b(G1201), .O(G1274) );
nand2 gate466( .a(G1105), .b(G1201), .O(G1275) );

  xor2  gate1037(.a(G1204), .b(G25), .O(gate467inter0));
  nand2 gate1038(.a(gate467inter0), .b(s_70), .O(gate467inter1));
  and2  gate1039(.a(G1204), .b(G25), .O(gate467inter2));
  inv1  gate1040(.a(s_70), .O(gate467inter3));
  inv1  gate1041(.a(s_71), .O(gate467inter4));
  nand2 gate1042(.a(gate467inter4), .b(gate467inter3), .O(gate467inter5));
  nor2  gate1043(.a(gate467inter5), .b(gate467inter2), .O(gate467inter6));
  inv1  gate1044(.a(G25), .O(gate467inter7));
  inv1  gate1045(.a(G1204), .O(gate467inter8));
  nand2 gate1046(.a(gate467inter8), .b(gate467inter7), .O(gate467inter9));
  nand2 gate1047(.a(s_71), .b(gate467inter3), .O(gate467inter10));
  nor2  gate1048(.a(gate467inter10), .b(gate467inter9), .O(gate467inter11));
  nor2  gate1049(.a(gate467inter11), .b(gate467inter6), .O(gate467inter12));
  nand2 gate1050(.a(gate467inter12), .b(gate467inter1), .O(G1276));
nand2 gate468( .a(G1108), .b(G1204), .O(G1277) );
nand2 gate469( .a(G26), .b(G1207), .O(G1278) );
nand2 gate470( .a(G1111), .b(G1207), .O(G1279) );
nand2 gate471( .a(G27), .b(G1210), .O(G1280) );
nand2 gate472( .a(G1114), .b(G1210), .O(G1281) );
nand2 gate473( .a(G28), .b(G1213), .O(G1282) );
nand2 gate474( .a(G1117), .b(G1213), .O(G1283) );
nand2 gate475( .a(G29), .b(G1216), .O(G1284) );
nand2 gate476( .a(G1120), .b(G1216), .O(G1285) );

  xor2  gate855(.a(G1219), .b(G30), .O(gate477inter0));
  nand2 gate856(.a(gate477inter0), .b(s_44), .O(gate477inter1));
  and2  gate857(.a(G1219), .b(G30), .O(gate477inter2));
  inv1  gate858(.a(s_44), .O(gate477inter3));
  inv1  gate859(.a(s_45), .O(gate477inter4));
  nand2 gate860(.a(gate477inter4), .b(gate477inter3), .O(gate477inter5));
  nor2  gate861(.a(gate477inter5), .b(gate477inter2), .O(gate477inter6));
  inv1  gate862(.a(G30), .O(gate477inter7));
  inv1  gate863(.a(G1219), .O(gate477inter8));
  nand2 gate864(.a(gate477inter8), .b(gate477inter7), .O(gate477inter9));
  nand2 gate865(.a(s_45), .b(gate477inter3), .O(gate477inter10));
  nor2  gate866(.a(gate477inter10), .b(gate477inter9), .O(gate477inter11));
  nor2  gate867(.a(gate477inter11), .b(gate477inter6), .O(gate477inter12));
  nand2 gate868(.a(gate477inter12), .b(gate477inter1), .O(G1286));

  xor2  gate2381(.a(G1219), .b(G1123), .O(gate478inter0));
  nand2 gate2382(.a(gate478inter0), .b(s_262), .O(gate478inter1));
  and2  gate2383(.a(G1219), .b(G1123), .O(gate478inter2));
  inv1  gate2384(.a(s_262), .O(gate478inter3));
  inv1  gate2385(.a(s_263), .O(gate478inter4));
  nand2 gate2386(.a(gate478inter4), .b(gate478inter3), .O(gate478inter5));
  nor2  gate2387(.a(gate478inter5), .b(gate478inter2), .O(gate478inter6));
  inv1  gate2388(.a(G1123), .O(gate478inter7));
  inv1  gate2389(.a(G1219), .O(gate478inter8));
  nand2 gate2390(.a(gate478inter8), .b(gate478inter7), .O(gate478inter9));
  nand2 gate2391(.a(s_263), .b(gate478inter3), .O(gate478inter10));
  nor2  gate2392(.a(gate478inter10), .b(gate478inter9), .O(gate478inter11));
  nor2  gate2393(.a(gate478inter11), .b(gate478inter6), .O(gate478inter12));
  nand2 gate2394(.a(gate478inter12), .b(gate478inter1), .O(G1287));

  xor2  gate2801(.a(G1222), .b(G31), .O(gate479inter0));
  nand2 gate2802(.a(gate479inter0), .b(s_322), .O(gate479inter1));
  and2  gate2803(.a(G1222), .b(G31), .O(gate479inter2));
  inv1  gate2804(.a(s_322), .O(gate479inter3));
  inv1  gate2805(.a(s_323), .O(gate479inter4));
  nand2 gate2806(.a(gate479inter4), .b(gate479inter3), .O(gate479inter5));
  nor2  gate2807(.a(gate479inter5), .b(gate479inter2), .O(gate479inter6));
  inv1  gate2808(.a(G31), .O(gate479inter7));
  inv1  gate2809(.a(G1222), .O(gate479inter8));
  nand2 gate2810(.a(gate479inter8), .b(gate479inter7), .O(gate479inter9));
  nand2 gate2811(.a(s_323), .b(gate479inter3), .O(gate479inter10));
  nor2  gate2812(.a(gate479inter10), .b(gate479inter9), .O(gate479inter11));
  nor2  gate2813(.a(gate479inter11), .b(gate479inter6), .O(gate479inter12));
  nand2 gate2814(.a(gate479inter12), .b(gate479inter1), .O(G1288));
nand2 gate480( .a(G1126), .b(G1222), .O(G1289) );
nand2 gate481( .a(G32), .b(G1225), .O(G1290) );
nand2 gate482( .a(G1129), .b(G1225), .O(G1291) );

  xor2  gate925(.a(G1229), .b(G1228), .O(gate483inter0));
  nand2 gate926(.a(gate483inter0), .b(s_54), .O(gate483inter1));
  and2  gate927(.a(G1229), .b(G1228), .O(gate483inter2));
  inv1  gate928(.a(s_54), .O(gate483inter3));
  inv1  gate929(.a(s_55), .O(gate483inter4));
  nand2 gate930(.a(gate483inter4), .b(gate483inter3), .O(gate483inter5));
  nor2  gate931(.a(gate483inter5), .b(gate483inter2), .O(gate483inter6));
  inv1  gate932(.a(G1228), .O(gate483inter7));
  inv1  gate933(.a(G1229), .O(gate483inter8));
  nand2 gate934(.a(gate483inter8), .b(gate483inter7), .O(gate483inter9));
  nand2 gate935(.a(s_55), .b(gate483inter3), .O(gate483inter10));
  nor2  gate936(.a(gate483inter10), .b(gate483inter9), .O(gate483inter11));
  nor2  gate937(.a(gate483inter11), .b(gate483inter6), .O(gate483inter12));
  nand2 gate938(.a(gate483inter12), .b(gate483inter1), .O(G1292));
nand2 gate484( .a(G1230), .b(G1231), .O(G1293) );
nand2 gate485( .a(G1232), .b(G1233), .O(G1294) );

  xor2  gate659(.a(G1235), .b(G1234), .O(gate486inter0));
  nand2 gate660(.a(gate486inter0), .b(s_16), .O(gate486inter1));
  and2  gate661(.a(G1235), .b(G1234), .O(gate486inter2));
  inv1  gate662(.a(s_16), .O(gate486inter3));
  inv1  gate663(.a(s_17), .O(gate486inter4));
  nand2 gate664(.a(gate486inter4), .b(gate486inter3), .O(gate486inter5));
  nor2  gate665(.a(gate486inter5), .b(gate486inter2), .O(gate486inter6));
  inv1  gate666(.a(G1234), .O(gate486inter7));
  inv1  gate667(.a(G1235), .O(gate486inter8));
  nand2 gate668(.a(gate486inter8), .b(gate486inter7), .O(gate486inter9));
  nand2 gate669(.a(s_17), .b(gate486inter3), .O(gate486inter10));
  nor2  gate670(.a(gate486inter10), .b(gate486inter9), .O(gate486inter11));
  nor2  gate671(.a(gate486inter11), .b(gate486inter6), .O(gate486inter12));
  nand2 gate672(.a(gate486inter12), .b(gate486inter1), .O(G1295));

  xor2  gate1331(.a(G1237), .b(G1236), .O(gate487inter0));
  nand2 gate1332(.a(gate487inter0), .b(s_112), .O(gate487inter1));
  and2  gate1333(.a(G1237), .b(G1236), .O(gate487inter2));
  inv1  gate1334(.a(s_112), .O(gate487inter3));
  inv1  gate1335(.a(s_113), .O(gate487inter4));
  nand2 gate1336(.a(gate487inter4), .b(gate487inter3), .O(gate487inter5));
  nor2  gate1337(.a(gate487inter5), .b(gate487inter2), .O(gate487inter6));
  inv1  gate1338(.a(G1236), .O(gate487inter7));
  inv1  gate1339(.a(G1237), .O(gate487inter8));
  nand2 gate1340(.a(gate487inter8), .b(gate487inter7), .O(gate487inter9));
  nand2 gate1341(.a(s_113), .b(gate487inter3), .O(gate487inter10));
  nor2  gate1342(.a(gate487inter10), .b(gate487inter9), .O(gate487inter11));
  nor2  gate1343(.a(gate487inter11), .b(gate487inter6), .O(gate487inter12));
  nand2 gate1344(.a(gate487inter12), .b(gate487inter1), .O(G1296));
nand2 gate488( .a(G1238), .b(G1239), .O(G1297) );

  xor2  gate575(.a(G1241), .b(G1240), .O(gate489inter0));
  nand2 gate576(.a(gate489inter0), .b(s_4), .O(gate489inter1));
  and2  gate577(.a(G1241), .b(G1240), .O(gate489inter2));
  inv1  gate578(.a(s_4), .O(gate489inter3));
  inv1  gate579(.a(s_5), .O(gate489inter4));
  nand2 gate580(.a(gate489inter4), .b(gate489inter3), .O(gate489inter5));
  nor2  gate581(.a(gate489inter5), .b(gate489inter2), .O(gate489inter6));
  inv1  gate582(.a(G1240), .O(gate489inter7));
  inv1  gate583(.a(G1241), .O(gate489inter8));
  nand2 gate584(.a(gate489inter8), .b(gate489inter7), .O(gate489inter9));
  nand2 gate585(.a(s_5), .b(gate489inter3), .O(gate489inter10));
  nor2  gate586(.a(gate489inter10), .b(gate489inter9), .O(gate489inter11));
  nor2  gate587(.a(gate489inter11), .b(gate489inter6), .O(gate489inter12));
  nand2 gate588(.a(gate489inter12), .b(gate489inter1), .O(G1298));
nand2 gate490( .a(G1242), .b(G1243), .O(G1299) );
nand2 gate491( .a(G1244), .b(G1245), .O(G1300) );
nand2 gate492( .a(G1246), .b(G1247), .O(G1301) );
nand2 gate493( .a(G1248), .b(G1249), .O(G1302) );
nand2 gate494( .a(G1250), .b(G1251), .O(G1303) );
nand2 gate495( .a(G1252), .b(G1253), .O(G1304) );

  xor2  gate2157(.a(G1255), .b(G1254), .O(gate496inter0));
  nand2 gate2158(.a(gate496inter0), .b(s_230), .O(gate496inter1));
  and2  gate2159(.a(G1255), .b(G1254), .O(gate496inter2));
  inv1  gate2160(.a(s_230), .O(gate496inter3));
  inv1  gate2161(.a(s_231), .O(gate496inter4));
  nand2 gate2162(.a(gate496inter4), .b(gate496inter3), .O(gate496inter5));
  nor2  gate2163(.a(gate496inter5), .b(gate496inter2), .O(gate496inter6));
  inv1  gate2164(.a(G1254), .O(gate496inter7));
  inv1  gate2165(.a(G1255), .O(gate496inter8));
  nand2 gate2166(.a(gate496inter8), .b(gate496inter7), .O(gate496inter9));
  nand2 gate2167(.a(s_231), .b(gate496inter3), .O(gate496inter10));
  nor2  gate2168(.a(gate496inter10), .b(gate496inter9), .O(gate496inter11));
  nor2  gate2169(.a(gate496inter11), .b(gate496inter6), .O(gate496inter12));
  nand2 gate2170(.a(gate496inter12), .b(gate496inter1), .O(G1305));
nand2 gate497( .a(G1256), .b(G1257), .O(G1306) );
nand2 gate498( .a(G1258), .b(G1259), .O(G1307) );
nand2 gate499( .a(G1260), .b(G1261), .O(G1308) );
nand2 gate500( .a(G1262), .b(G1263), .O(G1309) );
nand2 gate501( .a(G1264), .b(G1265), .O(G1310) );

  xor2  gate2423(.a(G1267), .b(G1266), .O(gate502inter0));
  nand2 gate2424(.a(gate502inter0), .b(s_268), .O(gate502inter1));
  and2  gate2425(.a(G1267), .b(G1266), .O(gate502inter2));
  inv1  gate2426(.a(s_268), .O(gate502inter3));
  inv1  gate2427(.a(s_269), .O(gate502inter4));
  nand2 gate2428(.a(gate502inter4), .b(gate502inter3), .O(gate502inter5));
  nor2  gate2429(.a(gate502inter5), .b(gate502inter2), .O(gate502inter6));
  inv1  gate2430(.a(G1266), .O(gate502inter7));
  inv1  gate2431(.a(G1267), .O(gate502inter8));
  nand2 gate2432(.a(gate502inter8), .b(gate502inter7), .O(gate502inter9));
  nand2 gate2433(.a(s_269), .b(gate502inter3), .O(gate502inter10));
  nor2  gate2434(.a(gate502inter10), .b(gate502inter9), .O(gate502inter11));
  nor2  gate2435(.a(gate502inter11), .b(gate502inter6), .O(gate502inter12));
  nand2 gate2436(.a(gate502inter12), .b(gate502inter1), .O(G1311));
nand2 gate503( .a(G1268), .b(G1269), .O(G1312) );

  xor2  gate1849(.a(G1271), .b(G1270), .O(gate504inter0));
  nand2 gate1850(.a(gate504inter0), .b(s_186), .O(gate504inter1));
  and2  gate1851(.a(G1271), .b(G1270), .O(gate504inter2));
  inv1  gate1852(.a(s_186), .O(gate504inter3));
  inv1  gate1853(.a(s_187), .O(gate504inter4));
  nand2 gate1854(.a(gate504inter4), .b(gate504inter3), .O(gate504inter5));
  nor2  gate1855(.a(gate504inter5), .b(gate504inter2), .O(gate504inter6));
  inv1  gate1856(.a(G1270), .O(gate504inter7));
  inv1  gate1857(.a(G1271), .O(gate504inter8));
  nand2 gate1858(.a(gate504inter8), .b(gate504inter7), .O(gate504inter9));
  nand2 gate1859(.a(s_187), .b(gate504inter3), .O(gate504inter10));
  nor2  gate1860(.a(gate504inter10), .b(gate504inter9), .O(gate504inter11));
  nor2  gate1861(.a(gate504inter11), .b(gate504inter6), .O(gate504inter12));
  nand2 gate1862(.a(gate504inter12), .b(gate504inter1), .O(G1313));
nand2 gate505( .a(G1272), .b(G1273), .O(G1314) );

  xor2  gate743(.a(G1275), .b(G1274), .O(gate506inter0));
  nand2 gate744(.a(gate506inter0), .b(s_28), .O(gate506inter1));
  and2  gate745(.a(G1275), .b(G1274), .O(gate506inter2));
  inv1  gate746(.a(s_28), .O(gate506inter3));
  inv1  gate747(.a(s_29), .O(gate506inter4));
  nand2 gate748(.a(gate506inter4), .b(gate506inter3), .O(gate506inter5));
  nor2  gate749(.a(gate506inter5), .b(gate506inter2), .O(gate506inter6));
  inv1  gate750(.a(G1274), .O(gate506inter7));
  inv1  gate751(.a(G1275), .O(gate506inter8));
  nand2 gate752(.a(gate506inter8), .b(gate506inter7), .O(gate506inter9));
  nand2 gate753(.a(s_29), .b(gate506inter3), .O(gate506inter10));
  nor2  gate754(.a(gate506inter10), .b(gate506inter9), .O(gate506inter11));
  nor2  gate755(.a(gate506inter11), .b(gate506inter6), .O(gate506inter12));
  nand2 gate756(.a(gate506inter12), .b(gate506inter1), .O(G1315));
nand2 gate507( .a(G1276), .b(G1277), .O(G1316) );

  xor2  gate589(.a(G1279), .b(G1278), .O(gate508inter0));
  nand2 gate590(.a(gate508inter0), .b(s_6), .O(gate508inter1));
  and2  gate591(.a(G1279), .b(G1278), .O(gate508inter2));
  inv1  gate592(.a(s_6), .O(gate508inter3));
  inv1  gate593(.a(s_7), .O(gate508inter4));
  nand2 gate594(.a(gate508inter4), .b(gate508inter3), .O(gate508inter5));
  nor2  gate595(.a(gate508inter5), .b(gate508inter2), .O(gate508inter6));
  inv1  gate596(.a(G1278), .O(gate508inter7));
  inv1  gate597(.a(G1279), .O(gate508inter8));
  nand2 gate598(.a(gate508inter8), .b(gate508inter7), .O(gate508inter9));
  nand2 gate599(.a(s_7), .b(gate508inter3), .O(gate508inter10));
  nor2  gate600(.a(gate508inter10), .b(gate508inter9), .O(gate508inter11));
  nor2  gate601(.a(gate508inter11), .b(gate508inter6), .O(gate508inter12));
  nand2 gate602(.a(gate508inter12), .b(gate508inter1), .O(G1317));
nand2 gate509( .a(G1280), .b(G1281), .O(G1318) );

  xor2  gate631(.a(G1283), .b(G1282), .O(gate510inter0));
  nand2 gate632(.a(gate510inter0), .b(s_12), .O(gate510inter1));
  and2  gate633(.a(G1283), .b(G1282), .O(gate510inter2));
  inv1  gate634(.a(s_12), .O(gate510inter3));
  inv1  gate635(.a(s_13), .O(gate510inter4));
  nand2 gate636(.a(gate510inter4), .b(gate510inter3), .O(gate510inter5));
  nor2  gate637(.a(gate510inter5), .b(gate510inter2), .O(gate510inter6));
  inv1  gate638(.a(G1282), .O(gate510inter7));
  inv1  gate639(.a(G1283), .O(gate510inter8));
  nand2 gate640(.a(gate510inter8), .b(gate510inter7), .O(gate510inter9));
  nand2 gate641(.a(s_13), .b(gate510inter3), .O(gate510inter10));
  nor2  gate642(.a(gate510inter10), .b(gate510inter9), .O(gate510inter11));
  nor2  gate643(.a(gate510inter11), .b(gate510inter6), .O(gate510inter12));
  nand2 gate644(.a(gate510inter12), .b(gate510inter1), .O(G1319));
nand2 gate511( .a(G1284), .b(G1285), .O(G1320) );

  xor2  gate2689(.a(G1287), .b(G1286), .O(gate512inter0));
  nand2 gate2690(.a(gate512inter0), .b(s_306), .O(gate512inter1));
  and2  gate2691(.a(G1287), .b(G1286), .O(gate512inter2));
  inv1  gate2692(.a(s_306), .O(gate512inter3));
  inv1  gate2693(.a(s_307), .O(gate512inter4));
  nand2 gate2694(.a(gate512inter4), .b(gate512inter3), .O(gate512inter5));
  nor2  gate2695(.a(gate512inter5), .b(gate512inter2), .O(gate512inter6));
  inv1  gate2696(.a(G1286), .O(gate512inter7));
  inv1  gate2697(.a(G1287), .O(gate512inter8));
  nand2 gate2698(.a(gate512inter8), .b(gate512inter7), .O(gate512inter9));
  nand2 gate2699(.a(s_307), .b(gate512inter3), .O(gate512inter10));
  nor2  gate2700(.a(gate512inter10), .b(gate512inter9), .O(gate512inter11));
  nor2  gate2701(.a(gate512inter11), .b(gate512inter6), .O(gate512inter12));
  nand2 gate2702(.a(gate512inter12), .b(gate512inter1), .O(G1321));
nand2 gate513( .a(G1288), .b(G1289), .O(G1322) );
nand2 gate514( .a(G1290), .b(G1291), .O(G1323) );
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule