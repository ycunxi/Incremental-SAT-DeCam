module c432 (N1,N4,N8,N11,N14,N17,N21,N24,N27,N30,
             N34,N37,N40,N43,N47,N50,N53,N56,N60,N63,
             N66,N69,N73,N76,N79,N82,N86,N89,N92,N95,
             N99,N102,N105,N108,N112,N115,N223,N329,N370,N421,
             N430,N431,N432);

input N1,N4,N8,N11,N14,N17,N21,N24,N27,N30,
      N34,N37,N40,N43,N47,N50,N53,N56,N60,N63,
      N66,N69,N73,N76,N79,N82,N86,N89,N92,N95,
      N99,N102,N105,N108,N112,N115;//RE__PI;

input s_0,s_1;//RE__ALLOW(00,01,10,11);
input s_2,s_3;//RE__ALLOW(00,01,10,11);
input s_4,s_5;//RE__ALLOW(00,01,10,11);
input s_6,s_7;//RE__ALLOW(00,01,10,11);
input s_8,s_9;//RE__ALLOW(00,01,10,11);
input s_10,s_11;//RE__ALLOW(00,01,10,11);
input s_12,s_13;//RE__ALLOW(00,01,10,11);
input s_14,s_15;//RE__ALLOW(00,01,10,11);
input s_16,s_17;//RE__ALLOW(00,01,10,11);
input s_18,s_19;//RE__ALLOW(00,01,10,11);
input s_20,s_21;//RE__ALLOW(00,01,10,11);
input s_22,s_23;//RE__ALLOW(00,01,10,11);
input s_24,s_25;//RE__ALLOW(00,01,10,11);
input s_26,s_27;//RE__ALLOW(00,01,10,11);
input s_28,s_29;//RE__ALLOW(00,01,10,11);
input s_30,s_31;//RE__ALLOW(00,01,10,11);
input s_32,s_33;//RE__ALLOW(00,01,10,11);
input s_34,s_35;//RE__ALLOW(00,01,10,11);
input s_36,s_37;//RE__ALLOW(00,01,10,11);
input s_38,s_39;//RE__ALLOW(00,01,10,11);
input s_40,s_41;//RE__ALLOW(00,01,10,11);
input s_42,s_43;//RE__ALLOW(00,01,10,11);
input s_44,s_45;//RE__ALLOW(00,01,10,11);
input s_46,s_47;//RE__ALLOW(00,01,10,11);
input s_48,s_49;//RE__ALLOW(00,01,10,11);
input s_50,s_51;//RE__ALLOW(00,01,10,11);
output N223,N329,N370,N421,N430,N431,N432;

wire N118,N119,N122,N123,N126,N127,N130,N131,N134,N135,
     N138,N139,N142,N143,N146,N147,N150,N151,N154,N157,
     N158,N159,N162,N165,N168,N171,N174,N177,N180,N183,
     N184,N185,N186,N187,N188,N189,N190,N191,N192,N193,
     N194,N195,N196,N197,N198,N199,N203,N213,N224,N227,
     N230,N233,N236,N239,N242,N243,N246,N247,N250,N251,
     N254,N255,N256,N257,N258,N259,N260,N263,N264,N267,
     N270,N273,N276,N279,N282,N285,N288,N289,N290,N291,
     N292,N293,N294,N295,N296,N300,N301,N302,N303,N304,
     N305,N306,N307,N308,N309,N319,N330,N331,N332,N333,
     N334,N335,N336,N337,N338,N339,N340,N341,N342,N343,
     N344,N345,N346,N347,N348,N349,N350,N351,N352,N353,
     N354,N355,N356,N357,N360,N371,N372,N373,N374,N375,
     N376,N377,N378,N379,N380,N381,N386,N393,N399,N404,
     N407,N411,N414,N415,N416,N417,N418,N419,N420,N422,
     N425,N428,N429, gate30inter0, gate30inter1, gate30inter2, gate30inter3, gate30inter4, gate30inter5, gate30inter6, gate30inter7, gate30inter8, gate30inter9, gate30inter10, gate30inter11, gate30inter12, gate71inter0, gate71inter1, gate71inter2, gate71inter3, gate71inter4, gate71inter5, gate71inter6, gate71inter7, gate71inter8, gate71inter9, gate71inter10, gate71inter11, gate71inter12, gate108inter0, gate108inter1, gate108inter2, gate108inter3, gate108inter4, gate108inter5, gate108inter6, gate108inter7, gate108inter8, gate108inter9, gate108inter10, gate108inter11, gate108inter12, gate114inter0, gate114inter1, gate114inter2, gate114inter3, gate114inter4, gate114inter5, gate114inter6, gate114inter7, gate114inter8, gate114inter9, gate114inter10, gate114inter11, gate114inter12, gate130inter0, gate130inter1, gate130inter2, gate130inter3, gate130inter4, gate130inter5, gate130inter6, gate130inter7, gate130inter8, gate130inter9, gate130inter10, gate130inter11, gate130inter12, gate72inter0, gate72inter1, gate72inter2, gate72inter3, gate72inter4, gate72inter5, gate72inter6, gate72inter7, gate72inter8, gate72inter9, gate72inter10, gate72inter11, gate72inter12, gate70inter0, gate70inter1, gate70inter2, gate70inter3, gate70inter4, gate70inter5, gate70inter6, gate70inter7, gate70inter8, gate70inter9, gate70inter10, gate70inter11, gate70inter12, gate36inter0, gate36inter1, gate36inter2, gate36inter3, gate36inter4, gate36inter5, gate36inter6, gate36inter7, gate36inter8, gate36inter9, gate36inter10, gate36inter11, gate36inter12, gate82inter0, gate82inter1, gate82inter2, gate82inter3, gate82inter4, gate82inter5, gate82inter6, gate82inter7, gate82inter8, gate82inter9, gate82inter10, gate82inter11, gate82inter12, gate42inter0, gate42inter1, gate42inter2, gate42inter3, gate42inter4, gate42inter5, gate42inter6, gate42inter7, gate42inter8, gate42inter9, gate42inter10, gate42inter11, gate42inter12, gate57inter0, gate57inter1, gate57inter2, gate57inter3, gate57inter4, gate57inter5, gate57inter6, gate57inter7, gate57inter8, gate57inter9, gate57inter10, gate57inter11, gate57inter12, gate116inter0, gate116inter1, gate116inter2, gate116inter3, gate116inter4, gate116inter5, gate116inter6, gate116inter7, gate116inter8, gate116inter9, gate116inter10, gate116inter11, gate116inter12, gate85inter0, gate85inter1, gate85inter2, gate85inter3, gate85inter4, gate85inter5, gate85inter6, gate85inter7, gate85inter8, gate85inter9, gate85inter10, gate85inter11, gate85inter12, gate59inter0, gate59inter1, gate59inter2, gate59inter3, gate59inter4, gate59inter5, gate59inter6, gate59inter7, gate59inter8, gate59inter9, gate59inter10, gate59inter11, gate59inter12, gate101inter0, gate101inter1, gate101inter2, gate101inter3, gate101inter4, gate101inter5, gate101inter6, gate101inter7, gate101inter8, gate101inter9, gate101inter10, gate101inter11, gate101inter12, gate37inter0, gate37inter1, gate37inter2, gate37inter3, gate37inter4, gate37inter5, gate37inter6, gate37inter7, gate37inter8, gate37inter9, gate37inter10, gate37inter11, gate37inter12, gate131inter0, gate131inter1, gate131inter2, gate131inter3, gate131inter4, gate131inter5, gate131inter6, gate131inter7, gate131inter8, gate131inter9, gate131inter10, gate131inter11, gate131inter12, gate132inter0, gate132inter1, gate132inter2, gate132inter3, gate132inter4, gate132inter5, gate132inter6, gate132inter7, gate132inter8, gate132inter9, gate132inter10, gate132inter11, gate132inter12, gate135inter0, gate135inter1, gate135inter2, gate135inter3, gate135inter4, gate135inter5, gate135inter6, gate135inter7, gate135inter8, gate135inter9, gate135inter10, gate135inter11, gate135inter12, gate28inter0, gate28inter1, gate28inter2, gate28inter3, gate28inter4, gate28inter5, gate28inter6, gate28inter7, gate28inter8, gate28inter9, gate28inter10, gate28inter11, gate28inter12, gate104inter0, gate104inter1, gate104inter2, gate104inter3, gate104inter4, gate104inter5, gate104inter6, gate104inter7, gate104inter8, gate104inter9, gate104inter10, gate104inter11, gate104inter12, gate65inter0, gate65inter1, gate65inter2, gate65inter3, gate65inter4, gate65inter5, gate65inter6, gate65inter7, gate65inter8, gate65inter9, gate65inter10, gate65inter11, gate65inter12, gate25inter0, gate25inter1, gate25inter2, gate25inter3, gate25inter4, gate25inter5, gate25inter6, gate25inter7, gate25inter8, gate25inter9, gate25inter10, gate25inter11, gate25inter12, gate154inter0, gate154inter1, gate154inter2, gate154inter3, gate154inter4, gate154inter5, gate154inter6, gate154inter7, gate154inter8, gate154inter9, gate154inter10, gate154inter11, gate154inter12, gate68inter0, gate68inter1, gate68inter2, gate68inter3, gate68inter4, gate68inter5, gate68inter6, gate68inter7, gate68inter8, gate68inter9, gate68inter10, gate68inter11, gate68inter12, gate41inter0, gate41inter1, gate41inter2, gate41inter3, gate41inter4, gate41inter5, gate41inter6, gate41inter7, gate41inter8, gate41inter9, gate41inter10, gate41inter11, gate41inter12;



inv1 gate1( .a(N1), .O(N118) );
inv1 gate2( .a(N4), .O(N119) );
inv1 gate3( .a(N11), .O(N122) );
inv1 gate4( .a(N17), .O(N123) );
inv1 gate5( .a(N24), .O(N126) );
inv1 gate6( .a(N30), .O(N127) );
inv1 gate7( .a(N37), .O(N130) );
inv1 gate8( .a(N43), .O(N131) );
inv1 gate9( .a(N50), .O(N134) );
inv1 gate10( .a(N56), .O(N135) );
inv1 gate11( .a(N63), .O(N138) );
inv1 gate12( .a(N69), .O(N139) );
inv1 gate13( .a(N76), .O(N142) );
inv1 gate14( .a(N82), .O(N143) );
inv1 gate15( .a(N89), .O(N146) );
inv1 gate16( .a(N95), .O(N147) );
inv1 gate17( .a(N102), .O(N150) );
inv1 gate18( .a(N108), .O(N151) );
nand2 gate19( .a(N118), .b(N4), .O(N154) );
nor2 gate20( .a(N8), .b(N119), .O(N157) );
nor2 gate21( .a(N14), .b(N119), .O(N158) );
nand2 gate22( .a(N122), .b(N17), .O(N159) );
nand2 gate23( .a(N126), .b(N30), .O(N162) );
nand2 gate24( .a(N130), .b(N43), .O(N165) );

  xor2  gate469(.a(N56), .b(N134), .O(gate25inter0));
  nand2 gate470(.a(gate25inter0), .b(s_44), .O(gate25inter1));
  and2  gate471(.a(N56), .b(N134), .O(gate25inter2));
  inv1  gate472(.a(s_44), .O(gate25inter3));
  inv1  gate473(.a(s_45), .O(gate25inter4));
  nand2 gate474(.a(gate25inter4), .b(gate25inter3), .O(gate25inter5));
  nor2  gate475(.a(gate25inter5), .b(gate25inter2), .O(gate25inter6));
  inv1  gate476(.a(N134), .O(gate25inter7));
  inv1  gate477(.a(N56), .O(gate25inter8));
  nand2 gate478(.a(gate25inter8), .b(gate25inter7), .O(gate25inter9));
  nand2 gate479(.a(s_45), .b(gate25inter3), .O(gate25inter10));
  nor2  gate480(.a(gate25inter10), .b(gate25inter9), .O(gate25inter11));
  nor2  gate481(.a(gate25inter11), .b(gate25inter6), .O(gate25inter12));
  nand2 gate482(.a(gate25inter12), .b(gate25inter1), .O(N168));
nand2 gate26( .a(N138), .b(N69), .O(N171) );
nand2 gate27( .a(N142), .b(N82), .O(N174) );

  xor2  gate427(.a(N95), .b(N146), .O(gate28inter0));
  nand2 gate428(.a(gate28inter0), .b(s_38), .O(gate28inter1));
  and2  gate429(.a(N95), .b(N146), .O(gate28inter2));
  inv1  gate430(.a(s_38), .O(gate28inter3));
  inv1  gate431(.a(s_39), .O(gate28inter4));
  nand2 gate432(.a(gate28inter4), .b(gate28inter3), .O(gate28inter5));
  nor2  gate433(.a(gate28inter5), .b(gate28inter2), .O(gate28inter6));
  inv1  gate434(.a(N146), .O(gate28inter7));
  inv1  gate435(.a(N95), .O(gate28inter8));
  nand2 gate436(.a(gate28inter8), .b(gate28inter7), .O(gate28inter9));
  nand2 gate437(.a(s_39), .b(gate28inter3), .O(gate28inter10));
  nor2  gate438(.a(gate28inter10), .b(gate28inter9), .O(gate28inter11));
  nor2  gate439(.a(gate28inter11), .b(gate28inter6), .O(gate28inter12));
  nand2 gate440(.a(gate28inter12), .b(gate28inter1), .O(N177));
nand2 gate29( .a(N150), .b(N108), .O(N180) );

  xor2  gate161(.a(N123), .b(N21), .O(gate30inter0));
  nand2 gate162(.a(gate30inter0), .b(s_0), .O(gate30inter1));
  and2  gate163(.a(N123), .b(N21), .O(gate30inter2));
  inv1  gate164(.a(s_0), .O(gate30inter3));
  inv1  gate165(.a(s_1), .O(gate30inter4));
  nand2 gate166(.a(gate30inter4), .b(gate30inter3), .O(gate30inter5));
  nor2  gate167(.a(gate30inter5), .b(gate30inter2), .O(gate30inter6));
  inv1  gate168(.a(N21), .O(gate30inter7));
  inv1  gate169(.a(N123), .O(gate30inter8));
  nand2 gate170(.a(gate30inter8), .b(gate30inter7), .O(gate30inter9));
  nand2 gate171(.a(s_1), .b(gate30inter3), .O(gate30inter10));
  nor2  gate172(.a(gate30inter10), .b(gate30inter9), .O(gate30inter11));
  nor2  gate173(.a(gate30inter11), .b(gate30inter6), .O(gate30inter12));
  nand2 gate174(.a(gate30inter12), .b(gate30inter1), .O(N183));
nor2 gate31( .a(N27), .b(N123), .O(N184) );
nor2 gate32( .a(N34), .b(N127), .O(N185) );
nor2 gate33( .a(N40), .b(N127), .O(N186) );
nor2 gate34( .a(N47), .b(N131), .O(N187) );
nor2 gate35( .a(N53), .b(N131), .O(N188) );

  xor2  gate259(.a(N135), .b(N60), .O(gate36inter0));
  nand2 gate260(.a(gate36inter0), .b(s_14), .O(gate36inter1));
  and2  gate261(.a(N135), .b(N60), .O(gate36inter2));
  inv1  gate262(.a(s_14), .O(gate36inter3));
  inv1  gate263(.a(s_15), .O(gate36inter4));
  nand2 gate264(.a(gate36inter4), .b(gate36inter3), .O(gate36inter5));
  nor2  gate265(.a(gate36inter5), .b(gate36inter2), .O(gate36inter6));
  inv1  gate266(.a(N60), .O(gate36inter7));
  inv1  gate267(.a(N135), .O(gate36inter8));
  nand2 gate268(.a(gate36inter8), .b(gate36inter7), .O(gate36inter9));
  nand2 gate269(.a(s_15), .b(gate36inter3), .O(gate36inter10));
  nor2  gate270(.a(gate36inter10), .b(gate36inter9), .O(gate36inter11));
  nor2  gate271(.a(gate36inter11), .b(gate36inter6), .O(gate36inter12));
  nand2 gate272(.a(gate36inter12), .b(gate36inter1), .O(N189));

  xor2  gate371(.a(N135), .b(N66), .O(gate37inter0));
  nand2 gate372(.a(gate37inter0), .b(s_30), .O(gate37inter1));
  and2  gate373(.a(N135), .b(N66), .O(gate37inter2));
  inv1  gate374(.a(s_30), .O(gate37inter3));
  inv1  gate375(.a(s_31), .O(gate37inter4));
  nand2 gate376(.a(gate37inter4), .b(gate37inter3), .O(gate37inter5));
  nor2  gate377(.a(gate37inter5), .b(gate37inter2), .O(gate37inter6));
  inv1  gate378(.a(N66), .O(gate37inter7));
  inv1  gate379(.a(N135), .O(gate37inter8));
  nand2 gate380(.a(gate37inter8), .b(gate37inter7), .O(gate37inter9));
  nand2 gate381(.a(s_31), .b(gate37inter3), .O(gate37inter10));
  nor2  gate382(.a(gate37inter10), .b(gate37inter9), .O(gate37inter11));
  nor2  gate383(.a(gate37inter11), .b(gate37inter6), .O(gate37inter12));
  nand2 gate384(.a(gate37inter12), .b(gate37inter1), .O(N190));
nor2 gate38( .a(N73), .b(N139), .O(N191) );
nor2 gate39( .a(N79), .b(N139), .O(N192) );
nor2 gate40( .a(N86), .b(N143), .O(N193) );

  xor2  gate511(.a(N143), .b(N92), .O(gate41inter0));
  nand2 gate512(.a(gate41inter0), .b(s_50), .O(gate41inter1));
  and2  gate513(.a(N143), .b(N92), .O(gate41inter2));
  inv1  gate514(.a(s_50), .O(gate41inter3));
  inv1  gate515(.a(s_51), .O(gate41inter4));
  nand2 gate516(.a(gate41inter4), .b(gate41inter3), .O(gate41inter5));
  nor2  gate517(.a(gate41inter5), .b(gate41inter2), .O(gate41inter6));
  inv1  gate518(.a(N92), .O(gate41inter7));
  inv1  gate519(.a(N143), .O(gate41inter8));
  nand2 gate520(.a(gate41inter8), .b(gate41inter7), .O(gate41inter9));
  nand2 gate521(.a(s_51), .b(gate41inter3), .O(gate41inter10));
  nor2  gate522(.a(gate41inter10), .b(gate41inter9), .O(gate41inter11));
  nor2  gate523(.a(gate41inter11), .b(gate41inter6), .O(gate41inter12));
  nand2 gate524(.a(gate41inter12), .b(gate41inter1), .O(N194));

  xor2  gate287(.a(N147), .b(N99), .O(gate42inter0));
  nand2 gate288(.a(gate42inter0), .b(s_18), .O(gate42inter1));
  and2  gate289(.a(N147), .b(N99), .O(gate42inter2));
  inv1  gate290(.a(s_18), .O(gate42inter3));
  inv1  gate291(.a(s_19), .O(gate42inter4));
  nand2 gate292(.a(gate42inter4), .b(gate42inter3), .O(gate42inter5));
  nor2  gate293(.a(gate42inter5), .b(gate42inter2), .O(gate42inter6));
  inv1  gate294(.a(N99), .O(gate42inter7));
  inv1  gate295(.a(N147), .O(gate42inter8));
  nand2 gate296(.a(gate42inter8), .b(gate42inter7), .O(gate42inter9));
  nand2 gate297(.a(s_19), .b(gate42inter3), .O(gate42inter10));
  nor2  gate298(.a(gate42inter10), .b(gate42inter9), .O(gate42inter11));
  nor2  gate299(.a(gate42inter11), .b(gate42inter6), .O(gate42inter12));
  nand2 gate300(.a(gate42inter12), .b(gate42inter1), .O(N195));
nor2 gate43( .a(N105), .b(N147), .O(N196) );
nor2 gate44( .a(N112), .b(N151), .O(N197) );
nor2 gate45( .a(N115), .b(N151), .O(N198) );
and9 gate46( .a(N154), .b(N159), .c(N162), .d(N165), .e(N168), .f(N171), .g(N174), .h(N177), .i(N180), .O(N199) );
inv1 gate47( .a(N199), .O(N203) );
inv1 gate48( .a(N199), .O(N213) );
inv1 gate49( .a(N199), .O(N223) );
xor2 gate50( .a(N203), .b(N154), .O(N224) );
xor2 gate51( .a(N203), .b(N159), .O(N227) );
xor2 gate52( .a(N203), .b(N162), .O(N230) );
xor2 gate53( .a(N203), .b(N165), .O(N233) );
xor2 gate54( .a(N203), .b(N168), .O(N236) );
xor2 gate55( .a(N203), .b(N171), .O(N239) );
nand2 gate56( .a(N1), .b(N213), .O(N242) );

  xor2  gate301(.a(N174), .b(N203), .O(gate57inter0));
  nand2 gate302(.a(gate57inter0), .b(s_20), .O(gate57inter1));
  and2  gate303(.a(N174), .b(N203), .O(gate57inter2));
  inv1  gate304(.a(s_20), .O(gate57inter3));
  inv1  gate305(.a(s_21), .O(gate57inter4));
  nand2 gate306(.a(gate57inter4), .b(gate57inter3), .O(gate57inter5));
  nor2  gate307(.a(gate57inter5), .b(gate57inter2), .O(gate57inter6));
  inv1  gate308(.a(N203), .O(gate57inter7));
  inv1  gate309(.a(N174), .O(gate57inter8));
  nand2 gate310(.a(gate57inter8), .b(gate57inter7), .O(gate57inter9));
  nand2 gate311(.a(s_21), .b(gate57inter3), .O(gate57inter10));
  nor2  gate312(.a(gate57inter10), .b(gate57inter9), .O(gate57inter11));
  nor2  gate313(.a(gate57inter11), .b(gate57inter6), .O(gate57inter12));
  nand2 gate314(.a(gate57inter12), .b(gate57inter1), .O(N243));
nand2 gate58( .a(N213), .b(N11), .O(N246) );

  xor2  gate343(.a(N177), .b(N203), .O(gate59inter0));
  nand2 gate344(.a(gate59inter0), .b(s_26), .O(gate59inter1));
  and2  gate345(.a(N177), .b(N203), .O(gate59inter2));
  inv1  gate346(.a(s_26), .O(gate59inter3));
  inv1  gate347(.a(s_27), .O(gate59inter4));
  nand2 gate348(.a(gate59inter4), .b(gate59inter3), .O(gate59inter5));
  nor2  gate349(.a(gate59inter5), .b(gate59inter2), .O(gate59inter6));
  inv1  gate350(.a(N203), .O(gate59inter7));
  inv1  gate351(.a(N177), .O(gate59inter8));
  nand2 gate352(.a(gate59inter8), .b(gate59inter7), .O(gate59inter9));
  nand2 gate353(.a(s_27), .b(gate59inter3), .O(gate59inter10));
  nor2  gate354(.a(gate59inter10), .b(gate59inter9), .O(gate59inter11));
  nor2  gate355(.a(gate59inter11), .b(gate59inter6), .O(gate59inter12));
  nand2 gate356(.a(gate59inter12), .b(gate59inter1), .O(N247));
nand2 gate60( .a(N213), .b(N24), .O(N250) );
xor2 gate61( .a(N203), .b(N180), .O(N251) );
nand2 gate62( .a(N213), .b(N37), .O(N254) );
nand2 gate63( .a(N213), .b(N50), .O(N255) );
nand2 gate64( .a(N213), .b(N63), .O(N256) );

  xor2  gate455(.a(N76), .b(N213), .O(gate65inter0));
  nand2 gate456(.a(gate65inter0), .b(s_42), .O(gate65inter1));
  and2  gate457(.a(N76), .b(N213), .O(gate65inter2));
  inv1  gate458(.a(s_42), .O(gate65inter3));
  inv1  gate459(.a(s_43), .O(gate65inter4));
  nand2 gate460(.a(gate65inter4), .b(gate65inter3), .O(gate65inter5));
  nor2  gate461(.a(gate65inter5), .b(gate65inter2), .O(gate65inter6));
  inv1  gate462(.a(N213), .O(gate65inter7));
  inv1  gate463(.a(N76), .O(gate65inter8));
  nand2 gate464(.a(gate65inter8), .b(gate65inter7), .O(gate65inter9));
  nand2 gate465(.a(s_43), .b(gate65inter3), .O(gate65inter10));
  nor2  gate466(.a(gate65inter10), .b(gate65inter9), .O(gate65inter11));
  nor2  gate467(.a(gate65inter11), .b(gate65inter6), .O(gate65inter12));
  nand2 gate468(.a(gate65inter12), .b(gate65inter1), .O(N257));
nand2 gate66( .a(N213), .b(N89), .O(N258) );
nand2 gate67( .a(N213), .b(N102), .O(N259) );

  xor2  gate497(.a(N157), .b(N224), .O(gate68inter0));
  nand2 gate498(.a(gate68inter0), .b(s_48), .O(gate68inter1));
  and2  gate499(.a(N157), .b(N224), .O(gate68inter2));
  inv1  gate500(.a(s_48), .O(gate68inter3));
  inv1  gate501(.a(s_49), .O(gate68inter4));
  nand2 gate502(.a(gate68inter4), .b(gate68inter3), .O(gate68inter5));
  nor2  gate503(.a(gate68inter5), .b(gate68inter2), .O(gate68inter6));
  inv1  gate504(.a(N224), .O(gate68inter7));
  inv1  gate505(.a(N157), .O(gate68inter8));
  nand2 gate506(.a(gate68inter8), .b(gate68inter7), .O(gate68inter9));
  nand2 gate507(.a(s_49), .b(gate68inter3), .O(gate68inter10));
  nor2  gate508(.a(gate68inter10), .b(gate68inter9), .O(gate68inter11));
  nor2  gate509(.a(gate68inter11), .b(gate68inter6), .O(gate68inter12));
  nand2 gate510(.a(gate68inter12), .b(gate68inter1), .O(N260));
nand2 gate69( .a(N224), .b(N158), .O(N263) );

  xor2  gate245(.a(N183), .b(N227), .O(gate70inter0));
  nand2 gate246(.a(gate70inter0), .b(s_12), .O(gate70inter1));
  and2  gate247(.a(N183), .b(N227), .O(gate70inter2));
  inv1  gate248(.a(s_12), .O(gate70inter3));
  inv1  gate249(.a(s_13), .O(gate70inter4));
  nand2 gate250(.a(gate70inter4), .b(gate70inter3), .O(gate70inter5));
  nor2  gate251(.a(gate70inter5), .b(gate70inter2), .O(gate70inter6));
  inv1  gate252(.a(N227), .O(gate70inter7));
  inv1  gate253(.a(N183), .O(gate70inter8));
  nand2 gate254(.a(gate70inter8), .b(gate70inter7), .O(gate70inter9));
  nand2 gate255(.a(s_13), .b(gate70inter3), .O(gate70inter10));
  nor2  gate256(.a(gate70inter10), .b(gate70inter9), .O(gate70inter11));
  nor2  gate257(.a(gate70inter11), .b(gate70inter6), .O(gate70inter12));
  nand2 gate258(.a(gate70inter12), .b(gate70inter1), .O(N264));

  xor2  gate175(.a(N185), .b(N230), .O(gate71inter0));
  nand2 gate176(.a(gate71inter0), .b(s_2), .O(gate71inter1));
  and2  gate177(.a(N185), .b(N230), .O(gate71inter2));
  inv1  gate178(.a(s_2), .O(gate71inter3));
  inv1  gate179(.a(s_3), .O(gate71inter4));
  nand2 gate180(.a(gate71inter4), .b(gate71inter3), .O(gate71inter5));
  nor2  gate181(.a(gate71inter5), .b(gate71inter2), .O(gate71inter6));
  inv1  gate182(.a(N230), .O(gate71inter7));
  inv1  gate183(.a(N185), .O(gate71inter8));
  nand2 gate184(.a(gate71inter8), .b(gate71inter7), .O(gate71inter9));
  nand2 gate185(.a(s_3), .b(gate71inter3), .O(gate71inter10));
  nor2  gate186(.a(gate71inter10), .b(gate71inter9), .O(gate71inter11));
  nor2  gate187(.a(gate71inter11), .b(gate71inter6), .O(gate71inter12));
  nand2 gate188(.a(gate71inter12), .b(gate71inter1), .O(N267));

  xor2  gate231(.a(N187), .b(N233), .O(gate72inter0));
  nand2 gate232(.a(gate72inter0), .b(s_10), .O(gate72inter1));
  and2  gate233(.a(N187), .b(N233), .O(gate72inter2));
  inv1  gate234(.a(s_10), .O(gate72inter3));
  inv1  gate235(.a(s_11), .O(gate72inter4));
  nand2 gate236(.a(gate72inter4), .b(gate72inter3), .O(gate72inter5));
  nor2  gate237(.a(gate72inter5), .b(gate72inter2), .O(gate72inter6));
  inv1  gate238(.a(N233), .O(gate72inter7));
  inv1  gate239(.a(N187), .O(gate72inter8));
  nand2 gate240(.a(gate72inter8), .b(gate72inter7), .O(gate72inter9));
  nand2 gate241(.a(s_11), .b(gate72inter3), .O(gate72inter10));
  nor2  gate242(.a(gate72inter10), .b(gate72inter9), .O(gate72inter11));
  nor2  gate243(.a(gate72inter11), .b(gate72inter6), .O(gate72inter12));
  nand2 gate244(.a(gate72inter12), .b(gate72inter1), .O(N270));
nand2 gate73( .a(N236), .b(N189), .O(N273) );
nand2 gate74( .a(N239), .b(N191), .O(N276) );
nand2 gate75( .a(N243), .b(N193), .O(N279) );
nand2 gate76( .a(N247), .b(N195), .O(N282) );
nand2 gate77( .a(N251), .b(N197), .O(N285) );
nand2 gate78( .a(N227), .b(N184), .O(N288) );
nand2 gate79( .a(N230), .b(N186), .O(N289) );
nand2 gate80( .a(N233), .b(N188), .O(N290) );
nand2 gate81( .a(N236), .b(N190), .O(N291) );

  xor2  gate273(.a(N192), .b(N239), .O(gate82inter0));
  nand2 gate274(.a(gate82inter0), .b(s_16), .O(gate82inter1));
  and2  gate275(.a(N192), .b(N239), .O(gate82inter2));
  inv1  gate276(.a(s_16), .O(gate82inter3));
  inv1  gate277(.a(s_17), .O(gate82inter4));
  nand2 gate278(.a(gate82inter4), .b(gate82inter3), .O(gate82inter5));
  nor2  gate279(.a(gate82inter5), .b(gate82inter2), .O(gate82inter6));
  inv1  gate280(.a(N239), .O(gate82inter7));
  inv1  gate281(.a(N192), .O(gate82inter8));
  nand2 gate282(.a(gate82inter8), .b(gate82inter7), .O(gate82inter9));
  nand2 gate283(.a(s_17), .b(gate82inter3), .O(gate82inter10));
  nor2  gate284(.a(gate82inter10), .b(gate82inter9), .O(gate82inter11));
  nor2  gate285(.a(gate82inter11), .b(gate82inter6), .O(gate82inter12));
  nand2 gate286(.a(gate82inter12), .b(gate82inter1), .O(N292));
nand2 gate83( .a(N243), .b(N194), .O(N293) );
nand2 gate84( .a(N247), .b(N196), .O(N294) );

  xor2  gate329(.a(N198), .b(N251), .O(gate85inter0));
  nand2 gate330(.a(gate85inter0), .b(s_24), .O(gate85inter1));
  and2  gate331(.a(N198), .b(N251), .O(gate85inter2));
  inv1  gate332(.a(s_24), .O(gate85inter3));
  inv1  gate333(.a(s_25), .O(gate85inter4));
  nand2 gate334(.a(gate85inter4), .b(gate85inter3), .O(gate85inter5));
  nor2  gate335(.a(gate85inter5), .b(gate85inter2), .O(gate85inter6));
  inv1  gate336(.a(N251), .O(gate85inter7));
  inv1  gate337(.a(N198), .O(gate85inter8));
  nand2 gate338(.a(gate85inter8), .b(gate85inter7), .O(gate85inter9));
  nand2 gate339(.a(s_25), .b(gate85inter3), .O(gate85inter10));
  nor2  gate340(.a(gate85inter10), .b(gate85inter9), .O(gate85inter11));
  nor2  gate341(.a(gate85inter11), .b(gate85inter6), .O(gate85inter12));
  nand2 gate342(.a(gate85inter12), .b(gate85inter1), .O(N295));
and9 gate86( .a(N260), .b(N264), .c(N267), .d(N270), .e(N273), .f(N276), .g(N279), .h(N282), .i(N285), .O(N296) );
inv1 gate87( .a(N263), .O(N300) );
inv1 gate88( .a(N288), .O(N301) );
inv1 gate89( .a(N289), .O(N302) );
inv1 gate90( .a(N290), .O(N303) );
inv1 gate91( .a(N291), .O(N304) );
inv1 gate92( .a(N292), .O(N305) );
inv1 gate93( .a(N293), .O(N306) );
inv1 gate94( .a(N294), .O(N307) );
inv1 gate95( .a(N295), .O(N308) );
inv1 gate96( .a(N296), .O(N309) );
inv1 gate97( .a(N296), .O(N319) );
inv1 gate98( .a(N296), .O(N329) );
xor2 gate99( .a(N309), .b(N260), .O(N330) );
xor2 gate100( .a(N309), .b(N264), .O(N331) );

  xor2  gate357(.a(N267), .b(N309), .O(gate101inter0));
  nand2 gate358(.a(gate101inter0), .b(s_28), .O(gate101inter1));
  and2  gate359(.a(N267), .b(N309), .O(gate101inter2));
  inv1  gate360(.a(s_28), .O(gate101inter3));
  inv1  gate361(.a(s_29), .O(gate101inter4));
  nand2 gate362(.a(gate101inter4), .b(gate101inter3), .O(gate101inter5));
  nor2  gate363(.a(gate101inter5), .b(gate101inter2), .O(gate101inter6));
  inv1  gate364(.a(N309), .O(gate101inter7));
  inv1  gate365(.a(N267), .O(gate101inter8));
  nand2 gate366(.a(gate101inter8), .b(gate101inter7), .O(gate101inter9));
  nand2 gate367(.a(s_29), .b(gate101inter3), .O(gate101inter10));
  nor2  gate368(.a(gate101inter10), .b(gate101inter9), .O(gate101inter11));
  nor2  gate369(.a(gate101inter11), .b(gate101inter6), .O(gate101inter12));
  nand2 gate370(.a(gate101inter12), .b(gate101inter1), .O(N332));
xor2 gate102( .a(N309), .b(N270), .O(N333) );
nand2 gate103( .a(N8), .b(N319), .O(N334) );

  xor2  gate441(.a(N273), .b(N309), .O(gate104inter0));
  nand2 gate442(.a(gate104inter0), .b(s_40), .O(gate104inter1));
  and2  gate443(.a(N273), .b(N309), .O(gate104inter2));
  inv1  gate444(.a(s_40), .O(gate104inter3));
  inv1  gate445(.a(s_41), .O(gate104inter4));
  nand2 gate446(.a(gate104inter4), .b(gate104inter3), .O(gate104inter5));
  nor2  gate447(.a(gate104inter5), .b(gate104inter2), .O(gate104inter6));
  inv1  gate448(.a(N309), .O(gate104inter7));
  inv1  gate449(.a(N273), .O(gate104inter8));
  nand2 gate450(.a(gate104inter8), .b(gate104inter7), .O(gate104inter9));
  nand2 gate451(.a(s_41), .b(gate104inter3), .O(gate104inter10));
  nor2  gate452(.a(gate104inter10), .b(gate104inter9), .O(gate104inter11));
  nor2  gate453(.a(gate104inter11), .b(gate104inter6), .O(gate104inter12));
  nand2 gate454(.a(gate104inter12), .b(gate104inter1), .O(N335));
nand2 gate105( .a(N319), .b(N21), .O(N336) );
xor2 gate106( .a(N309), .b(N276), .O(N337) );
nand2 gate107( .a(N319), .b(N34), .O(N338) );

  xor2  gate189(.a(N279), .b(N309), .O(gate108inter0));
  nand2 gate190(.a(gate108inter0), .b(s_4), .O(gate108inter1));
  and2  gate191(.a(N279), .b(N309), .O(gate108inter2));
  inv1  gate192(.a(s_4), .O(gate108inter3));
  inv1  gate193(.a(s_5), .O(gate108inter4));
  nand2 gate194(.a(gate108inter4), .b(gate108inter3), .O(gate108inter5));
  nor2  gate195(.a(gate108inter5), .b(gate108inter2), .O(gate108inter6));
  inv1  gate196(.a(N309), .O(gate108inter7));
  inv1  gate197(.a(N279), .O(gate108inter8));
  nand2 gate198(.a(gate108inter8), .b(gate108inter7), .O(gate108inter9));
  nand2 gate199(.a(s_5), .b(gate108inter3), .O(gate108inter10));
  nor2  gate200(.a(gate108inter10), .b(gate108inter9), .O(gate108inter11));
  nor2  gate201(.a(gate108inter11), .b(gate108inter6), .O(gate108inter12));
  nand2 gate202(.a(gate108inter12), .b(gate108inter1), .O(N339));
nand2 gate109( .a(N319), .b(N47), .O(N340) );
xor2 gate110( .a(N309), .b(N282), .O(N341) );
nand2 gate111( .a(N319), .b(N60), .O(N342) );
xor2 gate112( .a(N309), .b(N285), .O(N343) );
nand2 gate113( .a(N319), .b(N73), .O(N344) );

  xor2  gate203(.a(N86), .b(N319), .O(gate114inter0));
  nand2 gate204(.a(gate114inter0), .b(s_6), .O(gate114inter1));
  and2  gate205(.a(N86), .b(N319), .O(gate114inter2));
  inv1  gate206(.a(s_6), .O(gate114inter3));
  inv1  gate207(.a(s_7), .O(gate114inter4));
  nand2 gate208(.a(gate114inter4), .b(gate114inter3), .O(gate114inter5));
  nor2  gate209(.a(gate114inter5), .b(gate114inter2), .O(gate114inter6));
  inv1  gate210(.a(N319), .O(gate114inter7));
  inv1  gate211(.a(N86), .O(gate114inter8));
  nand2 gate212(.a(gate114inter8), .b(gate114inter7), .O(gate114inter9));
  nand2 gate213(.a(s_7), .b(gate114inter3), .O(gate114inter10));
  nor2  gate214(.a(gate114inter10), .b(gate114inter9), .O(gate114inter11));
  nor2  gate215(.a(gate114inter11), .b(gate114inter6), .O(gate114inter12));
  nand2 gate216(.a(gate114inter12), .b(gate114inter1), .O(N345));
nand2 gate115( .a(N319), .b(N99), .O(N346) );

  xor2  gate315(.a(N112), .b(N319), .O(gate116inter0));
  nand2 gate316(.a(gate116inter0), .b(s_22), .O(gate116inter1));
  and2  gate317(.a(N112), .b(N319), .O(gate116inter2));
  inv1  gate318(.a(s_22), .O(gate116inter3));
  inv1  gate319(.a(s_23), .O(gate116inter4));
  nand2 gate320(.a(gate116inter4), .b(gate116inter3), .O(gate116inter5));
  nor2  gate321(.a(gate116inter5), .b(gate116inter2), .O(gate116inter6));
  inv1  gate322(.a(N319), .O(gate116inter7));
  inv1  gate323(.a(N112), .O(gate116inter8));
  nand2 gate324(.a(gate116inter8), .b(gate116inter7), .O(gate116inter9));
  nand2 gate325(.a(s_23), .b(gate116inter3), .O(gate116inter10));
  nor2  gate326(.a(gate116inter10), .b(gate116inter9), .O(gate116inter11));
  nor2  gate327(.a(gate116inter11), .b(gate116inter6), .O(gate116inter12));
  nand2 gate328(.a(gate116inter12), .b(gate116inter1), .O(N347));
nand2 gate117( .a(N330), .b(N300), .O(N348) );
nand2 gate118( .a(N331), .b(N301), .O(N349) );
nand2 gate119( .a(N332), .b(N302), .O(N350) );
nand2 gate120( .a(N333), .b(N303), .O(N351) );
nand2 gate121( .a(N335), .b(N304), .O(N352) );
nand2 gate122( .a(N337), .b(N305), .O(N353) );
nand2 gate123( .a(N339), .b(N306), .O(N354) );
nand2 gate124( .a(N341), .b(N307), .O(N355) );
nand2 gate125( .a(N343), .b(N308), .O(N356) );
and9 gate126( .a(N348), .b(N349), .c(N350), .d(N351), .e(N352), .f(N353), .g(N354), .h(N355), .i(N356), .O(N357) );
inv1 gate127( .a(N357), .O(N360) );
inv1 gate128( .a(N357), .O(N370) );
nand2 gate129( .a(N14), .b(N360), .O(N371) );

  xor2  gate217(.a(N27), .b(N360), .O(gate130inter0));
  nand2 gate218(.a(gate130inter0), .b(s_8), .O(gate130inter1));
  and2  gate219(.a(N27), .b(N360), .O(gate130inter2));
  inv1  gate220(.a(s_8), .O(gate130inter3));
  inv1  gate221(.a(s_9), .O(gate130inter4));
  nand2 gate222(.a(gate130inter4), .b(gate130inter3), .O(gate130inter5));
  nor2  gate223(.a(gate130inter5), .b(gate130inter2), .O(gate130inter6));
  inv1  gate224(.a(N360), .O(gate130inter7));
  inv1  gate225(.a(N27), .O(gate130inter8));
  nand2 gate226(.a(gate130inter8), .b(gate130inter7), .O(gate130inter9));
  nand2 gate227(.a(s_9), .b(gate130inter3), .O(gate130inter10));
  nor2  gate228(.a(gate130inter10), .b(gate130inter9), .O(gate130inter11));
  nor2  gate229(.a(gate130inter11), .b(gate130inter6), .O(gate130inter12));
  nand2 gate230(.a(gate130inter12), .b(gate130inter1), .O(N372));

  xor2  gate385(.a(N40), .b(N360), .O(gate131inter0));
  nand2 gate386(.a(gate131inter0), .b(s_32), .O(gate131inter1));
  and2  gate387(.a(N40), .b(N360), .O(gate131inter2));
  inv1  gate388(.a(s_32), .O(gate131inter3));
  inv1  gate389(.a(s_33), .O(gate131inter4));
  nand2 gate390(.a(gate131inter4), .b(gate131inter3), .O(gate131inter5));
  nor2  gate391(.a(gate131inter5), .b(gate131inter2), .O(gate131inter6));
  inv1  gate392(.a(N360), .O(gate131inter7));
  inv1  gate393(.a(N40), .O(gate131inter8));
  nand2 gate394(.a(gate131inter8), .b(gate131inter7), .O(gate131inter9));
  nand2 gate395(.a(s_33), .b(gate131inter3), .O(gate131inter10));
  nor2  gate396(.a(gate131inter10), .b(gate131inter9), .O(gate131inter11));
  nor2  gate397(.a(gate131inter11), .b(gate131inter6), .O(gate131inter12));
  nand2 gate398(.a(gate131inter12), .b(gate131inter1), .O(N373));

  xor2  gate399(.a(N53), .b(N360), .O(gate132inter0));
  nand2 gate400(.a(gate132inter0), .b(s_34), .O(gate132inter1));
  and2  gate401(.a(N53), .b(N360), .O(gate132inter2));
  inv1  gate402(.a(s_34), .O(gate132inter3));
  inv1  gate403(.a(s_35), .O(gate132inter4));
  nand2 gate404(.a(gate132inter4), .b(gate132inter3), .O(gate132inter5));
  nor2  gate405(.a(gate132inter5), .b(gate132inter2), .O(gate132inter6));
  inv1  gate406(.a(N360), .O(gate132inter7));
  inv1  gate407(.a(N53), .O(gate132inter8));
  nand2 gate408(.a(gate132inter8), .b(gate132inter7), .O(gate132inter9));
  nand2 gate409(.a(s_35), .b(gate132inter3), .O(gate132inter10));
  nor2  gate410(.a(gate132inter10), .b(gate132inter9), .O(gate132inter11));
  nor2  gate411(.a(gate132inter11), .b(gate132inter6), .O(gate132inter12));
  nand2 gate412(.a(gate132inter12), .b(gate132inter1), .O(N374));
nand2 gate133( .a(N360), .b(N66), .O(N375) );
nand2 gate134( .a(N360), .b(N79), .O(N376) );

  xor2  gate413(.a(N92), .b(N360), .O(gate135inter0));
  nand2 gate414(.a(gate135inter0), .b(s_36), .O(gate135inter1));
  and2  gate415(.a(N92), .b(N360), .O(gate135inter2));
  inv1  gate416(.a(s_36), .O(gate135inter3));
  inv1  gate417(.a(s_37), .O(gate135inter4));
  nand2 gate418(.a(gate135inter4), .b(gate135inter3), .O(gate135inter5));
  nor2  gate419(.a(gate135inter5), .b(gate135inter2), .O(gate135inter6));
  inv1  gate420(.a(N360), .O(gate135inter7));
  inv1  gate421(.a(N92), .O(gate135inter8));
  nand2 gate422(.a(gate135inter8), .b(gate135inter7), .O(gate135inter9));
  nand2 gate423(.a(s_37), .b(gate135inter3), .O(gate135inter10));
  nor2  gate424(.a(gate135inter10), .b(gate135inter9), .O(gate135inter11));
  nor2  gate425(.a(gate135inter11), .b(gate135inter6), .O(gate135inter12));
  nand2 gate426(.a(gate135inter12), .b(gate135inter1), .O(N377));
nand2 gate136( .a(N360), .b(N105), .O(N378) );
nand2 gate137( .a(N360), .b(N115), .O(N379) );
nand4 gate138( .a(N4), .b(N242), .c(N334), .d(N371), .O(N380) );
nand4 gate139( .a(N246), .b(N336), .c(N372), .d(N17), .O(N381) );
nand4 gate140( .a(N250), .b(N338), .c(N373), .d(N30), .O(N386) );
nand4 gate141( .a(N254), .b(N340), .c(N374), .d(N43), .O(N393) );
nand4 gate142( .a(N255), .b(N342), .c(N375), .d(N56), .O(N399) );
nand4 gate143( .a(N256), .b(N344), .c(N376), .d(N69), .O(N404) );
nand4 gate144( .a(N257), .b(N345), .c(N377), .d(N82), .O(N407) );
nand4 gate145( .a(N258), .b(N346), .c(N378), .d(N95), .O(N411) );
nand4 gate146( .a(N259), .b(N347), .c(N379), .d(N108), .O(N414) );
inv1 gate147( .a(N380), .O(N415) );
and8 gate148( .a(N381), .b(N386), .c(N393), .d(N399), .e(N404), .f(N407), .g(N411), .h(N414), .O(N416) );
inv1 gate149( .a(N393), .O(N417) );
inv1 gate150( .a(N404), .O(N418) );
inv1 gate151( .a(N407), .O(N419) );
inv1 gate152( .a(N411), .O(N420) );
nor2 gate153( .a(N415), .b(N416), .O(N421) );

  xor2  gate483(.a(N417), .b(N386), .O(gate154inter0));
  nand2 gate484(.a(gate154inter0), .b(s_46), .O(gate154inter1));
  and2  gate485(.a(N417), .b(N386), .O(gate154inter2));
  inv1  gate486(.a(s_46), .O(gate154inter3));
  inv1  gate487(.a(s_47), .O(gate154inter4));
  nand2 gate488(.a(gate154inter4), .b(gate154inter3), .O(gate154inter5));
  nor2  gate489(.a(gate154inter5), .b(gate154inter2), .O(gate154inter6));
  inv1  gate490(.a(N386), .O(gate154inter7));
  inv1  gate491(.a(N417), .O(gate154inter8));
  nand2 gate492(.a(gate154inter8), .b(gate154inter7), .O(gate154inter9));
  nand2 gate493(.a(s_47), .b(gate154inter3), .O(gate154inter10));
  nor2  gate494(.a(gate154inter10), .b(gate154inter9), .O(gate154inter11));
  nor2  gate495(.a(gate154inter11), .b(gate154inter6), .O(gate154inter12));
  nand2 gate496(.a(gate154inter12), .b(gate154inter1), .O(N422));
nand4 gate155( .a(N386), .b(N393), .c(N418), .d(N399), .O(N425) );
nand3 gate156( .a(N399), .b(N393), .c(N419), .O(N428) );
nand4 gate157( .a(N386), .b(N393), .c(N407), .d(N420), .O(N429) );
nand4 gate158( .a(N381), .b(N386), .c(N422), .d(N399), .O(N430) );
nand4 gate159( .a(N381), .b(N386), .c(N425), .d(N428), .O(N431) );
nand4 gate160( .a(N381), .b(N422), .c(N425), .d(N429), .O(N432) );

endmodule