module c432 (N1,N4,N8,N11,N14,N17,N21,N24,N27,N30,
             N34,N37,N40,N43,N47,N50,N53,N56,N60,N63,
             N66,N69,N73,N76,N79,N82,N86,N89,N92,N95,
             N99,N102,N105,N108,N112,N115,N223,N329,N370,N421,
             N430,N431,N432);

input N1,N4,N8,N11,N14,N17,N21,N24,N27,N30,
      N34,N37,N40,N43,N47,N50,N53,N56,N60,N63,
      N66,N69,N73,N76,N79,N82,N86,N89,N92,N95,
      N99,N102,N105,N108,N112,N115;//RE__PI;

input s_0,s_1;//RE__ALLOW(00,01,10,11);
input s_2,s_3;//RE__ALLOW(00,01,10,11);
input s_4,s_5;//RE__ALLOW(00,01,10,11);
input s_6,s_7;//RE__ALLOW(00,01,10,11);
input s_8,s_9;//RE__ALLOW(00,01,10,11);
input s_10,s_11;//RE__ALLOW(00,01,10,11);
input s_12,s_13;//RE__ALLOW(00,01,10,11);
input s_14,s_15;//RE__ALLOW(00,01,10,11);
input s_16,s_17;//RE__ALLOW(00,01,10,11);
input s_18,s_19;//RE__ALLOW(00,01,10,11);
input s_20,s_21;//RE__ALLOW(00,01,10,11);
input s_22,s_23;//RE__ALLOW(00,01,10,11);
input s_24,s_25;//RE__ALLOW(00,01,10,11);
input s_26,s_27;//RE__ALLOW(00,01,10,11);
input s_28,s_29;//RE__ALLOW(00,01,10,11);
input s_30,s_31;//RE__ALLOW(00,01,10,11);
input s_32,s_33;//RE__ALLOW(00,01,10,11);
input s_34,s_35;//RE__ALLOW(00,01,10,11);
input s_36,s_37;//RE__ALLOW(00,01,10,11);
input s_38,s_39;//RE__ALLOW(00,01,10,11);
input s_40,s_41;//RE__ALLOW(00,01,10,11);
input s_42,s_43;//RE__ALLOW(00,01,10,11);
input s_44,s_45;//RE__ALLOW(00,01,10,11);
input s_46,s_47;//RE__ALLOW(00,01,10,11);
input s_48,s_49;//RE__ALLOW(00,01,10,11);
input s_50,s_51;//RE__ALLOW(00,01,10,11);
output N223,N329,N370,N421,N430,N431,N432;

wire N118,N119,N122,N123,N126,N127,N130,N131,N134,N135,
     N138,N139,N142,N143,N146,N147,N150,N151,N154,N157,
     N158,N159,N162,N165,N168,N171,N174,N177,N180,N183,
     N184,N185,N186,N187,N188,N189,N190,N191,N192,N193,
     N194,N195,N196,N197,N198,N199,N203,N213,N224,N227,
     N230,N233,N236,N239,N242,N243,N246,N247,N250,N251,
     N254,N255,N256,N257,N258,N259,N260,N263,N264,N267,
     N270,N273,N276,N279,N282,N285,N288,N289,N290,N291,
     N292,N293,N294,N295,N296,N300,N301,N302,N303,N304,
     N305,N306,N307,N308,N309,N319,N330,N331,N332,N333,
     N334,N335,N336,N337,N338,N339,N340,N341,N342,N343,
     N344,N345,N346,N347,N348,N349,N350,N351,N352,N353,
     N354,N355,N356,N357,N360,N371,N372,N373,N374,N375,
     N376,N377,N378,N379,N380,N381,N386,N393,N399,N404,
     N407,N411,N414,N415,N416,N417,N418,N419,N420,N422,
     N425,N428,N429, gate57inter0, gate57inter1, gate57inter2, gate57inter3, gate57inter4, gate57inter5, gate57inter6, gate57inter7, gate57inter8, gate57inter9, gate57inter10, gate57inter11, gate57inter12, gate58inter0, gate58inter1, gate58inter2, gate58inter3, gate58inter4, gate58inter5, gate58inter6, gate58inter7, gate58inter8, gate58inter9, gate58inter10, gate58inter11, gate58inter12, gate40inter0, gate40inter1, gate40inter2, gate40inter3, gate40inter4, gate40inter5, gate40inter6, gate40inter7, gate40inter8, gate40inter9, gate40inter10, gate40inter11, gate40inter12, gate154inter0, gate154inter1, gate154inter2, gate154inter3, gate154inter4, gate154inter5, gate154inter6, gate154inter7, gate154inter8, gate154inter9, gate154inter10, gate154inter11, gate154inter12, gate118inter0, gate118inter1, gate118inter2, gate118inter3, gate118inter4, gate118inter5, gate118inter6, gate118inter7, gate118inter8, gate118inter9, gate118inter10, gate118inter11, gate118inter12, gate123inter0, gate123inter1, gate123inter2, gate123inter3, gate123inter4, gate123inter5, gate123inter6, gate123inter7, gate123inter8, gate123inter9, gate123inter10, gate123inter11, gate123inter12, gate80inter0, gate80inter1, gate80inter2, gate80inter3, gate80inter4, gate80inter5, gate80inter6, gate80inter7, gate80inter8, gate80inter9, gate80inter10, gate80inter11, gate80inter12, gate32inter0, gate32inter1, gate32inter2, gate32inter3, gate32inter4, gate32inter5, gate32inter6, gate32inter7, gate32inter8, gate32inter9, gate32inter10, gate32inter11, gate32inter12, gate70inter0, gate70inter1, gate70inter2, gate70inter3, gate70inter4, gate70inter5, gate70inter6, gate70inter7, gate70inter8, gate70inter9, gate70inter10, gate70inter11, gate70inter12, gate20inter0, gate20inter1, gate20inter2, gate20inter3, gate20inter4, gate20inter5, gate20inter6, gate20inter7, gate20inter8, gate20inter9, gate20inter10, gate20inter11, gate20inter12, gate136inter0, gate136inter1, gate136inter2, gate136inter3, gate136inter4, gate136inter5, gate136inter6, gate136inter7, gate136inter8, gate136inter9, gate136inter10, gate136inter11, gate136inter12, gate113inter0, gate113inter1, gate113inter2, gate113inter3, gate113inter4, gate113inter5, gate113inter6, gate113inter7, gate113inter8, gate113inter9, gate113inter10, gate113inter11, gate113inter12, gate72inter0, gate72inter1, gate72inter2, gate72inter3, gate72inter4, gate72inter5, gate72inter6, gate72inter7, gate72inter8, gate72inter9, gate72inter10, gate72inter11, gate72inter12, gate77inter0, gate77inter1, gate77inter2, gate77inter3, gate77inter4, gate77inter5, gate77inter6, gate77inter7, gate77inter8, gate77inter9, gate77inter10, gate77inter11, gate77inter12, gate54inter0, gate54inter1, gate54inter2, gate54inter3, gate54inter4, gate54inter5, gate54inter6, gate54inter7, gate54inter8, gate54inter9, gate54inter10, gate54inter11, gate54inter12, gate43inter0, gate43inter1, gate43inter2, gate43inter3, gate43inter4, gate43inter5, gate43inter6, gate43inter7, gate43inter8, gate43inter9, gate43inter10, gate43inter11, gate43inter12, gate119inter0, gate119inter1, gate119inter2, gate119inter3, gate119inter4, gate119inter5, gate119inter6, gate119inter7, gate119inter8, gate119inter9, gate119inter10, gate119inter11, gate119inter12, gate24inter0, gate24inter1, gate24inter2, gate24inter3, gate24inter4, gate24inter5, gate24inter6, gate24inter7, gate24inter8, gate24inter9, gate24inter10, gate24inter11, gate24inter12, gate37inter0, gate37inter1, gate37inter2, gate37inter3, gate37inter4, gate37inter5, gate37inter6, gate37inter7, gate37inter8, gate37inter9, gate37inter10, gate37inter11, gate37inter12, gate129inter0, gate129inter1, gate129inter2, gate129inter3, gate129inter4, gate129inter5, gate129inter6, gate129inter7, gate129inter8, gate129inter9, gate129inter10, gate129inter11, gate129inter12, gate85inter0, gate85inter1, gate85inter2, gate85inter3, gate85inter4, gate85inter5, gate85inter6, gate85inter7, gate85inter8, gate85inter9, gate85inter10, gate85inter11, gate85inter12, gate75inter0, gate75inter1, gate75inter2, gate75inter3, gate75inter4, gate75inter5, gate75inter6, gate75inter7, gate75inter8, gate75inter9, gate75inter10, gate75inter11, gate75inter12, gate52inter0, gate52inter1, gate52inter2, gate52inter3, gate52inter4, gate52inter5, gate52inter6, gate52inter7, gate52inter8, gate52inter9, gate52inter10, gate52inter11, gate52inter12, gate111inter0, gate111inter1, gate111inter2, gate111inter3, gate111inter4, gate111inter5, gate111inter6, gate111inter7, gate111inter8, gate111inter9, gate111inter10, gate111inter11, gate111inter12, gate22inter0, gate22inter1, gate22inter2, gate22inter3, gate22inter4, gate22inter5, gate22inter6, gate22inter7, gate22inter8, gate22inter9, gate22inter10, gate22inter11, gate22inter12, gate62inter0, gate62inter1, gate62inter2, gate62inter3, gate62inter4, gate62inter5, gate62inter6, gate62inter7, gate62inter8, gate62inter9, gate62inter10, gate62inter11, gate62inter12;



inv1 gate1( .a(N1), .O(N118) );
inv1 gate2( .a(N4), .O(N119) );
inv1 gate3( .a(N11), .O(N122) );
inv1 gate4( .a(N17), .O(N123) );
inv1 gate5( .a(N24), .O(N126) );
inv1 gate6( .a(N30), .O(N127) );
inv1 gate7( .a(N37), .O(N130) );
inv1 gate8( .a(N43), .O(N131) );
inv1 gate9( .a(N50), .O(N134) );
inv1 gate10( .a(N56), .O(N135) );
inv1 gate11( .a(N63), .O(N138) );
inv1 gate12( .a(N69), .O(N139) );
inv1 gate13( .a(N76), .O(N142) );
inv1 gate14( .a(N82), .O(N143) );
inv1 gate15( .a(N89), .O(N146) );
inv1 gate16( .a(N95), .O(N147) );
inv1 gate17( .a(N102), .O(N150) );
inv1 gate18( .a(N108), .O(N151) );
nand2 gate19( .a(N118), .b(N4), .O(N154) );

  xor2  gate287(.a(N119), .b(N8), .O(gate20inter0));
  nand2 gate288(.a(gate20inter0), .b(s_18), .O(gate20inter1));
  and2  gate289(.a(N119), .b(N8), .O(gate20inter2));
  inv1  gate290(.a(s_18), .O(gate20inter3));
  inv1  gate291(.a(s_19), .O(gate20inter4));
  nand2 gate292(.a(gate20inter4), .b(gate20inter3), .O(gate20inter5));
  nor2  gate293(.a(gate20inter5), .b(gate20inter2), .O(gate20inter6));
  inv1  gate294(.a(N8), .O(gate20inter7));
  inv1  gate295(.a(N119), .O(gate20inter8));
  nand2 gate296(.a(gate20inter8), .b(gate20inter7), .O(gate20inter9));
  nand2 gate297(.a(s_19), .b(gate20inter3), .O(gate20inter10));
  nor2  gate298(.a(gate20inter10), .b(gate20inter9), .O(gate20inter11));
  nor2  gate299(.a(gate20inter11), .b(gate20inter6), .O(gate20inter12));
  nand2 gate300(.a(gate20inter12), .b(gate20inter1), .O(N157));
nor2 gate21( .a(N14), .b(N119), .O(N158) );

  xor2  gate497(.a(N17), .b(N122), .O(gate22inter0));
  nand2 gate498(.a(gate22inter0), .b(s_48), .O(gate22inter1));
  and2  gate499(.a(N17), .b(N122), .O(gate22inter2));
  inv1  gate500(.a(s_48), .O(gate22inter3));
  inv1  gate501(.a(s_49), .O(gate22inter4));
  nand2 gate502(.a(gate22inter4), .b(gate22inter3), .O(gate22inter5));
  nor2  gate503(.a(gate22inter5), .b(gate22inter2), .O(gate22inter6));
  inv1  gate504(.a(N122), .O(gate22inter7));
  inv1  gate505(.a(N17), .O(gate22inter8));
  nand2 gate506(.a(gate22inter8), .b(gate22inter7), .O(gate22inter9));
  nand2 gate507(.a(s_49), .b(gate22inter3), .O(gate22inter10));
  nor2  gate508(.a(gate22inter10), .b(gate22inter9), .O(gate22inter11));
  nor2  gate509(.a(gate22inter11), .b(gate22inter6), .O(gate22inter12));
  nand2 gate510(.a(gate22inter12), .b(gate22inter1), .O(N159));
nand2 gate23( .a(N126), .b(N30), .O(N162) );

  xor2  gate399(.a(N43), .b(N130), .O(gate24inter0));
  nand2 gate400(.a(gate24inter0), .b(s_34), .O(gate24inter1));
  and2  gate401(.a(N43), .b(N130), .O(gate24inter2));
  inv1  gate402(.a(s_34), .O(gate24inter3));
  inv1  gate403(.a(s_35), .O(gate24inter4));
  nand2 gate404(.a(gate24inter4), .b(gate24inter3), .O(gate24inter5));
  nor2  gate405(.a(gate24inter5), .b(gate24inter2), .O(gate24inter6));
  inv1  gate406(.a(N130), .O(gate24inter7));
  inv1  gate407(.a(N43), .O(gate24inter8));
  nand2 gate408(.a(gate24inter8), .b(gate24inter7), .O(gate24inter9));
  nand2 gate409(.a(s_35), .b(gate24inter3), .O(gate24inter10));
  nor2  gate410(.a(gate24inter10), .b(gate24inter9), .O(gate24inter11));
  nor2  gate411(.a(gate24inter11), .b(gate24inter6), .O(gate24inter12));
  nand2 gate412(.a(gate24inter12), .b(gate24inter1), .O(N165));
nand2 gate25( .a(N134), .b(N56), .O(N168) );
nand2 gate26( .a(N138), .b(N69), .O(N171) );
nand2 gate27( .a(N142), .b(N82), .O(N174) );
nand2 gate28( .a(N146), .b(N95), .O(N177) );
nand2 gate29( .a(N150), .b(N108), .O(N180) );
nor2 gate30( .a(N21), .b(N123), .O(N183) );
nor2 gate31( .a(N27), .b(N123), .O(N184) );

  xor2  gate259(.a(N127), .b(N34), .O(gate32inter0));
  nand2 gate260(.a(gate32inter0), .b(s_14), .O(gate32inter1));
  and2  gate261(.a(N127), .b(N34), .O(gate32inter2));
  inv1  gate262(.a(s_14), .O(gate32inter3));
  inv1  gate263(.a(s_15), .O(gate32inter4));
  nand2 gate264(.a(gate32inter4), .b(gate32inter3), .O(gate32inter5));
  nor2  gate265(.a(gate32inter5), .b(gate32inter2), .O(gate32inter6));
  inv1  gate266(.a(N34), .O(gate32inter7));
  inv1  gate267(.a(N127), .O(gate32inter8));
  nand2 gate268(.a(gate32inter8), .b(gate32inter7), .O(gate32inter9));
  nand2 gate269(.a(s_15), .b(gate32inter3), .O(gate32inter10));
  nor2  gate270(.a(gate32inter10), .b(gate32inter9), .O(gate32inter11));
  nor2  gate271(.a(gate32inter11), .b(gate32inter6), .O(gate32inter12));
  nand2 gate272(.a(gate32inter12), .b(gate32inter1), .O(N185));
nor2 gate33( .a(N40), .b(N127), .O(N186) );
nor2 gate34( .a(N47), .b(N131), .O(N187) );
nor2 gate35( .a(N53), .b(N131), .O(N188) );
nor2 gate36( .a(N60), .b(N135), .O(N189) );

  xor2  gate413(.a(N135), .b(N66), .O(gate37inter0));
  nand2 gate414(.a(gate37inter0), .b(s_36), .O(gate37inter1));
  and2  gate415(.a(N135), .b(N66), .O(gate37inter2));
  inv1  gate416(.a(s_36), .O(gate37inter3));
  inv1  gate417(.a(s_37), .O(gate37inter4));
  nand2 gate418(.a(gate37inter4), .b(gate37inter3), .O(gate37inter5));
  nor2  gate419(.a(gate37inter5), .b(gate37inter2), .O(gate37inter6));
  inv1  gate420(.a(N66), .O(gate37inter7));
  inv1  gate421(.a(N135), .O(gate37inter8));
  nand2 gate422(.a(gate37inter8), .b(gate37inter7), .O(gate37inter9));
  nand2 gate423(.a(s_37), .b(gate37inter3), .O(gate37inter10));
  nor2  gate424(.a(gate37inter10), .b(gate37inter9), .O(gate37inter11));
  nor2  gate425(.a(gate37inter11), .b(gate37inter6), .O(gate37inter12));
  nand2 gate426(.a(gate37inter12), .b(gate37inter1), .O(N190));
nor2 gate38( .a(N73), .b(N139), .O(N191) );
nor2 gate39( .a(N79), .b(N139), .O(N192) );

  xor2  gate189(.a(N143), .b(N86), .O(gate40inter0));
  nand2 gate190(.a(gate40inter0), .b(s_4), .O(gate40inter1));
  and2  gate191(.a(N143), .b(N86), .O(gate40inter2));
  inv1  gate192(.a(s_4), .O(gate40inter3));
  inv1  gate193(.a(s_5), .O(gate40inter4));
  nand2 gate194(.a(gate40inter4), .b(gate40inter3), .O(gate40inter5));
  nor2  gate195(.a(gate40inter5), .b(gate40inter2), .O(gate40inter6));
  inv1  gate196(.a(N86), .O(gate40inter7));
  inv1  gate197(.a(N143), .O(gate40inter8));
  nand2 gate198(.a(gate40inter8), .b(gate40inter7), .O(gate40inter9));
  nand2 gate199(.a(s_5), .b(gate40inter3), .O(gate40inter10));
  nor2  gate200(.a(gate40inter10), .b(gate40inter9), .O(gate40inter11));
  nor2  gate201(.a(gate40inter11), .b(gate40inter6), .O(gate40inter12));
  nand2 gate202(.a(gate40inter12), .b(gate40inter1), .O(N193));
nor2 gate41( .a(N92), .b(N143), .O(N194) );
nor2 gate42( .a(N99), .b(N147), .O(N195) );

  xor2  gate371(.a(N147), .b(N105), .O(gate43inter0));
  nand2 gate372(.a(gate43inter0), .b(s_30), .O(gate43inter1));
  and2  gate373(.a(N147), .b(N105), .O(gate43inter2));
  inv1  gate374(.a(s_30), .O(gate43inter3));
  inv1  gate375(.a(s_31), .O(gate43inter4));
  nand2 gate376(.a(gate43inter4), .b(gate43inter3), .O(gate43inter5));
  nor2  gate377(.a(gate43inter5), .b(gate43inter2), .O(gate43inter6));
  inv1  gate378(.a(N105), .O(gate43inter7));
  inv1  gate379(.a(N147), .O(gate43inter8));
  nand2 gate380(.a(gate43inter8), .b(gate43inter7), .O(gate43inter9));
  nand2 gate381(.a(s_31), .b(gate43inter3), .O(gate43inter10));
  nor2  gate382(.a(gate43inter10), .b(gate43inter9), .O(gate43inter11));
  nor2  gate383(.a(gate43inter11), .b(gate43inter6), .O(gate43inter12));
  nand2 gate384(.a(gate43inter12), .b(gate43inter1), .O(N196));
nor2 gate44( .a(N112), .b(N151), .O(N197) );
nor2 gate45( .a(N115), .b(N151), .O(N198) );
and9 gate46( .a(N154), .b(N159), .c(N162), .d(N165), .e(N168), .f(N171), .g(N174), .h(N177), .i(N180), .O(N199) );
inv1 gate47( .a(N199), .O(N203) );
inv1 gate48( .a(N199), .O(N213) );
inv1 gate49( .a(N199), .O(N223) );
xor2 gate50( .a(N203), .b(N154), .O(N224) );
xor2 gate51( .a(N203), .b(N159), .O(N227) );

  xor2  gate469(.a(N162), .b(N203), .O(gate52inter0));
  nand2 gate470(.a(gate52inter0), .b(s_44), .O(gate52inter1));
  and2  gate471(.a(N162), .b(N203), .O(gate52inter2));
  inv1  gate472(.a(s_44), .O(gate52inter3));
  inv1  gate473(.a(s_45), .O(gate52inter4));
  nand2 gate474(.a(gate52inter4), .b(gate52inter3), .O(gate52inter5));
  nor2  gate475(.a(gate52inter5), .b(gate52inter2), .O(gate52inter6));
  inv1  gate476(.a(N203), .O(gate52inter7));
  inv1  gate477(.a(N162), .O(gate52inter8));
  nand2 gate478(.a(gate52inter8), .b(gate52inter7), .O(gate52inter9));
  nand2 gate479(.a(s_45), .b(gate52inter3), .O(gate52inter10));
  nor2  gate480(.a(gate52inter10), .b(gate52inter9), .O(gate52inter11));
  nor2  gate481(.a(gate52inter11), .b(gate52inter6), .O(gate52inter12));
  nand2 gate482(.a(gate52inter12), .b(gate52inter1), .O(N230));
xor2 gate53( .a(N203), .b(N165), .O(N233) );

  xor2  gate357(.a(N168), .b(N203), .O(gate54inter0));
  nand2 gate358(.a(gate54inter0), .b(s_28), .O(gate54inter1));
  and2  gate359(.a(N168), .b(N203), .O(gate54inter2));
  inv1  gate360(.a(s_28), .O(gate54inter3));
  inv1  gate361(.a(s_29), .O(gate54inter4));
  nand2 gate362(.a(gate54inter4), .b(gate54inter3), .O(gate54inter5));
  nor2  gate363(.a(gate54inter5), .b(gate54inter2), .O(gate54inter6));
  inv1  gate364(.a(N203), .O(gate54inter7));
  inv1  gate365(.a(N168), .O(gate54inter8));
  nand2 gate366(.a(gate54inter8), .b(gate54inter7), .O(gate54inter9));
  nand2 gate367(.a(s_29), .b(gate54inter3), .O(gate54inter10));
  nor2  gate368(.a(gate54inter10), .b(gate54inter9), .O(gate54inter11));
  nor2  gate369(.a(gate54inter11), .b(gate54inter6), .O(gate54inter12));
  nand2 gate370(.a(gate54inter12), .b(gate54inter1), .O(N236));
xor2 gate55( .a(N203), .b(N171), .O(N239) );
nand2 gate56( .a(N1), .b(N213), .O(N242) );

  xor2  gate161(.a(N174), .b(N203), .O(gate57inter0));
  nand2 gate162(.a(gate57inter0), .b(s_0), .O(gate57inter1));
  and2  gate163(.a(N174), .b(N203), .O(gate57inter2));
  inv1  gate164(.a(s_0), .O(gate57inter3));
  inv1  gate165(.a(s_1), .O(gate57inter4));
  nand2 gate166(.a(gate57inter4), .b(gate57inter3), .O(gate57inter5));
  nor2  gate167(.a(gate57inter5), .b(gate57inter2), .O(gate57inter6));
  inv1  gate168(.a(N203), .O(gate57inter7));
  inv1  gate169(.a(N174), .O(gate57inter8));
  nand2 gate170(.a(gate57inter8), .b(gate57inter7), .O(gate57inter9));
  nand2 gate171(.a(s_1), .b(gate57inter3), .O(gate57inter10));
  nor2  gate172(.a(gate57inter10), .b(gate57inter9), .O(gate57inter11));
  nor2  gate173(.a(gate57inter11), .b(gate57inter6), .O(gate57inter12));
  nand2 gate174(.a(gate57inter12), .b(gate57inter1), .O(N243));

  xor2  gate175(.a(N11), .b(N213), .O(gate58inter0));
  nand2 gate176(.a(gate58inter0), .b(s_2), .O(gate58inter1));
  and2  gate177(.a(N11), .b(N213), .O(gate58inter2));
  inv1  gate178(.a(s_2), .O(gate58inter3));
  inv1  gate179(.a(s_3), .O(gate58inter4));
  nand2 gate180(.a(gate58inter4), .b(gate58inter3), .O(gate58inter5));
  nor2  gate181(.a(gate58inter5), .b(gate58inter2), .O(gate58inter6));
  inv1  gate182(.a(N213), .O(gate58inter7));
  inv1  gate183(.a(N11), .O(gate58inter8));
  nand2 gate184(.a(gate58inter8), .b(gate58inter7), .O(gate58inter9));
  nand2 gate185(.a(s_3), .b(gate58inter3), .O(gate58inter10));
  nor2  gate186(.a(gate58inter10), .b(gate58inter9), .O(gate58inter11));
  nor2  gate187(.a(gate58inter11), .b(gate58inter6), .O(gate58inter12));
  nand2 gate188(.a(gate58inter12), .b(gate58inter1), .O(N246));
xor2 gate59( .a(N203), .b(N177), .O(N247) );
nand2 gate60( .a(N213), .b(N24), .O(N250) );
xor2 gate61( .a(N203), .b(N180), .O(N251) );

  xor2  gate511(.a(N37), .b(N213), .O(gate62inter0));
  nand2 gate512(.a(gate62inter0), .b(s_50), .O(gate62inter1));
  and2  gate513(.a(N37), .b(N213), .O(gate62inter2));
  inv1  gate514(.a(s_50), .O(gate62inter3));
  inv1  gate515(.a(s_51), .O(gate62inter4));
  nand2 gate516(.a(gate62inter4), .b(gate62inter3), .O(gate62inter5));
  nor2  gate517(.a(gate62inter5), .b(gate62inter2), .O(gate62inter6));
  inv1  gate518(.a(N213), .O(gate62inter7));
  inv1  gate519(.a(N37), .O(gate62inter8));
  nand2 gate520(.a(gate62inter8), .b(gate62inter7), .O(gate62inter9));
  nand2 gate521(.a(s_51), .b(gate62inter3), .O(gate62inter10));
  nor2  gate522(.a(gate62inter10), .b(gate62inter9), .O(gate62inter11));
  nor2  gate523(.a(gate62inter11), .b(gate62inter6), .O(gate62inter12));
  nand2 gate524(.a(gate62inter12), .b(gate62inter1), .O(N254));
nand2 gate63( .a(N213), .b(N50), .O(N255) );
nand2 gate64( .a(N213), .b(N63), .O(N256) );
nand2 gate65( .a(N213), .b(N76), .O(N257) );
nand2 gate66( .a(N213), .b(N89), .O(N258) );
nand2 gate67( .a(N213), .b(N102), .O(N259) );
nand2 gate68( .a(N224), .b(N157), .O(N260) );
nand2 gate69( .a(N224), .b(N158), .O(N263) );

  xor2  gate273(.a(N183), .b(N227), .O(gate70inter0));
  nand2 gate274(.a(gate70inter0), .b(s_16), .O(gate70inter1));
  and2  gate275(.a(N183), .b(N227), .O(gate70inter2));
  inv1  gate276(.a(s_16), .O(gate70inter3));
  inv1  gate277(.a(s_17), .O(gate70inter4));
  nand2 gate278(.a(gate70inter4), .b(gate70inter3), .O(gate70inter5));
  nor2  gate279(.a(gate70inter5), .b(gate70inter2), .O(gate70inter6));
  inv1  gate280(.a(N227), .O(gate70inter7));
  inv1  gate281(.a(N183), .O(gate70inter8));
  nand2 gate282(.a(gate70inter8), .b(gate70inter7), .O(gate70inter9));
  nand2 gate283(.a(s_17), .b(gate70inter3), .O(gate70inter10));
  nor2  gate284(.a(gate70inter10), .b(gate70inter9), .O(gate70inter11));
  nor2  gate285(.a(gate70inter11), .b(gate70inter6), .O(gate70inter12));
  nand2 gate286(.a(gate70inter12), .b(gate70inter1), .O(N264));
nand2 gate71( .a(N230), .b(N185), .O(N267) );

  xor2  gate329(.a(N187), .b(N233), .O(gate72inter0));
  nand2 gate330(.a(gate72inter0), .b(s_24), .O(gate72inter1));
  and2  gate331(.a(N187), .b(N233), .O(gate72inter2));
  inv1  gate332(.a(s_24), .O(gate72inter3));
  inv1  gate333(.a(s_25), .O(gate72inter4));
  nand2 gate334(.a(gate72inter4), .b(gate72inter3), .O(gate72inter5));
  nor2  gate335(.a(gate72inter5), .b(gate72inter2), .O(gate72inter6));
  inv1  gate336(.a(N233), .O(gate72inter7));
  inv1  gate337(.a(N187), .O(gate72inter8));
  nand2 gate338(.a(gate72inter8), .b(gate72inter7), .O(gate72inter9));
  nand2 gate339(.a(s_25), .b(gate72inter3), .O(gate72inter10));
  nor2  gate340(.a(gate72inter10), .b(gate72inter9), .O(gate72inter11));
  nor2  gate341(.a(gate72inter11), .b(gate72inter6), .O(gate72inter12));
  nand2 gate342(.a(gate72inter12), .b(gate72inter1), .O(N270));
nand2 gate73( .a(N236), .b(N189), .O(N273) );
nand2 gate74( .a(N239), .b(N191), .O(N276) );

  xor2  gate455(.a(N193), .b(N243), .O(gate75inter0));
  nand2 gate456(.a(gate75inter0), .b(s_42), .O(gate75inter1));
  and2  gate457(.a(N193), .b(N243), .O(gate75inter2));
  inv1  gate458(.a(s_42), .O(gate75inter3));
  inv1  gate459(.a(s_43), .O(gate75inter4));
  nand2 gate460(.a(gate75inter4), .b(gate75inter3), .O(gate75inter5));
  nor2  gate461(.a(gate75inter5), .b(gate75inter2), .O(gate75inter6));
  inv1  gate462(.a(N243), .O(gate75inter7));
  inv1  gate463(.a(N193), .O(gate75inter8));
  nand2 gate464(.a(gate75inter8), .b(gate75inter7), .O(gate75inter9));
  nand2 gate465(.a(s_43), .b(gate75inter3), .O(gate75inter10));
  nor2  gate466(.a(gate75inter10), .b(gate75inter9), .O(gate75inter11));
  nor2  gate467(.a(gate75inter11), .b(gate75inter6), .O(gate75inter12));
  nand2 gate468(.a(gate75inter12), .b(gate75inter1), .O(N279));
nand2 gate76( .a(N247), .b(N195), .O(N282) );

  xor2  gate343(.a(N197), .b(N251), .O(gate77inter0));
  nand2 gate344(.a(gate77inter0), .b(s_26), .O(gate77inter1));
  and2  gate345(.a(N197), .b(N251), .O(gate77inter2));
  inv1  gate346(.a(s_26), .O(gate77inter3));
  inv1  gate347(.a(s_27), .O(gate77inter4));
  nand2 gate348(.a(gate77inter4), .b(gate77inter3), .O(gate77inter5));
  nor2  gate349(.a(gate77inter5), .b(gate77inter2), .O(gate77inter6));
  inv1  gate350(.a(N251), .O(gate77inter7));
  inv1  gate351(.a(N197), .O(gate77inter8));
  nand2 gate352(.a(gate77inter8), .b(gate77inter7), .O(gate77inter9));
  nand2 gate353(.a(s_27), .b(gate77inter3), .O(gate77inter10));
  nor2  gate354(.a(gate77inter10), .b(gate77inter9), .O(gate77inter11));
  nor2  gate355(.a(gate77inter11), .b(gate77inter6), .O(gate77inter12));
  nand2 gate356(.a(gate77inter12), .b(gate77inter1), .O(N285));
nand2 gate78( .a(N227), .b(N184), .O(N288) );
nand2 gate79( .a(N230), .b(N186), .O(N289) );

  xor2  gate245(.a(N188), .b(N233), .O(gate80inter0));
  nand2 gate246(.a(gate80inter0), .b(s_12), .O(gate80inter1));
  and2  gate247(.a(N188), .b(N233), .O(gate80inter2));
  inv1  gate248(.a(s_12), .O(gate80inter3));
  inv1  gate249(.a(s_13), .O(gate80inter4));
  nand2 gate250(.a(gate80inter4), .b(gate80inter3), .O(gate80inter5));
  nor2  gate251(.a(gate80inter5), .b(gate80inter2), .O(gate80inter6));
  inv1  gate252(.a(N233), .O(gate80inter7));
  inv1  gate253(.a(N188), .O(gate80inter8));
  nand2 gate254(.a(gate80inter8), .b(gate80inter7), .O(gate80inter9));
  nand2 gate255(.a(s_13), .b(gate80inter3), .O(gate80inter10));
  nor2  gate256(.a(gate80inter10), .b(gate80inter9), .O(gate80inter11));
  nor2  gate257(.a(gate80inter11), .b(gate80inter6), .O(gate80inter12));
  nand2 gate258(.a(gate80inter12), .b(gate80inter1), .O(N290));
nand2 gate81( .a(N236), .b(N190), .O(N291) );
nand2 gate82( .a(N239), .b(N192), .O(N292) );
nand2 gate83( .a(N243), .b(N194), .O(N293) );
nand2 gate84( .a(N247), .b(N196), .O(N294) );

  xor2  gate441(.a(N198), .b(N251), .O(gate85inter0));
  nand2 gate442(.a(gate85inter0), .b(s_40), .O(gate85inter1));
  and2  gate443(.a(N198), .b(N251), .O(gate85inter2));
  inv1  gate444(.a(s_40), .O(gate85inter3));
  inv1  gate445(.a(s_41), .O(gate85inter4));
  nand2 gate446(.a(gate85inter4), .b(gate85inter3), .O(gate85inter5));
  nor2  gate447(.a(gate85inter5), .b(gate85inter2), .O(gate85inter6));
  inv1  gate448(.a(N251), .O(gate85inter7));
  inv1  gate449(.a(N198), .O(gate85inter8));
  nand2 gate450(.a(gate85inter8), .b(gate85inter7), .O(gate85inter9));
  nand2 gate451(.a(s_41), .b(gate85inter3), .O(gate85inter10));
  nor2  gate452(.a(gate85inter10), .b(gate85inter9), .O(gate85inter11));
  nor2  gate453(.a(gate85inter11), .b(gate85inter6), .O(gate85inter12));
  nand2 gate454(.a(gate85inter12), .b(gate85inter1), .O(N295));
and9 gate86( .a(N260), .b(N264), .c(N267), .d(N270), .e(N273), .f(N276), .g(N279), .h(N282), .i(N285), .O(N296) );
inv1 gate87( .a(N263), .O(N300) );
inv1 gate88( .a(N288), .O(N301) );
inv1 gate89( .a(N289), .O(N302) );
inv1 gate90( .a(N290), .O(N303) );
inv1 gate91( .a(N291), .O(N304) );
inv1 gate92( .a(N292), .O(N305) );
inv1 gate93( .a(N293), .O(N306) );
inv1 gate94( .a(N294), .O(N307) );
inv1 gate95( .a(N295), .O(N308) );
inv1 gate96( .a(N296), .O(N309) );
inv1 gate97( .a(N296), .O(N319) );
inv1 gate98( .a(N296), .O(N329) );
xor2 gate99( .a(N309), .b(N260), .O(N330) );
xor2 gate100( .a(N309), .b(N264), .O(N331) );
xor2 gate101( .a(N309), .b(N267), .O(N332) );
xor2 gate102( .a(N309), .b(N270), .O(N333) );
nand2 gate103( .a(N8), .b(N319), .O(N334) );
xor2 gate104( .a(N309), .b(N273), .O(N335) );
nand2 gate105( .a(N319), .b(N21), .O(N336) );
xor2 gate106( .a(N309), .b(N276), .O(N337) );
nand2 gate107( .a(N319), .b(N34), .O(N338) );
xor2 gate108( .a(N309), .b(N279), .O(N339) );
nand2 gate109( .a(N319), .b(N47), .O(N340) );
xor2 gate110( .a(N309), .b(N282), .O(N341) );

  xor2  gate483(.a(N60), .b(N319), .O(gate111inter0));
  nand2 gate484(.a(gate111inter0), .b(s_46), .O(gate111inter1));
  and2  gate485(.a(N60), .b(N319), .O(gate111inter2));
  inv1  gate486(.a(s_46), .O(gate111inter3));
  inv1  gate487(.a(s_47), .O(gate111inter4));
  nand2 gate488(.a(gate111inter4), .b(gate111inter3), .O(gate111inter5));
  nor2  gate489(.a(gate111inter5), .b(gate111inter2), .O(gate111inter6));
  inv1  gate490(.a(N319), .O(gate111inter7));
  inv1  gate491(.a(N60), .O(gate111inter8));
  nand2 gate492(.a(gate111inter8), .b(gate111inter7), .O(gate111inter9));
  nand2 gate493(.a(s_47), .b(gate111inter3), .O(gate111inter10));
  nor2  gate494(.a(gate111inter10), .b(gate111inter9), .O(gate111inter11));
  nor2  gate495(.a(gate111inter11), .b(gate111inter6), .O(gate111inter12));
  nand2 gate496(.a(gate111inter12), .b(gate111inter1), .O(N342));
xor2 gate112( .a(N309), .b(N285), .O(N343) );

  xor2  gate315(.a(N73), .b(N319), .O(gate113inter0));
  nand2 gate316(.a(gate113inter0), .b(s_22), .O(gate113inter1));
  and2  gate317(.a(N73), .b(N319), .O(gate113inter2));
  inv1  gate318(.a(s_22), .O(gate113inter3));
  inv1  gate319(.a(s_23), .O(gate113inter4));
  nand2 gate320(.a(gate113inter4), .b(gate113inter3), .O(gate113inter5));
  nor2  gate321(.a(gate113inter5), .b(gate113inter2), .O(gate113inter6));
  inv1  gate322(.a(N319), .O(gate113inter7));
  inv1  gate323(.a(N73), .O(gate113inter8));
  nand2 gate324(.a(gate113inter8), .b(gate113inter7), .O(gate113inter9));
  nand2 gate325(.a(s_23), .b(gate113inter3), .O(gate113inter10));
  nor2  gate326(.a(gate113inter10), .b(gate113inter9), .O(gate113inter11));
  nor2  gate327(.a(gate113inter11), .b(gate113inter6), .O(gate113inter12));
  nand2 gate328(.a(gate113inter12), .b(gate113inter1), .O(N344));
nand2 gate114( .a(N319), .b(N86), .O(N345) );
nand2 gate115( .a(N319), .b(N99), .O(N346) );
nand2 gate116( .a(N319), .b(N112), .O(N347) );
nand2 gate117( .a(N330), .b(N300), .O(N348) );

  xor2  gate217(.a(N301), .b(N331), .O(gate118inter0));
  nand2 gate218(.a(gate118inter0), .b(s_8), .O(gate118inter1));
  and2  gate219(.a(N301), .b(N331), .O(gate118inter2));
  inv1  gate220(.a(s_8), .O(gate118inter3));
  inv1  gate221(.a(s_9), .O(gate118inter4));
  nand2 gate222(.a(gate118inter4), .b(gate118inter3), .O(gate118inter5));
  nor2  gate223(.a(gate118inter5), .b(gate118inter2), .O(gate118inter6));
  inv1  gate224(.a(N331), .O(gate118inter7));
  inv1  gate225(.a(N301), .O(gate118inter8));
  nand2 gate226(.a(gate118inter8), .b(gate118inter7), .O(gate118inter9));
  nand2 gate227(.a(s_9), .b(gate118inter3), .O(gate118inter10));
  nor2  gate228(.a(gate118inter10), .b(gate118inter9), .O(gate118inter11));
  nor2  gate229(.a(gate118inter11), .b(gate118inter6), .O(gate118inter12));
  nand2 gate230(.a(gate118inter12), .b(gate118inter1), .O(N349));

  xor2  gate385(.a(N302), .b(N332), .O(gate119inter0));
  nand2 gate386(.a(gate119inter0), .b(s_32), .O(gate119inter1));
  and2  gate387(.a(N302), .b(N332), .O(gate119inter2));
  inv1  gate388(.a(s_32), .O(gate119inter3));
  inv1  gate389(.a(s_33), .O(gate119inter4));
  nand2 gate390(.a(gate119inter4), .b(gate119inter3), .O(gate119inter5));
  nor2  gate391(.a(gate119inter5), .b(gate119inter2), .O(gate119inter6));
  inv1  gate392(.a(N332), .O(gate119inter7));
  inv1  gate393(.a(N302), .O(gate119inter8));
  nand2 gate394(.a(gate119inter8), .b(gate119inter7), .O(gate119inter9));
  nand2 gate395(.a(s_33), .b(gate119inter3), .O(gate119inter10));
  nor2  gate396(.a(gate119inter10), .b(gate119inter9), .O(gate119inter11));
  nor2  gate397(.a(gate119inter11), .b(gate119inter6), .O(gate119inter12));
  nand2 gate398(.a(gate119inter12), .b(gate119inter1), .O(N350));
nand2 gate120( .a(N333), .b(N303), .O(N351) );
nand2 gate121( .a(N335), .b(N304), .O(N352) );
nand2 gate122( .a(N337), .b(N305), .O(N353) );

  xor2  gate231(.a(N306), .b(N339), .O(gate123inter0));
  nand2 gate232(.a(gate123inter0), .b(s_10), .O(gate123inter1));
  and2  gate233(.a(N306), .b(N339), .O(gate123inter2));
  inv1  gate234(.a(s_10), .O(gate123inter3));
  inv1  gate235(.a(s_11), .O(gate123inter4));
  nand2 gate236(.a(gate123inter4), .b(gate123inter3), .O(gate123inter5));
  nor2  gate237(.a(gate123inter5), .b(gate123inter2), .O(gate123inter6));
  inv1  gate238(.a(N339), .O(gate123inter7));
  inv1  gate239(.a(N306), .O(gate123inter8));
  nand2 gate240(.a(gate123inter8), .b(gate123inter7), .O(gate123inter9));
  nand2 gate241(.a(s_11), .b(gate123inter3), .O(gate123inter10));
  nor2  gate242(.a(gate123inter10), .b(gate123inter9), .O(gate123inter11));
  nor2  gate243(.a(gate123inter11), .b(gate123inter6), .O(gate123inter12));
  nand2 gate244(.a(gate123inter12), .b(gate123inter1), .O(N354));
nand2 gate124( .a(N341), .b(N307), .O(N355) );
nand2 gate125( .a(N343), .b(N308), .O(N356) );
and9 gate126( .a(N348), .b(N349), .c(N350), .d(N351), .e(N352), .f(N353), .g(N354), .h(N355), .i(N356), .O(N357) );
inv1 gate127( .a(N357), .O(N360) );
inv1 gate128( .a(N357), .O(N370) );

  xor2  gate427(.a(N360), .b(N14), .O(gate129inter0));
  nand2 gate428(.a(gate129inter0), .b(s_38), .O(gate129inter1));
  and2  gate429(.a(N360), .b(N14), .O(gate129inter2));
  inv1  gate430(.a(s_38), .O(gate129inter3));
  inv1  gate431(.a(s_39), .O(gate129inter4));
  nand2 gate432(.a(gate129inter4), .b(gate129inter3), .O(gate129inter5));
  nor2  gate433(.a(gate129inter5), .b(gate129inter2), .O(gate129inter6));
  inv1  gate434(.a(N14), .O(gate129inter7));
  inv1  gate435(.a(N360), .O(gate129inter8));
  nand2 gate436(.a(gate129inter8), .b(gate129inter7), .O(gate129inter9));
  nand2 gate437(.a(s_39), .b(gate129inter3), .O(gate129inter10));
  nor2  gate438(.a(gate129inter10), .b(gate129inter9), .O(gate129inter11));
  nor2  gate439(.a(gate129inter11), .b(gate129inter6), .O(gate129inter12));
  nand2 gate440(.a(gate129inter12), .b(gate129inter1), .O(N371));
nand2 gate130( .a(N360), .b(N27), .O(N372) );
nand2 gate131( .a(N360), .b(N40), .O(N373) );
nand2 gate132( .a(N360), .b(N53), .O(N374) );
nand2 gate133( .a(N360), .b(N66), .O(N375) );
nand2 gate134( .a(N360), .b(N79), .O(N376) );
nand2 gate135( .a(N360), .b(N92), .O(N377) );

  xor2  gate301(.a(N105), .b(N360), .O(gate136inter0));
  nand2 gate302(.a(gate136inter0), .b(s_20), .O(gate136inter1));
  and2  gate303(.a(N105), .b(N360), .O(gate136inter2));
  inv1  gate304(.a(s_20), .O(gate136inter3));
  inv1  gate305(.a(s_21), .O(gate136inter4));
  nand2 gate306(.a(gate136inter4), .b(gate136inter3), .O(gate136inter5));
  nor2  gate307(.a(gate136inter5), .b(gate136inter2), .O(gate136inter6));
  inv1  gate308(.a(N360), .O(gate136inter7));
  inv1  gate309(.a(N105), .O(gate136inter8));
  nand2 gate310(.a(gate136inter8), .b(gate136inter7), .O(gate136inter9));
  nand2 gate311(.a(s_21), .b(gate136inter3), .O(gate136inter10));
  nor2  gate312(.a(gate136inter10), .b(gate136inter9), .O(gate136inter11));
  nor2  gate313(.a(gate136inter11), .b(gate136inter6), .O(gate136inter12));
  nand2 gate314(.a(gate136inter12), .b(gate136inter1), .O(N378));
nand2 gate137( .a(N360), .b(N115), .O(N379) );
nand4 gate138( .a(N4), .b(N242), .c(N334), .d(N371), .O(N380) );
nand4 gate139( .a(N246), .b(N336), .c(N372), .d(N17), .O(N381) );
nand4 gate140( .a(N250), .b(N338), .c(N373), .d(N30), .O(N386) );
nand4 gate141( .a(N254), .b(N340), .c(N374), .d(N43), .O(N393) );
nand4 gate142( .a(N255), .b(N342), .c(N375), .d(N56), .O(N399) );
nand4 gate143( .a(N256), .b(N344), .c(N376), .d(N69), .O(N404) );
nand4 gate144( .a(N257), .b(N345), .c(N377), .d(N82), .O(N407) );
nand4 gate145( .a(N258), .b(N346), .c(N378), .d(N95), .O(N411) );
nand4 gate146( .a(N259), .b(N347), .c(N379), .d(N108), .O(N414) );
inv1 gate147( .a(N380), .O(N415) );
and8 gate148( .a(N381), .b(N386), .c(N393), .d(N399), .e(N404), .f(N407), .g(N411), .h(N414), .O(N416) );
inv1 gate149( .a(N393), .O(N417) );
inv1 gate150( .a(N404), .O(N418) );
inv1 gate151( .a(N407), .O(N419) );
inv1 gate152( .a(N411), .O(N420) );
nor2 gate153( .a(N415), .b(N416), .O(N421) );

  xor2  gate203(.a(N417), .b(N386), .O(gate154inter0));
  nand2 gate204(.a(gate154inter0), .b(s_6), .O(gate154inter1));
  and2  gate205(.a(N417), .b(N386), .O(gate154inter2));
  inv1  gate206(.a(s_6), .O(gate154inter3));
  inv1  gate207(.a(s_7), .O(gate154inter4));
  nand2 gate208(.a(gate154inter4), .b(gate154inter3), .O(gate154inter5));
  nor2  gate209(.a(gate154inter5), .b(gate154inter2), .O(gate154inter6));
  inv1  gate210(.a(N386), .O(gate154inter7));
  inv1  gate211(.a(N417), .O(gate154inter8));
  nand2 gate212(.a(gate154inter8), .b(gate154inter7), .O(gate154inter9));
  nand2 gate213(.a(s_7), .b(gate154inter3), .O(gate154inter10));
  nor2  gate214(.a(gate154inter10), .b(gate154inter9), .O(gate154inter11));
  nor2  gate215(.a(gate154inter11), .b(gate154inter6), .O(gate154inter12));
  nand2 gate216(.a(gate154inter12), .b(gate154inter1), .O(N422));
nand4 gate155( .a(N386), .b(N393), .c(N418), .d(N399), .O(N425) );
nand3 gate156( .a(N399), .b(N393), .c(N419), .O(N428) );
nand4 gate157( .a(N386), .b(N393), .c(N407), .d(N420), .O(N429) );
nand4 gate158( .a(N381), .b(N386), .c(N422), .d(N399), .O(N430) );
nand4 gate159( .a(N381), .b(N386), .c(N425), .d(N428), .O(N431) );
nand4 gate160( .a(N381), .b(N422), .c(N425), .d(N429), .O(N432) );

endmodule