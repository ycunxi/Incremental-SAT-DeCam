module c432 (N1,N4,N8,N11,N14,N17,N21,N24,N27,N30,
             N34,N37,N40,N43,N47,N50,N53,N56,N60,N63,
             N66,N69,N73,N76,N79,N82,N86,N89,N92,N95,
             N99,N102,N105,N108,N112,N115,N223,N329,N370,N421,
             N430,N431,N432);

input N1,N4,N8,N11,N14,N17,N21,N24,N27,N30,
      N34,N37,N40,N43,N47,N50,N53,N56,N60,N63,
      N66,N69,N73,N76,N79,N82,N86,N89,N92,N95,
      N99,N102,N105,N108,N112,N115;//RE__PI;

input s_0,s_1;//RE__ALLOW(00,01,10,11);
input s_2,s_3;//RE__ALLOW(00,01,10,11);
input s_4,s_5;//RE__ALLOW(00,01,10,11);
input s_6,s_7;//RE__ALLOW(00,01,10,11);
input s_8,s_9;//RE__ALLOW(00,01,10,11);
input s_10,s_11;//RE__ALLOW(00,01,10,11);
input s_12,s_13;//RE__ALLOW(00,01,10,11);
input s_14,s_15;//RE__ALLOW(00,01,10,11);
input s_16,s_17;//RE__ALLOW(00,01,10,11);
input s_18,s_19;//RE__ALLOW(00,01,10,11);
input s_20,s_21;//RE__ALLOW(00,01,10,11);
input s_22,s_23;//RE__ALLOW(00,01,10,11);
input s_24,s_25;//RE__ALLOW(00,01,10,11);
input s_26,s_27;//RE__ALLOW(00,01,10,11);
input s_28,s_29;//RE__ALLOW(00,01,10,11);
input s_30,s_31;//RE__ALLOW(00,01,10,11);
input s_32,s_33;//RE__ALLOW(00,01,10,11);
input s_34,s_35;//RE__ALLOW(00,01,10,11);
input s_36,s_37;//RE__ALLOW(00,01,10,11);
input s_38,s_39;//RE__ALLOW(00,01,10,11);
input s_40,s_41;//RE__ALLOW(00,01,10,11);
input s_42,s_43;//RE__ALLOW(00,01,10,11);
input s_44,s_45;//RE__ALLOW(00,01,10,11);
input s_46,s_47;//RE__ALLOW(00,01,10,11);
input s_48,s_49;//RE__ALLOW(00,01,10,11);
input s_50,s_51;//RE__ALLOW(00,01,10,11);
output N223,N329,N370,N421,N430,N431,N432;

wire N118,N119,N122,N123,N126,N127,N130,N131,N134,N135,
     N138,N139,N142,N143,N146,N147,N150,N151,N154,N157,
     N158,N159,N162,N165,N168,N171,N174,N177,N180,N183,
     N184,N185,N186,N187,N188,N189,N190,N191,N192,N193,
     N194,N195,N196,N197,N198,N199,N203,N213,N224,N227,
     N230,N233,N236,N239,N242,N243,N246,N247,N250,N251,
     N254,N255,N256,N257,N258,N259,N260,N263,N264,N267,
     N270,N273,N276,N279,N282,N285,N288,N289,N290,N291,
     N292,N293,N294,N295,N296,N300,N301,N302,N303,N304,
     N305,N306,N307,N308,N309,N319,N330,N331,N332,N333,
     N334,N335,N336,N337,N338,N339,N340,N341,N342,N343,
     N344,N345,N346,N347,N348,N349,N350,N351,N352,N353,
     N354,N355,N356,N357,N360,N371,N372,N373,N374,N375,
     N376,N377,N378,N379,N380,N381,N386,N393,N399,N404,
     N407,N411,N414,N415,N416,N417,N418,N419,N420,N422,
     N425,N428,N429, gate23inter0, gate23inter1, gate23inter2, gate23inter3, gate23inter4, gate23inter5, gate23inter6, gate23inter7, gate23inter8, gate23inter9, gate23inter10, gate23inter11, gate23inter12, gate29inter0, gate29inter1, gate29inter2, gate29inter3, gate29inter4, gate29inter5, gate29inter6, gate29inter7, gate29inter8, gate29inter9, gate29inter10, gate29inter11, gate29inter12, gate25inter0, gate25inter1, gate25inter2, gate25inter3, gate25inter4, gate25inter5, gate25inter6, gate25inter7, gate25inter8, gate25inter9, gate25inter10, gate25inter11, gate25inter12, gate122inter0, gate122inter1, gate122inter2, gate122inter3, gate122inter4, gate122inter5, gate122inter6, gate122inter7, gate122inter8, gate122inter9, gate122inter10, gate122inter11, gate122inter12, gate83inter0, gate83inter1, gate83inter2, gate83inter3, gate83inter4, gate83inter5, gate83inter6, gate83inter7, gate83inter8, gate83inter9, gate83inter10, gate83inter11, gate83inter12, gate131inter0, gate131inter1, gate131inter2, gate131inter3, gate131inter4, gate131inter5, gate131inter6, gate131inter7, gate131inter8, gate131inter9, gate131inter10, gate131inter11, gate131inter12, gate52inter0, gate52inter1, gate52inter2, gate52inter3, gate52inter4, gate52inter5, gate52inter6, gate52inter7, gate52inter8, gate52inter9, gate52inter10, gate52inter11, gate52inter12, gate116inter0, gate116inter1, gate116inter2, gate116inter3, gate116inter4, gate116inter5, gate116inter6, gate116inter7, gate116inter8, gate116inter9, gate116inter10, gate116inter11, gate116inter12, gate103inter0, gate103inter1, gate103inter2, gate103inter3, gate103inter4, gate103inter5, gate103inter6, gate103inter7, gate103inter8, gate103inter9, gate103inter10, gate103inter11, gate103inter12, gate72inter0, gate72inter1, gate72inter2, gate72inter3, gate72inter4, gate72inter5, gate72inter6, gate72inter7, gate72inter8, gate72inter9, gate72inter10, gate72inter11, gate72inter12, gate117inter0, gate117inter1, gate117inter2, gate117inter3, gate117inter4, gate117inter5, gate117inter6, gate117inter7, gate117inter8, gate117inter9, gate117inter10, gate117inter11, gate117inter12, gate63inter0, gate63inter1, gate63inter2, gate63inter3, gate63inter4, gate63inter5, gate63inter6, gate63inter7, gate63inter8, gate63inter9, gate63inter10, gate63inter11, gate63inter12, gate77inter0, gate77inter1, gate77inter2, gate77inter3, gate77inter4, gate77inter5, gate77inter6, gate77inter7, gate77inter8, gate77inter9, gate77inter10, gate77inter11, gate77inter12, gate50inter0, gate50inter1, gate50inter2, gate50inter3, gate50inter4, gate50inter5, gate50inter6, gate50inter7, gate50inter8, gate50inter9, gate50inter10, gate50inter11, gate50inter12, gate120inter0, gate120inter1, gate120inter2, gate120inter3, gate120inter4, gate120inter5, gate120inter6, gate120inter7, gate120inter8, gate120inter9, gate120inter10, gate120inter11, gate120inter12, gate113inter0, gate113inter1, gate113inter2, gate113inter3, gate113inter4, gate113inter5, gate113inter6, gate113inter7, gate113inter8, gate113inter9, gate113inter10, gate113inter11, gate113inter12, gate26inter0, gate26inter1, gate26inter2, gate26inter3, gate26inter4, gate26inter5, gate26inter6, gate26inter7, gate26inter8, gate26inter9, gate26inter10, gate26inter11, gate26inter12, gate59inter0, gate59inter1, gate59inter2, gate59inter3, gate59inter4, gate59inter5, gate59inter6, gate59inter7, gate59inter8, gate59inter9, gate59inter10, gate59inter11, gate59inter12, gate57inter0, gate57inter1, gate57inter2, gate57inter3, gate57inter4, gate57inter5, gate57inter6, gate57inter7, gate57inter8, gate57inter9, gate57inter10, gate57inter11, gate57inter12, gate36inter0, gate36inter1, gate36inter2, gate36inter3, gate36inter4, gate36inter5, gate36inter6, gate36inter7, gate36inter8, gate36inter9, gate36inter10, gate36inter11, gate36inter12, gate71inter0, gate71inter1, gate71inter2, gate71inter3, gate71inter4, gate71inter5, gate71inter6, gate71inter7, gate71inter8, gate71inter9, gate71inter10, gate71inter11, gate71inter12, gate123inter0, gate123inter1, gate123inter2, gate123inter3, gate123inter4, gate123inter5, gate123inter6, gate123inter7, gate123inter8, gate123inter9, gate123inter10, gate123inter11, gate123inter12, gate65inter0, gate65inter1, gate65inter2, gate65inter3, gate65inter4, gate65inter5, gate65inter6, gate65inter7, gate65inter8, gate65inter9, gate65inter10, gate65inter11, gate65inter12, gate129inter0, gate129inter1, gate129inter2, gate129inter3, gate129inter4, gate129inter5, gate129inter6, gate129inter7, gate129inter8, gate129inter9, gate129inter10, gate129inter11, gate129inter12, gate70inter0, gate70inter1, gate70inter2, gate70inter3, gate70inter4, gate70inter5, gate70inter6, gate70inter7, gate70inter8, gate70inter9, gate70inter10, gate70inter11, gate70inter12, gate154inter0, gate154inter1, gate154inter2, gate154inter3, gate154inter4, gate154inter5, gate154inter6, gate154inter7, gate154inter8, gate154inter9, gate154inter10, gate154inter11, gate154inter12;



inv1 gate1( .a(N1), .O(N118) );
inv1 gate2( .a(N4), .O(N119) );
inv1 gate3( .a(N11), .O(N122) );
inv1 gate4( .a(N17), .O(N123) );
inv1 gate5( .a(N24), .O(N126) );
inv1 gate6( .a(N30), .O(N127) );
inv1 gate7( .a(N37), .O(N130) );
inv1 gate8( .a(N43), .O(N131) );
inv1 gate9( .a(N50), .O(N134) );
inv1 gate10( .a(N56), .O(N135) );
inv1 gate11( .a(N63), .O(N138) );
inv1 gate12( .a(N69), .O(N139) );
inv1 gate13( .a(N76), .O(N142) );
inv1 gate14( .a(N82), .O(N143) );
inv1 gate15( .a(N89), .O(N146) );
inv1 gate16( .a(N95), .O(N147) );
inv1 gate17( .a(N102), .O(N150) );
inv1 gate18( .a(N108), .O(N151) );
nand2 gate19( .a(N118), .b(N4), .O(N154) );
nor2 gate20( .a(N8), .b(N119), .O(N157) );
nor2 gate21( .a(N14), .b(N119), .O(N158) );
nand2 gate22( .a(N122), .b(N17), .O(N159) );

  xor2  gate161(.a(N30), .b(N126), .O(gate23inter0));
  nand2 gate162(.a(gate23inter0), .b(s_0), .O(gate23inter1));
  and2  gate163(.a(N30), .b(N126), .O(gate23inter2));
  inv1  gate164(.a(s_0), .O(gate23inter3));
  inv1  gate165(.a(s_1), .O(gate23inter4));
  nand2 gate166(.a(gate23inter4), .b(gate23inter3), .O(gate23inter5));
  nor2  gate167(.a(gate23inter5), .b(gate23inter2), .O(gate23inter6));
  inv1  gate168(.a(N126), .O(gate23inter7));
  inv1  gate169(.a(N30), .O(gate23inter8));
  nand2 gate170(.a(gate23inter8), .b(gate23inter7), .O(gate23inter9));
  nand2 gate171(.a(s_1), .b(gate23inter3), .O(gate23inter10));
  nor2  gate172(.a(gate23inter10), .b(gate23inter9), .O(gate23inter11));
  nor2  gate173(.a(gate23inter11), .b(gate23inter6), .O(gate23inter12));
  nand2 gate174(.a(gate23inter12), .b(gate23inter1), .O(N162));
nand2 gate24( .a(N130), .b(N43), .O(N165) );

  xor2  gate189(.a(N56), .b(N134), .O(gate25inter0));
  nand2 gate190(.a(gate25inter0), .b(s_4), .O(gate25inter1));
  and2  gate191(.a(N56), .b(N134), .O(gate25inter2));
  inv1  gate192(.a(s_4), .O(gate25inter3));
  inv1  gate193(.a(s_5), .O(gate25inter4));
  nand2 gate194(.a(gate25inter4), .b(gate25inter3), .O(gate25inter5));
  nor2  gate195(.a(gate25inter5), .b(gate25inter2), .O(gate25inter6));
  inv1  gate196(.a(N134), .O(gate25inter7));
  inv1  gate197(.a(N56), .O(gate25inter8));
  nand2 gate198(.a(gate25inter8), .b(gate25inter7), .O(gate25inter9));
  nand2 gate199(.a(s_5), .b(gate25inter3), .O(gate25inter10));
  nor2  gate200(.a(gate25inter10), .b(gate25inter9), .O(gate25inter11));
  nor2  gate201(.a(gate25inter11), .b(gate25inter6), .O(gate25inter12));
  nand2 gate202(.a(gate25inter12), .b(gate25inter1), .O(N168));

  xor2  gate385(.a(N69), .b(N138), .O(gate26inter0));
  nand2 gate386(.a(gate26inter0), .b(s_32), .O(gate26inter1));
  and2  gate387(.a(N69), .b(N138), .O(gate26inter2));
  inv1  gate388(.a(s_32), .O(gate26inter3));
  inv1  gate389(.a(s_33), .O(gate26inter4));
  nand2 gate390(.a(gate26inter4), .b(gate26inter3), .O(gate26inter5));
  nor2  gate391(.a(gate26inter5), .b(gate26inter2), .O(gate26inter6));
  inv1  gate392(.a(N138), .O(gate26inter7));
  inv1  gate393(.a(N69), .O(gate26inter8));
  nand2 gate394(.a(gate26inter8), .b(gate26inter7), .O(gate26inter9));
  nand2 gate395(.a(s_33), .b(gate26inter3), .O(gate26inter10));
  nor2  gate396(.a(gate26inter10), .b(gate26inter9), .O(gate26inter11));
  nor2  gate397(.a(gate26inter11), .b(gate26inter6), .O(gate26inter12));
  nand2 gate398(.a(gate26inter12), .b(gate26inter1), .O(N171));
nand2 gate27( .a(N142), .b(N82), .O(N174) );
nand2 gate28( .a(N146), .b(N95), .O(N177) );

  xor2  gate175(.a(N108), .b(N150), .O(gate29inter0));
  nand2 gate176(.a(gate29inter0), .b(s_2), .O(gate29inter1));
  and2  gate177(.a(N108), .b(N150), .O(gate29inter2));
  inv1  gate178(.a(s_2), .O(gate29inter3));
  inv1  gate179(.a(s_3), .O(gate29inter4));
  nand2 gate180(.a(gate29inter4), .b(gate29inter3), .O(gate29inter5));
  nor2  gate181(.a(gate29inter5), .b(gate29inter2), .O(gate29inter6));
  inv1  gate182(.a(N150), .O(gate29inter7));
  inv1  gate183(.a(N108), .O(gate29inter8));
  nand2 gate184(.a(gate29inter8), .b(gate29inter7), .O(gate29inter9));
  nand2 gate185(.a(s_3), .b(gate29inter3), .O(gate29inter10));
  nor2  gate186(.a(gate29inter10), .b(gate29inter9), .O(gate29inter11));
  nor2  gate187(.a(gate29inter11), .b(gate29inter6), .O(gate29inter12));
  nand2 gate188(.a(gate29inter12), .b(gate29inter1), .O(N180));
nor2 gate30( .a(N21), .b(N123), .O(N183) );
nor2 gate31( .a(N27), .b(N123), .O(N184) );
nor2 gate32( .a(N34), .b(N127), .O(N185) );
nor2 gate33( .a(N40), .b(N127), .O(N186) );
nor2 gate34( .a(N47), .b(N131), .O(N187) );
nor2 gate35( .a(N53), .b(N131), .O(N188) );

  xor2  gate427(.a(N135), .b(N60), .O(gate36inter0));
  nand2 gate428(.a(gate36inter0), .b(s_38), .O(gate36inter1));
  and2  gate429(.a(N135), .b(N60), .O(gate36inter2));
  inv1  gate430(.a(s_38), .O(gate36inter3));
  inv1  gate431(.a(s_39), .O(gate36inter4));
  nand2 gate432(.a(gate36inter4), .b(gate36inter3), .O(gate36inter5));
  nor2  gate433(.a(gate36inter5), .b(gate36inter2), .O(gate36inter6));
  inv1  gate434(.a(N60), .O(gate36inter7));
  inv1  gate435(.a(N135), .O(gate36inter8));
  nand2 gate436(.a(gate36inter8), .b(gate36inter7), .O(gate36inter9));
  nand2 gate437(.a(s_39), .b(gate36inter3), .O(gate36inter10));
  nor2  gate438(.a(gate36inter10), .b(gate36inter9), .O(gate36inter11));
  nor2  gate439(.a(gate36inter11), .b(gate36inter6), .O(gate36inter12));
  nand2 gate440(.a(gate36inter12), .b(gate36inter1), .O(N189));
nor2 gate37( .a(N66), .b(N135), .O(N190) );
nor2 gate38( .a(N73), .b(N139), .O(N191) );
nor2 gate39( .a(N79), .b(N139), .O(N192) );
nor2 gate40( .a(N86), .b(N143), .O(N193) );
nor2 gate41( .a(N92), .b(N143), .O(N194) );
nor2 gate42( .a(N99), .b(N147), .O(N195) );
nor2 gate43( .a(N105), .b(N147), .O(N196) );
nor2 gate44( .a(N112), .b(N151), .O(N197) );
nor2 gate45( .a(N115), .b(N151), .O(N198) );
and9 gate46( .a(N154), .b(N159), .c(N162), .d(N165), .e(N168), .f(N171), .g(N174), .h(N177), .i(N180), .O(N199) );
inv1 gate47( .a(N199), .O(N203) );
inv1 gate48( .a(N199), .O(N213) );
inv1 gate49( .a(N199), .O(N223) );

  xor2  gate343(.a(N154), .b(N203), .O(gate50inter0));
  nand2 gate344(.a(gate50inter0), .b(s_26), .O(gate50inter1));
  and2  gate345(.a(N154), .b(N203), .O(gate50inter2));
  inv1  gate346(.a(s_26), .O(gate50inter3));
  inv1  gate347(.a(s_27), .O(gate50inter4));
  nand2 gate348(.a(gate50inter4), .b(gate50inter3), .O(gate50inter5));
  nor2  gate349(.a(gate50inter5), .b(gate50inter2), .O(gate50inter6));
  inv1  gate350(.a(N203), .O(gate50inter7));
  inv1  gate351(.a(N154), .O(gate50inter8));
  nand2 gate352(.a(gate50inter8), .b(gate50inter7), .O(gate50inter9));
  nand2 gate353(.a(s_27), .b(gate50inter3), .O(gate50inter10));
  nor2  gate354(.a(gate50inter10), .b(gate50inter9), .O(gate50inter11));
  nor2  gate355(.a(gate50inter11), .b(gate50inter6), .O(gate50inter12));
  nand2 gate356(.a(gate50inter12), .b(gate50inter1), .O(N224));
xor2 gate51( .a(N203), .b(N159), .O(N227) );

  xor2  gate245(.a(N162), .b(N203), .O(gate52inter0));
  nand2 gate246(.a(gate52inter0), .b(s_12), .O(gate52inter1));
  and2  gate247(.a(N162), .b(N203), .O(gate52inter2));
  inv1  gate248(.a(s_12), .O(gate52inter3));
  inv1  gate249(.a(s_13), .O(gate52inter4));
  nand2 gate250(.a(gate52inter4), .b(gate52inter3), .O(gate52inter5));
  nor2  gate251(.a(gate52inter5), .b(gate52inter2), .O(gate52inter6));
  inv1  gate252(.a(N203), .O(gate52inter7));
  inv1  gate253(.a(N162), .O(gate52inter8));
  nand2 gate254(.a(gate52inter8), .b(gate52inter7), .O(gate52inter9));
  nand2 gate255(.a(s_13), .b(gate52inter3), .O(gate52inter10));
  nor2  gate256(.a(gate52inter10), .b(gate52inter9), .O(gate52inter11));
  nor2  gate257(.a(gate52inter11), .b(gate52inter6), .O(gate52inter12));
  nand2 gate258(.a(gate52inter12), .b(gate52inter1), .O(N230));
xor2 gate53( .a(N203), .b(N165), .O(N233) );
xor2 gate54( .a(N203), .b(N168), .O(N236) );
xor2 gate55( .a(N203), .b(N171), .O(N239) );
nand2 gate56( .a(N1), .b(N213), .O(N242) );

  xor2  gate413(.a(N174), .b(N203), .O(gate57inter0));
  nand2 gate414(.a(gate57inter0), .b(s_36), .O(gate57inter1));
  and2  gate415(.a(N174), .b(N203), .O(gate57inter2));
  inv1  gate416(.a(s_36), .O(gate57inter3));
  inv1  gate417(.a(s_37), .O(gate57inter4));
  nand2 gate418(.a(gate57inter4), .b(gate57inter3), .O(gate57inter5));
  nor2  gate419(.a(gate57inter5), .b(gate57inter2), .O(gate57inter6));
  inv1  gate420(.a(N203), .O(gate57inter7));
  inv1  gate421(.a(N174), .O(gate57inter8));
  nand2 gate422(.a(gate57inter8), .b(gate57inter7), .O(gate57inter9));
  nand2 gate423(.a(s_37), .b(gate57inter3), .O(gate57inter10));
  nor2  gate424(.a(gate57inter10), .b(gate57inter9), .O(gate57inter11));
  nor2  gate425(.a(gate57inter11), .b(gate57inter6), .O(gate57inter12));
  nand2 gate426(.a(gate57inter12), .b(gate57inter1), .O(N243));
nand2 gate58( .a(N213), .b(N11), .O(N246) );

  xor2  gate399(.a(N177), .b(N203), .O(gate59inter0));
  nand2 gate400(.a(gate59inter0), .b(s_34), .O(gate59inter1));
  and2  gate401(.a(N177), .b(N203), .O(gate59inter2));
  inv1  gate402(.a(s_34), .O(gate59inter3));
  inv1  gate403(.a(s_35), .O(gate59inter4));
  nand2 gate404(.a(gate59inter4), .b(gate59inter3), .O(gate59inter5));
  nor2  gate405(.a(gate59inter5), .b(gate59inter2), .O(gate59inter6));
  inv1  gate406(.a(N203), .O(gate59inter7));
  inv1  gate407(.a(N177), .O(gate59inter8));
  nand2 gate408(.a(gate59inter8), .b(gate59inter7), .O(gate59inter9));
  nand2 gate409(.a(s_35), .b(gate59inter3), .O(gate59inter10));
  nor2  gate410(.a(gate59inter10), .b(gate59inter9), .O(gate59inter11));
  nor2  gate411(.a(gate59inter11), .b(gate59inter6), .O(gate59inter12));
  nand2 gate412(.a(gate59inter12), .b(gate59inter1), .O(N247));
nand2 gate60( .a(N213), .b(N24), .O(N250) );
xor2 gate61( .a(N203), .b(N180), .O(N251) );
nand2 gate62( .a(N213), .b(N37), .O(N254) );

  xor2  gate315(.a(N50), .b(N213), .O(gate63inter0));
  nand2 gate316(.a(gate63inter0), .b(s_22), .O(gate63inter1));
  and2  gate317(.a(N50), .b(N213), .O(gate63inter2));
  inv1  gate318(.a(s_22), .O(gate63inter3));
  inv1  gate319(.a(s_23), .O(gate63inter4));
  nand2 gate320(.a(gate63inter4), .b(gate63inter3), .O(gate63inter5));
  nor2  gate321(.a(gate63inter5), .b(gate63inter2), .O(gate63inter6));
  inv1  gate322(.a(N213), .O(gate63inter7));
  inv1  gate323(.a(N50), .O(gate63inter8));
  nand2 gate324(.a(gate63inter8), .b(gate63inter7), .O(gate63inter9));
  nand2 gate325(.a(s_23), .b(gate63inter3), .O(gate63inter10));
  nor2  gate326(.a(gate63inter10), .b(gate63inter9), .O(gate63inter11));
  nor2  gate327(.a(gate63inter11), .b(gate63inter6), .O(gate63inter12));
  nand2 gate328(.a(gate63inter12), .b(gate63inter1), .O(N255));
nand2 gate64( .a(N213), .b(N63), .O(N256) );

  xor2  gate469(.a(N76), .b(N213), .O(gate65inter0));
  nand2 gate470(.a(gate65inter0), .b(s_44), .O(gate65inter1));
  and2  gate471(.a(N76), .b(N213), .O(gate65inter2));
  inv1  gate472(.a(s_44), .O(gate65inter3));
  inv1  gate473(.a(s_45), .O(gate65inter4));
  nand2 gate474(.a(gate65inter4), .b(gate65inter3), .O(gate65inter5));
  nor2  gate475(.a(gate65inter5), .b(gate65inter2), .O(gate65inter6));
  inv1  gate476(.a(N213), .O(gate65inter7));
  inv1  gate477(.a(N76), .O(gate65inter8));
  nand2 gate478(.a(gate65inter8), .b(gate65inter7), .O(gate65inter9));
  nand2 gate479(.a(s_45), .b(gate65inter3), .O(gate65inter10));
  nor2  gate480(.a(gate65inter10), .b(gate65inter9), .O(gate65inter11));
  nor2  gate481(.a(gate65inter11), .b(gate65inter6), .O(gate65inter12));
  nand2 gate482(.a(gate65inter12), .b(gate65inter1), .O(N257));
nand2 gate66( .a(N213), .b(N89), .O(N258) );
nand2 gate67( .a(N213), .b(N102), .O(N259) );
nand2 gate68( .a(N224), .b(N157), .O(N260) );
nand2 gate69( .a(N224), .b(N158), .O(N263) );

  xor2  gate497(.a(N183), .b(N227), .O(gate70inter0));
  nand2 gate498(.a(gate70inter0), .b(s_48), .O(gate70inter1));
  and2  gate499(.a(N183), .b(N227), .O(gate70inter2));
  inv1  gate500(.a(s_48), .O(gate70inter3));
  inv1  gate501(.a(s_49), .O(gate70inter4));
  nand2 gate502(.a(gate70inter4), .b(gate70inter3), .O(gate70inter5));
  nor2  gate503(.a(gate70inter5), .b(gate70inter2), .O(gate70inter6));
  inv1  gate504(.a(N227), .O(gate70inter7));
  inv1  gate505(.a(N183), .O(gate70inter8));
  nand2 gate506(.a(gate70inter8), .b(gate70inter7), .O(gate70inter9));
  nand2 gate507(.a(s_49), .b(gate70inter3), .O(gate70inter10));
  nor2  gate508(.a(gate70inter10), .b(gate70inter9), .O(gate70inter11));
  nor2  gate509(.a(gate70inter11), .b(gate70inter6), .O(gate70inter12));
  nand2 gate510(.a(gate70inter12), .b(gate70inter1), .O(N264));

  xor2  gate441(.a(N185), .b(N230), .O(gate71inter0));
  nand2 gate442(.a(gate71inter0), .b(s_40), .O(gate71inter1));
  and2  gate443(.a(N185), .b(N230), .O(gate71inter2));
  inv1  gate444(.a(s_40), .O(gate71inter3));
  inv1  gate445(.a(s_41), .O(gate71inter4));
  nand2 gate446(.a(gate71inter4), .b(gate71inter3), .O(gate71inter5));
  nor2  gate447(.a(gate71inter5), .b(gate71inter2), .O(gate71inter6));
  inv1  gate448(.a(N230), .O(gate71inter7));
  inv1  gate449(.a(N185), .O(gate71inter8));
  nand2 gate450(.a(gate71inter8), .b(gate71inter7), .O(gate71inter9));
  nand2 gate451(.a(s_41), .b(gate71inter3), .O(gate71inter10));
  nor2  gate452(.a(gate71inter10), .b(gate71inter9), .O(gate71inter11));
  nor2  gate453(.a(gate71inter11), .b(gate71inter6), .O(gate71inter12));
  nand2 gate454(.a(gate71inter12), .b(gate71inter1), .O(N267));

  xor2  gate287(.a(N187), .b(N233), .O(gate72inter0));
  nand2 gate288(.a(gate72inter0), .b(s_18), .O(gate72inter1));
  and2  gate289(.a(N187), .b(N233), .O(gate72inter2));
  inv1  gate290(.a(s_18), .O(gate72inter3));
  inv1  gate291(.a(s_19), .O(gate72inter4));
  nand2 gate292(.a(gate72inter4), .b(gate72inter3), .O(gate72inter5));
  nor2  gate293(.a(gate72inter5), .b(gate72inter2), .O(gate72inter6));
  inv1  gate294(.a(N233), .O(gate72inter7));
  inv1  gate295(.a(N187), .O(gate72inter8));
  nand2 gate296(.a(gate72inter8), .b(gate72inter7), .O(gate72inter9));
  nand2 gate297(.a(s_19), .b(gate72inter3), .O(gate72inter10));
  nor2  gate298(.a(gate72inter10), .b(gate72inter9), .O(gate72inter11));
  nor2  gate299(.a(gate72inter11), .b(gate72inter6), .O(gate72inter12));
  nand2 gate300(.a(gate72inter12), .b(gate72inter1), .O(N270));
nand2 gate73( .a(N236), .b(N189), .O(N273) );
nand2 gate74( .a(N239), .b(N191), .O(N276) );
nand2 gate75( .a(N243), .b(N193), .O(N279) );
nand2 gate76( .a(N247), .b(N195), .O(N282) );

  xor2  gate329(.a(N197), .b(N251), .O(gate77inter0));
  nand2 gate330(.a(gate77inter0), .b(s_24), .O(gate77inter1));
  and2  gate331(.a(N197), .b(N251), .O(gate77inter2));
  inv1  gate332(.a(s_24), .O(gate77inter3));
  inv1  gate333(.a(s_25), .O(gate77inter4));
  nand2 gate334(.a(gate77inter4), .b(gate77inter3), .O(gate77inter5));
  nor2  gate335(.a(gate77inter5), .b(gate77inter2), .O(gate77inter6));
  inv1  gate336(.a(N251), .O(gate77inter7));
  inv1  gate337(.a(N197), .O(gate77inter8));
  nand2 gate338(.a(gate77inter8), .b(gate77inter7), .O(gate77inter9));
  nand2 gate339(.a(s_25), .b(gate77inter3), .O(gate77inter10));
  nor2  gate340(.a(gate77inter10), .b(gate77inter9), .O(gate77inter11));
  nor2  gate341(.a(gate77inter11), .b(gate77inter6), .O(gate77inter12));
  nand2 gate342(.a(gate77inter12), .b(gate77inter1), .O(N285));
nand2 gate78( .a(N227), .b(N184), .O(N288) );
nand2 gate79( .a(N230), .b(N186), .O(N289) );
nand2 gate80( .a(N233), .b(N188), .O(N290) );
nand2 gate81( .a(N236), .b(N190), .O(N291) );
nand2 gate82( .a(N239), .b(N192), .O(N292) );

  xor2  gate217(.a(N194), .b(N243), .O(gate83inter0));
  nand2 gate218(.a(gate83inter0), .b(s_8), .O(gate83inter1));
  and2  gate219(.a(N194), .b(N243), .O(gate83inter2));
  inv1  gate220(.a(s_8), .O(gate83inter3));
  inv1  gate221(.a(s_9), .O(gate83inter4));
  nand2 gate222(.a(gate83inter4), .b(gate83inter3), .O(gate83inter5));
  nor2  gate223(.a(gate83inter5), .b(gate83inter2), .O(gate83inter6));
  inv1  gate224(.a(N243), .O(gate83inter7));
  inv1  gate225(.a(N194), .O(gate83inter8));
  nand2 gate226(.a(gate83inter8), .b(gate83inter7), .O(gate83inter9));
  nand2 gate227(.a(s_9), .b(gate83inter3), .O(gate83inter10));
  nor2  gate228(.a(gate83inter10), .b(gate83inter9), .O(gate83inter11));
  nor2  gate229(.a(gate83inter11), .b(gate83inter6), .O(gate83inter12));
  nand2 gate230(.a(gate83inter12), .b(gate83inter1), .O(N293));
nand2 gate84( .a(N247), .b(N196), .O(N294) );
nand2 gate85( .a(N251), .b(N198), .O(N295) );
and9 gate86( .a(N260), .b(N264), .c(N267), .d(N270), .e(N273), .f(N276), .g(N279), .h(N282), .i(N285), .O(N296) );
inv1 gate87( .a(N263), .O(N300) );
inv1 gate88( .a(N288), .O(N301) );
inv1 gate89( .a(N289), .O(N302) );
inv1 gate90( .a(N290), .O(N303) );
inv1 gate91( .a(N291), .O(N304) );
inv1 gate92( .a(N292), .O(N305) );
inv1 gate93( .a(N293), .O(N306) );
inv1 gate94( .a(N294), .O(N307) );
inv1 gate95( .a(N295), .O(N308) );
inv1 gate96( .a(N296), .O(N309) );
inv1 gate97( .a(N296), .O(N319) );
inv1 gate98( .a(N296), .O(N329) );
xor2 gate99( .a(N309), .b(N260), .O(N330) );
xor2 gate100( .a(N309), .b(N264), .O(N331) );
xor2 gate101( .a(N309), .b(N267), .O(N332) );
xor2 gate102( .a(N309), .b(N270), .O(N333) );

  xor2  gate273(.a(N319), .b(N8), .O(gate103inter0));
  nand2 gate274(.a(gate103inter0), .b(s_16), .O(gate103inter1));
  and2  gate275(.a(N319), .b(N8), .O(gate103inter2));
  inv1  gate276(.a(s_16), .O(gate103inter3));
  inv1  gate277(.a(s_17), .O(gate103inter4));
  nand2 gate278(.a(gate103inter4), .b(gate103inter3), .O(gate103inter5));
  nor2  gate279(.a(gate103inter5), .b(gate103inter2), .O(gate103inter6));
  inv1  gate280(.a(N8), .O(gate103inter7));
  inv1  gate281(.a(N319), .O(gate103inter8));
  nand2 gate282(.a(gate103inter8), .b(gate103inter7), .O(gate103inter9));
  nand2 gate283(.a(s_17), .b(gate103inter3), .O(gate103inter10));
  nor2  gate284(.a(gate103inter10), .b(gate103inter9), .O(gate103inter11));
  nor2  gate285(.a(gate103inter11), .b(gate103inter6), .O(gate103inter12));
  nand2 gate286(.a(gate103inter12), .b(gate103inter1), .O(N334));
xor2 gate104( .a(N309), .b(N273), .O(N335) );
nand2 gate105( .a(N319), .b(N21), .O(N336) );
xor2 gate106( .a(N309), .b(N276), .O(N337) );
nand2 gate107( .a(N319), .b(N34), .O(N338) );
xor2 gate108( .a(N309), .b(N279), .O(N339) );
nand2 gate109( .a(N319), .b(N47), .O(N340) );
xor2 gate110( .a(N309), .b(N282), .O(N341) );
nand2 gate111( .a(N319), .b(N60), .O(N342) );
xor2 gate112( .a(N309), .b(N285), .O(N343) );

  xor2  gate371(.a(N73), .b(N319), .O(gate113inter0));
  nand2 gate372(.a(gate113inter0), .b(s_30), .O(gate113inter1));
  and2  gate373(.a(N73), .b(N319), .O(gate113inter2));
  inv1  gate374(.a(s_30), .O(gate113inter3));
  inv1  gate375(.a(s_31), .O(gate113inter4));
  nand2 gate376(.a(gate113inter4), .b(gate113inter3), .O(gate113inter5));
  nor2  gate377(.a(gate113inter5), .b(gate113inter2), .O(gate113inter6));
  inv1  gate378(.a(N319), .O(gate113inter7));
  inv1  gate379(.a(N73), .O(gate113inter8));
  nand2 gate380(.a(gate113inter8), .b(gate113inter7), .O(gate113inter9));
  nand2 gate381(.a(s_31), .b(gate113inter3), .O(gate113inter10));
  nor2  gate382(.a(gate113inter10), .b(gate113inter9), .O(gate113inter11));
  nor2  gate383(.a(gate113inter11), .b(gate113inter6), .O(gate113inter12));
  nand2 gate384(.a(gate113inter12), .b(gate113inter1), .O(N344));
nand2 gate114( .a(N319), .b(N86), .O(N345) );
nand2 gate115( .a(N319), .b(N99), .O(N346) );

  xor2  gate259(.a(N112), .b(N319), .O(gate116inter0));
  nand2 gate260(.a(gate116inter0), .b(s_14), .O(gate116inter1));
  and2  gate261(.a(N112), .b(N319), .O(gate116inter2));
  inv1  gate262(.a(s_14), .O(gate116inter3));
  inv1  gate263(.a(s_15), .O(gate116inter4));
  nand2 gate264(.a(gate116inter4), .b(gate116inter3), .O(gate116inter5));
  nor2  gate265(.a(gate116inter5), .b(gate116inter2), .O(gate116inter6));
  inv1  gate266(.a(N319), .O(gate116inter7));
  inv1  gate267(.a(N112), .O(gate116inter8));
  nand2 gate268(.a(gate116inter8), .b(gate116inter7), .O(gate116inter9));
  nand2 gate269(.a(s_15), .b(gate116inter3), .O(gate116inter10));
  nor2  gate270(.a(gate116inter10), .b(gate116inter9), .O(gate116inter11));
  nor2  gate271(.a(gate116inter11), .b(gate116inter6), .O(gate116inter12));
  nand2 gate272(.a(gate116inter12), .b(gate116inter1), .O(N347));

  xor2  gate301(.a(N300), .b(N330), .O(gate117inter0));
  nand2 gate302(.a(gate117inter0), .b(s_20), .O(gate117inter1));
  and2  gate303(.a(N300), .b(N330), .O(gate117inter2));
  inv1  gate304(.a(s_20), .O(gate117inter3));
  inv1  gate305(.a(s_21), .O(gate117inter4));
  nand2 gate306(.a(gate117inter4), .b(gate117inter3), .O(gate117inter5));
  nor2  gate307(.a(gate117inter5), .b(gate117inter2), .O(gate117inter6));
  inv1  gate308(.a(N330), .O(gate117inter7));
  inv1  gate309(.a(N300), .O(gate117inter8));
  nand2 gate310(.a(gate117inter8), .b(gate117inter7), .O(gate117inter9));
  nand2 gate311(.a(s_21), .b(gate117inter3), .O(gate117inter10));
  nor2  gate312(.a(gate117inter10), .b(gate117inter9), .O(gate117inter11));
  nor2  gate313(.a(gate117inter11), .b(gate117inter6), .O(gate117inter12));
  nand2 gate314(.a(gate117inter12), .b(gate117inter1), .O(N348));
nand2 gate118( .a(N331), .b(N301), .O(N349) );
nand2 gate119( .a(N332), .b(N302), .O(N350) );

  xor2  gate357(.a(N303), .b(N333), .O(gate120inter0));
  nand2 gate358(.a(gate120inter0), .b(s_28), .O(gate120inter1));
  and2  gate359(.a(N303), .b(N333), .O(gate120inter2));
  inv1  gate360(.a(s_28), .O(gate120inter3));
  inv1  gate361(.a(s_29), .O(gate120inter4));
  nand2 gate362(.a(gate120inter4), .b(gate120inter3), .O(gate120inter5));
  nor2  gate363(.a(gate120inter5), .b(gate120inter2), .O(gate120inter6));
  inv1  gate364(.a(N333), .O(gate120inter7));
  inv1  gate365(.a(N303), .O(gate120inter8));
  nand2 gate366(.a(gate120inter8), .b(gate120inter7), .O(gate120inter9));
  nand2 gate367(.a(s_29), .b(gate120inter3), .O(gate120inter10));
  nor2  gate368(.a(gate120inter10), .b(gate120inter9), .O(gate120inter11));
  nor2  gate369(.a(gate120inter11), .b(gate120inter6), .O(gate120inter12));
  nand2 gate370(.a(gate120inter12), .b(gate120inter1), .O(N351));
nand2 gate121( .a(N335), .b(N304), .O(N352) );

  xor2  gate203(.a(N305), .b(N337), .O(gate122inter0));
  nand2 gate204(.a(gate122inter0), .b(s_6), .O(gate122inter1));
  and2  gate205(.a(N305), .b(N337), .O(gate122inter2));
  inv1  gate206(.a(s_6), .O(gate122inter3));
  inv1  gate207(.a(s_7), .O(gate122inter4));
  nand2 gate208(.a(gate122inter4), .b(gate122inter3), .O(gate122inter5));
  nor2  gate209(.a(gate122inter5), .b(gate122inter2), .O(gate122inter6));
  inv1  gate210(.a(N337), .O(gate122inter7));
  inv1  gate211(.a(N305), .O(gate122inter8));
  nand2 gate212(.a(gate122inter8), .b(gate122inter7), .O(gate122inter9));
  nand2 gate213(.a(s_7), .b(gate122inter3), .O(gate122inter10));
  nor2  gate214(.a(gate122inter10), .b(gate122inter9), .O(gate122inter11));
  nor2  gate215(.a(gate122inter11), .b(gate122inter6), .O(gate122inter12));
  nand2 gate216(.a(gate122inter12), .b(gate122inter1), .O(N353));

  xor2  gate455(.a(N306), .b(N339), .O(gate123inter0));
  nand2 gate456(.a(gate123inter0), .b(s_42), .O(gate123inter1));
  and2  gate457(.a(N306), .b(N339), .O(gate123inter2));
  inv1  gate458(.a(s_42), .O(gate123inter3));
  inv1  gate459(.a(s_43), .O(gate123inter4));
  nand2 gate460(.a(gate123inter4), .b(gate123inter3), .O(gate123inter5));
  nor2  gate461(.a(gate123inter5), .b(gate123inter2), .O(gate123inter6));
  inv1  gate462(.a(N339), .O(gate123inter7));
  inv1  gate463(.a(N306), .O(gate123inter8));
  nand2 gate464(.a(gate123inter8), .b(gate123inter7), .O(gate123inter9));
  nand2 gate465(.a(s_43), .b(gate123inter3), .O(gate123inter10));
  nor2  gate466(.a(gate123inter10), .b(gate123inter9), .O(gate123inter11));
  nor2  gate467(.a(gate123inter11), .b(gate123inter6), .O(gate123inter12));
  nand2 gate468(.a(gate123inter12), .b(gate123inter1), .O(N354));
nand2 gate124( .a(N341), .b(N307), .O(N355) );
nand2 gate125( .a(N343), .b(N308), .O(N356) );
and9 gate126( .a(N348), .b(N349), .c(N350), .d(N351), .e(N352), .f(N353), .g(N354), .h(N355), .i(N356), .O(N357) );
inv1 gate127( .a(N357), .O(N360) );
inv1 gate128( .a(N357), .O(N370) );

  xor2  gate483(.a(N360), .b(N14), .O(gate129inter0));
  nand2 gate484(.a(gate129inter0), .b(s_46), .O(gate129inter1));
  and2  gate485(.a(N360), .b(N14), .O(gate129inter2));
  inv1  gate486(.a(s_46), .O(gate129inter3));
  inv1  gate487(.a(s_47), .O(gate129inter4));
  nand2 gate488(.a(gate129inter4), .b(gate129inter3), .O(gate129inter5));
  nor2  gate489(.a(gate129inter5), .b(gate129inter2), .O(gate129inter6));
  inv1  gate490(.a(N14), .O(gate129inter7));
  inv1  gate491(.a(N360), .O(gate129inter8));
  nand2 gate492(.a(gate129inter8), .b(gate129inter7), .O(gate129inter9));
  nand2 gate493(.a(s_47), .b(gate129inter3), .O(gate129inter10));
  nor2  gate494(.a(gate129inter10), .b(gate129inter9), .O(gate129inter11));
  nor2  gate495(.a(gate129inter11), .b(gate129inter6), .O(gate129inter12));
  nand2 gate496(.a(gate129inter12), .b(gate129inter1), .O(N371));
nand2 gate130( .a(N360), .b(N27), .O(N372) );

  xor2  gate231(.a(N40), .b(N360), .O(gate131inter0));
  nand2 gate232(.a(gate131inter0), .b(s_10), .O(gate131inter1));
  and2  gate233(.a(N40), .b(N360), .O(gate131inter2));
  inv1  gate234(.a(s_10), .O(gate131inter3));
  inv1  gate235(.a(s_11), .O(gate131inter4));
  nand2 gate236(.a(gate131inter4), .b(gate131inter3), .O(gate131inter5));
  nor2  gate237(.a(gate131inter5), .b(gate131inter2), .O(gate131inter6));
  inv1  gate238(.a(N360), .O(gate131inter7));
  inv1  gate239(.a(N40), .O(gate131inter8));
  nand2 gate240(.a(gate131inter8), .b(gate131inter7), .O(gate131inter9));
  nand2 gate241(.a(s_11), .b(gate131inter3), .O(gate131inter10));
  nor2  gate242(.a(gate131inter10), .b(gate131inter9), .O(gate131inter11));
  nor2  gate243(.a(gate131inter11), .b(gate131inter6), .O(gate131inter12));
  nand2 gate244(.a(gate131inter12), .b(gate131inter1), .O(N373));
nand2 gate132( .a(N360), .b(N53), .O(N374) );
nand2 gate133( .a(N360), .b(N66), .O(N375) );
nand2 gate134( .a(N360), .b(N79), .O(N376) );
nand2 gate135( .a(N360), .b(N92), .O(N377) );
nand2 gate136( .a(N360), .b(N105), .O(N378) );
nand2 gate137( .a(N360), .b(N115), .O(N379) );
nand4 gate138( .a(N4), .b(N242), .c(N334), .d(N371), .O(N380) );
nand4 gate139( .a(N246), .b(N336), .c(N372), .d(N17), .O(N381) );
nand4 gate140( .a(N250), .b(N338), .c(N373), .d(N30), .O(N386) );
nand4 gate141( .a(N254), .b(N340), .c(N374), .d(N43), .O(N393) );
nand4 gate142( .a(N255), .b(N342), .c(N375), .d(N56), .O(N399) );
nand4 gate143( .a(N256), .b(N344), .c(N376), .d(N69), .O(N404) );
nand4 gate144( .a(N257), .b(N345), .c(N377), .d(N82), .O(N407) );
nand4 gate145( .a(N258), .b(N346), .c(N378), .d(N95), .O(N411) );
nand4 gate146( .a(N259), .b(N347), .c(N379), .d(N108), .O(N414) );
inv1 gate147( .a(N380), .O(N415) );
and8 gate148( .a(N381), .b(N386), .c(N393), .d(N399), .e(N404), .f(N407), .g(N411), .h(N414), .O(N416) );
inv1 gate149( .a(N393), .O(N417) );
inv1 gate150( .a(N404), .O(N418) );
inv1 gate151( .a(N407), .O(N419) );
inv1 gate152( .a(N411), .O(N420) );
nor2 gate153( .a(N415), .b(N416), .O(N421) );

  xor2  gate511(.a(N417), .b(N386), .O(gate154inter0));
  nand2 gate512(.a(gate154inter0), .b(s_50), .O(gate154inter1));
  and2  gate513(.a(N417), .b(N386), .O(gate154inter2));
  inv1  gate514(.a(s_50), .O(gate154inter3));
  inv1  gate515(.a(s_51), .O(gate154inter4));
  nand2 gate516(.a(gate154inter4), .b(gate154inter3), .O(gate154inter5));
  nor2  gate517(.a(gate154inter5), .b(gate154inter2), .O(gate154inter6));
  inv1  gate518(.a(N386), .O(gate154inter7));
  inv1  gate519(.a(N417), .O(gate154inter8));
  nand2 gate520(.a(gate154inter8), .b(gate154inter7), .O(gate154inter9));
  nand2 gate521(.a(s_51), .b(gate154inter3), .O(gate154inter10));
  nor2  gate522(.a(gate154inter10), .b(gate154inter9), .O(gate154inter11));
  nor2  gate523(.a(gate154inter11), .b(gate154inter6), .O(gate154inter12));
  nand2 gate524(.a(gate154inter12), .b(gate154inter1), .O(N422));
nand4 gate155( .a(N386), .b(N393), .c(N418), .d(N399), .O(N425) );
nand3 gate156( .a(N399), .b(N393), .c(N419), .O(N428) );
nand4 gate157( .a(N386), .b(N393), .c(N407), .d(N420), .O(N429) );
nand4 gate158( .a(N381), .b(N386), .c(N422), .d(N399), .O(N430) );
nand4 gate159( .a(N381), .b(N386), .c(N425), .d(N428), .O(N431) );
nand4 gate160( .a(N381), .b(N422), .c(N425), .d(N429), .O(N432) );

endmodule