module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);

input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;//RE__PI;

input s_0,s_1;//RE__ALLOW(00,01,10,11);
input s_2,s_3;//RE__ALLOW(00,01,10,11);
input s_4,s_5;//RE__ALLOW(00,01,10,11);
input s_6,s_7;//RE__ALLOW(00,01,10,11);
input s_8,s_9;//RE__ALLOW(00,01,10,11);
input s_10,s_11;//RE__ALLOW(00,01,10,11);
input s_12,s_13;//RE__ALLOW(00,01,10,11);
input s_14,s_15;//RE__ALLOW(00,01,10,11);
input s_16,s_17;//RE__ALLOW(00,01,10,11);
input s_18,s_19;//RE__ALLOW(00,01,10,11);
input s_20,s_21;//RE__ALLOW(00,01,10,11);
input s_22,s_23;//RE__ALLOW(00,01,10,11);
input s_24,s_25;//RE__ALLOW(00,01,10,11);
input s_26,s_27;//RE__ALLOW(00,01,10,11);
input s_28,s_29;//RE__ALLOW(00,01,10,11);
input s_30,s_31;//RE__ALLOW(00,01,10,11);
input s_32,s_33;//RE__ALLOW(00,01,10,11);
input s_34,s_35;//RE__ALLOW(00,01,10,11);
input s_36,s_37;//RE__ALLOW(00,01,10,11);
input s_38,s_39;//RE__ALLOW(00,01,10,11);
input s_40,s_41;//RE__ALLOW(00,01,10,11);
input s_42,s_43;//RE__ALLOW(00,01,10,11);
input s_44,s_45;//RE__ALLOW(00,01,10,11);
input s_46,s_47;//RE__ALLOW(00,01,10,11);
input s_48,s_49;//RE__ALLOW(00,01,10,11);
input s_50,s_51;//RE__ALLOW(00,01,10,11);
input s_52,s_53;//RE__ALLOW(00,01,10,11);
input s_54,s_55;//RE__ALLOW(00,01,10,11);
input s_56,s_57;//RE__ALLOW(00,01,10,11);
input s_58,s_59;//RE__ALLOW(00,01,10,11);
input s_60,s_61;//RE__ALLOW(00,01,10,11);
input s_62,s_63;//RE__ALLOW(00,01,10,11);
input s_64,s_65;//RE__ALLOW(00,01,10,11);
input s_66,s_67;//RE__ALLOW(00,01,10,11);
input s_68,s_69;//RE__ALLOW(00,01,10,11);
input s_70,s_71;//RE__ALLOW(00,01,10,11);
input s_72,s_73;//RE__ALLOW(00,01,10,11);
input s_74,s_75;//RE__ALLOW(00,01,10,11);
input s_76,s_77;//RE__ALLOW(00,01,10,11);
input s_78,s_79;//RE__ALLOW(00,01,10,11);
input s_80,s_81;//RE__ALLOW(00,01,10,11);
input s_82,s_83;//RE__ALLOW(00,01,10,11);
input s_84,s_85;//RE__ALLOW(00,01,10,11);
input s_86,s_87;//RE__ALLOW(00,01,10,11);
input s_88,s_89;//RE__ALLOW(00,01,10,11);
input s_90,s_91;//RE__ALLOW(00,01,10,11);
input s_92,s_93;//RE__ALLOW(00,01,10,11);
input s_94,s_95;//RE__ALLOW(00,01,10,11);
input s_96,s_97;//RE__ALLOW(00,01,10,11);
input s_98,s_99;//RE__ALLOW(00,01,10,11);
input s_100,s_101;//RE__ALLOW(00,01,10,11);
input s_102,s_103;//RE__ALLOW(00,01,10,11);
input s_104,s_105;//RE__ALLOW(00,01,10,11);
input s_106,s_107;//RE__ALLOW(00,01,10,11);
input s_108,s_109;//RE__ALLOW(00,01,10,11);
input s_110,s_111;//RE__ALLOW(00,01,10,11);
input s_112,s_113;//RE__ALLOW(00,01,10,11);
input s_114,s_115;//RE__ALLOW(00,01,10,11);
input s_116,s_117;//RE__ALLOW(00,01,10,11);
input s_118,s_119;//RE__ALLOW(00,01,10,11);
input s_120,s_121;//RE__ALLOW(00,01,10,11);
input s_122,s_123;//RE__ALLOW(00,01,10,11);
input s_124,s_125;//RE__ALLOW(00,01,10,11);
input s_126,s_127;//RE__ALLOW(00,01,10,11);
input s_128,s_129;//RE__ALLOW(00,01,10,11);
input s_130,s_131;//RE__ALLOW(00,01,10,11);
input s_132,s_133;//RE__ALLOW(00,01,10,11);
input s_134,s_135;//RE__ALLOW(00,01,10,11);
input s_136,s_137;//RE__ALLOW(00,01,10,11);
input s_138,s_139;//RE__ALLOW(00,01,10,11);
input s_140,s_141;//RE__ALLOW(00,01,10,11);
input s_142,s_143;//RE__ALLOW(00,01,10,11);
input s_144,s_145;//RE__ALLOW(00,01,10,11);
input s_146,s_147;//RE__ALLOW(00,01,10,11);
input s_148,s_149;//RE__ALLOW(00,01,10,11);
input s_150,s_151;//RE__ALLOW(00,01,10,11);
input s_152,s_153;//RE__ALLOW(00,01,10,11);
input s_154,s_155;//RE__ALLOW(00,01,10,11);
input s_156,s_157;//RE__ALLOW(00,01,10,11);
input s_158,s_159;//RE__ALLOW(00,01,10,11);
input s_160,s_161;//RE__ALLOW(00,01,10,11);
input s_162,s_163;//RE__ALLOW(00,01,10,11);
input s_164,s_165;//RE__ALLOW(00,01,10,11);
input s_166,s_167;//RE__ALLOW(00,01,10,11);
input s_168,s_169;//RE__ALLOW(00,01,10,11);
input s_170,s_171;//RE__ALLOW(00,01,10,11);
input s_172,s_173;//RE__ALLOW(00,01,10,11);
input s_174,s_175;//RE__ALLOW(00,01,10,11);
input s_176,s_177;//RE__ALLOW(00,01,10,11);
input s_178,s_179;//RE__ALLOW(00,01,10,11);
input s_180,s_181;//RE__ALLOW(00,01,10,11);
input s_182,s_183;//RE__ALLOW(00,01,10,11);
input s_184,s_185;//RE__ALLOW(00,01,10,11);
input s_186,s_187;//RE__ALLOW(00,01,10,11);
input s_188,s_189;//RE__ALLOW(00,01,10,11);
input s_190,s_191;//RE__ALLOW(00,01,10,11);
input s_192,s_193;//RE__ALLOW(00,01,10,11);
input s_194,s_195;//RE__ALLOW(00,01,10,11);
input s_196,s_197;//RE__ALLOW(00,01,10,11);
input s_198,s_199;//RE__ALLOW(00,01,10,11);
input s_200,s_201;//RE__ALLOW(00,01,10,11);
input s_202,s_203;//RE__ALLOW(00,01,10,11);
input s_204,s_205;//RE__ALLOW(00,01,10,11);
input s_206,s_207;//RE__ALLOW(00,01,10,11);
input s_208,s_209;//RE__ALLOW(00,01,10,11);
input s_210,s_211;//RE__ALLOW(00,01,10,11);
input s_212,s_213;//RE__ALLOW(00,01,10,11);
input s_214,s_215;//RE__ALLOW(00,01,10,11);
input s_216,s_217;//RE__ALLOW(00,01,10,11);
input s_218,s_219;//RE__ALLOW(00,01,10,11);
input s_220,s_221;//RE__ALLOW(00,01,10,11);
input s_222,s_223;//RE__ALLOW(00,01,10,11);
input s_224,s_225;//RE__ALLOW(00,01,10,11);
input s_226,s_227;//RE__ALLOW(00,01,10,11);
input s_228,s_229;//RE__ALLOW(00,01,10,11);
input s_230,s_231;//RE__ALLOW(00,01,10,11);
input s_232,s_233;//RE__ALLOW(00,01,10,11);
input s_234,s_235;//RE__ALLOW(00,01,10,11);
input s_236,s_237;//RE__ALLOW(00,01,10,11);
input s_238,s_239;//RE__ALLOW(00,01,10,11);
input s_240,s_241;//RE__ALLOW(00,01,10,11);
input s_242,s_243;//RE__ALLOW(00,01,10,11);
input s_244,s_245;//RE__ALLOW(00,01,10,11);
input s_246,s_247;//RE__ALLOW(00,01,10,11);
input s_248,s_249;//RE__ALLOW(00,01,10,11);
input s_250,s_251;//RE__ALLOW(00,01,10,11);
input s_252,s_253;//RE__ALLOW(00,01,10,11);
input s_254,s_255;//RE__ALLOW(00,01,10,11);
input s_256,s_257;//RE__ALLOW(00,01,10,11);
input s_258,s_259;//RE__ALLOW(00,01,10,11);
input s_260,s_261;//RE__ALLOW(00,01,10,11);
input s_262,s_263;//RE__ALLOW(00,01,10,11);
input s_264,s_265;//RE__ALLOW(00,01,10,11);
input s_266,s_267;//RE__ALLOW(00,01,10,11);
input s_268,s_269;//RE__ALLOW(00,01,10,11);
input s_270,s_271;//RE__ALLOW(00,01,10,11);
input s_272,s_273;//RE__ALLOW(00,01,10,11);
input s_274,s_275;//RE__ALLOW(00,01,10,11);
input s_276,s_277;//RE__ALLOW(00,01,10,11);
input s_278,s_279;//RE__ALLOW(00,01,10,11);
input s_280,s_281;//RE__ALLOW(00,01,10,11);
input s_282,s_283;//RE__ALLOW(00,01,10,11);
input s_284,s_285;//RE__ALLOW(00,01,10,11);
input s_286,s_287;//RE__ALLOW(00,01,10,11);
input s_288,s_289;//RE__ALLOW(00,01,10,11);
input s_290,s_291;//RE__ALLOW(00,01,10,11);
input s_292,s_293;//RE__ALLOW(00,01,10,11);
input s_294,s_295;//RE__ALLOW(00,01,10,11);
input s_296,s_297;//RE__ALLOW(00,01,10,11);
input s_298,s_299;//RE__ALLOW(00,01,10,11);
input s_300,s_301;//RE__ALLOW(00,01,10,11);
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;

  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate144inter0, gate144inter1, gate144inter2, gate144inter3, gate144inter4, gate144inter5, gate144inter6, gate144inter7, gate144inter8, gate144inter9, gate144inter10, gate144inter11, gate144inter12, gate295inter0, gate295inter1, gate295inter2, gate295inter3, gate295inter4, gate295inter5, gate295inter6, gate295inter7, gate295inter8, gate295inter9, gate295inter10, gate295inter11, gate295inter12, gate51inter0, gate51inter1, gate51inter2, gate51inter3, gate51inter4, gate51inter5, gate51inter6, gate51inter7, gate51inter8, gate51inter9, gate51inter10, gate51inter11, gate51inter12, gate212inter0, gate212inter1, gate212inter2, gate212inter3, gate212inter4, gate212inter5, gate212inter6, gate212inter7, gate212inter8, gate212inter9, gate212inter10, gate212inter11, gate212inter12, gate25inter0, gate25inter1, gate25inter2, gate25inter3, gate25inter4, gate25inter5, gate25inter6, gate25inter7, gate25inter8, gate25inter9, gate25inter10, gate25inter11, gate25inter12, gate106inter0, gate106inter1, gate106inter2, gate106inter3, gate106inter4, gate106inter5, gate106inter6, gate106inter7, gate106inter8, gate106inter9, gate106inter10, gate106inter11, gate106inter12, gate416inter0, gate416inter1, gate416inter2, gate416inter3, gate416inter4, gate416inter5, gate416inter6, gate416inter7, gate416inter8, gate416inter9, gate416inter10, gate416inter11, gate416inter12, gate99inter0, gate99inter1, gate99inter2, gate99inter3, gate99inter4, gate99inter5, gate99inter6, gate99inter7, gate99inter8, gate99inter9, gate99inter10, gate99inter11, gate99inter12, gate141inter0, gate141inter1, gate141inter2, gate141inter3, gate141inter4, gate141inter5, gate141inter6, gate141inter7, gate141inter8, gate141inter9, gate141inter10, gate141inter11, gate141inter12, gate438inter0, gate438inter1, gate438inter2, gate438inter3, gate438inter4, gate438inter5, gate438inter6, gate438inter7, gate438inter8, gate438inter9, gate438inter10, gate438inter11, gate438inter12, gate415inter0, gate415inter1, gate415inter2, gate415inter3, gate415inter4, gate415inter5, gate415inter6, gate415inter7, gate415inter8, gate415inter9, gate415inter10, gate415inter11, gate415inter12, gate81inter0, gate81inter1, gate81inter2, gate81inter3, gate81inter4, gate81inter5, gate81inter6, gate81inter7, gate81inter8, gate81inter9, gate81inter10, gate81inter11, gate81inter12, gate453inter0, gate453inter1, gate453inter2, gate453inter3, gate453inter4, gate453inter5, gate453inter6, gate453inter7, gate453inter8, gate453inter9, gate453inter10, gate453inter11, gate453inter12, gate421inter0, gate421inter1, gate421inter2, gate421inter3, gate421inter4, gate421inter5, gate421inter6, gate421inter7, gate421inter8, gate421inter9, gate421inter10, gate421inter11, gate421inter12, gate410inter0, gate410inter1, gate410inter2, gate410inter3, gate410inter4, gate410inter5, gate410inter6, gate410inter7, gate410inter8, gate410inter9, gate410inter10, gate410inter11, gate410inter12, gate67inter0, gate67inter1, gate67inter2, gate67inter3, gate67inter4, gate67inter5, gate67inter6, gate67inter7, gate67inter8, gate67inter9, gate67inter10, gate67inter11, gate67inter12, gate496inter0, gate496inter1, gate496inter2, gate496inter3, gate496inter4, gate496inter5, gate496inter6, gate496inter7, gate496inter8, gate496inter9, gate496inter10, gate496inter11, gate496inter12, gate277inter0, gate277inter1, gate277inter2, gate277inter3, gate277inter4, gate277inter5, gate277inter6, gate277inter7, gate277inter8, gate277inter9, gate277inter10, gate277inter11, gate277inter12, gate205inter0, gate205inter1, gate205inter2, gate205inter3, gate205inter4, gate205inter5, gate205inter6, gate205inter7, gate205inter8, gate205inter9, gate205inter10, gate205inter11, gate205inter12, gate50inter0, gate50inter1, gate50inter2, gate50inter3, gate50inter4, gate50inter5, gate50inter6, gate50inter7, gate50inter8, gate50inter9, gate50inter10, gate50inter11, gate50inter12, gate47inter0, gate47inter1, gate47inter2, gate47inter3, gate47inter4, gate47inter5, gate47inter6, gate47inter7, gate47inter8, gate47inter9, gate47inter10, gate47inter11, gate47inter12, gate223inter0, gate223inter1, gate223inter2, gate223inter3, gate223inter4, gate223inter5, gate223inter6, gate223inter7, gate223inter8, gate223inter9, gate223inter10, gate223inter11, gate223inter12, gate189inter0, gate189inter1, gate189inter2, gate189inter3, gate189inter4, gate189inter5, gate189inter6, gate189inter7, gate189inter8, gate189inter9, gate189inter10, gate189inter11, gate189inter12, gate165inter0, gate165inter1, gate165inter2, gate165inter3, gate165inter4, gate165inter5, gate165inter6, gate165inter7, gate165inter8, gate165inter9, gate165inter10, gate165inter11, gate165inter12, gate478inter0, gate478inter1, gate478inter2, gate478inter3, gate478inter4, gate478inter5, gate478inter6, gate478inter7, gate478inter8, gate478inter9, gate478inter10, gate478inter11, gate478inter12, gate221inter0, gate221inter1, gate221inter2, gate221inter3, gate221inter4, gate221inter5, gate221inter6, gate221inter7, gate221inter8, gate221inter9, gate221inter10, gate221inter11, gate221inter12, gate40inter0, gate40inter1, gate40inter2, gate40inter3, gate40inter4, gate40inter5, gate40inter6, gate40inter7, gate40inter8, gate40inter9, gate40inter10, gate40inter11, gate40inter12, gate72inter0, gate72inter1, gate72inter2, gate72inter3, gate72inter4, gate72inter5, gate72inter6, gate72inter7, gate72inter8, gate72inter9, gate72inter10, gate72inter11, gate72inter12, gate149inter0, gate149inter1, gate149inter2, gate149inter3, gate149inter4, gate149inter5, gate149inter6, gate149inter7, gate149inter8, gate149inter9, gate149inter10, gate149inter11, gate149inter12, gate107inter0, gate107inter1, gate107inter2, gate107inter3, gate107inter4, gate107inter5, gate107inter6, gate107inter7, gate107inter8, gate107inter9, gate107inter10, gate107inter11, gate107inter12, gate457inter0, gate457inter1, gate457inter2, gate457inter3, gate457inter4, gate457inter5, gate457inter6, gate457inter7, gate457inter8, gate457inter9, gate457inter10, gate457inter11, gate457inter12, gate430inter0, gate430inter1, gate430inter2, gate430inter3, gate430inter4, gate430inter5, gate430inter6, gate430inter7, gate430inter8, gate430inter9, gate430inter10, gate430inter11, gate430inter12, gate413inter0, gate413inter1, gate413inter2, gate413inter3, gate413inter4, gate413inter5, gate413inter6, gate413inter7, gate413inter8, gate413inter9, gate413inter10, gate413inter11, gate413inter12, gate472inter0, gate472inter1, gate472inter2, gate472inter3, gate472inter4, gate472inter5, gate472inter6, gate472inter7, gate472inter8, gate472inter9, gate472inter10, gate472inter11, gate472inter12, gate456inter0, gate456inter1, gate456inter2, gate456inter3, gate456inter4, gate456inter5, gate456inter6, gate456inter7, gate456inter8, gate456inter9, gate456inter10, gate456inter11, gate456inter12, gate437inter0, gate437inter1, gate437inter2, gate437inter3, gate437inter4, gate437inter5, gate437inter6, gate437inter7, gate437inter8, gate437inter9, gate437inter10, gate437inter11, gate437inter12, gate48inter0, gate48inter1, gate48inter2, gate48inter3, gate48inter4, gate48inter5, gate48inter6, gate48inter7, gate48inter8, gate48inter9, gate48inter10, gate48inter11, gate48inter12, gate119inter0, gate119inter1, gate119inter2, gate119inter3, gate119inter4, gate119inter5, gate119inter6, gate119inter7, gate119inter8, gate119inter9, gate119inter10, gate119inter11, gate119inter12, gate69inter0, gate69inter1, gate69inter2, gate69inter3, gate69inter4, gate69inter5, gate69inter6, gate69inter7, gate69inter8, gate69inter9, gate69inter10, gate69inter11, gate69inter12, gate211inter0, gate211inter1, gate211inter2, gate211inter3, gate211inter4, gate211inter5, gate211inter6, gate211inter7, gate211inter8, gate211inter9, gate211inter10, gate211inter11, gate211inter12, gate414inter0, gate414inter1, gate414inter2, gate414inter3, gate414inter4, gate414inter5, gate414inter6, gate414inter7, gate414inter8, gate414inter9, gate414inter10, gate414inter11, gate414inter12, gate216inter0, gate216inter1, gate216inter2, gate216inter3, gate216inter4, gate216inter5, gate216inter6, gate216inter7, gate216inter8, gate216inter9, gate216inter10, gate216inter11, gate216inter12, gate474inter0, gate474inter1, gate474inter2, gate474inter3, gate474inter4, gate474inter5, gate474inter6, gate474inter7, gate474inter8, gate474inter9, gate474inter10, gate474inter11, gate474inter12, gate62inter0, gate62inter1, gate62inter2, gate62inter3, gate62inter4, gate62inter5, gate62inter6, gate62inter7, gate62inter8, gate62inter9, gate62inter10, gate62inter11, gate62inter12, gate268inter0, gate268inter1, gate268inter2, gate268inter3, gate268inter4, gate268inter5, gate268inter6, gate268inter7, gate268inter8, gate268inter9, gate268inter10, gate268inter11, gate268inter12, gate466inter0, gate466inter1, gate466inter2, gate466inter3, gate466inter4, gate466inter5, gate466inter6, gate466inter7, gate466inter8, gate466inter9, gate466inter10, gate466inter11, gate466inter12, gate213inter0, gate213inter1, gate213inter2, gate213inter3, gate213inter4, gate213inter5, gate213inter6, gate213inter7, gate213inter8, gate213inter9, gate213inter10, gate213inter11, gate213inter12, gate483inter0, gate483inter1, gate483inter2, gate483inter3, gate483inter4, gate483inter5, gate483inter6, gate483inter7, gate483inter8, gate483inter9, gate483inter10, gate483inter11, gate483inter12, gate18inter0, gate18inter1, gate18inter2, gate18inter3, gate18inter4, gate18inter5, gate18inter6, gate18inter7, gate18inter8, gate18inter9, gate18inter10, gate18inter11, gate18inter12, gate41inter0, gate41inter1, gate41inter2, gate41inter3, gate41inter4, gate41inter5, gate41inter6, gate41inter7, gate41inter8, gate41inter9, gate41inter10, gate41inter11, gate41inter12, gate391inter0, gate391inter1, gate391inter2, gate391inter3, gate391inter4, gate391inter5, gate391inter6, gate391inter7, gate391inter8, gate391inter9, gate391inter10, gate391inter11, gate391inter12, gate278inter0, gate278inter1, gate278inter2, gate278inter3, gate278inter4, gate278inter5, gate278inter6, gate278inter7, gate278inter8, gate278inter9, gate278inter10, gate278inter11, gate278inter12, gate462inter0, gate462inter1, gate462inter2, gate462inter3, gate462inter4, gate462inter5, gate462inter6, gate462inter7, gate462inter8, gate462inter9, gate462inter10, gate462inter11, gate462inter12, gate53inter0, gate53inter1, gate53inter2, gate53inter3, gate53inter4, gate53inter5, gate53inter6, gate53inter7, gate53inter8, gate53inter9, gate53inter10, gate53inter11, gate53inter12, gate206inter0, gate206inter1, gate206inter2, gate206inter3, gate206inter4, gate206inter5, gate206inter6, gate206inter7, gate206inter8, gate206inter9, gate206inter10, gate206inter11, gate206inter12, gate282inter0, gate282inter1, gate282inter2, gate282inter3, gate282inter4, gate282inter5, gate282inter6, gate282inter7, gate282inter8, gate282inter9, gate282inter10, gate282inter11, gate282inter12, gate61inter0, gate61inter1, gate61inter2, gate61inter3, gate61inter4, gate61inter5, gate61inter6, gate61inter7, gate61inter8, gate61inter9, gate61inter10, gate61inter11, gate61inter12, gate503inter0, gate503inter1, gate503inter2, gate503inter3, gate503inter4, gate503inter5, gate503inter6, gate503inter7, gate503inter8, gate503inter9, gate503inter10, gate503inter11, gate503inter12, gate417inter0, gate417inter1, gate417inter2, gate417inter3, gate417inter4, gate417inter5, gate417inter6, gate417inter7, gate417inter8, gate417inter9, gate417inter10, gate417inter11, gate417inter12, gate271inter0, gate271inter1, gate271inter2, gate271inter3, gate271inter4, gate271inter5, gate271inter6, gate271inter7, gate271inter8, gate271inter9, gate271inter10, gate271inter11, gate271inter12, gate52inter0, gate52inter1, gate52inter2, gate52inter3, gate52inter4, gate52inter5, gate52inter6, gate52inter7, gate52inter8, gate52inter9, gate52inter10, gate52inter11, gate52inter12, gate252inter0, gate252inter1, gate252inter2, gate252inter3, gate252inter4, gate252inter5, gate252inter6, gate252inter7, gate252inter8, gate252inter9, gate252inter10, gate252inter11, gate252inter12, gate257inter0, gate257inter1, gate257inter2, gate257inter3, gate257inter4, gate257inter5, gate257inter6, gate257inter7, gate257inter8, gate257inter9, gate257inter10, gate257inter11, gate257inter12, gate234inter0, gate234inter1, gate234inter2, gate234inter3, gate234inter4, gate234inter5, gate234inter6, gate234inter7, gate234inter8, gate234inter9, gate234inter10, gate234inter11, gate234inter12, gate393inter0, gate393inter1, gate393inter2, gate393inter3, gate393inter4, gate393inter5, gate393inter6, gate393inter7, gate393inter8, gate393inter9, gate393inter10, gate393inter11, gate393inter12, gate442inter0, gate442inter1, gate442inter2, gate442inter3, gate442inter4, gate442inter5, gate442inter6, gate442inter7, gate442inter8, gate442inter9, gate442inter10, gate442inter11, gate442inter12, gate435inter0, gate435inter1, gate435inter2, gate435inter3, gate435inter4, gate435inter5, gate435inter6, gate435inter7, gate435inter8, gate435inter9, gate435inter10, gate435inter11, gate435inter12, gate481inter0, gate481inter1, gate481inter2, gate481inter3, gate481inter4, gate481inter5, gate481inter6, gate481inter7, gate481inter8, gate481inter9, gate481inter10, gate481inter11, gate481inter12, gate392inter0, gate392inter1, gate392inter2, gate392inter3, gate392inter4, gate392inter5, gate392inter6, gate392inter7, gate392inter8, gate392inter9, gate392inter10, gate392inter11, gate392inter12, gate27inter0, gate27inter1, gate27inter2, gate27inter3, gate27inter4, gate27inter5, gate27inter6, gate27inter7, gate27inter8, gate27inter9, gate27inter10, gate27inter11, gate27inter12, gate288inter0, gate288inter1, gate288inter2, gate288inter3, gate288inter4, gate288inter5, gate288inter6, gate288inter7, gate288inter8, gate288inter9, gate288inter10, gate288inter11, gate288inter12, gate464inter0, gate464inter1, gate464inter2, gate464inter3, gate464inter4, gate464inter5, gate464inter6, gate464inter7, gate464inter8, gate464inter9, gate464inter10, gate464inter11, gate464inter12, gate84inter0, gate84inter1, gate84inter2, gate84inter3, gate84inter4, gate84inter5, gate84inter6, gate84inter7, gate84inter8, gate84inter9, gate84inter10, gate84inter11, gate84inter12, gate394inter0, gate394inter1, gate394inter2, gate394inter3, gate394inter4, gate394inter5, gate394inter6, gate394inter7, gate394inter8, gate394inter9, gate394inter10, gate394inter11, gate394inter12, gate43inter0, gate43inter1, gate43inter2, gate43inter3, gate43inter4, gate43inter5, gate43inter6, gate43inter7, gate43inter8, gate43inter9, gate43inter10, gate43inter11, gate43inter12, gate260inter0, gate260inter1, gate260inter2, gate260inter3, gate260inter4, gate260inter5, gate260inter6, gate260inter7, gate260inter8, gate260inter9, gate260inter10, gate260inter11, gate260inter12, gate485inter0, gate485inter1, gate485inter2, gate485inter3, gate485inter4, gate485inter5, gate485inter6, gate485inter7, gate485inter8, gate485inter9, gate485inter10, gate485inter11, gate485inter12, gate388inter0, gate388inter1, gate388inter2, gate388inter3, gate388inter4, gate388inter5, gate388inter6, gate388inter7, gate388inter8, gate388inter9, gate388inter10, gate388inter11, gate388inter12, gate178inter0, gate178inter1, gate178inter2, gate178inter3, gate178inter4, gate178inter5, gate178inter6, gate178inter7, gate178inter8, gate178inter9, gate178inter10, gate178inter11, gate178inter12, gate181inter0, gate181inter1, gate181inter2, gate181inter3, gate181inter4, gate181inter5, gate181inter6, gate181inter7, gate181inter8, gate181inter9, gate181inter10, gate181inter11, gate181inter12, gate400inter0, gate400inter1, gate400inter2, gate400inter3, gate400inter4, gate400inter5, gate400inter6, gate400inter7, gate400inter8, gate400inter9, gate400inter10, gate400inter11, gate400inter12, gate251inter0, gate251inter1, gate251inter2, gate251inter3, gate251inter4, gate251inter5, gate251inter6, gate251inter7, gate251inter8, gate251inter9, gate251inter10, gate251inter11, gate251inter12, gate255inter0, gate255inter1, gate255inter2, gate255inter3, gate255inter4, gate255inter5, gate255inter6, gate255inter7, gate255inter8, gate255inter9, gate255inter10, gate255inter11, gate255inter12, gate158inter0, gate158inter1, gate158inter2, gate158inter3, gate158inter4, gate158inter5, gate158inter6, gate158inter7, gate158inter8, gate158inter9, gate158inter10, gate158inter11, gate158inter12, gate270inter0, gate270inter1, gate270inter2, gate270inter3, gate270inter4, gate270inter5, gate270inter6, gate270inter7, gate270inter8, gate270inter9, gate270inter10, gate270inter11, gate270inter12, gate73inter0, gate73inter1, gate73inter2, gate73inter3, gate73inter4, gate73inter5, gate73inter6, gate73inter7, gate73inter8, gate73inter9, gate73inter10, gate73inter11, gate73inter12, gate511inter0, gate511inter1, gate511inter2, gate511inter3, gate511inter4, gate511inter5, gate511inter6, gate511inter7, gate511inter8, gate511inter9, gate511inter10, gate511inter11, gate511inter12, gate74inter0, gate74inter1, gate74inter2, gate74inter3, gate74inter4, gate74inter5, gate74inter6, gate74inter7, gate74inter8, gate74inter9, gate74inter10, gate74inter11, gate74inter12, gate64inter0, gate64inter1, gate64inter2, gate64inter3, gate64inter4, gate64inter5, gate64inter6, gate64inter7, gate64inter8, gate64inter9, gate64inter10, gate64inter11, gate64inter12, gate192inter0, gate192inter1, gate192inter2, gate192inter3, gate192inter4, gate192inter5, gate192inter6, gate192inter7, gate192inter8, gate192inter9, gate192inter10, gate192inter11, gate192inter12, gate480inter0, gate480inter1, gate480inter2, gate480inter3, gate480inter4, gate480inter5, gate480inter6, gate480inter7, gate480inter8, gate480inter9, gate480inter10, gate480inter11, gate480inter12, gate228inter0, gate228inter1, gate228inter2, gate228inter3, gate228inter4, gate228inter5, gate228inter6, gate228inter7, gate228inter8, gate228inter9, gate228inter10, gate228inter11, gate228inter12, gate280inter0, gate280inter1, gate280inter2, gate280inter3, gate280inter4, gate280inter5, gate280inter6, gate280inter7, gate280inter8, gate280inter9, gate280inter10, gate280inter11, gate280inter12, gate155inter0, gate155inter1, gate155inter2, gate155inter3, gate155inter4, gate155inter5, gate155inter6, gate155inter7, gate155inter8, gate155inter9, gate155inter10, gate155inter11, gate155inter12, gate194inter0, gate194inter1, gate194inter2, gate194inter3, gate194inter4, gate194inter5, gate194inter6, gate194inter7, gate194inter8, gate194inter9, gate194inter10, gate194inter11, gate194inter12, gate115inter0, gate115inter1, gate115inter2, gate115inter3, gate115inter4, gate115inter5, gate115inter6, gate115inter7, gate115inter8, gate115inter9, gate115inter10, gate115inter11, gate115inter12, gate296inter0, gate296inter1, gate296inter2, gate296inter3, gate296inter4, gate296inter5, gate296inter6, gate296inter7, gate296inter8, gate296inter9, gate296inter10, gate296inter11, gate296inter12, gate88inter0, gate88inter1, gate88inter2, gate88inter3, gate88inter4, gate88inter5, gate88inter6, gate88inter7, gate88inter8, gate88inter9, gate88inter10, gate88inter11, gate88inter12, gate128inter0, gate128inter1, gate128inter2, gate128inter3, gate128inter4, gate128inter5, gate128inter6, gate128inter7, gate128inter8, gate128inter9, gate128inter10, gate128inter11, gate128inter12, gate157inter0, gate157inter1, gate157inter2, gate157inter3, gate157inter4, gate157inter5, gate157inter6, gate157inter7, gate157inter8, gate157inter9, gate157inter10, gate157inter11, gate157inter12, gate227inter0, gate227inter1, gate227inter2, gate227inter3, gate227inter4, gate227inter5, gate227inter6, gate227inter7, gate227inter8, gate227inter9, gate227inter10, gate227inter11, gate227inter12, gate461inter0, gate461inter1, gate461inter2, gate461inter3, gate461inter4, gate461inter5, gate461inter6, gate461inter7, gate461inter8, gate461inter9, gate461inter10, gate461inter11, gate461inter12, gate443inter0, gate443inter1, gate443inter2, gate443inter3, gate443inter4, gate443inter5, gate443inter6, gate443inter7, gate443inter8, gate443inter9, gate443inter10, gate443inter11, gate443inter12, gate126inter0, gate126inter1, gate126inter2, gate126inter3, gate126inter4, gate126inter5, gate126inter6, gate126inter7, gate126inter8, gate126inter9, gate126inter10, gate126inter11, gate126inter12, gate408inter0, gate408inter1, gate408inter2, gate408inter3, gate408inter4, gate408inter5, gate408inter6, gate408inter7, gate408inter8, gate408inter9, gate408inter10, gate408inter11, gate408inter12, gate407inter0, gate407inter1, gate407inter2, gate407inter3, gate407inter4, gate407inter5, gate407inter6, gate407inter7, gate407inter8, gate407inter9, gate407inter10, gate407inter11, gate407inter12, gate92inter0, gate92inter1, gate92inter2, gate92inter3, gate92inter4, gate92inter5, gate92inter6, gate92inter7, gate92inter8, gate92inter9, gate92inter10, gate92inter11, gate92inter12, gate293inter0, gate293inter1, gate293inter2, gate293inter3, gate293inter4, gate293inter5, gate293inter6, gate293inter7, gate293inter8, gate293inter9, gate293inter10, gate293inter11, gate293inter12, gate168inter0, gate168inter1, gate168inter2, gate168inter3, gate168inter4, gate168inter5, gate168inter6, gate168inter7, gate168inter8, gate168inter9, gate168inter10, gate168inter11, gate168inter12, gate446inter0, gate446inter1, gate446inter2, gate446inter3, gate446inter4, gate446inter5, gate446inter6, gate446inter7, gate446inter8, gate446inter9, gate446inter10, gate446inter11, gate446inter12, gate397inter0, gate397inter1, gate397inter2, gate397inter3, gate397inter4, gate397inter5, gate397inter6, gate397inter7, gate397inter8, gate397inter9, gate397inter10, gate397inter11, gate397inter12, gate98inter0, gate98inter1, gate98inter2, gate98inter3, gate98inter4, gate98inter5, gate98inter6, gate98inter7, gate98inter8, gate98inter9, gate98inter10, gate98inter11, gate98inter12, gate36inter0, gate36inter1, gate36inter2, gate36inter3, gate36inter4, gate36inter5, gate36inter6, gate36inter7, gate36inter8, gate36inter9, gate36inter10, gate36inter11, gate36inter12, gate188inter0, gate188inter1, gate188inter2, gate188inter3, gate188inter4, gate188inter5, gate188inter6, gate188inter7, gate188inter8, gate188inter9, gate188inter10, gate188inter11, gate188inter12, gate186inter0, gate186inter1, gate186inter2, gate186inter3, gate186inter4, gate186inter5, gate186inter6, gate186inter7, gate186inter8, gate186inter9, gate186inter10, gate186inter11, gate186inter12, gate22inter0, gate22inter1, gate22inter2, gate22inter3, gate22inter4, gate22inter5, gate22inter6, gate22inter7, gate22inter8, gate22inter9, gate22inter10, gate22inter11, gate22inter12, gate85inter0, gate85inter1, gate85inter2, gate85inter3, gate85inter4, gate85inter5, gate85inter6, gate85inter7, gate85inter8, gate85inter9, gate85inter10, gate85inter11, gate85inter12, gate512inter0, gate512inter1, gate512inter2, gate512inter3, gate512inter4, gate512inter5, gate512inter6, gate512inter7, gate512inter8, gate512inter9, gate512inter10, gate512inter11, gate512inter12, gate184inter0, gate184inter1, gate184inter2, gate184inter3, gate184inter4, gate184inter5, gate184inter6, gate184inter7, gate184inter8, gate184inter9, gate184inter10, gate184inter11, gate184inter12, gate195inter0, gate195inter1, gate195inter2, gate195inter3, gate195inter4, gate195inter5, gate195inter6, gate195inter7, gate195inter8, gate195inter9, gate195inter10, gate195inter11, gate195inter12, gate172inter0, gate172inter1, gate172inter2, gate172inter3, gate172inter4, gate172inter5, gate172inter6, gate172inter7, gate172inter8, gate172inter9, gate172inter10, gate172inter11, gate172inter12, gate123inter0, gate123inter1, gate123inter2, gate123inter3, gate123inter4, gate123inter5, gate123inter6, gate123inter7, gate123inter8, gate123inter9, gate123inter10, gate123inter11, gate123inter12, gate20inter0, gate20inter1, gate20inter2, gate20inter3, gate20inter4, gate20inter5, gate20inter6, gate20inter7, gate20inter8, gate20inter9, gate20inter10, gate20inter11, gate20inter12, gate484inter0, gate484inter1, gate484inter2, gate484inter3, gate484inter4, gate484inter5, gate484inter6, gate484inter7, gate484inter8, gate484inter9, gate484inter10, gate484inter11, gate484inter12, gate292inter0, gate292inter1, gate292inter2, gate292inter3, gate292inter4, gate292inter5, gate292inter6, gate292inter7, gate292inter8, gate292inter9, gate292inter10, gate292inter11, gate292inter12, gate265inter0, gate265inter1, gate265inter2, gate265inter3, gate265inter4, gate265inter5, gate265inter6, gate265inter7, gate265inter8, gate265inter9, gate265inter10, gate265inter11, gate265inter12, gate49inter0, gate49inter1, gate49inter2, gate49inter3, gate49inter4, gate49inter5, gate49inter6, gate49inter7, gate49inter8, gate49inter9, gate49inter10, gate49inter11, gate49inter12, gate439inter0, gate439inter1, gate439inter2, gate439inter3, gate439inter4, gate439inter5, gate439inter6, gate439inter7, gate439inter8, gate439inter9, gate439inter10, gate439inter11, gate439inter12, gate506inter0, gate506inter1, gate506inter2, gate506inter3, gate506inter4, gate506inter5, gate506inter6, gate506inter7, gate506inter8, gate506inter9, gate506inter10, gate506inter11, gate506inter12, gate44inter0, gate44inter1, gate44inter2, gate44inter3, gate44inter4, gate44inter5, gate44inter6, gate44inter7, gate44inter8, gate44inter9, gate44inter10, gate44inter11, gate44inter12, gate54inter0, gate54inter1, gate54inter2, gate54inter3, gate54inter4, gate54inter5, gate54inter6, gate54inter7, gate54inter8, gate54inter9, gate54inter10, gate54inter11, gate54inter12, gate56inter0, gate56inter1, gate56inter2, gate56inter3, gate56inter4, gate56inter5, gate56inter6, gate56inter7, gate56inter8, gate56inter9, gate56inter10, gate56inter11, gate56inter12, gate289inter0, gate289inter1, gate289inter2, gate289inter3, gate289inter4, gate289inter5, gate289inter6, gate289inter7, gate289inter8, gate289inter9, gate289inter10, gate289inter11, gate289inter12, gate493inter0, gate493inter1, gate493inter2, gate493inter3, gate493inter4, gate493inter5, gate493inter6, gate493inter7, gate493inter8, gate493inter9, gate493inter10, gate493inter11, gate493inter12, gate101inter0, gate101inter1, gate101inter2, gate101inter3, gate101inter4, gate101inter5, gate101inter6, gate101inter7, gate101inter8, gate101inter9, gate101inter10, gate101inter11, gate101inter12, gate140inter0, gate140inter1, gate140inter2, gate140inter3, gate140inter4, gate140inter5, gate140inter6, gate140inter7, gate140inter8, gate140inter9, gate140inter10, gate140inter11, gate140inter12, gate151inter0, gate151inter1, gate151inter2, gate151inter3, gate151inter4, gate151inter5, gate151inter6, gate151inter7, gate151inter8, gate151inter9, gate151inter10, gate151inter11, gate151inter12, gate447inter0, gate447inter1, gate447inter2, gate447inter3, gate447inter4, gate447inter5, gate447inter6, gate447inter7, gate447inter8, gate447inter9, gate447inter10, gate447inter11, gate447inter12, gate507inter0, gate507inter1, gate507inter2, gate507inter3, gate507inter4, gate507inter5, gate507inter6, gate507inter7, gate507inter8, gate507inter9, gate507inter10, gate507inter11, gate507inter12, gate276inter0, gate276inter1, gate276inter2, gate276inter3, gate276inter4, gate276inter5, gate276inter6, gate276inter7, gate276inter8, gate276inter9, gate276inter10, gate276inter11, gate276inter12, gate196inter0, gate196inter1, gate196inter2, gate196inter3, gate196inter4, gate196inter5, gate196inter6, gate196inter7, gate196inter8, gate196inter9, gate196inter10, gate196inter11, gate196inter12, gate387inter0, gate387inter1, gate387inter2, gate387inter3, gate387inter4, gate387inter5, gate387inter6, gate387inter7, gate387inter8, gate387inter9, gate387inter10, gate387inter11, gate387inter12, gate102inter0, gate102inter1, gate102inter2, gate102inter3, gate102inter4, gate102inter5, gate102inter6, gate102inter7, gate102inter8, gate102inter9, gate102inter10, gate102inter11, gate102inter12, gate491inter0, gate491inter1, gate491inter2, gate491inter3, gate491inter4, gate491inter5, gate491inter6, gate491inter7, gate491inter8, gate491inter9, gate491inter10, gate491inter11, gate491inter12, gate495inter0, gate495inter1, gate495inter2, gate495inter3, gate495inter4, gate495inter5, gate495inter6, gate495inter7, gate495inter8, gate495inter9, gate495inter10, gate495inter11, gate495inter12, gate169inter0, gate169inter1, gate169inter2, gate169inter3, gate169inter4, gate169inter5, gate169inter6, gate169inter7, gate169inter8, gate169inter9, gate169inter10, gate169inter11, gate169inter12, gate55inter0, gate55inter1, gate55inter2, gate55inter3, gate55inter4, gate55inter5, gate55inter6, gate55inter7, gate55inter8, gate55inter9, gate55inter10, gate55inter11, gate55inter12, gate32inter0, gate32inter1, gate32inter2, gate32inter3, gate32inter4, gate32inter5, gate32inter6, gate32inter7, gate32inter8, gate32inter9, gate32inter10, gate32inter11, gate32inter12, gate285inter0, gate285inter1, gate285inter2, gate285inter3, gate285inter4, gate285inter5, gate285inter6, gate285inter7, gate285inter8, gate285inter9, gate285inter10, gate285inter11, gate285inter12, gate139inter0, gate139inter1, gate139inter2, gate139inter3, gate139inter4, gate139inter5, gate139inter6, gate139inter7, gate139inter8, gate139inter9, gate139inter10, gate139inter11, gate139inter12, gate87inter0, gate87inter1, gate87inter2, gate87inter3, gate87inter4, gate87inter5, gate87inter6, gate87inter7, gate87inter8, gate87inter9, gate87inter10, gate87inter11, gate87inter12;



and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );
nand2 gate9( .a(G1), .b(G2), .O(G266) );
nand2 gate10( .a(G3), .b(G4), .O(G269) );
nand2 gate11( .a(G5), .b(G6), .O(G272) );
nand2 gate12( .a(G7), .b(G8), .O(G275) );
nand2 gate13( .a(G9), .b(G10), .O(G278) );
nand2 gate14( .a(G11), .b(G12), .O(G281) );
nand2 gate15( .a(G13), .b(G14), .O(G284) );
nand2 gate16( .a(G15), .b(G16), .O(G287) );
nand2 gate17( .a(G17), .b(G18), .O(G290) );

  xor2  gate1219(.a(G20), .b(G19), .O(gate18inter0));
  nand2 gate1220(.a(gate18inter0), .b(s_96), .O(gate18inter1));
  and2  gate1221(.a(G20), .b(G19), .O(gate18inter2));
  inv1  gate1222(.a(s_96), .O(gate18inter3));
  inv1  gate1223(.a(s_97), .O(gate18inter4));
  nand2 gate1224(.a(gate18inter4), .b(gate18inter3), .O(gate18inter5));
  nor2  gate1225(.a(gate18inter5), .b(gate18inter2), .O(gate18inter6));
  inv1  gate1226(.a(G19), .O(gate18inter7));
  inv1  gate1227(.a(G20), .O(gate18inter8));
  nand2 gate1228(.a(gate18inter8), .b(gate18inter7), .O(gate18inter9));
  nand2 gate1229(.a(s_97), .b(gate18inter3), .O(gate18inter10));
  nor2  gate1230(.a(gate18inter10), .b(gate18inter9), .O(gate18inter11));
  nor2  gate1231(.a(gate18inter11), .b(gate18inter6), .O(gate18inter12));
  nand2 gate1232(.a(gate18inter12), .b(gate18inter1), .O(G293));
nand2 gate19( .a(G21), .b(G22), .O(G296) );

  xor2  gate2255(.a(G24), .b(G23), .O(gate20inter0));
  nand2 gate2256(.a(gate20inter0), .b(s_244), .O(gate20inter1));
  and2  gate2257(.a(G24), .b(G23), .O(gate20inter2));
  inv1  gate2258(.a(s_244), .O(gate20inter3));
  inv1  gate2259(.a(s_245), .O(gate20inter4));
  nand2 gate2260(.a(gate20inter4), .b(gate20inter3), .O(gate20inter5));
  nor2  gate2261(.a(gate20inter5), .b(gate20inter2), .O(gate20inter6));
  inv1  gate2262(.a(G23), .O(gate20inter7));
  inv1  gate2263(.a(G24), .O(gate20inter8));
  nand2 gate2264(.a(gate20inter8), .b(gate20inter7), .O(gate20inter9));
  nand2 gate2265(.a(s_245), .b(gate20inter3), .O(gate20inter10));
  nor2  gate2266(.a(gate20inter10), .b(gate20inter9), .O(gate20inter11));
  nor2  gate2267(.a(gate20inter11), .b(gate20inter6), .O(gate20inter12));
  nand2 gate2268(.a(gate20inter12), .b(gate20inter1), .O(G299));
nand2 gate21( .a(G25), .b(G26), .O(G302) );

  xor2  gate2157(.a(G28), .b(G27), .O(gate22inter0));
  nand2 gate2158(.a(gate22inter0), .b(s_230), .O(gate22inter1));
  and2  gate2159(.a(G28), .b(G27), .O(gate22inter2));
  inv1  gate2160(.a(s_230), .O(gate22inter3));
  inv1  gate2161(.a(s_231), .O(gate22inter4));
  nand2 gate2162(.a(gate22inter4), .b(gate22inter3), .O(gate22inter5));
  nor2  gate2163(.a(gate22inter5), .b(gate22inter2), .O(gate22inter6));
  inv1  gate2164(.a(G27), .O(gate22inter7));
  inv1  gate2165(.a(G28), .O(gate22inter8));
  nand2 gate2166(.a(gate22inter8), .b(gate22inter7), .O(gate22inter9));
  nand2 gate2167(.a(s_231), .b(gate22inter3), .O(gate22inter10));
  nor2  gate2168(.a(gate22inter10), .b(gate22inter9), .O(gate22inter11));
  nor2  gate2169(.a(gate22inter11), .b(gate22inter6), .O(gate22inter12));
  nand2 gate2170(.a(gate22inter12), .b(gate22inter1), .O(G305));
nand2 gate23( .a(G29), .b(G30), .O(G308) );
nand2 gate24( .a(G31), .b(G32), .O(G311) );

  xor2  gate603(.a(G5), .b(G1), .O(gate25inter0));
  nand2 gate604(.a(gate25inter0), .b(s_8), .O(gate25inter1));
  and2  gate605(.a(G5), .b(G1), .O(gate25inter2));
  inv1  gate606(.a(s_8), .O(gate25inter3));
  inv1  gate607(.a(s_9), .O(gate25inter4));
  nand2 gate608(.a(gate25inter4), .b(gate25inter3), .O(gate25inter5));
  nor2  gate609(.a(gate25inter5), .b(gate25inter2), .O(gate25inter6));
  inv1  gate610(.a(G1), .O(gate25inter7));
  inv1  gate611(.a(G5), .O(gate25inter8));
  nand2 gate612(.a(gate25inter8), .b(gate25inter7), .O(gate25inter9));
  nand2 gate613(.a(s_9), .b(gate25inter3), .O(gate25inter10));
  nor2  gate614(.a(gate25inter10), .b(gate25inter9), .O(gate25inter11));
  nor2  gate615(.a(gate25inter11), .b(gate25inter6), .O(gate25inter12));
  nand2 gate616(.a(gate25inter12), .b(gate25inter1), .O(G314));
nand2 gate26( .a(G9), .b(G13), .O(G317) );

  xor2  gate1513(.a(G6), .b(G2), .O(gate27inter0));
  nand2 gate1514(.a(gate27inter0), .b(s_138), .O(gate27inter1));
  and2  gate1515(.a(G6), .b(G2), .O(gate27inter2));
  inv1  gate1516(.a(s_138), .O(gate27inter3));
  inv1  gate1517(.a(s_139), .O(gate27inter4));
  nand2 gate1518(.a(gate27inter4), .b(gate27inter3), .O(gate27inter5));
  nor2  gate1519(.a(gate27inter5), .b(gate27inter2), .O(gate27inter6));
  inv1  gate1520(.a(G2), .O(gate27inter7));
  inv1  gate1521(.a(G6), .O(gate27inter8));
  nand2 gate1522(.a(gate27inter8), .b(gate27inter7), .O(gate27inter9));
  nand2 gate1523(.a(s_139), .b(gate27inter3), .O(gate27inter10));
  nor2  gate1524(.a(gate27inter10), .b(gate27inter9), .O(gate27inter11));
  nor2  gate1525(.a(gate27inter11), .b(gate27inter6), .O(gate27inter12));
  nand2 gate1526(.a(gate27inter12), .b(gate27inter1), .O(G320));
nand2 gate28( .a(G10), .b(G14), .O(G323) );
nand2 gate29( .a(G3), .b(G7), .O(G326) );
nand2 gate30( .a(G11), .b(G15), .O(G329) );
nand2 gate31( .a(G4), .b(G8), .O(G332) );

  xor2  gate2605(.a(G16), .b(G12), .O(gate32inter0));
  nand2 gate2606(.a(gate32inter0), .b(s_294), .O(gate32inter1));
  and2  gate2607(.a(G16), .b(G12), .O(gate32inter2));
  inv1  gate2608(.a(s_294), .O(gate32inter3));
  inv1  gate2609(.a(s_295), .O(gate32inter4));
  nand2 gate2610(.a(gate32inter4), .b(gate32inter3), .O(gate32inter5));
  nor2  gate2611(.a(gate32inter5), .b(gate32inter2), .O(gate32inter6));
  inv1  gate2612(.a(G12), .O(gate32inter7));
  inv1  gate2613(.a(G16), .O(gate32inter8));
  nand2 gate2614(.a(gate32inter8), .b(gate32inter7), .O(gate32inter9));
  nand2 gate2615(.a(s_295), .b(gate32inter3), .O(gate32inter10));
  nor2  gate2616(.a(gate32inter10), .b(gate32inter9), .O(gate32inter11));
  nor2  gate2617(.a(gate32inter11), .b(gate32inter6), .O(gate32inter12));
  nand2 gate2618(.a(gate32inter12), .b(gate32inter1), .O(G335));
nand2 gate33( .a(G17), .b(G21), .O(G338) );
nand2 gate34( .a(G25), .b(G29), .O(G341) );
nand2 gate35( .a(G18), .b(G22), .O(G344) );

  xor2  gate2115(.a(G30), .b(G26), .O(gate36inter0));
  nand2 gate2116(.a(gate36inter0), .b(s_224), .O(gate36inter1));
  and2  gate2117(.a(G30), .b(G26), .O(gate36inter2));
  inv1  gate2118(.a(s_224), .O(gate36inter3));
  inv1  gate2119(.a(s_225), .O(gate36inter4));
  nand2 gate2120(.a(gate36inter4), .b(gate36inter3), .O(gate36inter5));
  nor2  gate2121(.a(gate36inter5), .b(gate36inter2), .O(gate36inter6));
  inv1  gate2122(.a(G26), .O(gate36inter7));
  inv1  gate2123(.a(G30), .O(gate36inter8));
  nand2 gate2124(.a(gate36inter8), .b(gate36inter7), .O(gate36inter9));
  nand2 gate2125(.a(s_225), .b(gate36inter3), .O(gate36inter10));
  nor2  gate2126(.a(gate36inter10), .b(gate36inter9), .O(gate36inter11));
  nor2  gate2127(.a(gate36inter11), .b(gate36inter6), .O(gate36inter12));
  nand2 gate2128(.a(gate36inter12), .b(gate36inter1), .O(G347));
nand2 gate37( .a(G19), .b(G23), .O(G350) );
nand2 gate38( .a(G27), .b(G31), .O(G353) );
nand2 gate39( .a(G20), .b(G24), .O(G356) );

  xor2  gate911(.a(G32), .b(G28), .O(gate40inter0));
  nand2 gate912(.a(gate40inter0), .b(s_52), .O(gate40inter1));
  and2  gate913(.a(G32), .b(G28), .O(gate40inter2));
  inv1  gate914(.a(s_52), .O(gate40inter3));
  inv1  gate915(.a(s_53), .O(gate40inter4));
  nand2 gate916(.a(gate40inter4), .b(gate40inter3), .O(gate40inter5));
  nor2  gate917(.a(gate40inter5), .b(gate40inter2), .O(gate40inter6));
  inv1  gate918(.a(G28), .O(gate40inter7));
  inv1  gate919(.a(G32), .O(gate40inter8));
  nand2 gate920(.a(gate40inter8), .b(gate40inter7), .O(gate40inter9));
  nand2 gate921(.a(s_53), .b(gate40inter3), .O(gate40inter10));
  nor2  gate922(.a(gate40inter10), .b(gate40inter9), .O(gate40inter11));
  nor2  gate923(.a(gate40inter11), .b(gate40inter6), .O(gate40inter12));
  nand2 gate924(.a(gate40inter12), .b(gate40inter1), .O(G359));

  xor2  gate1233(.a(G266), .b(G1), .O(gate41inter0));
  nand2 gate1234(.a(gate41inter0), .b(s_98), .O(gate41inter1));
  and2  gate1235(.a(G266), .b(G1), .O(gate41inter2));
  inv1  gate1236(.a(s_98), .O(gate41inter3));
  inv1  gate1237(.a(s_99), .O(gate41inter4));
  nand2 gate1238(.a(gate41inter4), .b(gate41inter3), .O(gate41inter5));
  nor2  gate1239(.a(gate41inter5), .b(gate41inter2), .O(gate41inter6));
  inv1  gate1240(.a(G1), .O(gate41inter7));
  inv1  gate1241(.a(G266), .O(gate41inter8));
  nand2 gate1242(.a(gate41inter8), .b(gate41inter7), .O(gate41inter9));
  nand2 gate1243(.a(s_99), .b(gate41inter3), .O(gate41inter10));
  nor2  gate1244(.a(gate41inter10), .b(gate41inter9), .O(gate41inter11));
  nor2  gate1245(.a(gate41inter11), .b(gate41inter6), .O(gate41inter12));
  nand2 gate1246(.a(gate41inter12), .b(gate41inter1), .O(G362));
nand2 gate42( .a(G2), .b(G266), .O(G363) );

  xor2  gate1583(.a(G269), .b(G3), .O(gate43inter0));
  nand2 gate1584(.a(gate43inter0), .b(s_148), .O(gate43inter1));
  and2  gate1585(.a(G269), .b(G3), .O(gate43inter2));
  inv1  gate1586(.a(s_148), .O(gate43inter3));
  inv1  gate1587(.a(s_149), .O(gate43inter4));
  nand2 gate1588(.a(gate43inter4), .b(gate43inter3), .O(gate43inter5));
  nor2  gate1589(.a(gate43inter5), .b(gate43inter2), .O(gate43inter6));
  inv1  gate1590(.a(G3), .O(gate43inter7));
  inv1  gate1591(.a(G269), .O(gate43inter8));
  nand2 gate1592(.a(gate43inter8), .b(gate43inter7), .O(gate43inter9));
  nand2 gate1593(.a(s_149), .b(gate43inter3), .O(gate43inter10));
  nor2  gate1594(.a(gate43inter10), .b(gate43inter9), .O(gate43inter11));
  nor2  gate1595(.a(gate43inter11), .b(gate43inter6), .O(gate43inter12));
  nand2 gate1596(.a(gate43inter12), .b(gate43inter1), .O(G364));

  xor2  gate2353(.a(G269), .b(G4), .O(gate44inter0));
  nand2 gate2354(.a(gate44inter0), .b(s_258), .O(gate44inter1));
  and2  gate2355(.a(G269), .b(G4), .O(gate44inter2));
  inv1  gate2356(.a(s_258), .O(gate44inter3));
  inv1  gate2357(.a(s_259), .O(gate44inter4));
  nand2 gate2358(.a(gate44inter4), .b(gate44inter3), .O(gate44inter5));
  nor2  gate2359(.a(gate44inter5), .b(gate44inter2), .O(gate44inter6));
  inv1  gate2360(.a(G4), .O(gate44inter7));
  inv1  gate2361(.a(G269), .O(gate44inter8));
  nand2 gate2362(.a(gate44inter8), .b(gate44inter7), .O(gate44inter9));
  nand2 gate2363(.a(s_259), .b(gate44inter3), .O(gate44inter10));
  nor2  gate2364(.a(gate44inter10), .b(gate44inter9), .O(gate44inter11));
  nor2  gate2365(.a(gate44inter11), .b(gate44inter6), .O(gate44inter12));
  nand2 gate2366(.a(gate44inter12), .b(gate44inter1), .O(G365));
nand2 gate45( .a(G5), .b(G272), .O(G366) );
nand2 gate46( .a(G6), .b(G272), .O(G367) );

  xor2  gate827(.a(G275), .b(G7), .O(gate47inter0));
  nand2 gate828(.a(gate47inter0), .b(s_40), .O(gate47inter1));
  and2  gate829(.a(G275), .b(G7), .O(gate47inter2));
  inv1  gate830(.a(s_40), .O(gate47inter3));
  inv1  gate831(.a(s_41), .O(gate47inter4));
  nand2 gate832(.a(gate47inter4), .b(gate47inter3), .O(gate47inter5));
  nor2  gate833(.a(gate47inter5), .b(gate47inter2), .O(gate47inter6));
  inv1  gate834(.a(G7), .O(gate47inter7));
  inv1  gate835(.a(G275), .O(gate47inter8));
  nand2 gate836(.a(gate47inter8), .b(gate47inter7), .O(gate47inter9));
  nand2 gate837(.a(s_41), .b(gate47inter3), .O(gate47inter10));
  nor2  gate838(.a(gate47inter10), .b(gate47inter9), .O(gate47inter11));
  nor2  gate839(.a(gate47inter11), .b(gate47inter6), .O(gate47inter12));
  nand2 gate840(.a(gate47inter12), .b(gate47inter1), .O(G368));

  xor2  gate1051(.a(G275), .b(G8), .O(gate48inter0));
  nand2 gate1052(.a(gate48inter0), .b(s_72), .O(gate48inter1));
  and2  gate1053(.a(G275), .b(G8), .O(gate48inter2));
  inv1  gate1054(.a(s_72), .O(gate48inter3));
  inv1  gate1055(.a(s_73), .O(gate48inter4));
  nand2 gate1056(.a(gate48inter4), .b(gate48inter3), .O(gate48inter5));
  nor2  gate1057(.a(gate48inter5), .b(gate48inter2), .O(gate48inter6));
  inv1  gate1058(.a(G8), .O(gate48inter7));
  inv1  gate1059(.a(G275), .O(gate48inter8));
  nand2 gate1060(.a(gate48inter8), .b(gate48inter7), .O(gate48inter9));
  nand2 gate1061(.a(s_73), .b(gate48inter3), .O(gate48inter10));
  nor2  gate1062(.a(gate48inter10), .b(gate48inter9), .O(gate48inter11));
  nor2  gate1063(.a(gate48inter11), .b(gate48inter6), .O(gate48inter12));
  nand2 gate1064(.a(gate48inter12), .b(gate48inter1), .O(G369));

  xor2  gate2311(.a(G278), .b(G9), .O(gate49inter0));
  nand2 gate2312(.a(gate49inter0), .b(s_252), .O(gate49inter1));
  and2  gate2313(.a(G278), .b(G9), .O(gate49inter2));
  inv1  gate2314(.a(s_252), .O(gate49inter3));
  inv1  gate2315(.a(s_253), .O(gate49inter4));
  nand2 gate2316(.a(gate49inter4), .b(gate49inter3), .O(gate49inter5));
  nor2  gate2317(.a(gate49inter5), .b(gate49inter2), .O(gate49inter6));
  inv1  gate2318(.a(G9), .O(gate49inter7));
  inv1  gate2319(.a(G278), .O(gate49inter8));
  nand2 gate2320(.a(gate49inter8), .b(gate49inter7), .O(gate49inter9));
  nand2 gate2321(.a(s_253), .b(gate49inter3), .O(gate49inter10));
  nor2  gate2322(.a(gate49inter10), .b(gate49inter9), .O(gate49inter11));
  nor2  gate2323(.a(gate49inter11), .b(gate49inter6), .O(gate49inter12));
  nand2 gate2324(.a(gate49inter12), .b(gate49inter1), .O(G370));

  xor2  gate813(.a(G278), .b(G10), .O(gate50inter0));
  nand2 gate814(.a(gate50inter0), .b(s_38), .O(gate50inter1));
  and2  gate815(.a(G278), .b(G10), .O(gate50inter2));
  inv1  gate816(.a(s_38), .O(gate50inter3));
  inv1  gate817(.a(s_39), .O(gate50inter4));
  nand2 gate818(.a(gate50inter4), .b(gate50inter3), .O(gate50inter5));
  nor2  gate819(.a(gate50inter5), .b(gate50inter2), .O(gate50inter6));
  inv1  gate820(.a(G10), .O(gate50inter7));
  inv1  gate821(.a(G278), .O(gate50inter8));
  nand2 gate822(.a(gate50inter8), .b(gate50inter7), .O(gate50inter9));
  nand2 gate823(.a(s_39), .b(gate50inter3), .O(gate50inter10));
  nor2  gate824(.a(gate50inter10), .b(gate50inter9), .O(gate50inter11));
  nor2  gate825(.a(gate50inter11), .b(gate50inter6), .O(gate50inter12));
  nand2 gate826(.a(gate50inter12), .b(gate50inter1), .O(G371));

  xor2  gate575(.a(G281), .b(G11), .O(gate51inter0));
  nand2 gate576(.a(gate51inter0), .b(s_4), .O(gate51inter1));
  and2  gate577(.a(G281), .b(G11), .O(gate51inter2));
  inv1  gate578(.a(s_4), .O(gate51inter3));
  inv1  gate579(.a(s_5), .O(gate51inter4));
  nand2 gate580(.a(gate51inter4), .b(gate51inter3), .O(gate51inter5));
  nor2  gate581(.a(gate51inter5), .b(gate51inter2), .O(gate51inter6));
  inv1  gate582(.a(G11), .O(gate51inter7));
  inv1  gate583(.a(G281), .O(gate51inter8));
  nand2 gate584(.a(gate51inter8), .b(gate51inter7), .O(gate51inter9));
  nand2 gate585(.a(s_5), .b(gate51inter3), .O(gate51inter10));
  nor2  gate586(.a(gate51inter10), .b(gate51inter9), .O(gate51inter11));
  nor2  gate587(.a(gate51inter11), .b(gate51inter6), .O(gate51inter12));
  nand2 gate588(.a(gate51inter12), .b(gate51inter1), .O(G372));

  xor2  gate1387(.a(G281), .b(G12), .O(gate52inter0));
  nand2 gate1388(.a(gate52inter0), .b(s_120), .O(gate52inter1));
  and2  gate1389(.a(G281), .b(G12), .O(gate52inter2));
  inv1  gate1390(.a(s_120), .O(gate52inter3));
  inv1  gate1391(.a(s_121), .O(gate52inter4));
  nand2 gate1392(.a(gate52inter4), .b(gate52inter3), .O(gate52inter5));
  nor2  gate1393(.a(gate52inter5), .b(gate52inter2), .O(gate52inter6));
  inv1  gate1394(.a(G12), .O(gate52inter7));
  inv1  gate1395(.a(G281), .O(gate52inter8));
  nand2 gate1396(.a(gate52inter8), .b(gate52inter7), .O(gate52inter9));
  nand2 gate1397(.a(s_121), .b(gate52inter3), .O(gate52inter10));
  nor2  gate1398(.a(gate52inter10), .b(gate52inter9), .O(gate52inter11));
  nor2  gate1399(.a(gate52inter11), .b(gate52inter6), .O(gate52inter12));
  nand2 gate1400(.a(gate52inter12), .b(gate52inter1), .O(G373));

  xor2  gate1289(.a(G284), .b(G13), .O(gate53inter0));
  nand2 gate1290(.a(gate53inter0), .b(s_106), .O(gate53inter1));
  and2  gate1291(.a(G284), .b(G13), .O(gate53inter2));
  inv1  gate1292(.a(s_106), .O(gate53inter3));
  inv1  gate1293(.a(s_107), .O(gate53inter4));
  nand2 gate1294(.a(gate53inter4), .b(gate53inter3), .O(gate53inter5));
  nor2  gate1295(.a(gate53inter5), .b(gate53inter2), .O(gate53inter6));
  inv1  gate1296(.a(G13), .O(gate53inter7));
  inv1  gate1297(.a(G284), .O(gate53inter8));
  nand2 gate1298(.a(gate53inter8), .b(gate53inter7), .O(gate53inter9));
  nand2 gate1299(.a(s_107), .b(gate53inter3), .O(gate53inter10));
  nor2  gate1300(.a(gate53inter10), .b(gate53inter9), .O(gate53inter11));
  nor2  gate1301(.a(gate53inter11), .b(gate53inter6), .O(gate53inter12));
  nand2 gate1302(.a(gate53inter12), .b(gate53inter1), .O(G374));

  xor2  gate2367(.a(G284), .b(G14), .O(gate54inter0));
  nand2 gate2368(.a(gate54inter0), .b(s_260), .O(gate54inter1));
  and2  gate2369(.a(G284), .b(G14), .O(gate54inter2));
  inv1  gate2370(.a(s_260), .O(gate54inter3));
  inv1  gate2371(.a(s_261), .O(gate54inter4));
  nand2 gate2372(.a(gate54inter4), .b(gate54inter3), .O(gate54inter5));
  nor2  gate2373(.a(gate54inter5), .b(gate54inter2), .O(gate54inter6));
  inv1  gate2374(.a(G14), .O(gate54inter7));
  inv1  gate2375(.a(G284), .O(gate54inter8));
  nand2 gate2376(.a(gate54inter8), .b(gate54inter7), .O(gate54inter9));
  nand2 gate2377(.a(s_261), .b(gate54inter3), .O(gate54inter10));
  nor2  gate2378(.a(gate54inter10), .b(gate54inter9), .O(gate54inter11));
  nor2  gate2379(.a(gate54inter11), .b(gate54inter6), .O(gate54inter12));
  nand2 gate2380(.a(gate54inter12), .b(gate54inter1), .O(G375));

  xor2  gate2591(.a(G287), .b(G15), .O(gate55inter0));
  nand2 gate2592(.a(gate55inter0), .b(s_292), .O(gate55inter1));
  and2  gate2593(.a(G287), .b(G15), .O(gate55inter2));
  inv1  gate2594(.a(s_292), .O(gate55inter3));
  inv1  gate2595(.a(s_293), .O(gate55inter4));
  nand2 gate2596(.a(gate55inter4), .b(gate55inter3), .O(gate55inter5));
  nor2  gate2597(.a(gate55inter5), .b(gate55inter2), .O(gate55inter6));
  inv1  gate2598(.a(G15), .O(gate55inter7));
  inv1  gate2599(.a(G287), .O(gate55inter8));
  nand2 gate2600(.a(gate55inter8), .b(gate55inter7), .O(gate55inter9));
  nand2 gate2601(.a(s_293), .b(gate55inter3), .O(gate55inter10));
  nor2  gate2602(.a(gate55inter10), .b(gate55inter9), .O(gate55inter11));
  nor2  gate2603(.a(gate55inter11), .b(gate55inter6), .O(gate55inter12));
  nand2 gate2604(.a(gate55inter12), .b(gate55inter1), .O(G376));

  xor2  gate2381(.a(G287), .b(G16), .O(gate56inter0));
  nand2 gate2382(.a(gate56inter0), .b(s_262), .O(gate56inter1));
  and2  gate2383(.a(G287), .b(G16), .O(gate56inter2));
  inv1  gate2384(.a(s_262), .O(gate56inter3));
  inv1  gate2385(.a(s_263), .O(gate56inter4));
  nand2 gate2386(.a(gate56inter4), .b(gate56inter3), .O(gate56inter5));
  nor2  gate2387(.a(gate56inter5), .b(gate56inter2), .O(gate56inter6));
  inv1  gate2388(.a(G16), .O(gate56inter7));
  inv1  gate2389(.a(G287), .O(gate56inter8));
  nand2 gate2390(.a(gate56inter8), .b(gate56inter7), .O(gate56inter9));
  nand2 gate2391(.a(s_263), .b(gate56inter3), .O(gate56inter10));
  nor2  gate2392(.a(gate56inter10), .b(gate56inter9), .O(gate56inter11));
  nor2  gate2393(.a(gate56inter11), .b(gate56inter6), .O(gate56inter12));
  nand2 gate2394(.a(gate56inter12), .b(gate56inter1), .O(G377));
nand2 gate57( .a(G17), .b(G290), .O(G378) );
nand2 gate58( .a(G18), .b(G290), .O(G379) );
nand2 gate59( .a(G19), .b(G293), .O(G380) );
nand2 gate60( .a(G20), .b(G293), .O(G381) );

  xor2  gate1331(.a(G296), .b(G21), .O(gate61inter0));
  nand2 gate1332(.a(gate61inter0), .b(s_112), .O(gate61inter1));
  and2  gate1333(.a(G296), .b(G21), .O(gate61inter2));
  inv1  gate1334(.a(s_112), .O(gate61inter3));
  inv1  gate1335(.a(s_113), .O(gate61inter4));
  nand2 gate1336(.a(gate61inter4), .b(gate61inter3), .O(gate61inter5));
  nor2  gate1337(.a(gate61inter5), .b(gate61inter2), .O(gate61inter6));
  inv1  gate1338(.a(G21), .O(gate61inter7));
  inv1  gate1339(.a(G296), .O(gate61inter8));
  nand2 gate1340(.a(gate61inter8), .b(gate61inter7), .O(gate61inter9));
  nand2 gate1341(.a(s_113), .b(gate61inter3), .O(gate61inter10));
  nor2  gate1342(.a(gate61inter10), .b(gate61inter9), .O(gate61inter11));
  nor2  gate1343(.a(gate61inter11), .b(gate61inter6), .O(gate61inter12));
  nand2 gate1344(.a(gate61inter12), .b(gate61inter1), .O(G382));

  xor2  gate1149(.a(G296), .b(G22), .O(gate62inter0));
  nand2 gate1150(.a(gate62inter0), .b(s_86), .O(gate62inter1));
  and2  gate1151(.a(G296), .b(G22), .O(gate62inter2));
  inv1  gate1152(.a(s_86), .O(gate62inter3));
  inv1  gate1153(.a(s_87), .O(gate62inter4));
  nand2 gate1154(.a(gate62inter4), .b(gate62inter3), .O(gate62inter5));
  nor2  gate1155(.a(gate62inter5), .b(gate62inter2), .O(gate62inter6));
  inv1  gate1156(.a(G22), .O(gate62inter7));
  inv1  gate1157(.a(G296), .O(gate62inter8));
  nand2 gate1158(.a(gate62inter8), .b(gate62inter7), .O(gate62inter9));
  nand2 gate1159(.a(s_87), .b(gate62inter3), .O(gate62inter10));
  nor2  gate1160(.a(gate62inter10), .b(gate62inter9), .O(gate62inter11));
  nor2  gate1161(.a(gate62inter11), .b(gate62inter6), .O(gate62inter12));
  nand2 gate1162(.a(gate62inter12), .b(gate62inter1), .O(G383));
nand2 gate63( .a(G23), .b(G299), .O(G384) );

  xor2  gate1779(.a(G299), .b(G24), .O(gate64inter0));
  nand2 gate1780(.a(gate64inter0), .b(s_176), .O(gate64inter1));
  and2  gate1781(.a(G299), .b(G24), .O(gate64inter2));
  inv1  gate1782(.a(s_176), .O(gate64inter3));
  inv1  gate1783(.a(s_177), .O(gate64inter4));
  nand2 gate1784(.a(gate64inter4), .b(gate64inter3), .O(gate64inter5));
  nor2  gate1785(.a(gate64inter5), .b(gate64inter2), .O(gate64inter6));
  inv1  gate1786(.a(G24), .O(gate64inter7));
  inv1  gate1787(.a(G299), .O(gate64inter8));
  nand2 gate1788(.a(gate64inter8), .b(gate64inter7), .O(gate64inter9));
  nand2 gate1789(.a(s_177), .b(gate64inter3), .O(gate64inter10));
  nor2  gate1790(.a(gate64inter10), .b(gate64inter9), .O(gate64inter11));
  nor2  gate1791(.a(gate64inter11), .b(gate64inter6), .O(gate64inter12));
  nand2 gate1792(.a(gate64inter12), .b(gate64inter1), .O(G385));
nand2 gate65( .a(G25), .b(G302), .O(G386) );
nand2 gate66( .a(G26), .b(G302), .O(G387) );

  xor2  gate757(.a(G305), .b(G27), .O(gate67inter0));
  nand2 gate758(.a(gate67inter0), .b(s_30), .O(gate67inter1));
  and2  gate759(.a(G305), .b(G27), .O(gate67inter2));
  inv1  gate760(.a(s_30), .O(gate67inter3));
  inv1  gate761(.a(s_31), .O(gate67inter4));
  nand2 gate762(.a(gate67inter4), .b(gate67inter3), .O(gate67inter5));
  nor2  gate763(.a(gate67inter5), .b(gate67inter2), .O(gate67inter6));
  inv1  gate764(.a(G27), .O(gate67inter7));
  inv1  gate765(.a(G305), .O(gate67inter8));
  nand2 gate766(.a(gate67inter8), .b(gate67inter7), .O(gate67inter9));
  nand2 gate767(.a(s_31), .b(gate67inter3), .O(gate67inter10));
  nor2  gate768(.a(gate67inter10), .b(gate67inter9), .O(gate67inter11));
  nor2  gate769(.a(gate67inter11), .b(gate67inter6), .O(gate67inter12));
  nand2 gate770(.a(gate67inter12), .b(gate67inter1), .O(G388));
nand2 gate68( .a(G28), .b(G305), .O(G389) );

  xor2  gate1079(.a(G308), .b(G29), .O(gate69inter0));
  nand2 gate1080(.a(gate69inter0), .b(s_76), .O(gate69inter1));
  and2  gate1081(.a(G308), .b(G29), .O(gate69inter2));
  inv1  gate1082(.a(s_76), .O(gate69inter3));
  inv1  gate1083(.a(s_77), .O(gate69inter4));
  nand2 gate1084(.a(gate69inter4), .b(gate69inter3), .O(gate69inter5));
  nor2  gate1085(.a(gate69inter5), .b(gate69inter2), .O(gate69inter6));
  inv1  gate1086(.a(G29), .O(gate69inter7));
  inv1  gate1087(.a(G308), .O(gate69inter8));
  nand2 gate1088(.a(gate69inter8), .b(gate69inter7), .O(gate69inter9));
  nand2 gate1089(.a(s_77), .b(gate69inter3), .O(gate69inter10));
  nor2  gate1090(.a(gate69inter10), .b(gate69inter9), .O(gate69inter11));
  nor2  gate1091(.a(gate69inter11), .b(gate69inter6), .O(gate69inter12));
  nand2 gate1092(.a(gate69inter12), .b(gate69inter1), .O(G390));
nand2 gate70( .a(G30), .b(G308), .O(G391) );
nand2 gate71( .a(G31), .b(G311), .O(G392) );

  xor2  gate925(.a(G311), .b(G32), .O(gate72inter0));
  nand2 gate926(.a(gate72inter0), .b(s_54), .O(gate72inter1));
  and2  gate927(.a(G311), .b(G32), .O(gate72inter2));
  inv1  gate928(.a(s_54), .O(gate72inter3));
  inv1  gate929(.a(s_55), .O(gate72inter4));
  nand2 gate930(.a(gate72inter4), .b(gate72inter3), .O(gate72inter5));
  nor2  gate931(.a(gate72inter5), .b(gate72inter2), .O(gate72inter6));
  inv1  gate932(.a(G32), .O(gate72inter7));
  inv1  gate933(.a(G311), .O(gate72inter8));
  nand2 gate934(.a(gate72inter8), .b(gate72inter7), .O(gate72inter9));
  nand2 gate935(.a(s_55), .b(gate72inter3), .O(gate72inter10));
  nor2  gate936(.a(gate72inter10), .b(gate72inter9), .O(gate72inter11));
  nor2  gate937(.a(gate72inter11), .b(gate72inter6), .O(gate72inter12));
  nand2 gate938(.a(gate72inter12), .b(gate72inter1), .O(G393));

  xor2  gate1737(.a(G314), .b(G1), .O(gate73inter0));
  nand2 gate1738(.a(gate73inter0), .b(s_170), .O(gate73inter1));
  and2  gate1739(.a(G314), .b(G1), .O(gate73inter2));
  inv1  gate1740(.a(s_170), .O(gate73inter3));
  inv1  gate1741(.a(s_171), .O(gate73inter4));
  nand2 gate1742(.a(gate73inter4), .b(gate73inter3), .O(gate73inter5));
  nor2  gate1743(.a(gate73inter5), .b(gate73inter2), .O(gate73inter6));
  inv1  gate1744(.a(G1), .O(gate73inter7));
  inv1  gate1745(.a(G314), .O(gate73inter8));
  nand2 gate1746(.a(gate73inter8), .b(gate73inter7), .O(gate73inter9));
  nand2 gate1747(.a(s_171), .b(gate73inter3), .O(gate73inter10));
  nor2  gate1748(.a(gate73inter10), .b(gate73inter9), .O(gate73inter11));
  nor2  gate1749(.a(gate73inter11), .b(gate73inter6), .O(gate73inter12));
  nand2 gate1750(.a(gate73inter12), .b(gate73inter1), .O(G394));

  xor2  gate1765(.a(G314), .b(G5), .O(gate74inter0));
  nand2 gate1766(.a(gate74inter0), .b(s_174), .O(gate74inter1));
  and2  gate1767(.a(G314), .b(G5), .O(gate74inter2));
  inv1  gate1768(.a(s_174), .O(gate74inter3));
  inv1  gate1769(.a(s_175), .O(gate74inter4));
  nand2 gate1770(.a(gate74inter4), .b(gate74inter3), .O(gate74inter5));
  nor2  gate1771(.a(gate74inter5), .b(gate74inter2), .O(gate74inter6));
  inv1  gate1772(.a(G5), .O(gate74inter7));
  inv1  gate1773(.a(G314), .O(gate74inter8));
  nand2 gate1774(.a(gate74inter8), .b(gate74inter7), .O(gate74inter9));
  nand2 gate1775(.a(s_175), .b(gate74inter3), .O(gate74inter10));
  nor2  gate1776(.a(gate74inter10), .b(gate74inter9), .O(gate74inter11));
  nor2  gate1777(.a(gate74inter11), .b(gate74inter6), .O(gate74inter12));
  nand2 gate1778(.a(gate74inter12), .b(gate74inter1), .O(G395));
nand2 gate75( .a(G9), .b(G317), .O(G396) );
nand2 gate76( .a(G13), .b(G317), .O(G397) );
nand2 gate77( .a(G2), .b(G320), .O(G398) );
nand2 gate78( .a(G6), .b(G320), .O(G399) );
nand2 gate79( .a(G10), .b(G323), .O(G400) );
nand2 gate80( .a(G14), .b(G323), .O(G401) );

  xor2  gate701(.a(G326), .b(G3), .O(gate81inter0));
  nand2 gate702(.a(gate81inter0), .b(s_22), .O(gate81inter1));
  and2  gate703(.a(G326), .b(G3), .O(gate81inter2));
  inv1  gate704(.a(s_22), .O(gate81inter3));
  inv1  gate705(.a(s_23), .O(gate81inter4));
  nand2 gate706(.a(gate81inter4), .b(gate81inter3), .O(gate81inter5));
  nor2  gate707(.a(gate81inter5), .b(gate81inter2), .O(gate81inter6));
  inv1  gate708(.a(G3), .O(gate81inter7));
  inv1  gate709(.a(G326), .O(gate81inter8));
  nand2 gate710(.a(gate81inter8), .b(gate81inter7), .O(gate81inter9));
  nand2 gate711(.a(s_23), .b(gate81inter3), .O(gate81inter10));
  nor2  gate712(.a(gate81inter10), .b(gate81inter9), .O(gate81inter11));
  nor2  gate713(.a(gate81inter11), .b(gate81inter6), .O(gate81inter12));
  nand2 gate714(.a(gate81inter12), .b(gate81inter1), .O(G402));
nand2 gate82( .a(G7), .b(G326), .O(G403) );
nand2 gate83( .a(G11), .b(G329), .O(G404) );

  xor2  gate1555(.a(G329), .b(G15), .O(gate84inter0));
  nand2 gate1556(.a(gate84inter0), .b(s_144), .O(gate84inter1));
  and2  gate1557(.a(G329), .b(G15), .O(gate84inter2));
  inv1  gate1558(.a(s_144), .O(gate84inter3));
  inv1  gate1559(.a(s_145), .O(gate84inter4));
  nand2 gate1560(.a(gate84inter4), .b(gate84inter3), .O(gate84inter5));
  nor2  gate1561(.a(gate84inter5), .b(gate84inter2), .O(gate84inter6));
  inv1  gate1562(.a(G15), .O(gate84inter7));
  inv1  gate1563(.a(G329), .O(gate84inter8));
  nand2 gate1564(.a(gate84inter8), .b(gate84inter7), .O(gate84inter9));
  nand2 gate1565(.a(s_145), .b(gate84inter3), .O(gate84inter10));
  nor2  gate1566(.a(gate84inter10), .b(gate84inter9), .O(gate84inter11));
  nor2  gate1567(.a(gate84inter11), .b(gate84inter6), .O(gate84inter12));
  nand2 gate1568(.a(gate84inter12), .b(gate84inter1), .O(G405));

  xor2  gate2171(.a(G332), .b(G4), .O(gate85inter0));
  nand2 gate2172(.a(gate85inter0), .b(s_232), .O(gate85inter1));
  and2  gate2173(.a(G332), .b(G4), .O(gate85inter2));
  inv1  gate2174(.a(s_232), .O(gate85inter3));
  inv1  gate2175(.a(s_233), .O(gate85inter4));
  nand2 gate2176(.a(gate85inter4), .b(gate85inter3), .O(gate85inter5));
  nor2  gate2177(.a(gate85inter5), .b(gate85inter2), .O(gate85inter6));
  inv1  gate2178(.a(G4), .O(gate85inter7));
  inv1  gate2179(.a(G332), .O(gate85inter8));
  nand2 gate2180(.a(gate85inter8), .b(gate85inter7), .O(gate85inter9));
  nand2 gate2181(.a(s_233), .b(gate85inter3), .O(gate85inter10));
  nor2  gate2182(.a(gate85inter10), .b(gate85inter9), .O(gate85inter11));
  nor2  gate2183(.a(gate85inter11), .b(gate85inter6), .O(gate85inter12));
  nand2 gate2184(.a(gate85inter12), .b(gate85inter1), .O(G406));
nand2 gate86( .a(G8), .b(G332), .O(G407) );

  xor2  gate2647(.a(G335), .b(G12), .O(gate87inter0));
  nand2 gate2648(.a(gate87inter0), .b(s_300), .O(gate87inter1));
  and2  gate2649(.a(G335), .b(G12), .O(gate87inter2));
  inv1  gate2650(.a(s_300), .O(gate87inter3));
  inv1  gate2651(.a(s_301), .O(gate87inter4));
  nand2 gate2652(.a(gate87inter4), .b(gate87inter3), .O(gate87inter5));
  nor2  gate2653(.a(gate87inter5), .b(gate87inter2), .O(gate87inter6));
  inv1  gate2654(.a(G12), .O(gate87inter7));
  inv1  gate2655(.a(G335), .O(gate87inter8));
  nand2 gate2656(.a(gate87inter8), .b(gate87inter7), .O(gate87inter9));
  nand2 gate2657(.a(s_301), .b(gate87inter3), .O(gate87inter10));
  nor2  gate2658(.a(gate87inter10), .b(gate87inter9), .O(gate87inter11));
  nor2  gate2659(.a(gate87inter11), .b(gate87inter6), .O(gate87inter12));
  nand2 gate2660(.a(gate87inter12), .b(gate87inter1), .O(G408));

  xor2  gate1905(.a(G335), .b(G16), .O(gate88inter0));
  nand2 gate1906(.a(gate88inter0), .b(s_194), .O(gate88inter1));
  and2  gate1907(.a(G335), .b(G16), .O(gate88inter2));
  inv1  gate1908(.a(s_194), .O(gate88inter3));
  inv1  gate1909(.a(s_195), .O(gate88inter4));
  nand2 gate1910(.a(gate88inter4), .b(gate88inter3), .O(gate88inter5));
  nor2  gate1911(.a(gate88inter5), .b(gate88inter2), .O(gate88inter6));
  inv1  gate1912(.a(G16), .O(gate88inter7));
  inv1  gate1913(.a(G335), .O(gate88inter8));
  nand2 gate1914(.a(gate88inter8), .b(gate88inter7), .O(gate88inter9));
  nand2 gate1915(.a(s_195), .b(gate88inter3), .O(gate88inter10));
  nor2  gate1916(.a(gate88inter10), .b(gate88inter9), .O(gate88inter11));
  nor2  gate1917(.a(gate88inter11), .b(gate88inter6), .O(gate88inter12));
  nand2 gate1918(.a(gate88inter12), .b(gate88inter1), .O(G409));
nand2 gate89( .a(G17), .b(G338), .O(G410) );
nand2 gate90( .a(G21), .b(G338), .O(G411) );
nand2 gate91( .a(G25), .b(G341), .O(G412) );

  xor2  gate2031(.a(G341), .b(G29), .O(gate92inter0));
  nand2 gate2032(.a(gate92inter0), .b(s_212), .O(gate92inter1));
  and2  gate2033(.a(G341), .b(G29), .O(gate92inter2));
  inv1  gate2034(.a(s_212), .O(gate92inter3));
  inv1  gate2035(.a(s_213), .O(gate92inter4));
  nand2 gate2036(.a(gate92inter4), .b(gate92inter3), .O(gate92inter5));
  nor2  gate2037(.a(gate92inter5), .b(gate92inter2), .O(gate92inter6));
  inv1  gate2038(.a(G29), .O(gate92inter7));
  inv1  gate2039(.a(G341), .O(gate92inter8));
  nand2 gate2040(.a(gate92inter8), .b(gate92inter7), .O(gate92inter9));
  nand2 gate2041(.a(s_213), .b(gate92inter3), .O(gate92inter10));
  nor2  gate2042(.a(gate92inter10), .b(gate92inter9), .O(gate92inter11));
  nor2  gate2043(.a(gate92inter11), .b(gate92inter6), .O(gate92inter12));
  nand2 gate2044(.a(gate92inter12), .b(gate92inter1), .O(G413));
nand2 gate93( .a(G18), .b(G344), .O(G414) );
nand2 gate94( .a(G22), .b(G344), .O(G415) );
nand2 gate95( .a(G26), .b(G347), .O(G416) );
nand2 gate96( .a(G30), .b(G347), .O(G417) );
nand2 gate97( .a(G19), .b(G350), .O(G418) );

  xor2  gate2101(.a(G350), .b(G23), .O(gate98inter0));
  nand2 gate2102(.a(gate98inter0), .b(s_222), .O(gate98inter1));
  and2  gate2103(.a(G350), .b(G23), .O(gate98inter2));
  inv1  gate2104(.a(s_222), .O(gate98inter3));
  inv1  gate2105(.a(s_223), .O(gate98inter4));
  nand2 gate2106(.a(gate98inter4), .b(gate98inter3), .O(gate98inter5));
  nor2  gate2107(.a(gate98inter5), .b(gate98inter2), .O(gate98inter6));
  inv1  gate2108(.a(G23), .O(gate98inter7));
  inv1  gate2109(.a(G350), .O(gate98inter8));
  nand2 gate2110(.a(gate98inter8), .b(gate98inter7), .O(gate98inter9));
  nand2 gate2111(.a(s_223), .b(gate98inter3), .O(gate98inter10));
  nor2  gate2112(.a(gate98inter10), .b(gate98inter9), .O(gate98inter11));
  nor2  gate2113(.a(gate98inter11), .b(gate98inter6), .O(gate98inter12));
  nand2 gate2114(.a(gate98inter12), .b(gate98inter1), .O(G419));

  xor2  gate645(.a(G353), .b(G27), .O(gate99inter0));
  nand2 gate646(.a(gate99inter0), .b(s_14), .O(gate99inter1));
  and2  gate647(.a(G353), .b(G27), .O(gate99inter2));
  inv1  gate648(.a(s_14), .O(gate99inter3));
  inv1  gate649(.a(s_15), .O(gate99inter4));
  nand2 gate650(.a(gate99inter4), .b(gate99inter3), .O(gate99inter5));
  nor2  gate651(.a(gate99inter5), .b(gate99inter2), .O(gate99inter6));
  inv1  gate652(.a(G27), .O(gate99inter7));
  inv1  gate653(.a(G353), .O(gate99inter8));
  nand2 gate654(.a(gate99inter8), .b(gate99inter7), .O(gate99inter9));
  nand2 gate655(.a(s_15), .b(gate99inter3), .O(gate99inter10));
  nor2  gate656(.a(gate99inter10), .b(gate99inter9), .O(gate99inter11));
  nor2  gate657(.a(gate99inter11), .b(gate99inter6), .O(gate99inter12));
  nand2 gate658(.a(gate99inter12), .b(gate99inter1), .O(G420));
nand2 gate100( .a(G31), .b(G353), .O(G421) );

  xor2  gate2423(.a(G356), .b(G20), .O(gate101inter0));
  nand2 gate2424(.a(gate101inter0), .b(s_268), .O(gate101inter1));
  and2  gate2425(.a(G356), .b(G20), .O(gate101inter2));
  inv1  gate2426(.a(s_268), .O(gate101inter3));
  inv1  gate2427(.a(s_269), .O(gate101inter4));
  nand2 gate2428(.a(gate101inter4), .b(gate101inter3), .O(gate101inter5));
  nor2  gate2429(.a(gate101inter5), .b(gate101inter2), .O(gate101inter6));
  inv1  gate2430(.a(G20), .O(gate101inter7));
  inv1  gate2431(.a(G356), .O(gate101inter8));
  nand2 gate2432(.a(gate101inter8), .b(gate101inter7), .O(gate101inter9));
  nand2 gate2433(.a(s_269), .b(gate101inter3), .O(gate101inter10));
  nor2  gate2434(.a(gate101inter10), .b(gate101inter9), .O(gate101inter11));
  nor2  gate2435(.a(gate101inter11), .b(gate101inter6), .O(gate101inter12));
  nand2 gate2436(.a(gate101inter12), .b(gate101inter1), .O(G422));

  xor2  gate2535(.a(G356), .b(G24), .O(gate102inter0));
  nand2 gate2536(.a(gate102inter0), .b(s_284), .O(gate102inter1));
  and2  gate2537(.a(G356), .b(G24), .O(gate102inter2));
  inv1  gate2538(.a(s_284), .O(gate102inter3));
  inv1  gate2539(.a(s_285), .O(gate102inter4));
  nand2 gate2540(.a(gate102inter4), .b(gate102inter3), .O(gate102inter5));
  nor2  gate2541(.a(gate102inter5), .b(gate102inter2), .O(gate102inter6));
  inv1  gate2542(.a(G24), .O(gate102inter7));
  inv1  gate2543(.a(G356), .O(gate102inter8));
  nand2 gate2544(.a(gate102inter8), .b(gate102inter7), .O(gate102inter9));
  nand2 gate2545(.a(s_285), .b(gate102inter3), .O(gate102inter10));
  nor2  gate2546(.a(gate102inter10), .b(gate102inter9), .O(gate102inter11));
  nor2  gate2547(.a(gate102inter11), .b(gate102inter6), .O(gate102inter12));
  nand2 gate2548(.a(gate102inter12), .b(gate102inter1), .O(G423));
nand2 gate103( .a(G28), .b(G359), .O(G424) );
nand2 gate104( .a(G32), .b(G359), .O(G425) );
nand2 gate105( .a(G362), .b(G363), .O(G426) );

  xor2  gate617(.a(G365), .b(G364), .O(gate106inter0));
  nand2 gate618(.a(gate106inter0), .b(s_10), .O(gate106inter1));
  and2  gate619(.a(G365), .b(G364), .O(gate106inter2));
  inv1  gate620(.a(s_10), .O(gate106inter3));
  inv1  gate621(.a(s_11), .O(gate106inter4));
  nand2 gate622(.a(gate106inter4), .b(gate106inter3), .O(gate106inter5));
  nor2  gate623(.a(gate106inter5), .b(gate106inter2), .O(gate106inter6));
  inv1  gate624(.a(G364), .O(gate106inter7));
  inv1  gate625(.a(G365), .O(gate106inter8));
  nand2 gate626(.a(gate106inter8), .b(gate106inter7), .O(gate106inter9));
  nand2 gate627(.a(s_11), .b(gate106inter3), .O(gate106inter10));
  nor2  gate628(.a(gate106inter10), .b(gate106inter9), .O(gate106inter11));
  nor2  gate629(.a(gate106inter11), .b(gate106inter6), .O(gate106inter12));
  nand2 gate630(.a(gate106inter12), .b(gate106inter1), .O(G429));

  xor2  gate953(.a(G367), .b(G366), .O(gate107inter0));
  nand2 gate954(.a(gate107inter0), .b(s_58), .O(gate107inter1));
  and2  gate955(.a(G367), .b(G366), .O(gate107inter2));
  inv1  gate956(.a(s_58), .O(gate107inter3));
  inv1  gate957(.a(s_59), .O(gate107inter4));
  nand2 gate958(.a(gate107inter4), .b(gate107inter3), .O(gate107inter5));
  nor2  gate959(.a(gate107inter5), .b(gate107inter2), .O(gate107inter6));
  inv1  gate960(.a(G366), .O(gate107inter7));
  inv1  gate961(.a(G367), .O(gate107inter8));
  nand2 gate962(.a(gate107inter8), .b(gate107inter7), .O(gate107inter9));
  nand2 gate963(.a(s_59), .b(gate107inter3), .O(gate107inter10));
  nor2  gate964(.a(gate107inter10), .b(gate107inter9), .O(gate107inter11));
  nor2  gate965(.a(gate107inter11), .b(gate107inter6), .O(gate107inter12));
  nand2 gate966(.a(gate107inter12), .b(gate107inter1), .O(G432));
nand2 gate108( .a(G368), .b(G369), .O(G435) );
nand2 gate109( .a(G370), .b(G371), .O(G438) );
nand2 gate110( .a(G372), .b(G373), .O(G441) );
nand2 gate111( .a(G374), .b(G375), .O(G444) );
nand2 gate112( .a(G376), .b(G377), .O(G447) );
nand2 gate113( .a(G378), .b(G379), .O(G450) );
nand2 gate114( .a(G380), .b(G381), .O(G453) );

  xor2  gate1877(.a(G383), .b(G382), .O(gate115inter0));
  nand2 gate1878(.a(gate115inter0), .b(s_190), .O(gate115inter1));
  and2  gate1879(.a(G383), .b(G382), .O(gate115inter2));
  inv1  gate1880(.a(s_190), .O(gate115inter3));
  inv1  gate1881(.a(s_191), .O(gate115inter4));
  nand2 gate1882(.a(gate115inter4), .b(gate115inter3), .O(gate115inter5));
  nor2  gate1883(.a(gate115inter5), .b(gate115inter2), .O(gate115inter6));
  inv1  gate1884(.a(G382), .O(gate115inter7));
  inv1  gate1885(.a(G383), .O(gate115inter8));
  nand2 gate1886(.a(gate115inter8), .b(gate115inter7), .O(gate115inter9));
  nand2 gate1887(.a(s_191), .b(gate115inter3), .O(gate115inter10));
  nor2  gate1888(.a(gate115inter10), .b(gate115inter9), .O(gate115inter11));
  nor2  gate1889(.a(gate115inter11), .b(gate115inter6), .O(gate115inter12));
  nand2 gate1890(.a(gate115inter12), .b(gate115inter1), .O(G456));
nand2 gate116( .a(G384), .b(G385), .O(G459) );
nand2 gate117( .a(G386), .b(G387), .O(G462) );
nand2 gate118( .a(G388), .b(G389), .O(G465) );

  xor2  gate1065(.a(G391), .b(G390), .O(gate119inter0));
  nand2 gate1066(.a(gate119inter0), .b(s_74), .O(gate119inter1));
  and2  gate1067(.a(G391), .b(G390), .O(gate119inter2));
  inv1  gate1068(.a(s_74), .O(gate119inter3));
  inv1  gate1069(.a(s_75), .O(gate119inter4));
  nand2 gate1070(.a(gate119inter4), .b(gate119inter3), .O(gate119inter5));
  nor2  gate1071(.a(gate119inter5), .b(gate119inter2), .O(gate119inter6));
  inv1  gate1072(.a(G390), .O(gate119inter7));
  inv1  gate1073(.a(G391), .O(gate119inter8));
  nand2 gate1074(.a(gate119inter8), .b(gate119inter7), .O(gate119inter9));
  nand2 gate1075(.a(s_75), .b(gate119inter3), .O(gate119inter10));
  nor2  gate1076(.a(gate119inter10), .b(gate119inter9), .O(gate119inter11));
  nor2  gate1077(.a(gate119inter11), .b(gate119inter6), .O(gate119inter12));
  nand2 gate1078(.a(gate119inter12), .b(gate119inter1), .O(G468));
nand2 gate120( .a(G392), .b(G393), .O(G471) );
nand2 gate121( .a(G394), .b(G395), .O(G474) );
nand2 gate122( .a(G396), .b(G397), .O(G477) );

  xor2  gate2241(.a(G399), .b(G398), .O(gate123inter0));
  nand2 gate2242(.a(gate123inter0), .b(s_242), .O(gate123inter1));
  and2  gate2243(.a(G399), .b(G398), .O(gate123inter2));
  inv1  gate2244(.a(s_242), .O(gate123inter3));
  inv1  gate2245(.a(s_243), .O(gate123inter4));
  nand2 gate2246(.a(gate123inter4), .b(gate123inter3), .O(gate123inter5));
  nor2  gate2247(.a(gate123inter5), .b(gate123inter2), .O(gate123inter6));
  inv1  gate2248(.a(G398), .O(gate123inter7));
  inv1  gate2249(.a(G399), .O(gate123inter8));
  nand2 gate2250(.a(gate123inter8), .b(gate123inter7), .O(gate123inter9));
  nand2 gate2251(.a(s_243), .b(gate123inter3), .O(gate123inter10));
  nor2  gate2252(.a(gate123inter10), .b(gate123inter9), .O(gate123inter11));
  nor2  gate2253(.a(gate123inter11), .b(gate123inter6), .O(gate123inter12));
  nand2 gate2254(.a(gate123inter12), .b(gate123inter1), .O(G480));
nand2 gate124( .a(G400), .b(G401), .O(G483) );
nand2 gate125( .a(G402), .b(G403), .O(G486) );

  xor2  gate1989(.a(G405), .b(G404), .O(gate126inter0));
  nand2 gate1990(.a(gate126inter0), .b(s_206), .O(gate126inter1));
  and2  gate1991(.a(G405), .b(G404), .O(gate126inter2));
  inv1  gate1992(.a(s_206), .O(gate126inter3));
  inv1  gate1993(.a(s_207), .O(gate126inter4));
  nand2 gate1994(.a(gate126inter4), .b(gate126inter3), .O(gate126inter5));
  nor2  gate1995(.a(gate126inter5), .b(gate126inter2), .O(gate126inter6));
  inv1  gate1996(.a(G404), .O(gate126inter7));
  inv1  gate1997(.a(G405), .O(gate126inter8));
  nand2 gate1998(.a(gate126inter8), .b(gate126inter7), .O(gate126inter9));
  nand2 gate1999(.a(s_207), .b(gate126inter3), .O(gate126inter10));
  nor2  gate2000(.a(gate126inter10), .b(gate126inter9), .O(gate126inter11));
  nor2  gate2001(.a(gate126inter11), .b(gate126inter6), .O(gate126inter12));
  nand2 gate2002(.a(gate126inter12), .b(gate126inter1), .O(G489));
nand2 gate127( .a(G406), .b(G407), .O(G492) );

  xor2  gate1919(.a(G409), .b(G408), .O(gate128inter0));
  nand2 gate1920(.a(gate128inter0), .b(s_196), .O(gate128inter1));
  and2  gate1921(.a(G409), .b(G408), .O(gate128inter2));
  inv1  gate1922(.a(s_196), .O(gate128inter3));
  inv1  gate1923(.a(s_197), .O(gate128inter4));
  nand2 gate1924(.a(gate128inter4), .b(gate128inter3), .O(gate128inter5));
  nor2  gate1925(.a(gate128inter5), .b(gate128inter2), .O(gate128inter6));
  inv1  gate1926(.a(G408), .O(gate128inter7));
  inv1  gate1927(.a(G409), .O(gate128inter8));
  nand2 gate1928(.a(gate128inter8), .b(gate128inter7), .O(gate128inter9));
  nand2 gate1929(.a(s_197), .b(gate128inter3), .O(gate128inter10));
  nor2  gate1930(.a(gate128inter10), .b(gate128inter9), .O(gate128inter11));
  nor2  gate1931(.a(gate128inter11), .b(gate128inter6), .O(gate128inter12));
  nand2 gate1932(.a(gate128inter12), .b(gate128inter1), .O(G495));
nand2 gate129( .a(G410), .b(G411), .O(G498) );
nand2 gate130( .a(G412), .b(G413), .O(G501) );
nand2 gate131( .a(G414), .b(G415), .O(G504) );
nand2 gate132( .a(G416), .b(G417), .O(G507) );
nand2 gate133( .a(G418), .b(G419), .O(G510) );
nand2 gate134( .a(G420), .b(G421), .O(G513) );
nand2 gate135( .a(G422), .b(G423), .O(G516) );
nand2 gate136( .a(G424), .b(G425), .O(G519) );
nand2 gate137( .a(G426), .b(G429), .O(G522) );
nand2 gate138( .a(G432), .b(G435), .O(G525) );

  xor2  gate2633(.a(G441), .b(G438), .O(gate139inter0));
  nand2 gate2634(.a(gate139inter0), .b(s_298), .O(gate139inter1));
  and2  gate2635(.a(G441), .b(G438), .O(gate139inter2));
  inv1  gate2636(.a(s_298), .O(gate139inter3));
  inv1  gate2637(.a(s_299), .O(gate139inter4));
  nand2 gate2638(.a(gate139inter4), .b(gate139inter3), .O(gate139inter5));
  nor2  gate2639(.a(gate139inter5), .b(gate139inter2), .O(gate139inter6));
  inv1  gate2640(.a(G438), .O(gate139inter7));
  inv1  gate2641(.a(G441), .O(gate139inter8));
  nand2 gate2642(.a(gate139inter8), .b(gate139inter7), .O(gate139inter9));
  nand2 gate2643(.a(s_299), .b(gate139inter3), .O(gate139inter10));
  nor2  gate2644(.a(gate139inter10), .b(gate139inter9), .O(gate139inter11));
  nor2  gate2645(.a(gate139inter11), .b(gate139inter6), .O(gate139inter12));
  nand2 gate2646(.a(gate139inter12), .b(gate139inter1), .O(G528));

  xor2  gate2437(.a(G447), .b(G444), .O(gate140inter0));
  nand2 gate2438(.a(gate140inter0), .b(s_270), .O(gate140inter1));
  and2  gate2439(.a(G447), .b(G444), .O(gate140inter2));
  inv1  gate2440(.a(s_270), .O(gate140inter3));
  inv1  gate2441(.a(s_271), .O(gate140inter4));
  nand2 gate2442(.a(gate140inter4), .b(gate140inter3), .O(gate140inter5));
  nor2  gate2443(.a(gate140inter5), .b(gate140inter2), .O(gate140inter6));
  inv1  gate2444(.a(G444), .O(gate140inter7));
  inv1  gate2445(.a(G447), .O(gate140inter8));
  nand2 gate2446(.a(gate140inter8), .b(gate140inter7), .O(gate140inter9));
  nand2 gate2447(.a(s_271), .b(gate140inter3), .O(gate140inter10));
  nor2  gate2448(.a(gate140inter10), .b(gate140inter9), .O(gate140inter11));
  nor2  gate2449(.a(gate140inter11), .b(gate140inter6), .O(gate140inter12));
  nand2 gate2450(.a(gate140inter12), .b(gate140inter1), .O(G531));

  xor2  gate659(.a(G453), .b(G450), .O(gate141inter0));
  nand2 gate660(.a(gate141inter0), .b(s_16), .O(gate141inter1));
  and2  gate661(.a(G453), .b(G450), .O(gate141inter2));
  inv1  gate662(.a(s_16), .O(gate141inter3));
  inv1  gate663(.a(s_17), .O(gate141inter4));
  nand2 gate664(.a(gate141inter4), .b(gate141inter3), .O(gate141inter5));
  nor2  gate665(.a(gate141inter5), .b(gate141inter2), .O(gate141inter6));
  inv1  gate666(.a(G450), .O(gate141inter7));
  inv1  gate667(.a(G453), .O(gate141inter8));
  nand2 gate668(.a(gate141inter8), .b(gate141inter7), .O(gate141inter9));
  nand2 gate669(.a(s_17), .b(gate141inter3), .O(gate141inter10));
  nor2  gate670(.a(gate141inter10), .b(gate141inter9), .O(gate141inter11));
  nor2  gate671(.a(gate141inter11), .b(gate141inter6), .O(gate141inter12));
  nand2 gate672(.a(gate141inter12), .b(gate141inter1), .O(G534));
nand2 gate142( .a(G456), .b(G459), .O(G537) );
nand2 gate143( .a(G462), .b(G465), .O(G540) );

  xor2  gate547(.a(G471), .b(G468), .O(gate144inter0));
  nand2 gate548(.a(gate144inter0), .b(s_0), .O(gate144inter1));
  and2  gate549(.a(G471), .b(G468), .O(gate144inter2));
  inv1  gate550(.a(s_0), .O(gate144inter3));
  inv1  gate551(.a(s_1), .O(gate144inter4));
  nand2 gate552(.a(gate144inter4), .b(gate144inter3), .O(gate144inter5));
  nor2  gate553(.a(gate144inter5), .b(gate144inter2), .O(gate144inter6));
  inv1  gate554(.a(G468), .O(gate144inter7));
  inv1  gate555(.a(G471), .O(gate144inter8));
  nand2 gate556(.a(gate144inter8), .b(gate144inter7), .O(gate144inter9));
  nand2 gate557(.a(s_1), .b(gate144inter3), .O(gate144inter10));
  nor2  gate558(.a(gate144inter10), .b(gate144inter9), .O(gate144inter11));
  nor2  gate559(.a(gate144inter11), .b(gate144inter6), .O(gate144inter12));
  nand2 gate560(.a(gate144inter12), .b(gate144inter1), .O(G543));
nand2 gate145( .a(G474), .b(G477), .O(G546) );
nand2 gate146( .a(G480), .b(G483), .O(G549) );
nand2 gate147( .a(G486), .b(G489), .O(G552) );
nand2 gate148( .a(G492), .b(G495), .O(G555) );

  xor2  gate939(.a(G501), .b(G498), .O(gate149inter0));
  nand2 gate940(.a(gate149inter0), .b(s_56), .O(gate149inter1));
  and2  gate941(.a(G501), .b(G498), .O(gate149inter2));
  inv1  gate942(.a(s_56), .O(gate149inter3));
  inv1  gate943(.a(s_57), .O(gate149inter4));
  nand2 gate944(.a(gate149inter4), .b(gate149inter3), .O(gate149inter5));
  nor2  gate945(.a(gate149inter5), .b(gate149inter2), .O(gate149inter6));
  inv1  gate946(.a(G498), .O(gate149inter7));
  inv1  gate947(.a(G501), .O(gate149inter8));
  nand2 gate948(.a(gate149inter8), .b(gate149inter7), .O(gate149inter9));
  nand2 gate949(.a(s_57), .b(gate149inter3), .O(gate149inter10));
  nor2  gate950(.a(gate149inter10), .b(gate149inter9), .O(gate149inter11));
  nor2  gate951(.a(gate149inter11), .b(gate149inter6), .O(gate149inter12));
  nand2 gate952(.a(gate149inter12), .b(gate149inter1), .O(G558));
nand2 gate150( .a(G504), .b(G507), .O(G561) );

  xor2  gate2451(.a(G513), .b(G510), .O(gate151inter0));
  nand2 gate2452(.a(gate151inter0), .b(s_272), .O(gate151inter1));
  and2  gate2453(.a(G513), .b(G510), .O(gate151inter2));
  inv1  gate2454(.a(s_272), .O(gate151inter3));
  inv1  gate2455(.a(s_273), .O(gate151inter4));
  nand2 gate2456(.a(gate151inter4), .b(gate151inter3), .O(gate151inter5));
  nor2  gate2457(.a(gate151inter5), .b(gate151inter2), .O(gate151inter6));
  inv1  gate2458(.a(G510), .O(gate151inter7));
  inv1  gate2459(.a(G513), .O(gate151inter8));
  nand2 gate2460(.a(gate151inter8), .b(gate151inter7), .O(gate151inter9));
  nand2 gate2461(.a(s_273), .b(gate151inter3), .O(gate151inter10));
  nor2  gate2462(.a(gate151inter10), .b(gate151inter9), .O(gate151inter11));
  nor2  gate2463(.a(gate151inter11), .b(gate151inter6), .O(gate151inter12));
  nand2 gate2464(.a(gate151inter12), .b(gate151inter1), .O(G564));
nand2 gate152( .a(G516), .b(G519), .O(G567) );
nand2 gate153( .a(G426), .b(G522), .O(G570) );
nand2 gate154( .a(G429), .b(G522), .O(G571) );

  xor2  gate1849(.a(G525), .b(G432), .O(gate155inter0));
  nand2 gate1850(.a(gate155inter0), .b(s_186), .O(gate155inter1));
  and2  gate1851(.a(G525), .b(G432), .O(gate155inter2));
  inv1  gate1852(.a(s_186), .O(gate155inter3));
  inv1  gate1853(.a(s_187), .O(gate155inter4));
  nand2 gate1854(.a(gate155inter4), .b(gate155inter3), .O(gate155inter5));
  nor2  gate1855(.a(gate155inter5), .b(gate155inter2), .O(gate155inter6));
  inv1  gate1856(.a(G432), .O(gate155inter7));
  inv1  gate1857(.a(G525), .O(gate155inter8));
  nand2 gate1858(.a(gate155inter8), .b(gate155inter7), .O(gate155inter9));
  nand2 gate1859(.a(s_187), .b(gate155inter3), .O(gate155inter10));
  nor2  gate1860(.a(gate155inter10), .b(gate155inter9), .O(gate155inter11));
  nor2  gate1861(.a(gate155inter11), .b(gate155inter6), .O(gate155inter12));
  nand2 gate1862(.a(gate155inter12), .b(gate155inter1), .O(G572));
nand2 gate156( .a(G435), .b(G525), .O(G573) );

  xor2  gate1933(.a(G528), .b(G438), .O(gate157inter0));
  nand2 gate1934(.a(gate157inter0), .b(s_198), .O(gate157inter1));
  and2  gate1935(.a(G528), .b(G438), .O(gate157inter2));
  inv1  gate1936(.a(s_198), .O(gate157inter3));
  inv1  gate1937(.a(s_199), .O(gate157inter4));
  nand2 gate1938(.a(gate157inter4), .b(gate157inter3), .O(gate157inter5));
  nor2  gate1939(.a(gate157inter5), .b(gate157inter2), .O(gate157inter6));
  inv1  gate1940(.a(G438), .O(gate157inter7));
  inv1  gate1941(.a(G528), .O(gate157inter8));
  nand2 gate1942(.a(gate157inter8), .b(gate157inter7), .O(gate157inter9));
  nand2 gate1943(.a(s_199), .b(gate157inter3), .O(gate157inter10));
  nor2  gate1944(.a(gate157inter10), .b(gate157inter9), .O(gate157inter11));
  nor2  gate1945(.a(gate157inter11), .b(gate157inter6), .O(gate157inter12));
  nand2 gate1946(.a(gate157inter12), .b(gate157inter1), .O(G574));

  xor2  gate1709(.a(G528), .b(G441), .O(gate158inter0));
  nand2 gate1710(.a(gate158inter0), .b(s_166), .O(gate158inter1));
  and2  gate1711(.a(G528), .b(G441), .O(gate158inter2));
  inv1  gate1712(.a(s_166), .O(gate158inter3));
  inv1  gate1713(.a(s_167), .O(gate158inter4));
  nand2 gate1714(.a(gate158inter4), .b(gate158inter3), .O(gate158inter5));
  nor2  gate1715(.a(gate158inter5), .b(gate158inter2), .O(gate158inter6));
  inv1  gate1716(.a(G441), .O(gate158inter7));
  inv1  gate1717(.a(G528), .O(gate158inter8));
  nand2 gate1718(.a(gate158inter8), .b(gate158inter7), .O(gate158inter9));
  nand2 gate1719(.a(s_167), .b(gate158inter3), .O(gate158inter10));
  nor2  gate1720(.a(gate158inter10), .b(gate158inter9), .O(gate158inter11));
  nor2  gate1721(.a(gate158inter11), .b(gate158inter6), .O(gate158inter12));
  nand2 gate1722(.a(gate158inter12), .b(gate158inter1), .O(G575));
nand2 gate159( .a(G444), .b(G531), .O(G576) );
nand2 gate160( .a(G447), .b(G531), .O(G577) );
nand2 gate161( .a(G450), .b(G534), .O(G578) );
nand2 gate162( .a(G453), .b(G534), .O(G579) );
nand2 gate163( .a(G456), .b(G537), .O(G580) );
nand2 gate164( .a(G459), .b(G537), .O(G581) );

  xor2  gate869(.a(G540), .b(G462), .O(gate165inter0));
  nand2 gate870(.a(gate165inter0), .b(s_46), .O(gate165inter1));
  and2  gate871(.a(G540), .b(G462), .O(gate165inter2));
  inv1  gate872(.a(s_46), .O(gate165inter3));
  inv1  gate873(.a(s_47), .O(gate165inter4));
  nand2 gate874(.a(gate165inter4), .b(gate165inter3), .O(gate165inter5));
  nor2  gate875(.a(gate165inter5), .b(gate165inter2), .O(gate165inter6));
  inv1  gate876(.a(G462), .O(gate165inter7));
  inv1  gate877(.a(G540), .O(gate165inter8));
  nand2 gate878(.a(gate165inter8), .b(gate165inter7), .O(gate165inter9));
  nand2 gate879(.a(s_47), .b(gate165inter3), .O(gate165inter10));
  nor2  gate880(.a(gate165inter10), .b(gate165inter9), .O(gate165inter11));
  nor2  gate881(.a(gate165inter11), .b(gate165inter6), .O(gate165inter12));
  nand2 gate882(.a(gate165inter12), .b(gate165inter1), .O(G582));
nand2 gate166( .a(G465), .b(G540), .O(G583) );
nand2 gate167( .a(G468), .b(G543), .O(G584) );

  xor2  gate2059(.a(G543), .b(G471), .O(gate168inter0));
  nand2 gate2060(.a(gate168inter0), .b(s_216), .O(gate168inter1));
  and2  gate2061(.a(G543), .b(G471), .O(gate168inter2));
  inv1  gate2062(.a(s_216), .O(gate168inter3));
  inv1  gate2063(.a(s_217), .O(gate168inter4));
  nand2 gate2064(.a(gate168inter4), .b(gate168inter3), .O(gate168inter5));
  nor2  gate2065(.a(gate168inter5), .b(gate168inter2), .O(gate168inter6));
  inv1  gate2066(.a(G471), .O(gate168inter7));
  inv1  gate2067(.a(G543), .O(gate168inter8));
  nand2 gate2068(.a(gate168inter8), .b(gate168inter7), .O(gate168inter9));
  nand2 gate2069(.a(s_217), .b(gate168inter3), .O(gate168inter10));
  nor2  gate2070(.a(gate168inter10), .b(gate168inter9), .O(gate168inter11));
  nor2  gate2071(.a(gate168inter11), .b(gate168inter6), .O(gate168inter12));
  nand2 gate2072(.a(gate168inter12), .b(gate168inter1), .O(G585));

  xor2  gate2577(.a(G546), .b(G474), .O(gate169inter0));
  nand2 gate2578(.a(gate169inter0), .b(s_290), .O(gate169inter1));
  and2  gate2579(.a(G546), .b(G474), .O(gate169inter2));
  inv1  gate2580(.a(s_290), .O(gate169inter3));
  inv1  gate2581(.a(s_291), .O(gate169inter4));
  nand2 gate2582(.a(gate169inter4), .b(gate169inter3), .O(gate169inter5));
  nor2  gate2583(.a(gate169inter5), .b(gate169inter2), .O(gate169inter6));
  inv1  gate2584(.a(G474), .O(gate169inter7));
  inv1  gate2585(.a(G546), .O(gate169inter8));
  nand2 gate2586(.a(gate169inter8), .b(gate169inter7), .O(gate169inter9));
  nand2 gate2587(.a(s_291), .b(gate169inter3), .O(gate169inter10));
  nor2  gate2588(.a(gate169inter10), .b(gate169inter9), .O(gate169inter11));
  nor2  gate2589(.a(gate169inter11), .b(gate169inter6), .O(gate169inter12));
  nand2 gate2590(.a(gate169inter12), .b(gate169inter1), .O(G586));
nand2 gate170( .a(G477), .b(G546), .O(G587) );
nand2 gate171( .a(G480), .b(G549), .O(G588) );

  xor2  gate2227(.a(G549), .b(G483), .O(gate172inter0));
  nand2 gate2228(.a(gate172inter0), .b(s_240), .O(gate172inter1));
  and2  gate2229(.a(G549), .b(G483), .O(gate172inter2));
  inv1  gate2230(.a(s_240), .O(gate172inter3));
  inv1  gate2231(.a(s_241), .O(gate172inter4));
  nand2 gate2232(.a(gate172inter4), .b(gate172inter3), .O(gate172inter5));
  nor2  gate2233(.a(gate172inter5), .b(gate172inter2), .O(gate172inter6));
  inv1  gate2234(.a(G483), .O(gate172inter7));
  inv1  gate2235(.a(G549), .O(gate172inter8));
  nand2 gate2236(.a(gate172inter8), .b(gate172inter7), .O(gate172inter9));
  nand2 gate2237(.a(s_241), .b(gate172inter3), .O(gate172inter10));
  nor2  gate2238(.a(gate172inter10), .b(gate172inter9), .O(gate172inter11));
  nor2  gate2239(.a(gate172inter11), .b(gate172inter6), .O(gate172inter12));
  nand2 gate2240(.a(gate172inter12), .b(gate172inter1), .O(G589));
nand2 gate173( .a(G486), .b(G552), .O(G590) );
nand2 gate174( .a(G489), .b(G552), .O(G591) );
nand2 gate175( .a(G492), .b(G555), .O(G592) );
nand2 gate176( .a(G495), .b(G555), .O(G593) );
nand2 gate177( .a(G498), .b(G558), .O(G594) );

  xor2  gate1639(.a(G558), .b(G501), .O(gate178inter0));
  nand2 gate1640(.a(gate178inter0), .b(s_156), .O(gate178inter1));
  and2  gate1641(.a(G558), .b(G501), .O(gate178inter2));
  inv1  gate1642(.a(s_156), .O(gate178inter3));
  inv1  gate1643(.a(s_157), .O(gate178inter4));
  nand2 gate1644(.a(gate178inter4), .b(gate178inter3), .O(gate178inter5));
  nor2  gate1645(.a(gate178inter5), .b(gate178inter2), .O(gate178inter6));
  inv1  gate1646(.a(G501), .O(gate178inter7));
  inv1  gate1647(.a(G558), .O(gate178inter8));
  nand2 gate1648(.a(gate178inter8), .b(gate178inter7), .O(gate178inter9));
  nand2 gate1649(.a(s_157), .b(gate178inter3), .O(gate178inter10));
  nor2  gate1650(.a(gate178inter10), .b(gate178inter9), .O(gate178inter11));
  nor2  gate1651(.a(gate178inter11), .b(gate178inter6), .O(gate178inter12));
  nand2 gate1652(.a(gate178inter12), .b(gate178inter1), .O(G595));
nand2 gate179( .a(G504), .b(G561), .O(G596) );
nand2 gate180( .a(G507), .b(G561), .O(G597) );

  xor2  gate1653(.a(G564), .b(G510), .O(gate181inter0));
  nand2 gate1654(.a(gate181inter0), .b(s_158), .O(gate181inter1));
  and2  gate1655(.a(G564), .b(G510), .O(gate181inter2));
  inv1  gate1656(.a(s_158), .O(gate181inter3));
  inv1  gate1657(.a(s_159), .O(gate181inter4));
  nand2 gate1658(.a(gate181inter4), .b(gate181inter3), .O(gate181inter5));
  nor2  gate1659(.a(gate181inter5), .b(gate181inter2), .O(gate181inter6));
  inv1  gate1660(.a(G510), .O(gate181inter7));
  inv1  gate1661(.a(G564), .O(gate181inter8));
  nand2 gate1662(.a(gate181inter8), .b(gate181inter7), .O(gate181inter9));
  nand2 gate1663(.a(s_159), .b(gate181inter3), .O(gate181inter10));
  nor2  gate1664(.a(gate181inter10), .b(gate181inter9), .O(gate181inter11));
  nor2  gate1665(.a(gate181inter11), .b(gate181inter6), .O(gate181inter12));
  nand2 gate1666(.a(gate181inter12), .b(gate181inter1), .O(G598));
nand2 gate182( .a(G513), .b(G564), .O(G599) );
nand2 gate183( .a(G516), .b(G567), .O(G600) );

  xor2  gate2199(.a(G567), .b(G519), .O(gate184inter0));
  nand2 gate2200(.a(gate184inter0), .b(s_236), .O(gate184inter1));
  and2  gate2201(.a(G567), .b(G519), .O(gate184inter2));
  inv1  gate2202(.a(s_236), .O(gate184inter3));
  inv1  gate2203(.a(s_237), .O(gate184inter4));
  nand2 gate2204(.a(gate184inter4), .b(gate184inter3), .O(gate184inter5));
  nor2  gate2205(.a(gate184inter5), .b(gate184inter2), .O(gate184inter6));
  inv1  gate2206(.a(G519), .O(gate184inter7));
  inv1  gate2207(.a(G567), .O(gate184inter8));
  nand2 gate2208(.a(gate184inter8), .b(gate184inter7), .O(gate184inter9));
  nand2 gate2209(.a(s_237), .b(gate184inter3), .O(gate184inter10));
  nor2  gate2210(.a(gate184inter10), .b(gate184inter9), .O(gate184inter11));
  nor2  gate2211(.a(gate184inter11), .b(gate184inter6), .O(gate184inter12));
  nand2 gate2212(.a(gate184inter12), .b(gate184inter1), .O(G601));
nand2 gate185( .a(G570), .b(G571), .O(G602) );

  xor2  gate2143(.a(G573), .b(G572), .O(gate186inter0));
  nand2 gate2144(.a(gate186inter0), .b(s_228), .O(gate186inter1));
  and2  gate2145(.a(G573), .b(G572), .O(gate186inter2));
  inv1  gate2146(.a(s_228), .O(gate186inter3));
  inv1  gate2147(.a(s_229), .O(gate186inter4));
  nand2 gate2148(.a(gate186inter4), .b(gate186inter3), .O(gate186inter5));
  nor2  gate2149(.a(gate186inter5), .b(gate186inter2), .O(gate186inter6));
  inv1  gate2150(.a(G572), .O(gate186inter7));
  inv1  gate2151(.a(G573), .O(gate186inter8));
  nand2 gate2152(.a(gate186inter8), .b(gate186inter7), .O(gate186inter9));
  nand2 gate2153(.a(s_229), .b(gate186inter3), .O(gate186inter10));
  nor2  gate2154(.a(gate186inter10), .b(gate186inter9), .O(gate186inter11));
  nor2  gate2155(.a(gate186inter11), .b(gate186inter6), .O(gate186inter12));
  nand2 gate2156(.a(gate186inter12), .b(gate186inter1), .O(G607));
nand2 gate187( .a(G574), .b(G575), .O(G612) );

  xor2  gate2129(.a(G577), .b(G576), .O(gate188inter0));
  nand2 gate2130(.a(gate188inter0), .b(s_226), .O(gate188inter1));
  and2  gate2131(.a(G577), .b(G576), .O(gate188inter2));
  inv1  gate2132(.a(s_226), .O(gate188inter3));
  inv1  gate2133(.a(s_227), .O(gate188inter4));
  nand2 gate2134(.a(gate188inter4), .b(gate188inter3), .O(gate188inter5));
  nor2  gate2135(.a(gate188inter5), .b(gate188inter2), .O(gate188inter6));
  inv1  gate2136(.a(G576), .O(gate188inter7));
  inv1  gate2137(.a(G577), .O(gate188inter8));
  nand2 gate2138(.a(gate188inter8), .b(gate188inter7), .O(gate188inter9));
  nand2 gate2139(.a(s_227), .b(gate188inter3), .O(gate188inter10));
  nor2  gate2140(.a(gate188inter10), .b(gate188inter9), .O(gate188inter11));
  nor2  gate2141(.a(gate188inter11), .b(gate188inter6), .O(gate188inter12));
  nand2 gate2142(.a(gate188inter12), .b(gate188inter1), .O(G617));

  xor2  gate855(.a(G579), .b(G578), .O(gate189inter0));
  nand2 gate856(.a(gate189inter0), .b(s_44), .O(gate189inter1));
  and2  gate857(.a(G579), .b(G578), .O(gate189inter2));
  inv1  gate858(.a(s_44), .O(gate189inter3));
  inv1  gate859(.a(s_45), .O(gate189inter4));
  nand2 gate860(.a(gate189inter4), .b(gate189inter3), .O(gate189inter5));
  nor2  gate861(.a(gate189inter5), .b(gate189inter2), .O(gate189inter6));
  inv1  gate862(.a(G578), .O(gate189inter7));
  inv1  gate863(.a(G579), .O(gate189inter8));
  nand2 gate864(.a(gate189inter8), .b(gate189inter7), .O(gate189inter9));
  nand2 gate865(.a(s_45), .b(gate189inter3), .O(gate189inter10));
  nor2  gate866(.a(gate189inter10), .b(gate189inter9), .O(gate189inter11));
  nor2  gate867(.a(gate189inter11), .b(gate189inter6), .O(gate189inter12));
  nand2 gate868(.a(gate189inter12), .b(gate189inter1), .O(G622));
nand2 gate190( .a(G580), .b(G581), .O(G627) );
nand2 gate191( .a(G582), .b(G583), .O(G632) );

  xor2  gate1793(.a(G585), .b(G584), .O(gate192inter0));
  nand2 gate1794(.a(gate192inter0), .b(s_178), .O(gate192inter1));
  and2  gate1795(.a(G585), .b(G584), .O(gate192inter2));
  inv1  gate1796(.a(s_178), .O(gate192inter3));
  inv1  gate1797(.a(s_179), .O(gate192inter4));
  nand2 gate1798(.a(gate192inter4), .b(gate192inter3), .O(gate192inter5));
  nor2  gate1799(.a(gate192inter5), .b(gate192inter2), .O(gate192inter6));
  inv1  gate1800(.a(G584), .O(gate192inter7));
  inv1  gate1801(.a(G585), .O(gate192inter8));
  nand2 gate1802(.a(gate192inter8), .b(gate192inter7), .O(gate192inter9));
  nand2 gate1803(.a(s_179), .b(gate192inter3), .O(gate192inter10));
  nor2  gate1804(.a(gate192inter10), .b(gate192inter9), .O(gate192inter11));
  nor2  gate1805(.a(gate192inter11), .b(gate192inter6), .O(gate192inter12));
  nand2 gate1806(.a(gate192inter12), .b(gate192inter1), .O(G637));
nand2 gate193( .a(G586), .b(G587), .O(G642) );

  xor2  gate1863(.a(G589), .b(G588), .O(gate194inter0));
  nand2 gate1864(.a(gate194inter0), .b(s_188), .O(gate194inter1));
  and2  gate1865(.a(G589), .b(G588), .O(gate194inter2));
  inv1  gate1866(.a(s_188), .O(gate194inter3));
  inv1  gate1867(.a(s_189), .O(gate194inter4));
  nand2 gate1868(.a(gate194inter4), .b(gate194inter3), .O(gate194inter5));
  nor2  gate1869(.a(gate194inter5), .b(gate194inter2), .O(gate194inter6));
  inv1  gate1870(.a(G588), .O(gate194inter7));
  inv1  gate1871(.a(G589), .O(gate194inter8));
  nand2 gate1872(.a(gate194inter8), .b(gate194inter7), .O(gate194inter9));
  nand2 gate1873(.a(s_189), .b(gate194inter3), .O(gate194inter10));
  nor2  gate1874(.a(gate194inter10), .b(gate194inter9), .O(gate194inter11));
  nor2  gate1875(.a(gate194inter11), .b(gate194inter6), .O(gate194inter12));
  nand2 gate1876(.a(gate194inter12), .b(gate194inter1), .O(G645));

  xor2  gate2213(.a(G591), .b(G590), .O(gate195inter0));
  nand2 gate2214(.a(gate195inter0), .b(s_238), .O(gate195inter1));
  and2  gate2215(.a(G591), .b(G590), .O(gate195inter2));
  inv1  gate2216(.a(s_238), .O(gate195inter3));
  inv1  gate2217(.a(s_239), .O(gate195inter4));
  nand2 gate2218(.a(gate195inter4), .b(gate195inter3), .O(gate195inter5));
  nor2  gate2219(.a(gate195inter5), .b(gate195inter2), .O(gate195inter6));
  inv1  gate2220(.a(G590), .O(gate195inter7));
  inv1  gate2221(.a(G591), .O(gate195inter8));
  nand2 gate2222(.a(gate195inter8), .b(gate195inter7), .O(gate195inter9));
  nand2 gate2223(.a(s_239), .b(gate195inter3), .O(gate195inter10));
  nor2  gate2224(.a(gate195inter10), .b(gate195inter9), .O(gate195inter11));
  nor2  gate2225(.a(gate195inter11), .b(gate195inter6), .O(gate195inter12));
  nand2 gate2226(.a(gate195inter12), .b(gate195inter1), .O(G648));

  xor2  gate2507(.a(G593), .b(G592), .O(gate196inter0));
  nand2 gate2508(.a(gate196inter0), .b(s_280), .O(gate196inter1));
  and2  gate2509(.a(G593), .b(G592), .O(gate196inter2));
  inv1  gate2510(.a(s_280), .O(gate196inter3));
  inv1  gate2511(.a(s_281), .O(gate196inter4));
  nand2 gate2512(.a(gate196inter4), .b(gate196inter3), .O(gate196inter5));
  nor2  gate2513(.a(gate196inter5), .b(gate196inter2), .O(gate196inter6));
  inv1  gate2514(.a(G592), .O(gate196inter7));
  inv1  gate2515(.a(G593), .O(gate196inter8));
  nand2 gate2516(.a(gate196inter8), .b(gate196inter7), .O(gate196inter9));
  nand2 gate2517(.a(s_281), .b(gate196inter3), .O(gate196inter10));
  nor2  gate2518(.a(gate196inter10), .b(gate196inter9), .O(gate196inter11));
  nor2  gate2519(.a(gate196inter11), .b(gate196inter6), .O(gate196inter12));
  nand2 gate2520(.a(gate196inter12), .b(gate196inter1), .O(G651));
nand2 gate197( .a(G594), .b(G595), .O(G654) );
nand2 gate198( .a(G596), .b(G597), .O(G657) );
nand2 gate199( .a(G598), .b(G599), .O(G660) );
nand2 gate200( .a(G600), .b(G601), .O(G663) );
nand2 gate201( .a(G602), .b(G607), .O(G666) );
nand2 gate202( .a(G612), .b(G617), .O(G669) );
nand2 gate203( .a(G602), .b(G612), .O(G672) );
nand2 gate204( .a(G607), .b(G617), .O(G675) );

  xor2  gate799(.a(G627), .b(G622), .O(gate205inter0));
  nand2 gate800(.a(gate205inter0), .b(s_36), .O(gate205inter1));
  and2  gate801(.a(G627), .b(G622), .O(gate205inter2));
  inv1  gate802(.a(s_36), .O(gate205inter3));
  inv1  gate803(.a(s_37), .O(gate205inter4));
  nand2 gate804(.a(gate205inter4), .b(gate205inter3), .O(gate205inter5));
  nor2  gate805(.a(gate205inter5), .b(gate205inter2), .O(gate205inter6));
  inv1  gate806(.a(G622), .O(gate205inter7));
  inv1  gate807(.a(G627), .O(gate205inter8));
  nand2 gate808(.a(gate205inter8), .b(gate205inter7), .O(gate205inter9));
  nand2 gate809(.a(s_37), .b(gate205inter3), .O(gate205inter10));
  nor2  gate810(.a(gate205inter10), .b(gate205inter9), .O(gate205inter11));
  nor2  gate811(.a(gate205inter11), .b(gate205inter6), .O(gate205inter12));
  nand2 gate812(.a(gate205inter12), .b(gate205inter1), .O(G678));

  xor2  gate1303(.a(G637), .b(G632), .O(gate206inter0));
  nand2 gate1304(.a(gate206inter0), .b(s_108), .O(gate206inter1));
  and2  gate1305(.a(G637), .b(G632), .O(gate206inter2));
  inv1  gate1306(.a(s_108), .O(gate206inter3));
  inv1  gate1307(.a(s_109), .O(gate206inter4));
  nand2 gate1308(.a(gate206inter4), .b(gate206inter3), .O(gate206inter5));
  nor2  gate1309(.a(gate206inter5), .b(gate206inter2), .O(gate206inter6));
  inv1  gate1310(.a(G632), .O(gate206inter7));
  inv1  gate1311(.a(G637), .O(gate206inter8));
  nand2 gate1312(.a(gate206inter8), .b(gate206inter7), .O(gate206inter9));
  nand2 gate1313(.a(s_109), .b(gate206inter3), .O(gate206inter10));
  nor2  gate1314(.a(gate206inter10), .b(gate206inter9), .O(gate206inter11));
  nor2  gate1315(.a(gate206inter11), .b(gate206inter6), .O(gate206inter12));
  nand2 gate1316(.a(gate206inter12), .b(gate206inter1), .O(G681));
nand2 gate207( .a(G622), .b(G632), .O(G684) );
nand2 gate208( .a(G627), .b(G637), .O(G687) );
nand2 gate209( .a(G602), .b(G666), .O(G690) );
nand2 gate210( .a(G607), .b(G666), .O(G691) );

  xor2  gate1093(.a(G669), .b(G612), .O(gate211inter0));
  nand2 gate1094(.a(gate211inter0), .b(s_78), .O(gate211inter1));
  and2  gate1095(.a(G669), .b(G612), .O(gate211inter2));
  inv1  gate1096(.a(s_78), .O(gate211inter3));
  inv1  gate1097(.a(s_79), .O(gate211inter4));
  nand2 gate1098(.a(gate211inter4), .b(gate211inter3), .O(gate211inter5));
  nor2  gate1099(.a(gate211inter5), .b(gate211inter2), .O(gate211inter6));
  inv1  gate1100(.a(G612), .O(gate211inter7));
  inv1  gate1101(.a(G669), .O(gate211inter8));
  nand2 gate1102(.a(gate211inter8), .b(gate211inter7), .O(gate211inter9));
  nand2 gate1103(.a(s_79), .b(gate211inter3), .O(gate211inter10));
  nor2  gate1104(.a(gate211inter10), .b(gate211inter9), .O(gate211inter11));
  nor2  gate1105(.a(gate211inter11), .b(gate211inter6), .O(gate211inter12));
  nand2 gate1106(.a(gate211inter12), .b(gate211inter1), .O(G692));

  xor2  gate589(.a(G669), .b(G617), .O(gate212inter0));
  nand2 gate590(.a(gate212inter0), .b(s_6), .O(gate212inter1));
  and2  gate591(.a(G669), .b(G617), .O(gate212inter2));
  inv1  gate592(.a(s_6), .O(gate212inter3));
  inv1  gate593(.a(s_7), .O(gate212inter4));
  nand2 gate594(.a(gate212inter4), .b(gate212inter3), .O(gate212inter5));
  nor2  gate595(.a(gate212inter5), .b(gate212inter2), .O(gate212inter6));
  inv1  gate596(.a(G617), .O(gate212inter7));
  inv1  gate597(.a(G669), .O(gate212inter8));
  nand2 gate598(.a(gate212inter8), .b(gate212inter7), .O(gate212inter9));
  nand2 gate599(.a(s_7), .b(gate212inter3), .O(gate212inter10));
  nor2  gate600(.a(gate212inter10), .b(gate212inter9), .O(gate212inter11));
  nor2  gate601(.a(gate212inter11), .b(gate212inter6), .O(gate212inter12));
  nand2 gate602(.a(gate212inter12), .b(gate212inter1), .O(G693));

  xor2  gate1191(.a(G672), .b(G602), .O(gate213inter0));
  nand2 gate1192(.a(gate213inter0), .b(s_92), .O(gate213inter1));
  and2  gate1193(.a(G672), .b(G602), .O(gate213inter2));
  inv1  gate1194(.a(s_92), .O(gate213inter3));
  inv1  gate1195(.a(s_93), .O(gate213inter4));
  nand2 gate1196(.a(gate213inter4), .b(gate213inter3), .O(gate213inter5));
  nor2  gate1197(.a(gate213inter5), .b(gate213inter2), .O(gate213inter6));
  inv1  gate1198(.a(G602), .O(gate213inter7));
  inv1  gate1199(.a(G672), .O(gate213inter8));
  nand2 gate1200(.a(gate213inter8), .b(gate213inter7), .O(gate213inter9));
  nand2 gate1201(.a(s_93), .b(gate213inter3), .O(gate213inter10));
  nor2  gate1202(.a(gate213inter10), .b(gate213inter9), .O(gate213inter11));
  nor2  gate1203(.a(gate213inter11), .b(gate213inter6), .O(gate213inter12));
  nand2 gate1204(.a(gate213inter12), .b(gate213inter1), .O(G694));
nand2 gate214( .a(G612), .b(G672), .O(G695) );
nand2 gate215( .a(G607), .b(G675), .O(G696) );

  xor2  gate1121(.a(G675), .b(G617), .O(gate216inter0));
  nand2 gate1122(.a(gate216inter0), .b(s_82), .O(gate216inter1));
  and2  gate1123(.a(G675), .b(G617), .O(gate216inter2));
  inv1  gate1124(.a(s_82), .O(gate216inter3));
  inv1  gate1125(.a(s_83), .O(gate216inter4));
  nand2 gate1126(.a(gate216inter4), .b(gate216inter3), .O(gate216inter5));
  nor2  gate1127(.a(gate216inter5), .b(gate216inter2), .O(gate216inter6));
  inv1  gate1128(.a(G617), .O(gate216inter7));
  inv1  gate1129(.a(G675), .O(gate216inter8));
  nand2 gate1130(.a(gate216inter8), .b(gate216inter7), .O(gate216inter9));
  nand2 gate1131(.a(s_83), .b(gate216inter3), .O(gate216inter10));
  nor2  gate1132(.a(gate216inter10), .b(gate216inter9), .O(gate216inter11));
  nor2  gate1133(.a(gate216inter11), .b(gate216inter6), .O(gate216inter12));
  nand2 gate1134(.a(gate216inter12), .b(gate216inter1), .O(G697));
nand2 gate217( .a(G622), .b(G678), .O(G698) );
nand2 gate218( .a(G627), .b(G678), .O(G699) );
nand2 gate219( .a(G632), .b(G681), .O(G700) );
nand2 gate220( .a(G637), .b(G681), .O(G701) );

  xor2  gate897(.a(G684), .b(G622), .O(gate221inter0));
  nand2 gate898(.a(gate221inter0), .b(s_50), .O(gate221inter1));
  and2  gate899(.a(G684), .b(G622), .O(gate221inter2));
  inv1  gate900(.a(s_50), .O(gate221inter3));
  inv1  gate901(.a(s_51), .O(gate221inter4));
  nand2 gate902(.a(gate221inter4), .b(gate221inter3), .O(gate221inter5));
  nor2  gate903(.a(gate221inter5), .b(gate221inter2), .O(gate221inter6));
  inv1  gate904(.a(G622), .O(gate221inter7));
  inv1  gate905(.a(G684), .O(gate221inter8));
  nand2 gate906(.a(gate221inter8), .b(gate221inter7), .O(gate221inter9));
  nand2 gate907(.a(s_51), .b(gate221inter3), .O(gate221inter10));
  nor2  gate908(.a(gate221inter10), .b(gate221inter9), .O(gate221inter11));
  nor2  gate909(.a(gate221inter11), .b(gate221inter6), .O(gate221inter12));
  nand2 gate910(.a(gate221inter12), .b(gate221inter1), .O(G702));
nand2 gate222( .a(G632), .b(G684), .O(G703) );

  xor2  gate841(.a(G687), .b(G627), .O(gate223inter0));
  nand2 gate842(.a(gate223inter0), .b(s_42), .O(gate223inter1));
  and2  gate843(.a(G687), .b(G627), .O(gate223inter2));
  inv1  gate844(.a(s_42), .O(gate223inter3));
  inv1  gate845(.a(s_43), .O(gate223inter4));
  nand2 gate846(.a(gate223inter4), .b(gate223inter3), .O(gate223inter5));
  nor2  gate847(.a(gate223inter5), .b(gate223inter2), .O(gate223inter6));
  inv1  gate848(.a(G627), .O(gate223inter7));
  inv1  gate849(.a(G687), .O(gate223inter8));
  nand2 gate850(.a(gate223inter8), .b(gate223inter7), .O(gate223inter9));
  nand2 gate851(.a(s_43), .b(gate223inter3), .O(gate223inter10));
  nor2  gate852(.a(gate223inter10), .b(gate223inter9), .O(gate223inter11));
  nor2  gate853(.a(gate223inter11), .b(gate223inter6), .O(gate223inter12));
  nand2 gate854(.a(gate223inter12), .b(gate223inter1), .O(G704));
nand2 gate224( .a(G637), .b(G687), .O(G705) );
nand2 gate225( .a(G690), .b(G691), .O(G706) );
nand2 gate226( .a(G692), .b(G693), .O(G709) );

  xor2  gate1947(.a(G695), .b(G694), .O(gate227inter0));
  nand2 gate1948(.a(gate227inter0), .b(s_200), .O(gate227inter1));
  and2  gate1949(.a(G695), .b(G694), .O(gate227inter2));
  inv1  gate1950(.a(s_200), .O(gate227inter3));
  inv1  gate1951(.a(s_201), .O(gate227inter4));
  nand2 gate1952(.a(gate227inter4), .b(gate227inter3), .O(gate227inter5));
  nor2  gate1953(.a(gate227inter5), .b(gate227inter2), .O(gate227inter6));
  inv1  gate1954(.a(G694), .O(gate227inter7));
  inv1  gate1955(.a(G695), .O(gate227inter8));
  nand2 gate1956(.a(gate227inter8), .b(gate227inter7), .O(gate227inter9));
  nand2 gate1957(.a(s_201), .b(gate227inter3), .O(gate227inter10));
  nor2  gate1958(.a(gate227inter10), .b(gate227inter9), .O(gate227inter11));
  nor2  gate1959(.a(gate227inter11), .b(gate227inter6), .O(gate227inter12));
  nand2 gate1960(.a(gate227inter12), .b(gate227inter1), .O(G712));

  xor2  gate1821(.a(G697), .b(G696), .O(gate228inter0));
  nand2 gate1822(.a(gate228inter0), .b(s_182), .O(gate228inter1));
  and2  gate1823(.a(G697), .b(G696), .O(gate228inter2));
  inv1  gate1824(.a(s_182), .O(gate228inter3));
  inv1  gate1825(.a(s_183), .O(gate228inter4));
  nand2 gate1826(.a(gate228inter4), .b(gate228inter3), .O(gate228inter5));
  nor2  gate1827(.a(gate228inter5), .b(gate228inter2), .O(gate228inter6));
  inv1  gate1828(.a(G696), .O(gate228inter7));
  inv1  gate1829(.a(G697), .O(gate228inter8));
  nand2 gate1830(.a(gate228inter8), .b(gate228inter7), .O(gate228inter9));
  nand2 gate1831(.a(s_183), .b(gate228inter3), .O(gate228inter10));
  nor2  gate1832(.a(gate228inter10), .b(gate228inter9), .O(gate228inter11));
  nor2  gate1833(.a(gate228inter11), .b(gate228inter6), .O(gate228inter12));
  nand2 gate1834(.a(gate228inter12), .b(gate228inter1), .O(G715));
nand2 gate229( .a(G698), .b(G699), .O(G718) );
nand2 gate230( .a(G700), .b(G701), .O(G721) );
nand2 gate231( .a(G702), .b(G703), .O(G724) );
nand2 gate232( .a(G704), .b(G705), .O(G727) );
nand2 gate233( .a(G242), .b(G718), .O(G730) );

  xor2  gate1429(.a(G721), .b(G245), .O(gate234inter0));
  nand2 gate1430(.a(gate234inter0), .b(s_126), .O(gate234inter1));
  and2  gate1431(.a(G721), .b(G245), .O(gate234inter2));
  inv1  gate1432(.a(s_126), .O(gate234inter3));
  inv1  gate1433(.a(s_127), .O(gate234inter4));
  nand2 gate1434(.a(gate234inter4), .b(gate234inter3), .O(gate234inter5));
  nor2  gate1435(.a(gate234inter5), .b(gate234inter2), .O(gate234inter6));
  inv1  gate1436(.a(G245), .O(gate234inter7));
  inv1  gate1437(.a(G721), .O(gate234inter8));
  nand2 gate1438(.a(gate234inter8), .b(gate234inter7), .O(gate234inter9));
  nand2 gate1439(.a(s_127), .b(gate234inter3), .O(gate234inter10));
  nor2  gate1440(.a(gate234inter10), .b(gate234inter9), .O(gate234inter11));
  nor2  gate1441(.a(gate234inter11), .b(gate234inter6), .O(gate234inter12));
  nand2 gate1442(.a(gate234inter12), .b(gate234inter1), .O(G733));
nand2 gate235( .a(G248), .b(G724), .O(G736) );
nand2 gate236( .a(G251), .b(G727), .O(G739) );
nand2 gate237( .a(G254), .b(G706), .O(G742) );
nand2 gate238( .a(G257), .b(G709), .O(G745) );
nand2 gate239( .a(G260), .b(G712), .O(G748) );
nand2 gate240( .a(G263), .b(G715), .O(G751) );
nand2 gate241( .a(G242), .b(G730), .O(G754) );
nand2 gate242( .a(G718), .b(G730), .O(G755) );
nand2 gate243( .a(G245), .b(G733), .O(G756) );
nand2 gate244( .a(G721), .b(G733), .O(G757) );
nand2 gate245( .a(G248), .b(G736), .O(G758) );
nand2 gate246( .a(G724), .b(G736), .O(G759) );
nand2 gate247( .a(G251), .b(G739), .O(G760) );
nand2 gate248( .a(G727), .b(G739), .O(G761) );
nand2 gate249( .a(G254), .b(G742), .O(G762) );
nand2 gate250( .a(G706), .b(G742), .O(G763) );

  xor2  gate1681(.a(G745), .b(G257), .O(gate251inter0));
  nand2 gate1682(.a(gate251inter0), .b(s_162), .O(gate251inter1));
  and2  gate1683(.a(G745), .b(G257), .O(gate251inter2));
  inv1  gate1684(.a(s_162), .O(gate251inter3));
  inv1  gate1685(.a(s_163), .O(gate251inter4));
  nand2 gate1686(.a(gate251inter4), .b(gate251inter3), .O(gate251inter5));
  nor2  gate1687(.a(gate251inter5), .b(gate251inter2), .O(gate251inter6));
  inv1  gate1688(.a(G257), .O(gate251inter7));
  inv1  gate1689(.a(G745), .O(gate251inter8));
  nand2 gate1690(.a(gate251inter8), .b(gate251inter7), .O(gate251inter9));
  nand2 gate1691(.a(s_163), .b(gate251inter3), .O(gate251inter10));
  nor2  gate1692(.a(gate251inter10), .b(gate251inter9), .O(gate251inter11));
  nor2  gate1693(.a(gate251inter11), .b(gate251inter6), .O(gate251inter12));
  nand2 gate1694(.a(gate251inter12), .b(gate251inter1), .O(G764));

  xor2  gate1401(.a(G745), .b(G709), .O(gate252inter0));
  nand2 gate1402(.a(gate252inter0), .b(s_122), .O(gate252inter1));
  and2  gate1403(.a(G745), .b(G709), .O(gate252inter2));
  inv1  gate1404(.a(s_122), .O(gate252inter3));
  inv1  gate1405(.a(s_123), .O(gate252inter4));
  nand2 gate1406(.a(gate252inter4), .b(gate252inter3), .O(gate252inter5));
  nor2  gate1407(.a(gate252inter5), .b(gate252inter2), .O(gate252inter6));
  inv1  gate1408(.a(G709), .O(gate252inter7));
  inv1  gate1409(.a(G745), .O(gate252inter8));
  nand2 gate1410(.a(gate252inter8), .b(gate252inter7), .O(gate252inter9));
  nand2 gate1411(.a(s_123), .b(gate252inter3), .O(gate252inter10));
  nor2  gate1412(.a(gate252inter10), .b(gate252inter9), .O(gate252inter11));
  nor2  gate1413(.a(gate252inter11), .b(gate252inter6), .O(gate252inter12));
  nand2 gate1414(.a(gate252inter12), .b(gate252inter1), .O(G765));
nand2 gate253( .a(G260), .b(G748), .O(G766) );
nand2 gate254( .a(G712), .b(G748), .O(G767) );

  xor2  gate1695(.a(G751), .b(G263), .O(gate255inter0));
  nand2 gate1696(.a(gate255inter0), .b(s_164), .O(gate255inter1));
  and2  gate1697(.a(G751), .b(G263), .O(gate255inter2));
  inv1  gate1698(.a(s_164), .O(gate255inter3));
  inv1  gate1699(.a(s_165), .O(gate255inter4));
  nand2 gate1700(.a(gate255inter4), .b(gate255inter3), .O(gate255inter5));
  nor2  gate1701(.a(gate255inter5), .b(gate255inter2), .O(gate255inter6));
  inv1  gate1702(.a(G263), .O(gate255inter7));
  inv1  gate1703(.a(G751), .O(gate255inter8));
  nand2 gate1704(.a(gate255inter8), .b(gate255inter7), .O(gate255inter9));
  nand2 gate1705(.a(s_165), .b(gate255inter3), .O(gate255inter10));
  nor2  gate1706(.a(gate255inter10), .b(gate255inter9), .O(gate255inter11));
  nor2  gate1707(.a(gate255inter11), .b(gate255inter6), .O(gate255inter12));
  nand2 gate1708(.a(gate255inter12), .b(gate255inter1), .O(G768));
nand2 gate256( .a(G715), .b(G751), .O(G769) );

  xor2  gate1415(.a(G755), .b(G754), .O(gate257inter0));
  nand2 gate1416(.a(gate257inter0), .b(s_124), .O(gate257inter1));
  and2  gate1417(.a(G755), .b(G754), .O(gate257inter2));
  inv1  gate1418(.a(s_124), .O(gate257inter3));
  inv1  gate1419(.a(s_125), .O(gate257inter4));
  nand2 gate1420(.a(gate257inter4), .b(gate257inter3), .O(gate257inter5));
  nor2  gate1421(.a(gate257inter5), .b(gate257inter2), .O(gate257inter6));
  inv1  gate1422(.a(G754), .O(gate257inter7));
  inv1  gate1423(.a(G755), .O(gate257inter8));
  nand2 gate1424(.a(gate257inter8), .b(gate257inter7), .O(gate257inter9));
  nand2 gate1425(.a(s_125), .b(gate257inter3), .O(gate257inter10));
  nor2  gate1426(.a(gate257inter10), .b(gate257inter9), .O(gate257inter11));
  nor2  gate1427(.a(gate257inter11), .b(gate257inter6), .O(gate257inter12));
  nand2 gate1428(.a(gate257inter12), .b(gate257inter1), .O(G770));
nand2 gate258( .a(G756), .b(G757), .O(G773) );
nand2 gate259( .a(G758), .b(G759), .O(G776) );

  xor2  gate1597(.a(G761), .b(G760), .O(gate260inter0));
  nand2 gate1598(.a(gate260inter0), .b(s_150), .O(gate260inter1));
  and2  gate1599(.a(G761), .b(G760), .O(gate260inter2));
  inv1  gate1600(.a(s_150), .O(gate260inter3));
  inv1  gate1601(.a(s_151), .O(gate260inter4));
  nand2 gate1602(.a(gate260inter4), .b(gate260inter3), .O(gate260inter5));
  nor2  gate1603(.a(gate260inter5), .b(gate260inter2), .O(gate260inter6));
  inv1  gate1604(.a(G760), .O(gate260inter7));
  inv1  gate1605(.a(G761), .O(gate260inter8));
  nand2 gate1606(.a(gate260inter8), .b(gate260inter7), .O(gate260inter9));
  nand2 gate1607(.a(s_151), .b(gate260inter3), .O(gate260inter10));
  nor2  gate1608(.a(gate260inter10), .b(gate260inter9), .O(gate260inter11));
  nor2  gate1609(.a(gate260inter11), .b(gate260inter6), .O(gate260inter12));
  nand2 gate1610(.a(gate260inter12), .b(gate260inter1), .O(G779));
nand2 gate261( .a(G762), .b(G763), .O(G782) );
nand2 gate262( .a(G764), .b(G765), .O(G785) );
nand2 gate263( .a(G766), .b(G767), .O(G788) );
nand2 gate264( .a(G768), .b(G769), .O(G791) );

  xor2  gate2297(.a(G770), .b(G642), .O(gate265inter0));
  nand2 gate2298(.a(gate265inter0), .b(s_250), .O(gate265inter1));
  and2  gate2299(.a(G770), .b(G642), .O(gate265inter2));
  inv1  gate2300(.a(s_250), .O(gate265inter3));
  inv1  gate2301(.a(s_251), .O(gate265inter4));
  nand2 gate2302(.a(gate265inter4), .b(gate265inter3), .O(gate265inter5));
  nor2  gate2303(.a(gate265inter5), .b(gate265inter2), .O(gate265inter6));
  inv1  gate2304(.a(G642), .O(gate265inter7));
  inv1  gate2305(.a(G770), .O(gate265inter8));
  nand2 gate2306(.a(gate265inter8), .b(gate265inter7), .O(gate265inter9));
  nand2 gate2307(.a(s_251), .b(gate265inter3), .O(gate265inter10));
  nor2  gate2308(.a(gate265inter10), .b(gate265inter9), .O(gate265inter11));
  nor2  gate2309(.a(gate265inter11), .b(gate265inter6), .O(gate265inter12));
  nand2 gate2310(.a(gate265inter12), .b(gate265inter1), .O(G794));
nand2 gate266( .a(G645), .b(G773), .O(G797) );
nand2 gate267( .a(G648), .b(G776), .O(G800) );

  xor2  gate1163(.a(G779), .b(G651), .O(gate268inter0));
  nand2 gate1164(.a(gate268inter0), .b(s_88), .O(gate268inter1));
  and2  gate1165(.a(G779), .b(G651), .O(gate268inter2));
  inv1  gate1166(.a(s_88), .O(gate268inter3));
  inv1  gate1167(.a(s_89), .O(gate268inter4));
  nand2 gate1168(.a(gate268inter4), .b(gate268inter3), .O(gate268inter5));
  nor2  gate1169(.a(gate268inter5), .b(gate268inter2), .O(gate268inter6));
  inv1  gate1170(.a(G651), .O(gate268inter7));
  inv1  gate1171(.a(G779), .O(gate268inter8));
  nand2 gate1172(.a(gate268inter8), .b(gate268inter7), .O(gate268inter9));
  nand2 gate1173(.a(s_89), .b(gate268inter3), .O(gate268inter10));
  nor2  gate1174(.a(gate268inter10), .b(gate268inter9), .O(gate268inter11));
  nor2  gate1175(.a(gate268inter11), .b(gate268inter6), .O(gate268inter12));
  nand2 gate1176(.a(gate268inter12), .b(gate268inter1), .O(G803));
nand2 gate269( .a(G654), .b(G782), .O(G806) );

  xor2  gate1723(.a(G785), .b(G657), .O(gate270inter0));
  nand2 gate1724(.a(gate270inter0), .b(s_168), .O(gate270inter1));
  and2  gate1725(.a(G785), .b(G657), .O(gate270inter2));
  inv1  gate1726(.a(s_168), .O(gate270inter3));
  inv1  gate1727(.a(s_169), .O(gate270inter4));
  nand2 gate1728(.a(gate270inter4), .b(gate270inter3), .O(gate270inter5));
  nor2  gate1729(.a(gate270inter5), .b(gate270inter2), .O(gate270inter6));
  inv1  gate1730(.a(G657), .O(gate270inter7));
  inv1  gate1731(.a(G785), .O(gate270inter8));
  nand2 gate1732(.a(gate270inter8), .b(gate270inter7), .O(gate270inter9));
  nand2 gate1733(.a(s_169), .b(gate270inter3), .O(gate270inter10));
  nor2  gate1734(.a(gate270inter10), .b(gate270inter9), .O(gate270inter11));
  nor2  gate1735(.a(gate270inter11), .b(gate270inter6), .O(gate270inter12));
  nand2 gate1736(.a(gate270inter12), .b(gate270inter1), .O(G809));

  xor2  gate1373(.a(G788), .b(G660), .O(gate271inter0));
  nand2 gate1374(.a(gate271inter0), .b(s_118), .O(gate271inter1));
  and2  gate1375(.a(G788), .b(G660), .O(gate271inter2));
  inv1  gate1376(.a(s_118), .O(gate271inter3));
  inv1  gate1377(.a(s_119), .O(gate271inter4));
  nand2 gate1378(.a(gate271inter4), .b(gate271inter3), .O(gate271inter5));
  nor2  gate1379(.a(gate271inter5), .b(gate271inter2), .O(gate271inter6));
  inv1  gate1380(.a(G660), .O(gate271inter7));
  inv1  gate1381(.a(G788), .O(gate271inter8));
  nand2 gate1382(.a(gate271inter8), .b(gate271inter7), .O(gate271inter9));
  nand2 gate1383(.a(s_119), .b(gate271inter3), .O(gate271inter10));
  nor2  gate1384(.a(gate271inter10), .b(gate271inter9), .O(gate271inter11));
  nor2  gate1385(.a(gate271inter11), .b(gate271inter6), .O(gate271inter12));
  nand2 gate1386(.a(gate271inter12), .b(gate271inter1), .O(G812));
nand2 gate272( .a(G663), .b(G791), .O(G815) );
nand2 gate273( .a(G642), .b(G794), .O(G818) );
nand2 gate274( .a(G770), .b(G794), .O(G819) );
nand2 gate275( .a(G645), .b(G797), .O(G820) );

  xor2  gate2493(.a(G797), .b(G773), .O(gate276inter0));
  nand2 gate2494(.a(gate276inter0), .b(s_278), .O(gate276inter1));
  and2  gate2495(.a(G797), .b(G773), .O(gate276inter2));
  inv1  gate2496(.a(s_278), .O(gate276inter3));
  inv1  gate2497(.a(s_279), .O(gate276inter4));
  nand2 gate2498(.a(gate276inter4), .b(gate276inter3), .O(gate276inter5));
  nor2  gate2499(.a(gate276inter5), .b(gate276inter2), .O(gate276inter6));
  inv1  gate2500(.a(G773), .O(gate276inter7));
  inv1  gate2501(.a(G797), .O(gate276inter8));
  nand2 gate2502(.a(gate276inter8), .b(gate276inter7), .O(gate276inter9));
  nand2 gate2503(.a(s_279), .b(gate276inter3), .O(gate276inter10));
  nor2  gate2504(.a(gate276inter10), .b(gate276inter9), .O(gate276inter11));
  nor2  gate2505(.a(gate276inter11), .b(gate276inter6), .O(gate276inter12));
  nand2 gate2506(.a(gate276inter12), .b(gate276inter1), .O(G821));

  xor2  gate785(.a(G800), .b(G648), .O(gate277inter0));
  nand2 gate786(.a(gate277inter0), .b(s_34), .O(gate277inter1));
  and2  gate787(.a(G800), .b(G648), .O(gate277inter2));
  inv1  gate788(.a(s_34), .O(gate277inter3));
  inv1  gate789(.a(s_35), .O(gate277inter4));
  nand2 gate790(.a(gate277inter4), .b(gate277inter3), .O(gate277inter5));
  nor2  gate791(.a(gate277inter5), .b(gate277inter2), .O(gate277inter6));
  inv1  gate792(.a(G648), .O(gate277inter7));
  inv1  gate793(.a(G800), .O(gate277inter8));
  nand2 gate794(.a(gate277inter8), .b(gate277inter7), .O(gate277inter9));
  nand2 gate795(.a(s_35), .b(gate277inter3), .O(gate277inter10));
  nor2  gate796(.a(gate277inter10), .b(gate277inter9), .O(gate277inter11));
  nor2  gate797(.a(gate277inter11), .b(gate277inter6), .O(gate277inter12));
  nand2 gate798(.a(gate277inter12), .b(gate277inter1), .O(G822));

  xor2  gate1261(.a(G800), .b(G776), .O(gate278inter0));
  nand2 gate1262(.a(gate278inter0), .b(s_102), .O(gate278inter1));
  and2  gate1263(.a(G800), .b(G776), .O(gate278inter2));
  inv1  gate1264(.a(s_102), .O(gate278inter3));
  inv1  gate1265(.a(s_103), .O(gate278inter4));
  nand2 gate1266(.a(gate278inter4), .b(gate278inter3), .O(gate278inter5));
  nor2  gate1267(.a(gate278inter5), .b(gate278inter2), .O(gate278inter6));
  inv1  gate1268(.a(G776), .O(gate278inter7));
  inv1  gate1269(.a(G800), .O(gate278inter8));
  nand2 gate1270(.a(gate278inter8), .b(gate278inter7), .O(gate278inter9));
  nand2 gate1271(.a(s_103), .b(gate278inter3), .O(gate278inter10));
  nor2  gate1272(.a(gate278inter10), .b(gate278inter9), .O(gate278inter11));
  nor2  gate1273(.a(gate278inter11), .b(gate278inter6), .O(gate278inter12));
  nand2 gate1274(.a(gate278inter12), .b(gate278inter1), .O(G823));
nand2 gate279( .a(G651), .b(G803), .O(G824) );

  xor2  gate1835(.a(G803), .b(G779), .O(gate280inter0));
  nand2 gate1836(.a(gate280inter0), .b(s_184), .O(gate280inter1));
  and2  gate1837(.a(G803), .b(G779), .O(gate280inter2));
  inv1  gate1838(.a(s_184), .O(gate280inter3));
  inv1  gate1839(.a(s_185), .O(gate280inter4));
  nand2 gate1840(.a(gate280inter4), .b(gate280inter3), .O(gate280inter5));
  nor2  gate1841(.a(gate280inter5), .b(gate280inter2), .O(gate280inter6));
  inv1  gate1842(.a(G779), .O(gate280inter7));
  inv1  gate1843(.a(G803), .O(gate280inter8));
  nand2 gate1844(.a(gate280inter8), .b(gate280inter7), .O(gate280inter9));
  nand2 gate1845(.a(s_185), .b(gate280inter3), .O(gate280inter10));
  nor2  gate1846(.a(gate280inter10), .b(gate280inter9), .O(gate280inter11));
  nor2  gate1847(.a(gate280inter11), .b(gate280inter6), .O(gate280inter12));
  nand2 gate1848(.a(gate280inter12), .b(gate280inter1), .O(G825));
nand2 gate281( .a(G654), .b(G806), .O(G826) );

  xor2  gate1317(.a(G806), .b(G782), .O(gate282inter0));
  nand2 gate1318(.a(gate282inter0), .b(s_110), .O(gate282inter1));
  and2  gate1319(.a(G806), .b(G782), .O(gate282inter2));
  inv1  gate1320(.a(s_110), .O(gate282inter3));
  inv1  gate1321(.a(s_111), .O(gate282inter4));
  nand2 gate1322(.a(gate282inter4), .b(gate282inter3), .O(gate282inter5));
  nor2  gate1323(.a(gate282inter5), .b(gate282inter2), .O(gate282inter6));
  inv1  gate1324(.a(G782), .O(gate282inter7));
  inv1  gate1325(.a(G806), .O(gate282inter8));
  nand2 gate1326(.a(gate282inter8), .b(gate282inter7), .O(gate282inter9));
  nand2 gate1327(.a(s_111), .b(gate282inter3), .O(gate282inter10));
  nor2  gate1328(.a(gate282inter10), .b(gate282inter9), .O(gate282inter11));
  nor2  gate1329(.a(gate282inter11), .b(gate282inter6), .O(gate282inter12));
  nand2 gate1330(.a(gate282inter12), .b(gate282inter1), .O(G827));
nand2 gate283( .a(G657), .b(G809), .O(G828) );
nand2 gate284( .a(G785), .b(G809), .O(G829) );

  xor2  gate2619(.a(G812), .b(G660), .O(gate285inter0));
  nand2 gate2620(.a(gate285inter0), .b(s_296), .O(gate285inter1));
  and2  gate2621(.a(G812), .b(G660), .O(gate285inter2));
  inv1  gate2622(.a(s_296), .O(gate285inter3));
  inv1  gate2623(.a(s_297), .O(gate285inter4));
  nand2 gate2624(.a(gate285inter4), .b(gate285inter3), .O(gate285inter5));
  nor2  gate2625(.a(gate285inter5), .b(gate285inter2), .O(gate285inter6));
  inv1  gate2626(.a(G660), .O(gate285inter7));
  inv1  gate2627(.a(G812), .O(gate285inter8));
  nand2 gate2628(.a(gate285inter8), .b(gate285inter7), .O(gate285inter9));
  nand2 gate2629(.a(s_297), .b(gate285inter3), .O(gate285inter10));
  nor2  gate2630(.a(gate285inter10), .b(gate285inter9), .O(gate285inter11));
  nor2  gate2631(.a(gate285inter11), .b(gate285inter6), .O(gate285inter12));
  nand2 gate2632(.a(gate285inter12), .b(gate285inter1), .O(G830));
nand2 gate286( .a(G788), .b(G812), .O(G831) );
nand2 gate287( .a(G663), .b(G815), .O(G832) );

  xor2  gate1527(.a(G815), .b(G791), .O(gate288inter0));
  nand2 gate1528(.a(gate288inter0), .b(s_140), .O(gate288inter1));
  and2  gate1529(.a(G815), .b(G791), .O(gate288inter2));
  inv1  gate1530(.a(s_140), .O(gate288inter3));
  inv1  gate1531(.a(s_141), .O(gate288inter4));
  nand2 gate1532(.a(gate288inter4), .b(gate288inter3), .O(gate288inter5));
  nor2  gate1533(.a(gate288inter5), .b(gate288inter2), .O(gate288inter6));
  inv1  gate1534(.a(G791), .O(gate288inter7));
  inv1  gate1535(.a(G815), .O(gate288inter8));
  nand2 gate1536(.a(gate288inter8), .b(gate288inter7), .O(gate288inter9));
  nand2 gate1537(.a(s_141), .b(gate288inter3), .O(gate288inter10));
  nor2  gate1538(.a(gate288inter10), .b(gate288inter9), .O(gate288inter11));
  nor2  gate1539(.a(gate288inter11), .b(gate288inter6), .O(gate288inter12));
  nand2 gate1540(.a(gate288inter12), .b(gate288inter1), .O(G833));

  xor2  gate2395(.a(G819), .b(G818), .O(gate289inter0));
  nand2 gate2396(.a(gate289inter0), .b(s_264), .O(gate289inter1));
  and2  gate2397(.a(G819), .b(G818), .O(gate289inter2));
  inv1  gate2398(.a(s_264), .O(gate289inter3));
  inv1  gate2399(.a(s_265), .O(gate289inter4));
  nand2 gate2400(.a(gate289inter4), .b(gate289inter3), .O(gate289inter5));
  nor2  gate2401(.a(gate289inter5), .b(gate289inter2), .O(gate289inter6));
  inv1  gate2402(.a(G818), .O(gate289inter7));
  inv1  gate2403(.a(G819), .O(gate289inter8));
  nand2 gate2404(.a(gate289inter8), .b(gate289inter7), .O(gate289inter9));
  nand2 gate2405(.a(s_265), .b(gate289inter3), .O(gate289inter10));
  nor2  gate2406(.a(gate289inter10), .b(gate289inter9), .O(gate289inter11));
  nor2  gate2407(.a(gate289inter11), .b(gate289inter6), .O(gate289inter12));
  nand2 gate2408(.a(gate289inter12), .b(gate289inter1), .O(G834));
nand2 gate290( .a(G820), .b(G821), .O(G847) );
nand2 gate291( .a(G822), .b(G823), .O(G860) );

  xor2  gate2283(.a(G825), .b(G824), .O(gate292inter0));
  nand2 gate2284(.a(gate292inter0), .b(s_248), .O(gate292inter1));
  and2  gate2285(.a(G825), .b(G824), .O(gate292inter2));
  inv1  gate2286(.a(s_248), .O(gate292inter3));
  inv1  gate2287(.a(s_249), .O(gate292inter4));
  nand2 gate2288(.a(gate292inter4), .b(gate292inter3), .O(gate292inter5));
  nor2  gate2289(.a(gate292inter5), .b(gate292inter2), .O(gate292inter6));
  inv1  gate2290(.a(G824), .O(gate292inter7));
  inv1  gate2291(.a(G825), .O(gate292inter8));
  nand2 gate2292(.a(gate292inter8), .b(gate292inter7), .O(gate292inter9));
  nand2 gate2293(.a(s_249), .b(gate292inter3), .O(gate292inter10));
  nor2  gate2294(.a(gate292inter10), .b(gate292inter9), .O(gate292inter11));
  nor2  gate2295(.a(gate292inter11), .b(gate292inter6), .O(gate292inter12));
  nand2 gate2296(.a(gate292inter12), .b(gate292inter1), .O(G873));

  xor2  gate2045(.a(G829), .b(G828), .O(gate293inter0));
  nand2 gate2046(.a(gate293inter0), .b(s_214), .O(gate293inter1));
  and2  gate2047(.a(G829), .b(G828), .O(gate293inter2));
  inv1  gate2048(.a(s_214), .O(gate293inter3));
  inv1  gate2049(.a(s_215), .O(gate293inter4));
  nand2 gate2050(.a(gate293inter4), .b(gate293inter3), .O(gate293inter5));
  nor2  gate2051(.a(gate293inter5), .b(gate293inter2), .O(gate293inter6));
  inv1  gate2052(.a(G828), .O(gate293inter7));
  inv1  gate2053(.a(G829), .O(gate293inter8));
  nand2 gate2054(.a(gate293inter8), .b(gate293inter7), .O(gate293inter9));
  nand2 gate2055(.a(s_215), .b(gate293inter3), .O(gate293inter10));
  nor2  gate2056(.a(gate293inter10), .b(gate293inter9), .O(gate293inter11));
  nor2  gate2057(.a(gate293inter11), .b(gate293inter6), .O(gate293inter12));
  nand2 gate2058(.a(gate293inter12), .b(gate293inter1), .O(G886));
nand2 gate294( .a(G832), .b(G833), .O(G899) );

  xor2  gate561(.a(G831), .b(G830), .O(gate295inter0));
  nand2 gate562(.a(gate295inter0), .b(s_2), .O(gate295inter1));
  and2  gate563(.a(G831), .b(G830), .O(gate295inter2));
  inv1  gate564(.a(s_2), .O(gate295inter3));
  inv1  gate565(.a(s_3), .O(gate295inter4));
  nand2 gate566(.a(gate295inter4), .b(gate295inter3), .O(gate295inter5));
  nor2  gate567(.a(gate295inter5), .b(gate295inter2), .O(gate295inter6));
  inv1  gate568(.a(G830), .O(gate295inter7));
  inv1  gate569(.a(G831), .O(gate295inter8));
  nand2 gate570(.a(gate295inter8), .b(gate295inter7), .O(gate295inter9));
  nand2 gate571(.a(s_3), .b(gate295inter3), .O(gate295inter10));
  nor2  gate572(.a(gate295inter10), .b(gate295inter9), .O(gate295inter11));
  nor2  gate573(.a(gate295inter11), .b(gate295inter6), .O(gate295inter12));
  nand2 gate574(.a(gate295inter12), .b(gate295inter1), .O(G912));

  xor2  gate1891(.a(G827), .b(G826), .O(gate296inter0));
  nand2 gate1892(.a(gate296inter0), .b(s_192), .O(gate296inter1));
  and2  gate1893(.a(G827), .b(G826), .O(gate296inter2));
  inv1  gate1894(.a(s_192), .O(gate296inter3));
  inv1  gate1895(.a(s_193), .O(gate296inter4));
  nand2 gate1896(.a(gate296inter4), .b(gate296inter3), .O(gate296inter5));
  nor2  gate1897(.a(gate296inter5), .b(gate296inter2), .O(gate296inter6));
  inv1  gate1898(.a(G826), .O(gate296inter7));
  inv1  gate1899(.a(G827), .O(gate296inter8));
  nand2 gate1900(.a(gate296inter8), .b(gate296inter7), .O(gate296inter9));
  nand2 gate1901(.a(s_193), .b(gate296inter3), .O(gate296inter10));
  nor2  gate1902(.a(gate296inter10), .b(gate296inter9), .O(gate296inter11));
  nor2  gate1903(.a(gate296inter11), .b(gate296inter6), .O(gate296inter12));
  nand2 gate1904(.a(gate296inter12), .b(gate296inter1), .O(G925));
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );

  xor2  gate2521(.a(G1036), .b(G1), .O(gate387inter0));
  nand2 gate2522(.a(gate387inter0), .b(s_282), .O(gate387inter1));
  and2  gate2523(.a(G1036), .b(G1), .O(gate387inter2));
  inv1  gate2524(.a(s_282), .O(gate387inter3));
  inv1  gate2525(.a(s_283), .O(gate387inter4));
  nand2 gate2526(.a(gate387inter4), .b(gate387inter3), .O(gate387inter5));
  nor2  gate2527(.a(gate387inter5), .b(gate387inter2), .O(gate387inter6));
  inv1  gate2528(.a(G1), .O(gate387inter7));
  inv1  gate2529(.a(G1036), .O(gate387inter8));
  nand2 gate2530(.a(gate387inter8), .b(gate387inter7), .O(gate387inter9));
  nand2 gate2531(.a(s_283), .b(gate387inter3), .O(gate387inter10));
  nor2  gate2532(.a(gate387inter10), .b(gate387inter9), .O(gate387inter11));
  nor2  gate2533(.a(gate387inter11), .b(gate387inter6), .O(gate387inter12));
  nand2 gate2534(.a(gate387inter12), .b(gate387inter1), .O(G1132));

  xor2  gate1625(.a(G1039), .b(G2), .O(gate388inter0));
  nand2 gate1626(.a(gate388inter0), .b(s_154), .O(gate388inter1));
  and2  gate1627(.a(G1039), .b(G2), .O(gate388inter2));
  inv1  gate1628(.a(s_154), .O(gate388inter3));
  inv1  gate1629(.a(s_155), .O(gate388inter4));
  nand2 gate1630(.a(gate388inter4), .b(gate388inter3), .O(gate388inter5));
  nor2  gate1631(.a(gate388inter5), .b(gate388inter2), .O(gate388inter6));
  inv1  gate1632(.a(G2), .O(gate388inter7));
  inv1  gate1633(.a(G1039), .O(gate388inter8));
  nand2 gate1634(.a(gate388inter8), .b(gate388inter7), .O(gate388inter9));
  nand2 gate1635(.a(s_155), .b(gate388inter3), .O(gate388inter10));
  nor2  gate1636(.a(gate388inter10), .b(gate388inter9), .O(gate388inter11));
  nor2  gate1637(.a(gate388inter11), .b(gate388inter6), .O(gate388inter12));
  nand2 gate1638(.a(gate388inter12), .b(gate388inter1), .O(G1135));
nand2 gate389( .a(G3), .b(G1042), .O(G1138) );
nand2 gate390( .a(G4), .b(G1045), .O(G1141) );

  xor2  gate1247(.a(G1048), .b(G5), .O(gate391inter0));
  nand2 gate1248(.a(gate391inter0), .b(s_100), .O(gate391inter1));
  and2  gate1249(.a(G1048), .b(G5), .O(gate391inter2));
  inv1  gate1250(.a(s_100), .O(gate391inter3));
  inv1  gate1251(.a(s_101), .O(gate391inter4));
  nand2 gate1252(.a(gate391inter4), .b(gate391inter3), .O(gate391inter5));
  nor2  gate1253(.a(gate391inter5), .b(gate391inter2), .O(gate391inter6));
  inv1  gate1254(.a(G5), .O(gate391inter7));
  inv1  gate1255(.a(G1048), .O(gate391inter8));
  nand2 gate1256(.a(gate391inter8), .b(gate391inter7), .O(gate391inter9));
  nand2 gate1257(.a(s_101), .b(gate391inter3), .O(gate391inter10));
  nor2  gate1258(.a(gate391inter10), .b(gate391inter9), .O(gate391inter11));
  nor2  gate1259(.a(gate391inter11), .b(gate391inter6), .O(gate391inter12));
  nand2 gate1260(.a(gate391inter12), .b(gate391inter1), .O(G1144));

  xor2  gate1499(.a(G1051), .b(G6), .O(gate392inter0));
  nand2 gate1500(.a(gate392inter0), .b(s_136), .O(gate392inter1));
  and2  gate1501(.a(G1051), .b(G6), .O(gate392inter2));
  inv1  gate1502(.a(s_136), .O(gate392inter3));
  inv1  gate1503(.a(s_137), .O(gate392inter4));
  nand2 gate1504(.a(gate392inter4), .b(gate392inter3), .O(gate392inter5));
  nor2  gate1505(.a(gate392inter5), .b(gate392inter2), .O(gate392inter6));
  inv1  gate1506(.a(G6), .O(gate392inter7));
  inv1  gate1507(.a(G1051), .O(gate392inter8));
  nand2 gate1508(.a(gate392inter8), .b(gate392inter7), .O(gate392inter9));
  nand2 gate1509(.a(s_137), .b(gate392inter3), .O(gate392inter10));
  nor2  gate1510(.a(gate392inter10), .b(gate392inter9), .O(gate392inter11));
  nor2  gate1511(.a(gate392inter11), .b(gate392inter6), .O(gate392inter12));
  nand2 gate1512(.a(gate392inter12), .b(gate392inter1), .O(G1147));

  xor2  gate1443(.a(G1054), .b(G7), .O(gate393inter0));
  nand2 gate1444(.a(gate393inter0), .b(s_128), .O(gate393inter1));
  and2  gate1445(.a(G1054), .b(G7), .O(gate393inter2));
  inv1  gate1446(.a(s_128), .O(gate393inter3));
  inv1  gate1447(.a(s_129), .O(gate393inter4));
  nand2 gate1448(.a(gate393inter4), .b(gate393inter3), .O(gate393inter5));
  nor2  gate1449(.a(gate393inter5), .b(gate393inter2), .O(gate393inter6));
  inv1  gate1450(.a(G7), .O(gate393inter7));
  inv1  gate1451(.a(G1054), .O(gate393inter8));
  nand2 gate1452(.a(gate393inter8), .b(gate393inter7), .O(gate393inter9));
  nand2 gate1453(.a(s_129), .b(gate393inter3), .O(gate393inter10));
  nor2  gate1454(.a(gate393inter10), .b(gate393inter9), .O(gate393inter11));
  nor2  gate1455(.a(gate393inter11), .b(gate393inter6), .O(gate393inter12));
  nand2 gate1456(.a(gate393inter12), .b(gate393inter1), .O(G1150));

  xor2  gate1569(.a(G1057), .b(G8), .O(gate394inter0));
  nand2 gate1570(.a(gate394inter0), .b(s_146), .O(gate394inter1));
  and2  gate1571(.a(G1057), .b(G8), .O(gate394inter2));
  inv1  gate1572(.a(s_146), .O(gate394inter3));
  inv1  gate1573(.a(s_147), .O(gate394inter4));
  nand2 gate1574(.a(gate394inter4), .b(gate394inter3), .O(gate394inter5));
  nor2  gate1575(.a(gate394inter5), .b(gate394inter2), .O(gate394inter6));
  inv1  gate1576(.a(G8), .O(gate394inter7));
  inv1  gate1577(.a(G1057), .O(gate394inter8));
  nand2 gate1578(.a(gate394inter8), .b(gate394inter7), .O(gate394inter9));
  nand2 gate1579(.a(s_147), .b(gate394inter3), .O(gate394inter10));
  nor2  gate1580(.a(gate394inter10), .b(gate394inter9), .O(gate394inter11));
  nor2  gate1581(.a(gate394inter11), .b(gate394inter6), .O(gate394inter12));
  nand2 gate1582(.a(gate394inter12), .b(gate394inter1), .O(G1153));
nand2 gate395( .a(G9), .b(G1060), .O(G1156) );
nand2 gate396( .a(G10), .b(G1063), .O(G1159) );

  xor2  gate2087(.a(G1066), .b(G11), .O(gate397inter0));
  nand2 gate2088(.a(gate397inter0), .b(s_220), .O(gate397inter1));
  and2  gate2089(.a(G1066), .b(G11), .O(gate397inter2));
  inv1  gate2090(.a(s_220), .O(gate397inter3));
  inv1  gate2091(.a(s_221), .O(gate397inter4));
  nand2 gate2092(.a(gate397inter4), .b(gate397inter3), .O(gate397inter5));
  nor2  gate2093(.a(gate397inter5), .b(gate397inter2), .O(gate397inter6));
  inv1  gate2094(.a(G11), .O(gate397inter7));
  inv1  gate2095(.a(G1066), .O(gate397inter8));
  nand2 gate2096(.a(gate397inter8), .b(gate397inter7), .O(gate397inter9));
  nand2 gate2097(.a(s_221), .b(gate397inter3), .O(gate397inter10));
  nor2  gate2098(.a(gate397inter10), .b(gate397inter9), .O(gate397inter11));
  nor2  gate2099(.a(gate397inter11), .b(gate397inter6), .O(gate397inter12));
  nand2 gate2100(.a(gate397inter12), .b(gate397inter1), .O(G1162));
nand2 gate398( .a(G12), .b(G1069), .O(G1165) );
nand2 gate399( .a(G13), .b(G1072), .O(G1168) );

  xor2  gate1667(.a(G1075), .b(G14), .O(gate400inter0));
  nand2 gate1668(.a(gate400inter0), .b(s_160), .O(gate400inter1));
  and2  gate1669(.a(G1075), .b(G14), .O(gate400inter2));
  inv1  gate1670(.a(s_160), .O(gate400inter3));
  inv1  gate1671(.a(s_161), .O(gate400inter4));
  nand2 gate1672(.a(gate400inter4), .b(gate400inter3), .O(gate400inter5));
  nor2  gate1673(.a(gate400inter5), .b(gate400inter2), .O(gate400inter6));
  inv1  gate1674(.a(G14), .O(gate400inter7));
  inv1  gate1675(.a(G1075), .O(gate400inter8));
  nand2 gate1676(.a(gate400inter8), .b(gate400inter7), .O(gate400inter9));
  nand2 gate1677(.a(s_161), .b(gate400inter3), .O(gate400inter10));
  nor2  gate1678(.a(gate400inter10), .b(gate400inter9), .O(gate400inter11));
  nor2  gate1679(.a(gate400inter11), .b(gate400inter6), .O(gate400inter12));
  nand2 gate1680(.a(gate400inter12), .b(gate400inter1), .O(G1171));
nand2 gate401( .a(G15), .b(G1078), .O(G1174) );
nand2 gate402( .a(G16), .b(G1081), .O(G1177) );
nand2 gate403( .a(G17), .b(G1084), .O(G1180) );
nand2 gate404( .a(G18), .b(G1087), .O(G1183) );
nand2 gate405( .a(G19), .b(G1090), .O(G1186) );
nand2 gate406( .a(G20), .b(G1093), .O(G1189) );

  xor2  gate2017(.a(G1096), .b(G21), .O(gate407inter0));
  nand2 gate2018(.a(gate407inter0), .b(s_210), .O(gate407inter1));
  and2  gate2019(.a(G1096), .b(G21), .O(gate407inter2));
  inv1  gate2020(.a(s_210), .O(gate407inter3));
  inv1  gate2021(.a(s_211), .O(gate407inter4));
  nand2 gate2022(.a(gate407inter4), .b(gate407inter3), .O(gate407inter5));
  nor2  gate2023(.a(gate407inter5), .b(gate407inter2), .O(gate407inter6));
  inv1  gate2024(.a(G21), .O(gate407inter7));
  inv1  gate2025(.a(G1096), .O(gate407inter8));
  nand2 gate2026(.a(gate407inter8), .b(gate407inter7), .O(gate407inter9));
  nand2 gate2027(.a(s_211), .b(gate407inter3), .O(gate407inter10));
  nor2  gate2028(.a(gate407inter10), .b(gate407inter9), .O(gate407inter11));
  nor2  gate2029(.a(gate407inter11), .b(gate407inter6), .O(gate407inter12));
  nand2 gate2030(.a(gate407inter12), .b(gate407inter1), .O(G1192));

  xor2  gate2003(.a(G1099), .b(G22), .O(gate408inter0));
  nand2 gate2004(.a(gate408inter0), .b(s_208), .O(gate408inter1));
  and2  gate2005(.a(G1099), .b(G22), .O(gate408inter2));
  inv1  gate2006(.a(s_208), .O(gate408inter3));
  inv1  gate2007(.a(s_209), .O(gate408inter4));
  nand2 gate2008(.a(gate408inter4), .b(gate408inter3), .O(gate408inter5));
  nor2  gate2009(.a(gate408inter5), .b(gate408inter2), .O(gate408inter6));
  inv1  gate2010(.a(G22), .O(gate408inter7));
  inv1  gate2011(.a(G1099), .O(gate408inter8));
  nand2 gate2012(.a(gate408inter8), .b(gate408inter7), .O(gate408inter9));
  nand2 gate2013(.a(s_209), .b(gate408inter3), .O(gate408inter10));
  nor2  gate2014(.a(gate408inter10), .b(gate408inter9), .O(gate408inter11));
  nor2  gate2015(.a(gate408inter11), .b(gate408inter6), .O(gate408inter12));
  nand2 gate2016(.a(gate408inter12), .b(gate408inter1), .O(G1195));
nand2 gate409( .a(G23), .b(G1102), .O(G1198) );

  xor2  gate743(.a(G1105), .b(G24), .O(gate410inter0));
  nand2 gate744(.a(gate410inter0), .b(s_28), .O(gate410inter1));
  and2  gate745(.a(G1105), .b(G24), .O(gate410inter2));
  inv1  gate746(.a(s_28), .O(gate410inter3));
  inv1  gate747(.a(s_29), .O(gate410inter4));
  nand2 gate748(.a(gate410inter4), .b(gate410inter3), .O(gate410inter5));
  nor2  gate749(.a(gate410inter5), .b(gate410inter2), .O(gate410inter6));
  inv1  gate750(.a(G24), .O(gate410inter7));
  inv1  gate751(.a(G1105), .O(gate410inter8));
  nand2 gate752(.a(gate410inter8), .b(gate410inter7), .O(gate410inter9));
  nand2 gate753(.a(s_29), .b(gate410inter3), .O(gate410inter10));
  nor2  gate754(.a(gate410inter10), .b(gate410inter9), .O(gate410inter11));
  nor2  gate755(.a(gate410inter11), .b(gate410inter6), .O(gate410inter12));
  nand2 gate756(.a(gate410inter12), .b(gate410inter1), .O(G1201));
nand2 gate411( .a(G25), .b(G1108), .O(G1204) );
nand2 gate412( .a(G26), .b(G1111), .O(G1207) );

  xor2  gate995(.a(G1114), .b(G27), .O(gate413inter0));
  nand2 gate996(.a(gate413inter0), .b(s_64), .O(gate413inter1));
  and2  gate997(.a(G1114), .b(G27), .O(gate413inter2));
  inv1  gate998(.a(s_64), .O(gate413inter3));
  inv1  gate999(.a(s_65), .O(gate413inter4));
  nand2 gate1000(.a(gate413inter4), .b(gate413inter3), .O(gate413inter5));
  nor2  gate1001(.a(gate413inter5), .b(gate413inter2), .O(gate413inter6));
  inv1  gate1002(.a(G27), .O(gate413inter7));
  inv1  gate1003(.a(G1114), .O(gate413inter8));
  nand2 gate1004(.a(gate413inter8), .b(gate413inter7), .O(gate413inter9));
  nand2 gate1005(.a(s_65), .b(gate413inter3), .O(gate413inter10));
  nor2  gate1006(.a(gate413inter10), .b(gate413inter9), .O(gate413inter11));
  nor2  gate1007(.a(gate413inter11), .b(gate413inter6), .O(gate413inter12));
  nand2 gate1008(.a(gate413inter12), .b(gate413inter1), .O(G1210));

  xor2  gate1107(.a(G1117), .b(G28), .O(gate414inter0));
  nand2 gate1108(.a(gate414inter0), .b(s_80), .O(gate414inter1));
  and2  gate1109(.a(G1117), .b(G28), .O(gate414inter2));
  inv1  gate1110(.a(s_80), .O(gate414inter3));
  inv1  gate1111(.a(s_81), .O(gate414inter4));
  nand2 gate1112(.a(gate414inter4), .b(gate414inter3), .O(gate414inter5));
  nor2  gate1113(.a(gate414inter5), .b(gate414inter2), .O(gate414inter6));
  inv1  gate1114(.a(G28), .O(gate414inter7));
  inv1  gate1115(.a(G1117), .O(gate414inter8));
  nand2 gate1116(.a(gate414inter8), .b(gate414inter7), .O(gate414inter9));
  nand2 gate1117(.a(s_81), .b(gate414inter3), .O(gate414inter10));
  nor2  gate1118(.a(gate414inter10), .b(gate414inter9), .O(gate414inter11));
  nor2  gate1119(.a(gate414inter11), .b(gate414inter6), .O(gate414inter12));
  nand2 gate1120(.a(gate414inter12), .b(gate414inter1), .O(G1213));

  xor2  gate687(.a(G1120), .b(G29), .O(gate415inter0));
  nand2 gate688(.a(gate415inter0), .b(s_20), .O(gate415inter1));
  and2  gate689(.a(G1120), .b(G29), .O(gate415inter2));
  inv1  gate690(.a(s_20), .O(gate415inter3));
  inv1  gate691(.a(s_21), .O(gate415inter4));
  nand2 gate692(.a(gate415inter4), .b(gate415inter3), .O(gate415inter5));
  nor2  gate693(.a(gate415inter5), .b(gate415inter2), .O(gate415inter6));
  inv1  gate694(.a(G29), .O(gate415inter7));
  inv1  gate695(.a(G1120), .O(gate415inter8));
  nand2 gate696(.a(gate415inter8), .b(gate415inter7), .O(gate415inter9));
  nand2 gate697(.a(s_21), .b(gate415inter3), .O(gate415inter10));
  nor2  gate698(.a(gate415inter10), .b(gate415inter9), .O(gate415inter11));
  nor2  gate699(.a(gate415inter11), .b(gate415inter6), .O(gate415inter12));
  nand2 gate700(.a(gate415inter12), .b(gate415inter1), .O(G1216));

  xor2  gate631(.a(G1123), .b(G30), .O(gate416inter0));
  nand2 gate632(.a(gate416inter0), .b(s_12), .O(gate416inter1));
  and2  gate633(.a(G1123), .b(G30), .O(gate416inter2));
  inv1  gate634(.a(s_12), .O(gate416inter3));
  inv1  gate635(.a(s_13), .O(gate416inter4));
  nand2 gate636(.a(gate416inter4), .b(gate416inter3), .O(gate416inter5));
  nor2  gate637(.a(gate416inter5), .b(gate416inter2), .O(gate416inter6));
  inv1  gate638(.a(G30), .O(gate416inter7));
  inv1  gate639(.a(G1123), .O(gate416inter8));
  nand2 gate640(.a(gate416inter8), .b(gate416inter7), .O(gate416inter9));
  nand2 gate641(.a(s_13), .b(gate416inter3), .O(gate416inter10));
  nor2  gate642(.a(gate416inter10), .b(gate416inter9), .O(gate416inter11));
  nor2  gate643(.a(gate416inter11), .b(gate416inter6), .O(gate416inter12));
  nand2 gate644(.a(gate416inter12), .b(gate416inter1), .O(G1219));

  xor2  gate1359(.a(G1126), .b(G31), .O(gate417inter0));
  nand2 gate1360(.a(gate417inter0), .b(s_116), .O(gate417inter1));
  and2  gate1361(.a(G1126), .b(G31), .O(gate417inter2));
  inv1  gate1362(.a(s_116), .O(gate417inter3));
  inv1  gate1363(.a(s_117), .O(gate417inter4));
  nand2 gate1364(.a(gate417inter4), .b(gate417inter3), .O(gate417inter5));
  nor2  gate1365(.a(gate417inter5), .b(gate417inter2), .O(gate417inter6));
  inv1  gate1366(.a(G31), .O(gate417inter7));
  inv1  gate1367(.a(G1126), .O(gate417inter8));
  nand2 gate1368(.a(gate417inter8), .b(gate417inter7), .O(gate417inter9));
  nand2 gate1369(.a(s_117), .b(gate417inter3), .O(gate417inter10));
  nor2  gate1370(.a(gate417inter10), .b(gate417inter9), .O(gate417inter11));
  nor2  gate1371(.a(gate417inter11), .b(gate417inter6), .O(gate417inter12));
  nand2 gate1372(.a(gate417inter12), .b(gate417inter1), .O(G1222));
nand2 gate418( .a(G32), .b(G1129), .O(G1225) );
nand2 gate419( .a(G1), .b(G1132), .O(G1228) );
nand2 gate420( .a(G1036), .b(G1132), .O(G1229) );

  xor2  gate729(.a(G1135), .b(G2), .O(gate421inter0));
  nand2 gate730(.a(gate421inter0), .b(s_26), .O(gate421inter1));
  and2  gate731(.a(G1135), .b(G2), .O(gate421inter2));
  inv1  gate732(.a(s_26), .O(gate421inter3));
  inv1  gate733(.a(s_27), .O(gate421inter4));
  nand2 gate734(.a(gate421inter4), .b(gate421inter3), .O(gate421inter5));
  nor2  gate735(.a(gate421inter5), .b(gate421inter2), .O(gate421inter6));
  inv1  gate736(.a(G2), .O(gate421inter7));
  inv1  gate737(.a(G1135), .O(gate421inter8));
  nand2 gate738(.a(gate421inter8), .b(gate421inter7), .O(gate421inter9));
  nand2 gate739(.a(s_27), .b(gate421inter3), .O(gate421inter10));
  nor2  gate740(.a(gate421inter10), .b(gate421inter9), .O(gate421inter11));
  nor2  gate741(.a(gate421inter11), .b(gate421inter6), .O(gate421inter12));
  nand2 gate742(.a(gate421inter12), .b(gate421inter1), .O(G1230));
nand2 gate422( .a(G1039), .b(G1135), .O(G1231) );
nand2 gate423( .a(G3), .b(G1138), .O(G1232) );
nand2 gate424( .a(G1042), .b(G1138), .O(G1233) );
nand2 gate425( .a(G4), .b(G1141), .O(G1234) );
nand2 gate426( .a(G1045), .b(G1141), .O(G1235) );
nand2 gate427( .a(G5), .b(G1144), .O(G1236) );
nand2 gate428( .a(G1048), .b(G1144), .O(G1237) );
nand2 gate429( .a(G6), .b(G1147), .O(G1238) );

  xor2  gate981(.a(G1147), .b(G1051), .O(gate430inter0));
  nand2 gate982(.a(gate430inter0), .b(s_62), .O(gate430inter1));
  and2  gate983(.a(G1147), .b(G1051), .O(gate430inter2));
  inv1  gate984(.a(s_62), .O(gate430inter3));
  inv1  gate985(.a(s_63), .O(gate430inter4));
  nand2 gate986(.a(gate430inter4), .b(gate430inter3), .O(gate430inter5));
  nor2  gate987(.a(gate430inter5), .b(gate430inter2), .O(gate430inter6));
  inv1  gate988(.a(G1051), .O(gate430inter7));
  inv1  gate989(.a(G1147), .O(gate430inter8));
  nand2 gate990(.a(gate430inter8), .b(gate430inter7), .O(gate430inter9));
  nand2 gate991(.a(s_63), .b(gate430inter3), .O(gate430inter10));
  nor2  gate992(.a(gate430inter10), .b(gate430inter9), .O(gate430inter11));
  nor2  gate993(.a(gate430inter11), .b(gate430inter6), .O(gate430inter12));
  nand2 gate994(.a(gate430inter12), .b(gate430inter1), .O(G1239));
nand2 gate431( .a(G7), .b(G1150), .O(G1240) );
nand2 gate432( .a(G1054), .b(G1150), .O(G1241) );
nand2 gate433( .a(G8), .b(G1153), .O(G1242) );
nand2 gate434( .a(G1057), .b(G1153), .O(G1243) );

  xor2  gate1471(.a(G1156), .b(G9), .O(gate435inter0));
  nand2 gate1472(.a(gate435inter0), .b(s_132), .O(gate435inter1));
  and2  gate1473(.a(G1156), .b(G9), .O(gate435inter2));
  inv1  gate1474(.a(s_132), .O(gate435inter3));
  inv1  gate1475(.a(s_133), .O(gate435inter4));
  nand2 gate1476(.a(gate435inter4), .b(gate435inter3), .O(gate435inter5));
  nor2  gate1477(.a(gate435inter5), .b(gate435inter2), .O(gate435inter6));
  inv1  gate1478(.a(G9), .O(gate435inter7));
  inv1  gate1479(.a(G1156), .O(gate435inter8));
  nand2 gate1480(.a(gate435inter8), .b(gate435inter7), .O(gate435inter9));
  nand2 gate1481(.a(s_133), .b(gate435inter3), .O(gate435inter10));
  nor2  gate1482(.a(gate435inter10), .b(gate435inter9), .O(gate435inter11));
  nor2  gate1483(.a(gate435inter11), .b(gate435inter6), .O(gate435inter12));
  nand2 gate1484(.a(gate435inter12), .b(gate435inter1), .O(G1244));
nand2 gate436( .a(G1060), .b(G1156), .O(G1245) );

  xor2  gate1037(.a(G1159), .b(G10), .O(gate437inter0));
  nand2 gate1038(.a(gate437inter0), .b(s_70), .O(gate437inter1));
  and2  gate1039(.a(G1159), .b(G10), .O(gate437inter2));
  inv1  gate1040(.a(s_70), .O(gate437inter3));
  inv1  gate1041(.a(s_71), .O(gate437inter4));
  nand2 gate1042(.a(gate437inter4), .b(gate437inter3), .O(gate437inter5));
  nor2  gate1043(.a(gate437inter5), .b(gate437inter2), .O(gate437inter6));
  inv1  gate1044(.a(G10), .O(gate437inter7));
  inv1  gate1045(.a(G1159), .O(gate437inter8));
  nand2 gate1046(.a(gate437inter8), .b(gate437inter7), .O(gate437inter9));
  nand2 gate1047(.a(s_71), .b(gate437inter3), .O(gate437inter10));
  nor2  gate1048(.a(gate437inter10), .b(gate437inter9), .O(gate437inter11));
  nor2  gate1049(.a(gate437inter11), .b(gate437inter6), .O(gate437inter12));
  nand2 gate1050(.a(gate437inter12), .b(gate437inter1), .O(G1246));

  xor2  gate673(.a(G1159), .b(G1063), .O(gate438inter0));
  nand2 gate674(.a(gate438inter0), .b(s_18), .O(gate438inter1));
  and2  gate675(.a(G1159), .b(G1063), .O(gate438inter2));
  inv1  gate676(.a(s_18), .O(gate438inter3));
  inv1  gate677(.a(s_19), .O(gate438inter4));
  nand2 gate678(.a(gate438inter4), .b(gate438inter3), .O(gate438inter5));
  nor2  gate679(.a(gate438inter5), .b(gate438inter2), .O(gate438inter6));
  inv1  gate680(.a(G1063), .O(gate438inter7));
  inv1  gate681(.a(G1159), .O(gate438inter8));
  nand2 gate682(.a(gate438inter8), .b(gate438inter7), .O(gate438inter9));
  nand2 gate683(.a(s_19), .b(gate438inter3), .O(gate438inter10));
  nor2  gate684(.a(gate438inter10), .b(gate438inter9), .O(gate438inter11));
  nor2  gate685(.a(gate438inter11), .b(gate438inter6), .O(gate438inter12));
  nand2 gate686(.a(gate438inter12), .b(gate438inter1), .O(G1247));

  xor2  gate2325(.a(G1162), .b(G11), .O(gate439inter0));
  nand2 gate2326(.a(gate439inter0), .b(s_254), .O(gate439inter1));
  and2  gate2327(.a(G1162), .b(G11), .O(gate439inter2));
  inv1  gate2328(.a(s_254), .O(gate439inter3));
  inv1  gate2329(.a(s_255), .O(gate439inter4));
  nand2 gate2330(.a(gate439inter4), .b(gate439inter3), .O(gate439inter5));
  nor2  gate2331(.a(gate439inter5), .b(gate439inter2), .O(gate439inter6));
  inv1  gate2332(.a(G11), .O(gate439inter7));
  inv1  gate2333(.a(G1162), .O(gate439inter8));
  nand2 gate2334(.a(gate439inter8), .b(gate439inter7), .O(gate439inter9));
  nand2 gate2335(.a(s_255), .b(gate439inter3), .O(gate439inter10));
  nor2  gate2336(.a(gate439inter10), .b(gate439inter9), .O(gate439inter11));
  nor2  gate2337(.a(gate439inter11), .b(gate439inter6), .O(gate439inter12));
  nand2 gate2338(.a(gate439inter12), .b(gate439inter1), .O(G1248));
nand2 gate440( .a(G1066), .b(G1162), .O(G1249) );
nand2 gate441( .a(G12), .b(G1165), .O(G1250) );

  xor2  gate1457(.a(G1165), .b(G1069), .O(gate442inter0));
  nand2 gate1458(.a(gate442inter0), .b(s_130), .O(gate442inter1));
  and2  gate1459(.a(G1165), .b(G1069), .O(gate442inter2));
  inv1  gate1460(.a(s_130), .O(gate442inter3));
  inv1  gate1461(.a(s_131), .O(gate442inter4));
  nand2 gate1462(.a(gate442inter4), .b(gate442inter3), .O(gate442inter5));
  nor2  gate1463(.a(gate442inter5), .b(gate442inter2), .O(gate442inter6));
  inv1  gate1464(.a(G1069), .O(gate442inter7));
  inv1  gate1465(.a(G1165), .O(gate442inter8));
  nand2 gate1466(.a(gate442inter8), .b(gate442inter7), .O(gate442inter9));
  nand2 gate1467(.a(s_131), .b(gate442inter3), .O(gate442inter10));
  nor2  gate1468(.a(gate442inter10), .b(gate442inter9), .O(gate442inter11));
  nor2  gate1469(.a(gate442inter11), .b(gate442inter6), .O(gate442inter12));
  nand2 gate1470(.a(gate442inter12), .b(gate442inter1), .O(G1251));

  xor2  gate1975(.a(G1168), .b(G13), .O(gate443inter0));
  nand2 gate1976(.a(gate443inter0), .b(s_204), .O(gate443inter1));
  and2  gate1977(.a(G1168), .b(G13), .O(gate443inter2));
  inv1  gate1978(.a(s_204), .O(gate443inter3));
  inv1  gate1979(.a(s_205), .O(gate443inter4));
  nand2 gate1980(.a(gate443inter4), .b(gate443inter3), .O(gate443inter5));
  nor2  gate1981(.a(gate443inter5), .b(gate443inter2), .O(gate443inter6));
  inv1  gate1982(.a(G13), .O(gate443inter7));
  inv1  gate1983(.a(G1168), .O(gate443inter8));
  nand2 gate1984(.a(gate443inter8), .b(gate443inter7), .O(gate443inter9));
  nand2 gate1985(.a(s_205), .b(gate443inter3), .O(gate443inter10));
  nor2  gate1986(.a(gate443inter10), .b(gate443inter9), .O(gate443inter11));
  nor2  gate1987(.a(gate443inter11), .b(gate443inter6), .O(gate443inter12));
  nand2 gate1988(.a(gate443inter12), .b(gate443inter1), .O(G1252));
nand2 gate444( .a(G1072), .b(G1168), .O(G1253) );
nand2 gate445( .a(G14), .b(G1171), .O(G1254) );

  xor2  gate2073(.a(G1171), .b(G1075), .O(gate446inter0));
  nand2 gate2074(.a(gate446inter0), .b(s_218), .O(gate446inter1));
  and2  gate2075(.a(G1171), .b(G1075), .O(gate446inter2));
  inv1  gate2076(.a(s_218), .O(gate446inter3));
  inv1  gate2077(.a(s_219), .O(gate446inter4));
  nand2 gate2078(.a(gate446inter4), .b(gate446inter3), .O(gate446inter5));
  nor2  gate2079(.a(gate446inter5), .b(gate446inter2), .O(gate446inter6));
  inv1  gate2080(.a(G1075), .O(gate446inter7));
  inv1  gate2081(.a(G1171), .O(gate446inter8));
  nand2 gate2082(.a(gate446inter8), .b(gate446inter7), .O(gate446inter9));
  nand2 gate2083(.a(s_219), .b(gate446inter3), .O(gate446inter10));
  nor2  gate2084(.a(gate446inter10), .b(gate446inter9), .O(gate446inter11));
  nor2  gate2085(.a(gate446inter11), .b(gate446inter6), .O(gate446inter12));
  nand2 gate2086(.a(gate446inter12), .b(gate446inter1), .O(G1255));

  xor2  gate2465(.a(G1174), .b(G15), .O(gate447inter0));
  nand2 gate2466(.a(gate447inter0), .b(s_274), .O(gate447inter1));
  and2  gate2467(.a(G1174), .b(G15), .O(gate447inter2));
  inv1  gate2468(.a(s_274), .O(gate447inter3));
  inv1  gate2469(.a(s_275), .O(gate447inter4));
  nand2 gate2470(.a(gate447inter4), .b(gate447inter3), .O(gate447inter5));
  nor2  gate2471(.a(gate447inter5), .b(gate447inter2), .O(gate447inter6));
  inv1  gate2472(.a(G15), .O(gate447inter7));
  inv1  gate2473(.a(G1174), .O(gate447inter8));
  nand2 gate2474(.a(gate447inter8), .b(gate447inter7), .O(gate447inter9));
  nand2 gate2475(.a(s_275), .b(gate447inter3), .O(gate447inter10));
  nor2  gate2476(.a(gate447inter10), .b(gate447inter9), .O(gate447inter11));
  nor2  gate2477(.a(gate447inter11), .b(gate447inter6), .O(gate447inter12));
  nand2 gate2478(.a(gate447inter12), .b(gate447inter1), .O(G1256));
nand2 gate448( .a(G1078), .b(G1174), .O(G1257) );
nand2 gate449( .a(G16), .b(G1177), .O(G1258) );
nand2 gate450( .a(G1081), .b(G1177), .O(G1259) );
nand2 gate451( .a(G17), .b(G1180), .O(G1260) );
nand2 gate452( .a(G1084), .b(G1180), .O(G1261) );

  xor2  gate715(.a(G1183), .b(G18), .O(gate453inter0));
  nand2 gate716(.a(gate453inter0), .b(s_24), .O(gate453inter1));
  and2  gate717(.a(G1183), .b(G18), .O(gate453inter2));
  inv1  gate718(.a(s_24), .O(gate453inter3));
  inv1  gate719(.a(s_25), .O(gate453inter4));
  nand2 gate720(.a(gate453inter4), .b(gate453inter3), .O(gate453inter5));
  nor2  gate721(.a(gate453inter5), .b(gate453inter2), .O(gate453inter6));
  inv1  gate722(.a(G18), .O(gate453inter7));
  inv1  gate723(.a(G1183), .O(gate453inter8));
  nand2 gate724(.a(gate453inter8), .b(gate453inter7), .O(gate453inter9));
  nand2 gate725(.a(s_25), .b(gate453inter3), .O(gate453inter10));
  nor2  gate726(.a(gate453inter10), .b(gate453inter9), .O(gate453inter11));
  nor2  gate727(.a(gate453inter11), .b(gate453inter6), .O(gate453inter12));
  nand2 gate728(.a(gate453inter12), .b(gate453inter1), .O(G1262));
nand2 gate454( .a(G1087), .b(G1183), .O(G1263) );
nand2 gate455( .a(G19), .b(G1186), .O(G1264) );

  xor2  gate1023(.a(G1186), .b(G1090), .O(gate456inter0));
  nand2 gate1024(.a(gate456inter0), .b(s_68), .O(gate456inter1));
  and2  gate1025(.a(G1186), .b(G1090), .O(gate456inter2));
  inv1  gate1026(.a(s_68), .O(gate456inter3));
  inv1  gate1027(.a(s_69), .O(gate456inter4));
  nand2 gate1028(.a(gate456inter4), .b(gate456inter3), .O(gate456inter5));
  nor2  gate1029(.a(gate456inter5), .b(gate456inter2), .O(gate456inter6));
  inv1  gate1030(.a(G1090), .O(gate456inter7));
  inv1  gate1031(.a(G1186), .O(gate456inter8));
  nand2 gate1032(.a(gate456inter8), .b(gate456inter7), .O(gate456inter9));
  nand2 gate1033(.a(s_69), .b(gate456inter3), .O(gate456inter10));
  nor2  gate1034(.a(gate456inter10), .b(gate456inter9), .O(gate456inter11));
  nor2  gate1035(.a(gate456inter11), .b(gate456inter6), .O(gate456inter12));
  nand2 gate1036(.a(gate456inter12), .b(gate456inter1), .O(G1265));

  xor2  gate967(.a(G1189), .b(G20), .O(gate457inter0));
  nand2 gate968(.a(gate457inter0), .b(s_60), .O(gate457inter1));
  and2  gate969(.a(G1189), .b(G20), .O(gate457inter2));
  inv1  gate970(.a(s_60), .O(gate457inter3));
  inv1  gate971(.a(s_61), .O(gate457inter4));
  nand2 gate972(.a(gate457inter4), .b(gate457inter3), .O(gate457inter5));
  nor2  gate973(.a(gate457inter5), .b(gate457inter2), .O(gate457inter6));
  inv1  gate974(.a(G20), .O(gate457inter7));
  inv1  gate975(.a(G1189), .O(gate457inter8));
  nand2 gate976(.a(gate457inter8), .b(gate457inter7), .O(gate457inter9));
  nand2 gate977(.a(s_61), .b(gate457inter3), .O(gate457inter10));
  nor2  gate978(.a(gate457inter10), .b(gate457inter9), .O(gate457inter11));
  nor2  gate979(.a(gate457inter11), .b(gate457inter6), .O(gate457inter12));
  nand2 gate980(.a(gate457inter12), .b(gate457inter1), .O(G1266));
nand2 gate458( .a(G1093), .b(G1189), .O(G1267) );
nand2 gate459( .a(G21), .b(G1192), .O(G1268) );
nand2 gate460( .a(G1096), .b(G1192), .O(G1269) );

  xor2  gate1961(.a(G1195), .b(G22), .O(gate461inter0));
  nand2 gate1962(.a(gate461inter0), .b(s_202), .O(gate461inter1));
  and2  gate1963(.a(G1195), .b(G22), .O(gate461inter2));
  inv1  gate1964(.a(s_202), .O(gate461inter3));
  inv1  gate1965(.a(s_203), .O(gate461inter4));
  nand2 gate1966(.a(gate461inter4), .b(gate461inter3), .O(gate461inter5));
  nor2  gate1967(.a(gate461inter5), .b(gate461inter2), .O(gate461inter6));
  inv1  gate1968(.a(G22), .O(gate461inter7));
  inv1  gate1969(.a(G1195), .O(gate461inter8));
  nand2 gate1970(.a(gate461inter8), .b(gate461inter7), .O(gate461inter9));
  nand2 gate1971(.a(s_203), .b(gate461inter3), .O(gate461inter10));
  nor2  gate1972(.a(gate461inter10), .b(gate461inter9), .O(gate461inter11));
  nor2  gate1973(.a(gate461inter11), .b(gate461inter6), .O(gate461inter12));
  nand2 gate1974(.a(gate461inter12), .b(gate461inter1), .O(G1270));

  xor2  gate1275(.a(G1195), .b(G1099), .O(gate462inter0));
  nand2 gate1276(.a(gate462inter0), .b(s_104), .O(gate462inter1));
  and2  gate1277(.a(G1195), .b(G1099), .O(gate462inter2));
  inv1  gate1278(.a(s_104), .O(gate462inter3));
  inv1  gate1279(.a(s_105), .O(gate462inter4));
  nand2 gate1280(.a(gate462inter4), .b(gate462inter3), .O(gate462inter5));
  nor2  gate1281(.a(gate462inter5), .b(gate462inter2), .O(gate462inter6));
  inv1  gate1282(.a(G1099), .O(gate462inter7));
  inv1  gate1283(.a(G1195), .O(gate462inter8));
  nand2 gate1284(.a(gate462inter8), .b(gate462inter7), .O(gate462inter9));
  nand2 gate1285(.a(s_105), .b(gate462inter3), .O(gate462inter10));
  nor2  gate1286(.a(gate462inter10), .b(gate462inter9), .O(gate462inter11));
  nor2  gate1287(.a(gate462inter11), .b(gate462inter6), .O(gate462inter12));
  nand2 gate1288(.a(gate462inter12), .b(gate462inter1), .O(G1271));
nand2 gate463( .a(G23), .b(G1198), .O(G1272) );

  xor2  gate1541(.a(G1198), .b(G1102), .O(gate464inter0));
  nand2 gate1542(.a(gate464inter0), .b(s_142), .O(gate464inter1));
  and2  gate1543(.a(G1198), .b(G1102), .O(gate464inter2));
  inv1  gate1544(.a(s_142), .O(gate464inter3));
  inv1  gate1545(.a(s_143), .O(gate464inter4));
  nand2 gate1546(.a(gate464inter4), .b(gate464inter3), .O(gate464inter5));
  nor2  gate1547(.a(gate464inter5), .b(gate464inter2), .O(gate464inter6));
  inv1  gate1548(.a(G1102), .O(gate464inter7));
  inv1  gate1549(.a(G1198), .O(gate464inter8));
  nand2 gate1550(.a(gate464inter8), .b(gate464inter7), .O(gate464inter9));
  nand2 gate1551(.a(s_143), .b(gate464inter3), .O(gate464inter10));
  nor2  gate1552(.a(gate464inter10), .b(gate464inter9), .O(gate464inter11));
  nor2  gate1553(.a(gate464inter11), .b(gate464inter6), .O(gate464inter12));
  nand2 gate1554(.a(gate464inter12), .b(gate464inter1), .O(G1273));
nand2 gate465( .a(G24), .b(G1201), .O(G1274) );

  xor2  gate1177(.a(G1201), .b(G1105), .O(gate466inter0));
  nand2 gate1178(.a(gate466inter0), .b(s_90), .O(gate466inter1));
  and2  gate1179(.a(G1201), .b(G1105), .O(gate466inter2));
  inv1  gate1180(.a(s_90), .O(gate466inter3));
  inv1  gate1181(.a(s_91), .O(gate466inter4));
  nand2 gate1182(.a(gate466inter4), .b(gate466inter3), .O(gate466inter5));
  nor2  gate1183(.a(gate466inter5), .b(gate466inter2), .O(gate466inter6));
  inv1  gate1184(.a(G1105), .O(gate466inter7));
  inv1  gate1185(.a(G1201), .O(gate466inter8));
  nand2 gate1186(.a(gate466inter8), .b(gate466inter7), .O(gate466inter9));
  nand2 gate1187(.a(s_91), .b(gate466inter3), .O(gate466inter10));
  nor2  gate1188(.a(gate466inter10), .b(gate466inter9), .O(gate466inter11));
  nor2  gate1189(.a(gate466inter11), .b(gate466inter6), .O(gate466inter12));
  nand2 gate1190(.a(gate466inter12), .b(gate466inter1), .O(G1275));
nand2 gate467( .a(G25), .b(G1204), .O(G1276) );
nand2 gate468( .a(G1108), .b(G1204), .O(G1277) );
nand2 gate469( .a(G26), .b(G1207), .O(G1278) );
nand2 gate470( .a(G1111), .b(G1207), .O(G1279) );
nand2 gate471( .a(G27), .b(G1210), .O(G1280) );

  xor2  gate1009(.a(G1210), .b(G1114), .O(gate472inter0));
  nand2 gate1010(.a(gate472inter0), .b(s_66), .O(gate472inter1));
  and2  gate1011(.a(G1210), .b(G1114), .O(gate472inter2));
  inv1  gate1012(.a(s_66), .O(gate472inter3));
  inv1  gate1013(.a(s_67), .O(gate472inter4));
  nand2 gate1014(.a(gate472inter4), .b(gate472inter3), .O(gate472inter5));
  nor2  gate1015(.a(gate472inter5), .b(gate472inter2), .O(gate472inter6));
  inv1  gate1016(.a(G1114), .O(gate472inter7));
  inv1  gate1017(.a(G1210), .O(gate472inter8));
  nand2 gate1018(.a(gate472inter8), .b(gate472inter7), .O(gate472inter9));
  nand2 gate1019(.a(s_67), .b(gate472inter3), .O(gate472inter10));
  nor2  gate1020(.a(gate472inter10), .b(gate472inter9), .O(gate472inter11));
  nor2  gate1021(.a(gate472inter11), .b(gate472inter6), .O(gate472inter12));
  nand2 gate1022(.a(gate472inter12), .b(gate472inter1), .O(G1281));
nand2 gate473( .a(G28), .b(G1213), .O(G1282) );

  xor2  gate1135(.a(G1213), .b(G1117), .O(gate474inter0));
  nand2 gate1136(.a(gate474inter0), .b(s_84), .O(gate474inter1));
  and2  gate1137(.a(G1213), .b(G1117), .O(gate474inter2));
  inv1  gate1138(.a(s_84), .O(gate474inter3));
  inv1  gate1139(.a(s_85), .O(gate474inter4));
  nand2 gate1140(.a(gate474inter4), .b(gate474inter3), .O(gate474inter5));
  nor2  gate1141(.a(gate474inter5), .b(gate474inter2), .O(gate474inter6));
  inv1  gate1142(.a(G1117), .O(gate474inter7));
  inv1  gate1143(.a(G1213), .O(gate474inter8));
  nand2 gate1144(.a(gate474inter8), .b(gate474inter7), .O(gate474inter9));
  nand2 gate1145(.a(s_85), .b(gate474inter3), .O(gate474inter10));
  nor2  gate1146(.a(gate474inter10), .b(gate474inter9), .O(gate474inter11));
  nor2  gate1147(.a(gate474inter11), .b(gate474inter6), .O(gate474inter12));
  nand2 gate1148(.a(gate474inter12), .b(gate474inter1), .O(G1283));
nand2 gate475( .a(G29), .b(G1216), .O(G1284) );
nand2 gate476( .a(G1120), .b(G1216), .O(G1285) );
nand2 gate477( .a(G30), .b(G1219), .O(G1286) );

  xor2  gate883(.a(G1219), .b(G1123), .O(gate478inter0));
  nand2 gate884(.a(gate478inter0), .b(s_48), .O(gate478inter1));
  and2  gate885(.a(G1219), .b(G1123), .O(gate478inter2));
  inv1  gate886(.a(s_48), .O(gate478inter3));
  inv1  gate887(.a(s_49), .O(gate478inter4));
  nand2 gate888(.a(gate478inter4), .b(gate478inter3), .O(gate478inter5));
  nor2  gate889(.a(gate478inter5), .b(gate478inter2), .O(gate478inter6));
  inv1  gate890(.a(G1123), .O(gate478inter7));
  inv1  gate891(.a(G1219), .O(gate478inter8));
  nand2 gate892(.a(gate478inter8), .b(gate478inter7), .O(gate478inter9));
  nand2 gate893(.a(s_49), .b(gate478inter3), .O(gate478inter10));
  nor2  gate894(.a(gate478inter10), .b(gate478inter9), .O(gate478inter11));
  nor2  gate895(.a(gate478inter11), .b(gate478inter6), .O(gate478inter12));
  nand2 gate896(.a(gate478inter12), .b(gate478inter1), .O(G1287));
nand2 gate479( .a(G31), .b(G1222), .O(G1288) );

  xor2  gate1807(.a(G1222), .b(G1126), .O(gate480inter0));
  nand2 gate1808(.a(gate480inter0), .b(s_180), .O(gate480inter1));
  and2  gate1809(.a(G1222), .b(G1126), .O(gate480inter2));
  inv1  gate1810(.a(s_180), .O(gate480inter3));
  inv1  gate1811(.a(s_181), .O(gate480inter4));
  nand2 gate1812(.a(gate480inter4), .b(gate480inter3), .O(gate480inter5));
  nor2  gate1813(.a(gate480inter5), .b(gate480inter2), .O(gate480inter6));
  inv1  gate1814(.a(G1126), .O(gate480inter7));
  inv1  gate1815(.a(G1222), .O(gate480inter8));
  nand2 gate1816(.a(gate480inter8), .b(gate480inter7), .O(gate480inter9));
  nand2 gate1817(.a(s_181), .b(gate480inter3), .O(gate480inter10));
  nor2  gate1818(.a(gate480inter10), .b(gate480inter9), .O(gate480inter11));
  nor2  gate1819(.a(gate480inter11), .b(gate480inter6), .O(gate480inter12));
  nand2 gate1820(.a(gate480inter12), .b(gate480inter1), .O(G1289));

  xor2  gate1485(.a(G1225), .b(G32), .O(gate481inter0));
  nand2 gate1486(.a(gate481inter0), .b(s_134), .O(gate481inter1));
  and2  gate1487(.a(G1225), .b(G32), .O(gate481inter2));
  inv1  gate1488(.a(s_134), .O(gate481inter3));
  inv1  gate1489(.a(s_135), .O(gate481inter4));
  nand2 gate1490(.a(gate481inter4), .b(gate481inter3), .O(gate481inter5));
  nor2  gate1491(.a(gate481inter5), .b(gate481inter2), .O(gate481inter6));
  inv1  gate1492(.a(G32), .O(gate481inter7));
  inv1  gate1493(.a(G1225), .O(gate481inter8));
  nand2 gate1494(.a(gate481inter8), .b(gate481inter7), .O(gate481inter9));
  nand2 gate1495(.a(s_135), .b(gate481inter3), .O(gate481inter10));
  nor2  gate1496(.a(gate481inter10), .b(gate481inter9), .O(gate481inter11));
  nor2  gate1497(.a(gate481inter11), .b(gate481inter6), .O(gate481inter12));
  nand2 gate1498(.a(gate481inter12), .b(gate481inter1), .O(G1290));
nand2 gate482( .a(G1129), .b(G1225), .O(G1291) );

  xor2  gate1205(.a(G1229), .b(G1228), .O(gate483inter0));
  nand2 gate1206(.a(gate483inter0), .b(s_94), .O(gate483inter1));
  and2  gate1207(.a(G1229), .b(G1228), .O(gate483inter2));
  inv1  gate1208(.a(s_94), .O(gate483inter3));
  inv1  gate1209(.a(s_95), .O(gate483inter4));
  nand2 gate1210(.a(gate483inter4), .b(gate483inter3), .O(gate483inter5));
  nor2  gate1211(.a(gate483inter5), .b(gate483inter2), .O(gate483inter6));
  inv1  gate1212(.a(G1228), .O(gate483inter7));
  inv1  gate1213(.a(G1229), .O(gate483inter8));
  nand2 gate1214(.a(gate483inter8), .b(gate483inter7), .O(gate483inter9));
  nand2 gate1215(.a(s_95), .b(gate483inter3), .O(gate483inter10));
  nor2  gate1216(.a(gate483inter10), .b(gate483inter9), .O(gate483inter11));
  nor2  gate1217(.a(gate483inter11), .b(gate483inter6), .O(gate483inter12));
  nand2 gate1218(.a(gate483inter12), .b(gate483inter1), .O(G1292));

  xor2  gate2269(.a(G1231), .b(G1230), .O(gate484inter0));
  nand2 gate2270(.a(gate484inter0), .b(s_246), .O(gate484inter1));
  and2  gate2271(.a(G1231), .b(G1230), .O(gate484inter2));
  inv1  gate2272(.a(s_246), .O(gate484inter3));
  inv1  gate2273(.a(s_247), .O(gate484inter4));
  nand2 gate2274(.a(gate484inter4), .b(gate484inter3), .O(gate484inter5));
  nor2  gate2275(.a(gate484inter5), .b(gate484inter2), .O(gate484inter6));
  inv1  gate2276(.a(G1230), .O(gate484inter7));
  inv1  gate2277(.a(G1231), .O(gate484inter8));
  nand2 gate2278(.a(gate484inter8), .b(gate484inter7), .O(gate484inter9));
  nand2 gate2279(.a(s_247), .b(gate484inter3), .O(gate484inter10));
  nor2  gate2280(.a(gate484inter10), .b(gate484inter9), .O(gate484inter11));
  nor2  gate2281(.a(gate484inter11), .b(gate484inter6), .O(gate484inter12));
  nand2 gate2282(.a(gate484inter12), .b(gate484inter1), .O(G1293));

  xor2  gate1611(.a(G1233), .b(G1232), .O(gate485inter0));
  nand2 gate1612(.a(gate485inter0), .b(s_152), .O(gate485inter1));
  and2  gate1613(.a(G1233), .b(G1232), .O(gate485inter2));
  inv1  gate1614(.a(s_152), .O(gate485inter3));
  inv1  gate1615(.a(s_153), .O(gate485inter4));
  nand2 gate1616(.a(gate485inter4), .b(gate485inter3), .O(gate485inter5));
  nor2  gate1617(.a(gate485inter5), .b(gate485inter2), .O(gate485inter6));
  inv1  gate1618(.a(G1232), .O(gate485inter7));
  inv1  gate1619(.a(G1233), .O(gate485inter8));
  nand2 gate1620(.a(gate485inter8), .b(gate485inter7), .O(gate485inter9));
  nand2 gate1621(.a(s_153), .b(gate485inter3), .O(gate485inter10));
  nor2  gate1622(.a(gate485inter10), .b(gate485inter9), .O(gate485inter11));
  nor2  gate1623(.a(gate485inter11), .b(gate485inter6), .O(gate485inter12));
  nand2 gate1624(.a(gate485inter12), .b(gate485inter1), .O(G1294));
nand2 gate486( .a(G1234), .b(G1235), .O(G1295) );
nand2 gate487( .a(G1236), .b(G1237), .O(G1296) );
nand2 gate488( .a(G1238), .b(G1239), .O(G1297) );
nand2 gate489( .a(G1240), .b(G1241), .O(G1298) );
nand2 gate490( .a(G1242), .b(G1243), .O(G1299) );

  xor2  gate2549(.a(G1245), .b(G1244), .O(gate491inter0));
  nand2 gate2550(.a(gate491inter0), .b(s_286), .O(gate491inter1));
  and2  gate2551(.a(G1245), .b(G1244), .O(gate491inter2));
  inv1  gate2552(.a(s_286), .O(gate491inter3));
  inv1  gate2553(.a(s_287), .O(gate491inter4));
  nand2 gate2554(.a(gate491inter4), .b(gate491inter3), .O(gate491inter5));
  nor2  gate2555(.a(gate491inter5), .b(gate491inter2), .O(gate491inter6));
  inv1  gate2556(.a(G1244), .O(gate491inter7));
  inv1  gate2557(.a(G1245), .O(gate491inter8));
  nand2 gate2558(.a(gate491inter8), .b(gate491inter7), .O(gate491inter9));
  nand2 gate2559(.a(s_287), .b(gate491inter3), .O(gate491inter10));
  nor2  gate2560(.a(gate491inter10), .b(gate491inter9), .O(gate491inter11));
  nor2  gate2561(.a(gate491inter11), .b(gate491inter6), .O(gate491inter12));
  nand2 gate2562(.a(gate491inter12), .b(gate491inter1), .O(G1300));
nand2 gate492( .a(G1246), .b(G1247), .O(G1301) );

  xor2  gate2409(.a(G1249), .b(G1248), .O(gate493inter0));
  nand2 gate2410(.a(gate493inter0), .b(s_266), .O(gate493inter1));
  and2  gate2411(.a(G1249), .b(G1248), .O(gate493inter2));
  inv1  gate2412(.a(s_266), .O(gate493inter3));
  inv1  gate2413(.a(s_267), .O(gate493inter4));
  nand2 gate2414(.a(gate493inter4), .b(gate493inter3), .O(gate493inter5));
  nor2  gate2415(.a(gate493inter5), .b(gate493inter2), .O(gate493inter6));
  inv1  gate2416(.a(G1248), .O(gate493inter7));
  inv1  gate2417(.a(G1249), .O(gate493inter8));
  nand2 gate2418(.a(gate493inter8), .b(gate493inter7), .O(gate493inter9));
  nand2 gate2419(.a(s_267), .b(gate493inter3), .O(gate493inter10));
  nor2  gate2420(.a(gate493inter10), .b(gate493inter9), .O(gate493inter11));
  nor2  gate2421(.a(gate493inter11), .b(gate493inter6), .O(gate493inter12));
  nand2 gate2422(.a(gate493inter12), .b(gate493inter1), .O(G1302));
nand2 gate494( .a(G1250), .b(G1251), .O(G1303) );

  xor2  gate2563(.a(G1253), .b(G1252), .O(gate495inter0));
  nand2 gate2564(.a(gate495inter0), .b(s_288), .O(gate495inter1));
  and2  gate2565(.a(G1253), .b(G1252), .O(gate495inter2));
  inv1  gate2566(.a(s_288), .O(gate495inter3));
  inv1  gate2567(.a(s_289), .O(gate495inter4));
  nand2 gate2568(.a(gate495inter4), .b(gate495inter3), .O(gate495inter5));
  nor2  gate2569(.a(gate495inter5), .b(gate495inter2), .O(gate495inter6));
  inv1  gate2570(.a(G1252), .O(gate495inter7));
  inv1  gate2571(.a(G1253), .O(gate495inter8));
  nand2 gate2572(.a(gate495inter8), .b(gate495inter7), .O(gate495inter9));
  nand2 gate2573(.a(s_289), .b(gate495inter3), .O(gate495inter10));
  nor2  gate2574(.a(gate495inter10), .b(gate495inter9), .O(gate495inter11));
  nor2  gate2575(.a(gate495inter11), .b(gate495inter6), .O(gate495inter12));
  nand2 gate2576(.a(gate495inter12), .b(gate495inter1), .O(G1304));

  xor2  gate771(.a(G1255), .b(G1254), .O(gate496inter0));
  nand2 gate772(.a(gate496inter0), .b(s_32), .O(gate496inter1));
  and2  gate773(.a(G1255), .b(G1254), .O(gate496inter2));
  inv1  gate774(.a(s_32), .O(gate496inter3));
  inv1  gate775(.a(s_33), .O(gate496inter4));
  nand2 gate776(.a(gate496inter4), .b(gate496inter3), .O(gate496inter5));
  nor2  gate777(.a(gate496inter5), .b(gate496inter2), .O(gate496inter6));
  inv1  gate778(.a(G1254), .O(gate496inter7));
  inv1  gate779(.a(G1255), .O(gate496inter8));
  nand2 gate780(.a(gate496inter8), .b(gate496inter7), .O(gate496inter9));
  nand2 gate781(.a(s_33), .b(gate496inter3), .O(gate496inter10));
  nor2  gate782(.a(gate496inter10), .b(gate496inter9), .O(gate496inter11));
  nor2  gate783(.a(gate496inter11), .b(gate496inter6), .O(gate496inter12));
  nand2 gate784(.a(gate496inter12), .b(gate496inter1), .O(G1305));
nand2 gate497( .a(G1256), .b(G1257), .O(G1306) );
nand2 gate498( .a(G1258), .b(G1259), .O(G1307) );
nand2 gate499( .a(G1260), .b(G1261), .O(G1308) );
nand2 gate500( .a(G1262), .b(G1263), .O(G1309) );
nand2 gate501( .a(G1264), .b(G1265), .O(G1310) );
nand2 gate502( .a(G1266), .b(G1267), .O(G1311) );

  xor2  gate1345(.a(G1269), .b(G1268), .O(gate503inter0));
  nand2 gate1346(.a(gate503inter0), .b(s_114), .O(gate503inter1));
  and2  gate1347(.a(G1269), .b(G1268), .O(gate503inter2));
  inv1  gate1348(.a(s_114), .O(gate503inter3));
  inv1  gate1349(.a(s_115), .O(gate503inter4));
  nand2 gate1350(.a(gate503inter4), .b(gate503inter3), .O(gate503inter5));
  nor2  gate1351(.a(gate503inter5), .b(gate503inter2), .O(gate503inter6));
  inv1  gate1352(.a(G1268), .O(gate503inter7));
  inv1  gate1353(.a(G1269), .O(gate503inter8));
  nand2 gate1354(.a(gate503inter8), .b(gate503inter7), .O(gate503inter9));
  nand2 gate1355(.a(s_115), .b(gate503inter3), .O(gate503inter10));
  nor2  gate1356(.a(gate503inter10), .b(gate503inter9), .O(gate503inter11));
  nor2  gate1357(.a(gate503inter11), .b(gate503inter6), .O(gate503inter12));
  nand2 gate1358(.a(gate503inter12), .b(gate503inter1), .O(G1312));
nand2 gate504( .a(G1270), .b(G1271), .O(G1313) );
nand2 gate505( .a(G1272), .b(G1273), .O(G1314) );

  xor2  gate2339(.a(G1275), .b(G1274), .O(gate506inter0));
  nand2 gate2340(.a(gate506inter0), .b(s_256), .O(gate506inter1));
  and2  gate2341(.a(G1275), .b(G1274), .O(gate506inter2));
  inv1  gate2342(.a(s_256), .O(gate506inter3));
  inv1  gate2343(.a(s_257), .O(gate506inter4));
  nand2 gate2344(.a(gate506inter4), .b(gate506inter3), .O(gate506inter5));
  nor2  gate2345(.a(gate506inter5), .b(gate506inter2), .O(gate506inter6));
  inv1  gate2346(.a(G1274), .O(gate506inter7));
  inv1  gate2347(.a(G1275), .O(gate506inter8));
  nand2 gate2348(.a(gate506inter8), .b(gate506inter7), .O(gate506inter9));
  nand2 gate2349(.a(s_257), .b(gate506inter3), .O(gate506inter10));
  nor2  gate2350(.a(gate506inter10), .b(gate506inter9), .O(gate506inter11));
  nor2  gate2351(.a(gate506inter11), .b(gate506inter6), .O(gate506inter12));
  nand2 gate2352(.a(gate506inter12), .b(gate506inter1), .O(G1315));

  xor2  gate2479(.a(G1277), .b(G1276), .O(gate507inter0));
  nand2 gate2480(.a(gate507inter0), .b(s_276), .O(gate507inter1));
  and2  gate2481(.a(G1277), .b(G1276), .O(gate507inter2));
  inv1  gate2482(.a(s_276), .O(gate507inter3));
  inv1  gate2483(.a(s_277), .O(gate507inter4));
  nand2 gate2484(.a(gate507inter4), .b(gate507inter3), .O(gate507inter5));
  nor2  gate2485(.a(gate507inter5), .b(gate507inter2), .O(gate507inter6));
  inv1  gate2486(.a(G1276), .O(gate507inter7));
  inv1  gate2487(.a(G1277), .O(gate507inter8));
  nand2 gate2488(.a(gate507inter8), .b(gate507inter7), .O(gate507inter9));
  nand2 gate2489(.a(s_277), .b(gate507inter3), .O(gate507inter10));
  nor2  gate2490(.a(gate507inter10), .b(gate507inter9), .O(gate507inter11));
  nor2  gate2491(.a(gate507inter11), .b(gate507inter6), .O(gate507inter12));
  nand2 gate2492(.a(gate507inter12), .b(gate507inter1), .O(G1316));
nand2 gate508( .a(G1278), .b(G1279), .O(G1317) );
nand2 gate509( .a(G1280), .b(G1281), .O(G1318) );
nand2 gate510( .a(G1282), .b(G1283), .O(G1319) );

  xor2  gate1751(.a(G1285), .b(G1284), .O(gate511inter0));
  nand2 gate1752(.a(gate511inter0), .b(s_172), .O(gate511inter1));
  and2  gate1753(.a(G1285), .b(G1284), .O(gate511inter2));
  inv1  gate1754(.a(s_172), .O(gate511inter3));
  inv1  gate1755(.a(s_173), .O(gate511inter4));
  nand2 gate1756(.a(gate511inter4), .b(gate511inter3), .O(gate511inter5));
  nor2  gate1757(.a(gate511inter5), .b(gate511inter2), .O(gate511inter6));
  inv1  gate1758(.a(G1284), .O(gate511inter7));
  inv1  gate1759(.a(G1285), .O(gate511inter8));
  nand2 gate1760(.a(gate511inter8), .b(gate511inter7), .O(gate511inter9));
  nand2 gate1761(.a(s_173), .b(gate511inter3), .O(gate511inter10));
  nor2  gate1762(.a(gate511inter10), .b(gate511inter9), .O(gate511inter11));
  nor2  gate1763(.a(gate511inter11), .b(gate511inter6), .O(gate511inter12));
  nand2 gate1764(.a(gate511inter12), .b(gate511inter1), .O(G1320));

  xor2  gate2185(.a(G1287), .b(G1286), .O(gate512inter0));
  nand2 gate2186(.a(gate512inter0), .b(s_234), .O(gate512inter1));
  and2  gate2187(.a(G1287), .b(G1286), .O(gate512inter2));
  inv1  gate2188(.a(s_234), .O(gate512inter3));
  inv1  gate2189(.a(s_235), .O(gate512inter4));
  nand2 gate2190(.a(gate512inter4), .b(gate512inter3), .O(gate512inter5));
  nor2  gate2191(.a(gate512inter5), .b(gate512inter2), .O(gate512inter6));
  inv1  gate2192(.a(G1286), .O(gate512inter7));
  inv1  gate2193(.a(G1287), .O(gate512inter8));
  nand2 gate2194(.a(gate512inter8), .b(gate512inter7), .O(gate512inter9));
  nand2 gate2195(.a(s_235), .b(gate512inter3), .O(gate512inter10));
  nor2  gate2196(.a(gate512inter10), .b(gate512inter9), .O(gate512inter11));
  nor2  gate2197(.a(gate512inter11), .b(gate512inter6), .O(gate512inter12));
  nand2 gate2198(.a(gate512inter12), .b(gate512inter1), .O(G1321));
nand2 gate513( .a(G1288), .b(G1289), .O(G1322) );
nand2 gate514( .a(G1290), .b(G1291), .O(G1323) );
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule