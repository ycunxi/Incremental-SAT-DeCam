module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);

input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;//RE__PI;

input s_0,s_1;//RE__ALLOW(00,01,10,11);
input s_2,s_3;//RE__ALLOW(00,01,10,11);
input s_4,s_5;//RE__ALLOW(00,01,10,11);
input s_6,s_7;//RE__ALLOW(00,01,10,11);
input s_8,s_9;//RE__ALLOW(00,01,10,11);
input s_10,s_11;//RE__ALLOW(00,01,10,11);
input s_12,s_13;//RE__ALLOW(00,01,10,11);
input s_14,s_15;//RE__ALLOW(00,01,10,11);
input s_16,s_17;//RE__ALLOW(00,01,10,11);
input s_18,s_19;//RE__ALLOW(00,01,10,11);
input s_20,s_21;//RE__ALLOW(00,01,10,11);
input s_22,s_23;//RE__ALLOW(00,01,10,11);
input s_24,s_25;//RE__ALLOW(00,01,10,11);
input s_26,s_27;//RE__ALLOW(00,01,10,11);
input s_28,s_29;//RE__ALLOW(00,01,10,11);
input s_30,s_31;//RE__ALLOW(00,01,10,11);
input s_32,s_33;//RE__ALLOW(00,01,10,11);
input s_34,s_35;//RE__ALLOW(00,01,10,11);
input s_36,s_37;//RE__ALLOW(00,01,10,11);
input s_38,s_39;//RE__ALLOW(00,01,10,11);
input s_40,s_41;//RE__ALLOW(00,01,10,11);
input s_42,s_43;//RE__ALLOW(00,01,10,11);
input s_44,s_45;//RE__ALLOW(00,01,10,11);
input s_46,s_47;//RE__ALLOW(00,01,10,11);
input s_48,s_49;//RE__ALLOW(00,01,10,11);
input s_50,s_51;//RE__ALLOW(00,01,10,11);
input s_52,s_53;//RE__ALLOW(00,01,10,11);
input s_54,s_55;//RE__ALLOW(00,01,10,11);
input s_56,s_57;//RE__ALLOW(00,01,10,11);
input s_58,s_59;//RE__ALLOW(00,01,10,11);
input s_60,s_61;//RE__ALLOW(00,01,10,11);
input s_62,s_63;//RE__ALLOW(00,01,10,11);
input s_64,s_65;//RE__ALLOW(00,01,10,11);
input s_66,s_67;//RE__ALLOW(00,01,10,11);
input s_68,s_69;//RE__ALLOW(00,01,10,11);
input s_70,s_71;//RE__ALLOW(00,01,10,11);
input s_72,s_73;//RE__ALLOW(00,01,10,11);
input s_74,s_75;//RE__ALLOW(00,01,10,11);
input s_76,s_77;//RE__ALLOW(00,01,10,11);
input s_78,s_79;//RE__ALLOW(00,01,10,11);
input s_80,s_81;//RE__ALLOW(00,01,10,11);
input s_82,s_83;//RE__ALLOW(00,01,10,11);
input s_84,s_85;//RE__ALLOW(00,01,10,11);
input s_86,s_87;//RE__ALLOW(00,01,10,11);
input s_88,s_89;//RE__ALLOW(00,01,10,11);
input s_90,s_91;//RE__ALLOW(00,01,10,11);
input s_92,s_93;//RE__ALLOW(00,01,10,11);
input s_94,s_95;//RE__ALLOW(00,01,10,11);
input s_96,s_97;//RE__ALLOW(00,01,10,11);
input s_98,s_99;//RE__ALLOW(00,01,10,11);
input s_100,s_101;//RE__ALLOW(00,01,10,11);
input s_102,s_103;//RE__ALLOW(00,01,10,11);
input s_104,s_105;//RE__ALLOW(00,01,10,11);
input s_106,s_107;//RE__ALLOW(00,01,10,11);
input s_108,s_109;//RE__ALLOW(00,01,10,11);
input s_110,s_111;//RE__ALLOW(00,01,10,11);
input s_112,s_113;//RE__ALLOW(00,01,10,11);
input s_114,s_115;//RE__ALLOW(00,01,10,11);
input s_116,s_117;//RE__ALLOW(00,01,10,11);
input s_118,s_119;//RE__ALLOW(00,01,10,11);
input s_120,s_121;//RE__ALLOW(00,01,10,11);
input s_122,s_123;//RE__ALLOW(00,01,10,11);
input s_124,s_125;//RE__ALLOW(00,01,10,11);
input s_126,s_127;//RE__ALLOW(00,01,10,11);
input s_128,s_129;//RE__ALLOW(00,01,10,11);
input s_130,s_131;//RE__ALLOW(00,01,10,11);
input s_132,s_133;//RE__ALLOW(00,01,10,11);
input s_134,s_135;//RE__ALLOW(00,01,10,11);
input s_136,s_137;//RE__ALLOW(00,01,10,11);
input s_138,s_139;//RE__ALLOW(00,01,10,11);
input s_140,s_141;//RE__ALLOW(00,01,10,11);
input s_142,s_143;//RE__ALLOW(00,01,10,11);
input s_144,s_145;//RE__ALLOW(00,01,10,11);
input s_146,s_147;//RE__ALLOW(00,01,10,11);
input s_148,s_149;//RE__ALLOW(00,01,10,11);
input s_150,s_151;//RE__ALLOW(00,01,10,11);
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;

  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate16inter0, gate16inter1, gate16inter2, gate16inter3, gate16inter4, gate16inter5, gate16inter6, gate16inter7, gate16inter8, gate16inter9, gate16inter10, gate16inter11, gate16inter12, gate402inter0, gate402inter1, gate402inter2, gate402inter3, gate402inter4, gate402inter5, gate402inter6, gate402inter7, gate402inter8, gate402inter9, gate402inter10, gate402inter11, gate402inter12, gate137inter0, gate137inter1, gate137inter2, gate137inter3, gate137inter4, gate137inter5, gate137inter6, gate137inter7, gate137inter8, gate137inter9, gate137inter10, gate137inter11, gate137inter12, gate461inter0, gate461inter1, gate461inter2, gate461inter3, gate461inter4, gate461inter5, gate461inter6, gate461inter7, gate461inter8, gate461inter9, gate461inter10, gate461inter11, gate461inter12, gate431inter0, gate431inter1, gate431inter2, gate431inter3, gate431inter4, gate431inter5, gate431inter6, gate431inter7, gate431inter8, gate431inter9, gate431inter10, gate431inter11, gate431inter12, gate191inter0, gate191inter1, gate191inter2, gate191inter3, gate191inter4, gate191inter5, gate191inter6, gate191inter7, gate191inter8, gate191inter9, gate191inter10, gate191inter11, gate191inter12, gate64inter0, gate64inter1, gate64inter2, gate64inter3, gate64inter4, gate64inter5, gate64inter6, gate64inter7, gate64inter8, gate64inter9, gate64inter10, gate64inter11, gate64inter12, gate196inter0, gate196inter1, gate196inter2, gate196inter3, gate196inter4, gate196inter5, gate196inter6, gate196inter7, gate196inter8, gate196inter9, gate196inter10, gate196inter11, gate196inter12, gate127inter0, gate127inter1, gate127inter2, gate127inter3, gate127inter4, gate127inter5, gate127inter6, gate127inter7, gate127inter8, gate127inter9, gate127inter10, gate127inter11, gate127inter12, gate12inter0, gate12inter1, gate12inter2, gate12inter3, gate12inter4, gate12inter5, gate12inter6, gate12inter7, gate12inter8, gate12inter9, gate12inter10, gate12inter11, gate12inter12, gate233inter0, gate233inter1, gate233inter2, gate233inter3, gate233inter4, gate233inter5, gate233inter6, gate233inter7, gate233inter8, gate233inter9, gate233inter10, gate233inter11, gate233inter12, gate144inter0, gate144inter1, gate144inter2, gate144inter3, gate144inter4, gate144inter5, gate144inter6, gate144inter7, gate144inter8, gate144inter9, gate144inter10, gate144inter11, gate144inter12, gate15inter0, gate15inter1, gate15inter2, gate15inter3, gate15inter4, gate15inter5, gate15inter6, gate15inter7, gate15inter8, gate15inter9, gate15inter10, gate15inter11, gate15inter12, gate169inter0, gate169inter1, gate169inter2, gate169inter3, gate169inter4, gate169inter5, gate169inter6, gate169inter7, gate169inter8, gate169inter9, gate169inter10, gate169inter11, gate169inter12, gate173inter0, gate173inter1, gate173inter2, gate173inter3, gate173inter4, gate173inter5, gate173inter6, gate173inter7, gate173inter8, gate173inter9, gate173inter10, gate173inter11, gate173inter12, gate99inter0, gate99inter1, gate99inter2, gate99inter3, gate99inter4, gate99inter5, gate99inter6, gate99inter7, gate99inter8, gate99inter9, gate99inter10, gate99inter11, gate99inter12, gate118inter0, gate118inter1, gate118inter2, gate118inter3, gate118inter4, gate118inter5, gate118inter6, gate118inter7, gate118inter8, gate118inter9, gate118inter10, gate118inter11, gate118inter12, gate211inter0, gate211inter1, gate211inter2, gate211inter3, gate211inter4, gate211inter5, gate211inter6, gate211inter7, gate211inter8, gate211inter9, gate211inter10, gate211inter11, gate211inter12, gate77inter0, gate77inter1, gate77inter2, gate77inter3, gate77inter4, gate77inter5, gate77inter6, gate77inter7, gate77inter8, gate77inter9, gate77inter10, gate77inter11, gate77inter12, gate391inter0, gate391inter1, gate391inter2, gate391inter3, gate391inter4, gate391inter5, gate391inter6, gate391inter7, gate391inter8, gate391inter9, gate391inter10, gate391inter11, gate391inter12, gate221inter0, gate221inter1, gate221inter2, gate221inter3, gate221inter4, gate221inter5, gate221inter6, gate221inter7, gate221inter8, gate221inter9, gate221inter10, gate221inter11, gate221inter12, gate132inter0, gate132inter1, gate132inter2, gate132inter3, gate132inter4, gate132inter5, gate132inter6, gate132inter7, gate132inter8, gate132inter9, gate132inter10, gate132inter11, gate132inter12, gate117inter0, gate117inter1, gate117inter2, gate117inter3, gate117inter4, gate117inter5, gate117inter6, gate117inter7, gate117inter8, gate117inter9, gate117inter10, gate117inter11, gate117inter12, gate243inter0, gate243inter1, gate243inter2, gate243inter3, gate243inter4, gate243inter5, gate243inter6, gate243inter7, gate243inter8, gate243inter9, gate243inter10, gate243inter11, gate243inter12, gate441inter0, gate441inter1, gate441inter2, gate441inter3, gate441inter4, gate441inter5, gate441inter6, gate441inter7, gate441inter8, gate441inter9, gate441inter10, gate441inter11, gate441inter12, gate208inter0, gate208inter1, gate208inter2, gate208inter3, gate208inter4, gate208inter5, gate208inter6, gate208inter7, gate208inter8, gate208inter9, gate208inter10, gate208inter11, gate208inter12, gate86inter0, gate86inter1, gate86inter2, gate86inter3, gate86inter4, gate86inter5, gate86inter6, gate86inter7, gate86inter8, gate86inter9, gate86inter10, gate86inter11, gate86inter12, gate497inter0, gate497inter1, gate497inter2, gate497inter3, gate497inter4, gate497inter5, gate497inter6, gate497inter7, gate497inter8, gate497inter9, gate497inter10, gate497inter11, gate497inter12, gate444inter0, gate444inter1, gate444inter2, gate444inter3, gate444inter4, gate444inter5, gate444inter6, gate444inter7, gate444inter8, gate444inter9, gate444inter10, gate444inter11, gate444inter12, gate395inter0, gate395inter1, gate395inter2, gate395inter3, gate395inter4, gate395inter5, gate395inter6, gate395inter7, gate395inter8, gate395inter9, gate395inter10, gate395inter11, gate395inter12, gate220inter0, gate220inter1, gate220inter2, gate220inter3, gate220inter4, gate220inter5, gate220inter6, gate220inter7, gate220inter8, gate220inter9, gate220inter10, gate220inter11, gate220inter12, gate410inter0, gate410inter1, gate410inter2, gate410inter3, gate410inter4, gate410inter5, gate410inter6, gate410inter7, gate410inter8, gate410inter9, gate410inter10, gate410inter11, gate410inter12, gate456inter0, gate456inter1, gate456inter2, gate456inter3, gate456inter4, gate456inter5, gate456inter6, gate456inter7, gate456inter8, gate456inter9, gate456inter10, gate456inter11, gate456inter12, gate239inter0, gate239inter1, gate239inter2, gate239inter3, gate239inter4, gate239inter5, gate239inter6, gate239inter7, gate239inter8, gate239inter9, gate239inter10, gate239inter11, gate239inter12, gate153inter0, gate153inter1, gate153inter2, gate153inter3, gate153inter4, gate153inter5, gate153inter6, gate153inter7, gate153inter8, gate153inter9, gate153inter10, gate153inter11, gate153inter12, gate296inter0, gate296inter1, gate296inter2, gate296inter3, gate296inter4, gate296inter5, gate296inter6, gate296inter7, gate296inter8, gate296inter9, gate296inter10, gate296inter11, gate296inter12, gate416inter0, gate416inter1, gate416inter2, gate416inter3, gate416inter4, gate416inter5, gate416inter6, gate416inter7, gate416inter8, gate416inter9, gate416inter10, gate416inter11, gate416inter12, gate156inter0, gate156inter1, gate156inter2, gate156inter3, gate156inter4, gate156inter5, gate156inter6, gate156inter7, gate156inter8, gate156inter9, gate156inter10, gate156inter11, gate156inter12, gate390inter0, gate390inter1, gate390inter2, gate390inter3, gate390inter4, gate390inter5, gate390inter6, gate390inter7, gate390inter8, gate390inter9, gate390inter10, gate390inter11, gate390inter12, gate78inter0, gate78inter1, gate78inter2, gate78inter3, gate78inter4, gate78inter5, gate78inter6, gate78inter7, gate78inter8, gate78inter9, gate78inter10, gate78inter11, gate78inter12, gate56inter0, gate56inter1, gate56inter2, gate56inter3, gate56inter4, gate56inter5, gate56inter6, gate56inter7, gate56inter8, gate56inter9, gate56inter10, gate56inter11, gate56inter12, gate274inter0, gate274inter1, gate274inter2, gate274inter3, gate274inter4, gate274inter5, gate274inter6, gate274inter7, gate274inter8, gate274inter9, gate274inter10, gate274inter11, gate274inter12, gate415inter0, gate415inter1, gate415inter2, gate415inter3, gate415inter4, gate415inter5, gate415inter6, gate415inter7, gate415inter8, gate415inter9, gate415inter10, gate415inter11, gate415inter12, gate473inter0, gate473inter1, gate473inter2, gate473inter3, gate473inter4, gate473inter5, gate473inter6, gate473inter7, gate473inter8, gate473inter9, gate473inter10, gate473inter11, gate473inter12, gate271inter0, gate271inter1, gate271inter2, gate271inter3, gate271inter4, gate271inter5, gate271inter6, gate271inter7, gate271inter8, gate271inter9, gate271inter10, gate271inter11, gate271inter12, gate447inter0, gate447inter1, gate447inter2, gate447inter3, gate447inter4, gate447inter5, gate447inter6, gate447inter7, gate447inter8, gate447inter9, gate447inter10, gate447inter11, gate447inter12, gate493inter0, gate493inter1, gate493inter2, gate493inter3, gate493inter4, gate493inter5, gate493inter6, gate493inter7, gate493inter8, gate493inter9, gate493inter10, gate493inter11, gate493inter12, gate417inter0, gate417inter1, gate417inter2, gate417inter3, gate417inter4, gate417inter5, gate417inter6, gate417inter7, gate417inter8, gate417inter9, gate417inter10, gate417inter11, gate417inter12, gate283inter0, gate283inter1, gate283inter2, gate283inter3, gate283inter4, gate283inter5, gate283inter6, gate283inter7, gate283inter8, gate283inter9, gate283inter10, gate283inter11, gate283inter12, gate237inter0, gate237inter1, gate237inter2, gate237inter3, gate237inter4, gate237inter5, gate237inter6, gate237inter7, gate237inter8, gate237inter9, gate237inter10, gate237inter11, gate237inter12, gate433inter0, gate433inter1, gate433inter2, gate433inter3, gate433inter4, gate433inter5, gate433inter6, gate433inter7, gate433inter8, gate433inter9, gate433inter10, gate433inter11, gate433inter12, gate136inter0, gate136inter1, gate136inter2, gate136inter3, gate136inter4, gate136inter5, gate136inter6, gate136inter7, gate136inter8, gate136inter9, gate136inter10, gate136inter11, gate136inter12, gate234inter0, gate234inter1, gate234inter2, gate234inter3, gate234inter4, gate234inter5, gate234inter6, gate234inter7, gate234inter8, gate234inter9, gate234inter10, gate234inter11, gate234inter12, gate40inter0, gate40inter1, gate40inter2, gate40inter3, gate40inter4, gate40inter5, gate40inter6, gate40inter7, gate40inter8, gate40inter9, gate40inter10, gate40inter11, gate40inter12, gate419inter0, gate419inter1, gate419inter2, gate419inter3, gate419inter4, gate419inter5, gate419inter6, gate419inter7, gate419inter8, gate419inter9, gate419inter10, gate419inter11, gate419inter12, gate66inter0, gate66inter1, gate66inter2, gate66inter3, gate66inter4, gate66inter5, gate66inter6, gate66inter7, gate66inter8, gate66inter9, gate66inter10, gate66inter11, gate66inter12, gate227inter0, gate227inter1, gate227inter2, gate227inter3, gate227inter4, gate227inter5, gate227inter6, gate227inter7, gate227inter8, gate227inter9, gate227inter10, gate227inter11, gate227inter12, gate278inter0, gate278inter1, gate278inter2, gate278inter3, gate278inter4, gate278inter5, gate278inter6, gate278inter7, gate278inter8, gate278inter9, gate278inter10, gate278inter11, gate278inter12, gate108inter0, gate108inter1, gate108inter2, gate108inter3, gate108inter4, gate108inter5, gate108inter6, gate108inter7, gate108inter8, gate108inter9, gate108inter10, gate108inter11, gate108inter12, gate286inter0, gate286inter1, gate286inter2, gate286inter3, gate286inter4, gate286inter5, gate286inter6, gate286inter7, gate286inter8, gate286inter9, gate286inter10, gate286inter11, gate286inter12, gate147inter0, gate147inter1, gate147inter2, gate147inter3, gate147inter4, gate147inter5, gate147inter6, gate147inter7, gate147inter8, gate147inter9, gate147inter10, gate147inter11, gate147inter12, gate93inter0, gate93inter1, gate93inter2, gate93inter3, gate93inter4, gate93inter5, gate93inter6, gate93inter7, gate93inter8, gate93inter9, gate93inter10, gate93inter11, gate93inter12, gate19inter0, gate19inter1, gate19inter2, gate19inter3, gate19inter4, gate19inter5, gate19inter6, gate19inter7, gate19inter8, gate19inter9, gate19inter10, gate19inter11, gate19inter12, gate135inter0, gate135inter1, gate135inter2, gate135inter3, gate135inter4, gate135inter5, gate135inter6, gate135inter7, gate135inter8, gate135inter9, gate135inter10, gate135inter11, gate135inter12, gate158inter0, gate158inter1, gate158inter2, gate158inter3, gate158inter4, gate158inter5, gate158inter6, gate158inter7, gate158inter8, gate158inter9, gate158inter10, gate158inter11, gate158inter12, gate405inter0, gate405inter1, gate405inter2, gate405inter3, gate405inter4, gate405inter5, gate405inter6, gate405inter7, gate405inter8, gate405inter9, gate405inter10, gate405inter11, gate405inter12, gate261inter0, gate261inter1, gate261inter2, gate261inter3, gate261inter4, gate261inter5, gate261inter6, gate261inter7, gate261inter8, gate261inter9, gate261inter10, gate261inter11, gate261inter12, gate489inter0, gate489inter1, gate489inter2, gate489inter3, gate489inter4, gate489inter5, gate489inter6, gate489inter7, gate489inter8, gate489inter9, gate489inter10, gate489inter11, gate489inter12, gate513inter0, gate513inter1, gate513inter2, gate513inter3, gate513inter4, gate513inter5, gate513inter6, gate513inter7, gate513inter8, gate513inter9, gate513inter10, gate513inter11, gate513inter12, gate187inter0, gate187inter1, gate187inter2, gate187inter3, gate187inter4, gate187inter5, gate187inter6, gate187inter7, gate187inter8, gate187inter9, gate187inter10, gate187inter11, gate187inter12, gate418inter0, gate418inter1, gate418inter2, gate418inter3, gate418inter4, gate418inter5, gate418inter6, gate418inter7, gate418inter8, gate418inter9, gate418inter10, gate418inter11, gate418inter12, gate131inter0, gate131inter1, gate131inter2, gate131inter3, gate131inter4, gate131inter5, gate131inter6, gate131inter7, gate131inter8, gate131inter9, gate131inter10, gate131inter11, gate131inter12, gate103inter0, gate103inter1, gate103inter2, gate103inter3, gate103inter4, gate103inter5, gate103inter6, gate103inter7, gate103inter8, gate103inter9, gate103inter10, gate103inter11, gate103inter12, gate425inter0, gate425inter1, gate425inter2, gate425inter3, gate425inter4, gate425inter5, gate425inter6, gate425inter7, gate425inter8, gate425inter9, gate425inter10, gate425inter11, gate425inter12, gate294inter0, gate294inter1, gate294inter2, gate294inter3, gate294inter4, gate294inter5, gate294inter6, gate294inter7, gate294inter8, gate294inter9, gate294inter10, gate294inter11, gate294inter12, gate62inter0, gate62inter1, gate62inter2, gate62inter3, gate62inter4, gate62inter5, gate62inter6, gate62inter7, gate62inter8, gate62inter9, gate62inter10, gate62inter11, gate62inter12;



and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );
nand2 gate9( .a(G1), .b(G2), .O(G266) );
nand2 gate10( .a(G3), .b(G4), .O(G269) );
nand2 gate11( .a(G5), .b(G6), .O(G272) );

  xor2  gate673(.a(G8), .b(G7), .O(gate12inter0));
  nand2 gate674(.a(gate12inter0), .b(s_18), .O(gate12inter1));
  and2  gate675(.a(G8), .b(G7), .O(gate12inter2));
  inv1  gate676(.a(s_18), .O(gate12inter3));
  inv1  gate677(.a(s_19), .O(gate12inter4));
  nand2 gate678(.a(gate12inter4), .b(gate12inter3), .O(gate12inter5));
  nor2  gate679(.a(gate12inter5), .b(gate12inter2), .O(gate12inter6));
  inv1  gate680(.a(G7), .O(gate12inter7));
  inv1  gate681(.a(G8), .O(gate12inter8));
  nand2 gate682(.a(gate12inter8), .b(gate12inter7), .O(gate12inter9));
  nand2 gate683(.a(s_19), .b(gate12inter3), .O(gate12inter10));
  nor2  gate684(.a(gate12inter10), .b(gate12inter9), .O(gate12inter11));
  nor2  gate685(.a(gate12inter11), .b(gate12inter6), .O(gate12inter12));
  nand2 gate686(.a(gate12inter12), .b(gate12inter1), .O(G275));
nand2 gate13( .a(G9), .b(G10), .O(G278) );
nand2 gate14( .a(G11), .b(G12), .O(G281) );

  xor2  gate715(.a(G14), .b(G13), .O(gate15inter0));
  nand2 gate716(.a(gate15inter0), .b(s_24), .O(gate15inter1));
  and2  gate717(.a(G14), .b(G13), .O(gate15inter2));
  inv1  gate718(.a(s_24), .O(gate15inter3));
  inv1  gate719(.a(s_25), .O(gate15inter4));
  nand2 gate720(.a(gate15inter4), .b(gate15inter3), .O(gate15inter5));
  nor2  gate721(.a(gate15inter5), .b(gate15inter2), .O(gate15inter6));
  inv1  gate722(.a(G13), .O(gate15inter7));
  inv1  gate723(.a(G14), .O(gate15inter8));
  nand2 gate724(.a(gate15inter8), .b(gate15inter7), .O(gate15inter9));
  nand2 gate725(.a(s_25), .b(gate15inter3), .O(gate15inter10));
  nor2  gate726(.a(gate15inter10), .b(gate15inter9), .O(gate15inter11));
  nor2  gate727(.a(gate15inter11), .b(gate15inter6), .O(gate15inter12));
  nand2 gate728(.a(gate15inter12), .b(gate15inter1), .O(G284));

  xor2  gate547(.a(G16), .b(G15), .O(gate16inter0));
  nand2 gate548(.a(gate16inter0), .b(s_0), .O(gate16inter1));
  and2  gate549(.a(G16), .b(G15), .O(gate16inter2));
  inv1  gate550(.a(s_0), .O(gate16inter3));
  inv1  gate551(.a(s_1), .O(gate16inter4));
  nand2 gate552(.a(gate16inter4), .b(gate16inter3), .O(gate16inter5));
  nor2  gate553(.a(gate16inter5), .b(gate16inter2), .O(gate16inter6));
  inv1  gate554(.a(G15), .O(gate16inter7));
  inv1  gate555(.a(G16), .O(gate16inter8));
  nand2 gate556(.a(gate16inter8), .b(gate16inter7), .O(gate16inter9));
  nand2 gate557(.a(s_1), .b(gate16inter3), .O(gate16inter10));
  nor2  gate558(.a(gate16inter10), .b(gate16inter9), .O(gate16inter11));
  nor2  gate559(.a(gate16inter11), .b(gate16inter6), .O(gate16inter12));
  nand2 gate560(.a(gate16inter12), .b(gate16inter1), .O(G287));
nand2 gate17( .a(G17), .b(G18), .O(G290) );
nand2 gate18( .a(G19), .b(G20), .O(G293) );

  xor2  gate1415(.a(G22), .b(G21), .O(gate19inter0));
  nand2 gate1416(.a(gate19inter0), .b(s_124), .O(gate19inter1));
  and2  gate1417(.a(G22), .b(G21), .O(gate19inter2));
  inv1  gate1418(.a(s_124), .O(gate19inter3));
  inv1  gate1419(.a(s_125), .O(gate19inter4));
  nand2 gate1420(.a(gate19inter4), .b(gate19inter3), .O(gate19inter5));
  nor2  gate1421(.a(gate19inter5), .b(gate19inter2), .O(gate19inter6));
  inv1  gate1422(.a(G21), .O(gate19inter7));
  inv1  gate1423(.a(G22), .O(gate19inter8));
  nand2 gate1424(.a(gate19inter8), .b(gate19inter7), .O(gate19inter9));
  nand2 gate1425(.a(s_125), .b(gate19inter3), .O(gate19inter10));
  nor2  gate1426(.a(gate19inter10), .b(gate19inter9), .O(gate19inter11));
  nor2  gate1427(.a(gate19inter11), .b(gate19inter6), .O(gate19inter12));
  nand2 gate1428(.a(gate19inter12), .b(gate19inter1), .O(G296));
nand2 gate20( .a(G23), .b(G24), .O(G299) );
nand2 gate21( .a(G25), .b(G26), .O(G302) );
nand2 gate22( .a(G27), .b(G28), .O(G305) );
nand2 gate23( .a(G29), .b(G30), .O(G308) );
nand2 gate24( .a(G31), .b(G32), .O(G311) );
nand2 gate25( .a(G1), .b(G5), .O(G314) );
nand2 gate26( .a(G9), .b(G13), .O(G317) );
nand2 gate27( .a(G2), .b(G6), .O(G320) );
nand2 gate28( .a(G10), .b(G14), .O(G323) );
nand2 gate29( .a(G3), .b(G7), .O(G326) );
nand2 gate30( .a(G11), .b(G15), .O(G329) );
nand2 gate31( .a(G4), .b(G8), .O(G332) );
nand2 gate32( .a(G12), .b(G16), .O(G335) );
nand2 gate33( .a(G17), .b(G21), .O(G338) );
nand2 gate34( .a(G25), .b(G29), .O(G341) );
nand2 gate35( .a(G18), .b(G22), .O(G344) );
nand2 gate36( .a(G26), .b(G30), .O(G347) );
nand2 gate37( .a(G19), .b(G23), .O(G350) );
nand2 gate38( .a(G27), .b(G31), .O(G353) );
nand2 gate39( .a(G20), .b(G24), .O(G356) );

  xor2  gate1289(.a(G32), .b(G28), .O(gate40inter0));
  nand2 gate1290(.a(gate40inter0), .b(s_106), .O(gate40inter1));
  and2  gate1291(.a(G32), .b(G28), .O(gate40inter2));
  inv1  gate1292(.a(s_106), .O(gate40inter3));
  inv1  gate1293(.a(s_107), .O(gate40inter4));
  nand2 gate1294(.a(gate40inter4), .b(gate40inter3), .O(gate40inter5));
  nor2  gate1295(.a(gate40inter5), .b(gate40inter2), .O(gate40inter6));
  inv1  gate1296(.a(G28), .O(gate40inter7));
  inv1  gate1297(.a(G32), .O(gate40inter8));
  nand2 gate1298(.a(gate40inter8), .b(gate40inter7), .O(gate40inter9));
  nand2 gate1299(.a(s_107), .b(gate40inter3), .O(gate40inter10));
  nor2  gate1300(.a(gate40inter10), .b(gate40inter9), .O(gate40inter11));
  nor2  gate1301(.a(gate40inter11), .b(gate40inter6), .O(gate40inter12));
  nand2 gate1302(.a(gate40inter12), .b(gate40inter1), .O(G359));
nand2 gate41( .a(G1), .b(G266), .O(G362) );
nand2 gate42( .a(G2), .b(G266), .O(G363) );
nand2 gate43( .a(G3), .b(G269), .O(G364) );
nand2 gate44( .a(G4), .b(G269), .O(G365) );
nand2 gate45( .a(G5), .b(G272), .O(G366) );
nand2 gate46( .a(G6), .b(G272), .O(G367) );
nand2 gate47( .a(G7), .b(G275), .O(G368) );
nand2 gate48( .a(G8), .b(G275), .O(G369) );
nand2 gate49( .a(G9), .b(G278), .O(G370) );
nand2 gate50( .a(G10), .b(G278), .O(G371) );
nand2 gate51( .a(G11), .b(G281), .O(G372) );
nand2 gate52( .a(G12), .b(G281), .O(G373) );
nand2 gate53( .a(G13), .b(G284), .O(G374) );
nand2 gate54( .a(G14), .b(G284), .O(G375) );
nand2 gate55( .a(G15), .b(G287), .O(G376) );

  xor2  gate1107(.a(G287), .b(G16), .O(gate56inter0));
  nand2 gate1108(.a(gate56inter0), .b(s_80), .O(gate56inter1));
  and2  gate1109(.a(G287), .b(G16), .O(gate56inter2));
  inv1  gate1110(.a(s_80), .O(gate56inter3));
  inv1  gate1111(.a(s_81), .O(gate56inter4));
  nand2 gate1112(.a(gate56inter4), .b(gate56inter3), .O(gate56inter5));
  nor2  gate1113(.a(gate56inter5), .b(gate56inter2), .O(gate56inter6));
  inv1  gate1114(.a(G16), .O(gate56inter7));
  inv1  gate1115(.a(G287), .O(gate56inter8));
  nand2 gate1116(.a(gate56inter8), .b(gate56inter7), .O(gate56inter9));
  nand2 gate1117(.a(s_81), .b(gate56inter3), .O(gate56inter10));
  nor2  gate1118(.a(gate56inter10), .b(gate56inter9), .O(gate56inter11));
  nor2  gate1119(.a(gate56inter11), .b(gate56inter6), .O(gate56inter12));
  nand2 gate1120(.a(gate56inter12), .b(gate56inter1), .O(G377));
nand2 gate57( .a(G17), .b(G290), .O(G378) );
nand2 gate58( .a(G18), .b(G290), .O(G379) );
nand2 gate59( .a(G19), .b(G293), .O(G380) );
nand2 gate60( .a(G20), .b(G293), .O(G381) );
nand2 gate61( .a(G21), .b(G296), .O(G382) );

  xor2  gate1597(.a(G296), .b(G22), .O(gate62inter0));
  nand2 gate1598(.a(gate62inter0), .b(s_150), .O(gate62inter1));
  and2  gate1599(.a(G296), .b(G22), .O(gate62inter2));
  inv1  gate1600(.a(s_150), .O(gate62inter3));
  inv1  gate1601(.a(s_151), .O(gate62inter4));
  nand2 gate1602(.a(gate62inter4), .b(gate62inter3), .O(gate62inter5));
  nor2  gate1603(.a(gate62inter5), .b(gate62inter2), .O(gate62inter6));
  inv1  gate1604(.a(G22), .O(gate62inter7));
  inv1  gate1605(.a(G296), .O(gate62inter8));
  nand2 gate1606(.a(gate62inter8), .b(gate62inter7), .O(gate62inter9));
  nand2 gate1607(.a(s_151), .b(gate62inter3), .O(gate62inter10));
  nor2  gate1608(.a(gate62inter10), .b(gate62inter9), .O(gate62inter11));
  nor2  gate1609(.a(gate62inter11), .b(gate62inter6), .O(gate62inter12));
  nand2 gate1610(.a(gate62inter12), .b(gate62inter1), .O(G383));
nand2 gate63( .a(G23), .b(G299), .O(G384) );

  xor2  gate631(.a(G299), .b(G24), .O(gate64inter0));
  nand2 gate632(.a(gate64inter0), .b(s_12), .O(gate64inter1));
  and2  gate633(.a(G299), .b(G24), .O(gate64inter2));
  inv1  gate634(.a(s_12), .O(gate64inter3));
  inv1  gate635(.a(s_13), .O(gate64inter4));
  nand2 gate636(.a(gate64inter4), .b(gate64inter3), .O(gate64inter5));
  nor2  gate637(.a(gate64inter5), .b(gate64inter2), .O(gate64inter6));
  inv1  gate638(.a(G24), .O(gate64inter7));
  inv1  gate639(.a(G299), .O(gate64inter8));
  nand2 gate640(.a(gate64inter8), .b(gate64inter7), .O(gate64inter9));
  nand2 gate641(.a(s_13), .b(gate64inter3), .O(gate64inter10));
  nor2  gate642(.a(gate64inter10), .b(gate64inter9), .O(gate64inter11));
  nor2  gate643(.a(gate64inter11), .b(gate64inter6), .O(gate64inter12));
  nand2 gate644(.a(gate64inter12), .b(gate64inter1), .O(G385));
nand2 gate65( .a(G25), .b(G302), .O(G386) );

  xor2  gate1317(.a(G302), .b(G26), .O(gate66inter0));
  nand2 gate1318(.a(gate66inter0), .b(s_110), .O(gate66inter1));
  and2  gate1319(.a(G302), .b(G26), .O(gate66inter2));
  inv1  gate1320(.a(s_110), .O(gate66inter3));
  inv1  gate1321(.a(s_111), .O(gate66inter4));
  nand2 gate1322(.a(gate66inter4), .b(gate66inter3), .O(gate66inter5));
  nor2  gate1323(.a(gate66inter5), .b(gate66inter2), .O(gate66inter6));
  inv1  gate1324(.a(G26), .O(gate66inter7));
  inv1  gate1325(.a(G302), .O(gate66inter8));
  nand2 gate1326(.a(gate66inter8), .b(gate66inter7), .O(gate66inter9));
  nand2 gate1327(.a(s_111), .b(gate66inter3), .O(gate66inter10));
  nor2  gate1328(.a(gate66inter10), .b(gate66inter9), .O(gate66inter11));
  nor2  gate1329(.a(gate66inter11), .b(gate66inter6), .O(gate66inter12));
  nand2 gate1330(.a(gate66inter12), .b(gate66inter1), .O(G387));
nand2 gate67( .a(G27), .b(G305), .O(G388) );
nand2 gate68( .a(G28), .b(G305), .O(G389) );
nand2 gate69( .a(G29), .b(G308), .O(G390) );
nand2 gate70( .a(G30), .b(G308), .O(G391) );
nand2 gate71( .a(G31), .b(G311), .O(G392) );
nand2 gate72( .a(G32), .b(G311), .O(G393) );
nand2 gate73( .a(G1), .b(G314), .O(G394) );
nand2 gate74( .a(G5), .b(G314), .O(G395) );
nand2 gate75( .a(G9), .b(G317), .O(G396) );
nand2 gate76( .a(G13), .b(G317), .O(G397) );

  xor2  gate799(.a(G320), .b(G2), .O(gate77inter0));
  nand2 gate800(.a(gate77inter0), .b(s_36), .O(gate77inter1));
  and2  gate801(.a(G320), .b(G2), .O(gate77inter2));
  inv1  gate802(.a(s_36), .O(gate77inter3));
  inv1  gate803(.a(s_37), .O(gate77inter4));
  nand2 gate804(.a(gate77inter4), .b(gate77inter3), .O(gate77inter5));
  nor2  gate805(.a(gate77inter5), .b(gate77inter2), .O(gate77inter6));
  inv1  gate806(.a(G2), .O(gate77inter7));
  inv1  gate807(.a(G320), .O(gate77inter8));
  nand2 gate808(.a(gate77inter8), .b(gate77inter7), .O(gate77inter9));
  nand2 gate809(.a(s_37), .b(gate77inter3), .O(gate77inter10));
  nor2  gate810(.a(gate77inter10), .b(gate77inter9), .O(gate77inter11));
  nor2  gate811(.a(gate77inter11), .b(gate77inter6), .O(gate77inter12));
  nand2 gate812(.a(gate77inter12), .b(gate77inter1), .O(G398));

  xor2  gate1093(.a(G320), .b(G6), .O(gate78inter0));
  nand2 gate1094(.a(gate78inter0), .b(s_78), .O(gate78inter1));
  and2  gate1095(.a(G320), .b(G6), .O(gate78inter2));
  inv1  gate1096(.a(s_78), .O(gate78inter3));
  inv1  gate1097(.a(s_79), .O(gate78inter4));
  nand2 gate1098(.a(gate78inter4), .b(gate78inter3), .O(gate78inter5));
  nor2  gate1099(.a(gate78inter5), .b(gate78inter2), .O(gate78inter6));
  inv1  gate1100(.a(G6), .O(gate78inter7));
  inv1  gate1101(.a(G320), .O(gate78inter8));
  nand2 gate1102(.a(gate78inter8), .b(gate78inter7), .O(gate78inter9));
  nand2 gate1103(.a(s_79), .b(gate78inter3), .O(gate78inter10));
  nor2  gate1104(.a(gate78inter10), .b(gate78inter9), .O(gate78inter11));
  nor2  gate1105(.a(gate78inter11), .b(gate78inter6), .O(gate78inter12));
  nand2 gate1106(.a(gate78inter12), .b(gate78inter1), .O(G399));
nand2 gate79( .a(G10), .b(G323), .O(G400) );
nand2 gate80( .a(G14), .b(G323), .O(G401) );
nand2 gate81( .a(G3), .b(G326), .O(G402) );
nand2 gate82( .a(G7), .b(G326), .O(G403) );
nand2 gate83( .a(G11), .b(G329), .O(G404) );
nand2 gate84( .a(G15), .b(G329), .O(G405) );
nand2 gate85( .a(G4), .b(G332), .O(G406) );

  xor2  gate911(.a(G332), .b(G8), .O(gate86inter0));
  nand2 gate912(.a(gate86inter0), .b(s_52), .O(gate86inter1));
  and2  gate913(.a(G332), .b(G8), .O(gate86inter2));
  inv1  gate914(.a(s_52), .O(gate86inter3));
  inv1  gate915(.a(s_53), .O(gate86inter4));
  nand2 gate916(.a(gate86inter4), .b(gate86inter3), .O(gate86inter5));
  nor2  gate917(.a(gate86inter5), .b(gate86inter2), .O(gate86inter6));
  inv1  gate918(.a(G8), .O(gate86inter7));
  inv1  gate919(.a(G332), .O(gate86inter8));
  nand2 gate920(.a(gate86inter8), .b(gate86inter7), .O(gate86inter9));
  nand2 gate921(.a(s_53), .b(gate86inter3), .O(gate86inter10));
  nor2  gate922(.a(gate86inter10), .b(gate86inter9), .O(gate86inter11));
  nor2  gate923(.a(gate86inter11), .b(gate86inter6), .O(gate86inter12));
  nand2 gate924(.a(gate86inter12), .b(gate86inter1), .O(G407));
nand2 gate87( .a(G12), .b(G335), .O(G408) );
nand2 gate88( .a(G16), .b(G335), .O(G409) );
nand2 gate89( .a(G17), .b(G338), .O(G410) );
nand2 gate90( .a(G21), .b(G338), .O(G411) );
nand2 gate91( .a(G25), .b(G341), .O(G412) );
nand2 gate92( .a(G29), .b(G341), .O(G413) );

  xor2  gate1401(.a(G344), .b(G18), .O(gate93inter0));
  nand2 gate1402(.a(gate93inter0), .b(s_122), .O(gate93inter1));
  and2  gate1403(.a(G344), .b(G18), .O(gate93inter2));
  inv1  gate1404(.a(s_122), .O(gate93inter3));
  inv1  gate1405(.a(s_123), .O(gate93inter4));
  nand2 gate1406(.a(gate93inter4), .b(gate93inter3), .O(gate93inter5));
  nor2  gate1407(.a(gate93inter5), .b(gate93inter2), .O(gate93inter6));
  inv1  gate1408(.a(G18), .O(gate93inter7));
  inv1  gate1409(.a(G344), .O(gate93inter8));
  nand2 gate1410(.a(gate93inter8), .b(gate93inter7), .O(gate93inter9));
  nand2 gate1411(.a(s_123), .b(gate93inter3), .O(gate93inter10));
  nor2  gate1412(.a(gate93inter10), .b(gate93inter9), .O(gate93inter11));
  nor2  gate1413(.a(gate93inter11), .b(gate93inter6), .O(gate93inter12));
  nand2 gate1414(.a(gate93inter12), .b(gate93inter1), .O(G414));
nand2 gate94( .a(G22), .b(G344), .O(G415) );
nand2 gate95( .a(G26), .b(G347), .O(G416) );
nand2 gate96( .a(G30), .b(G347), .O(G417) );
nand2 gate97( .a(G19), .b(G350), .O(G418) );
nand2 gate98( .a(G23), .b(G350), .O(G419) );

  xor2  gate757(.a(G353), .b(G27), .O(gate99inter0));
  nand2 gate758(.a(gate99inter0), .b(s_30), .O(gate99inter1));
  and2  gate759(.a(G353), .b(G27), .O(gate99inter2));
  inv1  gate760(.a(s_30), .O(gate99inter3));
  inv1  gate761(.a(s_31), .O(gate99inter4));
  nand2 gate762(.a(gate99inter4), .b(gate99inter3), .O(gate99inter5));
  nor2  gate763(.a(gate99inter5), .b(gate99inter2), .O(gate99inter6));
  inv1  gate764(.a(G27), .O(gate99inter7));
  inv1  gate765(.a(G353), .O(gate99inter8));
  nand2 gate766(.a(gate99inter8), .b(gate99inter7), .O(gate99inter9));
  nand2 gate767(.a(s_31), .b(gate99inter3), .O(gate99inter10));
  nor2  gate768(.a(gate99inter10), .b(gate99inter9), .O(gate99inter11));
  nor2  gate769(.a(gate99inter11), .b(gate99inter6), .O(gate99inter12));
  nand2 gate770(.a(gate99inter12), .b(gate99inter1), .O(G420));
nand2 gate100( .a(G31), .b(G353), .O(G421) );
nand2 gate101( .a(G20), .b(G356), .O(G422) );
nand2 gate102( .a(G24), .b(G356), .O(G423) );

  xor2  gate1555(.a(G359), .b(G28), .O(gate103inter0));
  nand2 gate1556(.a(gate103inter0), .b(s_144), .O(gate103inter1));
  and2  gate1557(.a(G359), .b(G28), .O(gate103inter2));
  inv1  gate1558(.a(s_144), .O(gate103inter3));
  inv1  gate1559(.a(s_145), .O(gate103inter4));
  nand2 gate1560(.a(gate103inter4), .b(gate103inter3), .O(gate103inter5));
  nor2  gate1561(.a(gate103inter5), .b(gate103inter2), .O(gate103inter6));
  inv1  gate1562(.a(G28), .O(gate103inter7));
  inv1  gate1563(.a(G359), .O(gate103inter8));
  nand2 gate1564(.a(gate103inter8), .b(gate103inter7), .O(gate103inter9));
  nand2 gate1565(.a(s_145), .b(gate103inter3), .O(gate103inter10));
  nor2  gate1566(.a(gate103inter10), .b(gate103inter9), .O(gate103inter11));
  nor2  gate1567(.a(gate103inter11), .b(gate103inter6), .O(gate103inter12));
  nand2 gate1568(.a(gate103inter12), .b(gate103inter1), .O(G424));
nand2 gate104( .a(G32), .b(G359), .O(G425) );
nand2 gate105( .a(G362), .b(G363), .O(G426) );
nand2 gate106( .a(G364), .b(G365), .O(G429) );
nand2 gate107( .a(G366), .b(G367), .O(G432) );

  xor2  gate1359(.a(G369), .b(G368), .O(gate108inter0));
  nand2 gate1360(.a(gate108inter0), .b(s_116), .O(gate108inter1));
  and2  gate1361(.a(G369), .b(G368), .O(gate108inter2));
  inv1  gate1362(.a(s_116), .O(gate108inter3));
  inv1  gate1363(.a(s_117), .O(gate108inter4));
  nand2 gate1364(.a(gate108inter4), .b(gate108inter3), .O(gate108inter5));
  nor2  gate1365(.a(gate108inter5), .b(gate108inter2), .O(gate108inter6));
  inv1  gate1366(.a(G368), .O(gate108inter7));
  inv1  gate1367(.a(G369), .O(gate108inter8));
  nand2 gate1368(.a(gate108inter8), .b(gate108inter7), .O(gate108inter9));
  nand2 gate1369(.a(s_117), .b(gate108inter3), .O(gate108inter10));
  nor2  gate1370(.a(gate108inter10), .b(gate108inter9), .O(gate108inter11));
  nor2  gate1371(.a(gate108inter11), .b(gate108inter6), .O(gate108inter12));
  nand2 gate1372(.a(gate108inter12), .b(gate108inter1), .O(G435));
nand2 gate109( .a(G370), .b(G371), .O(G438) );
nand2 gate110( .a(G372), .b(G373), .O(G441) );
nand2 gate111( .a(G374), .b(G375), .O(G444) );
nand2 gate112( .a(G376), .b(G377), .O(G447) );
nand2 gate113( .a(G378), .b(G379), .O(G450) );
nand2 gate114( .a(G380), .b(G381), .O(G453) );
nand2 gate115( .a(G382), .b(G383), .O(G456) );
nand2 gate116( .a(G384), .b(G385), .O(G459) );

  xor2  gate855(.a(G387), .b(G386), .O(gate117inter0));
  nand2 gate856(.a(gate117inter0), .b(s_44), .O(gate117inter1));
  and2  gate857(.a(G387), .b(G386), .O(gate117inter2));
  inv1  gate858(.a(s_44), .O(gate117inter3));
  inv1  gate859(.a(s_45), .O(gate117inter4));
  nand2 gate860(.a(gate117inter4), .b(gate117inter3), .O(gate117inter5));
  nor2  gate861(.a(gate117inter5), .b(gate117inter2), .O(gate117inter6));
  inv1  gate862(.a(G386), .O(gate117inter7));
  inv1  gate863(.a(G387), .O(gate117inter8));
  nand2 gate864(.a(gate117inter8), .b(gate117inter7), .O(gate117inter9));
  nand2 gate865(.a(s_45), .b(gate117inter3), .O(gate117inter10));
  nor2  gate866(.a(gate117inter10), .b(gate117inter9), .O(gate117inter11));
  nor2  gate867(.a(gate117inter11), .b(gate117inter6), .O(gate117inter12));
  nand2 gate868(.a(gate117inter12), .b(gate117inter1), .O(G462));

  xor2  gate771(.a(G389), .b(G388), .O(gate118inter0));
  nand2 gate772(.a(gate118inter0), .b(s_32), .O(gate118inter1));
  and2  gate773(.a(G389), .b(G388), .O(gate118inter2));
  inv1  gate774(.a(s_32), .O(gate118inter3));
  inv1  gate775(.a(s_33), .O(gate118inter4));
  nand2 gate776(.a(gate118inter4), .b(gate118inter3), .O(gate118inter5));
  nor2  gate777(.a(gate118inter5), .b(gate118inter2), .O(gate118inter6));
  inv1  gate778(.a(G388), .O(gate118inter7));
  inv1  gate779(.a(G389), .O(gate118inter8));
  nand2 gate780(.a(gate118inter8), .b(gate118inter7), .O(gate118inter9));
  nand2 gate781(.a(s_33), .b(gate118inter3), .O(gate118inter10));
  nor2  gate782(.a(gate118inter10), .b(gate118inter9), .O(gate118inter11));
  nor2  gate783(.a(gate118inter11), .b(gate118inter6), .O(gate118inter12));
  nand2 gate784(.a(gate118inter12), .b(gate118inter1), .O(G465));
nand2 gate119( .a(G390), .b(G391), .O(G468) );
nand2 gate120( .a(G392), .b(G393), .O(G471) );
nand2 gate121( .a(G394), .b(G395), .O(G474) );
nand2 gate122( .a(G396), .b(G397), .O(G477) );
nand2 gate123( .a(G398), .b(G399), .O(G480) );
nand2 gate124( .a(G400), .b(G401), .O(G483) );
nand2 gate125( .a(G402), .b(G403), .O(G486) );
nand2 gate126( .a(G404), .b(G405), .O(G489) );

  xor2  gate659(.a(G407), .b(G406), .O(gate127inter0));
  nand2 gate660(.a(gate127inter0), .b(s_16), .O(gate127inter1));
  and2  gate661(.a(G407), .b(G406), .O(gate127inter2));
  inv1  gate662(.a(s_16), .O(gate127inter3));
  inv1  gate663(.a(s_17), .O(gate127inter4));
  nand2 gate664(.a(gate127inter4), .b(gate127inter3), .O(gate127inter5));
  nor2  gate665(.a(gate127inter5), .b(gate127inter2), .O(gate127inter6));
  inv1  gate666(.a(G406), .O(gate127inter7));
  inv1  gate667(.a(G407), .O(gate127inter8));
  nand2 gate668(.a(gate127inter8), .b(gate127inter7), .O(gate127inter9));
  nand2 gate669(.a(s_17), .b(gate127inter3), .O(gate127inter10));
  nor2  gate670(.a(gate127inter10), .b(gate127inter9), .O(gate127inter11));
  nor2  gate671(.a(gate127inter11), .b(gate127inter6), .O(gate127inter12));
  nand2 gate672(.a(gate127inter12), .b(gate127inter1), .O(G492));
nand2 gate128( .a(G408), .b(G409), .O(G495) );
nand2 gate129( .a(G410), .b(G411), .O(G498) );
nand2 gate130( .a(G412), .b(G413), .O(G501) );

  xor2  gate1541(.a(G415), .b(G414), .O(gate131inter0));
  nand2 gate1542(.a(gate131inter0), .b(s_142), .O(gate131inter1));
  and2  gate1543(.a(G415), .b(G414), .O(gate131inter2));
  inv1  gate1544(.a(s_142), .O(gate131inter3));
  inv1  gate1545(.a(s_143), .O(gate131inter4));
  nand2 gate1546(.a(gate131inter4), .b(gate131inter3), .O(gate131inter5));
  nor2  gate1547(.a(gate131inter5), .b(gate131inter2), .O(gate131inter6));
  inv1  gate1548(.a(G414), .O(gate131inter7));
  inv1  gate1549(.a(G415), .O(gate131inter8));
  nand2 gate1550(.a(gate131inter8), .b(gate131inter7), .O(gate131inter9));
  nand2 gate1551(.a(s_143), .b(gate131inter3), .O(gate131inter10));
  nor2  gate1552(.a(gate131inter10), .b(gate131inter9), .O(gate131inter11));
  nor2  gate1553(.a(gate131inter11), .b(gate131inter6), .O(gate131inter12));
  nand2 gate1554(.a(gate131inter12), .b(gate131inter1), .O(G504));

  xor2  gate841(.a(G417), .b(G416), .O(gate132inter0));
  nand2 gate842(.a(gate132inter0), .b(s_42), .O(gate132inter1));
  and2  gate843(.a(G417), .b(G416), .O(gate132inter2));
  inv1  gate844(.a(s_42), .O(gate132inter3));
  inv1  gate845(.a(s_43), .O(gate132inter4));
  nand2 gate846(.a(gate132inter4), .b(gate132inter3), .O(gate132inter5));
  nor2  gate847(.a(gate132inter5), .b(gate132inter2), .O(gate132inter6));
  inv1  gate848(.a(G416), .O(gate132inter7));
  inv1  gate849(.a(G417), .O(gate132inter8));
  nand2 gate850(.a(gate132inter8), .b(gate132inter7), .O(gate132inter9));
  nand2 gate851(.a(s_43), .b(gate132inter3), .O(gate132inter10));
  nor2  gate852(.a(gate132inter10), .b(gate132inter9), .O(gate132inter11));
  nor2  gate853(.a(gate132inter11), .b(gate132inter6), .O(gate132inter12));
  nand2 gate854(.a(gate132inter12), .b(gate132inter1), .O(G507));
nand2 gate133( .a(G418), .b(G419), .O(G510) );
nand2 gate134( .a(G420), .b(G421), .O(G513) );

  xor2  gate1429(.a(G423), .b(G422), .O(gate135inter0));
  nand2 gate1430(.a(gate135inter0), .b(s_126), .O(gate135inter1));
  and2  gate1431(.a(G423), .b(G422), .O(gate135inter2));
  inv1  gate1432(.a(s_126), .O(gate135inter3));
  inv1  gate1433(.a(s_127), .O(gate135inter4));
  nand2 gate1434(.a(gate135inter4), .b(gate135inter3), .O(gate135inter5));
  nor2  gate1435(.a(gate135inter5), .b(gate135inter2), .O(gate135inter6));
  inv1  gate1436(.a(G422), .O(gate135inter7));
  inv1  gate1437(.a(G423), .O(gate135inter8));
  nand2 gate1438(.a(gate135inter8), .b(gate135inter7), .O(gate135inter9));
  nand2 gate1439(.a(s_127), .b(gate135inter3), .O(gate135inter10));
  nor2  gate1440(.a(gate135inter10), .b(gate135inter9), .O(gate135inter11));
  nor2  gate1441(.a(gate135inter11), .b(gate135inter6), .O(gate135inter12));
  nand2 gate1442(.a(gate135inter12), .b(gate135inter1), .O(G516));

  xor2  gate1261(.a(G425), .b(G424), .O(gate136inter0));
  nand2 gate1262(.a(gate136inter0), .b(s_102), .O(gate136inter1));
  and2  gate1263(.a(G425), .b(G424), .O(gate136inter2));
  inv1  gate1264(.a(s_102), .O(gate136inter3));
  inv1  gate1265(.a(s_103), .O(gate136inter4));
  nand2 gate1266(.a(gate136inter4), .b(gate136inter3), .O(gate136inter5));
  nor2  gate1267(.a(gate136inter5), .b(gate136inter2), .O(gate136inter6));
  inv1  gate1268(.a(G424), .O(gate136inter7));
  inv1  gate1269(.a(G425), .O(gate136inter8));
  nand2 gate1270(.a(gate136inter8), .b(gate136inter7), .O(gate136inter9));
  nand2 gate1271(.a(s_103), .b(gate136inter3), .O(gate136inter10));
  nor2  gate1272(.a(gate136inter10), .b(gate136inter9), .O(gate136inter11));
  nor2  gate1273(.a(gate136inter11), .b(gate136inter6), .O(gate136inter12));
  nand2 gate1274(.a(gate136inter12), .b(gate136inter1), .O(G519));

  xor2  gate575(.a(G429), .b(G426), .O(gate137inter0));
  nand2 gate576(.a(gate137inter0), .b(s_4), .O(gate137inter1));
  and2  gate577(.a(G429), .b(G426), .O(gate137inter2));
  inv1  gate578(.a(s_4), .O(gate137inter3));
  inv1  gate579(.a(s_5), .O(gate137inter4));
  nand2 gate580(.a(gate137inter4), .b(gate137inter3), .O(gate137inter5));
  nor2  gate581(.a(gate137inter5), .b(gate137inter2), .O(gate137inter6));
  inv1  gate582(.a(G426), .O(gate137inter7));
  inv1  gate583(.a(G429), .O(gate137inter8));
  nand2 gate584(.a(gate137inter8), .b(gate137inter7), .O(gate137inter9));
  nand2 gate585(.a(s_5), .b(gate137inter3), .O(gate137inter10));
  nor2  gate586(.a(gate137inter10), .b(gate137inter9), .O(gate137inter11));
  nor2  gate587(.a(gate137inter11), .b(gate137inter6), .O(gate137inter12));
  nand2 gate588(.a(gate137inter12), .b(gate137inter1), .O(G522));
nand2 gate138( .a(G432), .b(G435), .O(G525) );
nand2 gate139( .a(G438), .b(G441), .O(G528) );
nand2 gate140( .a(G444), .b(G447), .O(G531) );
nand2 gate141( .a(G450), .b(G453), .O(G534) );
nand2 gate142( .a(G456), .b(G459), .O(G537) );
nand2 gate143( .a(G462), .b(G465), .O(G540) );

  xor2  gate701(.a(G471), .b(G468), .O(gate144inter0));
  nand2 gate702(.a(gate144inter0), .b(s_22), .O(gate144inter1));
  and2  gate703(.a(G471), .b(G468), .O(gate144inter2));
  inv1  gate704(.a(s_22), .O(gate144inter3));
  inv1  gate705(.a(s_23), .O(gate144inter4));
  nand2 gate706(.a(gate144inter4), .b(gate144inter3), .O(gate144inter5));
  nor2  gate707(.a(gate144inter5), .b(gate144inter2), .O(gate144inter6));
  inv1  gate708(.a(G468), .O(gate144inter7));
  inv1  gate709(.a(G471), .O(gate144inter8));
  nand2 gate710(.a(gate144inter8), .b(gate144inter7), .O(gate144inter9));
  nand2 gate711(.a(s_23), .b(gate144inter3), .O(gate144inter10));
  nor2  gate712(.a(gate144inter10), .b(gate144inter9), .O(gate144inter11));
  nor2  gate713(.a(gate144inter11), .b(gate144inter6), .O(gate144inter12));
  nand2 gate714(.a(gate144inter12), .b(gate144inter1), .O(G543));
nand2 gate145( .a(G474), .b(G477), .O(G546) );
nand2 gate146( .a(G480), .b(G483), .O(G549) );

  xor2  gate1387(.a(G489), .b(G486), .O(gate147inter0));
  nand2 gate1388(.a(gate147inter0), .b(s_120), .O(gate147inter1));
  and2  gate1389(.a(G489), .b(G486), .O(gate147inter2));
  inv1  gate1390(.a(s_120), .O(gate147inter3));
  inv1  gate1391(.a(s_121), .O(gate147inter4));
  nand2 gate1392(.a(gate147inter4), .b(gate147inter3), .O(gate147inter5));
  nor2  gate1393(.a(gate147inter5), .b(gate147inter2), .O(gate147inter6));
  inv1  gate1394(.a(G486), .O(gate147inter7));
  inv1  gate1395(.a(G489), .O(gate147inter8));
  nand2 gate1396(.a(gate147inter8), .b(gate147inter7), .O(gate147inter9));
  nand2 gate1397(.a(s_121), .b(gate147inter3), .O(gate147inter10));
  nor2  gate1398(.a(gate147inter10), .b(gate147inter9), .O(gate147inter11));
  nor2  gate1399(.a(gate147inter11), .b(gate147inter6), .O(gate147inter12));
  nand2 gate1400(.a(gate147inter12), .b(gate147inter1), .O(G552));
nand2 gate148( .a(G492), .b(G495), .O(G555) );
nand2 gate149( .a(G498), .b(G501), .O(G558) );
nand2 gate150( .a(G504), .b(G507), .O(G561) );
nand2 gate151( .a(G510), .b(G513), .O(G564) );
nand2 gate152( .a(G516), .b(G519), .O(G567) );

  xor2  gate1023(.a(G522), .b(G426), .O(gate153inter0));
  nand2 gate1024(.a(gate153inter0), .b(s_68), .O(gate153inter1));
  and2  gate1025(.a(G522), .b(G426), .O(gate153inter2));
  inv1  gate1026(.a(s_68), .O(gate153inter3));
  inv1  gate1027(.a(s_69), .O(gate153inter4));
  nand2 gate1028(.a(gate153inter4), .b(gate153inter3), .O(gate153inter5));
  nor2  gate1029(.a(gate153inter5), .b(gate153inter2), .O(gate153inter6));
  inv1  gate1030(.a(G426), .O(gate153inter7));
  inv1  gate1031(.a(G522), .O(gate153inter8));
  nand2 gate1032(.a(gate153inter8), .b(gate153inter7), .O(gate153inter9));
  nand2 gate1033(.a(s_69), .b(gate153inter3), .O(gate153inter10));
  nor2  gate1034(.a(gate153inter10), .b(gate153inter9), .O(gate153inter11));
  nor2  gate1035(.a(gate153inter11), .b(gate153inter6), .O(gate153inter12));
  nand2 gate1036(.a(gate153inter12), .b(gate153inter1), .O(G570));
nand2 gate154( .a(G429), .b(G522), .O(G571) );
nand2 gate155( .a(G432), .b(G525), .O(G572) );

  xor2  gate1065(.a(G525), .b(G435), .O(gate156inter0));
  nand2 gate1066(.a(gate156inter0), .b(s_74), .O(gate156inter1));
  and2  gate1067(.a(G525), .b(G435), .O(gate156inter2));
  inv1  gate1068(.a(s_74), .O(gate156inter3));
  inv1  gate1069(.a(s_75), .O(gate156inter4));
  nand2 gate1070(.a(gate156inter4), .b(gate156inter3), .O(gate156inter5));
  nor2  gate1071(.a(gate156inter5), .b(gate156inter2), .O(gate156inter6));
  inv1  gate1072(.a(G435), .O(gate156inter7));
  inv1  gate1073(.a(G525), .O(gate156inter8));
  nand2 gate1074(.a(gate156inter8), .b(gate156inter7), .O(gate156inter9));
  nand2 gate1075(.a(s_75), .b(gate156inter3), .O(gate156inter10));
  nor2  gate1076(.a(gate156inter10), .b(gate156inter9), .O(gate156inter11));
  nor2  gate1077(.a(gate156inter11), .b(gate156inter6), .O(gate156inter12));
  nand2 gate1078(.a(gate156inter12), .b(gate156inter1), .O(G573));
nand2 gate157( .a(G438), .b(G528), .O(G574) );

  xor2  gate1443(.a(G528), .b(G441), .O(gate158inter0));
  nand2 gate1444(.a(gate158inter0), .b(s_128), .O(gate158inter1));
  and2  gate1445(.a(G528), .b(G441), .O(gate158inter2));
  inv1  gate1446(.a(s_128), .O(gate158inter3));
  inv1  gate1447(.a(s_129), .O(gate158inter4));
  nand2 gate1448(.a(gate158inter4), .b(gate158inter3), .O(gate158inter5));
  nor2  gate1449(.a(gate158inter5), .b(gate158inter2), .O(gate158inter6));
  inv1  gate1450(.a(G441), .O(gate158inter7));
  inv1  gate1451(.a(G528), .O(gate158inter8));
  nand2 gate1452(.a(gate158inter8), .b(gate158inter7), .O(gate158inter9));
  nand2 gate1453(.a(s_129), .b(gate158inter3), .O(gate158inter10));
  nor2  gate1454(.a(gate158inter10), .b(gate158inter9), .O(gate158inter11));
  nor2  gate1455(.a(gate158inter11), .b(gate158inter6), .O(gate158inter12));
  nand2 gate1456(.a(gate158inter12), .b(gate158inter1), .O(G575));
nand2 gate159( .a(G444), .b(G531), .O(G576) );
nand2 gate160( .a(G447), .b(G531), .O(G577) );
nand2 gate161( .a(G450), .b(G534), .O(G578) );
nand2 gate162( .a(G453), .b(G534), .O(G579) );
nand2 gate163( .a(G456), .b(G537), .O(G580) );
nand2 gate164( .a(G459), .b(G537), .O(G581) );
nand2 gate165( .a(G462), .b(G540), .O(G582) );
nand2 gate166( .a(G465), .b(G540), .O(G583) );
nand2 gate167( .a(G468), .b(G543), .O(G584) );
nand2 gate168( .a(G471), .b(G543), .O(G585) );

  xor2  gate729(.a(G546), .b(G474), .O(gate169inter0));
  nand2 gate730(.a(gate169inter0), .b(s_26), .O(gate169inter1));
  and2  gate731(.a(G546), .b(G474), .O(gate169inter2));
  inv1  gate732(.a(s_26), .O(gate169inter3));
  inv1  gate733(.a(s_27), .O(gate169inter4));
  nand2 gate734(.a(gate169inter4), .b(gate169inter3), .O(gate169inter5));
  nor2  gate735(.a(gate169inter5), .b(gate169inter2), .O(gate169inter6));
  inv1  gate736(.a(G474), .O(gate169inter7));
  inv1  gate737(.a(G546), .O(gate169inter8));
  nand2 gate738(.a(gate169inter8), .b(gate169inter7), .O(gate169inter9));
  nand2 gate739(.a(s_27), .b(gate169inter3), .O(gate169inter10));
  nor2  gate740(.a(gate169inter10), .b(gate169inter9), .O(gate169inter11));
  nor2  gate741(.a(gate169inter11), .b(gate169inter6), .O(gate169inter12));
  nand2 gate742(.a(gate169inter12), .b(gate169inter1), .O(G586));
nand2 gate170( .a(G477), .b(G546), .O(G587) );
nand2 gate171( .a(G480), .b(G549), .O(G588) );
nand2 gate172( .a(G483), .b(G549), .O(G589) );

  xor2  gate743(.a(G552), .b(G486), .O(gate173inter0));
  nand2 gate744(.a(gate173inter0), .b(s_28), .O(gate173inter1));
  and2  gate745(.a(G552), .b(G486), .O(gate173inter2));
  inv1  gate746(.a(s_28), .O(gate173inter3));
  inv1  gate747(.a(s_29), .O(gate173inter4));
  nand2 gate748(.a(gate173inter4), .b(gate173inter3), .O(gate173inter5));
  nor2  gate749(.a(gate173inter5), .b(gate173inter2), .O(gate173inter6));
  inv1  gate750(.a(G486), .O(gate173inter7));
  inv1  gate751(.a(G552), .O(gate173inter8));
  nand2 gate752(.a(gate173inter8), .b(gate173inter7), .O(gate173inter9));
  nand2 gate753(.a(s_29), .b(gate173inter3), .O(gate173inter10));
  nor2  gate754(.a(gate173inter10), .b(gate173inter9), .O(gate173inter11));
  nor2  gate755(.a(gate173inter11), .b(gate173inter6), .O(gate173inter12));
  nand2 gate756(.a(gate173inter12), .b(gate173inter1), .O(G590));
nand2 gate174( .a(G489), .b(G552), .O(G591) );
nand2 gate175( .a(G492), .b(G555), .O(G592) );
nand2 gate176( .a(G495), .b(G555), .O(G593) );
nand2 gate177( .a(G498), .b(G558), .O(G594) );
nand2 gate178( .a(G501), .b(G558), .O(G595) );
nand2 gate179( .a(G504), .b(G561), .O(G596) );
nand2 gate180( .a(G507), .b(G561), .O(G597) );
nand2 gate181( .a(G510), .b(G564), .O(G598) );
nand2 gate182( .a(G513), .b(G564), .O(G599) );
nand2 gate183( .a(G516), .b(G567), .O(G600) );
nand2 gate184( .a(G519), .b(G567), .O(G601) );
nand2 gate185( .a(G570), .b(G571), .O(G602) );
nand2 gate186( .a(G572), .b(G573), .O(G607) );

  xor2  gate1513(.a(G575), .b(G574), .O(gate187inter0));
  nand2 gate1514(.a(gate187inter0), .b(s_138), .O(gate187inter1));
  and2  gate1515(.a(G575), .b(G574), .O(gate187inter2));
  inv1  gate1516(.a(s_138), .O(gate187inter3));
  inv1  gate1517(.a(s_139), .O(gate187inter4));
  nand2 gate1518(.a(gate187inter4), .b(gate187inter3), .O(gate187inter5));
  nor2  gate1519(.a(gate187inter5), .b(gate187inter2), .O(gate187inter6));
  inv1  gate1520(.a(G574), .O(gate187inter7));
  inv1  gate1521(.a(G575), .O(gate187inter8));
  nand2 gate1522(.a(gate187inter8), .b(gate187inter7), .O(gate187inter9));
  nand2 gate1523(.a(s_139), .b(gate187inter3), .O(gate187inter10));
  nor2  gate1524(.a(gate187inter10), .b(gate187inter9), .O(gate187inter11));
  nor2  gate1525(.a(gate187inter11), .b(gate187inter6), .O(gate187inter12));
  nand2 gate1526(.a(gate187inter12), .b(gate187inter1), .O(G612));
nand2 gate188( .a(G576), .b(G577), .O(G617) );
nand2 gate189( .a(G578), .b(G579), .O(G622) );
nand2 gate190( .a(G580), .b(G581), .O(G627) );

  xor2  gate617(.a(G583), .b(G582), .O(gate191inter0));
  nand2 gate618(.a(gate191inter0), .b(s_10), .O(gate191inter1));
  and2  gate619(.a(G583), .b(G582), .O(gate191inter2));
  inv1  gate620(.a(s_10), .O(gate191inter3));
  inv1  gate621(.a(s_11), .O(gate191inter4));
  nand2 gate622(.a(gate191inter4), .b(gate191inter3), .O(gate191inter5));
  nor2  gate623(.a(gate191inter5), .b(gate191inter2), .O(gate191inter6));
  inv1  gate624(.a(G582), .O(gate191inter7));
  inv1  gate625(.a(G583), .O(gate191inter8));
  nand2 gate626(.a(gate191inter8), .b(gate191inter7), .O(gate191inter9));
  nand2 gate627(.a(s_11), .b(gate191inter3), .O(gate191inter10));
  nor2  gate628(.a(gate191inter10), .b(gate191inter9), .O(gate191inter11));
  nor2  gate629(.a(gate191inter11), .b(gate191inter6), .O(gate191inter12));
  nand2 gate630(.a(gate191inter12), .b(gate191inter1), .O(G632));
nand2 gate192( .a(G584), .b(G585), .O(G637) );
nand2 gate193( .a(G586), .b(G587), .O(G642) );
nand2 gate194( .a(G588), .b(G589), .O(G645) );
nand2 gate195( .a(G590), .b(G591), .O(G648) );

  xor2  gate645(.a(G593), .b(G592), .O(gate196inter0));
  nand2 gate646(.a(gate196inter0), .b(s_14), .O(gate196inter1));
  and2  gate647(.a(G593), .b(G592), .O(gate196inter2));
  inv1  gate648(.a(s_14), .O(gate196inter3));
  inv1  gate649(.a(s_15), .O(gate196inter4));
  nand2 gate650(.a(gate196inter4), .b(gate196inter3), .O(gate196inter5));
  nor2  gate651(.a(gate196inter5), .b(gate196inter2), .O(gate196inter6));
  inv1  gate652(.a(G592), .O(gate196inter7));
  inv1  gate653(.a(G593), .O(gate196inter8));
  nand2 gate654(.a(gate196inter8), .b(gate196inter7), .O(gate196inter9));
  nand2 gate655(.a(s_15), .b(gate196inter3), .O(gate196inter10));
  nor2  gate656(.a(gate196inter10), .b(gate196inter9), .O(gate196inter11));
  nor2  gate657(.a(gate196inter11), .b(gate196inter6), .O(gate196inter12));
  nand2 gate658(.a(gate196inter12), .b(gate196inter1), .O(G651));
nand2 gate197( .a(G594), .b(G595), .O(G654) );
nand2 gate198( .a(G596), .b(G597), .O(G657) );
nand2 gate199( .a(G598), .b(G599), .O(G660) );
nand2 gate200( .a(G600), .b(G601), .O(G663) );
nand2 gate201( .a(G602), .b(G607), .O(G666) );
nand2 gate202( .a(G612), .b(G617), .O(G669) );
nand2 gate203( .a(G602), .b(G612), .O(G672) );
nand2 gate204( .a(G607), .b(G617), .O(G675) );
nand2 gate205( .a(G622), .b(G627), .O(G678) );
nand2 gate206( .a(G632), .b(G637), .O(G681) );
nand2 gate207( .a(G622), .b(G632), .O(G684) );

  xor2  gate897(.a(G637), .b(G627), .O(gate208inter0));
  nand2 gate898(.a(gate208inter0), .b(s_50), .O(gate208inter1));
  and2  gate899(.a(G637), .b(G627), .O(gate208inter2));
  inv1  gate900(.a(s_50), .O(gate208inter3));
  inv1  gate901(.a(s_51), .O(gate208inter4));
  nand2 gate902(.a(gate208inter4), .b(gate208inter3), .O(gate208inter5));
  nor2  gate903(.a(gate208inter5), .b(gate208inter2), .O(gate208inter6));
  inv1  gate904(.a(G627), .O(gate208inter7));
  inv1  gate905(.a(G637), .O(gate208inter8));
  nand2 gate906(.a(gate208inter8), .b(gate208inter7), .O(gate208inter9));
  nand2 gate907(.a(s_51), .b(gate208inter3), .O(gate208inter10));
  nor2  gate908(.a(gate208inter10), .b(gate208inter9), .O(gate208inter11));
  nor2  gate909(.a(gate208inter11), .b(gate208inter6), .O(gate208inter12));
  nand2 gate910(.a(gate208inter12), .b(gate208inter1), .O(G687));
nand2 gate209( .a(G602), .b(G666), .O(G690) );
nand2 gate210( .a(G607), .b(G666), .O(G691) );

  xor2  gate785(.a(G669), .b(G612), .O(gate211inter0));
  nand2 gate786(.a(gate211inter0), .b(s_34), .O(gate211inter1));
  and2  gate787(.a(G669), .b(G612), .O(gate211inter2));
  inv1  gate788(.a(s_34), .O(gate211inter3));
  inv1  gate789(.a(s_35), .O(gate211inter4));
  nand2 gate790(.a(gate211inter4), .b(gate211inter3), .O(gate211inter5));
  nor2  gate791(.a(gate211inter5), .b(gate211inter2), .O(gate211inter6));
  inv1  gate792(.a(G612), .O(gate211inter7));
  inv1  gate793(.a(G669), .O(gate211inter8));
  nand2 gate794(.a(gate211inter8), .b(gate211inter7), .O(gate211inter9));
  nand2 gate795(.a(s_35), .b(gate211inter3), .O(gate211inter10));
  nor2  gate796(.a(gate211inter10), .b(gate211inter9), .O(gate211inter11));
  nor2  gate797(.a(gate211inter11), .b(gate211inter6), .O(gate211inter12));
  nand2 gate798(.a(gate211inter12), .b(gate211inter1), .O(G692));
nand2 gate212( .a(G617), .b(G669), .O(G693) );
nand2 gate213( .a(G602), .b(G672), .O(G694) );
nand2 gate214( .a(G612), .b(G672), .O(G695) );
nand2 gate215( .a(G607), .b(G675), .O(G696) );
nand2 gate216( .a(G617), .b(G675), .O(G697) );
nand2 gate217( .a(G622), .b(G678), .O(G698) );
nand2 gate218( .a(G627), .b(G678), .O(G699) );
nand2 gate219( .a(G632), .b(G681), .O(G700) );

  xor2  gate967(.a(G681), .b(G637), .O(gate220inter0));
  nand2 gate968(.a(gate220inter0), .b(s_60), .O(gate220inter1));
  and2  gate969(.a(G681), .b(G637), .O(gate220inter2));
  inv1  gate970(.a(s_60), .O(gate220inter3));
  inv1  gate971(.a(s_61), .O(gate220inter4));
  nand2 gate972(.a(gate220inter4), .b(gate220inter3), .O(gate220inter5));
  nor2  gate973(.a(gate220inter5), .b(gate220inter2), .O(gate220inter6));
  inv1  gate974(.a(G637), .O(gate220inter7));
  inv1  gate975(.a(G681), .O(gate220inter8));
  nand2 gate976(.a(gate220inter8), .b(gate220inter7), .O(gate220inter9));
  nand2 gate977(.a(s_61), .b(gate220inter3), .O(gate220inter10));
  nor2  gate978(.a(gate220inter10), .b(gate220inter9), .O(gate220inter11));
  nor2  gate979(.a(gate220inter11), .b(gate220inter6), .O(gate220inter12));
  nand2 gate980(.a(gate220inter12), .b(gate220inter1), .O(G701));

  xor2  gate827(.a(G684), .b(G622), .O(gate221inter0));
  nand2 gate828(.a(gate221inter0), .b(s_40), .O(gate221inter1));
  and2  gate829(.a(G684), .b(G622), .O(gate221inter2));
  inv1  gate830(.a(s_40), .O(gate221inter3));
  inv1  gate831(.a(s_41), .O(gate221inter4));
  nand2 gate832(.a(gate221inter4), .b(gate221inter3), .O(gate221inter5));
  nor2  gate833(.a(gate221inter5), .b(gate221inter2), .O(gate221inter6));
  inv1  gate834(.a(G622), .O(gate221inter7));
  inv1  gate835(.a(G684), .O(gate221inter8));
  nand2 gate836(.a(gate221inter8), .b(gate221inter7), .O(gate221inter9));
  nand2 gate837(.a(s_41), .b(gate221inter3), .O(gate221inter10));
  nor2  gate838(.a(gate221inter10), .b(gate221inter9), .O(gate221inter11));
  nor2  gate839(.a(gate221inter11), .b(gate221inter6), .O(gate221inter12));
  nand2 gate840(.a(gate221inter12), .b(gate221inter1), .O(G702));
nand2 gate222( .a(G632), .b(G684), .O(G703) );
nand2 gate223( .a(G627), .b(G687), .O(G704) );
nand2 gate224( .a(G637), .b(G687), .O(G705) );
nand2 gate225( .a(G690), .b(G691), .O(G706) );
nand2 gate226( .a(G692), .b(G693), .O(G709) );

  xor2  gate1331(.a(G695), .b(G694), .O(gate227inter0));
  nand2 gate1332(.a(gate227inter0), .b(s_112), .O(gate227inter1));
  and2  gate1333(.a(G695), .b(G694), .O(gate227inter2));
  inv1  gate1334(.a(s_112), .O(gate227inter3));
  inv1  gate1335(.a(s_113), .O(gate227inter4));
  nand2 gate1336(.a(gate227inter4), .b(gate227inter3), .O(gate227inter5));
  nor2  gate1337(.a(gate227inter5), .b(gate227inter2), .O(gate227inter6));
  inv1  gate1338(.a(G694), .O(gate227inter7));
  inv1  gate1339(.a(G695), .O(gate227inter8));
  nand2 gate1340(.a(gate227inter8), .b(gate227inter7), .O(gate227inter9));
  nand2 gate1341(.a(s_113), .b(gate227inter3), .O(gate227inter10));
  nor2  gate1342(.a(gate227inter10), .b(gate227inter9), .O(gate227inter11));
  nor2  gate1343(.a(gate227inter11), .b(gate227inter6), .O(gate227inter12));
  nand2 gate1344(.a(gate227inter12), .b(gate227inter1), .O(G712));
nand2 gate228( .a(G696), .b(G697), .O(G715) );
nand2 gate229( .a(G698), .b(G699), .O(G718) );
nand2 gate230( .a(G700), .b(G701), .O(G721) );
nand2 gate231( .a(G702), .b(G703), .O(G724) );
nand2 gate232( .a(G704), .b(G705), .O(G727) );

  xor2  gate687(.a(G718), .b(G242), .O(gate233inter0));
  nand2 gate688(.a(gate233inter0), .b(s_20), .O(gate233inter1));
  and2  gate689(.a(G718), .b(G242), .O(gate233inter2));
  inv1  gate690(.a(s_20), .O(gate233inter3));
  inv1  gate691(.a(s_21), .O(gate233inter4));
  nand2 gate692(.a(gate233inter4), .b(gate233inter3), .O(gate233inter5));
  nor2  gate693(.a(gate233inter5), .b(gate233inter2), .O(gate233inter6));
  inv1  gate694(.a(G242), .O(gate233inter7));
  inv1  gate695(.a(G718), .O(gate233inter8));
  nand2 gate696(.a(gate233inter8), .b(gate233inter7), .O(gate233inter9));
  nand2 gate697(.a(s_21), .b(gate233inter3), .O(gate233inter10));
  nor2  gate698(.a(gate233inter10), .b(gate233inter9), .O(gate233inter11));
  nor2  gate699(.a(gate233inter11), .b(gate233inter6), .O(gate233inter12));
  nand2 gate700(.a(gate233inter12), .b(gate233inter1), .O(G730));

  xor2  gate1275(.a(G721), .b(G245), .O(gate234inter0));
  nand2 gate1276(.a(gate234inter0), .b(s_104), .O(gate234inter1));
  and2  gate1277(.a(G721), .b(G245), .O(gate234inter2));
  inv1  gate1278(.a(s_104), .O(gate234inter3));
  inv1  gate1279(.a(s_105), .O(gate234inter4));
  nand2 gate1280(.a(gate234inter4), .b(gate234inter3), .O(gate234inter5));
  nor2  gate1281(.a(gate234inter5), .b(gate234inter2), .O(gate234inter6));
  inv1  gate1282(.a(G245), .O(gate234inter7));
  inv1  gate1283(.a(G721), .O(gate234inter8));
  nand2 gate1284(.a(gate234inter8), .b(gate234inter7), .O(gate234inter9));
  nand2 gate1285(.a(s_105), .b(gate234inter3), .O(gate234inter10));
  nor2  gate1286(.a(gate234inter10), .b(gate234inter9), .O(gate234inter11));
  nor2  gate1287(.a(gate234inter11), .b(gate234inter6), .O(gate234inter12));
  nand2 gate1288(.a(gate234inter12), .b(gate234inter1), .O(G733));
nand2 gate235( .a(G248), .b(G724), .O(G736) );
nand2 gate236( .a(G251), .b(G727), .O(G739) );

  xor2  gate1233(.a(G706), .b(G254), .O(gate237inter0));
  nand2 gate1234(.a(gate237inter0), .b(s_98), .O(gate237inter1));
  and2  gate1235(.a(G706), .b(G254), .O(gate237inter2));
  inv1  gate1236(.a(s_98), .O(gate237inter3));
  inv1  gate1237(.a(s_99), .O(gate237inter4));
  nand2 gate1238(.a(gate237inter4), .b(gate237inter3), .O(gate237inter5));
  nor2  gate1239(.a(gate237inter5), .b(gate237inter2), .O(gate237inter6));
  inv1  gate1240(.a(G254), .O(gate237inter7));
  inv1  gate1241(.a(G706), .O(gate237inter8));
  nand2 gate1242(.a(gate237inter8), .b(gate237inter7), .O(gate237inter9));
  nand2 gate1243(.a(s_99), .b(gate237inter3), .O(gate237inter10));
  nor2  gate1244(.a(gate237inter10), .b(gate237inter9), .O(gate237inter11));
  nor2  gate1245(.a(gate237inter11), .b(gate237inter6), .O(gate237inter12));
  nand2 gate1246(.a(gate237inter12), .b(gate237inter1), .O(G742));
nand2 gate238( .a(G257), .b(G709), .O(G745) );

  xor2  gate1009(.a(G712), .b(G260), .O(gate239inter0));
  nand2 gate1010(.a(gate239inter0), .b(s_66), .O(gate239inter1));
  and2  gate1011(.a(G712), .b(G260), .O(gate239inter2));
  inv1  gate1012(.a(s_66), .O(gate239inter3));
  inv1  gate1013(.a(s_67), .O(gate239inter4));
  nand2 gate1014(.a(gate239inter4), .b(gate239inter3), .O(gate239inter5));
  nor2  gate1015(.a(gate239inter5), .b(gate239inter2), .O(gate239inter6));
  inv1  gate1016(.a(G260), .O(gate239inter7));
  inv1  gate1017(.a(G712), .O(gate239inter8));
  nand2 gate1018(.a(gate239inter8), .b(gate239inter7), .O(gate239inter9));
  nand2 gate1019(.a(s_67), .b(gate239inter3), .O(gate239inter10));
  nor2  gate1020(.a(gate239inter10), .b(gate239inter9), .O(gate239inter11));
  nor2  gate1021(.a(gate239inter11), .b(gate239inter6), .O(gate239inter12));
  nand2 gate1022(.a(gate239inter12), .b(gate239inter1), .O(G748));
nand2 gate240( .a(G263), .b(G715), .O(G751) );
nand2 gate241( .a(G242), .b(G730), .O(G754) );
nand2 gate242( .a(G718), .b(G730), .O(G755) );

  xor2  gate869(.a(G733), .b(G245), .O(gate243inter0));
  nand2 gate870(.a(gate243inter0), .b(s_46), .O(gate243inter1));
  and2  gate871(.a(G733), .b(G245), .O(gate243inter2));
  inv1  gate872(.a(s_46), .O(gate243inter3));
  inv1  gate873(.a(s_47), .O(gate243inter4));
  nand2 gate874(.a(gate243inter4), .b(gate243inter3), .O(gate243inter5));
  nor2  gate875(.a(gate243inter5), .b(gate243inter2), .O(gate243inter6));
  inv1  gate876(.a(G245), .O(gate243inter7));
  inv1  gate877(.a(G733), .O(gate243inter8));
  nand2 gate878(.a(gate243inter8), .b(gate243inter7), .O(gate243inter9));
  nand2 gate879(.a(s_47), .b(gate243inter3), .O(gate243inter10));
  nor2  gate880(.a(gate243inter10), .b(gate243inter9), .O(gate243inter11));
  nor2  gate881(.a(gate243inter11), .b(gate243inter6), .O(gate243inter12));
  nand2 gate882(.a(gate243inter12), .b(gate243inter1), .O(G756));
nand2 gate244( .a(G721), .b(G733), .O(G757) );
nand2 gate245( .a(G248), .b(G736), .O(G758) );
nand2 gate246( .a(G724), .b(G736), .O(G759) );
nand2 gate247( .a(G251), .b(G739), .O(G760) );
nand2 gate248( .a(G727), .b(G739), .O(G761) );
nand2 gate249( .a(G254), .b(G742), .O(G762) );
nand2 gate250( .a(G706), .b(G742), .O(G763) );
nand2 gate251( .a(G257), .b(G745), .O(G764) );
nand2 gate252( .a(G709), .b(G745), .O(G765) );
nand2 gate253( .a(G260), .b(G748), .O(G766) );
nand2 gate254( .a(G712), .b(G748), .O(G767) );
nand2 gate255( .a(G263), .b(G751), .O(G768) );
nand2 gate256( .a(G715), .b(G751), .O(G769) );
nand2 gate257( .a(G754), .b(G755), .O(G770) );
nand2 gate258( .a(G756), .b(G757), .O(G773) );
nand2 gate259( .a(G758), .b(G759), .O(G776) );
nand2 gate260( .a(G760), .b(G761), .O(G779) );

  xor2  gate1471(.a(G763), .b(G762), .O(gate261inter0));
  nand2 gate1472(.a(gate261inter0), .b(s_132), .O(gate261inter1));
  and2  gate1473(.a(G763), .b(G762), .O(gate261inter2));
  inv1  gate1474(.a(s_132), .O(gate261inter3));
  inv1  gate1475(.a(s_133), .O(gate261inter4));
  nand2 gate1476(.a(gate261inter4), .b(gate261inter3), .O(gate261inter5));
  nor2  gate1477(.a(gate261inter5), .b(gate261inter2), .O(gate261inter6));
  inv1  gate1478(.a(G762), .O(gate261inter7));
  inv1  gate1479(.a(G763), .O(gate261inter8));
  nand2 gate1480(.a(gate261inter8), .b(gate261inter7), .O(gate261inter9));
  nand2 gate1481(.a(s_133), .b(gate261inter3), .O(gate261inter10));
  nor2  gate1482(.a(gate261inter10), .b(gate261inter9), .O(gate261inter11));
  nor2  gate1483(.a(gate261inter11), .b(gate261inter6), .O(gate261inter12));
  nand2 gate1484(.a(gate261inter12), .b(gate261inter1), .O(G782));
nand2 gate262( .a(G764), .b(G765), .O(G785) );
nand2 gate263( .a(G766), .b(G767), .O(G788) );
nand2 gate264( .a(G768), .b(G769), .O(G791) );
nand2 gate265( .a(G642), .b(G770), .O(G794) );
nand2 gate266( .a(G645), .b(G773), .O(G797) );
nand2 gate267( .a(G648), .b(G776), .O(G800) );
nand2 gate268( .a(G651), .b(G779), .O(G803) );
nand2 gate269( .a(G654), .b(G782), .O(G806) );
nand2 gate270( .a(G657), .b(G785), .O(G809) );

  xor2  gate1163(.a(G788), .b(G660), .O(gate271inter0));
  nand2 gate1164(.a(gate271inter0), .b(s_88), .O(gate271inter1));
  and2  gate1165(.a(G788), .b(G660), .O(gate271inter2));
  inv1  gate1166(.a(s_88), .O(gate271inter3));
  inv1  gate1167(.a(s_89), .O(gate271inter4));
  nand2 gate1168(.a(gate271inter4), .b(gate271inter3), .O(gate271inter5));
  nor2  gate1169(.a(gate271inter5), .b(gate271inter2), .O(gate271inter6));
  inv1  gate1170(.a(G660), .O(gate271inter7));
  inv1  gate1171(.a(G788), .O(gate271inter8));
  nand2 gate1172(.a(gate271inter8), .b(gate271inter7), .O(gate271inter9));
  nand2 gate1173(.a(s_89), .b(gate271inter3), .O(gate271inter10));
  nor2  gate1174(.a(gate271inter10), .b(gate271inter9), .O(gate271inter11));
  nor2  gate1175(.a(gate271inter11), .b(gate271inter6), .O(gate271inter12));
  nand2 gate1176(.a(gate271inter12), .b(gate271inter1), .O(G812));
nand2 gate272( .a(G663), .b(G791), .O(G815) );
nand2 gate273( .a(G642), .b(G794), .O(G818) );

  xor2  gate1121(.a(G794), .b(G770), .O(gate274inter0));
  nand2 gate1122(.a(gate274inter0), .b(s_82), .O(gate274inter1));
  and2  gate1123(.a(G794), .b(G770), .O(gate274inter2));
  inv1  gate1124(.a(s_82), .O(gate274inter3));
  inv1  gate1125(.a(s_83), .O(gate274inter4));
  nand2 gate1126(.a(gate274inter4), .b(gate274inter3), .O(gate274inter5));
  nor2  gate1127(.a(gate274inter5), .b(gate274inter2), .O(gate274inter6));
  inv1  gate1128(.a(G770), .O(gate274inter7));
  inv1  gate1129(.a(G794), .O(gate274inter8));
  nand2 gate1130(.a(gate274inter8), .b(gate274inter7), .O(gate274inter9));
  nand2 gate1131(.a(s_83), .b(gate274inter3), .O(gate274inter10));
  nor2  gate1132(.a(gate274inter10), .b(gate274inter9), .O(gate274inter11));
  nor2  gate1133(.a(gate274inter11), .b(gate274inter6), .O(gate274inter12));
  nand2 gate1134(.a(gate274inter12), .b(gate274inter1), .O(G819));
nand2 gate275( .a(G645), .b(G797), .O(G820) );
nand2 gate276( .a(G773), .b(G797), .O(G821) );
nand2 gate277( .a(G648), .b(G800), .O(G822) );

  xor2  gate1345(.a(G800), .b(G776), .O(gate278inter0));
  nand2 gate1346(.a(gate278inter0), .b(s_114), .O(gate278inter1));
  and2  gate1347(.a(G800), .b(G776), .O(gate278inter2));
  inv1  gate1348(.a(s_114), .O(gate278inter3));
  inv1  gate1349(.a(s_115), .O(gate278inter4));
  nand2 gate1350(.a(gate278inter4), .b(gate278inter3), .O(gate278inter5));
  nor2  gate1351(.a(gate278inter5), .b(gate278inter2), .O(gate278inter6));
  inv1  gate1352(.a(G776), .O(gate278inter7));
  inv1  gate1353(.a(G800), .O(gate278inter8));
  nand2 gate1354(.a(gate278inter8), .b(gate278inter7), .O(gate278inter9));
  nand2 gate1355(.a(s_115), .b(gate278inter3), .O(gate278inter10));
  nor2  gate1356(.a(gate278inter10), .b(gate278inter9), .O(gate278inter11));
  nor2  gate1357(.a(gate278inter11), .b(gate278inter6), .O(gate278inter12));
  nand2 gate1358(.a(gate278inter12), .b(gate278inter1), .O(G823));
nand2 gate279( .a(G651), .b(G803), .O(G824) );
nand2 gate280( .a(G779), .b(G803), .O(G825) );
nand2 gate281( .a(G654), .b(G806), .O(G826) );
nand2 gate282( .a(G782), .b(G806), .O(G827) );

  xor2  gate1219(.a(G809), .b(G657), .O(gate283inter0));
  nand2 gate1220(.a(gate283inter0), .b(s_96), .O(gate283inter1));
  and2  gate1221(.a(G809), .b(G657), .O(gate283inter2));
  inv1  gate1222(.a(s_96), .O(gate283inter3));
  inv1  gate1223(.a(s_97), .O(gate283inter4));
  nand2 gate1224(.a(gate283inter4), .b(gate283inter3), .O(gate283inter5));
  nor2  gate1225(.a(gate283inter5), .b(gate283inter2), .O(gate283inter6));
  inv1  gate1226(.a(G657), .O(gate283inter7));
  inv1  gate1227(.a(G809), .O(gate283inter8));
  nand2 gate1228(.a(gate283inter8), .b(gate283inter7), .O(gate283inter9));
  nand2 gate1229(.a(s_97), .b(gate283inter3), .O(gate283inter10));
  nor2  gate1230(.a(gate283inter10), .b(gate283inter9), .O(gate283inter11));
  nor2  gate1231(.a(gate283inter11), .b(gate283inter6), .O(gate283inter12));
  nand2 gate1232(.a(gate283inter12), .b(gate283inter1), .O(G828));
nand2 gate284( .a(G785), .b(G809), .O(G829) );
nand2 gate285( .a(G660), .b(G812), .O(G830) );

  xor2  gate1373(.a(G812), .b(G788), .O(gate286inter0));
  nand2 gate1374(.a(gate286inter0), .b(s_118), .O(gate286inter1));
  and2  gate1375(.a(G812), .b(G788), .O(gate286inter2));
  inv1  gate1376(.a(s_118), .O(gate286inter3));
  inv1  gate1377(.a(s_119), .O(gate286inter4));
  nand2 gate1378(.a(gate286inter4), .b(gate286inter3), .O(gate286inter5));
  nor2  gate1379(.a(gate286inter5), .b(gate286inter2), .O(gate286inter6));
  inv1  gate1380(.a(G788), .O(gate286inter7));
  inv1  gate1381(.a(G812), .O(gate286inter8));
  nand2 gate1382(.a(gate286inter8), .b(gate286inter7), .O(gate286inter9));
  nand2 gate1383(.a(s_119), .b(gate286inter3), .O(gate286inter10));
  nor2  gate1384(.a(gate286inter10), .b(gate286inter9), .O(gate286inter11));
  nor2  gate1385(.a(gate286inter11), .b(gate286inter6), .O(gate286inter12));
  nand2 gate1386(.a(gate286inter12), .b(gate286inter1), .O(G831));
nand2 gate287( .a(G663), .b(G815), .O(G832) );
nand2 gate288( .a(G791), .b(G815), .O(G833) );
nand2 gate289( .a(G818), .b(G819), .O(G834) );
nand2 gate290( .a(G820), .b(G821), .O(G847) );
nand2 gate291( .a(G822), .b(G823), .O(G860) );
nand2 gate292( .a(G824), .b(G825), .O(G873) );
nand2 gate293( .a(G828), .b(G829), .O(G886) );

  xor2  gate1583(.a(G833), .b(G832), .O(gate294inter0));
  nand2 gate1584(.a(gate294inter0), .b(s_148), .O(gate294inter1));
  and2  gate1585(.a(G833), .b(G832), .O(gate294inter2));
  inv1  gate1586(.a(s_148), .O(gate294inter3));
  inv1  gate1587(.a(s_149), .O(gate294inter4));
  nand2 gate1588(.a(gate294inter4), .b(gate294inter3), .O(gate294inter5));
  nor2  gate1589(.a(gate294inter5), .b(gate294inter2), .O(gate294inter6));
  inv1  gate1590(.a(G832), .O(gate294inter7));
  inv1  gate1591(.a(G833), .O(gate294inter8));
  nand2 gate1592(.a(gate294inter8), .b(gate294inter7), .O(gate294inter9));
  nand2 gate1593(.a(s_149), .b(gate294inter3), .O(gate294inter10));
  nor2  gate1594(.a(gate294inter10), .b(gate294inter9), .O(gate294inter11));
  nor2  gate1595(.a(gate294inter11), .b(gate294inter6), .O(gate294inter12));
  nand2 gate1596(.a(gate294inter12), .b(gate294inter1), .O(G899));
nand2 gate295( .a(G830), .b(G831), .O(G912) );

  xor2  gate1037(.a(G827), .b(G826), .O(gate296inter0));
  nand2 gate1038(.a(gate296inter0), .b(s_70), .O(gate296inter1));
  and2  gate1039(.a(G827), .b(G826), .O(gate296inter2));
  inv1  gate1040(.a(s_70), .O(gate296inter3));
  inv1  gate1041(.a(s_71), .O(gate296inter4));
  nand2 gate1042(.a(gate296inter4), .b(gate296inter3), .O(gate296inter5));
  nor2  gate1043(.a(gate296inter5), .b(gate296inter2), .O(gate296inter6));
  inv1  gate1044(.a(G826), .O(gate296inter7));
  inv1  gate1045(.a(G827), .O(gate296inter8));
  nand2 gate1046(.a(gate296inter8), .b(gate296inter7), .O(gate296inter9));
  nand2 gate1047(.a(s_71), .b(gate296inter3), .O(gate296inter10));
  nor2  gate1048(.a(gate296inter10), .b(gate296inter9), .O(gate296inter11));
  nor2  gate1049(.a(gate296inter11), .b(gate296inter6), .O(gate296inter12));
  nand2 gate1050(.a(gate296inter12), .b(gate296inter1), .O(G925));
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );
nand2 gate387( .a(G1), .b(G1036), .O(G1132) );
nand2 gate388( .a(G2), .b(G1039), .O(G1135) );
nand2 gate389( .a(G3), .b(G1042), .O(G1138) );

  xor2  gate1079(.a(G1045), .b(G4), .O(gate390inter0));
  nand2 gate1080(.a(gate390inter0), .b(s_76), .O(gate390inter1));
  and2  gate1081(.a(G1045), .b(G4), .O(gate390inter2));
  inv1  gate1082(.a(s_76), .O(gate390inter3));
  inv1  gate1083(.a(s_77), .O(gate390inter4));
  nand2 gate1084(.a(gate390inter4), .b(gate390inter3), .O(gate390inter5));
  nor2  gate1085(.a(gate390inter5), .b(gate390inter2), .O(gate390inter6));
  inv1  gate1086(.a(G4), .O(gate390inter7));
  inv1  gate1087(.a(G1045), .O(gate390inter8));
  nand2 gate1088(.a(gate390inter8), .b(gate390inter7), .O(gate390inter9));
  nand2 gate1089(.a(s_77), .b(gate390inter3), .O(gate390inter10));
  nor2  gate1090(.a(gate390inter10), .b(gate390inter9), .O(gate390inter11));
  nor2  gate1091(.a(gate390inter11), .b(gate390inter6), .O(gate390inter12));
  nand2 gate1092(.a(gate390inter12), .b(gate390inter1), .O(G1141));

  xor2  gate813(.a(G1048), .b(G5), .O(gate391inter0));
  nand2 gate814(.a(gate391inter0), .b(s_38), .O(gate391inter1));
  and2  gate815(.a(G1048), .b(G5), .O(gate391inter2));
  inv1  gate816(.a(s_38), .O(gate391inter3));
  inv1  gate817(.a(s_39), .O(gate391inter4));
  nand2 gate818(.a(gate391inter4), .b(gate391inter3), .O(gate391inter5));
  nor2  gate819(.a(gate391inter5), .b(gate391inter2), .O(gate391inter6));
  inv1  gate820(.a(G5), .O(gate391inter7));
  inv1  gate821(.a(G1048), .O(gate391inter8));
  nand2 gate822(.a(gate391inter8), .b(gate391inter7), .O(gate391inter9));
  nand2 gate823(.a(s_39), .b(gate391inter3), .O(gate391inter10));
  nor2  gate824(.a(gate391inter10), .b(gate391inter9), .O(gate391inter11));
  nor2  gate825(.a(gate391inter11), .b(gate391inter6), .O(gate391inter12));
  nand2 gate826(.a(gate391inter12), .b(gate391inter1), .O(G1144));
nand2 gate392( .a(G6), .b(G1051), .O(G1147) );
nand2 gate393( .a(G7), .b(G1054), .O(G1150) );
nand2 gate394( .a(G8), .b(G1057), .O(G1153) );

  xor2  gate953(.a(G1060), .b(G9), .O(gate395inter0));
  nand2 gate954(.a(gate395inter0), .b(s_58), .O(gate395inter1));
  and2  gate955(.a(G1060), .b(G9), .O(gate395inter2));
  inv1  gate956(.a(s_58), .O(gate395inter3));
  inv1  gate957(.a(s_59), .O(gate395inter4));
  nand2 gate958(.a(gate395inter4), .b(gate395inter3), .O(gate395inter5));
  nor2  gate959(.a(gate395inter5), .b(gate395inter2), .O(gate395inter6));
  inv1  gate960(.a(G9), .O(gate395inter7));
  inv1  gate961(.a(G1060), .O(gate395inter8));
  nand2 gate962(.a(gate395inter8), .b(gate395inter7), .O(gate395inter9));
  nand2 gate963(.a(s_59), .b(gate395inter3), .O(gate395inter10));
  nor2  gate964(.a(gate395inter10), .b(gate395inter9), .O(gate395inter11));
  nor2  gate965(.a(gate395inter11), .b(gate395inter6), .O(gate395inter12));
  nand2 gate966(.a(gate395inter12), .b(gate395inter1), .O(G1156));
nand2 gate396( .a(G10), .b(G1063), .O(G1159) );
nand2 gate397( .a(G11), .b(G1066), .O(G1162) );
nand2 gate398( .a(G12), .b(G1069), .O(G1165) );
nand2 gate399( .a(G13), .b(G1072), .O(G1168) );
nand2 gate400( .a(G14), .b(G1075), .O(G1171) );
nand2 gate401( .a(G15), .b(G1078), .O(G1174) );

  xor2  gate561(.a(G1081), .b(G16), .O(gate402inter0));
  nand2 gate562(.a(gate402inter0), .b(s_2), .O(gate402inter1));
  and2  gate563(.a(G1081), .b(G16), .O(gate402inter2));
  inv1  gate564(.a(s_2), .O(gate402inter3));
  inv1  gate565(.a(s_3), .O(gate402inter4));
  nand2 gate566(.a(gate402inter4), .b(gate402inter3), .O(gate402inter5));
  nor2  gate567(.a(gate402inter5), .b(gate402inter2), .O(gate402inter6));
  inv1  gate568(.a(G16), .O(gate402inter7));
  inv1  gate569(.a(G1081), .O(gate402inter8));
  nand2 gate570(.a(gate402inter8), .b(gate402inter7), .O(gate402inter9));
  nand2 gate571(.a(s_3), .b(gate402inter3), .O(gate402inter10));
  nor2  gate572(.a(gate402inter10), .b(gate402inter9), .O(gate402inter11));
  nor2  gate573(.a(gate402inter11), .b(gate402inter6), .O(gate402inter12));
  nand2 gate574(.a(gate402inter12), .b(gate402inter1), .O(G1177));
nand2 gate403( .a(G17), .b(G1084), .O(G1180) );
nand2 gate404( .a(G18), .b(G1087), .O(G1183) );

  xor2  gate1457(.a(G1090), .b(G19), .O(gate405inter0));
  nand2 gate1458(.a(gate405inter0), .b(s_130), .O(gate405inter1));
  and2  gate1459(.a(G1090), .b(G19), .O(gate405inter2));
  inv1  gate1460(.a(s_130), .O(gate405inter3));
  inv1  gate1461(.a(s_131), .O(gate405inter4));
  nand2 gate1462(.a(gate405inter4), .b(gate405inter3), .O(gate405inter5));
  nor2  gate1463(.a(gate405inter5), .b(gate405inter2), .O(gate405inter6));
  inv1  gate1464(.a(G19), .O(gate405inter7));
  inv1  gate1465(.a(G1090), .O(gate405inter8));
  nand2 gate1466(.a(gate405inter8), .b(gate405inter7), .O(gate405inter9));
  nand2 gate1467(.a(s_131), .b(gate405inter3), .O(gate405inter10));
  nor2  gate1468(.a(gate405inter10), .b(gate405inter9), .O(gate405inter11));
  nor2  gate1469(.a(gate405inter11), .b(gate405inter6), .O(gate405inter12));
  nand2 gate1470(.a(gate405inter12), .b(gate405inter1), .O(G1186));
nand2 gate406( .a(G20), .b(G1093), .O(G1189) );
nand2 gate407( .a(G21), .b(G1096), .O(G1192) );
nand2 gate408( .a(G22), .b(G1099), .O(G1195) );
nand2 gate409( .a(G23), .b(G1102), .O(G1198) );

  xor2  gate981(.a(G1105), .b(G24), .O(gate410inter0));
  nand2 gate982(.a(gate410inter0), .b(s_62), .O(gate410inter1));
  and2  gate983(.a(G1105), .b(G24), .O(gate410inter2));
  inv1  gate984(.a(s_62), .O(gate410inter3));
  inv1  gate985(.a(s_63), .O(gate410inter4));
  nand2 gate986(.a(gate410inter4), .b(gate410inter3), .O(gate410inter5));
  nor2  gate987(.a(gate410inter5), .b(gate410inter2), .O(gate410inter6));
  inv1  gate988(.a(G24), .O(gate410inter7));
  inv1  gate989(.a(G1105), .O(gate410inter8));
  nand2 gate990(.a(gate410inter8), .b(gate410inter7), .O(gate410inter9));
  nand2 gate991(.a(s_63), .b(gate410inter3), .O(gate410inter10));
  nor2  gate992(.a(gate410inter10), .b(gate410inter9), .O(gate410inter11));
  nor2  gate993(.a(gate410inter11), .b(gate410inter6), .O(gate410inter12));
  nand2 gate994(.a(gate410inter12), .b(gate410inter1), .O(G1201));
nand2 gate411( .a(G25), .b(G1108), .O(G1204) );
nand2 gate412( .a(G26), .b(G1111), .O(G1207) );
nand2 gate413( .a(G27), .b(G1114), .O(G1210) );
nand2 gate414( .a(G28), .b(G1117), .O(G1213) );

  xor2  gate1135(.a(G1120), .b(G29), .O(gate415inter0));
  nand2 gate1136(.a(gate415inter0), .b(s_84), .O(gate415inter1));
  and2  gate1137(.a(G1120), .b(G29), .O(gate415inter2));
  inv1  gate1138(.a(s_84), .O(gate415inter3));
  inv1  gate1139(.a(s_85), .O(gate415inter4));
  nand2 gate1140(.a(gate415inter4), .b(gate415inter3), .O(gate415inter5));
  nor2  gate1141(.a(gate415inter5), .b(gate415inter2), .O(gate415inter6));
  inv1  gate1142(.a(G29), .O(gate415inter7));
  inv1  gate1143(.a(G1120), .O(gate415inter8));
  nand2 gate1144(.a(gate415inter8), .b(gate415inter7), .O(gate415inter9));
  nand2 gate1145(.a(s_85), .b(gate415inter3), .O(gate415inter10));
  nor2  gate1146(.a(gate415inter10), .b(gate415inter9), .O(gate415inter11));
  nor2  gate1147(.a(gate415inter11), .b(gate415inter6), .O(gate415inter12));
  nand2 gate1148(.a(gate415inter12), .b(gate415inter1), .O(G1216));

  xor2  gate1051(.a(G1123), .b(G30), .O(gate416inter0));
  nand2 gate1052(.a(gate416inter0), .b(s_72), .O(gate416inter1));
  and2  gate1053(.a(G1123), .b(G30), .O(gate416inter2));
  inv1  gate1054(.a(s_72), .O(gate416inter3));
  inv1  gate1055(.a(s_73), .O(gate416inter4));
  nand2 gate1056(.a(gate416inter4), .b(gate416inter3), .O(gate416inter5));
  nor2  gate1057(.a(gate416inter5), .b(gate416inter2), .O(gate416inter6));
  inv1  gate1058(.a(G30), .O(gate416inter7));
  inv1  gate1059(.a(G1123), .O(gate416inter8));
  nand2 gate1060(.a(gate416inter8), .b(gate416inter7), .O(gate416inter9));
  nand2 gate1061(.a(s_73), .b(gate416inter3), .O(gate416inter10));
  nor2  gate1062(.a(gate416inter10), .b(gate416inter9), .O(gate416inter11));
  nor2  gate1063(.a(gate416inter11), .b(gate416inter6), .O(gate416inter12));
  nand2 gate1064(.a(gate416inter12), .b(gate416inter1), .O(G1219));

  xor2  gate1205(.a(G1126), .b(G31), .O(gate417inter0));
  nand2 gate1206(.a(gate417inter0), .b(s_94), .O(gate417inter1));
  and2  gate1207(.a(G1126), .b(G31), .O(gate417inter2));
  inv1  gate1208(.a(s_94), .O(gate417inter3));
  inv1  gate1209(.a(s_95), .O(gate417inter4));
  nand2 gate1210(.a(gate417inter4), .b(gate417inter3), .O(gate417inter5));
  nor2  gate1211(.a(gate417inter5), .b(gate417inter2), .O(gate417inter6));
  inv1  gate1212(.a(G31), .O(gate417inter7));
  inv1  gate1213(.a(G1126), .O(gate417inter8));
  nand2 gate1214(.a(gate417inter8), .b(gate417inter7), .O(gate417inter9));
  nand2 gate1215(.a(s_95), .b(gate417inter3), .O(gate417inter10));
  nor2  gate1216(.a(gate417inter10), .b(gate417inter9), .O(gate417inter11));
  nor2  gate1217(.a(gate417inter11), .b(gate417inter6), .O(gate417inter12));
  nand2 gate1218(.a(gate417inter12), .b(gate417inter1), .O(G1222));

  xor2  gate1527(.a(G1129), .b(G32), .O(gate418inter0));
  nand2 gate1528(.a(gate418inter0), .b(s_140), .O(gate418inter1));
  and2  gate1529(.a(G1129), .b(G32), .O(gate418inter2));
  inv1  gate1530(.a(s_140), .O(gate418inter3));
  inv1  gate1531(.a(s_141), .O(gate418inter4));
  nand2 gate1532(.a(gate418inter4), .b(gate418inter3), .O(gate418inter5));
  nor2  gate1533(.a(gate418inter5), .b(gate418inter2), .O(gate418inter6));
  inv1  gate1534(.a(G32), .O(gate418inter7));
  inv1  gate1535(.a(G1129), .O(gate418inter8));
  nand2 gate1536(.a(gate418inter8), .b(gate418inter7), .O(gate418inter9));
  nand2 gate1537(.a(s_141), .b(gate418inter3), .O(gate418inter10));
  nor2  gate1538(.a(gate418inter10), .b(gate418inter9), .O(gate418inter11));
  nor2  gate1539(.a(gate418inter11), .b(gate418inter6), .O(gate418inter12));
  nand2 gate1540(.a(gate418inter12), .b(gate418inter1), .O(G1225));

  xor2  gate1303(.a(G1132), .b(G1), .O(gate419inter0));
  nand2 gate1304(.a(gate419inter0), .b(s_108), .O(gate419inter1));
  and2  gate1305(.a(G1132), .b(G1), .O(gate419inter2));
  inv1  gate1306(.a(s_108), .O(gate419inter3));
  inv1  gate1307(.a(s_109), .O(gate419inter4));
  nand2 gate1308(.a(gate419inter4), .b(gate419inter3), .O(gate419inter5));
  nor2  gate1309(.a(gate419inter5), .b(gate419inter2), .O(gate419inter6));
  inv1  gate1310(.a(G1), .O(gate419inter7));
  inv1  gate1311(.a(G1132), .O(gate419inter8));
  nand2 gate1312(.a(gate419inter8), .b(gate419inter7), .O(gate419inter9));
  nand2 gate1313(.a(s_109), .b(gate419inter3), .O(gate419inter10));
  nor2  gate1314(.a(gate419inter10), .b(gate419inter9), .O(gate419inter11));
  nor2  gate1315(.a(gate419inter11), .b(gate419inter6), .O(gate419inter12));
  nand2 gate1316(.a(gate419inter12), .b(gate419inter1), .O(G1228));
nand2 gate420( .a(G1036), .b(G1132), .O(G1229) );
nand2 gate421( .a(G2), .b(G1135), .O(G1230) );
nand2 gate422( .a(G1039), .b(G1135), .O(G1231) );
nand2 gate423( .a(G3), .b(G1138), .O(G1232) );
nand2 gate424( .a(G1042), .b(G1138), .O(G1233) );

  xor2  gate1569(.a(G1141), .b(G4), .O(gate425inter0));
  nand2 gate1570(.a(gate425inter0), .b(s_146), .O(gate425inter1));
  and2  gate1571(.a(G1141), .b(G4), .O(gate425inter2));
  inv1  gate1572(.a(s_146), .O(gate425inter3));
  inv1  gate1573(.a(s_147), .O(gate425inter4));
  nand2 gate1574(.a(gate425inter4), .b(gate425inter3), .O(gate425inter5));
  nor2  gate1575(.a(gate425inter5), .b(gate425inter2), .O(gate425inter6));
  inv1  gate1576(.a(G4), .O(gate425inter7));
  inv1  gate1577(.a(G1141), .O(gate425inter8));
  nand2 gate1578(.a(gate425inter8), .b(gate425inter7), .O(gate425inter9));
  nand2 gate1579(.a(s_147), .b(gate425inter3), .O(gate425inter10));
  nor2  gate1580(.a(gate425inter10), .b(gate425inter9), .O(gate425inter11));
  nor2  gate1581(.a(gate425inter11), .b(gate425inter6), .O(gate425inter12));
  nand2 gate1582(.a(gate425inter12), .b(gate425inter1), .O(G1234));
nand2 gate426( .a(G1045), .b(G1141), .O(G1235) );
nand2 gate427( .a(G5), .b(G1144), .O(G1236) );
nand2 gate428( .a(G1048), .b(G1144), .O(G1237) );
nand2 gate429( .a(G6), .b(G1147), .O(G1238) );
nand2 gate430( .a(G1051), .b(G1147), .O(G1239) );

  xor2  gate603(.a(G1150), .b(G7), .O(gate431inter0));
  nand2 gate604(.a(gate431inter0), .b(s_8), .O(gate431inter1));
  and2  gate605(.a(G1150), .b(G7), .O(gate431inter2));
  inv1  gate606(.a(s_8), .O(gate431inter3));
  inv1  gate607(.a(s_9), .O(gate431inter4));
  nand2 gate608(.a(gate431inter4), .b(gate431inter3), .O(gate431inter5));
  nor2  gate609(.a(gate431inter5), .b(gate431inter2), .O(gate431inter6));
  inv1  gate610(.a(G7), .O(gate431inter7));
  inv1  gate611(.a(G1150), .O(gate431inter8));
  nand2 gate612(.a(gate431inter8), .b(gate431inter7), .O(gate431inter9));
  nand2 gate613(.a(s_9), .b(gate431inter3), .O(gate431inter10));
  nor2  gate614(.a(gate431inter10), .b(gate431inter9), .O(gate431inter11));
  nor2  gate615(.a(gate431inter11), .b(gate431inter6), .O(gate431inter12));
  nand2 gate616(.a(gate431inter12), .b(gate431inter1), .O(G1240));
nand2 gate432( .a(G1054), .b(G1150), .O(G1241) );

  xor2  gate1247(.a(G1153), .b(G8), .O(gate433inter0));
  nand2 gate1248(.a(gate433inter0), .b(s_100), .O(gate433inter1));
  and2  gate1249(.a(G1153), .b(G8), .O(gate433inter2));
  inv1  gate1250(.a(s_100), .O(gate433inter3));
  inv1  gate1251(.a(s_101), .O(gate433inter4));
  nand2 gate1252(.a(gate433inter4), .b(gate433inter3), .O(gate433inter5));
  nor2  gate1253(.a(gate433inter5), .b(gate433inter2), .O(gate433inter6));
  inv1  gate1254(.a(G8), .O(gate433inter7));
  inv1  gate1255(.a(G1153), .O(gate433inter8));
  nand2 gate1256(.a(gate433inter8), .b(gate433inter7), .O(gate433inter9));
  nand2 gate1257(.a(s_101), .b(gate433inter3), .O(gate433inter10));
  nor2  gate1258(.a(gate433inter10), .b(gate433inter9), .O(gate433inter11));
  nor2  gate1259(.a(gate433inter11), .b(gate433inter6), .O(gate433inter12));
  nand2 gate1260(.a(gate433inter12), .b(gate433inter1), .O(G1242));
nand2 gate434( .a(G1057), .b(G1153), .O(G1243) );
nand2 gate435( .a(G9), .b(G1156), .O(G1244) );
nand2 gate436( .a(G1060), .b(G1156), .O(G1245) );
nand2 gate437( .a(G10), .b(G1159), .O(G1246) );
nand2 gate438( .a(G1063), .b(G1159), .O(G1247) );
nand2 gate439( .a(G11), .b(G1162), .O(G1248) );
nand2 gate440( .a(G1066), .b(G1162), .O(G1249) );

  xor2  gate883(.a(G1165), .b(G12), .O(gate441inter0));
  nand2 gate884(.a(gate441inter0), .b(s_48), .O(gate441inter1));
  and2  gate885(.a(G1165), .b(G12), .O(gate441inter2));
  inv1  gate886(.a(s_48), .O(gate441inter3));
  inv1  gate887(.a(s_49), .O(gate441inter4));
  nand2 gate888(.a(gate441inter4), .b(gate441inter3), .O(gate441inter5));
  nor2  gate889(.a(gate441inter5), .b(gate441inter2), .O(gate441inter6));
  inv1  gate890(.a(G12), .O(gate441inter7));
  inv1  gate891(.a(G1165), .O(gate441inter8));
  nand2 gate892(.a(gate441inter8), .b(gate441inter7), .O(gate441inter9));
  nand2 gate893(.a(s_49), .b(gate441inter3), .O(gate441inter10));
  nor2  gate894(.a(gate441inter10), .b(gate441inter9), .O(gate441inter11));
  nor2  gate895(.a(gate441inter11), .b(gate441inter6), .O(gate441inter12));
  nand2 gate896(.a(gate441inter12), .b(gate441inter1), .O(G1250));
nand2 gate442( .a(G1069), .b(G1165), .O(G1251) );
nand2 gate443( .a(G13), .b(G1168), .O(G1252) );

  xor2  gate939(.a(G1168), .b(G1072), .O(gate444inter0));
  nand2 gate940(.a(gate444inter0), .b(s_56), .O(gate444inter1));
  and2  gate941(.a(G1168), .b(G1072), .O(gate444inter2));
  inv1  gate942(.a(s_56), .O(gate444inter3));
  inv1  gate943(.a(s_57), .O(gate444inter4));
  nand2 gate944(.a(gate444inter4), .b(gate444inter3), .O(gate444inter5));
  nor2  gate945(.a(gate444inter5), .b(gate444inter2), .O(gate444inter6));
  inv1  gate946(.a(G1072), .O(gate444inter7));
  inv1  gate947(.a(G1168), .O(gate444inter8));
  nand2 gate948(.a(gate444inter8), .b(gate444inter7), .O(gate444inter9));
  nand2 gate949(.a(s_57), .b(gate444inter3), .O(gate444inter10));
  nor2  gate950(.a(gate444inter10), .b(gate444inter9), .O(gate444inter11));
  nor2  gate951(.a(gate444inter11), .b(gate444inter6), .O(gate444inter12));
  nand2 gate952(.a(gate444inter12), .b(gate444inter1), .O(G1253));
nand2 gate445( .a(G14), .b(G1171), .O(G1254) );
nand2 gate446( .a(G1075), .b(G1171), .O(G1255) );

  xor2  gate1177(.a(G1174), .b(G15), .O(gate447inter0));
  nand2 gate1178(.a(gate447inter0), .b(s_90), .O(gate447inter1));
  and2  gate1179(.a(G1174), .b(G15), .O(gate447inter2));
  inv1  gate1180(.a(s_90), .O(gate447inter3));
  inv1  gate1181(.a(s_91), .O(gate447inter4));
  nand2 gate1182(.a(gate447inter4), .b(gate447inter3), .O(gate447inter5));
  nor2  gate1183(.a(gate447inter5), .b(gate447inter2), .O(gate447inter6));
  inv1  gate1184(.a(G15), .O(gate447inter7));
  inv1  gate1185(.a(G1174), .O(gate447inter8));
  nand2 gate1186(.a(gate447inter8), .b(gate447inter7), .O(gate447inter9));
  nand2 gate1187(.a(s_91), .b(gate447inter3), .O(gate447inter10));
  nor2  gate1188(.a(gate447inter10), .b(gate447inter9), .O(gate447inter11));
  nor2  gate1189(.a(gate447inter11), .b(gate447inter6), .O(gate447inter12));
  nand2 gate1190(.a(gate447inter12), .b(gate447inter1), .O(G1256));
nand2 gate448( .a(G1078), .b(G1174), .O(G1257) );
nand2 gate449( .a(G16), .b(G1177), .O(G1258) );
nand2 gate450( .a(G1081), .b(G1177), .O(G1259) );
nand2 gate451( .a(G17), .b(G1180), .O(G1260) );
nand2 gate452( .a(G1084), .b(G1180), .O(G1261) );
nand2 gate453( .a(G18), .b(G1183), .O(G1262) );
nand2 gate454( .a(G1087), .b(G1183), .O(G1263) );
nand2 gate455( .a(G19), .b(G1186), .O(G1264) );

  xor2  gate995(.a(G1186), .b(G1090), .O(gate456inter0));
  nand2 gate996(.a(gate456inter0), .b(s_64), .O(gate456inter1));
  and2  gate997(.a(G1186), .b(G1090), .O(gate456inter2));
  inv1  gate998(.a(s_64), .O(gate456inter3));
  inv1  gate999(.a(s_65), .O(gate456inter4));
  nand2 gate1000(.a(gate456inter4), .b(gate456inter3), .O(gate456inter5));
  nor2  gate1001(.a(gate456inter5), .b(gate456inter2), .O(gate456inter6));
  inv1  gate1002(.a(G1090), .O(gate456inter7));
  inv1  gate1003(.a(G1186), .O(gate456inter8));
  nand2 gate1004(.a(gate456inter8), .b(gate456inter7), .O(gate456inter9));
  nand2 gate1005(.a(s_65), .b(gate456inter3), .O(gate456inter10));
  nor2  gate1006(.a(gate456inter10), .b(gate456inter9), .O(gate456inter11));
  nor2  gate1007(.a(gate456inter11), .b(gate456inter6), .O(gate456inter12));
  nand2 gate1008(.a(gate456inter12), .b(gate456inter1), .O(G1265));
nand2 gate457( .a(G20), .b(G1189), .O(G1266) );
nand2 gate458( .a(G1093), .b(G1189), .O(G1267) );
nand2 gate459( .a(G21), .b(G1192), .O(G1268) );
nand2 gate460( .a(G1096), .b(G1192), .O(G1269) );

  xor2  gate589(.a(G1195), .b(G22), .O(gate461inter0));
  nand2 gate590(.a(gate461inter0), .b(s_6), .O(gate461inter1));
  and2  gate591(.a(G1195), .b(G22), .O(gate461inter2));
  inv1  gate592(.a(s_6), .O(gate461inter3));
  inv1  gate593(.a(s_7), .O(gate461inter4));
  nand2 gate594(.a(gate461inter4), .b(gate461inter3), .O(gate461inter5));
  nor2  gate595(.a(gate461inter5), .b(gate461inter2), .O(gate461inter6));
  inv1  gate596(.a(G22), .O(gate461inter7));
  inv1  gate597(.a(G1195), .O(gate461inter8));
  nand2 gate598(.a(gate461inter8), .b(gate461inter7), .O(gate461inter9));
  nand2 gate599(.a(s_7), .b(gate461inter3), .O(gate461inter10));
  nor2  gate600(.a(gate461inter10), .b(gate461inter9), .O(gate461inter11));
  nor2  gate601(.a(gate461inter11), .b(gate461inter6), .O(gate461inter12));
  nand2 gate602(.a(gate461inter12), .b(gate461inter1), .O(G1270));
nand2 gate462( .a(G1099), .b(G1195), .O(G1271) );
nand2 gate463( .a(G23), .b(G1198), .O(G1272) );
nand2 gate464( .a(G1102), .b(G1198), .O(G1273) );
nand2 gate465( .a(G24), .b(G1201), .O(G1274) );
nand2 gate466( .a(G1105), .b(G1201), .O(G1275) );
nand2 gate467( .a(G25), .b(G1204), .O(G1276) );
nand2 gate468( .a(G1108), .b(G1204), .O(G1277) );
nand2 gate469( .a(G26), .b(G1207), .O(G1278) );
nand2 gate470( .a(G1111), .b(G1207), .O(G1279) );
nand2 gate471( .a(G27), .b(G1210), .O(G1280) );
nand2 gate472( .a(G1114), .b(G1210), .O(G1281) );

  xor2  gate1149(.a(G1213), .b(G28), .O(gate473inter0));
  nand2 gate1150(.a(gate473inter0), .b(s_86), .O(gate473inter1));
  and2  gate1151(.a(G1213), .b(G28), .O(gate473inter2));
  inv1  gate1152(.a(s_86), .O(gate473inter3));
  inv1  gate1153(.a(s_87), .O(gate473inter4));
  nand2 gate1154(.a(gate473inter4), .b(gate473inter3), .O(gate473inter5));
  nor2  gate1155(.a(gate473inter5), .b(gate473inter2), .O(gate473inter6));
  inv1  gate1156(.a(G28), .O(gate473inter7));
  inv1  gate1157(.a(G1213), .O(gate473inter8));
  nand2 gate1158(.a(gate473inter8), .b(gate473inter7), .O(gate473inter9));
  nand2 gate1159(.a(s_87), .b(gate473inter3), .O(gate473inter10));
  nor2  gate1160(.a(gate473inter10), .b(gate473inter9), .O(gate473inter11));
  nor2  gate1161(.a(gate473inter11), .b(gate473inter6), .O(gate473inter12));
  nand2 gate1162(.a(gate473inter12), .b(gate473inter1), .O(G1282));
nand2 gate474( .a(G1117), .b(G1213), .O(G1283) );
nand2 gate475( .a(G29), .b(G1216), .O(G1284) );
nand2 gate476( .a(G1120), .b(G1216), .O(G1285) );
nand2 gate477( .a(G30), .b(G1219), .O(G1286) );
nand2 gate478( .a(G1123), .b(G1219), .O(G1287) );
nand2 gate479( .a(G31), .b(G1222), .O(G1288) );
nand2 gate480( .a(G1126), .b(G1222), .O(G1289) );
nand2 gate481( .a(G32), .b(G1225), .O(G1290) );
nand2 gate482( .a(G1129), .b(G1225), .O(G1291) );
nand2 gate483( .a(G1228), .b(G1229), .O(G1292) );
nand2 gate484( .a(G1230), .b(G1231), .O(G1293) );
nand2 gate485( .a(G1232), .b(G1233), .O(G1294) );
nand2 gate486( .a(G1234), .b(G1235), .O(G1295) );
nand2 gate487( .a(G1236), .b(G1237), .O(G1296) );
nand2 gate488( .a(G1238), .b(G1239), .O(G1297) );

  xor2  gate1485(.a(G1241), .b(G1240), .O(gate489inter0));
  nand2 gate1486(.a(gate489inter0), .b(s_134), .O(gate489inter1));
  and2  gate1487(.a(G1241), .b(G1240), .O(gate489inter2));
  inv1  gate1488(.a(s_134), .O(gate489inter3));
  inv1  gate1489(.a(s_135), .O(gate489inter4));
  nand2 gate1490(.a(gate489inter4), .b(gate489inter3), .O(gate489inter5));
  nor2  gate1491(.a(gate489inter5), .b(gate489inter2), .O(gate489inter6));
  inv1  gate1492(.a(G1240), .O(gate489inter7));
  inv1  gate1493(.a(G1241), .O(gate489inter8));
  nand2 gate1494(.a(gate489inter8), .b(gate489inter7), .O(gate489inter9));
  nand2 gate1495(.a(s_135), .b(gate489inter3), .O(gate489inter10));
  nor2  gate1496(.a(gate489inter10), .b(gate489inter9), .O(gate489inter11));
  nor2  gate1497(.a(gate489inter11), .b(gate489inter6), .O(gate489inter12));
  nand2 gate1498(.a(gate489inter12), .b(gate489inter1), .O(G1298));
nand2 gate490( .a(G1242), .b(G1243), .O(G1299) );
nand2 gate491( .a(G1244), .b(G1245), .O(G1300) );
nand2 gate492( .a(G1246), .b(G1247), .O(G1301) );

  xor2  gate1191(.a(G1249), .b(G1248), .O(gate493inter0));
  nand2 gate1192(.a(gate493inter0), .b(s_92), .O(gate493inter1));
  and2  gate1193(.a(G1249), .b(G1248), .O(gate493inter2));
  inv1  gate1194(.a(s_92), .O(gate493inter3));
  inv1  gate1195(.a(s_93), .O(gate493inter4));
  nand2 gate1196(.a(gate493inter4), .b(gate493inter3), .O(gate493inter5));
  nor2  gate1197(.a(gate493inter5), .b(gate493inter2), .O(gate493inter6));
  inv1  gate1198(.a(G1248), .O(gate493inter7));
  inv1  gate1199(.a(G1249), .O(gate493inter8));
  nand2 gate1200(.a(gate493inter8), .b(gate493inter7), .O(gate493inter9));
  nand2 gate1201(.a(s_93), .b(gate493inter3), .O(gate493inter10));
  nor2  gate1202(.a(gate493inter10), .b(gate493inter9), .O(gate493inter11));
  nor2  gate1203(.a(gate493inter11), .b(gate493inter6), .O(gate493inter12));
  nand2 gate1204(.a(gate493inter12), .b(gate493inter1), .O(G1302));
nand2 gate494( .a(G1250), .b(G1251), .O(G1303) );
nand2 gate495( .a(G1252), .b(G1253), .O(G1304) );
nand2 gate496( .a(G1254), .b(G1255), .O(G1305) );

  xor2  gate925(.a(G1257), .b(G1256), .O(gate497inter0));
  nand2 gate926(.a(gate497inter0), .b(s_54), .O(gate497inter1));
  and2  gate927(.a(G1257), .b(G1256), .O(gate497inter2));
  inv1  gate928(.a(s_54), .O(gate497inter3));
  inv1  gate929(.a(s_55), .O(gate497inter4));
  nand2 gate930(.a(gate497inter4), .b(gate497inter3), .O(gate497inter5));
  nor2  gate931(.a(gate497inter5), .b(gate497inter2), .O(gate497inter6));
  inv1  gate932(.a(G1256), .O(gate497inter7));
  inv1  gate933(.a(G1257), .O(gate497inter8));
  nand2 gate934(.a(gate497inter8), .b(gate497inter7), .O(gate497inter9));
  nand2 gate935(.a(s_55), .b(gate497inter3), .O(gate497inter10));
  nor2  gate936(.a(gate497inter10), .b(gate497inter9), .O(gate497inter11));
  nor2  gate937(.a(gate497inter11), .b(gate497inter6), .O(gate497inter12));
  nand2 gate938(.a(gate497inter12), .b(gate497inter1), .O(G1306));
nand2 gate498( .a(G1258), .b(G1259), .O(G1307) );
nand2 gate499( .a(G1260), .b(G1261), .O(G1308) );
nand2 gate500( .a(G1262), .b(G1263), .O(G1309) );
nand2 gate501( .a(G1264), .b(G1265), .O(G1310) );
nand2 gate502( .a(G1266), .b(G1267), .O(G1311) );
nand2 gate503( .a(G1268), .b(G1269), .O(G1312) );
nand2 gate504( .a(G1270), .b(G1271), .O(G1313) );
nand2 gate505( .a(G1272), .b(G1273), .O(G1314) );
nand2 gate506( .a(G1274), .b(G1275), .O(G1315) );
nand2 gate507( .a(G1276), .b(G1277), .O(G1316) );
nand2 gate508( .a(G1278), .b(G1279), .O(G1317) );
nand2 gate509( .a(G1280), .b(G1281), .O(G1318) );
nand2 gate510( .a(G1282), .b(G1283), .O(G1319) );
nand2 gate511( .a(G1284), .b(G1285), .O(G1320) );
nand2 gate512( .a(G1286), .b(G1287), .O(G1321) );

  xor2  gate1499(.a(G1289), .b(G1288), .O(gate513inter0));
  nand2 gate1500(.a(gate513inter0), .b(s_136), .O(gate513inter1));
  and2  gate1501(.a(G1289), .b(G1288), .O(gate513inter2));
  inv1  gate1502(.a(s_136), .O(gate513inter3));
  inv1  gate1503(.a(s_137), .O(gate513inter4));
  nand2 gate1504(.a(gate513inter4), .b(gate513inter3), .O(gate513inter5));
  nor2  gate1505(.a(gate513inter5), .b(gate513inter2), .O(gate513inter6));
  inv1  gate1506(.a(G1288), .O(gate513inter7));
  inv1  gate1507(.a(G1289), .O(gate513inter8));
  nand2 gate1508(.a(gate513inter8), .b(gate513inter7), .O(gate513inter9));
  nand2 gate1509(.a(s_137), .b(gate513inter3), .O(gate513inter10));
  nor2  gate1510(.a(gate513inter10), .b(gate513inter9), .O(gate513inter11));
  nor2  gate1511(.a(gate513inter11), .b(gate513inter6), .O(gate513inter12));
  nand2 gate1512(.a(gate513inter12), .b(gate513inter1), .O(G1322));
nand2 gate514( .a(G1290), .b(G1291), .O(G1323) );
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule