module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);

input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;//RE__PI;

input s_0,s_1;//RE__ALLOW(00,01,10,11);
input s_2,s_3;//RE__ALLOW(00,01,10,11);
input s_4,s_5;//RE__ALLOW(00,01,10,11);
input s_6,s_7;//RE__ALLOW(00,01,10,11);
input s_8,s_9;//RE__ALLOW(00,01,10,11);
input s_10,s_11;//RE__ALLOW(00,01,10,11);
input s_12,s_13;//RE__ALLOW(00,01,10,11);
input s_14,s_15;//RE__ALLOW(00,01,10,11);
input s_16,s_17;//RE__ALLOW(00,01,10,11);
input s_18,s_19;//RE__ALLOW(00,01,10,11);
input s_20,s_21;//RE__ALLOW(00,01,10,11);
input s_22,s_23;//RE__ALLOW(00,01,10,11);
input s_24,s_25;//RE__ALLOW(00,01,10,11);
input s_26,s_27;//RE__ALLOW(00,01,10,11);
input s_28,s_29;//RE__ALLOW(00,01,10,11);
input s_30,s_31;//RE__ALLOW(00,01,10,11);
input s_32,s_33;//RE__ALLOW(00,01,10,11);
input s_34,s_35;//RE__ALLOW(00,01,10,11);
input s_36,s_37;//RE__ALLOW(00,01,10,11);
input s_38,s_39;//RE__ALLOW(00,01,10,11);
input s_40,s_41;//RE__ALLOW(00,01,10,11);
input s_42,s_43;//RE__ALLOW(00,01,10,11);
input s_44,s_45;//RE__ALLOW(00,01,10,11);
input s_46,s_47;//RE__ALLOW(00,01,10,11);
input s_48,s_49;//RE__ALLOW(00,01,10,11);
input s_50,s_51;//RE__ALLOW(00,01,10,11);
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;

  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate183inter0, gate183inter1, gate183inter2, gate183inter3, gate183inter4, gate183inter5, gate183inter6, gate183inter7, gate183inter8, gate183inter9, gate183inter10, gate183inter11, gate183inter12, gate20inter0, gate20inter1, gate20inter2, gate20inter3, gate20inter4, gate20inter5, gate20inter6, gate20inter7, gate20inter8, gate20inter9, gate20inter10, gate20inter11, gate20inter12, gate395inter0, gate395inter1, gate395inter2, gate395inter3, gate395inter4, gate395inter5, gate395inter6, gate395inter7, gate395inter8, gate395inter9, gate395inter10, gate395inter11, gate395inter12, gate54inter0, gate54inter1, gate54inter2, gate54inter3, gate54inter4, gate54inter5, gate54inter6, gate54inter7, gate54inter8, gate54inter9, gate54inter10, gate54inter11, gate54inter12, gate117inter0, gate117inter1, gate117inter2, gate117inter3, gate117inter4, gate117inter5, gate117inter6, gate117inter7, gate117inter8, gate117inter9, gate117inter10, gate117inter11, gate117inter12, gate24inter0, gate24inter1, gate24inter2, gate24inter3, gate24inter4, gate24inter5, gate24inter6, gate24inter7, gate24inter8, gate24inter9, gate24inter10, gate24inter11, gate24inter12, gate115inter0, gate115inter1, gate115inter2, gate115inter3, gate115inter4, gate115inter5, gate115inter6, gate115inter7, gate115inter8, gate115inter9, gate115inter10, gate115inter11, gate115inter12, gate11inter0, gate11inter1, gate11inter2, gate11inter3, gate11inter4, gate11inter5, gate11inter6, gate11inter7, gate11inter8, gate11inter9, gate11inter10, gate11inter11, gate11inter12, gate285inter0, gate285inter1, gate285inter2, gate285inter3, gate285inter4, gate285inter5, gate285inter6, gate285inter7, gate285inter8, gate285inter9, gate285inter10, gate285inter11, gate285inter12, gate241inter0, gate241inter1, gate241inter2, gate241inter3, gate241inter4, gate241inter5, gate241inter6, gate241inter7, gate241inter8, gate241inter9, gate241inter10, gate241inter11, gate241inter12, gate279inter0, gate279inter1, gate279inter2, gate279inter3, gate279inter4, gate279inter5, gate279inter6, gate279inter7, gate279inter8, gate279inter9, gate279inter10, gate279inter11, gate279inter12, gate289inter0, gate289inter1, gate289inter2, gate289inter3, gate289inter4, gate289inter5, gate289inter6, gate289inter7, gate289inter8, gate289inter9, gate289inter10, gate289inter11, gate289inter12, gate52inter0, gate52inter1, gate52inter2, gate52inter3, gate52inter4, gate52inter5, gate52inter6, gate52inter7, gate52inter8, gate52inter9, gate52inter10, gate52inter11, gate52inter12, gate472inter0, gate472inter1, gate472inter2, gate472inter3, gate472inter4, gate472inter5, gate472inter6, gate472inter7, gate472inter8, gate472inter9, gate472inter10, gate472inter11, gate472inter12, gate406inter0, gate406inter1, gate406inter2, gate406inter3, gate406inter4, gate406inter5, gate406inter6, gate406inter7, gate406inter8, gate406inter9, gate406inter10, gate406inter11, gate406inter12, gate265inter0, gate265inter1, gate265inter2, gate265inter3, gate265inter4, gate265inter5, gate265inter6, gate265inter7, gate265inter8, gate265inter9, gate265inter10, gate265inter11, gate265inter12, gate15inter0, gate15inter1, gate15inter2, gate15inter3, gate15inter4, gate15inter5, gate15inter6, gate15inter7, gate15inter8, gate15inter9, gate15inter10, gate15inter11, gate15inter12, gate26inter0, gate26inter1, gate26inter2, gate26inter3, gate26inter4, gate26inter5, gate26inter6, gate26inter7, gate26inter8, gate26inter9, gate26inter10, gate26inter11, gate26inter12, gate156inter0, gate156inter1, gate156inter2, gate156inter3, gate156inter4, gate156inter5, gate156inter6, gate156inter7, gate156inter8, gate156inter9, gate156inter10, gate156inter11, gate156inter12, gate48inter0, gate48inter1, gate48inter2, gate48inter3, gate48inter4, gate48inter5, gate48inter6, gate48inter7, gate48inter8, gate48inter9, gate48inter10, gate48inter11, gate48inter12, gate211inter0, gate211inter1, gate211inter2, gate211inter3, gate211inter4, gate211inter5, gate211inter6, gate211inter7, gate211inter8, gate211inter9, gate211inter10, gate211inter11, gate211inter12, gate9inter0, gate9inter1, gate9inter2, gate9inter3, gate9inter4, gate9inter5, gate9inter6, gate9inter7, gate9inter8, gate9inter9, gate9inter10, gate9inter11, gate9inter12, gate149inter0, gate149inter1, gate149inter2, gate149inter3, gate149inter4, gate149inter5, gate149inter6, gate149inter7, gate149inter8, gate149inter9, gate149inter10, gate149inter11, gate149inter12, gate436inter0, gate436inter1, gate436inter2, gate436inter3, gate436inter4, gate436inter5, gate436inter6, gate436inter7, gate436inter8, gate436inter9, gate436inter10, gate436inter11, gate436inter12, gate269inter0, gate269inter1, gate269inter2, gate269inter3, gate269inter4, gate269inter5, gate269inter6, gate269inter7, gate269inter8, gate269inter9, gate269inter10, gate269inter11, gate269inter12, gate195inter0, gate195inter1, gate195inter2, gate195inter3, gate195inter4, gate195inter5, gate195inter6, gate195inter7, gate195inter8, gate195inter9, gate195inter10, gate195inter11, gate195inter12;



and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );

  xor2  gate841(.a(G2), .b(G1), .O(gate9inter0));
  nand2 gate842(.a(gate9inter0), .b(s_42), .O(gate9inter1));
  and2  gate843(.a(G2), .b(G1), .O(gate9inter2));
  inv1  gate844(.a(s_42), .O(gate9inter3));
  inv1  gate845(.a(s_43), .O(gate9inter4));
  nand2 gate846(.a(gate9inter4), .b(gate9inter3), .O(gate9inter5));
  nor2  gate847(.a(gate9inter5), .b(gate9inter2), .O(gate9inter6));
  inv1  gate848(.a(G1), .O(gate9inter7));
  inv1  gate849(.a(G2), .O(gate9inter8));
  nand2 gate850(.a(gate9inter8), .b(gate9inter7), .O(gate9inter9));
  nand2 gate851(.a(s_43), .b(gate9inter3), .O(gate9inter10));
  nor2  gate852(.a(gate9inter10), .b(gate9inter9), .O(gate9inter11));
  nor2  gate853(.a(gate9inter11), .b(gate9inter6), .O(gate9inter12));
  nand2 gate854(.a(gate9inter12), .b(gate9inter1), .O(G266));
nand2 gate10( .a(G3), .b(G4), .O(G269) );

  xor2  gate645(.a(G6), .b(G5), .O(gate11inter0));
  nand2 gate646(.a(gate11inter0), .b(s_14), .O(gate11inter1));
  and2  gate647(.a(G6), .b(G5), .O(gate11inter2));
  inv1  gate648(.a(s_14), .O(gate11inter3));
  inv1  gate649(.a(s_15), .O(gate11inter4));
  nand2 gate650(.a(gate11inter4), .b(gate11inter3), .O(gate11inter5));
  nor2  gate651(.a(gate11inter5), .b(gate11inter2), .O(gate11inter6));
  inv1  gate652(.a(G5), .O(gate11inter7));
  inv1  gate653(.a(G6), .O(gate11inter8));
  nand2 gate654(.a(gate11inter8), .b(gate11inter7), .O(gate11inter9));
  nand2 gate655(.a(s_15), .b(gate11inter3), .O(gate11inter10));
  nor2  gate656(.a(gate11inter10), .b(gate11inter9), .O(gate11inter11));
  nor2  gate657(.a(gate11inter11), .b(gate11inter6), .O(gate11inter12));
  nand2 gate658(.a(gate11inter12), .b(gate11inter1), .O(G272));
nand2 gate12( .a(G7), .b(G8), .O(G275) );
nand2 gate13( .a(G9), .b(G10), .O(G278) );
nand2 gate14( .a(G11), .b(G12), .O(G281) );

  xor2  gate771(.a(G14), .b(G13), .O(gate15inter0));
  nand2 gate772(.a(gate15inter0), .b(s_32), .O(gate15inter1));
  and2  gate773(.a(G14), .b(G13), .O(gate15inter2));
  inv1  gate774(.a(s_32), .O(gate15inter3));
  inv1  gate775(.a(s_33), .O(gate15inter4));
  nand2 gate776(.a(gate15inter4), .b(gate15inter3), .O(gate15inter5));
  nor2  gate777(.a(gate15inter5), .b(gate15inter2), .O(gate15inter6));
  inv1  gate778(.a(G13), .O(gate15inter7));
  inv1  gate779(.a(G14), .O(gate15inter8));
  nand2 gate780(.a(gate15inter8), .b(gate15inter7), .O(gate15inter9));
  nand2 gate781(.a(s_33), .b(gate15inter3), .O(gate15inter10));
  nor2  gate782(.a(gate15inter10), .b(gate15inter9), .O(gate15inter11));
  nor2  gate783(.a(gate15inter11), .b(gate15inter6), .O(gate15inter12));
  nand2 gate784(.a(gate15inter12), .b(gate15inter1), .O(G284));
nand2 gate16( .a(G15), .b(G16), .O(G287) );
nand2 gate17( .a(G17), .b(G18), .O(G290) );
nand2 gate18( .a(G19), .b(G20), .O(G293) );
nand2 gate19( .a(G21), .b(G22), .O(G296) );

  xor2  gate561(.a(G24), .b(G23), .O(gate20inter0));
  nand2 gate562(.a(gate20inter0), .b(s_2), .O(gate20inter1));
  and2  gate563(.a(G24), .b(G23), .O(gate20inter2));
  inv1  gate564(.a(s_2), .O(gate20inter3));
  inv1  gate565(.a(s_3), .O(gate20inter4));
  nand2 gate566(.a(gate20inter4), .b(gate20inter3), .O(gate20inter5));
  nor2  gate567(.a(gate20inter5), .b(gate20inter2), .O(gate20inter6));
  inv1  gate568(.a(G23), .O(gate20inter7));
  inv1  gate569(.a(G24), .O(gate20inter8));
  nand2 gate570(.a(gate20inter8), .b(gate20inter7), .O(gate20inter9));
  nand2 gate571(.a(s_3), .b(gate20inter3), .O(gate20inter10));
  nor2  gate572(.a(gate20inter10), .b(gate20inter9), .O(gate20inter11));
  nor2  gate573(.a(gate20inter11), .b(gate20inter6), .O(gate20inter12));
  nand2 gate574(.a(gate20inter12), .b(gate20inter1), .O(G299));
nand2 gate21( .a(G25), .b(G26), .O(G302) );
nand2 gate22( .a(G27), .b(G28), .O(G305) );
nand2 gate23( .a(G29), .b(G30), .O(G308) );

  xor2  gate617(.a(G32), .b(G31), .O(gate24inter0));
  nand2 gate618(.a(gate24inter0), .b(s_10), .O(gate24inter1));
  and2  gate619(.a(G32), .b(G31), .O(gate24inter2));
  inv1  gate620(.a(s_10), .O(gate24inter3));
  inv1  gate621(.a(s_11), .O(gate24inter4));
  nand2 gate622(.a(gate24inter4), .b(gate24inter3), .O(gate24inter5));
  nor2  gate623(.a(gate24inter5), .b(gate24inter2), .O(gate24inter6));
  inv1  gate624(.a(G31), .O(gate24inter7));
  inv1  gate625(.a(G32), .O(gate24inter8));
  nand2 gate626(.a(gate24inter8), .b(gate24inter7), .O(gate24inter9));
  nand2 gate627(.a(s_11), .b(gate24inter3), .O(gate24inter10));
  nor2  gate628(.a(gate24inter10), .b(gate24inter9), .O(gate24inter11));
  nor2  gate629(.a(gate24inter11), .b(gate24inter6), .O(gate24inter12));
  nand2 gate630(.a(gate24inter12), .b(gate24inter1), .O(G311));
nand2 gate25( .a(G1), .b(G5), .O(G314) );

  xor2  gate785(.a(G13), .b(G9), .O(gate26inter0));
  nand2 gate786(.a(gate26inter0), .b(s_34), .O(gate26inter1));
  and2  gate787(.a(G13), .b(G9), .O(gate26inter2));
  inv1  gate788(.a(s_34), .O(gate26inter3));
  inv1  gate789(.a(s_35), .O(gate26inter4));
  nand2 gate790(.a(gate26inter4), .b(gate26inter3), .O(gate26inter5));
  nor2  gate791(.a(gate26inter5), .b(gate26inter2), .O(gate26inter6));
  inv1  gate792(.a(G9), .O(gate26inter7));
  inv1  gate793(.a(G13), .O(gate26inter8));
  nand2 gate794(.a(gate26inter8), .b(gate26inter7), .O(gate26inter9));
  nand2 gate795(.a(s_35), .b(gate26inter3), .O(gate26inter10));
  nor2  gate796(.a(gate26inter10), .b(gate26inter9), .O(gate26inter11));
  nor2  gate797(.a(gate26inter11), .b(gate26inter6), .O(gate26inter12));
  nand2 gate798(.a(gate26inter12), .b(gate26inter1), .O(G317));
nand2 gate27( .a(G2), .b(G6), .O(G320) );
nand2 gate28( .a(G10), .b(G14), .O(G323) );
nand2 gate29( .a(G3), .b(G7), .O(G326) );
nand2 gate30( .a(G11), .b(G15), .O(G329) );
nand2 gate31( .a(G4), .b(G8), .O(G332) );
nand2 gate32( .a(G12), .b(G16), .O(G335) );
nand2 gate33( .a(G17), .b(G21), .O(G338) );
nand2 gate34( .a(G25), .b(G29), .O(G341) );
nand2 gate35( .a(G18), .b(G22), .O(G344) );
nand2 gate36( .a(G26), .b(G30), .O(G347) );
nand2 gate37( .a(G19), .b(G23), .O(G350) );
nand2 gate38( .a(G27), .b(G31), .O(G353) );
nand2 gate39( .a(G20), .b(G24), .O(G356) );
nand2 gate40( .a(G28), .b(G32), .O(G359) );
nand2 gate41( .a(G1), .b(G266), .O(G362) );
nand2 gate42( .a(G2), .b(G266), .O(G363) );
nand2 gate43( .a(G3), .b(G269), .O(G364) );
nand2 gate44( .a(G4), .b(G269), .O(G365) );
nand2 gate45( .a(G5), .b(G272), .O(G366) );
nand2 gate46( .a(G6), .b(G272), .O(G367) );
nand2 gate47( .a(G7), .b(G275), .O(G368) );

  xor2  gate813(.a(G275), .b(G8), .O(gate48inter0));
  nand2 gate814(.a(gate48inter0), .b(s_38), .O(gate48inter1));
  and2  gate815(.a(G275), .b(G8), .O(gate48inter2));
  inv1  gate816(.a(s_38), .O(gate48inter3));
  inv1  gate817(.a(s_39), .O(gate48inter4));
  nand2 gate818(.a(gate48inter4), .b(gate48inter3), .O(gate48inter5));
  nor2  gate819(.a(gate48inter5), .b(gate48inter2), .O(gate48inter6));
  inv1  gate820(.a(G8), .O(gate48inter7));
  inv1  gate821(.a(G275), .O(gate48inter8));
  nand2 gate822(.a(gate48inter8), .b(gate48inter7), .O(gate48inter9));
  nand2 gate823(.a(s_39), .b(gate48inter3), .O(gate48inter10));
  nor2  gate824(.a(gate48inter10), .b(gate48inter9), .O(gate48inter11));
  nor2  gate825(.a(gate48inter11), .b(gate48inter6), .O(gate48inter12));
  nand2 gate826(.a(gate48inter12), .b(gate48inter1), .O(G369));
nand2 gate49( .a(G9), .b(G278), .O(G370) );
nand2 gate50( .a(G10), .b(G278), .O(G371) );
nand2 gate51( .a(G11), .b(G281), .O(G372) );

  xor2  gate715(.a(G281), .b(G12), .O(gate52inter0));
  nand2 gate716(.a(gate52inter0), .b(s_24), .O(gate52inter1));
  and2  gate717(.a(G281), .b(G12), .O(gate52inter2));
  inv1  gate718(.a(s_24), .O(gate52inter3));
  inv1  gate719(.a(s_25), .O(gate52inter4));
  nand2 gate720(.a(gate52inter4), .b(gate52inter3), .O(gate52inter5));
  nor2  gate721(.a(gate52inter5), .b(gate52inter2), .O(gate52inter6));
  inv1  gate722(.a(G12), .O(gate52inter7));
  inv1  gate723(.a(G281), .O(gate52inter8));
  nand2 gate724(.a(gate52inter8), .b(gate52inter7), .O(gate52inter9));
  nand2 gate725(.a(s_25), .b(gate52inter3), .O(gate52inter10));
  nor2  gate726(.a(gate52inter10), .b(gate52inter9), .O(gate52inter11));
  nor2  gate727(.a(gate52inter11), .b(gate52inter6), .O(gate52inter12));
  nand2 gate728(.a(gate52inter12), .b(gate52inter1), .O(G373));
nand2 gate53( .a(G13), .b(G284), .O(G374) );

  xor2  gate589(.a(G284), .b(G14), .O(gate54inter0));
  nand2 gate590(.a(gate54inter0), .b(s_6), .O(gate54inter1));
  and2  gate591(.a(G284), .b(G14), .O(gate54inter2));
  inv1  gate592(.a(s_6), .O(gate54inter3));
  inv1  gate593(.a(s_7), .O(gate54inter4));
  nand2 gate594(.a(gate54inter4), .b(gate54inter3), .O(gate54inter5));
  nor2  gate595(.a(gate54inter5), .b(gate54inter2), .O(gate54inter6));
  inv1  gate596(.a(G14), .O(gate54inter7));
  inv1  gate597(.a(G284), .O(gate54inter8));
  nand2 gate598(.a(gate54inter8), .b(gate54inter7), .O(gate54inter9));
  nand2 gate599(.a(s_7), .b(gate54inter3), .O(gate54inter10));
  nor2  gate600(.a(gate54inter10), .b(gate54inter9), .O(gate54inter11));
  nor2  gate601(.a(gate54inter11), .b(gate54inter6), .O(gate54inter12));
  nand2 gate602(.a(gate54inter12), .b(gate54inter1), .O(G375));
nand2 gate55( .a(G15), .b(G287), .O(G376) );
nand2 gate56( .a(G16), .b(G287), .O(G377) );
nand2 gate57( .a(G17), .b(G290), .O(G378) );
nand2 gate58( .a(G18), .b(G290), .O(G379) );
nand2 gate59( .a(G19), .b(G293), .O(G380) );
nand2 gate60( .a(G20), .b(G293), .O(G381) );
nand2 gate61( .a(G21), .b(G296), .O(G382) );
nand2 gate62( .a(G22), .b(G296), .O(G383) );
nand2 gate63( .a(G23), .b(G299), .O(G384) );
nand2 gate64( .a(G24), .b(G299), .O(G385) );
nand2 gate65( .a(G25), .b(G302), .O(G386) );
nand2 gate66( .a(G26), .b(G302), .O(G387) );
nand2 gate67( .a(G27), .b(G305), .O(G388) );
nand2 gate68( .a(G28), .b(G305), .O(G389) );
nand2 gate69( .a(G29), .b(G308), .O(G390) );
nand2 gate70( .a(G30), .b(G308), .O(G391) );
nand2 gate71( .a(G31), .b(G311), .O(G392) );
nand2 gate72( .a(G32), .b(G311), .O(G393) );
nand2 gate73( .a(G1), .b(G314), .O(G394) );
nand2 gate74( .a(G5), .b(G314), .O(G395) );
nand2 gate75( .a(G9), .b(G317), .O(G396) );
nand2 gate76( .a(G13), .b(G317), .O(G397) );
nand2 gate77( .a(G2), .b(G320), .O(G398) );
nand2 gate78( .a(G6), .b(G320), .O(G399) );
nand2 gate79( .a(G10), .b(G323), .O(G400) );
nand2 gate80( .a(G14), .b(G323), .O(G401) );
nand2 gate81( .a(G3), .b(G326), .O(G402) );
nand2 gate82( .a(G7), .b(G326), .O(G403) );
nand2 gate83( .a(G11), .b(G329), .O(G404) );
nand2 gate84( .a(G15), .b(G329), .O(G405) );
nand2 gate85( .a(G4), .b(G332), .O(G406) );
nand2 gate86( .a(G8), .b(G332), .O(G407) );
nand2 gate87( .a(G12), .b(G335), .O(G408) );
nand2 gate88( .a(G16), .b(G335), .O(G409) );
nand2 gate89( .a(G17), .b(G338), .O(G410) );
nand2 gate90( .a(G21), .b(G338), .O(G411) );
nand2 gate91( .a(G25), .b(G341), .O(G412) );
nand2 gate92( .a(G29), .b(G341), .O(G413) );
nand2 gate93( .a(G18), .b(G344), .O(G414) );
nand2 gate94( .a(G22), .b(G344), .O(G415) );
nand2 gate95( .a(G26), .b(G347), .O(G416) );
nand2 gate96( .a(G30), .b(G347), .O(G417) );
nand2 gate97( .a(G19), .b(G350), .O(G418) );
nand2 gate98( .a(G23), .b(G350), .O(G419) );
nand2 gate99( .a(G27), .b(G353), .O(G420) );
nand2 gate100( .a(G31), .b(G353), .O(G421) );
nand2 gate101( .a(G20), .b(G356), .O(G422) );
nand2 gate102( .a(G24), .b(G356), .O(G423) );
nand2 gate103( .a(G28), .b(G359), .O(G424) );
nand2 gate104( .a(G32), .b(G359), .O(G425) );
nand2 gate105( .a(G362), .b(G363), .O(G426) );
nand2 gate106( .a(G364), .b(G365), .O(G429) );
nand2 gate107( .a(G366), .b(G367), .O(G432) );
nand2 gate108( .a(G368), .b(G369), .O(G435) );
nand2 gate109( .a(G370), .b(G371), .O(G438) );
nand2 gate110( .a(G372), .b(G373), .O(G441) );
nand2 gate111( .a(G374), .b(G375), .O(G444) );
nand2 gate112( .a(G376), .b(G377), .O(G447) );
nand2 gate113( .a(G378), .b(G379), .O(G450) );
nand2 gate114( .a(G380), .b(G381), .O(G453) );

  xor2  gate631(.a(G383), .b(G382), .O(gate115inter0));
  nand2 gate632(.a(gate115inter0), .b(s_12), .O(gate115inter1));
  and2  gate633(.a(G383), .b(G382), .O(gate115inter2));
  inv1  gate634(.a(s_12), .O(gate115inter3));
  inv1  gate635(.a(s_13), .O(gate115inter4));
  nand2 gate636(.a(gate115inter4), .b(gate115inter3), .O(gate115inter5));
  nor2  gate637(.a(gate115inter5), .b(gate115inter2), .O(gate115inter6));
  inv1  gate638(.a(G382), .O(gate115inter7));
  inv1  gate639(.a(G383), .O(gate115inter8));
  nand2 gate640(.a(gate115inter8), .b(gate115inter7), .O(gate115inter9));
  nand2 gate641(.a(s_13), .b(gate115inter3), .O(gate115inter10));
  nor2  gate642(.a(gate115inter10), .b(gate115inter9), .O(gate115inter11));
  nor2  gate643(.a(gate115inter11), .b(gate115inter6), .O(gate115inter12));
  nand2 gate644(.a(gate115inter12), .b(gate115inter1), .O(G456));
nand2 gate116( .a(G384), .b(G385), .O(G459) );

  xor2  gate603(.a(G387), .b(G386), .O(gate117inter0));
  nand2 gate604(.a(gate117inter0), .b(s_8), .O(gate117inter1));
  and2  gate605(.a(G387), .b(G386), .O(gate117inter2));
  inv1  gate606(.a(s_8), .O(gate117inter3));
  inv1  gate607(.a(s_9), .O(gate117inter4));
  nand2 gate608(.a(gate117inter4), .b(gate117inter3), .O(gate117inter5));
  nor2  gate609(.a(gate117inter5), .b(gate117inter2), .O(gate117inter6));
  inv1  gate610(.a(G386), .O(gate117inter7));
  inv1  gate611(.a(G387), .O(gate117inter8));
  nand2 gate612(.a(gate117inter8), .b(gate117inter7), .O(gate117inter9));
  nand2 gate613(.a(s_9), .b(gate117inter3), .O(gate117inter10));
  nor2  gate614(.a(gate117inter10), .b(gate117inter9), .O(gate117inter11));
  nor2  gate615(.a(gate117inter11), .b(gate117inter6), .O(gate117inter12));
  nand2 gate616(.a(gate117inter12), .b(gate117inter1), .O(G462));
nand2 gate118( .a(G388), .b(G389), .O(G465) );
nand2 gate119( .a(G390), .b(G391), .O(G468) );
nand2 gate120( .a(G392), .b(G393), .O(G471) );
nand2 gate121( .a(G394), .b(G395), .O(G474) );
nand2 gate122( .a(G396), .b(G397), .O(G477) );
nand2 gate123( .a(G398), .b(G399), .O(G480) );
nand2 gate124( .a(G400), .b(G401), .O(G483) );
nand2 gate125( .a(G402), .b(G403), .O(G486) );
nand2 gate126( .a(G404), .b(G405), .O(G489) );
nand2 gate127( .a(G406), .b(G407), .O(G492) );
nand2 gate128( .a(G408), .b(G409), .O(G495) );
nand2 gate129( .a(G410), .b(G411), .O(G498) );
nand2 gate130( .a(G412), .b(G413), .O(G501) );
nand2 gate131( .a(G414), .b(G415), .O(G504) );
nand2 gate132( .a(G416), .b(G417), .O(G507) );
nand2 gate133( .a(G418), .b(G419), .O(G510) );
nand2 gate134( .a(G420), .b(G421), .O(G513) );
nand2 gate135( .a(G422), .b(G423), .O(G516) );
nand2 gate136( .a(G424), .b(G425), .O(G519) );
nand2 gate137( .a(G426), .b(G429), .O(G522) );
nand2 gate138( .a(G432), .b(G435), .O(G525) );
nand2 gate139( .a(G438), .b(G441), .O(G528) );
nand2 gate140( .a(G444), .b(G447), .O(G531) );
nand2 gate141( .a(G450), .b(G453), .O(G534) );
nand2 gate142( .a(G456), .b(G459), .O(G537) );
nand2 gate143( .a(G462), .b(G465), .O(G540) );
nand2 gate144( .a(G468), .b(G471), .O(G543) );
nand2 gate145( .a(G474), .b(G477), .O(G546) );
nand2 gate146( .a(G480), .b(G483), .O(G549) );
nand2 gate147( .a(G486), .b(G489), .O(G552) );
nand2 gate148( .a(G492), .b(G495), .O(G555) );

  xor2  gate855(.a(G501), .b(G498), .O(gate149inter0));
  nand2 gate856(.a(gate149inter0), .b(s_44), .O(gate149inter1));
  and2  gate857(.a(G501), .b(G498), .O(gate149inter2));
  inv1  gate858(.a(s_44), .O(gate149inter3));
  inv1  gate859(.a(s_45), .O(gate149inter4));
  nand2 gate860(.a(gate149inter4), .b(gate149inter3), .O(gate149inter5));
  nor2  gate861(.a(gate149inter5), .b(gate149inter2), .O(gate149inter6));
  inv1  gate862(.a(G498), .O(gate149inter7));
  inv1  gate863(.a(G501), .O(gate149inter8));
  nand2 gate864(.a(gate149inter8), .b(gate149inter7), .O(gate149inter9));
  nand2 gate865(.a(s_45), .b(gate149inter3), .O(gate149inter10));
  nor2  gate866(.a(gate149inter10), .b(gate149inter9), .O(gate149inter11));
  nor2  gate867(.a(gate149inter11), .b(gate149inter6), .O(gate149inter12));
  nand2 gate868(.a(gate149inter12), .b(gate149inter1), .O(G558));
nand2 gate150( .a(G504), .b(G507), .O(G561) );
nand2 gate151( .a(G510), .b(G513), .O(G564) );
nand2 gate152( .a(G516), .b(G519), .O(G567) );
nand2 gate153( .a(G426), .b(G522), .O(G570) );
nand2 gate154( .a(G429), .b(G522), .O(G571) );
nand2 gate155( .a(G432), .b(G525), .O(G572) );

  xor2  gate799(.a(G525), .b(G435), .O(gate156inter0));
  nand2 gate800(.a(gate156inter0), .b(s_36), .O(gate156inter1));
  and2  gate801(.a(G525), .b(G435), .O(gate156inter2));
  inv1  gate802(.a(s_36), .O(gate156inter3));
  inv1  gate803(.a(s_37), .O(gate156inter4));
  nand2 gate804(.a(gate156inter4), .b(gate156inter3), .O(gate156inter5));
  nor2  gate805(.a(gate156inter5), .b(gate156inter2), .O(gate156inter6));
  inv1  gate806(.a(G435), .O(gate156inter7));
  inv1  gate807(.a(G525), .O(gate156inter8));
  nand2 gate808(.a(gate156inter8), .b(gate156inter7), .O(gate156inter9));
  nand2 gate809(.a(s_37), .b(gate156inter3), .O(gate156inter10));
  nor2  gate810(.a(gate156inter10), .b(gate156inter9), .O(gate156inter11));
  nor2  gate811(.a(gate156inter11), .b(gate156inter6), .O(gate156inter12));
  nand2 gate812(.a(gate156inter12), .b(gate156inter1), .O(G573));
nand2 gate157( .a(G438), .b(G528), .O(G574) );
nand2 gate158( .a(G441), .b(G528), .O(G575) );
nand2 gate159( .a(G444), .b(G531), .O(G576) );
nand2 gate160( .a(G447), .b(G531), .O(G577) );
nand2 gate161( .a(G450), .b(G534), .O(G578) );
nand2 gate162( .a(G453), .b(G534), .O(G579) );
nand2 gate163( .a(G456), .b(G537), .O(G580) );
nand2 gate164( .a(G459), .b(G537), .O(G581) );
nand2 gate165( .a(G462), .b(G540), .O(G582) );
nand2 gate166( .a(G465), .b(G540), .O(G583) );
nand2 gate167( .a(G468), .b(G543), .O(G584) );
nand2 gate168( .a(G471), .b(G543), .O(G585) );
nand2 gate169( .a(G474), .b(G546), .O(G586) );
nand2 gate170( .a(G477), .b(G546), .O(G587) );
nand2 gate171( .a(G480), .b(G549), .O(G588) );
nand2 gate172( .a(G483), .b(G549), .O(G589) );
nand2 gate173( .a(G486), .b(G552), .O(G590) );
nand2 gate174( .a(G489), .b(G552), .O(G591) );
nand2 gate175( .a(G492), .b(G555), .O(G592) );
nand2 gate176( .a(G495), .b(G555), .O(G593) );
nand2 gate177( .a(G498), .b(G558), .O(G594) );
nand2 gate178( .a(G501), .b(G558), .O(G595) );
nand2 gate179( .a(G504), .b(G561), .O(G596) );
nand2 gate180( .a(G507), .b(G561), .O(G597) );
nand2 gate181( .a(G510), .b(G564), .O(G598) );
nand2 gate182( .a(G513), .b(G564), .O(G599) );

  xor2  gate547(.a(G567), .b(G516), .O(gate183inter0));
  nand2 gate548(.a(gate183inter0), .b(s_0), .O(gate183inter1));
  and2  gate549(.a(G567), .b(G516), .O(gate183inter2));
  inv1  gate550(.a(s_0), .O(gate183inter3));
  inv1  gate551(.a(s_1), .O(gate183inter4));
  nand2 gate552(.a(gate183inter4), .b(gate183inter3), .O(gate183inter5));
  nor2  gate553(.a(gate183inter5), .b(gate183inter2), .O(gate183inter6));
  inv1  gate554(.a(G516), .O(gate183inter7));
  inv1  gate555(.a(G567), .O(gate183inter8));
  nand2 gate556(.a(gate183inter8), .b(gate183inter7), .O(gate183inter9));
  nand2 gate557(.a(s_1), .b(gate183inter3), .O(gate183inter10));
  nor2  gate558(.a(gate183inter10), .b(gate183inter9), .O(gate183inter11));
  nor2  gate559(.a(gate183inter11), .b(gate183inter6), .O(gate183inter12));
  nand2 gate560(.a(gate183inter12), .b(gate183inter1), .O(G600));
nand2 gate184( .a(G519), .b(G567), .O(G601) );
nand2 gate185( .a(G570), .b(G571), .O(G602) );
nand2 gate186( .a(G572), .b(G573), .O(G607) );
nand2 gate187( .a(G574), .b(G575), .O(G612) );
nand2 gate188( .a(G576), .b(G577), .O(G617) );
nand2 gate189( .a(G578), .b(G579), .O(G622) );
nand2 gate190( .a(G580), .b(G581), .O(G627) );
nand2 gate191( .a(G582), .b(G583), .O(G632) );
nand2 gate192( .a(G584), .b(G585), .O(G637) );
nand2 gate193( .a(G586), .b(G587), .O(G642) );
nand2 gate194( .a(G588), .b(G589), .O(G645) );

  xor2  gate897(.a(G591), .b(G590), .O(gate195inter0));
  nand2 gate898(.a(gate195inter0), .b(s_50), .O(gate195inter1));
  and2  gate899(.a(G591), .b(G590), .O(gate195inter2));
  inv1  gate900(.a(s_50), .O(gate195inter3));
  inv1  gate901(.a(s_51), .O(gate195inter4));
  nand2 gate902(.a(gate195inter4), .b(gate195inter3), .O(gate195inter5));
  nor2  gate903(.a(gate195inter5), .b(gate195inter2), .O(gate195inter6));
  inv1  gate904(.a(G590), .O(gate195inter7));
  inv1  gate905(.a(G591), .O(gate195inter8));
  nand2 gate906(.a(gate195inter8), .b(gate195inter7), .O(gate195inter9));
  nand2 gate907(.a(s_51), .b(gate195inter3), .O(gate195inter10));
  nor2  gate908(.a(gate195inter10), .b(gate195inter9), .O(gate195inter11));
  nor2  gate909(.a(gate195inter11), .b(gate195inter6), .O(gate195inter12));
  nand2 gate910(.a(gate195inter12), .b(gate195inter1), .O(G648));
nand2 gate196( .a(G592), .b(G593), .O(G651) );
nand2 gate197( .a(G594), .b(G595), .O(G654) );
nand2 gate198( .a(G596), .b(G597), .O(G657) );
nand2 gate199( .a(G598), .b(G599), .O(G660) );
nand2 gate200( .a(G600), .b(G601), .O(G663) );
nand2 gate201( .a(G602), .b(G607), .O(G666) );
nand2 gate202( .a(G612), .b(G617), .O(G669) );
nand2 gate203( .a(G602), .b(G612), .O(G672) );
nand2 gate204( .a(G607), .b(G617), .O(G675) );
nand2 gate205( .a(G622), .b(G627), .O(G678) );
nand2 gate206( .a(G632), .b(G637), .O(G681) );
nand2 gate207( .a(G622), .b(G632), .O(G684) );
nand2 gate208( .a(G627), .b(G637), .O(G687) );
nand2 gate209( .a(G602), .b(G666), .O(G690) );
nand2 gate210( .a(G607), .b(G666), .O(G691) );

  xor2  gate827(.a(G669), .b(G612), .O(gate211inter0));
  nand2 gate828(.a(gate211inter0), .b(s_40), .O(gate211inter1));
  and2  gate829(.a(G669), .b(G612), .O(gate211inter2));
  inv1  gate830(.a(s_40), .O(gate211inter3));
  inv1  gate831(.a(s_41), .O(gate211inter4));
  nand2 gate832(.a(gate211inter4), .b(gate211inter3), .O(gate211inter5));
  nor2  gate833(.a(gate211inter5), .b(gate211inter2), .O(gate211inter6));
  inv1  gate834(.a(G612), .O(gate211inter7));
  inv1  gate835(.a(G669), .O(gate211inter8));
  nand2 gate836(.a(gate211inter8), .b(gate211inter7), .O(gate211inter9));
  nand2 gate837(.a(s_41), .b(gate211inter3), .O(gate211inter10));
  nor2  gate838(.a(gate211inter10), .b(gate211inter9), .O(gate211inter11));
  nor2  gate839(.a(gate211inter11), .b(gate211inter6), .O(gate211inter12));
  nand2 gate840(.a(gate211inter12), .b(gate211inter1), .O(G692));
nand2 gate212( .a(G617), .b(G669), .O(G693) );
nand2 gate213( .a(G602), .b(G672), .O(G694) );
nand2 gate214( .a(G612), .b(G672), .O(G695) );
nand2 gate215( .a(G607), .b(G675), .O(G696) );
nand2 gate216( .a(G617), .b(G675), .O(G697) );
nand2 gate217( .a(G622), .b(G678), .O(G698) );
nand2 gate218( .a(G627), .b(G678), .O(G699) );
nand2 gate219( .a(G632), .b(G681), .O(G700) );
nand2 gate220( .a(G637), .b(G681), .O(G701) );
nand2 gate221( .a(G622), .b(G684), .O(G702) );
nand2 gate222( .a(G632), .b(G684), .O(G703) );
nand2 gate223( .a(G627), .b(G687), .O(G704) );
nand2 gate224( .a(G637), .b(G687), .O(G705) );
nand2 gate225( .a(G690), .b(G691), .O(G706) );
nand2 gate226( .a(G692), .b(G693), .O(G709) );
nand2 gate227( .a(G694), .b(G695), .O(G712) );
nand2 gate228( .a(G696), .b(G697), .O(G715) );
nand2 gate229( .a(G698), .b(G699), .O(G718) );
nand2 gate230( .a(G700), .b(G701), .O(G721) );
nand2 gate231( .a(G702), .b(G703), .O(G724) );
nand2 gate232( .a(G704), .b(G705), .O(G727) );
nand2 gate233( .a(G242), .b(G718), .O(G730) );
nand2 gate234( .a(G245), .b(G721), .O(G733) );
nand2 gate235( .a(G248), .b(G724), .O(G736) );
nand2 gate236( .a(G251), .b(G727), .O(G739) );
nand2 gate237( .a(G254), .b(G706), .O(G742) );
nand2 gate238( .a(G257), .b(G709), .O(G745) );
nand2 gate239( .a(G260), .b(G712), .O(G748) );
nand2 gate240( .a(G263), .b(G715), .O(G751) );

  xor2  gate673(.a(G730), .b(G242), .O(gate241inter0));
  nand2 gate674(.a(gate241inter0), .b(s_18), .O(gate241inter1));
  and2  gate675(.a(G730), .b(G242), .O(gate241inter2));
  inv1  gate676(.a(s_18), .O(gate241inter3));
  inv1  gate677(.a(s_19), .O(gate241inter4));
  nand2 gate678(.a(gate241inter4), .b(gate241inter3), .O(gate241inter5));
  nor2  gate679(.a(gate241inter5), .b(gate241inter2), .O(gate241inter6));
  inv1  gate680(.a(G242), .O(gate241inter7));
  inv1  gate681(.a(G730), .O(gate241inter8));
  nand2 gate682(.a(gate241inter8), .b(gate241inter7), .O(gate241inter9));
  nand2 gate683(.a(s_19), .b(gate241inter3), .O(gate241inter10));
  nor2  gate684(.a(gate241inter10), .b(gate241inter9), .O(gate241inter11));
  nor2  gate685(.a(gate241inter11), .b(gate241inter6), .O(gate241inter12));
  nand2 gate686(.a(gate241inter12), .b(gate241inter1), .O(G754));
nand2 gate242( .a(G718), .b(G730), .O(G755) );
nand2 gate243( .a(G245), .b(G733), .O(G756) );
nand2 gate244( .a(G721), .b(G733), .O(G757) );
nand2 gate245( .a(G248), .b(G736), .O(G758) );
nand2 gate246( .a(G724), .b(G736), .O(G759) );
nand2 gate247( .a(G251), .b(G739), .O(G760) );
nand2 gate248( .a(G727), .b(G739), .O(G761) );
nand2 gate249( .a(G254), .b(G742), .O(G762) );
nand2 gate250( .a(G706), .b(G742), .O(G763) );
nand2 gate251( .a(G257), .b(G745), .O(G764) );
nand2 gate252( .a(G709), .b(G745), .O(G765) );
nand2 gate253( .a(G260), .b(G748), .O(G766) );
nand2 gate254( .a(G712), .b(G748), .O(G767) );
nand2 gate255( .a(G263), .b(G751), .O(G768) );
nand2 gate256( .a(G715), .b(G751), .O(G769) );
nand2 gate257( .a(G754), .b(G755), .O(G770) );
nand2 gate258( .a(G756), .b(G757), .O(G773) );
nand2 gate259( .a(G758), .b(G759), .O(G776) );
nand2 gate260( .a(G760), .b(G761), .O(G779) );
nand2 gate261( .a(G762), .b(G763), .O(G782) );
nand2 gate262( .a(G764), .b(G765), .O(G785) );
nand2 gate263( .a(G766), .b(G767), .O(G788) );
nand2 gate264( .a(G768), .b(G769), .O(G791) );

  xor2  gate757(.a(G770), .b(G642), .O(gate265inter0));
  nand2 gate758(.a(gate265inter0), .b(s_30), .O(gate265inter1));
  and2  gate759(.a(G770), .b(G642), .O(gate265inter2));
  inv1  gate760(.a(s_30), .O(gate265inter3));
  inv1  gate761(.a(s_31), .O(gate265inter4));
  nand2 gate762(.a(gate265inter4), .b(gate265inter3), .O(gate265inter5));
  nor2  gate763(.a(gate265inter5), .b(gate265inter2), .O(gate265inter6));
  inv1  gate764(.a(G642), .O(gate265inter7));
  inv1  gate765(.a(G770), .O(gate265inter8));
  nand2 gate766(.a(gate265inter8), .b(gate265inter7), .O(gate265inter9));
  nand2 gate767(.a(s_31), .b(gate265inter3), .O(gate265inter10));
  nor2  gate768(.a(gate265inter10), .b(gate265inter9), .O(gate265inter11));
  nor2  gate769(.a(gate265inter11), .b(gate265inter6), .O(gate265inter12));
  nand2 gate770(.a(gate265inter12), .b(gate265inter1), .O(G794));
nand2 gate266( .a(G645), .b(G773), .O(G797) );
nand2 gate267( .a(G648), .b(G776), .O(G800) );
nand2 gate268( .a(G651), .b(G779), .O(G803) );

  xor2  gate883(.a(G782), .b(G654), .O(gate269inter0));
  nand2 gate884(.a(gate269inter0), .b(s_48), .O(gate269inter1));
  and2  gate885(.a(G782), .b(G654), .O(gate269inter2));
  inv1  gate886(.a(s_48), .O(gate269inter3));
  inv1  gate887(.a(s_49), .O(gate269inter4));
  nand2 gate888(.a(gate269inter4), .b(gate269inter3), .O(gate269inter5));
  nor2  gate889(.a(gate269inter5), .b(gate269inter2), .O(gate269inter6));
  inv1  gate890(.a(G654), .O(gate269inter7));
  inv1  gate891(.a(G782), .O(gate269inter8));
  nand2 gate892(.a(gate269inter8), .b(gate269inter7), .O(gate269inter9));
  nand2 gate893(.a(s_49), .b(gate269inter3), .O(gate269inter10));
  nor2  gate894(.a(gate269inter10), .b(gate269inter9), .O(gate269inter11));
  nor2  gate895(.a(gate269inter11), .b(gate269inter6), .O(gate269inter12));
  nand2 gate896(.a(gate269inter12), .b(gate269inter1), .O(G806));
nand2 gate270( .a(G657), .b(G785), .O(G809) );
nand2 gate271( .a(G660), .b(G788), .O(G812) );
nand2 gate272( .a(G663), .b(G791), .O(G815) );
nand2 gate273( .a(G642), .b(G794), .O(G818) );
nand2 gate274( .a(G770), .b(G794), .O(G819) );
nand2 gate275( .a(G645), .b(G797), .O(G820) );
nand2 gate276( .a(G773), .b(G797), .O(G821) );
nand2 gate277( .a(G648), .b(G800), .O(G822) );
nand2 gate278( .a(G776), .b(G800), .O(G823) );

  xor2  gate687(.a(G803), .b(G651), .O(gate279inter0));
  nand2 gate688(.a(gate279inter0), .b(s_20), .O(gate279inter1));
  and2  gate689(.a(G803), .b(G651), .O(gate279inter2));
  inv1  gate690(.a(s_20), .O(gate279inter3));
  inv1  gate691(.a(s_21), .O(gate279inter4));
  nand2 gate692(.a(gate279inter4), .b(gate279inter3), .O(gate279inter5));
  nor2  gate693(.a(gate279inter5), .b(gate279inter2), .O(gate279inter6));
  inv1  gate694(.a(G651), .O(gate279inter7));
  inv1  gate695(.a(G803), .O(gate279inter8));
  nand2 gate696(.a(gate279inter8), .b(gate279inter7), .O(gate279inter9));
  nand2 gate697(.a(s_21), .b(gate279inter3), .O(gate279inter10));
  nor2  gate698(.a(gate279inter10), .b(gate279inter9), .O(gate279inter11));
  nor2  gate699(.a(gate279inter11), .b(gate279inter6), .O(gate279inter12));
  nand2 gate700(.a(gate279inter12), .b(gate279inter1), .O(G824));
nand2 gate280( .a(G779), .b(G803), .O(G825) );
nand2 gate281( .a(G654), .b(G806), .O(G826) );
nand2 gate282( .a(G782), .b(G806), .O(G827) );
nand2 gate283( .a(G657), .b(G809), .O(G828) );
nand2 gate284( .a(G785), .b(G809), .O(G829) );

  xor2  gate659(.a(G812), .b(G660), .O(gate285inter0));
  nand2 gate660(.a(gate285inter0), .b(s_16), .O(gate285inter1));
  and2  gate661(.a(G812), .b(G660), .O(gate285inter2));
  inv1  gate662(.a(s_16), .O(gate285inter3));
  inv1  gate663(.a(s_17), .O(gate285inter4));
  nand2 gate664(.a(gate285inter4), .b(gate285inter3), .O(gate285inter5));
  nor2  gate665(.a(gate285inter5), .b(gate285inter2), .O(gate285inter6));
  inv1  gate666(.a(G660), .O(gate285inter7));
  inv1  gate667(.a(G812), .O(gate285inter8));
  nand2 gate668(.a(gate285inter8), .b(gate285inter7), .O(gate285inter9));
  nand2 gate669(.a(s_17), .b(gate285inter3), .O(gate285inter10));
  nor2  gate670(.a(gate285inter10), .b(gate285inter9), .O(gate285inter11));
  nor2  gate671(.a(gate285inter11), .b(gate285inter6), .O(gate285inter12));
  nand2 gate672(.a(gate285inter12), .b(gate285inter1), .O(G830));
nand2 gate286( .a(G788), .b(G812), .O(G831) );
nand2 gate287( .a(G663), .b(G815), .O(G832) );
nand2 gate288( .a(G791), .b(G815), .O(G833) );

  xor2  gate701(.a(G819), .b(G818), .O(gate289inter0));
  nand2 gate702(.a(gate289inter0), .b(s_22), .O(gate289inter1));
  and2  gate703(.a(G819), .b(G818), .O(gate289inter2));
  inv1  gate704(.a(s_22), .O(gate289inter3));
  inv1  gate705(.a(s_23), .O(gate289inter4));
  nand2 gate706(.a(gate289inter4), .b(gate289inter3), .O(gate289inter5));
  nor2  gate707(.a(gate289inter5), .b(gate289inter2), .O(gate289inter6));
  inv1  gate708(.a(G818), .O(gate289inter7));
  inv1  gate709(.a(G819), .O(gate289inter8));
  nand2 gate710(.a(gate289inter8), .b(gate289inter7), .O(gate289inter9));
  nand2 gate711(.a(s_23), .b(gate289inter3), .O(gate289inter10));
  nor2  gate712(.a(gate289inter10), .b(gate289inter9), .O(gate289inter11));
  nor2  gate713(.a(gate289inter11), .b(gate289inter6), .O(gate289inter12));
  nand2 gate714(.a(gate289inter12), .b(gate289inter1), .O(G834));
nand2 gate290( .a(G820), .b(G821), .O(G847) );
nand2 gate291( .a(G822), .b(G823), .O(G860) );
nand2 gate292( .a(G824), .b(G825), .O(G873) );
nand2 gate293( .a(G828), .b(G829), .O(G886) );
nand2 gate294( .a(G832), .b(G833), .O(G899) );
nand2 gate295( .a(G830), .b(G831), .O(G912) );
nand2 gate296( .a(G826), .b(G827), .O(G925) );
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );
nand2 gate387( .a(G1), .b(G1036), .O(G1132) );
nand2 gate388( .a(G2), .b(G1039), .O(G1135) );
nand2 gate389( .a(G3), .b(G1042), .O(G1138) );
nand2 gate390( .a(G4), .b(G1045), .O(G1141) );
nand2 gate391( .a(G5), .b(G1048), .O(G1144) );
nand2 gate392( .a(G6), .b(G1051), .O(G1147) );
nand2 gate393( .a(G7), .b(G1054), .O(G1150) );
nand2 gate394( .a(G8), .b(G1057), .O(G1153) );

  xor2  gate575(.a(G1060), .b(G9), .O(gate395inter0));
  nand2 gate576(.a(gate395inter0), .b(s_4), .O(gate395inter1));
  and2  gate577(.a(G1060), .b(G9), .O(gate395inter2));
  inv1  gate578(.a(s_4), .O(gate395inter3));
  inv1  gate579(.a(s_5), .O(gate395inter4));
  nand2 gate580(.a(gate395inter4), .b(gate395inter3), .O(gate395inter5));
  nor2  gate581(.a(gate395inter5), .b(gate395inter2), .O(gate395inter6));
  inv1  gate582(.a(G9), .O(gate395inter7));
  inv1  gate583(.a(G1060), .O(gate395inter8));
  nand2 gate584(.a(gate395inter8), .b(gate395inter7), .O(gate395inter9));
  nand2 gate585(.a(s_5), .b(gate395inter3), .O(gate395inter10));
  nor2  gate586(.a(gate395inter10), .b(gate395inter9), .O(gate395inter11));
  nor2  gate587(.a(gate395inter11), .b(gate395inter6), .O(gate395inter12));
  nand2 gate588(.a(gate395inter12), .b(gate395inter1), .O(G1156));
nand2 gate396( .a(G10), .b(G1063), .O(G1159) );
nand2 gate397( .a(G11), .b(G1066), .O(G1162) );
nand2 gate398( .a(G12), .b(G1069), .O(G1165) );
nand2 gate399( .a(G13), .b(G1072), .O(G1168) );
nand2 gate400( .a(G14), .b(G1075), .O(G1171) );
nand2 gate401( .a(G15), .b(G1078), .O(G1174) );
nand2 gate402( .a(G16), .b(G1081), .O(G1177) );
nand2 gate403( .a(G17), .b(G1084), .O(G1180) );
nand2 gate404( .a(G18), .b(G1087), .O(G1183) );
nand2 gate405( .a(G19), .b(G1090), .O(G1186) );

  xor2  gate743(.a(G1093), .b(G20), .O(gate406inter0));
  nand2 gate744(.a(gate406inter0), .b(s_28), .O(gate406inter1));
  and2  gate745(.a(G1093), .b(G20), .O(gate406inter2));
  inv1  gate746(.a(s_28), .O(gate406inter3));
  inv1  gate747(.a(s_29), .O(gate406inter4));
  nand2 gate748(.a(gate406inter4), .b(gate406inter3), .O(gate406inter5));
  nor2  gate749(.a(gate406inter5), .b(gate406inter2), .O(gate406inter6));
  inv1  gate750(.a(G20), .O(gate406inter7));
  inv1  gate751(.a(G1093), .O(gate406inter8));
  nand2 gate752(.a(gate406inter8), .b(gate406inter7), .O(gate406inter9));
  nand2 gate753(.a(s_29), .b(gate406inter3), .O(gate406inter10));
  nor2  gate754(.a(gate406inter10), .b(gate406inter9), .O(gate406inter11));
  nor2  gate755(.a(gate406inter11), .b(gate406inter6), .O(gate406inter12));
  nand2 gate756(.a(gate406inter12), .b(gate406inter1), .O(G1189));
nand2 gate407( .a(G21), .b(G1096), .O(G1192) );
nand2 gate408( .a(G22), .b(G1099), .O(G1195) );
nand2 gate409( .a(G23), .b(G1102), .O(G1198) );
nand2 gate410( .a(G24), .b(G1105), .O(G1201) );
nand2 gate411( .a(G25), .b(G1108), .O(G1204) );
nand2 gate412( .a(G26), .b(G1111), .O(G1207) );
nand2 gate413( .a(G27), .b(G1114), .O(G1210) );
nand2 gate414( .a(G28), .b(G1117), .O(G1213) );
nand2 gate415( .a(G29), .b(G1120), .O(G1216) );
nand2 gate416( .a(G30), .b(G1123), .O(G1219) );
nand2 gate417( .a(G31), .b(G1126), .O(G1222) );
nand2 gate418( .a(G32), .b(G1129), .O(G1225) );
nand2 gate419( .a(G1), .b(G1132), .O(G1228) );
nand2 gate420( .a(G1036), .b(G1132), .O(G1229) );
nand2 gate421( .a(G2), .b(G1135), .O(G1230) );
nand2 gate422( .a(G1039), .b(G1135), .O(G1231) );
nand2 gate423( .a(G3), .b(G1138), .O(G1232) );
nand2 gate424( .a(G1042), .b(G1138), .O(G1233) );
nand2 gate425( .a(G4), .b(G1141), .O(G1234) );
nand2 gate426( .a(G1045), .b(G1141), .O(G1235) );
nand2 gate427( .a(G5), .b(G1144), .O(G1236) );
nand2 gate428( .a(G1048), .b(G1144), .O(G1237) );
nand2 gate429( .a(G6), .b(G1147), .O(G1238) );
nand2 gate430( .a(G1051), .b(G1147), .O(G1239) );
nand2 gate431( .a(G7), .b(G1150), .O(G1240) );
nand2 gate432( .a(G1054), .b(G1150), .O(G1241) );
nand2 gate433( .a(G8), .b(G1153), .O(G1242) );
nand2 gate434( .a(G1057), .b(G1153), .O(G1243) );
nand2 gate435( .a(G9), .b(G1156), .O(G1244) );

  xor2  gate869(.a(G1156), .b(G1060), .O(gate436inter0));
  nand2 gate870(.a(gate436inter0), .b(s_46), .O(gate436inter1));
  and2  gate871(.a(G1156), .b(G1060), .O(gate436inter2));
  inv1  gate872(.a(s_46), .O(gate436inter3));
  inv1  gate873(.a(s_47), .O(gate436inter4));
  nand2 gate874(.a(gate436inter4), .b(gate436inter3), .O(gate436inter5));
  nor2  gate875(.a(gate436inter5), .b(gate436inter2), .O(gate436inter6));
  inv1  gate876(.a(G1060), .O(gate436inter7));
  inv1  gate877(.a(G1156), .O(gate436inter8));
  nand2 gate878(.a(gate436inter8), .b(gate436inter7), .O(gate436inter9));
  nand2 gate879(.a(s_47), .b(gate436inter3), .O(gate436inter10));
  nor2  gate880(.a(gate436inter10), .b(gate436inter9), .O(gate436inter11));
  nor2  gate881(.a(gate436inter11), .b(gate436inter6), .O(gate436inter12));
  nand2 gate882(.a(gate436inter12), .b(gate436inter1), .O(G1245));
nand2 gate437( .a(G10), .b(G1159), .O(G1246) );
nand2 gate438( .a(G1063), .b(G1159), .O(G1247) );
nand2 gate439( .a(G11), .b(G1162), .O(G1248) );
nand2 gate440( .a(G1066), .b(G1162), .O(G1249) );
nand2 gate441( .a(G12), .b(G1165), .O(G1250) );
nand2 gate442( .a(G1069), .b(G1165), .O(G1251) );
nand2 gate443( .a(G13), .b(G1168), .O(G1252) );
nand2 gate444( .a(G1072), .b(G1168), .O(G1253) );
nand2 gate445( .a(G14), .b(G1171), .O(G1254) );
nand2 gate446( .a(G1075), .b(G1171), .O(G1255) );
nand2 gate447( .a(G15), .b(G1174), .O(G1256) );
nand2 gate448( .a(G1078), .b(G1174), .O(G1257) );
nand2 gate449( .a(G16), .b(G1177), .O(G1258) );
nand2 gate450( .a(G1081), .b(G1177), .O(G1259) );
nand2 gate451( .a(G17), .b(G1180), .O(G1260) );
nand2 gate452( .a(G1084), .b(G1180), .O(G1261) );
nand2 gate453( .a(G18), .b(G1183), .O(G1262) );
nand2 gate454( .a(G1087), .b(G1183), .O(G1263) );
nand2 gate455( .a(G19), .b(G1186), .O(G1264) );
nand2 gate456( .a(G1090), .b(G1186), .O(G1265) );
nand2 gate457( .a(G20), .b(G1189), .O(G1266) );
nand2 gate458( .a(G1093), .b(G1189), .O(G1267) );
nand2 gate459( .a(G21), .b(G1192), .O(G1268) );
nand2 gate460( .a(G1096), .b(G1192), .O(G1269) );
nand2 gate461( .a(G22), .b(G1195), .O(G1270) );
nand2 gate462( .a(G1099), .b(G1195), .O(G1271) );
nand2 gate463( .a(G23), .b(G1198), .O(G1272) );
nand2 gate464( .a(G1102), .b(G1198), .O(G1273) );
nand2 gate465( .a(G24), .b(G1201), .O(G1274) );
nand2 gate466( .a(G1105), .b(G1201), .O(G1275) );
nand2 gate467( .a(G25), .b(G1204), .O(G1276) );
nand2 gate468( .a(G1108), .b(G1204), .O(G1277) );
nand2 gate469( .a(G26), .b(G1207), .O(G1278) );
nand2 gate470( .a(G1111), .b(G1207), .O(G1279) );
nand2 gate471( .a(G27), .b(G1210), .O(G1280) );

  xor2  gate729(.a(G1210), .b(G1114), .O(gate472inter0));
  nand2 gate730(.a(gate472inter0), .b(s_26), .O(gate472inter1));
  and2  gate731(.a(G1210), .b(G1114), .O(gate472inter2));
  inv1  gate732(.a(s_26), .O(gate472inter3));
  inv1  gate733(.a(s_27), .O(gate472inter4));
  nand2 gate734(.a(gate472inter4), .b(gate472inter3), .O(gate472inter5));
  nor2  gate735(.a(gate472inter5), .b(gate472inter2), .O(gate472inter6));
  inv1  gate736(.a(G1114), .O(gate472inter7));
  inv1  gate737(.a(G1210), .O(gate472inter8));
  nand2 gate738(.a(gate472inter8), .b(gate472inter7), .O(gate472inter9));
  nand2 gate739(.a(s_27), .b(gate472inter3), .O(gate472inter10));
  nor2  gate740(.a(gate472inter10), .b(gate472inter9), .O(gate472inter11));
  nor2  gate741(.a(gate472inter11), .b(gate472inter6), .O(gate472inter12));
  nand2 gate742(.a(gate472inter12), .b(gate472inter1), .O(G1281));
nand2 gate473( .a(G28), .b(G1213), .O(G1282) );
nand2 gate474( .a(G1117), .b(G1213), .O(G1283) );
nand2 gate475( .a(G29), .b(G1216), .O(G1284) );
nand2 gate476( .a(G1120), .b(G1216), .O(G1285) );
nand2 gate477( .a(G30), .b(G1219), .O(G1286) );
nand2 gate478( .a(G1123), .b(G1219), .O(G1287) );
nand2 gate479( .a(G31), .b(G1222), .O(G1288) );
nand2 gate480( .a(G1126), .b(G1222), .O(G1289) );
nand2 gate481( .a(G32), .b(G1225), .O(G1290) );
nand2 gate482( .a(G1129), .b(G1225), .O(G1291) );
nand2 gate483( .a(G1228), .b(G1229), .O(G1292) );
nand2 gate484( .a(G1230), .b(G1231), .O(G1293) );
nand2 gate485( .a(G1232), .b(G1233), .O(G1294) );
nand2 gate486( .a(G1234), .b(G1235), .O(G1295) );
nand2 gate487( .a(G1236), .b(G1237), .O(G1296) );
nand2 gate488( .a(G1238), .b(G1239), .O(G1297) );
nand2 gate489( .a(G1240), .b(G1241), .O(G1298) );
nand2 gate490( .a(G1242), .b(G1243), .O(G1299) );
nand2 gate491( .a(G1244), .b(G1245), .O(G1300) );
nand2 gate492( .a(G1246), .b(G1247), .O(G1301) );
nand2 gate493( .a(G1248), .b(G1249), .O(G1302) );
nand2 gate494( .a(G1250), .b(G1251), .O(G1303) );
nand2 gate495( .a(G1252), .b(G1253), .O(G1304) );
nand2 gate496( .a(G1254), .b(G1255), .O(G1305) );
nand2 gate497( .a(G1256), .b(G1257), .O(G1306) );
nand2 gate498( .a(G1258), .b(G1259), .O(G1307) );
nand2 gate499( .a(G1260), .b(G1261), .O(G1308) );
nand2 gate500( .a(G1262), .b(G1263), .O(G1309) );
nand2 gate501( .a(G1264), .b(G1265), .O(G1310) );
nand2 gate502( .a(G1266), .b(G1267), .O(G1311) );
nand2 gate503( .a(G1268), .b(G1269), .O(G1312) );
nand2 gate504( .a(G1270), .b(G1271), .O(G1313) );
nand2 gate505( .a(G1272), .b(G1273), .O(G1314) );
nand2 gate506( .a(G1274), .b(G1275), .O(G1315) );
nand2 gate507( .a(G1276), .b(G1277), .O(G1316) );
nand2 gate508( .a(G1278), .b(G1279), .O(G1317) );
nand2 gate509( .a(G1280), .b(G1281), .O(G1318) );
nand2 gate510( .a(G1282), .b(G1283), .O(G1319) );
nand2 gate511( .a(G1284), .b(G1285), .O(G1320) );
nand2 gate512( .a(G1286), .b(G1287), .O(G1321) );
nand2 gate513( .a(G1288), .b(G1289), .O(G1322) );
nand2 gate514( .a(G1290), .b(G1291), .O(G1323) );
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule