module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);

input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;//RE__PI;

input s_0,s_1;//RE__ALLOW(00,01,10,11);
input s_2,s_3;//RE__ALLOW(00,01,10,11);
input s_4,s_5;//RE__ALLOW(00,01,10,11);
input s_6,s_7;//RE__ALLOW(00,01,10,11);
input s_8,s_9;//RE__ALLOW(00,01,10,11);
input s_10,s_11;//RE__ALLOW(00,01,10,11);
input s_12,s_13;//RE__ALLOW(00,01,10,11);
input s_14,s_15;//RE__ALLOW(00,01,10,11);
input s_16,s_17;//RE__ALLOW(00,01,10,11);
input s_18,s_19;//RE__ALLOW(00,01,10,11);
input s_20,s_21;//RE__ALLOW(00,01,10,11);
input s_22,s_23;//RE__ALLOW(00,01,10,11);
input s_24,s_25;//RE__ALLOW(00,01,10,11);
input s_26,s_27;//RE__ALLOW(00,01,10,11);
input s_28,s_29;//RE__ALLOW(00,01,10,11);
input s_30,s_31;//RE__ALLOW(00,01,10,11);
input s_32,s_33;//RE__ALLOW(00,01,10,11);
input s_34,s_35;//RE__ALLOW(00,01,10,11);
input s_36,s_37;//RE__ALLOW(00,01,10,11);
input s_38,s_39;//RE__ALLOW(00,01,10,11);
input s_40,s_41;//RE__ALLOW(00,01,10,11);
input s_42,s_43;//RE__ALLOW(00,01,10,11);
input s_44,s_45;//RE__ALLOW(00,01,10,11);
input s_46,s_47;//RE__ALLOW(00,01,10,11);
input s_48,s_49;//RE__ALLOW(00,01,10,11);
input s_50,s_51;//RE__ALLOW(00,01,10,11);
input s_52,s_53;//RE__ALLOW(00,01,10,11);
input s_54,s_55;//RE__ALLOW(00,01,10,11);
input s_56,s_57;//RE__ALLOW(00,01,10,11);
input s_58,s_59;//RE__ALLOW(00,01,10,11);
input s_60,s_61;//RE__ALLOW(00,01,10,11);
input s_62,s_63;//RE__ALLOW(00,01,10,11);
input s_64,s_65;//RE__ALLOW(00,01,10,11);
input s_66,s_67;//RE__ALLOW(00,01,10,11);
input s_68,s_69;//RE__ALLOW(00,01,10,11);
input s_70,s_71;//RE__ALLOW(00,01,10,11);
input s_72,s_73;//RE__ALLOW(00,01,10,11);
input s_74,s_75;//RE__ALLOW(00,01,10,11);
input s_76,s_77;//RE__ALLOW(00,01,10,11);
input s_78,s_79;//RE__ALLOW(00,01,10,11);
input s_80,s_81;//RE__ALLOW(00,01,10,11);
input s_82,s_83;//RE__ALLOW(00,01,10,11);
input s_84,s_85;//RE__ALLOW(00,01,10,11);
input s_86,s_87;//RE__ALLOW(00,01,10,11);
input s_88,s_89;//RE__ALLOW(00,01,10,11);
input s_90,s_91;//RE__ALLOW(00,01,10,11);
input s_92,s_93;//RE__ALLOW(00,01,10,11);
input s_94,s_95;//RE__ALLOW(00,01,10,11);
input s_96,s_97;//RE__ALLOW(00,01,10,11);
input s_98,s_99;//RE__ALLOW(00,01,10,11);
input s_100,s_101;//RE__ALLOW(00,01,10,11);
input s_102,s_103;//RE__ALLOW(00,01,10,11);
input s_104,s_105;//RE__ALLOW(00,01,10,11);
input s_106,s_107;//RE__ALLOW(00,01,10,11);
input s_108,s_109;//RE__ALLOW(00,01,10,11);
input s_110,s_111;//RE__ALLOW(00,01,10,11);
input s_112,s_113;//RE__ALLOW(00,01,10,11);
input s_114,s_115;//RE__ALLOW(00,01,10,11);
input s_116,s_117;//RE__ALLOW(00,01,10,11);
input s_118,s_119;//RE__ALLOW(00,01,10,11);
input s_120,s_121;//RE__ALLOW(00,01,10,11);
input s_122,s_123;//RE__ALLOW(00,01,10,11);
input s_124,s_125;//RE__ALLOW(00,01,10,11);
input s_126,s_127;//RE__ALLOW(00,01,10,11);
input s_128,s_129;//RE__ALLOW(00,01,10,11);
input s_130,s_131;//RE__ALLOW(00,01,10,11);
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;

  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate419inter0, gate419inter1, gate419inter2, gate419inter3, gate419inter4, gate419inter5, gate419inter6, gate419inter7, gate419inter8, gate419inter9, gate419inter10, gate419inter11, gate419inter12, gate277inter0, gate277inter1, gate277inter2, gate277inter3, gate277inter4, gate277inter5, gate277inter6, gate277inter7, gate277inter8, gate277inter9, gate277inter10, gate277inter11, gate277inter12, gate506inter0, gate506inter1, gate506inter2, gate506inter3, gate506inter4, gate506inter5, gate506inter6, gate506inter7, gate506inter8, gate506inter9, gate506inter10, gate506inter11, gate506inter12, gate215inter0, gate215inter1, gate215inter2, gate215inter3, gate215inter4, gate215inter5, gate215inter6, gate215inter7, gate215inter8, gate215inter9, gate215inter10, gate215inter11, gate215inter12, gate428inter0, gate428inter1, gate428inter2, gate428inter3, gate428inter4, gate428inter5, gate428inter6, gate428inter7, gate428inter8, gate428inter9, gate428inter10, gate428inter11, gate428inter12, gate417inter0, gate417inter1, gate417inter2, gate417inter3, gate417inter4, gate417inter5, gate417inter6, gate417inter7, gate417inter8, gate417inter9, gate417inter10, gate417inter11, gate417inter12, gate236inter0, gate236inter1, gate236inter2, gate236inter3, gate236inter4, gate236inter5, gate236inter6, gate236inter7, gate236inter8, gate236inter9, gate236inter10, gate236inter11, gate236inter12, gate291inter0, gate291inter1, gate291inter2, gate291inter3, gate291inter4, gate291inter5, gate291inter6, gate291inter7, gate291inter8, gate291inter9, gate291inter10, gate291inter11, gate291inter12, gate93inter0, gate93inter1, gate93inter2, gate93inter3, gate93inter4, gate93inter5, gate93inter6, gate93inter7, gate93inter8, gate93inter9, gate93inter10, gate93inter11, gate93inter12, gate104inter0, gate104inter1, gate104inter2, gate104inter3, gate104inter4, gate104inter5, gate104inter6, gate104inter7, gate104inter8, gate104inter9, gate104inter10, gate104inter11, gate104inter12, gate78inter0, gate78inter1, gate78inter2, gate78inter3, gate78inter4, gate78inter5, gate78inter6, gate78inter7, gate78inter8, gate78inter9, gate78inter10, gate78inter11, gate78inter12, gate17inter0, gate17inter1, gate17inter2, gate17inter3, gate17inter4, gate17inter5, gate17inter6, gate17inter7, gate17inter8, gate17inter9, gate17inter10, gate17inter11, gate17inter12, gate473inter0, gate473inter1, gate473inter2, gate473inter3, gate473inter4, gate473inter5, gate473inter6, gate473inter7, gate473inter8, gate473inter9, gate473inter10, gate473inter11, gate473inter12, gate289inter0, gate289inter1, gate289inter2, gate289inter3, gate289inter4, gate289inter5, gate289inter6, gate289inter7, gate289inter8, gate289inter9, gate289inter10, gate289inter11, gate289inter12, gate250inter0, gate250inter1, gate250inter2, gate250inter3, gate250inter4, gate250inter5, gate250inter6, gate250inter7, gate250inter8, gate250inter9, gate250inter10, gate250inter11, gate250inter12, gate415inter0, gate415inter1, gate415inter2, gate415inter3, gate415inter4, gate415inter5, gate415inter6, gate415inter7, gate415inter8, gate415inter9, gate415inter10, gate415inter11, gate415inter12, gate193inter0, gate193inter1, gate193inter2, gate193inter3, gate193inter4, gate193inter5, gate193inter6, gate193inter7, gate193inter8, gate193inter9, gate193inter10, gate193inter11, gate193inter12, gate287inter0, gate287inter1, gate287inter2, gate287inter3, gate287inter4, gate287inter5, gate287inter6, gate287inter7, gate287inter8, gate287inter9, gate287inter10, gate287inter11, gate287inter12, gate135inter0, gate135inter1, gate135inter2, gate135inter3, gate135inter4, gate135inter5, gate135inter6, gate135inter7, gate135inter8, gate135inter9, gate135inter10, gate135inter11, gate135inter12, gate449inter0, gate449inter1, gate449inter2, gate449inter3, gate449inter4, gate449inter5, gate449inter6, gate449inter7, gate449inter8, gate449inter9, gate449inter10, gate449inter11, gate449inter12, gate407inter0, gate407inter1, gate407inter2, gate407inter3, gate407inter4, gate407inter5, gate407inter6, gate407inter7, gate407inter8, gate407inter9, gate407inter10, gate407inter11, gate407inter12, gate79inter0, gate79inter1, gate79inter2, gate79inter3, gate79inter4, gate79inter5, gate79inter6, gate79inter7, gate79inter8, gate79inter9, gate79inter10, gate79inter11, gate79inter12, gate445inter0, gate445inter1, gate445inter2, gate445inter3, gate445inter4, gate445inter5, gate445inter6, gate445inter7, gate445inter8, gate445inter9, gate445inter10, gate445inter11, gate445inter12, gate471inter0, gate471inter1, gate471inter2, gate471inter3, gate471inter4, gate471inter5, gate471inter6, gate471inter7, gate471inter8, gate471inter9, gate471inter10, gate471inter11, gate471inter12, gate121inter0, gate121inter1, gate121inter2, gate121inter3, gate121inter4, gate121inter5, gate121inter6, gate121inter7, gate121inter8, gate121inter9, gate121inter10, gate121inter11, gate121inter12, gate65inter0, gate65inter1, gate65inter2, gate65inter3, gate65inter4, gate65inter5, gate65inter6, gate65inter7, gate65inter8, gate65inter9, gate65inter10, gate65inter11, gate65inter12, gate390inter0, gate390inter1, gate390inter2, gate390inter3, gate390inter4, gate390inter5, gate390inter6, gate390inter7, gate390inter8, gate390inter9, gate390inter10, gate390inter11, gate390inter12, gate254inter0, gate254inter1, gate254inter2, gate254inter3, gate254inter4, gate254inter5, gate254inter6, gate254inter7, gate254inter8, gate254inter9, gate254inter10, gate254inter11, gate254inter12, gate457inter0, gate457inter1, gate457inter2, gate457inter3, gate457inter4, gate457inter5, gate457inter6, gate457inter7, gate457inter8, gate457inter9, gate457inter10, gate457inter11, gate457inter12, gate30inter0, gate30inter1, gate30inter2, gate30inter3, gate30inter4, gate30inter5, gate30inter6, gate30inter7, gate30inter8, gate30inter9, gate30inter10, gate30inter11, gate30inter12, gate458inter0, gate458inter1, gate458inter2, gate458inter3, gate458inter4, gate458inter5, gate458inter6, gate458inter7, gate458inter8, gate458inter9, gate458inter10, gate458inter11, gate458inter12, gate153inter0, gate153inter1, gate153inter2, gate153inter3, gate153inter4, gate153inter5, gate153inter6, gate153inter7, gate153inter8, gate153inter9, gate153inter10, gate153inter11, gate153inter12, gate460inter0, gate460inter1, gate460inter2, gate460inter3, gate460inter4, gate460inter5, gate460inter6, gate460inter7, gate460inter8, gate460inter9, gate460inter10, gate460inter11, gate460inter12, gate444inter0, gate444inter1, gate444inter2, gate444inter3, gate444inter4, gate444inter5, gate444inter6, gate444inter7, gate444inter8, gate444inter9, gate444inter10, gate444inter11, gate444inter12, gate139inter0, gate139inter1, gate139inter2, gate139inter3, gate139inter4, gate139inter5, gate139inter6, gate139inter7, gate139inter8, gate139inter9, gate139inter10, gate139inter11, gate139inter12, gate448inter0, gate448inter1, gate448inter2, gate448inter3, gate448inter4, gate448inter5, gate448inter6, gate448inter7, gate448inter8, gate448inter9, gate448inter10, gate448inter11, gate448inter12, gate465inter0, gate465inter1, gate465inter2, gate465inter3, gate465inter4, gate465inter5, gate465inter6, gate465inter7, gate465inter8, gate465inter9, gate465inter10, gate465inter11, gate465inter12, gate127inter0, gate127inter1, gate127inter2, gate127inter3, gate127inter4, gate127inter5, gate127inter6, gate127inter7, gate127inter8, gate127inter9, gate127inter10, gate127inter11, gate127inter12, gate159inter0, gate159inter1, gate159inter2, gate159inter3, gate159inter4, gate159inter5, gate159inter6, gate159inter7, gate159inter8, gate159inter9, gate159inter10, gate159inter11, gate159inter12, gate27inter0, gate27inter1, gate27inter2, gate27inter3, gate27inter4, gate27inter5, gate27inter6, gate27inter7, gate27inter8, gate27inter9, gate27inter10, gate27inter11, gate27inter12, gate256inter0, gate256inter1, gate256inter2, gate256inter3, gate256inter4, gate256inter5, gate256inter6, gate256inter7, gate256inter8, gate256inter9, gate256inter10, gate256inter11, gate256inter12, gate491inter0, gate491inter1, gate491inter2, gate491inter3, gate491inter4, gate491inter5, gate491inter6, gate491inter7, gate491inter8, gate491inter9, gate491inter10, gate491inter11, gate491inter12, gate44inter0, gate44inter1, gate44inter2, gate44inter3, gate44inter4, gate44inter5, gate44inter6, gate44inter7, gate44inter8, gate44inter9, gate44inter10, gate44inter11, gate44inter12, gate18inter0, gate18inter1, gate18inter2, gate18inter3, gate18inter4, gate18inter5, gate18inter6, gate18inter7, gate18inter8, gate18inter9, gate18inter10, gate18inter11, gate18inter12, gate467inter0, gate467inter1, gate467inter2, gate467inter3, gate467inter4, gate467inter5, gate467inter6, gate467inter7, gate467inter8, gate467inter9, gate467inter10, gate467inter11, gate467inter12, gate32inter0, gate32inter1, gate32inter2, gate32inter3, gate32inter4, gate32inter5, gate32inter6, gate32inter7, gate32inter8, gate32inter9, gate32inter10, gate32inter11, gate32inter12, gate177inter0, gate177inter1, gate177inter2, gate177inter3, gate177inter4, gate177inter5, gate177inter6, gate177inter7, gate177inter8, gate177inter9, gate177inter10, gate177inter11, gate177inter12, gate242inter0, gate242inter1, gate242inter2, gate242inter3, gate242inter4, gate242inter5, gate242inter6, gate242inter7, gate242inter8, gate242inter9, gate242inter10, gate242inter11, gate242inter12, gate469inter0, gate469inter1, gate469inter2, gate469inter3, gate469inter4, gate469inter5, gate469inter6, gate469inter7, gate469inter8, gate469inter9, gate469inter10, gate469inter11, gate469inter12, gate432inter0, gate432inter1, gate432inter2, gate432inter3, gate432inter4, gate432inter5, gate432inter6, gate432inter7, gate432inter8, gate432inter9, gate432inter10, gate432inter11, gate432inter12, gate282inter0, gate282inter1, gate282inter2, gate282inter3, gate282inter4, gate282inter5, gate282inter6, gate282inter7, gate282inter8, gate282inter9, gate282inter10, gate282inter11, gate282inter12, gate403inter0, gate403inter1, gate403inter2, gate403inter3, gate403inter4, gate403inter5, gate403inter6, gate403inter7, gate403inter8, gate403inter9, gate403inter10, gate403inter11, gate403inter12, gate278inter0, gate278inter1, gate278inter2, gate278inter3, gate278inter4, gate278inter5, gate278inter6, gate278inter7, gate278inter8, gate278inter9, gate278inter10, gate278inter11, gate278inter12, gate113inter0, gate113inter1, gate113inter2, gate113inter3, gate113inter4, gate113inter5, gate113inter6, gate113inter7, gate113inter8, gate113inter9, gate113inter10, gate113inter11, gate113inter12, gate69inter0, gate69inter1, gate69inter2, gate69inter3, gate69inter4, gate69inter5, gate69inter6, gate69inter7, gate69inter8, gate69inter9, gate69inter10, gate69inter11, gate69inter12, gate55inter0, gate55inter1, gate55inter2, gate55inter3, gate55inter4, gate55inter5, gate55inter6, gate55inter7, gate55inter8, gate55inter9, gate55inter10, gate55inter11, gate55inter12, gate393inter0, gate393inter1, gate393inter2, gate393inter3, gate393inter4, gate393inter5, gate393inter6, gate393inter7, gate393inter8, gate393inter9, gate393inter10, gate393inter11, gate393inter12, gate200inter0, gate200inter1, gate200inter2, gate200inter3, gate200inter4, gate200inter5, gate200inter6, gate200inter7, gate200inter8, gate200inter9, gate200inter10, gate200inter11, gate200inter12, gate513inter0, gate513inter1, gate513inter2, gate513inter3, gate513inter4, gate513inter5, gate513inter6, gate513inter7, gate513inter8, gate513inter9, gate513inter10, gate513inter11, gate513inter12, gate204inter0, gate204inter1, gate204inter2, gate204inter3, gate204inter4, gate204inter5, gate204inter6, gate204inter7, gate204inter8, gate204inter9, gate204inter10, gate204inter11, gate204inter12, gate100inter0, gate100inter1, gate100inter2, gate100inter3, gate100inter4, gate100inter5, gate100inter6, gate100inter7, gate100inter8, gate100inter9, gate100inter10, gate100inter11, gate100inter12, gate272inter0, gate272inter1, gate272inter2, gate272inter3, gate272inter4, gate272inter5, gate272inter6, gate272inter7, gate272inter8, gate272inter9, gate272inter10, gate272inter11, gate272inter12, gate179inter0, gate179inter1, gate179inter2, gate179inter3, gate179inter4, gate179inter5, gate179inter6, gate179inter7, gate179inter8, gate179inter9, gate179inter10, gate179inter11, gate179inter12, gate151inter0, gate151inter1, gate151inter2, gate151inter3, gate151inter4, gate151inter5, gate151inter6, gate151inter7, gate151inter8, gate151inter9, gate151inter10, gate151inter11, gate151inter12, gate35inter0, gate35inter1, gate35inter2, gate35inter3, gate35inter4, gate35inter5, gate35inter6, gate35inter7, gate35inter8, gate35inter9, gate35inter10, gate35inter11, gate35inter12, gate99inter0, gate99inter1, gate99inter2, gate99inter3, gate99inter4, gate99inter5, gate99inter6, gate99inter7, gate99inter8, gate99inter9, gate99inter10, gate99inter11, gate99inter12;



and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );
nand2 gate9( .a(G1), .b(G2), .O(G266) );
nand2 gate10( .a(G3), .b(G4), .O(G269) );
nand2 gate11( .a(G5), .b(G6), .O(G272) );
nand2 gate12( .a(G7), .b(G8), .O(G275) );
nand2 gate13( .a(G9), .b(G10), .O(G278) );
nand2 gate14( .a(G11), .b(G12), .O(G281) );
nand2 gate15( .a(G13), .b(G14), .O(G284) );
nand2 gate16( .a(G15), .b(G16), .O(G287) );

  xor2  gate701(.a(G18), .b(G17), .O(gate17inter0));
  nand2 gate702(.a(gate17inter0), .b(s_22), .O(gate17inter1));
  and2  gate703(.a(G18), .b(G17), .O(gate17inter2));
  inv1  gate704(.a(s_22), .O(gate17inter3));
  inv1  gate705(.a(s_23), .O(gate17inter4));
  nand2 gate706(.a(gate17inter4), .b(gate17inter3), .O(gate17inter5));
  nor2  gate707(.a(gate17inter5), .b(gate17inter2), .O(gate17inter6));
  inv1  gate708(.a(G17), .O(gate17inter7));
  inv1  gate709(.a(G18), .O(gate17inter8));
  nand2 gate710(.a(gate17inter8), .b(gate17inter7), .O(gate17inter9));
  nand2 gate711(.a(s_23), .b(gate17inter3), .O(gate17inter10));
  nor2  gate712(.a(gate17inter10), .b(gate17inter9), .O(gate17inter11));
  nor2  gate713(.a(gate17inter11), .b(gate17inter6), .O(gate17inter12));
  nand2 gate714(.a(gate17inter12), .b(gate17inter1), .O(G290));

  xor2  gate1149(.a(G20), .b(G19), .O(gate18inter0));
  nand2 gate1150(.a(gate18inter0), .b(s_86), .O(gate18inter1));
  and2  gate1151(.a(G20), .b(G19), .O(gate18inter2));
  inv1  gate1152(.a(s_86), .O(gate18inter3));
  inv1  gate1153(.a(s_87), .O(gate18inter4));
  nand2 gate1154(.a(gate18inter4), .b(gate18inter3), .O(gate18inter5));
  nor2  gate1155(.a(gate18inter5), .b(gate18inter2), .O(gate18inter6));
  inv1  gate1156(.a(G19), .O(gate18inter7));
  inv1  gate1157(.a(G20), .O(gate18inter8));
  nand2 gate1158(.a(gate18inter8), .b(gate18inter7), .O(gate18inter9));
  nand2 gate1159(.a(s_87), .b(gate18inter3), .O(gate18inter10));
  nor2  gate1160(.a(gate18inter10), .b(gate18inter9), .O(gate18inter11));
  nor2  gate1161(.a(gate18inter11), .b(gate18inter6), .O(gate18inter12));
  nand2 gate1162(.a(gate18inter12), .b(gate18inter1), .O(G293));
nand2 gate19( .a(G21), .b(G22), .O(G296) );
nand2 gate20( .a(G23), .b(G24), .O(G299) );
nand2 gate21( .a(G25), .b(G26), .O(G302) );
nand2 gate22( .a(G27), .b(G28), .O(G305) );
nand2 gate23( .a(G29), .b(G30), .O(G308) );
nand2 gate24( .a(G31), .b(G32), .O(G311) );
nand2 gate25( .a(G1), .b(G5), .O(G314) );
nand2 gate26( .a(G9), .b(G13), .O(G317) );

  xor2  gate1093(.a(G6), .b(G2), .O(gate27inter0));
  nand2 gate1094(.a(gate27inter0), .b(s_78), .O(gate27inter1));
  and2  gate1095(.a(G6), .b(G2), .O(gate27inter2));
  inv1  gate1096(.a(s_78), .O(gate27inter3));
  inv1  gate1097(.a(s_79), .O(gate27inter4));
  nand2 gate1098(.a(gate27inter4), .b(gate27inter3), .O(gate27inter5));
  nor2  gate1099(.a(gate27inter5), .b(gate27inter2), .O(gate27inter6));
  inv1  gate1100(.a(G2), .O(gate27inter7));
  inv1  gate1101(.a(G6), .O(gate27inter8));
  nand2 gate1102(.a(gate27inter8), .b(gate27inter7), .O(gate27inter9));
  nand2 gate1103(.a(s_79), .b(gate27inter3), .O(gate27inter10));
  nor2  gate1104(.a(gate27inter10), .b(gate27inter9), .O(gate27inter11));
  nor2  gate1105(.a(gate27inter11), .b(gate27inter6), .O(gate27inter12));
  nand2 gate1106(.a(gate27inter12), .b(gate27inter1), .O(G320));
nand2 gate28( .a(G10), .b(G14), .O(G323) );
nand2 gate29( .a(G3), .b(G7), .O(G326) );

  xor2  gate953(.a(G15), .b(G11), .O(gate30inter0));
  nand2 gate954(.a(gate30inter0), .b(s_58), .O(gate30inter1));
  and2  gate955(.a(G15), .b(G11), .O(gate30inter2));
  inv1  gate956(.a(s_58), .O(gate30inter3));
  inv1  gate957(.a(s_59), .O(gate30inter4));
  nand2 gate958(.a(gate30inter4), .b(gate30inter3), .O(gate30inter5));
  nor2  gate959(.a(gate30inter5), .b(gate30inter2), .O(gate30inter6));
  inv1  gate960(.a(G11), .O(gate30inter7));
  inv1  gate961(.a(G15), .O(gate30inter8));
  nand2 gate962(.a(gate30inter8), .b(gate30inter7), .O(gate30inter9));
  nand2 gate963(.a(s_59), .b(gate30inter3), .O(gate30inter10));
  nor2  gate964(.a(gate30inter10), .b(gate30inter9), .O(gate30inter11));
  nor2  gate965(.a(gate30inter11), .b(gate30inter6), .O(gate30inter12));
  nand2 gate966(.a(gate30inter12), .b(gate30inter1), .O(G329));
nand2 gate31( .a(G4), .b(G8), .O(G332) );

  xor2  gate1177(.a(G16), .b(G12), .O(gate32inter0));
  nand2 gate1178(.a(gate32inter0), .b(s_90), .O(gate32inter1));
  and2  gate1179(.a(G16), .b(G12), .O(gate32inter2));
  inv1  gate1180(.a(s_90), .O(gate32inter3));
  inv1  gate1181(.a(s_91), .O(gate32inter4));
  nand2 gate1182(.a(gate32inter4), .b(gate32inter3), .O(gate32inter5));
  nor2  gate1183(.a(gate32inter5), .b(gate32inter2), .O(gate32inter6));
  inv1  gate1184(.a(G12), .O(gate32inter7));
  inv1  gate1185(.a(G16), .O(gate32inter8));
  nand2 gate1186(.a(gate32inter8), .b(gate32inter7), .O(gate32inter9));
  nand2 gate1187(.a(s_91), .b(gate32inter3), .O(gate32inter10));
  nor2  gate1188(.a(gate32inter10), .b(gate32inter9), .O(gate32inter11));
  nor2  gate1189(.a(gate32inter11), .b(gate32inter6), .O(gate32inter12));
  nand2 gate1190(.a(gate32inter12), .b(gate32inter1), .O(G335));
nand2 gate33( .a(G17), .b(G21), .O(G338) );
nand2 gate34( .a(G25), .b(G29), .O(G341) );

  xor2  gate1443(.a(G22), .b(G18), .O(gate35inter0));
  nand2 gate1444(.a(gate35inter0), .b(s_128), .O(gate35inter1));
  and2  gate1445(.a(G22), .b(G18), .O(gate35inter2));
  inv1  gate1446(.a(s_128), .O(gate35inter3));
  inv1  gate1447(.a(s_129), .O(gate35inter4));
  nand2 gate1448(.a(gate35inter4), .b(gate35inter3), .O(gate35inter5));
  nor2  gate1449(.a(gate35inter5), .b(gate35inter2), .O(gate35inter6));
  inv1  gate1450(.a(G18), .O(gate35inter7));
  inv1  gate1451(.a(G22), .O(gate35inter8));
  nand2 gate1452(.a(gate35inter8), .b(gate35inter7), .O(gate35inter9));
  nand2 gate1453(.a(s_129), .b(gate35inter3), .O(gate35inter10));
  nor2  gate1454(.a(gate35inter10), .b(gate35inter9), .O(gate35inter11));
  nor2  gate1455(.a(gate35inter11), .b(gate35inter6), .O(gate35inter12));
  nand2 gate1456(.a(gate35inter12), .b(gate35inter1), .O(G344));
nand2 gate36( .a(G26), .b(G30), .O(G347) );
nand2 gate37( .a(G19), .b(G23), .O(G350) );
nand2 gate38( .a(G27), .b(G31), .O(G353) );
nand2 gate39( .a(G20), .b(G24), .O(G356) );
nand2 gate40( .a(G28), .b(G32), .O(G359) );
nand2 gate41( .a(G1), .b(G266), .O(G362) );
nand2 gate42( .a(G2), .b(G266), .O(G363) );
nand2 gate43( .a(G3), .b(G269), .O(G364) );

  xor2  gate1135(.a(G269), .b(G4), .O(gate44inter0));
  nand2 gate1136(.a(gate44inter0), .b(s_84), .O(gate44inter1));
  and2  gate1137(.a(G269), .b(G4), .O(gate44inter2));
  inv1  gate1138(.a(s_84), .O(gate44inter3));
  inv1  gate1139(.a(s_85), .O(gate44inter4));
  nand2 gate1140(.a(gate44inter4), .b(gate44inter3), .O(gate44inter5));
  nor2  gate1141(.a(gate44inter5), .b(gate44inter2), .O(gate44inter6));
  inv1  gate1142(.a(G4), .O(gate44inter7));
  inv1  gate1143(.a(G269), .O(gate44inter8));
  nand2 gate1144(.a(gate44inter8), .b(gate44inter7), .O(gate44inter9));
  nand2 gate1145(.a(s_85), .b(gate44inter3), .O(gate44inter10));
  nor2  gate1146(.a(gate44inter10), .b(gate44inter9), .O(gate44inter11));
  nor2  gate1147(.a(gate44inter11), .b(gate44inter6), .O(gate44inter12));
  nand2 gate1148(.a(gate44inter12), .b(gate44inter1), .O(G365));
nand2 gate45( .a(G5), .b(G272), .O(G366) );
nand2 gate46( .a(G6), .b(G272), .O(G367) );
nand2 gate47( .a(G7), .b(G275), .O(G368) );
nand2 gate48( .a(G8), .b(G275), .O(G369) );
nand2 gate49( .a(G9), .b(G278), .O(G370) );
nand2 gate50( .a(G10), .b(G278), .O(G371) );
nand2 gate51( .a(G11), .b(G281), .O(G372) );
nand2 gate52( .a(G12), .b(G281), .O(G373) );
nand2 gate53( .a(G13), .b(G284), .O(G374) );
nand2 gate54( .a(G14), .b(G284), .O(G375) );

  xor2  gate1317(.a(G287), .b(G15), .O(gate55inter0));
  nand2 gate1318(.a(gate55inter0), .b(s_110), .O(gate55inter1));
  and2  gate1319(.a(G287), .b(G15), .O(gate55inter2));
  inv1  gate1320(.a(s_110), .O(gate55inter3));
  inv1  gate1321(.a(s_111), .O(gate55inter4));
  nand2 gate1322(.a(gate55inter4), .b(gate55inter3), .O(gate55inter5));
  nor2  gate1323(.a(gate55inter5), .b(gate55inter2), .O(gate55inter6));
  inv1  gate1324(.a(G15), .O(gate55inter7));
  inv1  gate1325(.a(G287), .O(gate55inter8));
  nand2 gate1326(.a(gate55inter8), .b(gate55inter7), .O(gate55inter9));
  nand2 gate1327(.a(s_111), .b(gate55inter3), .O(gate55inter10));
  nor2  gate1328(.a(gate55inter10), .b(gate55inter9), .O(gate55inter11));
  nor2  gate1329(.a(gate55inter11), .b(gate55inter6), .O(gate55inter12));
  nand2 gate1330(.a(gate55inter12), .b(gate55inter1), .O(G376));
nand2 gate56( .a(G16), .b(G287), .O(G377) );
nand2 gate57( .a(G17), .b(G290), .O(G378) );
nand2 gate58( .a(G18), .b(G290), .O(G379) );
nand2 gate59( .a(G19), .b(G293), .O(G380) );
nand2 gate60( .a(G20), .b(G293), .O(G381) );
nand2 gate61( .a(G21), .b(G296), .O(G382) );
nand2 gate62( .a(G22), .b(G296), .O(G383) );
nand2 gate63( .a(G23), .b(G299), .O(G384) );
nand2 gate64( .a(G24), .b(G299), .O(G385) );

  xor2  gate897(.a(G302), .b(G25), .O(gate65inter0));
  nand2 gate898(.a(gate65inter0), .b(s_50), .O(gate65inter1));
  and2  gate899(.a(G302), .b(G25), .O(gate65inter2));
  inv1  gate900(.a(s_50), .O(gate65inter3));
  inv1  gate901(.a(s_51), .O(gate65inter4));
  nand2 gate902(.a(gate65inter4), .b(gate65inter3), .O(gate65inter5));
  nor2  gate903(.a(gate65inter5), .b(gate65inter2), .O(gate65inter6));
  inv1  gate904(.a(G25), .O(gate65inter7));
  inv1  gate905(.a(G302), .O(gate65inter8));
  nand2 gate906(.a(gate65inter8), .b(gate65inter7), .O(gate65inter9));
  nand2 gate907(.a(s_51), .b(gate65inter3), .O(gate65inter10));
  nor2  gate908(.a(gate65inter10), .b(gate65inter9), .O(gate65inter11));
  nor2  gate909(.a(gate65inter11), .b(gate65inter6), .O(gate65inter12));
  nand2 gate910(.a(gate65inter12), .b(gate65inter1), .O(G386));
nand2 gate66( .a(G26), .b(G302), .O(G387) );
nand2 gate67( .a(G27), .b(G305), .O(G388) );
nand2 gate68( .a(G28), .b(G305), .O(G389) );

  xor2  gate1303(.a(G308), .b(G29), .O(gate69inter0));
  nand2 gate1304(.a(gate69inter0), .b(s_108), .O(gate69inter1));
  and2  gate1305(.a(G308), .b(G29), .O(gate69inter2));
  inv1  gate1306(.a(s_108), .O(gate69inter3));
  inv1  gate1307(.a(s_109), .O(gate69inter4));
  nand2 gate1308(.a(gate69inter4), .b(gate69inter3), .O(gate69inter5));
  nor2  gate1309(.a(gate69inter5), .b(gate69inter2), .O(gate69inter6));
  inv1  gate1310(.a(G29), .O(gate69inter7));
  inv1  gate1311(.a(G308), .O(gate69inter8));
  nand2 gate1312(.a(gate69inter8), .b(gate69inter7), .O(gate69inter9));
  nand2 gate1313(.a(s_109), .b(gate69inter3), .O(gate69inter10));
  nor2  gate1314(.a(gate69inter10), .b(gate69inter9), .O(gate69inter11));
  nor2  gate1315(.a(gate69inter11), .b(gate69inter6), .O(gate69inter12));
  nand2 gate1316(.a(gate69inter12), .b(gate69inter1), .O(G390));
nand2 gate70( .a(G30), .b(G308), .O(G391) );
nand2 gate71( .a(G31), .b(G311), .O(G392) );
nand2 gate72( .a(G32), .b(G311), .O(G393) );
nand2 gate73( .a(G1), .b(G314), .O(G394) );
nand2 gate74( .a(G5), .b(G314), .O(G395) );
nand2 gate75( .a(G9), .b(G317), .O(G396) );
nand2 gate76( .a(G13), .b(G317), .O(G397) );
nand2 gate77( .a(G2), .b(G320), .O(G398) );

  xor2  gate687(.a(G320), .b(G6), .O(gate78inter0));
  nand2 gate688(.a(gate78inter0), .b(s_20), .O(gate78inter1));
  and2  gate689(.a(G320), .b(G6), .O(gate78inter2));
  inv1  gate690(.a(s_20), .O(gate78inter3));
  inv1  gate691(.a(s_21), .O(gate78inter4));
  nand2 gate692(.a(gate78inter4), .b(gate78inter3), .O(gate78inter5));
  nor2  gate693(.a(gate78inter5), .b(gate78inter2), .O(gate78inter6));
  inv1  gate694(.a(G6), .O(gate78inter7));
  inv1  gate695(.a(G320), .O(gate78inter8));
  nand2 gate696(.a(gate78inter8), .b(gate78inter7), .O(gate78inter9));
  nand2 gate697(.a(s_21), .b(gate78inter3), .O(gate78inter10));
  nor2  gate698(.a(gate78inter10), .b(gate78inter9), .O(gate78inter11));
  nor2  gate699(.a(gate78inter11), .b(gate78inter6), .O(gate78inter12));
  nand2 gate700(.a(gate78inter12), .b(gate78inter1), .O(G399));

  xor2  gate841(.a(G323), .b(G10), .O(gate79inter0));
  nand2 gate842(.a(gate79inter0), .b(s_42), .O(gate79inter1));
  and2  gate843(.a(G323), .b(G10), .O(gate79inter2));
  inv1  gate844(.a(s_42), .O(gate79inter3));
  inv1  gate845(.a(s_43), .O(gate79inter4));
  nand2 gate846(.a(gate79inter4), .b(gate79inter3), .O(gate79inter5));
  nor2  gate847(.a(gate79inter5), .b(gate79inter2), .O(gate79inter6));
  inv1  gate848(.a(G10), .O(gate79inter7));
  inv1  gate849(.a(G323), .O(gate79inter8));
  nand2 gate850(.a(gate79inter8), .b(gate79inter7), .O(gate79inter9));
  nand2 gate851(.a(s_43), .b(gate79inter3), .O(gate79inter10));
  nor2  gate852(.a(gate79inter10), .b(gate79inter9), .O(gate79inter11));
  nor2  gate853(.a(gate79inter11), .b(gate79inter6), .O(gate79inter12));
  nand2 gate854(.a(gate79inter12), .b(gate79inter1), .O(G400));
nand2 gate80( .a(G14), .b(G323), .O(G401) );
nand2 gate81( .a(G3), .b(G326), .O(G402) );
nand2 gate82( .a(G7), .b(G326), .O(G403) );
nand2 gate83( .a(G11), .b(G329), .O(G404) );
nand2 gate84( .a(G15), .b(G329), .O(G405) );
nand2 gate85( .a(G4), .b(G332), .O(G406) );
nand2 gate86( .a(G8), .b(G332), .O(G407) );
nand2 gate87( .a(G12), .b(G335), .O(G408) );
nand2 gate88( .a(G16), .b(G335), .O(G409) );
nand2 gate89( .a(G17), .b(G338), .O(G410) );
nand2 gate90( .a(G21), .b(G338), .O(G411) );
nand2 gate91( .a(G25), .b(G341), .O(G412) );
nand2 gate92( .a(G29), .b(G341), .O(G413) );

  xor2  gate659(.a(G344), .b(G18), .O(gate93inter0));
  nand2 gate660(.a(gate93inter0), .b(s_16), .O(gate93inter1));
  and2  gate661(.a(G344), .b(G18), .O(gate93inter2));
  inv1  gate662(.a(s_16), .O(gate93inter3));
  inv1  gate663(.a(s_17), .O(gate93inter4));
  nand2 gate664(.a(gate93inter4), .b(gate93inter3), .O(gate93inter5));
  nor2  gate665(.a(gate93inter5), .b(gate93inter2), .O(gate93inter6));
  inv1  gate666(.a(G18), .O(gate93inter7));
  inv1  gate667(.a(G344), .O(gate93inter8));
  nand2 gate668(.a(gate93inter8), .b(gate93inter7), .O(gate93inter9));
  nand2 gate669(.a(s_17), .b(gate93inter3), .O(gate93inter10));
  nor2  gate670(.a(gate93inter10), .b(gate93inter9), .O(gate93inter11));
  nor2  gate671(.a(gate93inter11), .b(gate93inter6), .O(gate93inter12));
  nand2 gate672(.a(gate93inter12), .b(gate93inter1), .O(G414));
nand2 gate94( .a(G22), .b(G344), .O(G415) );
nand2 gate95( .a(G26), .b(G347), .O(G416) );
nand2 gate96( .a(G30), .b(G347), .O(G417) );
nand2 gate97( .a(G19), .b(G350), .O(G418) );
nand2 gate98( .a(G23), .b(G350), .O(G419) );

  xor2  gate1457(.a(G353), .b(G27), .O(gate99inter0));
  nand2 gate1458(.a(gate99inter0), .b(s_130), .O(gate99inter1));
  and2  gate1459(.a(G353), .b(G27), .O(gate99inter2));
  inv1  gate1460(.a(s_130), .O(gate99inter3));
  inv1  gate1461(.a(s_131), .O(gate99inter4));
  nand2 gate1462(.a(gate99inter4), .b(gate99inter3), .O(gate99inter5));
  nor2  gate1463(.a(gate99inter5), .b(gate99inter2), .O(gate99inter6));
  inv1  gate1464(.a(G27), .O(gate99inter7));
  inv1  gate1465(.a(G353), .O(gate99inter8));
  nand2 gate1466(.a(gate99inter8), .b(gate99inter7), .O(gate99inter9));
  nand2 gate1467(.a(s_131), .b(gate99inter3), .O(gate99inter10));
  nor2  gate1468(.a(gate99inter10), .b(gate99inter9), .O(gate99inter11));
  nor2  gate1469(.a(gate99inter11), .b(gate99inter6), .O(gate99inter12));
  nand2 gate1470(.a(gate99inter12), .b(gate99inter1), .O(G420));

  xor2  gate1387(.a(G353), .b(G31), .O(gate100inter0));
  nand2 gate1388(.a(gate100inter0), .b(s_120), .O(gate100inter1));
  and2  gate1389(.a(G353), .b(G31), .O(gate100inter2));
  inv1  gate1390(.a(s_120), .O(gate100inter3));
  inv1  gate1391(.a(s_121), .O(gate100inter4));
  nand2 gate1392(.a(gate100inter4), .b(gate100inter3), .O(gate100inter5));
  nor2  gate1393(.a(gate100inter5), .b(gate100inter2), .O(gate100inter6));
  inv1  gate1394(.a(G31), .O(gate100inter7));
  inv1  gate1395(.a(G353), .O(gate100inter8));
  nand2 gate1396(.a(gate100inter8), .b(gate100inter7), .O(gate100inter9));
  nand2 gate1397(.a(s_121), .b(gate100inter3), .O(gate100inter10));
  nor2  gate1398(.a(gate100inter10), .b(gate100inter9), .O(gate100inter11));
  nor2  gate1399(.a(gate100inter11), .b(gate100inter6), .O(gate100inter12));
  nand2 gate1400(.a(gate100inter12), .b(gate100inter1), .O(G421));
nand2 gate101( .a(G20), .b(G356), .O(G422) );
nand2 gate102( .a(G24), .b(G356), .O(G423) );
nand2 gate103( .a(G28), .b(G359), .O(G424) );

  xor2  gate673(.a(G359), .b(G32), .O(gate104inter0));
  nand2 gate674(.a(gate104inter0), .b(s_18), .O(gate104inter1));
  and2  gate675(.a(G359), .b(G32), .O(gate104inter2));
  inv1  gate676(.a(s_18), .O(gate104inter3));
  inv1  gate677(.a(s_19), .O(gate104inter4));
  nand2 gate678(.a(gate104inter4), .b(gate104inter3), .O(gate104inter5));
  nor2  gate679(.a(gate104inter5), .b(gate104inter2), .O(gate104inter6));
  inv1  gate680(.a(G32), .O(gate104inter7));
  inv1  gate681(.a(G359), .O(gate104inter8));
  nand2 gate682(.a(gate104inter8), .b(gate104inter7), .O(gate104inter9));
  nand2 gate683(.a(s_19), .b(gate104inter3), .O(gate104inter10));
  nor2  gate684(.a(gate104inter10), .b(gate104inter9), .O(gate104inter11));
  nor2  gate685(.a(gate104inter11), .b(gate104inter6), .O(gate104inter12));
  nand2 gate686(.a(gate104inter12), .b(gate104inter1), .O(G425));
nand2 gate105( .a(G362), .b(G363), .O(G426) );
nand2 gate106( .a(G364), .b(G365), .O(G429) );
nand2 gate107( .a(G366), .b(G367), .O(G432) );
nand2 gate108( .a(G368), .b(G369), .O(G435) );
nand2 gate109( .a(G370), .b(G371), .O(G438) );
nand2 gate110( .a(G372), .b(G373), .O(G441) );
nand2 gate111( .a(G374), .b(G375), .O(G444) );
nand2 gate112( .a(G376), .b(G377), .O(G447) );

  xor2  gate1289(.a(G379), .b(G378), .O(gate113inter0));
  nand2 gate1290(.a(gate113inter0), .b(s_106), .O(gate113inter1));
  and2  gate1291(.a(G379), .b(G378), .O(gate113inter2));
  inv1  gate1292(.a(s_106), .O(gate113inter3));
  inv1  gate1293(.a(s_107), .O(gate113inter4));
  nand2 gate1294(.a(gate113inter4), .b(gate113inter3), .O(gate113inter5));
  nor2  gate1295(.a(gate113inter5), .b(gate113inter2), .O(gate113inter6));
  inv1  gate1296(.a(G378), .O(gate113inter7));
  inv1  gate1297(.a(G379), .O(gate113inter8));
  nand2 gate1298(.a(gate113inter8), .b(gate113inter7), .O(gate113inter9));
  nand2 gate1299(.a(s_107), .b(gate113inter3), .O(gate113inter10));
  nor2  gate1300(.a(gate113inter10), .b(gate113inter9), .O(gate113inter11));
  nor2  gate1301(.a(gate113inter11), .b(gate113inter6), .O(gate113inter12));
  nand2 gate1302(.a(gate113inter12), .b(gate113inter1), .O(G450));
nand2 gate114( .a(G380), .b(G381), .O(G453) );
nand2 gate115( .a(G382), .b(G383), .O(G456) );
nand2 gate116( .a(G384), .b(G385), .O(G459) );
nand2 gate117( .a(G386), .b(G387), .O(G462) );
nand2 gate118( .a(G388), .b(G389), .O(G465) );
nand2 gate119( .a(G390), .b(G391), .O(G468) );
nand2 gate120( .a(G392), .b(G393), .O(G471) );

  xor2  gate883(.a(G395), .b(G394), .O(gate121inter0));
  nand2 gate884(.a(gate121inter0), .b(s_48), .O(gate121inter1));
  and2  gate885(.a(G395), .b(G394), .O(gate121inter2));
  inv1  gate886(.a(s_48), .O(gate121inter3));
  inv1  gate887(.a(s_49), .O(gate121inter4));
  nand2 gate888(.a(gate121inter4), .b(gate121inter3), .O(gate121inter5));
  nor2  gate889(.a(gate121inter5), .b(gate121inter2), .O(gate121inter6));
  inv1  gate890(.a(G394), .O(gate121inter7));
  inv1  gate891(.a(G395), .O(gate121inter8));
  nand2 gate892(.a(gate121inter8), .b(gate121inter7), .O(gate121inter9));
  nand2 gate893(.a(s_49), .b(gate121inter3), .O(gate121inter10));
  nor2  gate894(.a(gate121inter10), .b(gate121inter9), .O(gate121inter11));
  nor2  gate895(.a(gate121inter11), .b(gate121inter6), .O(gate121inter12));
  nand2 gate896(.a(gate121inter12), .b(gate121inter1), .O(G474));
nand2 gate122( .a(G396), .b(G397), .O(G477) );
nand2 gate123( .a(G398), .b(G399), .O(G480) );
nand2 gate124( .a(G400), .b(G401), .O(G483) );
nand2 gate125( .a(G402), .b(G403), .O(G486) );
nand2 gate126( .a(G404), .b(G405), .O(G489) );

  xor2  gate1065(.a(G407), .b(G406), .O(gate127inter0));
  nand2 gate1066(.a(gate127inter0), .b(s_74), .O(gate127inter1));
  and2  gate1067(.a(G407), .b(G406), .O(gate127inter2));
  inv1  gate1068(.a(s_74), .O(gate127inter3));
  inv1  gate1069(.a(s_75), .O(gate127inter4));
  nand2 gate1070(.a(gate127inter4), .b(gate127inter3), .O(gate127inter5));
  nor2  gate1071(.a(gate127inter5), .b(gate127inter2), .O(gate127inter6));
  inv1  gate1072(.a(G406), .O(gate127inter7));
  inv1  gate1073(.a(G407), .O(gate127inter8));
  nand2 gate1074(.a(gate127inter8), .b(gate127inter7), .O(gate127inter9));
  nand2 gate1075(.a(s_75), .b(gate127inter3), .O(gate127inter10));
  nor2  gate1076(.a(gate127inter10), .b(gate127inter9), .O(gate127inter11));
  nor2  gate1077(.a(gate127inter11), .b(gate127inter6), .O(gate127inter12));
  nand2 gate1078(.a(gate127inter12), .b(gate127inter1), .O(G492));
nand2 gate128( .a(G408), .b(G409), .O(G495) );
nand2 gate129( .a(G410), .b(G411), .O(G498) );
nand2 gate130( .a(G412), .b(G413), .O(G501) );
nand2 gate131( .a(G414), .b(G415), .O(G504) );
nand2 gate132( .a(G416), .b(G417), .O(G507) );
nand2 gate133( .a(G418), .b(G419), .O(G510) );
nand2 gate134( .a(G420), .b(G421), .O(G513) );

  xor2  gate799(.a(G423), .b(G422), .O(gate135inter0));
  nand2 gate800(.a(gate135inter0), .b(s_36), .O(gate135inter1));
  and2  gate801(.a(G423), .b(G422), .O(gate135inter2));
  inv1  gate802(.a(s_36), .O(gate135inter3));
  inv1  gate803(.a(s_37), .O(gate135inter4));
  nand2 gate804(.a(gate135inter4), .b(gate135inter3), .O(gate135inter5));
  nor2  gate805(.a(gate135inter5), .b(gate135inter2), .O(gate135inter6));
  inv1  gate806(.a(G422), .O(gate135inter7));
  inv1  gate807(.a(G423), .O(gate135inter8));
  nand2 gate808(.a(gate135inter8), .b(gate135inter7), .O(gate135inter9));
  nand2 gate809(.a(s_37), .b(gate135inter3), .O(gate135inter10));
  nor2  gate810(.a(gate135inter10), .b(gate135inter9), .O(gate135inter11));
  nor2  gate811(.a(gate135inter11), .b(gate135inter6), .O(gate135inter12));
  nand2 gate812(.a(gate135inter12), .b(gate135inter1), .O(G516));
nand2 gate136( .a(G424), .b(G425), .O(G519) );
nand2 gate137( .a(G426), .b(G429), .O(G522) );
nand2 gate138( .a(G432), .b(G435), .O(G525) );

  xor2  gate1023(.a(G441), .b(G438), .O(gate139inter0));
  nand2 gate1024(.a(gate139inter0), .b(s_68), .O(gate139inter1));
  and2  gate1025(.a(G441), .b(G438), .O(gate139inter2));
  inv1  gate1026(.a(s_68), .O(gate139inter3));
  inv1  gate1027(.a(s_69), .O(gate139inter4));
  nand2 gate1028(.a(gate139inter4), .b(gate139inter3), .O(gate139inter5));
  nor2  gate1029(.a(gate139inter5), .b(gate139inter2), .O(gate139inter6));
  inv1  gate1030(.a(G438), .O(gate139inter7));
  inv1  gate1031(.a(G441), .O(gate139inter8));
  nand2 gate1032(.a(gate139inter8), .b(gate139inter7), .O(gate139inter9));
  nand2 gate1033(.a(s_69), .b(gate139inter3), .O(gate139inter10));
  nor2  gate1034(.a(gate139inter10), .b(gate139inter9), .O(gate139inter11));
  nor2  gate1035(.a(gate139inter11), .b(gate139inter6), .O(gate139inter12));
  nand2 gate1036(.a(gate139inter12), .b(gate139inter1), .O(G528));
nand2 gate140( .a(G444), .b(G447), .O(G531) );
nand2 gate141( .a(G450), .b(G453), .O(G534) );
nand2 gate142( .a(G456), .b(G459), .O(G537) );
nand2 gate143( .a(G462), .b(G465), .O(G540) );
nand2 gate144( .a(G468), .b(G471), .O(G543) );
nand2 gate145( .a(G474), .b(G477), .O(G546) );
nand2 gate146( .a(G480), .b(G483), .O(G549) );
nand2 gate147( .a(G486), .b(G489), .O(G552) );
nand2 gate148( .a(G492), .b(G495), .O(G555) );
nand2 gate149( .a(G498), .b(G501), .O(G558) );
nand2 gate150( .a(G504), .b(G507), .O(G561) );

  xor2  gate1429(.a(G513), .b(G510), .O(gate151inter0));
  nand2 gate1430(.a(gate151inter0), .b(s_126), .O(gate151inter1));
  and2  gate1431(.a(G513), .b(G510), .O(gate151inter2));
  inv1  gate1432(.a(s_126), .O(gate151inter3));
  inv1  gate1433(.a(s_127), .O(gate151inter4));
  nand2 gate1434(.a(gate151inter4), .b(gate151inter3), .O(gate151inter5));
  nor2  gate1435(.a(gate151inter5), .b(gate151inter2), .O(gate151inter6));
  inv1  gate1436(.a(G510), .O(gate151inter7));
  inv1  gate1437(.a(G513), .O(gate151inter8));
  nand2 gate1438(.a(gate151inter8), .b(gate151inter7), .O(gate151inter9));
  nand2 gate1439(.a(s_127), .b(gate151inter3), .O(gate151inter10));
  nor2  gate1440(.a(gate151inter10), .b(gate151inter9), .O(gate151inter11));
  nor2  gate1441(.a(gate151inter11), .b(gate151inter6), .O(gate151inter12));
  nand2 gate1442(.a(gate151inter12), .b(gate151inter1), .O(G564));
nand2 gate152( .a(G516), .b(G519), .O(G567) );

  xor2  gate981(.a(G522), .b(G426), .O(gate153inter0));
  nand2 gate982(.a(gate153inter0), .b(s_62), .O(gate153inter1));
  and2  gate983(.a(G522), .b(G426), .O(gate153inter2));
  inv1  gate984(.a(s_62), .O(gate153inter3));
  inv1  gate985(.a(s_63), .O(gate153inter4));
  nand2 gate986(.a(gate153inter4), .b(gate153inter3), .O(gate153inter5));
  nor2  gate987(.a(gate153inter5), .b(gate153inter2), .O(gate153inter6));
  inv1  gate988(.a(G426), .O(gate153inter7));
  inv1  gate989(.a(G522), .O(gate153inter8));
  nand2 gate990(.a(gate153inter8), .b(gate153inter7), .O(gate153inter9));
  nand2 gate991(.a(s_63), .b(gate153inter3), .O(gate153inter10));
  nor2  gate992(.a(gate153inter10), .b(gate153inter9), .O(gate153inter11));
  nor2  gate993(.a(gate153inter11), .b(gate153inter6), .O(gate153inter12));
  nand2 gate994(.a(gate153inter12), .b(gate153inter1), .O(G570));
nand2 gate154( .a(G429), .b(G522), .O(G571) );
nand2 gate155( .a(G432), .b(G525), .O(G572) );
nand2 gate156( .a(G435), .b(G525), .O(G573) );
nand2 gate157( .a(G438), .b(G528), .O(G574) );
nand2 gate158( .a(G441), .b(G528), .O(G575) );

  xor2  gate1079(.a(G531), .b(G444), .O(gate159inter0));
  nand2 gate1080(.a(gate159inter0), .b(s_76), .O(gate159inter1));
  and2  gate1081(.a(G531), .b(G444), .O(gate159inter2));
  inv1  gate1082(.a(s_76), .O(gate159inter3));
  inv1  gate1083(.a(s_77), .O(gate159inter4));
  nand2 gate1084(.a(gate159inter4), .b(gate159inter3), .O(gate159inter5));
  nor2  gate1085(.a(gate159inter5), .b(gate159inter2), .O(gate159inter6));
  inv1  gate1086(.a(G444), .O(gate159inter7));
  inv1  gate1087(.a(G531), .O(gate159inter8));
  nand2 gate1088(.a(gate159inter8), .b(gate159inter7), .O(gate159inter9));
  nand2 gate1089(.a(s_77), .b(gate159inter3), .O(gate159inter10));
  nor2  gate1090(.a(gate159inter10), .b(gate159inter9), .O(gate159inter11));
  nor2  gate1091(.a(gate159inter11), .b(gate159inter6), .O(gate159inter12));
  nand2 gate1092(.a(gate159inter12), .b(gate159inter1), .O(G576));
nand2 gate160( .a(G447), .b(G531), .O(G577) );
nand2 gate161( .a(G450), .b(G534), .O(G578) );
nand2 gate162( .a(G453), .b(G534), .O(G579) );
nand2 gate163( .a(G456), .b(G537), .O(G580) );
nand2 gate164( .a(G459), .b(G537), .O(G581) );
nand2 gate165( .a(G462), .b(G540), .O(G582) );
nand2 gate166( .a(G465), .b(G540), .O(G583) );
nand2 gate167( .a(G468), .b(G543), .O(G584) );
nand2 gate168( .a(G471), .b(G543), .O(G585) );
nand2 gate169( .a(G474), .b(G546), .O(G586) );
nand2 gate170( .a(G477), .b(G546), .O(G587) );
nand2 gate171( .a(G480), .b(G549), .O(G588) );
nand2 gate172( .a(G483), .b(G549), .O(G589) );
nand2 gate173( .a(G486), .b(G552), .O(G590) );
nand2 gate174( .a(G489), .b(G552), .O(G591) );
nand2 gate175( .a(G492), .b(G555), .O(G592) );
nand2 gate176( .a(G495), .b(G555), .O(G593) );

  xor2  gate1191(.a(G558), .b(G498), .O(gate177inter0));
  nand2 gate1192(.a(gate177inter0), .b(s_92), .O(gate177inter1));
  and2  gate1193(.a(G558), .b(G498), .O(gate177inter2));
  inv1  gate1194(.a(s_92), .O(gate177inter3));
  inv1  gate1195(.a(s_93), .O(gate177inter4));
  nand2 gate1196(.a(gate177inter4), .b(gate177inter3), .O(gate177inter5));
  nor2  gate1197(.a(gate177inter5), .b(gate177inter2), .O(gate177inter6));
  inv1  gate1198(.a(G498), .O(gate177inter7));
  inv1  gate1199(.a(G558), .O(gate177inter8));
  nand2 gate1200(.a(gate177inter8), .b(gate177inter7), .O(gate177inter9));
  nand2 gate1201(.a(s_93), .b(gate177inter3), .O(gate177inter10));
  nor2  gate1202(.a(gate177inter10), .b(gate177inter9), .O(gate177inter11));
  nor2  gate1203(.a(gate177inter11), .b(gate177inter6), .O(gate177inter12));
  nand2 gate1204(.a(gate177inter12), .b(gate177inter1), .O(G594));
nand2 gate178( .a(G501), .b(G558), .O(G595) );

  xor2  gate1415(.a(G561), .b(G504), .O(gate179inter0));
  nand2 gate1416(.a(gate179inter0), .b(s_124), .O(gate179inter1));
  and2  gate1417(.a(G561), .b(G504), .O(gate179inter2));
  inv1  gate1418(.a(s_124), .O(gate179inter3));
  inv1  gate1419(.a(s_125), .O(gate179inter4));
  nand2 gate1420(.a(gate179inter4), .b(gate179inter3), .O(gate179inter5));
  nor2  gate1421(.a(gate179inter5), .b(gate179inter2), .O(gate179inter6));
  inv1  gate1422(.a(G504), .O(gate179inter7));
  inv1  gate1423(.a(G561), .O(gate179inter8));
  nand2 gate1424(.a(gate179inter8), .b(gate179inter7), .O(gate179inter9));
  nand2 gate1425(.a(s_125), .b(gate179inter3), .O(gate179inter10));
  nor2  gate1426(.a(gate179inter10), .b(gate179inter9), .O(gate179inter11));
  nor2  gate1427(.a(gate179inter11), .b(gate179inter6), .O(gate179inter12));
  nand2 gate1428(.a(gate179inter12), .b(gate179inter1), .O(G596));
nand2 gate180( .a(G507), .b(G561), .O(G597) );
nand2 gate181( .a(G510), .b(G564), .O(G598) );
nand2 gate182( .a(G513), .b(G564), .O(G599) );
nand2 gate183( .a(G516), .b(G567), .O(G600) );
nand2 gate184( .a(G519), .b(G567), .O(G601) );
nand2 gate185( .a(G570), .b(G571), .O(G602) );
nand2 gate186( .a(G572), .b(G573), .O(G607) );
nand2 gate187( .a(G574), .b(G575), .O(G612) );
nand2 gate188( .a(G576), .b(G577), .O(G617) );
nand2 gate189( .a(G578), .b(G579), .O(G622) );
nand2 gate190( .a(G580), .b(G581), .O(G627) );
nand2 gate191( .a(G582), .b(G583), .O(G632) );
nand2 gate192( .a(G584), .b(G585), .O(G637) );

  xor2  gate771(.a(G587), .b(G586), .O(gate193inter0));
  nand2 gate772(.a(gate193inter0), .b(s_32), .O(gate193inter1));
  and2  gate773(.a(G587), .b(G586), .O(gate193inter2));
  inv1  gate774(.a(s_32), .O(gate193inter3));
  inv1  gate775(.a(s_33), .O(gate193inter4));
  nand2 gate776(.a(gate193inter4), .b(gate193inter3), .O(gate193inter5));
  nor2  gate777(.a(gate193inter5), .b(gate193inter2), .O(gate193inter6));
  inv1  gate778(.a(G586), .O(gate193inter7));
  inv1  gate779(.a(G587), .O(gate193inter8));
  nand2 gate780(.a(gate193inter8), .b(gate193inter7), .O(gate193inter9));
  nand2 gate781(.a(s_33), .b(gate193inter3), .O(gate193inter10));
  nor2  gate782(.a(gate193inter10), .b(gate193inter9), .O(gate193inter11));
  nor2  gate783(.a(gate193inter11), .b(gate193inter6), .O(gate193inter12));
  nand2 gate784(.a(gate193inter12), .b(gate193inter1), .O(G642));
nand2 gate194( .a(G588), .b(G589), .O(G645) );
nand2 gate195( .a(G590), .b(G591), .O(G648) );
nand2 gate196( .a(G592), .b(G593), .O(G651) );
nand2 gate197( .a(G594), .b(G595), .O(G654) );
nand2 gate198( .a(G596), .b(G597), .O(G657) );
nand2 gate199( .a(G598), .b(G599), .O(G660) );

  xor2  gate1345(.a(G601), .b(G600), .O(gate200inter0));
  nand2 gate1346(.a(gate200inter0), .b(s_114), .O(gate200inter1));
  and2  gate1347(.a(G601), .b(G600), .O(gate200inter2));
  inv1  gate1348(.a(s_114), .O(gate200inter3));
  inv1  gate1349(.a(s_115), .O(gate200inter4));
  nand2 gate1350(.a(gate200inter4), .b(gate200inter3), .O(gate200inter5));
  nor2  gate1351(.a(gate200inter5), .b(gate200inter2), .O(gate200inter6));
  inv1  gate1352(.a(G600), .O(gate200inter7));
  inv1  gate1353(.a(G601), .O(gate200inter8));
  nand2 gate1354(.a(gate200inter8), .b(gate200inter7), .O(gate200inter9));
  nand2 gate1355(.a(s_115), .b(gate200inter3), .O(gate200inter10));
  nor2  gate1356(.a(gate200inter10), .b(gate200inter9), .O(gate200inter11));
  nor2  gate1357(.a(gate200inter11), .b(gate200inter6), .O(gate200inter12));
  nand2 gate1358(.a(gate200inter12), .b(gate200inter1), .O(G663));
nand2 gate201( .a(G602), .b(G607), .O(G666) );
nand2 gate202( .a(G612), .b(G617), .O(G669) );
nand2 gate203( .a(G602), .b(G612), .O(G672) );

  xor2  gate1373(.a(G617), .b(G607), .O(gate204inter0));
  nand2 gate1374(.a(gate204inter0), .b(s_118), .O(gate204inter1));
  and2  gate1375(.a(G617), .b(G607), .O(gate204inter2));
  inv1  gate1376(.a(s_118), .O(gate204inter3));
  inv1  gate1377(.a(s_119), .O(gate204inter4));
  nand2 gate1378(.a(gate204inter4), .b(gate204inter3), .O(gate204inter5));
  nor2  gate1379(.a(gate204inter5), .b(gate204inter2), .O(gate204inter6));
  inv1  gate1380(.a(G607), .O(gate204inter7));
  inv1  gate1381(.a(G617), .O(gate204inter8));
  nand2 gate1382(.a(gate204inter8), .b(gate204inter7), .O(gate204inter9));
  nand2 gate1383(.a(s_119), .b(gate204inter3), .O(gate204inter10));
  nor2  gate1384(.a(gate204inter10), .b(gate204inter9), .O(gate204inter11));
  nor2  gate1385(.a(gate204inter11), .b(gate204inter6), .O(gate204inter12));
  nand2 gate1386(.a(gate204inter12), .b(gate204inter1), .O(G675));
nand2 gate205( .a(G622), .b(G627), .O(G678) );
nand2 gate206( .a(G632), .b(G637), .O(G681) );
nand2 gate207( .a(G622), .b(G632), .O(G684) );
nand2 gate208( .a(G627), .b(G637), .O(G687) );
nand2 gate209( .a(G602), .b(G666), .O(G690) );
nand2 gate210( .a(G607), .b(G666), .O(G691) );
nand2 gate211( .a(G612), .b(G669), .O(G692) );
nand2 gate212( .a(G617), .b(G669), .O(G693) );
nand2 gate213( .a(G602), .b(G672), .O(G694) );
nand2 gate214( .a(G612), .b(G672), .O(G695) );

  xor2  gate589(.a(G675), .b(G607), .O(gate215inter0));
  nand2 gate590(.a(gate215inter0), .b(s_6), .O(gate215inter1));
  and2  gate591(.a(G675), .b(G607), .O(gate215inter2));
  inv1  gate592(.a(s_6), .O(gate215inter3));
  inv1  gate593(.a(s_7), .O(gate215inter4));
  nand2 gate594(.a(gate215inter4), .b(gate215inter3), .O(gate215inter5));
  nor2  gate595(.a(gate215inter5), .b(gate215inter2), .O(gate215inter6));
  inv1  gate596(.a(G607), .O(gate215inter7));
  inv1  gate597(.a(G675), .O(gate215inter8));
  nand2 gate598(.a(gate215inter8), .b(gate215inter7), .O(gate215inter9));
  nand2 gate599(.a(s_7), .b(gate215inter3), .O(gate215inter10));
  nor2  gate600(.a(gate215inter10), .b(gate215inter9), .O(gate215inter11));
  nor2  gate601(.a(gate215inter11), .b(gate215inter6), .O(gate215inter12));
  nand2 gate602(.a(gate215inter12), .b(gate215inter1), .O(G696));
nand2 gate216( .a(G617), .b(G675), .O(G697) );
nand2 gate217( .a(G622), .b(G678), .O(G698) );
nand2 gate218( .a(G627), .b(G678), .O(G699) );
nand2 gate219( .a(G632), .b(G681), .O(G700) );
nand2 gate220( .a(G637), .b(G681), .O(G701) );
nand2 gate221( .a(G622), .b(G684), .O(G702) );
nand2 gate222( .a(G632), .b(G684), .O(G703) );
nand2 gate223( .a(G627), .b(G687), .O(G704) );
nand2 gate224( .a(G637), .b(G687), .O(G705) );
nand2 gate225( .a(G690), .b(G691), .O(G706) );
nand2 gate226( .a(G692), .b(G693), .O(G709) );
nand2 gate227( .a(G694), .b(G695), .O(G712) );
nand2 gate228( .a(G696), .b(G697), .O(G715) );
nand2 gate229( .a(G698), .b(G699), .O(G718) );
nand2 gate230( .a(G700), .b(G701), .O(G721) );
nand2 gate231( .a(G702), .b(G703), .O(G724) );
nand2 gate232( .a(G704), .b(G705), .O(G727) );
nand2 gate233( .a(G242), .b(G718), .O(G730) );
nand2 gate234( .a(G245), .b(G721), .O(G733) );
nand2 gate235( .a(G248), .b(G724), .O(G736) );

  xor2  gate631(.a(G727), .b(G251), .O(gate236inter0));
  nand2 gate632(.a(gate236inter0), .b(s_12), .O(gate236inter1));
  and2  gate633(.a(G727), .b(G251), .O(gate236inter2));
  inv1  gate634(.a(s_12), .O(gate236inter3));
  inv1  gate635(.a(s_13), .O(gate236inter4));
  nand2 gate636(.a(gate236inter4), .b(gate236inter3), .O(gate236inter5));
  nor2  gate637(.a(gate236inter5), .b(gate236inter2), .O(gate236inter6));
  inv1  gate638(.a(G251), .O(gate236inter7));
  inv1  gate639(.a(G727), .O(gate236inter8));
  nand2 gate640(.a(gate236inter8), .b(gate236inter7), .O(gate236inter9));
  nand2 gate641(.a(s_13), .b(gate236inter3), .O(gate236inter10));
  nor2  gate642(.a(gate236inter10), .b(gate236inter9), .O(gate236inter11));
  nor2  gate643(.a(gate236inter11), .b(gate236inter6), .O(gate236inter12));
  nand2 gate644(.a(gate236inter12), .b(gate236inter1), .O(G739));
nand2 gate237( .a(G254), .b(G706), .O(G742) );
nand2 gate238( .a(G257), .b(G709), .O(G745) );
nand2 gate239( .a(G260), .b(G712), .O(G748) );
nand2 gate240( .a(G263), .b(G715), .O(G751) );
nand2 gate241( .a(G242), .b(G730), .O(G754) );

  xor2  gate1205(.a(G730), .b(G718), .O(gate242inter0));
  nand2 gate1206(.a(gate242inter0), .b(s_94), .O(gate242inter1));
  and2  gate1207(.a(G730), .b(G718), .O(gate242inter2));
  inv1  gate1208(.a(s_94), .O(gate242inter3));
  inv1  gate1209(.a(s_95), .O(gate242inter4));
  nand2 gate1210(.a(gate242inter4), .b(gate242inter3), .O(gate242inter5));
  nor2  gate1211(.a(gate242inter5), .b(gate242inter2), .O(gate242inter6));
  inv1  gate1212(.a(G718), .O(gate242inter7));
  inv1  gate1213(.a(G730), .O(gate242inter8));
  nand2 gate1214(.a(gate242inter8), .b(gate242inter7), .O(gate242inter9));
  nand2 gate1215(.a(s_95), .b(gate242inter3), .O(gate242inter10));
  nor2  gate1216(.a(gate242inter10), .b(gate242inter9), .O(gate242inter11));
  nor2  gate1217(.a(gate242inter11), .b(gate242inter6), .O(gate242inter12));
  nand2 gate1218(.a(gate242inter12), .b(gate242inter1), .O(G755));
nand2 gate243( .a(G245), .b(G733), .O(G756) );
nand2 gate244( .a(G721), .b(G733), .O(G757) );
nand2 gate245( .a(G248), .b(G736), .O(G758) );
nand2 gate246( .a(G724), .b(G736), .O(G759) );
nand2 gate247( .a(G251), .b(G739), .O(G760) );
nand2 gate248( .a(G727), .b(G739), .O(G761) );
nand2 gate249( .a(G254), .b(G742), .O(G762) );

  xor2  gate743(.a(G742), .b(G706), .O(gate250inter0));
  nand2 gate744(.a(gate250inter0), .b(s_28), .O(gate250inter1));
  and2  gate745(.a(G742), .b(G706), .O(gate250inter2));
  inv1  gate746(.a(s_28), .O(gate250inter3));
  inv1  gate747(.a(s_29), .O(gate250inter4));
  nand2 gate748(.a(gate250inter4), .b(gate250inter3), .O(gate250inter5));
  nor2  gate749(.a(gate250inter5), .b(gate250inter2), .O(gate250inter6));
  inv1  gate750(.a(G706), .O(gate250inter7));
  inv1  gate751(.a(G742), .O(gate250inter8));
  nand2 gate752(.a(gate250inter8), .b(gate250inter7), .O(gate250inter9));
  nand2 gate753(.a(s_29), .b(gate250inter3), .O(gate250inter10));
  nor2  gate754(.a(gate250inter10), .b(gate250inter9), .O(gate250inter11));
  nor2  gate755(.a(gate250inter11), .b(gate250inter6), .O(gate250inter12));
  nand2 gate756(.a(gate250inter12), .b(gate250inter1), .O(G763));
nand2 gate251( .a(G257), .b(G745), .O(G764) );
nand2 gate252( .a(G709), .b(G745), .O(G765) );
nand2 gate253( .a(G260), .b(G748), .O(G766) );

  xor2  gate925(.a(G748), .b(G712), .O(gate254inter0));
  nand2 gate926(.a(gate254inter0), .b(s_54), .O(gate254inter1));
  and2  gate927(.a(G748), .b(G712), .O(gate254inter2));
  inv1  gate928(.a(s_54), .O(gate254inter3));
  inv1  gate929(.a(s_55), .O(gate254inter4));
  nand2 gate930(.a(gate254inter4), .b(gate254inter3), .O(gate254inter5));
  nor2  gate931(.a(gate254inter5), .b(gate254inter2), .O(gate254inter6));
  inv1  gate932(.a(G712), .O(gate254inter7));
  inv1  gate933(.a(G748), .O(gate254inter8));
  nand2 gate934(.a(gate254inter8), .b(gate254inter7), .O(gate254inter9));
  nand2 gate935(.a(s_55), .b(gate254inter3), .O(gate254inter10));
  nor2  gate936(.a(gate254inter10), .b(gate254inter9), .O(gate254inter11));
  nor2  gate937(.a(gate254inter11), .b(gate254inter6), .O(gate254inter12));
  nand2 gate938(.a(gate254inter12), .b(gate254inter1), .O(G767));
nand2 gate255( .a(G263), .b(G751), .O(G768) );

  xor2  gate1107(.a(G751), .b(G715), .O(gate256inter0));
  nand2 gate1108(.a(gate256inter0), .b(s_80), .O(gate256inter1));
  and2  gate1109(.a(G751), .b(G715), .O(gate256inter2));
  inv1  gate1110(.a(s_80), .O(gate256inter3));
  inv1  gate1111(.a(s_81), .O(gate256inter4));
  nand2 gate1112(.a(gate256inter4), .b(gate256inter3), .O(gate256inter5));
  nor2  gate1113(.a(gate256inter5), .b(gate256inter2), .O(gate256inter6));
  inv1  gate1114(.a(G715), .O(gate256inter7));
  inv1  gate1115(.a(G751), .O(gate256inter8));
  nand2 gate1116(.a(gate256inter8), .b(gate256inter7), .O(gate256inter9));
  nand2 gate1117(.a(s_81), .b(gate256inter3), .O(gate256inter10));
  nor2  gate1118(.a(gate256inter10), .b(gate256inter9), .O(gate256inter11));
  nor2  gate1119(.a(gate256inter11), .b(gate256inter6), .O(gate256inter12));
  nand2 gate1120(.a(gate256inter12), .b(gate256inter1), .O(G769));
nand2 gate257( .a(G754), .b(G755), .O(G770) );
nand2 gate258( .a(G756), .b(G757), .O(G773) );
nand2 gate259( .a(G758), .b(G759), .O(G776) );
nand2 gate260( .a(G760), .b(G761), .O(G779) );
nand2 gate261( .a(G762), .b(G763), .O(G782) );
nand2 gate262( .a(G764), .b(G765), .O(G785) );
nand2 gate263( .a(G766), .b(G767), .O(G788) );
nand2 gate264( .a(G768), .b(G769), .O(G791) );
nand2 gate265( .a(G642), .b(G770), .O(G794) );
nand2 gate266( .a(G645), .b(G773), .O(G797) );
nand2 gate267( .a(G648), .b(G776), .O(G800) );
nand2 gate268( .a(G651), .b(G779), .O(G803) );
nand2 gate269( .a(G654), .b(G782), .O(G806) );
nand2 gate270( .a(G657), .b(G785), .O(G809) );
nand2 gate271( .a(G660), .b(G788), .O(G812) );

  xor2  gate1401(.a(G791), .b(G663), .O(gate272inter0));
  nand2 gate1402(.a(gate272inter0), .b(s_122), .O(gate272inter1));
  and2  gate1403(.a(G791), .b(G663), .O(gate272inter2));
  inv1  gate1404(.a(s_122), .O(gate272inter3));
  inv1  gate1405(.a(s_123), .O(gate272inter4));
  nand2 gate1406(.a(gate272inter4), .b(gate272inter3), .O(gate272inter5));
  nor2  gate1407(.a(gate272inter5), .b(gate272inter2), .O(gate272inter6));
  inv1  gate1408(.a(G663), .O(gate272inter7));
  inv1  gate1409(.a(G791), .O(gate272inter8));
  nand2 gate1410(.a(gate272inter8), .b(gate272inter7), .O(gate272inter9));
  nand2 gate1411(.a(s_123), .b(gate272inter3), .O(gate272inter10));
  nor2  gate1412(.a(gate272inter10), .b(gate272inter9), .O(gate272inter11));
  nor2  gate1413(.a(gate272inter11), .b(gate272inter6), .O(gate272inter12));
  nand2 gate1414(.a(gate272inter12), .b(gate272inter1), .O(G815));
nand2 gate273( .a(G642), .b(G794), .O(G818) );
nand2 gate274( .a(G770), .b(G794), .O(G819) );
nand2 gate275( .a(G645), .b(G797), .O(G820) );
nand2 gate276( .a(G773), .b(G797), .O(G821) );

  xor2  gate561(.a(G800), .b(G648), .O(gate277inter0));
  nand2 gate562(.a(gate277inter0), .b(s_2), .O(gate277inter1));
  and2  gate563(.a(G800), .b(G648), .O(gate277inter2));
  inv1  gate564(.a(s_2), .O(gate277inter3));
  inv1  gate565(.a(s_3), .O(gate277inter4));
  nand2 gate566(.a(gate277inter4), .b(gate277inter3), .O(gate277inter5));
  nor2  gate567(.a(gate277inter5), .b(gate277inter2), .O(gate277inter6));
  inv1  gate568(.a(G648), .O(gate277inter7));
  inv1  gate569(.a(G800), .O(gate277inter8));
  nand2 gate570(.a(gate277inter8), .b(gate277inter7), .O(gate277inter9));
  nand2 gate571(.a(s_3), .b(gate277inter3), .O(gate277inter10));
  nor2  gate572(.a(gate277inter10), .b(gate277inter9), .O(gate277inter11));
  nor2  gate573(.a(gate277inter11), .b(gate277inter6), .O(gate277inter12));
  nand2 gate574(.a(gate277inter12), .b(gate277inter1), .O(G822));

  xor2  gate1275(.a(G800), .b(G776), .O(gate278inter0));
  nand2 gate1276(.a(gate278inter0), .b(s_104), .O(gate278inter1));
  and2  gate1277(.a(G800), .b(G776), .O(gate278inter2));
  inv1  gate1278(.a(s_104), .O(gate278inter3));
  inv1  gate1279(.a(s_105), .O(gate278inter4));
  nand2 gate1280(.a(gate278inter4), .b(gate278inter3), .O(gate278inter5));
  nor2  gate1281(.a(gate278inter5), .b(gate278inter2), .O(gate278inter6));
  inv1  gate1282(.a(G776), .O(gate278inter7));
  inv1  gate1283(.a(G800), .O(gate278inter8));
  nand2 gate1284(.a(gate278inter8), .b(gate278inter7), .O(gate278inter9));
  nand2 gate1285(.a(s_105), .b(gate278inter3), .O(gate278inter10));
  nor2  gate1286(.a(gate278inter10), .b(gate278inter9), .O(gate278inter11));
  nor2  gate1287(.a(gate278inter11), .b(gate278inter6), .O(gate278inter12));
  nand2 gate1288(.a(gate278inter12), .b(gate278inter1), .O(G823));
nand2 gate279( .a(G651), .b(G803), .O(G824) );
nand2 gate280( .a(G779), .b(G803), .O(G825) );
nand2 gate281( .a(G654), .b(G806), .O(G826) );

  xor2  gate1247(.a(G806), .b(G782), .O(gate282inter0));
  nand2 gate1248(.a(gate282inter0), .b(s_100), .O(gate282inter1));
  and2  gate1249(.a(G806), .b(G782), .O(gate282inter2));
  inv1  gate1250(.a(s_100), .O(gate282inter3));
  inv1  gate1251(.a(s_101), .O(gate282inter4));
  nand2 gate1252(.a(gate282inter4), .b(gate282inter3), .O(gate282inter5));
  nor2  gate1253(.a(gate282inter5), .b(gate282inter2), .O(gate282inter6));
  inv1  gate1254(.a(G782), .O(gate282inter7));
  inv1  gate1255(.a(G806), .O(gate282inter8));
  nand2 gate1256(.a(gate282inter8), .b(gate282inter7), .O(gate282inter9));
  nand2 gate1257(.a(s_101), .b(gate282inter3), .O(gate282inter10));
  nor2  gate1258(.a(gate282inter10), .b(gate282inter9), .O(gate282inter11));
  nor2  gate1259(.a(gate282inter11), .b(gate282inter6), .O(gate282inter12));
  nand2 gate1260(.a(gate282inter12), .b(gate282inter1), .O(G827));
nand2 gate283( .a(G657), .b(G809), .O(G828) );
nand2 gate284( .a(G785), .b(G809), .O(G829) );
nand2 gate285( .a(G660), .b(G812), .O(G830) );
nand2 gate286( .a(G788), .b(G812), .O(G831) );

  xor2  gate785(.a(G815), .b(G663), .O(gate287inter0));
  nand2 gate786(.a(gate287inter0), .b(s_34), .O(gate287inter1));
  and2  gate787(.a(G815), .b(G663), .O(gate287inter2));
  inv1  gate788(.a(s_34), .O(gate287inter3));
  inv1  gate789(.a(s_35), .O(gate287inter4));
  nand2 gate790(.a(gate287inter4), .b(gate287inter3), .O(gate287inter5));
  nor2  gate791(.a(gate287inter5), .b(gate287inter2), .O(gate287inter6));
  inv1  gate792(.a(G663), .O(gate287inter7));
  inv1  gate793(.a(G815), .O(gate287inter8));
  nand2 gate794(.a(gate287inter8), .b(gate287inter7), .O(gate287inter9));
  nand2 gate795(.a(s_35), .b(gate287inter3), .O(gate287inter10));
  nor2  gate796(.a(gate287inter10), .b(gate287inter9), .O(gate287inter11));
  nor2  gate797(.a(gate287inter11), .b(gate287inter6), .O(gate287inter12));
  nand2 gate798(.a(gate287inter12), .b(gate287inter1), .O(G832));
nand2 gate288( .a(G791), .b(G815), .O(G833) );

  xor2  gate729(.a(G819), .b(G818), .O(gate289inter0));
  nand2 gate730(.a(gate289inter0), .b(s_26), .O(gate289inter1));
  and2  gate731(.a(G819), .b(G818), .O(gate289inter2));
  inv1  gate732(.a(s_26), .O(gate289inter3));
  inv1  gate733(.a(s_27), .O(gate289inter4));
  nand2 gate734(.a(gate289inter4), .b(gate289inter3), .O(gate289inter5));
  nor2  gate735(.a(gate289inter5), .b(gate289inter2), .O(gate289inter6));
  inv1  gate736(.a(G818), .O(gate289inter7));
  inv1  gate737(.a(G819), .O(gate289inter8));
  nand2 gate738(.a(gate289inter8), .b(gate289inter7), .O(gate289inter9));
  nand2 gate739(.a(s_27), .b(gate289inter3), .O(gate289inter10));
  nor2  gate740(.a(gate289inter10), .b(gate289inter9), .O(gate289inter11));
  nor2  gate741(.a(gate289inter11), .b(gate289inter6), .O(gate289inter12));
  nand2 gate742(.a(gate289inter12), .b(gate289inter1), .O(G834));
nand2 gate290( .a(G820), .b(G821), .O(G847) );

  xor2  gate645(.a(G823), .b(G822), .O(gate291inter0));
  nand2 gate646(.a(gate291inter0), .b(s_14), .O(gate291inter1));
  and2  gate647(.a(G823), .b(G822), .O(gate291inter2));
  inv1  gate648(.a(s_14), .O(gate291inter3));
  inv1  gate649(.a(s_15), .O(gate291inter4));
  nand2 gate650(.a(gate291inter4), .b(gate291inter3), .O(gate291inter5));
  nor2  gate651(.a(gate291inter5), .b(gate291inter2), .O(gate291inter6));
  inv1  gate652(.a(G822), .O(gate291inter7));
  inv1  gate653(.a(G823), .O(gate291inter8));
  nand2 gate654(.a(gate291inter8), .b(gate291inter7), .O(gate291inter9));
  nand2 gate655(.a(s_15), .b(gate291inter3), .O(gate291inter10));
  nor2  gate656(.a(gate291inter10), .b(gate291inter9), .O(gate291inter11));
  nor2  gate657(.a(gate291inter11), .b(gate291inter6), .O(gate291inter12));
  nand2 gate658(.a(gate291inter12), .b(gate291inter1), .O(G860));
nand2 gate292( .a(G824), .b(G825), .O(G873) );
nand2 gate293( .a(G828), .b(G829), .O(G886) );
nand2 gate294( .a(G832), .b(G833), .O(G899) );
nand2 gate295( .a(G830), .b(G831), .O(G912) );
nand2 gate296( .a(G826), .b(G827), .O(G925) );
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );
nand2 gate387( .a(G1), .b(G1036), .O(G1132) );
nand2 gate388( .a(G2), .b(G1039), .O(G1135) );
nand2 gate389( .a(G3), .b(G1042), .O(G1138) );

  xor2  gate911(.a(G1045), .b(G4), .O(gate390inter0));
  nand2 gate912(.a(gate390inter0), .b(s_52), .O(gate390inter1));
  and2  gate913(.a(G1045), .b(G4), .O(gate390inter2));
  inv1  gate914(.a(s_52), .O(gate390inter3));
  inv1  gate915(.a(s_53), .O(gate390inter4));
  nand2 gate916(.a(gate390inter4), .b(gate390inter3), .O(gate390inter5));
  nor2  gate917(.a(gate390inter5), .b(gate390inter2), .O(gate390inter6));
  inv1  gate918(.a(G4), .O(gate390inter7));
  inv1  gate919(.a(G1045), .O(gate390inter8));
  nand2 gate920(.a(gate390inter8), .b(gate390inter7), .O(gate390inter9));
  nand2 gate921(.a(s_53), .b(gate390inter3), .O(gate390inter10));
  nor2  gate922(.a(gate390inter10), .b(gate390inter9), .O(gate390inter11));
  nor2  gate923(.a(gate390inter11), .b(gate390inter6), .O(gate390inter12));
  nand2 gate924(.a(gate390inter12), .b(gate390inter1), .O(G1141));
nand2 gate391( .a(G5), .b(G1048), .O(G1144) );
nand2 gate392( .a(G6), .b(G1051), .O(G1147) );

  xor2  gate1331(.a(G1054), .b(G7), .O(gate393inter0));
  nand2 gate1332(.a(gate393inter0), .b(s_112), .O(gate393inter1));
  and2  gate1333(.a(G1054), .b(G7), .O(gate393inter2));
  inv1  gate1334(.a(s_112), .O(gate393inter3));
  inv1  gate1335(.a(s_113), .O(gate393inter4));
  nand2 gate1336(.a(gate393inter4), .b(gate393inter3), .O(gate393inter5));
  nor2  gate1337(.a(gate393inter5), .b(gate393inter2), .O(gate393inter6));
  inv1  gate1338(.a(G7), .O(gate393inter7));
  inv1  gate1339(.a(G1054), .O(gate393inter8));
  nand2 gate1340(.a(gate393inter8), .b(gate393inter7), .O(gate393inter9));
  nand2 gate1341(.a(s_113), .b(gate393inter3), .O(gate393inter10));
  nor2  gate1342(.a(gate393inter10), .b(gate393inter9), .O(gate393inter11));
  nor2  gate1343(.a(gate393inter11), .b(gate393inter6), .O(gate393inter12));
  nand2 gate1344(.a(gate393inter12), .b(gate393inter1), .O(G1150));
nand2 gate394( .a(G8), .b(G1057), .O(G1153) );
nand2 gate395( .a(G9), .b(G1060), .O(G1156) );
nand2 gate396( .a(G10), .b(G1063), .O(G1159) );
nand2 gate397( .a(G11), .b(G1066), .O(G1162) );
nand2 gate398( .a(G12), .b(G1069), .O(G1165) );
nand2 gate399( .a(G13), .b(G1072), .O(G1168) );
nand2 gate400( .a(G14), .b(G1075), .O(G1171) );
nand2 gate401( .a(G15), .b(G1078), .O(G1174) );
nand2 gate402( .a(G16), .b(G1081), .O(G1177) );

  xor2  gate1261(.a(G1084), .b(G17), .O(gate403inter0));
  nand2 gate1262(.a(gate403inter0), .b(s_102), .O(gate403inter1));
  and2  gate1263(.a(G1084), .b(G17), .O(gate403inter2));
  inv1  gate1264(.a(s_102), .O(gate403inter3));
  inv1  gate1265(.a(s_103), .O(gate403inter4));
  nand2 gate1266(.a(gate403inter4), .b(gate403inter3), .O(gate403inter5));
  nor2  gate1267(.a(gate403inter5), .b(gate403inter2), .O(gate403inter6));
  inv1  gate1268(.a(G17), .O(gate403inter7));
  inv1  gate1269(.a(G1084), .O(gate403inter8));
  nand2 gate1270(.a(gate403inter8), .b(gate403inter7), .O(gate403inter9));
  nand2 gate1271(.a(s_103), .b(gate403inter3), .O(gate403inter10));
  nor2  gate1272(.a(gate403inter10), .b(gate403inter9), .O(gate403inter11));
  nor2  gate1273(.a(gate403inter11), .b(gate403inter6), .O(gate403inter12));
  nand2 gate1274(.a(gate403inter12), .b(gate403inter1), .O(G1180));
nand2 gate404( .a(G18), .b(G1087), .O(G1183) );
nand2 gate405( .a(G19), .b(G1090), .O(G1186) );
nand2 gate406( .a(G20), .b(G1093), .O(G1189) );

  xor2  gate827(.a(G1096), .b(G21), .O(gate407inter0));
  nand2 gate828(.a(gate407inter0), .b(s_40), .O(gate407inter1));
  and2  gate829(.a(G1096), .b(G21), .O(gate407inter2));
  inv1  gate830(.a(s_40), .O(gate407inter3));
  inv1  gate831(.a(s_41), .O(gate407inter4));
  nand2 gate832(.a(gate407inter4), .b(gate407inter3), .O(gate407inter5));
  nor2  gate833(.a(gate407inter5), .b(gate407inter2), .O(gate407inter6));
  inv1  gate834(.a(G21), .O(gate407inter7));
  inv1  gate835(.a(G1096), .O(gate407inter8));
  nand2 gate836(.a(gate407inter8), .b(gate407inter7), .O(gate407inter9));
  nand2 gate837(.a(s_41), .b(gate407inter3), .O(gate407inter10));
  nor2  gate838(.a(gate407inter10), .b(gate407inter9), .O(gate407inter11));
  nor2  gate839(.a(gate407inter11), .b(gate407inter6), .O(gate407inter12));
  nand2 gate840(.a(gate407inter12), .b(gate407inter1), .O(G1192));
nand2 gate408( .a(G22), .b(G1099), .O(G1195) );
nand2 gate409( .a(G23), .b(G1102), .O(G1198) );
nand2 gate410( .a(G24), .b(G1105), .O(G1201) );
nand2 gate411( .a(G25), .b(G1108), .O(G1204) );
nand2 gate412( .a(G26), .b(G1111), .O(G1207) );
nand2 gate413( .a(G27), .b(G1114), .O(G1210) );
nand2 gate414( .a(G28), .b(G1117), .O(G1213) );

  xor2  gate757(.a(G1120), .b(G29), .O(gate415inter0));
  nand2 gate758(.a(gate415inter0), .b(s_30), .O(gate415inter1));
  and2  gate759(.a(G1120), .b(G29), .O(gate415inter2));
  inv1  gate760(.a(s_30), .O(gate415inter3));
  inv1  gate761(.a(s_31), .O(gate415inter4));
  nand2 gate762(.a(gate415inter4), .b(gate415inter3), .O(gate415inter5));
  nor2  gate763(.a(gate415inter5), .b(gate415inter2), .O(gate415inter6));
  inv1  gate764(.a(G29), .O(gate415inter7));
  inv1  gate765(.a(G1120), .O(gate415inter8));
  nand2 gate766(.a(gate415inter8), .b(gate415inter7), .O(gate415inter9));
  nand2 gate767(.a(s_31), .b(gate415inter3), .O(gate415inter10));
  nor2  gate768(.a(gate415inter10), .b(gate415inter9), .O(gate415inter11));
  nor2  gate769(.a(gate415inter11), .b(gate415inter6), .O(gate415inter12));
  nand2 gate770(.a(gate415inter12), .b(gate415inter1), .O(G1216));
nand2 gate416( .a(G30), .b(G1123), .O(G1219) );

  xor2  gate617(.a(G1126), .b(G31), .O(gate417inter0));
  nand2 gate618(.a(gate417inter0), .b(s_10), .O(gate417inter1));
  and2  gate619(.a(G1126), .b(G31), .O(gate417inter2));
  inv1  gate620(.a(s_10), .O(gate417inter3));
  inv1  gate621(.a(s_11), .O(gate417inter4));
  nand2 gate622(.a(gate417inter4), .b(gate417inter3), .O(gate417inter5));
  nor2  gate623(.a(gate417inter5), .b(gate417inter2), .O(gate417inter6));
  inv1  gate624(.a(G31), .O(gate417inter7));
  inv1  gate625(.a(G1126), .O(gate417inter8));
  nand2 gate626(.a(gate417inter8), .b(gate417inter7), .O(gate417inter9));
  nand2 gate627(.a(s_11), .b(gate417inter3), .O(gate417inter10));
  nor2  gate628(.a(gate417inter10), .b(gate417inter9), .O(gate417inter11));
  nor2  gate629(.a(gate417inter11), .b(gate417inter6), .O(gate417inter12));
  nand2 gate630(.a(gate417inter12), .b(gate417inter1), .O(G1222));
nand2 gate418( .a(G32), .b(G1129), .O(G1225) );

  xor2  gate547(.a(G1132), .b(G1), .O(gate419inter0));
  nand2 gate548(.a(gate419inter0), .b(s_0), .O(gate419inter1));
  and2  gate549(.a(G1132), .b(G1), .O(gate419inter2));
  inv1  gate550(.a(s_0), .O(gate419inter3));
  inv1  gate551(.a(s_1), .O(gate419inter4));
  nand2 gate552(.a(gate419inter4), .b(gate419inter3), .O(gate419inter5));
  nor2  gate553(.a(gate419inter5), .b(gate419inter2), .O(gate419inter6));
  inv1  gate554(.a(G1), .O(gate419inter7));
  inv1  gate555(.a(G1132), .O(gate419inter8));
  nand2 gate556(.a(gate419inter8), .b(gate419inter7), .O(gate419inter9));
  nand2 gate557(.a(s_1), .b(gate419inter3), .O(gate419inter10));
  nor2  gate558(.a(gate419inter10), .b(gate419inter9), .O(gate419inter11));
  nor2  gate559(.a(gate419inter11), .b(gate419inter6), .O(gate419inter12));
  nand2 gate560(.a(gate419inter12), .b(gate419inter1), .O(G1228));
nand2 gate420( .a(G1036), .b(G1132), .O(G1229) );
nand2 gate421( .a(G2), .b(G1135), .O(G1230) );
nand2 gate422( .a(G1039), .b(G1135), .O(G1231) );
nand2 gate423( .a(G3), .b(G1138), .O(G1232) );
nand2 gate424( .a(G1042), .b(G1138), .O(G1233) );
nand2 gate425( .a(G4), .b(G1141), .O(G1234) );
nand2 gate426( .a(G1045), .b(G1141), .O(G1235) );
nand2 gate427( .a(G5), .b(G1144), .O(G1236) );

  xor2  gate603(.a(G1144), .b(G1048), .O(gate428inter0));
  nand2 gate604(.a(gate428inter0), .b(s_8), .O(gate428inter1));
  and2  gate605(.a(G1144), .b(G1048), .O(gate428inter2));
  inv1  gate606(.a(s_8), .O(gate428inter3));
  inv1  gate607(.a(s_9), .O(gate428inter4));
  nand2 gate608(.a(gate428inter4), .b(gate428inter3), .O(gate428inter5));
  nor2  gate609(.a(gate428inter5), .b(gate428inter2), .O(gate428inter6));
  inv1  gate610(.a(G1048), .O(gate428inter7));
  inv1  gate611(.a(G1144), .O(gate428inter8));
  nand2 gate612(.a(gate428inter8), .b(gate428inter7), .O(gate428inter9));
  nand2 gate613(.a(s_9), .b(gate428inter3), .O(gate428inter10));
  nor2  gate614(.a(gate428inter10), .b(gate428inter9), .O(gate428inter11));
  nor2  gate615(.a(gate428inter11), .b(gate428inter6), .O(gate428inter12));
  nand2 gate616(.a(gate428inter12), .b(gate428inter1), .O(G1237));
nand2 gate429( .a(G6), .b(G1147), .O(G1238) );
nand2 gate430( .a(G1051), .b(G1147), .O(G1239) );
nand2 gate431( .a(G7), .b(G1150), .O(G1240) );

  xor2  gate1233(.a(G1150), .b(G1054), .O(gate432inter0));
  nand2 gate1234(.a(gate432inter0), .b(s_98), .O(gate432inter1));
  and2  gate1235(.a(G1150), .b(G1054), .O(gate432inter2));
  inv1  gate1236(.a(s_98), .O(gate432inter3));
  inv1  gate1237(.a(s_99), .O(gate432inter4));
  nand2 gate1238(.a(gate432inter4), .b(gate432inter3), .O(gate432inter5));
  nor2  gate1239(.a(gate432inter5), .b(gate432inter2), .O(gate432inter6));
  inv1  gate1240(.a(G1054), .O(gate432inter7));
  inv1  gate1241(.a(G1150), .O(gate432inter8));
  nand2 gate1242(.a(gate432inter8), .b(gate432inter7), .O(gate432inter9));
  nand2 gate1243(.a(s_99), .b(gate432inter3), .O(gate432inter10));
  nor2  gate1244(.a(gate432inter10), .b(gate432inter9), .O(gate432inter11));
  nor2  gate1245(.a(gate432inter11), .b(gate432inter6), .O(gate432inter12));
  nand2 gate1246(.a(gate432inter12), .b(gate432inter1), .O(G1241));
nand2 gate433( .a(G8), .b(G1153), .O(G1242) );
nand2 gate434( .a(G1057), .b(G1153), .O(G1243) );
nand2 gate435( .a(G9), .b(G1156), .O(G1244) );
nand2 gate436( .a(G1060), .b(G1156), .O(G1245) );
nand2 gate437( .a(G10), .b(G1159), .O(G1246) );
nand2 gate438( .a(G1063), .b(G1159), .O(G1247) );
nand2 gate439( .a(G11), .b(G1162), .O(G1248) );
nand2 gate440( .a(G1066), .b(G1162), .O(G1249) );
nand2 gate441( .a(G12), .b(G1165), .O(G1250) );
nand2 gate442( .a(G1069), .b(G1165), .O(G1251) );
nand2 gate443( .a(G13), .b(G1168), .O(G1252) );

  xor2  gate1009(.a(G1168), .b(G1072), .O(gate444inter0));
  nand2 gate1010(.a(gate444inter0), .b(s_66), .O(gate444inter1));
  and2  gate1011(.a(G1168), .b(G1072), .O(gate444inter2));
  inv1  gate1012(.a(s_66), .O(gate444inter3));
  inv1  gate1013(.a(s_67), .O(gate444inter4));
  nand2 gate1014(.a(gate444inter4), .b(gate444inter3), .O(gate444inter5));
  nor2  gate1015(.a(gate444inter5), .b(gate444inter2), .O(gate444inter6));
  inv1  gate1016(.a(G1072), .O(gate444inter7));
  inv1  gate1017(.a(G1168), .O(gate444inter8));
  nand2 gate1018(.a(gate444inter8), .b(gate444inter7), .O(gate444inter9));
  nand2 gate1019(.a(s_67), .b(gate444inter3), .O(gate444inter10));
  nor2  gate1020(.a(gate444inter10), .b(gate444inter9), .O(gate444inter11));
  nor2  gate1021(.a(gate444inter11), .b(gate444inter6), .O(gate444inter12));
  nand2 gate1022(.a(gate444inter12), .b(gate444inter1), .O(G1253));

  xor2  gate855(.a(G1171), .b(G14), .O(gate445inter0));
  nand2 gate856(.a(gate445inter0), .b(s_44), .O(gate445inter1));
  and2  gate857(.a(G1171), .b(G14), .O(gate445inter2));
  inv1  gate858(.a(s_44), .O(gate445inter3));
  inv1  gate859(.a(s_45), .O(gate445inter4));
  nand2 gate860(.a(gate445inter4), .b(gate445inter3), .O(gate445inter5));
  nor2  gate861(.a(gate445inter5), .b(gate445inter2), .O(gate445inter6));
  inv1  gate862(.a(G14), .O(gate445inter7));
  inv1  gate863(.a(G1171), .O(gate445inter8));
  nand2 gate864(.a(gate445inter8), .b(gate445inter7), .O(gate445inter9));
  nand2 gate865(.a(s_45), .b(gate445inter3), .O(gate445inter10));
  nor2  gate866(.a(gate445inter10), .b(gate445inter9), .O(gate445inter11));
  nor2  gate867(.a(gate445inter11), .b(gate445inter6), .O(gate445inter12));
  nand2 gate868(.a(gate445inter12), .b(gate445inter1), .O(G1254));
nand2 gate446( .a(G1075), .b(G1171), .O(G1255) );
nand2 gate447( .a(G15), .b(G1174), .O(G1256) );

  xor2  gate1037(.a(G1174), .b(G1078), .O(gate448inter0));
  nand2 gate1038(.a(gate448inter0), .b(s_70), .O(gate448inter1));
  and2  gate1039(.a(G1174), .b(G1078), .O(gate448inter2));
  inv1  gate1040(.a(s_70), .O(gate448inter3));
  inv1  gate1041(.a(s_71), .O(gate448inter4));
  nand2 gate1042(.a(gate448inter4), .b(gate448inter3), .O(gate448inter5));
  nor2  gate1043(.a(gate448inter5), .b(gate448inter2), .O(gate448inter6));
  inv1  gate1044(.a(G1078), .O(gate448inter7));
  inv1  gate1045(.a(G1174), .O(gate448inter8));
  nand2 gate1046(.a(gate448inter8), .b(gate448inter7), .O(gate448inter9));
  nand2 gate1047(.a(s_71), .b(gate448inter3), .O(gate448inter10));
  nor2  gate1048(.a(gate448inter10), .b(gate448inter9), .O(gate448inter11));
  nor2  gate1049(.a(gate448inter11), .b(gate448inter6), .O(gate448inter12));
  nand2 gate1050(.a(gate448inter12), .b(gate448inter1), .O(G1257));

  xor2  gate813(.a(G1177), .b(G16), .O(gate449inter0));
  nand2 gate814(.a(gate449inter0), .b(s_38), .O(gate449inter1));
  and2  gate815(.a(G1177), .b(G16), .O(gate449inter2));
  inv1  gate816(.a(s_38), .O(gate449inter3));
  inv1  gate817(.a(s_39), .O(gate449inter4));
  nand2 gate818(.a(gate449inter4), .b(gate449inter3), .O(gate449inter5));
  nor2  gate819(.a(gate449inter5), .b(gate449inter2), .O(gate449inter6));
  inv1  gate820(.a(G16), .O(gate449inter7));
  inv1  gate821(.a(G1177), .O(gate449inter8));
  nand2 gate822(.a(gate449inter8), .b(gate449inter7), .O(gate449inter9));
  nand2 gate823(.a(s_39), .b(gate449inter3), .O(gate449inter10));
  nor2  gate824(.a(gate449inter10), .b(gate449inter9), .O(gate449inter11));
  nor2  gate825(.a(gate449inter11), .b(gate449inter6), .O(gate449inter12));
  nand2 gate826(.a(gate449inter12), .b(gate449inter1), .O(G1258));
nand2 gate450( .a(G1081), .b(G1177), .O(G1259) );
nand2 gate451( .a(G17), .b(G1180), .O(G1260) );
nand2 gate452( .a(G1084), .b(G1180), .O(G1261) );
nand2 gate453( .a(G18), .b(G1183), .O(G1262) );
nand2 gate454( .a(G1087), .b(G1183), .O(G1263) );
nand2 gate455( .a(G19), .b(G1186), .O(G1264) );
nand2 gate456( .a(G1090), .b(G1186), .O(G1265) );

  xor2  gate939(.a(G1189), .b(G20), .O(gate457inter0));
  nand2 gate940(.a(gate457inter0), .b(s_56), .O(gate457inter1));
  and2  gate941(.a(G1189), .b(G20), .O(gate457inter2));
  inv1  gate942(.a(s_56), .O(gate457inter3));
  inv1  gate943(.a(s_57), .O(gate457inter4));
  nand2 gate944(.a(gate457inter4), .b(gate457inter3), .O(gate457inter5));
  nor2  gate945(.a(gate457inter5), .b(gate457inter2), .O(gate457inter6));
  inv1  gate946(.a(G20), .O(gate457inter7));
  inv1  gate947(.a(G1189), .O(gate457inter8));
  nand2 gate948(.a(gate457inter8), .b(gate457inter7), .O(gate457inter9));
  nand2 gate949(.a(s_57), .b(gate457inter3), .O(gate457inter10));
  nor2  gate950(.a(gate457inter10), .b(gate457inter9), .O(gate457inter11));
  nor2  gate951(.a(gate457inter11), .b(gate457inter6), .O(gate457inter12));
  nand2 gate952(.a(gate457inter12), .b(gate457inter1), .O(G1266));

  xor2  gate967(.a(G1189), .b(G1093), .O(gate458inter0));
  nand2 gate968(.a(gate458inter0), .b(s_60), .O(gate458inter1));
  and2  gate969(.a(G1189), .b(G1093), .O(gate458inter2));
  inv1  gate970(.a(s_60), .O(gate458inter3));
  inv1  gate971(.a(s_61), .O(gate458inter4));
  nand2 gate972(.a(gate458inter4), .b(gate458inter3), .O(gate458inter5));
  nor2  gate973(.a(gate458inter5), .b(gate458inter2), .O(gate458inter6));
  inv1  gate974(.a(G1093), .O(gate458inter7));
  inv1  gate975(.a(G1189), .O(gate458inter8));
  nand2 gate976(.a(gate458inter8), .b(gate458inter7), .O(gate458inter9));
  nand2 gate977(.a(s_61), .b(gate458inter3), .O(gate458inter10));
  nor2  gate978(.a(gate458inter10), .b(gate458inter9), .O(gate458inter11));
  nor2  gate979(.a(gate458inter11), .b(gate458inter6), .O(gate458inter12));
  nand2 gate980(.a(gate458inter12), .b(gate458inter1), .O(G1267));
nand2 gate459( .a(G21), .b(G1192), .O(G1268) );

  xor2  gate995(.a(G1192), .b(G1096), .O(gate460inter0));
  nand2 gate996(.a(gate460inter0), .b(s_64), .O(gate460inter1));
  and2  gate997(.a(G1192), .b(G1096), .O(gate460inter2));
  inv1  gate998(.a(s_64), .O(gate460inter3));
  inv1  gate999(.a(s_65), .O(gate460inter4));
  nand2 gate1000(.a(gate460inter4), .b(gate460inter3), .O(gate460inter5));
  nor2  gate1001(.a(gate460inter5), .b(gate460inter2), .O(gate460inter6));
  inv1  gate1002(.a(G1096), .O(gate460inter7));
  inv1  gate1003(.a(G1192), .O(gate460inter8));
  nand2 gate1004(.a(gate460inter8), .b(gate460inter7), .O(gate460inter9));
  nand2 gate1005(.a(s_65), .b(gate460inter3), .O(gate460inter10));
  nor2  gate1006(.a(gate460inter10), .b(gate460inter9), .O(gate460inter11));
  nor2  gate1007(.a(gate460inter11), .b(gate460inter6), .O(gate460inter12));
  nand2 gate1008(.a(gate460inter12), .b(gate460inter1), .O(G1269));
nand2 gate461( .a(G22), .b(G1195), .O(G1270) );
nand2 gate462( .a(G1099), .b(G1195), .O(G1271) );
nand2 gate463( .a(G23), .b(G1198), .O(G1272) );
nand2 gate464( .a(G1102), .b(G1198), .O(G1273) );

  xor2  gate1051(.a(G1201), .b(G24), .O(gate465inter0));
  nand2 gate1052(.a(gate465inter0), .b(s_72), .O(gate465inter1));
  and2  gate1053(.a(G1201), .b(G24), .O(gate465inter2));
  inv1  gate1054(.a(s_72), .O(gate465inter3));
  inv1  gate1055(.a(s_73), .O(gate465inter4));
  nand2 gate1056(.a(gate465inter4), .b(gate465inter3), .O(gate465inter5));
  nor2  gate1057(.a(gate465inter5), .b(gate465inter2), .O(gate465inter6));
  inv1  gate1058(.a(G24), .O(gate465inter7));
  inv1  gate1059(.a(G1201), .O(gate465inter8));
  nand2 gate1060(.a(gate465inter8), .b(gate465inter7), .O(gate465inter9));
  nand2 gate1061(.a(s_73), .b(gate465inter3), .O(gate465inter10));
  nor2  gate1062(.a(gate465inter10), .b(gate465inter9), .O(gate465inter11));
  nor2  gate1063(.a(gate465inter11), .b(gate465inter6), .O(gate465inter12));
  nand2 gate1064(.a(gate465inter12), .b(gate465inter1), .O(G1274));
nand2 gate466( .a(G1105), .b(G1201), .O(G1275) );

  xor2  gate1163(.a(G1204), .b(G25), .O(gate467inter0));
  nand2 gate1164(.a(gate467inter0), .b(s_88), .O(gate467inter1));
  and2  gate1165(.a(G1204), .b(G25), .O(gate467inter2));
  inv1  gate1166(.a(s_88), .O(gate467inter3));
  inv1  gate1167(.a(s_89), .O(gate467inter4));
  nand2 gate1168(.a(gate467inter4), .b(gate467inter3), .O(gate467inter5));
  nor2  gate1169(.a(gate467inter5), .b(gate467inter2), .O(gate467inter6));
  inv1  gate1170(.a(G25), .O(gate467inter7));
  inv1  gate1171(.a(G1204), .O(gate467inter8));
  nand2 gate1172(.a(gate467inter8), .b(gate467inter7), .O(gate467inter9));
  nand2 gate1173(.a(s_89), .b(gate467inter3), .O(gate467inter10));
  nor2  gate1174(.a(gate467inter10), .b(gate467inter9), .O(gate467inter11));
  nor2  gate1175(.a(gate467inter11), .b(gate467inter6), .O(gate467inter12));
  nand2 gate1176(.a(gate467inter12), .b(gate467inter1), .O(G1276));
nand2 gate468( .a(G1108), .b(G1204), .O(G1277) );

  xor2  gate1219(.a(G1207), .b(G26), .O(gate469inter0));
  nand2 gate1220(.a(gate469inter0), .b(s_96), .O(gate469inter1));
  and2  gate1221(.a(G1207), .b(G26), .O(gate469inter2));
  inv1  gate1222(.a(s_96), .O(gate469inter3));
  inv1  gate1223(.a(s_97), .O(gate469inter4));
  nand2 gate1224(.a(gate469inter4), .b(gate469inter3), .O(gate469inter5));
  nor2  gate1225(.a(gate469inter5), .b(gate469inter2), .O(gate469inter6));
  inv1  gate1226(.a(G26), .O(gate469inter7));
  inv1  gate1227(.a(G1207), .O(gate469inter8));
  nand2 gate1228(.a(gate469inter8), .b(gate469inter7), .O(gate469inter9));
  nand2 gate1229(.a(s_97), .b(gate469inter3), .O(gate469inter10));
  nor2  gate1230(.a(gate469inter10), .b(gate469inter9), .O(gate469inter11));
  nor2  gate1231(.a(gate469inter11), .b(gate469inter6), .O(gate469inter12));
  nand2 gate1232(.a(gate469inter12), .b(gate469inter1), .O(G1278));
nand2 gate470( .a(G1111), .b(G1207), .O(G1279) );

  xor2  gate869(.a(G1210), .b(G27), .O(gate471inter0));
  nand2 gate870(.a(gate471inter0), .b(s_46), .O(gate471inter1));
  and2  gate871(.a(G1210), .b(G27), .O(gate471inter2));
  inv1  gate872(.a(s_46), .O(gate471inter3));
  inv1  gate873(.a(s_47), .O(gate471inter4));
  nand2 gate874(.a(gate471inter4), .b(gate471inter3), .O(gate471inter5));
  nor2  gate875(.a(gate471inter5), .b(gate471inter2), .O(gate471inter6));
  inv1  gate876(.a(G27), .O(gate471inter7));
  inv1  gate877(.a(G1210), .O(gate471inter8));
  nand2 gate878(.a(gate471inter8), .b(gate471inter7), .O(gate471inter9));
  nand2 gate879(.a(s_47), .b(gate471inter3), .O(gate471inter10));
  nor2  gate880(.a(gate471inter10), .b(gate471inter9), .O(gate471inter11));
  nor2  gate881(.a(gate471inter11), .b(gate471inter6), .O(gate471inter12));
  nand2 gate882(.a(gate471inter12), .b(gate471inter1), .O(G1280));
nand2 gate472( .a(G1114), .b(G1210), .O(G1281) );

  xor2  gate715(.a(G1213), .b(G28), .O(gate473inter0));
  nand2 gate716(.a(gate473inter0), .b(s_24), .O(gate473inter1));
  and2  gate717(.a(G1213), .b(G28), .O(gate473inter2));
  inv1  gate718(.a(s_24), .O(gate473inter3));
  inv1  gate719(.a(s_25), .O(gate473inter4));
  nand2 gate720(.a(gate473inter4), .b(gate473inter3), .O(gate473inter5));
  nor2  gate721(.a(gate473inter5), .b(gate473inter2), .O(gate473inter6));
  inv1  gate722(.a(G28), .O(gate473inter7));
  inv1  gate723(.a(G1213), .O(gate473inter8));
  nand2 gate724(.a(gate473inter8), .b(gate473inter7), .O(gate473inter9));
  nand2 gate725(.a(s_25), .b(gate473inter3), .O(gate473inter10));
  nor2  gate726(.a(gate473inter10), .b(gate473inter9), .O(gate473inter11));
  nor2  gate727(.a(gate473inter11), .b(gate473inter6), .O(gate473inter12));
  nand2 gate728(.a(gate473inter12), .b(gate473inter1), .O(G1282));
nand2 gate474( .a(G1117), .b(G1213), .O(G1283) );
nand2 gate475( .a(G29), .b(G1216), .O(G1284) );
nand2 gate476( .a(G1120), .b(G1216), .O(G1285) );
nand2 gate477( .a(G30), .b(G1219), .O(G1286) );
nand2 gate478( .a(G1123), .b(G1219), .O(G1287) );
nand2 gate479( .a(G31), .b(G1222), .O(G1288) );
nand2 gate480( .a(G1126), .b(G1222), .O(G1289) );
nand2 gate481( .a(G32), .b(G1225), .O(G1290) );
nand2 gate482( .a(G1129), .b(G1225), .O(G1291) );
nand2 gate483( .a(G1228), .b(G1229), .O(G1292) );
nand2 gate484( .a(G1230), .b(G1231), .O(G1293) );
nand2 gate485( .a(G1232), .b(G1233), .O(G1294) );
nand2 gate486( .a(G1234), .b(G1235), .O(G1295) );
nand2 gate487( .a(G1236), .b(G1237), .O(G1296) );
nand2 gate488( .a(G1238), .b(G1239), .O(G1297) );
nand2 gate489( .a(G1240), .b(G1241), .O(G1298) );
nand2 gate490( .a(G1242), .b(G1243), .O(G1299) );

  xor2  gate1121(.a(G1245), .b(G1244), .O(gate491inter0));
  nand2 gate1122(.a(gate491inter0), .b(s_82), .O(gate491inter1));
  and2  gate1123(.a(G1245), .b(G1244), .O(gate491inter2));
  inv1  gate1124(.a(s_82), .O(gate491inter3));
  inv1  gate1125(.a(s_83), .O(gate491inter4));
  nand2 gate1126(.a(gate491inter4), .b(gate491inter3), .O(gate491inter5));
  nor2  gate1127(.a(gate491inter5), .b(gate491inter2), .O(gate491inter6));
  inv1  gate1128(.a(G1244), .O(gate491inter7));
  inv1  gate1129(.a(G1245), .O(gate491inter8));
  nand2 gate1130(.a(gate491inter8), .b(gate491inter7), .O(gate491inter9));
  nand2 gate1131(.a(s_83), .b(gate491inter3), .O(gate491inter10));
  nor2  gate1132(.a(gate491inter10), .b(gate491inter9), .O(gate491inter11));
  nor2  gate1133(.a(gate491inter11), .b(gate491inter6), .O(gate491inter12));
  nand2 gate1134(.a(gate491inter12), .b(gate491inter1), .O(G1300));
nand2 gate492( .a(G1246), .b(G1247), .O(G1301) );
nand2 gate493( .a(G1248), .b(G1249), .O(G1302) );
nand2 gate494( .a(G1250), .b(G1251), .O(G1303) );
nand2 gate495( .a(G1252), .b(G1253), .O(G1304) );
nand2 gate496( .a(G1254), .b(G1255), .O(G1305) );
nand2 gate497( .a(G1256), .b(G1257), .O(G1306) );
nand2 gate498( .a(G1258), .b(G1259), .O(G1307) );
nand2 gate499( .a(G1260), .b(G1261), .O(G1308) );
nand2 gate500( .a(G1262), .b(G1263), .O(G1309) );
nand2 gate501( .a(G1264), .b(G1265), .O(G1310) );
nand2 gate502( .a(G1266), .b(G1267), .O(G1311) );
nand2 gate503( .a(G1268), .b(G1269), .O(G1312) );
nand2 gate504( .a(G1270), .b(G1271), .O(G1313) );
nand2 gate505( .a(G1272), .b(G1273), .O(G1314) );

  xor2  gate575(.a(G1275), .b(G1274), .O(gate506inter0));
  nand2 gate576(.a(gate506inter0), .b(s_4), .O(gate506inter1));
  and2  gate577(.a(G1275), .b(G1274), .O(gate506inter2));
  inv1  gate578(.a(s_4), .O(gate506inter3));
  inv1  gate579(.a(s_5), .O(gate506inter4));
  nand2 gate580(.a(gate506inter4), .b(gate506inter3), .O(gate506inter5));
  nor2  gate581(.a(gate506inter5), .b(gate506inter2), .O(gate506inter6));
  inv1  gate582(.a(G1274), .O(gate506inter7));
  inv1  gate583(.a(G1275), .O(gate506inter8));
  nand2 gate584(.a(gate506inter8), .b(gate506inter7), .O(gate506inter9));
  nand2 gate585(.a(s_5), .b(gate506inter3), .O(gate506inter10));
  nor2  gate586(.a(gate506inter10), .b(gate506inter9), .O(gate506inter11));
  nor2  gate587(.a(gate506inter11), .b(gate506inter6), .O(gate506inter12));
  nand2 gate588(.a(gate506inter12), .b(gate506inter1), .O(G1315));
nand2 gate507( .a(G1276), .b(G1277), .O(G1316) );
nand2 gate508( .a(G1278), .b(G1279), .O(G1317) );
nand2 gate509( .a(G1280), .b(G1281), .O(G1318) );
nand2 gate510( .a(G1282), .b(G1283), .O(G1319) );
nand2 gate511( .a(G1284), .b(G1285), .O(G1320) );
nand2 gate512( .a(G1286), .b(G1287), .O(G1321) );

  xor2  gate1359(.a(G1289), .b(G1288), .O(gate513inter0));
  nand2 gate1360(.a(gate513inter0), .b(s_116), .O(gate513inter1));
  and2  gate1361(.a(G1289), .b(G1288), .O(gate513inter2));
  inv1  gate1362(.a(s_116), .O(gate513inter3));
  inv1  gate1363(.a(s_117), .O(gate513inter4));
  nand2 gate1364(.a(gate513inter4), .b(gate513inter3), .O(gate513inter5));
  nor2  gate1365(.a(gate513inter5), .b(gate513inter2), .O(gate513inter6));
  inv1  gate1366(.a(G1288), .O(gate513inter7));
  inv1  gate1367(.a(G1289), .O(gate513inter8));
  nand2 gate1368(.a(gate513inter8), .b(gate513inter7), .O(gate513inter9));
  nand2 gate1369(.a(s_117), .b(gate513inter3), .O(gate513inter10));
  nor2  gate1370(.a(gate513inter10), .b(gate513inter9), .O(gate513inter11));
  nor2  gate1371(.a(gate513inter11), .b(gate513inter6), .O(gate513inter12));
  nand2 gate1372(.a(gate513inter12), .b(gate513inter1), .O(G1322));
nand2 gate514( .a(G1290), .b(G1291), .O(G1323) );
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule