module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);

input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;//RE__PI;

input s_0,s_1;//RE__ALLOW(00,01,10,11);
input s_2,s_3;//RE__ALLOW(00,01,10,11);
input s_4,s_5;//RE__ALLOW(00,01,10,11);
input s_6,s_7;//RE__ALLOW(00,01,10,11);
input s_8,s_9;//RE__ALLOW(00,01,10,11);
input s_10,s_11;//RE__ALLOW(00,01,10,11);
input s_12,s_13;//RE__ALLOW(00,01,10,11);
input s_14,s_15;//RE__ALLOW(00,01,10,11);
input s_16,s_17;//RE__ALLOW(00,01,10,11);
input s_18,s_19;//RE__ALLOW(00,01,10,11);
input s_20,s_21;//RE__ALLOW(00,01,10,11);
input s_22,s_23;//RE__ALLOW(00,01,10,11);
input s_24,s_25;//RE__ALLOW(00,01,10,11);
input s_26,s_27;//RE__ALLOW(00,01,10,11);
input s_28,s_29;//RE__ALLOW(00,01,10,11);
input s_30,s_31;//RE__ALLOW(00,01,10,11);
input s_32,s_33;//RE__ALLOW(00,01,10,11);
input s_34,s_35;//RE__ALLOW(00,01,10,11);
input s_36,s_37;//RE__ALLOW(00,01,10,11);
input s_38,s_39;//RE__ALLOW(00,01,10,11);
input s_40,s_41;//RE__ALLOW(00,01,10,11);
input s_42,s_43;//RE__ALLOW(00,01,10,11);
input s_44,s_45;//RE__ALLOW(00,01,10,11);
input s_46,s_47;//RE__ALLOW(00,01,10,11);
input s_48,s_49;//RE__ALLOW(00,01,10,11);
input s_50,s_51;//RE__ALLOW(00,01,10,11);
input s_52,s_53;//RE__ALLOW(00,01,10,11);
input s_54,s_55;//RE__ALLOW(00,01,10,11);
input s_56,s_57;//RE__ALLOW(00,01,10,11);
input s_58,s_59;//RE__ALLOW(00,01,10,11);
input s_60,s_61;//RE__ALLOW(00,01,10,11);
input s_62,s_63;//RE__ALLOW(00,01,10,11);
input s_64,s_65;//RE__ALLOW(00,01,10,11);
input s_66,s_67;//RE__ALLOW(00,01,10,11);
input s_68,s_69;//RE__ALLOW(00,01,10,11);
input s_70,s_71;//RE__ALLOW(00,01,10,11);
input s_72,s_73;//RE__ALLOW(00,01,10,11);
input s_74,s_75;//RE__ALLOW(00,01,10,11);
input s_76,s_77;//RE__ALLOW(00,01,10,11);
input s_78,s_79;//RE__ALLOW(00,01,10,11);
input s_80,s_81;//RE__ALLOW(00,01,10,11);
input s_82,s_83;//RE__ALLOW(00,01,10,11);
input s_84,s_85;//RE__ALLOW(00,01,10,11);
input s_86,s_87;//RE__ALLOW(00,01,10,11);
input s_88,s_89;//RE__ALLOW(00,01,10,11);
input s_90,s_91;//RE__ALLOW(00,01,10,11);
input s_92,s_93;//RE__ALLOW(00,01,10,11);
input s_94,s_95;//RE__ALLOW(00,01,10,11);
input s_96,s_97;//RE__ALLOW(00,01,10,11);
input s_98,s_99;//RE__ALLOW(00,01,10,11);
input s_100,s_101;//RE__ALLOW(00,01,10,11);
input s_102,s_103;//RE__ALLOW(00,01,10,11);
input s_104,s_105;//RE__ALLOW(00,01,10,11);
input s_106,s_107;//RE__ALLOW(00,01,10,11);
input s_108,s_109;//RE__ALLOW(00,01,10,11);
input s_110,s_111;//RE__ALLOW(00,01,10,11);
input s_112,s_113;//RE__ALLOW(00,01,10,11);
input s_114,s_115;//RE__ALLOW(00,01,10,11);
input s_116,s_117;//RE__ALLOW(00,01,10,11);
input s_118,s_119;//RE__ALLOW(00,01,10,11);
input s_120,s_121;//RE__ALLOW(00,01,10,11);
input s_122,s_123;//RE__ALLOW(00,01,10,11);
input s_124,s_125;//RE__ALLOW(00,01,10,11);
input s_126,s_127;//RE__ALLOW(00,01,10,11);
input s_128,s_129;//RE__ALLOW(00,01,10,11);
input s_130,s_131;//RE__ALLOW(00,01,10,11);
input s_132,s_133;//RE__ALLOW(00,01,10,11);
input s_134,s_135;//RE__ALLOW(00,01,10,11);
input s_136,s_137;//RE__ALLOW(00,01,10,11);
input s_138,s_139;//RE__ALLOW(00,01,10,11);
input s_140,s_141;//RE__ALLOW(00,01,10,11);
input s_142,s_143;//RE__ALLOW(00,01,10,11);
input s_144,s_145;//RE__ALLOW(00,01,10,11);
input s_146,s_147;//RE__ALLOW(00,01,10,11);
input s_148,s_149;//RE__ALLOW(00,01,10,11);
input s_150,s_151;//RE__ALLOW(00,01,10,11);
input s_152,s_153;//RE__ALLOW(00,01,10,11);
input s_154,s_155;//RE__ALLOW(00,01,10,11);
input s_156,s_157;//RE__ALLOW(00,01,10,11);
input s_158,s_159;//RE__ALLOW(00,01,10,11);
input s_160,s_161;//RE__ALLOW(00,01,10,11);
input s_162,s_163;//RE__ALLOW(00,01,10,11);
input s_164,s_165;//RE__ALLOW(00,01,10,11);
input s_166,s_167;//RE__ALLOW(00,01,10,11);
input s_168,s_169;//RE__ALLOW(00,01,10,11);
input s_170,s_171;//RE__ALLOW(00,01,10,11);
input s_172,s_173;//RE__ALLOW(00,01,10,11);
input s_174,s_175;//RE__ALLOW(00,01,10,11);
input s_176,s_177;//RE__ALLOW(00,01,10,11);
input s_178,s_179;//RE__ALLOW(00,01,10,11);
input s_180,s_181;//RE__ALLOW(00,01,10,11);
input s_182,s_183;//RE__ALLOW(00,01,10,11);
input s_184,s_185;//RE__ALLOW(00,01,10,11);
input s_186,s_187;//RE__ALLOW(00,01,10,11);
input s_188,s_189;//RE__ALLOW(00,01,10,11);
input s_190,s_191;//RE__ALLOW(00,01,10,11);
input s_192,s_193;//RE__ALLOW(00,01,10,11);
input s_194,s_195;//RE__ALLOW(00,01,10,11);
input s_196,s_197;//RE__ALLOW(00,01,10,11);
input s_198,s_199;//RE__ALLOW(00,01,10,11);
input s_200,s_201;//RE__ALLOW(00,01,10,11);
input s_202,s_203;//RE__ALLOW(00,01,10,11);
input s_204,s_205;//RE__ALLOW(00,01,10,11);
input s_206,s_207;//RE__ALLOW(00,01,10,11);
input s_208,s_209;//RE__ALLOW(00,01,10,11);
input s_210,s_211;//RE__ALLOW(00,01,10,11);
input s_212,s_213;//RE__ALLOW(00,01,10,11);
input s_214,s_215;//RE__ALLOW(00,01,10,11);
input s_216,s_217;//RE__ALLOW(00,01,10,11);
input s_218,s_219;//RE__ALLOW(00,01,10,11);
input s_220,s_221;//RE__ALLOW(00,01,10,11);
input s_222,s_223;//RE__ALLOW(00,01,10,11);
input s_224,s_225;//RE__ALLOW(00,01,10,11);
input s_226,s_227;//RE__ALLOW(00,01,10,11);
input s_228,s_229;//RE__ALLOW(00,01,10,11);
input s_230,s_231;//RE__ALLOW(00,01,10,11);
input s_232,s_233;//RE__ALLOW(00,01,10,11);
input s_234,s_235;//RE__ALLOW(00,01,10,11);
input s_236,s_237;//RE__ALLOW(00,01,10,11);
input s_238,s_239;//RE__ALLOW(00,01,10,11);
input s_240,s_241;//RE__ALLOW(00,01,10,11);
input s_242,s_243;//RE__ALLOW(00,01,10,11);
input s_244,s_245;//RE__ALLOW(00,01,10,11);
input s_246,s_247;//RE__ALLOW(00,01,10,11);
input s_248,s_249;//RE__ALLOW(00,01,10,11);
input s_250,s_251;//RE__ALLOW(00,01,10,11);
input s_252,s_253;//RE__ALLOW(00,01,10,11);
input s_254,s_255;//RE__ALLOW(00,01,10,11);
input s_256,s_257;//RE__ALLOW(00,01,10,11);
input s_258,s_259;//RE__ALLOW(00,01,10,11);
input s_260,s_261;//RE__ALLOW(00,01,10,11);
input s_262,s_263;//RE__ALLOW(00,01,10,11);
input s_264,s_265;//RE__ALLOW(00,01,10,11);
input s_266,s_267;//RE__ALLOW(00,01,10,11);
input s_268,s_269;//RE__ALLOW(00,01,10,11);
input s_270,s_271;//RE__ALLOW(00,01,10,11);
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;

  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate454inter0, gate454inter1, gate454inter2, gate454inter3, gate454inter4, gate454inter5, gate454inter6, gate454inter7, gate454inter8, gate454inter9, gate454inter10, gate454inter11, gate454inter12, gate58inter0, gate58inter1, gate58inter2, gate58inter3, gate58inter4, gate58inter5, gate58inter6, gate58inter7, gate58inter8, gate58inter9, gate58inter10, gate58inter11, gate58inter12, gate217inter0, gate217inter1, gate217inter2, gate217inter3, gate217inter4, gate217inter5, gate217inter6, gate217inter7, gate217inter8, gate217inter9, gate217inter10, gate217inter11, gate217inter12, gate209inter0, gate209inter1, gate209inter2, gate209inter3, gate209inter4, gate209inter5, gate209inter6, gate209inter7, gate209inter8, gate209inter9, gate209inter10, gate209inter11, gate209inter12, gate260inter0, gate260inter1, gate260inter2, gate260inter3, gate260inter4, gate260inter5, gate260inter6, gate260inter7, gate260inter8, gate260inter9, gate260inter10, gate260inter11, gate260inter12, gate9inter0, gate9inter1, gate9inter2, gate9inter3, gate9inter4, gate9inter5, gate9inter6, gate9inter7, gate9inter8, gate9inter9, gate9inter10, gate9inter11, gate9inter12, gate141inter0, gate141inter1, gate141inter2, gate141inter3, gate141inter4, gate141inter5, gate141inter6, gate141inter7, gate141inter8, gate141inter9, gate141inter10, gate141inter11, gate141inter12, gate245inter0, gate245inter1, gate245inter2, gate245inter3, gate245inter4, gate245inter5, gate245inter6, gate245inter7, gate245inter8, gate245inter9, gate245inter10, gate245inter11, gate245inter12, gate126inter0, gate126inter1, gate126inter2, gate126inter3, gate126inter4, gate126inter5, gate126inter6, gate126inter7, gate126inter8, gate126inter9, gate126inter10, gate126inter11, gate126inter12, gate121inter0, gate121inter1, gate121inter2, gate121inter3, gate121inter4, gate121inter5, gate121inter6, gate121inter7, gate121inter8, gate121inter9, gate121inter10, gate121inter11, gate121inter12, gate390inter0, gate390inter1, gate390inter2, gate390inter3, gate390inter4, gate390inter5, gate390inter6, gate390inter7, gate390inter8, gate390inter9, gate390inter10, gate390inter11, gate390inter12, gate270inter0, gate270inter1, gate270inter2, gate270inter3, gate270inter4, gate270inter5, gate270inter6, gate270inter7, gate270inter8, gate270inter9, gate270inter10, gate270inter11, gate270inter12, gate465inter0, gate465inter1, gate465inter2, gate465inter3, gate465inter4, gate465inter5, gate465inter6, gate465inter7, gate465inter8, gate465inter9, gate465inter10, gate465inter11, gate465inter12, gate46inter0, gate46inter1, gate46inter2, gate46inter3, gate46inter4, gate46inter5, gate46inter6, gate46inter7, gate46inter8, gate46inter9, gate46inter10, gate46inter11, gate46inter12, gate216inter0, gate216inter1, gate216inter2, gate216inter3, gate216inter4, gate216inter5, gate216inter6, gate216inter7, gate216inter8, gate216inter9, gate216inter10, gate216inter11, gate216inter12, gate289inter0, gate289inter1, gate289inter2, gate289inter3, gate289inter4, gate289inter5, gate289inter6, gate289inter7, gate289inter8, gate289inter9, gate289inter10, gate289inter11, gate289inter12, gate63inter0, gate63inter1, gate63inter2, gate63inter3, gate63inter4, gate63inter5, gate63inter6, gate63inter7, gate63inter8, gate63inter9, gate63inter10, gate63inter11, gate63inter12, gate467inter0, gate467inter1, gate467inter2, gate467inter3, gate467inter4, gate467inter5, gate467inter6, gate467inter7, gate467inter8, gate467inter9, gate467inter10, gate467inter11, gate467inter12, gate59inter0, gate59inter1, gate59inter2, gate59inter3, gate59inter4, gate59inter5, gate59inter6, gate59inter7, gate59inter8, gate59inter9, gate59inter10, gate59inter11, gate59inter12, gate17inter0, gate17inter1, gate17inter2, gate17inter3, gate17inter4, gate17inter5, gate17inter6, gate17inter7, gate17inter8, gate17inter9, gate17inter10, gate17inter11, gate17inter12, gate70inter0, gate70inter1, gate70inter2, gate70inter3, gate70inter4, gate70inter5, gate70inter6, gate70inter7, gate70inter8, gate70inter9, gate70inter10, gate70inter11, gate70inter12, gate492inter0, gate492inter1, gate492inter2, gate492inter3, gate492inter4, gate492inter5, gate492inter6, gate492inter7, gate492inter8, gate492inter9, gate492inter10, gate492inter11, gate492inter12, gate73inter0, gate73inter1, gate73inter2, gate73inter3, gate73inter4, gate73inter5, gate73inter6, gate73inter7, gate73inter8, gate73inter9, gate73inter10, gate73inter11, gate73inter12, gate11inter0, gate11inter1, gate11inter2, gate11inter3, gate11inter4, gate11inter5, gate11inter6, gate11inter7, gate11inter8, gate11inter9, gate11inter10, gate11inter11, gate11inter12, gate428inter0, gate428inter1, gate428inter2, gate428inter3, gate428inter4, gate428inter5, gate428inter6, gate428inter7, gate428inter8, gate428inter9, gate428inter10, gate428inter11, gate428inter12, gate143inter0, gate143inter1, gate143inter2, gate143inter3, gate143inter4, gate143inter5, gate143inter6, gate143inter7, gate143inter8, gate143inter9, gate143inter10, gate143inter11, gate143inter12, gate468inter0, gate468inter1, gate468inter2, gate468inter3, gate468inter4, gate468inter5, gate468inter6, gate468inter7, gate468inter8, gate468inter9, gate468inter10, gate468inter11, gate468inter12, gate483inter0, gate483inter1, gate483inter2, gate483inter3, gate483inter4, gate483inter5, gate483inter6, gate483inter7, gate483inter8, gate483inter9, gate483inter10, gate483inter11, gate483inter12, gate111inter0, gate111inter1, gate111inter2, gate111inter3, gate111inter4, gate111inter5, gate111inter6, gate111inter7, gate111inter8, gate111inter9, gate111inter10, gate111inter11, gate111inter12, gate231inter0, gate231inter1, gate231inter2, gate231inter3, gate231inter4, gate231inter5, gate231inter6, gate231inter7, gate231inter8, gate231inter9, gate231inter10, gate231inter11, gate231inter12, gate222inter0, gate222inter1, gate222inter2, gate222inter3, gate222inter4, gate222inter5, gate222inter6, gate222inter7, gate222inter8, gate222inter9, gate222inter10, gate222inter11, gate222inter12, gate192inter0, gate192inter1, gate192inter2, gate192inter3, gate192inter4, gate192inter5, gate192inter6, gate192inter7, gate192inter8, gate192inter9, gate192inter10, gate192inter11, gate192inter12, gate211inter0, gate211inter1, gate211inter2, gate211inter3, gate211inter4, gate211inter5, gate211inter6, gate211inter7, gate211inter8, gate211inter9, gate211inter10, gate211inter11, gate211inter12, gate86inter0, gate86inter1, gate86inter2, gate86inter3, gate86inter4, gate86inter5, gate86inter6, gate86inter7, gate86inter8, gate86inter9, gate86inter10, gate86inter11, gate86inter12, gate18inter0, gate18inter1, gate18inter2, gate18inter3, gate18inter4, gate18inter5, gate18inter6, gate18inter7, gate18inter8, gate18inter9, gate18inter10, gate18inter11, gate18inter12, gate109inter0, gate109inter1, gate109inter2, gate109inter3, gate109inter4, gate109inter5, gate109inter6, gate109inter7, gate109inter8, gate109inter9, gate109inter10, gate109inter11, gate109inter12, gate138inter0, gate138inter1, gate138inter2, gate138inter3, gate138inter4, gate138inter5, gate138inter6, gate138inter7, gate138inter8, gate138inter9, gate138inter10, gate138inter11, gate138inter12, gate159inter0, gate159inter1, gate159inter2, gate159inter3, gate159inter4, gate159inter5, gate159inter6, gate159inter7, gate159inter8, gate159inter9, gate159inter10, gate159inter11, gate159inter12, gate153inter0, gate153inter1, gate153inter2, gate153inter3, gate153inter4, gate153inter5, gate153inter6, gate153inter7, gate153inter8, gate153inter9, gate153inter10, gate153inter11, gate153inter12, gate513inter0, gate513inter1, gate513inter2, gate513inter3, gate513inter4, gate513inter5, gate513inter6, gate513inter7, gate513inter8, gate513inter9, gate513inter10, gate513inter11, gate513inter12, gate204inter0, gate204inter1, gate204inter2, gate204inter3, gate204inter4, gate204inter5, gate204inter6, gate204inter7, gate204inter8, gate204inter9, gate204inter10, gate204inter11, gate204inter12, gate39inter0, gate39inter1, gate39inter2, gate39inter3, gate39inter4, gate39inter5, gate39inter6, gate39inter7, gate39inter8, gate39inter9, gate39inter10, gate39inter11, gate39inter12, gate110inter0, gate110inter1, gate110inter2, gate110inter3, gate110inter4, gate110inter5, gate110inter6, gate110inter7, gate110inter8, gate110inter9, gate110inter10, gate110inter11, gate110inter12, gate435inter0, gate435inter1, gate435inter2, gate435inter3, gate435inter4, gate435inter5, gate435inter6, gate435inter7, gate435inter8, gate435inter9, gate435inter10, gate435inter11, gate435inter12, gate254inter0, gate254inter1, gate254inter2, gate254inter3, gate254inter4, gate254inter5, gate254inter6, gate254inter7, gate254inter8, gate254inter9, gate254inter10, gate254inter11, gate254inter12, gate200inter0, gate200inter1, gate200inter2, gate200inter3, gate200inter4, gate200inter5, gate200inter6, gate200inter7, gate200inter8, gate200inter9, gate200inter10, gate200inter11, gate200inter12, gate52inter0, gate52inter1, gate52inter2, gate52inter3, gate52inter4, gate52inter5, gate52inter6, gate52inter7, gate52inter8, gate52inter9, gate52inter10, gate52inter11, gate52inter12, gate511inter0, gate511inter1, gate511inter2, gate511inter3, gate511inter4, gate511inter5, gate511inter6, gate511inter7, gate511inter8, gate511inter9, gate511inter10, gate511inter11, gate511inter12, gate491inter0, gate491inter1, gate491inter2, gate491inter3, gate491inter4, gate491inter5, gate491inter6, gate491inter7, gate491inter8, gate491inter9, gate491inter10, gate491inter11, gate491inter12, gate173inter0, gate173inter1, gate173inter2, gate173inter3, gate173inter4, gate173inter5, gate173inter6, gate173inter7, gate173inter8, gate173inter9, gate173inter10, gate173inter11, gate173inter12, gate122inter0, gate122inter1, gate122inter2, gate122inter3, gate122inter4, gate122inter5, gate122inter6, gate122inter7, gate122inter8, gate122inter9, gate122inter10, gate122inter11, gate122inter12, gate482inter0, gate482inter1, gate482inter2, gate482inter3, gate482inter4, gate482inter5, gate482inter6, gate482inter7, gate482inter8, gate482inter9, gate482inter10, gate482inter11, gate482inter12, gate32inter0, gate32inter1, gate32inter2, gate32inter3, gate32inter4, gate32inter5, gate32inter6, gate32inter7, gate32inter8, gate32inter9, gate32inter10, gate32inter11, gate32inter12, gate434inter0, gate434inter1, gate434inter2, gate434inter3, gate434inter4, gate434inter5, gate434inter6, gate434inter7, gate434inter8, gate434inter9, gate434inter10, gate434inter11, gate434inter12, gate197inter0, gate197inter1, gate197inter2, gate197inter3, gate197inter4, gate197inter5, gate197inter6, gate197inter7, gate197inter8, gate197inter9, gate197inter10, gate197inter11, gate197inter12, gate66inter0, gate66inter1, gate66inter2, gate66inter3, gate66inter4, gate66inter5, gate66inter6, gate66inter7, gate66inter8, gate66inter9, gate66inter10, gate66inter11, gate66inter12, gate210inter0, gate210inter1, gate210inter2, gate210inter3, gate210inter4, gate210inter5, gate210inter6, gate210inter7, gate210inter8, gate210inter9, gate210inter10, gate210inter11, gate210inter12, gate56inter0, gate56inter1, gate56inter2, gate56inter3, gate56inter4, gate56inter5, gate56inter6, gate56inter7, gate56inter8, gate56inter9, gate56inter10, gate56inter11, gate56inter12, gate55inter0, gate55inter1, gate55inter2, gate55inter3, gate55inter4, gate55inter5, gate55inter6, gate55inter7, gate55inter8, gate55inter9, gate55inter10, gate55inter11, gate55inter12, gate161inter0, gate161inter1, gate161inter2, gate161inter3, gate161inter4, gate161inter5, gate161inter6, gate161inter7, gate161inter8, gate161inter9, gate161inter10, gate161inter11, gate161inter12, gate388inter0, gate388inter1, gate388inter2, gate388inter3, gate388inter4, gate388inter5, gate388inter6, gate388inter7, gate388inter8, gate388inter9, gate388inter10, gate388inter11, gate388inter12, gate237inter0, gate237inter1, gate237inter2, gate237inter3, gate237inter4, gate237inter5, gate237inter6, gate237inter7, gate237inter8, gate237inter9, gate237inter10, gate237inter11, gate237inter12, gate94inter0, gate94inter1, gate94inter2, gate94inter3, gate94inter4, gate94inter5, gate94inter6, gate94inter7, gate94inter8, gate94inter9, gate94inter10, gate94inter11, gate94inter12, gate142inter0, gate142inter1, gate142inter2, gate142inter3, gate142inter4, gate142inter5, gate142inter6, gate142inter7, gate142inter8, gate142inter9, gate142inter10, gate142inter11, gate142inter12, gate414inter0, gate414inter1, gate414inter2, gate414inter3, gate414inter4, gate414inter5, gate414inter6, gate414inter7, gate414inter8, gate414inter9, gate414inter10, gate414inter11, gate414inter12, gate432inter0, gate432inter1, gate432inter2, gate432inter3, gate432inter4, gate432inter5, gate432inter6, gate432inter7, gate432inter8, gate432inter9, gate432inter10, gate432inter11, gate432inter12, gate463inter0, gate463inter1, gate463inter2, gate463inter3, gate463inter4, gate463inter5, gate463inter6, gate463inter7, gate463inter8, gate463inter9, gate463inter10, gate463inter11, gate463inter12, gate43inter0, gate43inter1, gate43inter2, gate43inter3, gate43inter4, gate43inter5, gate43inter6, gate43inter7, gate43inter8, gate43inter9, gate43inter10, gate43inter11, gate43inter12, gate190inter0, gate190inter1, gate190inter2, gate190inter3, gate190inter4, gate190inter5, gate190inter6, gate190inter7, gate190inter8, gate190inter9, gate190inter10, gate190inter11, gate190inter12, gate477inter0, gate477inter1, gate477inter2, gate477inter3, gate477inter4, gate477inter5, gate477inter6, gate477inter7, gate477inter8, gate477inter9, gate477inter10, gate477inter11, gate477inter12, gate144inter0, gate144inter1, gate144inter2, gate144inter3, gate144inter4, gate144inter5, gate144inter6, gate144inter7, gate144inter8, gate144inter9, gate144inter10, gate144inter11, gate144inter12, gate445inter0, gate445inter1, gate445inter2, gate445inter3, gate445inter4, gate445inter5, gate445inter6, gate445inter7, gate445inter8, gate445inter9, gate445inter10, gate445inter11, gate445inter12, gate436inter0, gate436inter1, gate436inter2, gate436inter3, gate436inter4, gate436inter5, gate436inter6, gate436inter7, gate436inter8, gate436inter9, gate436inter10, gate436inter11, gate436inter12, gate514inter0, gate514inter1, gate514inter2, gate514inter3, gate514inter4, gate514inter5, gate514inter6, gate514inter7, gate514inter8, gate514inter9, gate514inter10, gate514inter11, gate514inter12, gate187inter0, gate187inter1, gate187inter2, gate187inter3, gate187inter4, gate187inter5, gate187inter6, gate187inter7, gate187inter8, gate187inter9, gate187inter10, gate187inter11, gate187inter12, gate252inter0, gate252inter1, gate252inter2, gate252inter3, gate252inter4, gate252inter5, gate252inter6, gate252inter7, gate252inter8, gate252inter9, gate252inter10, gate252inter11, gate252inter12, gate175inter0, gate175inter1, gate175inter2, gate175inter3, gate175inter4, gate175inter5, gate175inter6, gate175inter7, gate175inter8, gate175inter9, gate175inter10, gate175inter11, gate175inter12, gate403inter0, gate403inter1, gate403inter2, gate403inter3, gate403inter4, gate403inter5, gate403inter6, gate403inter7, gate403inter8, gate403inter9, gate403inter10, gate403inter11, gate403inter12, gate54inter0, gate54inter1, gate54inter2, gate54inter3, gate54inter4, gate54inter5, gate54inter6, gate54inter7, gate54inter8, gate54inter9, gate54inter10, gate54inter11, gate54inter12, gate233inter0, gate233inter1, gate233inter2, gate233inter3, gate233inter4, gate233inter5, gate233inter6, gate233inter7, gate233inter8, gate233inter9, gate233inter10, gate233inter11, gate233inter12, gate83inter0, gate83inter1, gate83inter2, gate83inter3, gate83inter4, gate83inter5, gate83inter6, gate83inter7, gate83inter8, gate83inter9, gate83inter10, gate83inter11, gate83inter12, gate137inter0, gate137inter1, gate137inter2, gate137inter3, gate137inter4, gate137inter5, gate137inter6, gate137inter7, gate137inter8, gate137inter9, gate137inter10, gate137inter11, gate137inter12, gate87inter0, gate87inter1, gate87inter2, gate87inter3, gate87inter4, gate87inter5, gate87inter6, gate87inter7, gate87inter8, gate87inter9, gate87inter10, gate87inter11, gate87inter12, gate31inter0, gate31inter1, gate31inter2, gate31inter3, gate31inter4, gate31inter5, gate31inter6, gate31inter7, gate31inter8, gate31inter9, gate31inter10, gate31inter11, gate31inter12, gate164inter0, gate164inter1, gate164inter2, gate164inter3, gate164inter4, gate164inter5, gate164inter6, gate164inter7, gate164inter8, gate164inter9, gate164inter10, gate164inter11, gate164inter12, gate154inter0, gate154inter1, gate154inter2, gate154inter3, gate154inter4, gate154inter5, gate154inter6, gate154inter7, gate154inter8, gate154inter9, gate154inter10, gate154inter11, gate154inter12, gate487inter0, gate487inter1, gate487inter2, gate487inter3, gate487inter4, gate487inter5, gate487inter6, gate487inter7, gate487inter8, gate487inter9, gate487inter10, gate487inter11, gate487inter12, gate439inter0, gate439inter1, gate439inter2, gate439inter3, gate439inter4, gate439inter5, gate439inter6, gate439inter7, gate439inter8, gate439inter9, gate439inter10, gate439inter11, gate439inter12, gate389inter0, gate389inter1, gate389inter2, gate389inter3, gate389inter4, gate389inter5, gate389inter6, gate389inter7, gate389inter8, gate389inter9, gate389inter10, gate389inter11, gate389inter12, gate168inter0, gate168inter1, gate168inter2, gate168inter3, gate168inter4, gate168inter5, gate168inter6, gate168inter7, gate168inter8, gate168inter9, gate168inter10, gate168inter11, gate168inter12, gate494inter0, gate494inter1, gate494inter2, gate494inter3, gate494inter4, gate494inter5, gate494inter6, gate494inter7, gate494inter8, gate494inter9, gate494inter10, gate494inter11, gate494inter12, gate395inter0, gate395inter1, gate395inter2, gate395inter3, gate395inter4, gate395inter5, gate395inter6, gate395inter7, gate395inter8, gate395inter9, gate395inter10, gate395inter11, gate395inter12, gate205inter0, gate205inter1, gate205inter2, gate205inter3, gate205inter4, gate205inter5, gate205inter6, gate205inter7, gate205inter8, gate205inter9, gate205inter10, gate205inter11, gate205inter12, gate219inter0, gate219inter1, gate219inter2, gate219inter3, gate219inter4, gate219inter5, gate219inter6, gate219inter7, gate219inter8, gate219inter9, gate219inter10, gate219inter11, gate219inter12, gate440inter0, gate440inter1, gate440inter2, gate440inter3, gate440inter4, gate440inter5, gate440inter6, gate440inter7, gate440inter8, gate440inter9, gate440inter10, gate440inter11, gate440inter12, gate106inter0, gate106inter1, gate106inter2, gate106inter3, gate106inter4, gate106inter5, gate106inter6, gate106inter7, gate106inter8, gate106inter9, gate106inter10, gate106inter11, gate106inter12, gate500inter0, gate500inter1, gate500inter2, gate500inter3, gate500inter4, gate500inter5, gate500inter6, gate500inter7, gate500inter8, gate500inter9, gate500inter10, gate500inter11, gate500inter12, gate234inter0, gate234inter1, gate234inter2, gate234inter3, gate234inter4, gate234inter5, gate234inter6, gate234inter7, gate234inter8, gate234inter9, gate234inter10, gate234inter11, gate234inter12, gate512inter0, gate512inter1, gate512inter2, gate512inter3, gate512inter4, gate512inter5, gate512inter6, gate512inter7, gate512inter8, gate512inter9, gate512inter10, gate512inter11, gate512inter12, gate189inter0, gate189inter1, gate189inter2, gate189inter3, gate189inter4, gate189inter5, gate189inter6, gate189inter7, gate189inter8, gate189inter9, gate189inter10, gate189inter11, gate189inter12, gate212inter0, gate212inter1, gate212inter2, gate212inter3, gate212inter4, gate212inter5, gate212inter6, gate212inter7, gate212inter8, gate212inter9, gate212inter10, gate212inter11, gate212inter12, gate459inter0, gate459inter1, gate459inter2, gate459inter3, gate459inter4, gate459inter5, gate459inter6, gate459inter7, gate459inter8, gate459inter9, gate459inter10, gate459inter11, gate459inter12, gate256inter0, gate256inter1, gate256inter2, gate256inter3, gate256inter4, gate256inter5, gate256inter6, gate256inter7, gate256inter8, gate256inter9, gate256inter10, gate256inter11, gate256inter12, gate507inter0, gate507inter1, gate507inter2, gate507inter3, gate507inter4, gate507inter5, gate507inter6, gate507inter7, gate507inter8, gate507inter9, gate507inter10, gate507inter11, gate507inter12, gate49inter0, gate49inter1, gate49inter2, gate49inter3, gate49inter4, gate49inter5, gate49inter6, gate49inter7, gate49inter8, gate49inter9, gate49inter10, gate49inter11, gate49inter12, gate246inter0, gate246inter1, gate246inter2, gate246inter3, gate246inter4, gate246inter5, gate246inter6, gate246inter7, gate246inter8, gate246inter9, gate246inter10, gate246inter11, gate246inter12, gate262inter0, gate262inter1, gate262inter2, gate262inter3, gate262inter4, gate262inter5, gate262inter6, gate262inter7, gate262inter8, gate262inter9, gate262inter10, gate262inter11, gate262inter12, gate131inter0, gate131inter1, gate131inter2, gate131inter3, gate131inter4, gate131inter5, gate131inter6, gate131inter7, gate131inter8, gate131inter9, gate131inter10, gate131inter11, gate131inter12, gate119inter0, gate119inter1, gate119inter2, gate119inter3, gate119inter4, gate119inter5, gate119inter6, gate119inter7, gate119inter8, gate119inter9, gate119inter10, gate119inter11, gate119inter12, gate10inter0, gate10inter1, gate10inter2, gate10inter3, gate10inter4, gate10inter5, gate10inter6, gate10inter7, gate10inter8, gate10inter9, gate10inter10, gate10inter11, gate10inter12, gate201inter0, gate201inter1, gate201inter2, gate201inter3, gate201inter4, gate201inter5, gate201inter6, gate201inter7, gate201inter8, gate201inter9, gate201inter10, gate201inter11, gate201inter12, gate253inter0, gate253inter1, gate253inter2, gate253inter3, gate253inter4, gate253inter5, gate253inter6, gate253inter7, gate253inter8, gate253inter9, gate253inter10, gate253inter11, gate253inter12, gate165inter0, gate165inter1, gate165inter2, gate165inter3, gate165inter4, gate165inter5, gate165inter6, gate165inter7, gate165inter8, gate165inter9, gate165inter10, gate165inter11, gate165inter12, gate80inter0, gate80inter1, gate80inter2, gate80inter3, gate80inter4, gate80inter5, gate80inter6, gate80inter7, gate80inter8, gate80inter9, gate80inter10, gate80inter11, gate80inter12, gate37inter0, gate37inter1, gate37inter2, gate37inter3, gate37inter4, gate37inter5, gate37inter6, gate37inter7, gate37inter8, gate37inter9, gate37inter10, gate37inter11, gate37inter12, gate238inter0, gate238inter1, gate238inter2, gate238inter3, gate238inter4, gate238inter5, gate238inter6, gate238inter7, gate238inter8, gate238inter9, gate238inter10, gate238inter11, gate238inter12, gate291inter0, gate291inter1, gate291inter2, gate291inter3, gate291inter4, gate291inter5, gate291inter6, gate291inter7, gate291inter8, gate291inter9, gate291inter10, gate291inter11, gate291inter12, gate29inter0, gate29inter1, gate29inter2, gate29inter3, gate29inter4, gate29inter5, gate29inter6, gate29inter7, gate29inter8, gate29inter9, gate29inter10, gate29inter11, gate29inter12, gate421inter0, gate421inter1, gate421inter2, gate421inter3, gate421inter4, gate421inter5, gate421inter6, gate421inter7, gate421inter8, gate421inter9, gate421inter10, gate421inter11, gate421inter12, gate407inter0, gate407inter1, gate407inter2, gate407inter3, gate407inter4, gate407inter5, gate407inter6, gate407inter7, gate407inter8, gate407inter9, gate407inter10, gate407inter11, gate407inter12, gate426inter0, gate426inter1, gate426inter2, gate426inter3, gate426inter4, gate426inter5, gate426inter6, gate426inter7, gate426inter8, gate426inter9, gate426inter10, gate426inter11, gate426inter12, gate38inter0, gate38inter1, gate38inter2, gate38inter3, gate38inter4, gate38inter5, gate38inter6, gate38inter7, gate38inter8, gate38inter9, gate38inter10, gate38inter11, gate38inter12, gate258inter0, gate258inter1, gate258inter2, gate258inter3, gate258inter4, gate258inter5, gate258inter6, gate258inter7, gate258inter8, gate258inter9, gate258inter10, gate258inter11, gate258inter12, gate493inter0, gate493inter1, gate493inter2, gate493inter3, gate493inter4, gate493inter5, gate493inter6, gate493inter7, gate493inter8, gate493inter9, gate493inter10, gate493inter11, gate493inter12, gate453inter0, gate453inter1, gate453inter2, gate453inter3, gate453inter4, gate453inter5, gate453inter6, gate453inter7, gate453inter8, gate453inter9, gate453inter10, gate453inter11, gate453inter12, gate248inter0, gate248inter1, gate248inter2, gate248inter3, gate248inter4, gate248inter5, gate248inter6, gate248inter7, gate248inter8, gate248inter9, gate248inter10, gate248inter11, gate248inter12, gate146inter0, gate146inter1, gate146inter2, gate146inter3, gate146inter4, gate146inter5, gate146inter6, gate146inter7, gate146inter8, gate146inter9, gate146inter10, gate146inter11, gate146inter12, gate150inter0, gate150inter1, gate150inter2, gate150inter3, gate150inter4, gate150inter5, gate150inter6, gate150inter7, gate150inter8, gate150inter9, gate150inter10, gate150inter11, gate150inter12, gate472inter0, gate472inter1, gate472inter2, gate472inter3, gate472inter4, gate472inter5, gate472inter6, gate472inter7, gate472inter8, gate472inter9, gate472inter10, gate472inter11, gate472inter12, gate294inter0, gate294inter1, gate294inter2, gate294inter3, gate294inter4, gate294inter5, gate294inter6, gate294inter7, gate294inter8, gate294inter9, gate294inter10, gate294inter11, gate294inter12, gate404inter0, gate404inter1, gate404inter2, gate404inter3, gate404inter4, gate404inter5, gate404inter6, gate404inter7, gate404inter8, gate404inter9, gate404inter10, gate404inter11, gate404inter12, gate41inter0, gate41inter1, gate41inter2, gate41inter3, gate41inter4, gate41inter5, gate41inter6, gate41inter7, gate41inter8, gate41inter9, gate41inter10, gate41inter11, gate41inter12, gate401inter0, gate401inter1, gate401inter2, gate401inter3, gate401inter4, gate401inter5, gate401inter6, gate401inter7, gate401inter8, gate401inter9, gate401inter10, gate401inter11, gate401inter12, gate127inter0, gate127inter1, gate127inter2, gate127inter3, gate127inter4, gate127inter5, gate127inter6, gate127inter7, gate127inter8, gate127inter9, gate127inter10, gate127inter11, gate127inter12, gate218inter0, gate218inter1, gate218inter2, gate218inter3, gate218inter4, gate218inter5, gate218inter6, gate218inter7, gate218inter8, gate218inter9, gate218inter10, gate218inter11, gate218inter12, gate391inter0, gate391inter1, gate391inter2, gate391inter3, gate391inter4, gate391inter5, gate391inter6, gate391inter7, gate391inter8, gate391inter9, gate391inter10, gate391inter11, gate391inter12;



and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );

  xor2  gate617(.a(G2), .b(G1), .O(gate9inter0));
  nand2 gate618(.a(gate9inter0), .b(s_10), .O(gate9inter1));
  and2  gate619(.a(G2), .b(G1), .O(gate9inter2));
  inv1  gate620(.a(s_10), .O(gate9inter3));
  inv1  gate621(.a(s_11), .O(gate9inter4));
  nand2 gate622(.a(gate9inter4), .b(gate9inter3), .O(gate9inter5));
  nor2  gate623(.a(gate9inter5), .b(gate9inter2), .O(gate9inter6));
  inv1  gate624(.a(G1), .O(gate9inter7));
  inv1  gate625(.a(G2), .O(gate9inter8));
  nand2 gate626(.a(gate9inter8), .b(gate9inter7), .O(gate9inter9));
  nand2 gate627(.a(s_11), .b(gate9inter3), .O(gate9inter10));
  nor2  gate628(.a(gate9inter10), .b(gate9inter9), .O(gate9inter11));
  nor2  gate629(.a(gate9inter11), .b(gate9inter6), .O(gate9inter12));
  nand2 gate630(.a(gate9inter12), .b(gate9inter1), .O(G266));

  xor2  gate2073(.a(G4), .b(G3), .O(gate10inter0));
  nand2 gate2074(.a(gate10inter0), .b(s_218), .O(gate10inter1));
  and2  gate2075(.a(G4), .b(G3), .O(gate10inter2));
  inv1  gate2076(.a(s_218), .O(gate10inter3));
  inv1  gate2077(.a(s_219), .O(gate10inter4));
  nand2 gate2078(.a(gate10inter4), .b(gate10inter3), .O(gate10inter5));
  nor2  gate2079(.a(gate10inter5), .b(gate10inter2), .O(gate10inter6));
  inv1  gate2080(.a(G3), .O(gate10inter7));
  inv1  gate2081(.a(G4), .O(gate10inter8));
  nand2 gate2082(.a(gate10inter8), .b(gate10inter7), .O(gate10inter9));
  nand2 gate2083(.a(s_219), .b(gate10inter3), .O(gate10inter10));
  nor2  gate2084(.a(gate10inter10), .b(gate10inter9), .O(gate10inter11));
  nor2  gate2085(.a(gate10inter11), .b(gate10inter6), .O(gate10inter12));
  nand2 gate2086(.a(gate10inter12), .b(gate10inter1), .O(G269));

  xor2  gate869(.a(G6), .b(G5), .O(gate11inter0));
  nand2 gate870(.a(gate11inter0), .b(s_46), .O(gate11inter1));
  and2  gate871(.a(G6), .b(G5), .O(gate11inter2));
  inv1  gate872(.a(s_46), .O(gate11inter3));
  inv1  gate873(.a(s_47), .O(gate11inter4));
  nand2 gate874(.a(gate11inter4), .b(gate11inter3), .O(gate11inter5));
  nor2  gate875(.a(gate11inter5), .b(gate11inter2), .O(gate11inter6));
  inv1  gate876(.a(G5), .O(gate11inter7));
  inv1  gate877(.a(G6), .O(gate11inter8));
  nand2 gate878(.a(gate11inter8), .b(gate11inter7), .O(gate11inter9));
  nand2 gate879(.a(s_47), .b(gate11inter3), .O(gate11inter10));
  nor2  gate880(.a(gate11inter10), .b(gate11inter9), .O(gate11inter11));
  nor2  gate881(.a(gate11inter11), .b(gate11inter6), .O(gate11inter12));
  nand2 gate882(.a(gate11inter12), .b(gate11inter1), .O(G272));
nand2 gate12( .a(G7), .b(G8), .O(G275) );
nand2 gate13( .a(G9), .b(G10), .O(G278) );
nand2 gate14( .a(G11), .b(G12), .O(G281) );
nand2 gate15( .a(G13), .b(G14), .O(G284) );
nand2 gate16( .a(G15), .b(G16), .O(G287) );

  xor2  gate813(.a(G18), .b(G17), .O(gate17inter0));
  nand2 gate814(.a(gate17inter0), .b(s_38), .O(gate17inter1));
  and2  gate815(.a(G18), .b(G17), .O(gate17inter2));
  inv1  gate816(.a(s_38), .O(gate17inter3));
  inv1  gate817(.a(s_39), .O(gate17inter4));
  nand2 gate818(.a(gate17inter4), .b(gate17inter3), .O(gate17inter5));
  nor2  gate819(.a(gate17inter5), .b(gate17inter2), .O(gate17inter6));
  inv1  gate820(.a(G17), .O(gate17inter7));
  inv1  gate821(.a(G18), .O(gate17inter8));
  nand2 gate822(.a(gate17inter8), .b(gate17inter7), .O(gate17inter9));
  nand2 gate823(.a(s_39), .b(gate17inter3), .O(gate17inter10));
  nor2  gate824(.a(gate17inter10), .b(gate17inter9), .O(gate17inter11));
  nor2  gate825(.a(gate17inter11), .b(gate17inter6), .O(gate17inter12));
  nand2 gate826(.a(gate17inter12), .b(gate17inter1), .O(G290));

  xor2  gate1023(.a(G20), .b(G19), .O(gate18inter0));
  nand2 gate1024(.a(gate18inter0), .b(s_68), .O(gate18inter1));
  and2  gate1025(.a(G20), .b(G19), .O(gate18inter2));
  inv1  gate1026(.a(s_68), .O(gate18inter3));
  inv1  gate1027(.a(s_69), .O(gate18inter4));
  nand2 gate1028(.a(gate18inter4), .b(gate18inter3), .O(gate18inter5));
  nor2  gate1029(.a(gate18inter5), .b(gate18inter2), .O(gate18inter6));
  inv1  gate1030(.a(G19), .O(gate18inter7));
  inv1  gate1031(.a(G20), .O(gate18inter8));
  nand2 gate1032(.a(gate18inter8), .b(gate18inter7), .O(gate18inter9));
  nand2 gate1033(.a(s_69), .b(gate18inter3), .O(gate18inter10));
  nor2  gate1034(.a(gate18inter10), .b(gate18inter9), .O(gate18inter11));
  nor2  gate1035(.a(gate18inter11), .b(gate18inter6), .O(gate18inter12));
  nand2 gate1036(.a(gate18inter12), .b(gate18inter1), .O(G293));
nand2 gate19( .a(G21), .b(G22), .O(G296) );
nand2 gate20( .a(G23), .b(G24), .O(G299) );
nand2 gate21( .a(G25), .b(G26), .O(G302) );
nand2 gate22( .a(G27), .b(G28), .O(G305) );
nand2 gate23( .a(G29), .b(G30), .O(G308) );
nand2 gate24( .a(G31), .b(G32), .O(G311) );
nand2 gate25( .a(G1), .b(G5), .O(G314) );
nand2 gate26( .a(G9), .b(G13), .O(G317) );
nand2 gate27( .a(G2), .b(G6), .O(G320) );
nand2 gate28( .a(G10), .b(G14), .O(G323) );

  xor2  gate2185(.a(G7), .b(G3), .O(gate29inter0));
  nand2 gate2186(.a(gate29inter0), .b(s_234), .O(gate29inter1));
  and2  gate2187(.a(G7), .b(G3), .O(gate29inter2));
  inv1  gate2188(.a(s_234), .O(gate29inter3));
  inv1  gate2189(.a(s_235), .O(gate29inter4));
  nand2 gate2190(.a(gate29inter4), .b(gate29inter3), .O(gate29inter5));
  nor2  gate2191(.a(gate29inter5), .b(gate29inter2), .O(gate29inter6));
  inv1  gate2192(.a(G3), .O(gate29inter7));
  inv1  gate2193(.a(G7), .O(gate29inter8));
  nand2 gate2194(.a(gate29inter8), .b(gate29inter7), .O(gate29inter9));
  nand2 gate2195(.a(s_235), .b(gate29inter3), .O(gate29inter10));
  nor2  gate2196(.a(gate29inter10), .b(gate29inter9), .O(gate29inter11));
  nor2  gate2197(.a(gate29inter11), .b(gate29inter6), .O(gate29inter12));
  nand2 gate2198(.a(gate29inter12), .b(gate29inter1), .O(G326));
nand2 gate30( .a(G11), .b(G15), .O(G329) );

  xor2  gate1709(.a(G8), .b(G4), .O(gate31inter0));
  nand2 gate1710(.a(gate31inter0), .b(s_166), .O(gate31inter1));
  and2  gate1711(.a(G8), .b(G4), .O(gate31inter2));
  inv1  gate1712(.a(s_166), .O(gate31inter3));
  inv1  gate1713(.a(s_167), .O(gate31inter4));
  nand2 gate1714(.a(gate31inter4), .b(gate31inter3), .O(gate31inter5));
  nor2  gate1715(.a(gate31inter5), .b(gate31inter2), .O(gate31inter6));
  inv1  gate1716(.a(G4), .O(gate31inter7));
  inv1  gate1717(.a(G8), .O(gate31inter8));
  nand2 gate1718(.a(gate31inter8), .b(gate31inter7), .O(gate31inter9));
  nand2 gate1719(.a(s_167), .b(gate31inter3), .O(gate31inter10));
  nor2  gate1720(.a(gate31inter10), .b(gate31inter9), .O(gate31inter11));
  nor2  gate1721(.a(gate31inter11), .b(gate31inter6), .O(gate31inter12));
  nand2 gate1722(.a(gate31inter12), .b(gate31inter1), .O(G332));

  xor2  gate1275(.a(G16), .b(G12), .O(gate32inter0));
  nand2 gate1276(.a(gate32inter0), .b(s_104), .O(gate32inter1));
  and2  gate1277(.a(G16), .b(G12), .O(gate32inter2));
  inv1  gate1278(.a(s_104), .O(gate32inter3));
  inv1  gate1279(.a(s_105), .O(gate32inter4));
  nand2 gate1280(.a(gate32inter4), .b(gate32inter3), .O(gate32inter5));
  nor2  gate1281(.a(gate32inter5), .b(gate32inter2), .O(gate32inter6));
  inv1  gate1282(.a(G12), .O(gate32inter7));
  inv1  gate1283(.a(G16), .O(gate32inter8));
  nand2 gate1284(.a(gate32inter8), .b(gate32inter7), .O(gate32inter9));
  nand2 gate1285(.a(s_105), .b(gate32inter3), .O(gate32inter10));
  nor2  gate1286(.a(gate32inter10), .b(gate32inter9), .O(gate32inter11));
  nor2  gate1287(.a(gate32inter11), .b(gate32inter6), .O(gate32inter12));
  nand2 gate1288(.a(gate32inter12), .b(gate32inter1), .O(G335));
nand2 gate33( .a(G17), .b(G21), .O(G338) );
nand2 gate34( .a(G25), .b(G29), .O(G341) );
nand2 gate35( .a(G18), .b(G22), .O(G344) );
nand2 gate36( .a(G26), .b(G30), .O(G347) );

  xor2  gate2143(.a(G23), .b(G19), .O(gate37inter0));
  nand2 gate2144(.a(gate37inter0), .b(s_228), .O(gate37inter1));
  and2  gate2145(.a(G23), .b(G19), .O(gate37inter2));
  inv1  gate2146(.a(s_228), .O(gate37inter3));
  inv1  gate2147(.a(s_229), .O(gate37inter4));
  nand2 gate2148(.a(gate37inter4), .b(gate37inter3), .O(gate37inter5));
  nor2  gate2149(.a(gate37inter5), .b(gate37inter2), .O(gate37inter6));
  inv1  gate2150(.a(G19), .O(gate37inter7));
  inv1  gate2151(.a(G23), .O(gate37inter8));
  nand2 gate2152(.a(gate37inter8), .b(gate37inter7), .O(gate37inter9));
  nand2 gate2153(.a(s_229), .b(gate37inter3), .O(gate37inter10));
  nor2  gate2154(.a(gate37inter10), .b(gate37inter9), .O(gate37inter11));
  nor2  gate2155(.a(gate37inter11), .b(gate37inter6), .O(gate37inter12));
  nand2 gate2156(.a(gate37inter12), .b(gate37inter1), .O(G350));

  xor2  gate2241(.a(G31), .b(G27), .O(gate38inter0));
  nand2 gate2242(.a(gate38inter0), .b(s_242), .O(gate38inter1));
  and2  gate2243(.a(G31), .b(G27), .O(gate38inter2));
  inv1  gate2244(.a(s_242), .O(gate38inter3));
  inv1  gate2245(.a(s_243), .O(gate38inter4));
  nand2 gate2246(.a(gate38inter4), .b(gate38inter3), .O(gate38inter5));
  nor2  gate2247(.a(gate38inter5), .b(gate38inter2), .O(gate38inter6));
  inv1  gate2248(.a(G27), .O(gate38inter7));
  inv1  gate2249(.a(G31), .O(gate38inter8));
  nand2 gate2250(.a(gate38inter8), .b(gate38inter7), .O(gate38inter9));
  nand2 gate2251(.a(s_243), .b(gate38inter3), .O(gate38inter10));
  nor2  gate2252(.a(gate38inter10), .b(gate38inter9), .O(gate38inter11));
  nor2  gate2253(.a(gate38inter11), .b(gate38inter6), .O(gate38inter12));
  nand2 gate2254(.a(gate38inter12), .b(gate38inter1), .O(G353));

  xor2  gate1121(.a(G24), .b(G20), .O(gate39inter0));
  nand2 gate1122(.a(gate39inter0), .b(s_82), .O(gate39inter1));
  and2  gate1123(.a(G24), .b(G20), .O(gate39inter2));
  inv1  gate1124(.a(s_82), .O(gate39inter3));
  inv1  gate1125(.a(s_83), .O(gate39inter4));
  nand2 gate1126(.a(gate39inter4), .b(gate39inter3), .O(gate39inter5));
  nor2  gate1127(.a(gate39inter5), .b(gate39inter2), .O(gate39inter6));
  inv1  gate1128(.a(G20), .O(gate39inter7));
  inv1  gate1129(.a(G24), .O(gate39inter8));
  nand2 gate1130(.a(gate39inter8), .b(gate39inter7), .O(gate39inter9));
  nand2 gate1131(.a(s_83), .b(gate39inter3), .O(gate39inter10));
  nor2  gate1132(.a(gate39inter10), .b(gate39inter9), .O(gate39inter11));
  nor2  gate1133(.a(gate39inter11), .b(gate39inter6), .O(gate39inter12));
  nand2 gate1134(.a(gate39inter12), .b(gate39inter1), .O(G356));
nand2 gate40( .a(G28), .b(G32), .O(G359) );

  xor2  gate2381(.a(G266), .b(G1), .O(gate41inter0));
  nand2 gate2382(.a(gate41inter0), .b(s_262), .O(gate41inter1));
  and2  gate2383(.a(G266), .b(G1), .O(gate41inter2));
  inv1  gate2384(.a(s_262), .O(gate41inter3));
  inv1  gate2385(.a(s_263), .O(gate41inter4));
  nand2 gate2386(.a(gate41inter4), .b(gate41inter3), .O(gate41inter5));
  nor2  gate2387(.a(gate41inter5), .b(gate41inter2), .O(gate41inter6));
  inv1  gate2388(.a(G1), .O(gate41inter7));
  inv1  gate2389(.a(G266), .O(gate41inter8));
  nand2 gate2390(.a(gate41inter8), .b(gate41inter7), .O(gate41inter9));
  nand2 gate2391(.a(s_263), .b(gate41inter3), .O(gate41inter10));
  nor2  gate2392(.a(gate41inter10), .b(gate41inter9), .O(gate41inter11));
  nor2  gate2393(.a(gate41inter11), .b(gate41inter6), .O(gate41inter12));
  nand2 gate2394(.a(gate41inter12), .b(gate41inter1), .O(G362));
nand2 gate42( .a(G2), .b(G266), .O(G363) );

  xor2  gate1485(.a(G269), .b(G3), .O(gate43inter0));
  nand2 gate1486(.a(gate43inter0), .b(s_134), .O(gate43inter1));
  and2  gate1487(.a(G269), .b(G3), .O(gate43inter2));
  inv1  gate1488(.a(s_134), .O(gate43inter3));
  inv1  gate1489(.a(s_135), .O(gate43inter4));
  nand2 gate1490(.a(gate43inter4), .b(gate43inter3), .O(gate43inter5));
  nor2  gate1491(.a(gate43inter5), .b(gate43inter2), .O(gate43inter6));
  inv1  gate1492(.a(G3), .O(gate43inter7));
  inv1  gate1493(.a(G269), .O(gate43inter8));
  nand2 gate1494(.a(gate43inter8), .b(gate43inter7), .O(gate43inter9));
  nand2 gate1495(.a(s_135), .b(gate43inter3), .O(gate43inter10));
  nor2  gate1496(.a(gate43inter10), .b(gate43inter9), .O(gate43inter11));
  nor2  gate1497(.a(gate43inter11), .b(gate43inter6), .O(gate43inter12));
  nand2 gate1498(.a(gate43inter12), .b(gate43inter1), .O(G364));
nand2 gate44( .a(G4), .b(G269), .O(G365) );
nand2 gate45( .a(G5), .b(G272), .O(G366) );

  xor2  gate729(.a(G272), .b(G6), .O(gate46inter0));
  nand2 gate730(.a(gate46inter0), .b(s_26), .O(gate46inter1));
  and2  gate731(.a(G272), .b(G6), .O(gate46inter2));
  inv1  gate732(.a(s_26), .O(gate46inter3));
  inv1  gate733(.a(s_27), .O(gate46inter4));
  nand2 gate734(.a(gate46inter4), .b(gate46inter3), .O(gate46inter5));
  nor2  gate735(.a(gate46inter5), .b(gate46inter2), .O(gate46inter6));
  inv1  gate736(.a(G6), .O(gate46inter7));
  inv1  gate737(.a(G272), .O(gate46inter8));
  nand2 gate738(.a(gate46inter8), .b(gate46inter7), .O(gate46inter9));
  nand2 gate739(.a(s_27), .b(gate46inter3), .O(gate46inter10));
  nor2  gate740(.a(gate46inter10), .b(gate46inter9), .O(gate46inter11));
  nor2  gate741(.a(gate46inter11), .b(gate46inter6), .O(gate46inter12));
  nand2 gate742(.a(gate46inter12), .b(gate46inter1), .O(G367));
nand2 gate47( .a(G7), .b(G275), .O(G368) );
nand2 gate48( .a(G8), .b(G275), .O(G369) );

  xor2  gate2003(.a(G278), .b(G9), .O(gate49inter0));
  nand2 gate2004(.a(gate49inter0), .b(s_208), .O(gate49inter1));
  and2  gate2005(.a(G278), .b(G9), .O(gate49inter2));
  inv1  gate2006(.a(s_208), .O(gate49inter3));
  inv1  gate2007(.a(s_209), .O(gate49inter4));
  nand2 gate2008(.a(gate49inter4), .b(gate49inter3), .O(gate49inter5));
  nor2  gate2009(.a(gate49inter5), .b(gate49inter2), .O(gate49inter6));
  inv1  gate2010(.a(G9), .O(gate49inter7));
  inv1  gate2011(.a(G278), .O(gate49inter8));
  nand2 gate2012(.a(gate49inter8), .b(gate49inter7), .O(gate49inter9));
  nand2 gate2013(.a(s_209), .b(gate49inter3), .O(gate49inter10));
  nor2  gate2014(.a(gate49inter10), .b(gate49inter9), .O(gate49inter11));
  nor2  gate2015(.a(gate49inter11), .b(gate49inter6), .O(gate49inter12));
  nand2 gate2016(.a(gate49inter12), .b(gate49inter1), .O(G370));
nand2 gate50( .a(G10), .b(G278), .O(G371) );
nand2 gate51( .a(G11), .b(G281), .O(G372) );

  xor2  gate1191(.a(G281), .b(G12), .O(gate52inter0));
  nand2 gate1192(.a(gate52inter0), .b(s_92), .O(gate52inter1));
  and2  gate1193(.a(G281), .b(G12), .O(gate52inter2));
  inv1  gate1194(.a(s_92), .O(gate52inter3));
  inv1  gate1195(.a(s_93), .O(gate52inter4));
  nand2 gate1196(.a(gate52inter4), .b(gate52inter3), .O(gate52inter5));
  nor2  gate1197(.a(gate52inter5), .b(gate52inter2), .O(gate52inter6));
  inv1  gate1198(.a(G12), .O(gate52inter7));
  inv1  gate1199(.a(G281), .O(gate52inter8));
  nand2 gate1200(.a(gate52inter8), .b(gate52inter7), .O(gate52inter9));
  nand2 gate1201(.a(s_93), .b(gate52inter3), .O(gate52inter10));
  nor2  gate1202(.a(gate52inter10), .b(gate52inter9), .O(gate52inter11));
  nor2  gate1203(.a(gate52inter11), .b(gate52inter6), .O(gate52inter12));
  nand2 gate1204(.a(gate52inter12), .b(gate52inter1), .O(G373));
nand2 gate53( .a(G13), .b(G284), .O(G374) );

  xor2  gate1639(.a(G284), .b(G14), .O(gate54inter0));
  nand2 gate1640(.a(gate54inter0), .b(s_156), .O(gate54inter1));
  and2  gate1641(.a(G284), .b(G14), .O(gate54inter2));
  inv1  gate1642(.a(s_156), .O(gate54inter3));
  inv1  gate1643(.a(s_157), .O(gate54inter4));
  nand2 gate1644(.a(gate54inter4), .b(gate54inter3), .O(gate54inter5));
  nor2  gate1645(.a(gate54inter5), .b(gate54inter2), .O(gate54inter6));
  inv1  gate1646(.a(G14), .O(gate54inter7));
  inv1  gate1647(.a(G284), .O(gate54inter8));
  nand2 gate1648(.a(gate54inter8), .b(gate54inter7), .O(gate54inter9));
  nand2 gate1649(.a(s_157), .b(gate54inter3), .O(gate54inter10));
  nor2  gate1650(.a(gate54inter10), .b(gate54inter9), .O(gate54inter11));
  nor2  gate1651(.a(gate54inter11), .b(gate54inter6), .O(gate54inter12));
  nand2 gate1652(.a(gate54inter12), .b(gate54inter1), .O(G375));

  xor2  gate1359(.a(G287), .b(G15), .O(gate55inter0));
  nand2 gate1360(.a(gate55inter0), .b(s_116), .O(gate55inter1));
  and2  gate1361(.a(G287), .b(G15), .O(gate55inter2));
  inv1  gate1362(.a(s_116), .O(gate55inter3));
  inv1  gate1363(.a(s_117), .O(gate55inter4));
  nand2 gate1364(.a(gate55inter4), .b(gate55inter3), .O(gate55inter5));
  nor2  gate1365(.a(gate55inter5), .b(gate55inter2), .O(gate55inter6));
  inv1  gate1366(.a(G15), .O(gate55inter7));
  inv1  gate1367(.a(G287), .O(gate55inter8));
  nand2 gate1368(.a(gate55inter8), .b(gate55inter7), .O(gate55inter9));
  nand2 gate1369(.a(s_117), .b(gate55inter3), .O(gate55inter10));
  nor2  gate1370(.a(gate55inter10), .b(gate55inter9), .O(gate55inter11));
  nor2  gate1371(.a(gate55inter11), .b(gate55inter6), .O(gate55inter12));
  nand2 gate1372(.a(gate55inter12), .b(gate55inter1), .O(G376));

  xor2  gate1345(.a(G287), .b(G16), .O(gate56inter0));
  nand2 gate1346(.a(gate56inter0), .b(s_114), .O(gate56inter1));
  and2  gate1347(.a(G287), .b(G16), .O(gate56inter2));
  inv1  gate1348(.a(s_114), .O(gate56inter3));
  inv1  gate1349(.a(s_115), .O(gate56inter4));
  nand2 gate1350(.a(gate56inter4), .b(gate56inter3), .O(gate56inter5));
  nor2  gate1351(.a(gate56inter5), .b(gate56inter2), .O(gate56inter6));
  inv1  gate1352(.a(G16), .O(gate56inter7));
  inv1  gate1353(.a(G287), .O(gate56inter8));
  nand2 gate1354(.a(gate56inter8), .b(gate56inter7), .O(gate56inter9));
  nand2 gate1355(.a(s_115), .b(gate56inter3), .O(gate56inter10));
  nor2  gate1356(.a(gate56inter10), .b(gate56inter9), .O(gate56inter11));
  nor2  gate1357(.a(gate56inter11), .b(gate56inter6), .O(gate56inter12));
  nand2 gate1358(.a(gate56inter12), .b(gate56inter1), .O(G377));
nand2 gate57( .a(G17), .b(G290), .O(G378) );

  xor2  gate561(.a(G290), .b(G18), .O(gate58inter0));
  nand2 gate562(.a(gate58inter0), .b(s_2), .O(gate58inter1));
  and2  gate563(.a(G290), .b(G18), .O(gate58inter2));
  inv1  gate564(.a(s_2), .O(gate58inter3));
  inv1  gate565(.a(s_3), .O(gate58inter4));
  nand2 gate566(.a(gate58inter4), .b(gate58inter3), .O(gate58inter5));
  nor2  gate567(.a(gate58inter5), .b(gate58inter2), .O(gate58inter6));
  inv1  gate568(.a(G18), .O(gate58inter7));
  inv1  gate569(.a(G290), .O(gate58inter8));
  nand2 gate570(.a(gate58inter8), .b(gate58inter7), .O(gate58inter9));
  nand2 gate571(.a(s_3), .b(gate58inter3), .O(gate58inter10));
  nor2  gate572(.a(gate58inter10), .b(gate58inter9), .O(gate58inter11));
  nor2  gate573(.a(gate58inter11), .b(gate58inter6), .O(gate58inter12));
  nand2 gate574(.a(gate58inter12), .b(gate58inter1), .O(G379));

  xor2  gate799(.a(G293), .b(G19), .O(gate59inter0));
  nand2 gate800(.a(gate59inter0), .b(s_36), .O(gate59inter1));
  and2  gate801(.a(G293), .b(G19), .O(gate59inter2));
  inv1  gate802(.a(s_36), .O(gate59inter3));
  inv1  gate803(.a(s_37), .O(gate59inter4));
  nand2 gate804(.a(gate59inter4), .b(gate59inter3), .O(gate59inter5));
  nor2  gate805(.a(gate59inter5), .b(gate59inter2), .O(gate59inter6));
  inv1  gate806(.a(G19), .O(gate59inter7));
  inv1  gate807(.a(G293), .O(gate59inter8));
  nand2 gate808(.a(gate59inter8), .b(gate59inter7), .O(gate59inter9));
  nand2 gate809(.a(s_37), .b(gate59inter3), .O(gate59inter10));
  nor2  gate810(.a(gate59inter10), .b(gate59inter9), .O(gate59inter11));
  nor2  gate811(.a(gate59inter11), .b(gate59inter6), .O(gate59inter12));
  nand2 gate812(.a(gate59inter12), .b(gate59inter1), .O(G380));
nand2 gate60( .a(G20), .b(G293), .O(G381) );
nand2 gate61( .a(G21), .b(G296), .O(G382) );
nand2 gate62( .a(G22), .b(G296), .O(G383) );

  xor2  gate771(.a(G299), .b(G23), .O(gate63inter0));
  nand2 gate772(.a(gate63inter0), .b(s_32), .O(gate63inter1));
  and2  gate773(.a(G299), .b(G23), .O(gate63inter2));
  inv1  gate774(.a(s_32), .O(gate63inter3));
  inv1  gate775(.a(s_33), .O(gate63inter4));
  nand2 gate776(.a(gate63inter4), .b(gate63inter3), .O(gate63inter5));
  nor2  gate777(.a(gate63inter5), .b(gate63inter2), .O(gate63inter6));
  inv1  gate778(.a(G23), .O(gate63inter7));
  inv1  gate779(.a(G299), .O(gate63inter8));
  nand2 gate780(.a(gate63inter8), .b(gate63inter7), .O(gate63inter9));
  nand2 gate781(.a(s_33), .b(gate63inter3), .O(gate63inter10));
  nor2  gate782(.a(gate63inter10), .b(gate63inter9), .O(gate63inter11));
  nor2  gate783(.a(gate63inter11), .b(gate63inter6), .O(gate63inter12));
  nand2 gate784(.a(gate63inter12), .b(gate63inter1), .O(G384));
nand2 gate64( .a(G24), .b(G299), .O(G385) );
nand2 gate65( .a(G25), .b(G302), .O(G386) );

  xor2  gate1317(.a(G302), .b(G26), .O(gate66inter0));
  nand2 gate1318(.a(gate66inter0), .b(s_110), .O(gate66inter1));
  and2  gate1319(.a(G302), .b(G26), .O(gate66inter2));
  inv1  gate1320(.a(s_110), .O(gate66inter3));
  inv1  gate1321(.a(s_111), .O(gate66inter4));
  nand2 gate1322(.a(gate66inter4), .b(gate66inter3), .O(gate66inter5));
  nor2  gate1323(.a(gate66inter5), .b(gate66inter2), .O(gate66inter6));
  inv1  gate1324(.a(G26), .O(gate66inter7));
  inv1  gate1325(.a(G302), .O(gate66inter8));
  nand2 gate1326(.a(gate66inter8), .b(gate66inter7), .O(gate66inter9));
  nand2 gate1327(.a(s_111), .b(gate66inter3), .O(gate66inter10));
  nor2  gate1328(.a(gate66inter10), .b(gate66inter9), .O(gate66inter11));
  nor2  gate1329(.a(gate66inter11), .b(gate66inter6), .O(gate66inter12));
  nand2 gate1330(.a(gate66inter12), .b(gate66inter1), .O(G387));
nand2 gate67( .a(G27), .b(G305), .O(G388) );
nand2 gate68( .a(G28), .b(G305), .O(G389) );
nand2 gate69( .a(G29), .b(G308), .O(G390) );

  xor2  gate827(.a(G308), .b(G30), .O(gate70inter0));
  nand2 gate828(.a(gate70inter0), .b(s_40), .O(gate70inter1));
  and2  gate829(.a(G308), .b(G30), .O(gate70inter2));
  inv1  gate830(.a(s_40), .O(gate70inter3));
  inv1  gate831(.a(s_41), .O(gate70inter4));
  nand2 gate832(.a(gate70inter4), .b(gate70inter3), .O(gate70inter5));
  nor2  gate833(.a(gate70inter5), .b(gate70inter2), .O(gate70inter6));
  inv1  gate834(.a(G30), .O(gate70inter7));
  inv1  gate835(.a(G308), .O(gate70inter8));
  nand2 gate836(.a(gate70inter8), .b(gate70inter7), .O(gate70inter9));
  nand2 gate837(.a(s_41), .b(gate70inter3), .O(gate70inter10));
  nor2  gate838(.a(gate70inter10), .b(gate70inter9), .O(gate70inter11));
  nor2  gate839(.a(gate70inter11), .b(gate70inter6), .O(gate70inter12));
  nand2 gate840(.a(gate70inter12), .b(gate70inter1), .O(G391));
nand2 gate71( .a(G31), .b(G311), .O(G392) );
nand2 gate72( .a(G32), .b(G311), .O(G393) );

  xor2  gate855(.a(G314), .b(G1), .O(gate73inter0));
  nand2 gate856(.a(gate73inter0), .b(s_44), .O(gate73inter1));
  and2  gate857(.a(G314), .b(G1), .O(gate73inter2));
  inv1  gate858(.a(s_44), .O(gate73inter3));
  inv1  gate859(.a(s_45), .O(gate73inter4));
  nand2 gate860(.a(gate73inter4), .b(gate73inter3), .O(gate73inter5));
  nor2  gate861(.a(gate73inter5), .b(gate73inter2), .O(gate73inter6));
  inv1  gate862(.a(G1), .O(gate73inter7));
  inv1  gate863(.a(G314), .O(gate73inter8));
  nand2 gate864(.a(gate73inter8), .b(gate73inter7), .O(gate73inter9));
  nand2 gate865(.a(s_45), .b(gate73inter3), .O(gate73inter10));
  nor2  gate866(.a(gate73inter10), .b(gate73inter9), .O(gate73inter11));
  nor2  gate867(.a(gate73inter11), .b(gate73inter6), .O(gate73inter12));
  nand2 gate868(.a(gate73inter12), .b(gate73inter1), .O(G394));
nand2 gate74( .a(G5), .b(G314), .O(G395) );
nand2 gate75( .a(G9), .b(G317), .O(G396) );
nand2 gate76( .a(G13), .b(G317), .O(G397) );
nand2 gate77( .a(G2), .b(G320), .O(G398) );
nand2 gate78( .a(G6), .b(G320), .O(G399) );
nand2 gate79( .a(G10), .b(G323), .O(G400) );

  xor2  gate2129(.a(G323), .b(G14), .O(gate80inter0));
  nand2 gate2130(.a(gate80inter0), .b(s_226), .O(gate80inter1));
  and2  gate2131(.a(G323), .b(G14), .O(gate80inter2));
  inv1  gate2132(.a(s_226), .O(gate80inter3));
  inv1  gate2133(.a(s_227), .O(gate80inter4));
  nand2 gate2134(.a(gate80inter4), .b(gate80inter3), .O(gate80inter5));
  nor2  gate2135(.a(gate80inter5), .b(gate80inter2), .O(gate80inter6));
  inv1  gate2136(.a(G14), .O(gate80inter7));
  inv1  gate2137(.a(G323), .O(gate80inter8));
  nand2 gate2138(.a(gate80inter8), .b(gate80inter7), .O(gate80inter9));
  nand2 gate2139(.a(s_227), .b(gate80inter3), .O(gate80inter10));
  nor2  gate2140(.a(gate80inter10), .b(gate80inter9), .O(gate80inter11));
  nor2  gate2141(.a(gate80inter11), .b(gate80inter6), .O(gate80inter12));
  nand2 gate2142(.a(gate80inter12), .b(gate80inter1), .O(G401));
nand2 gate81( .a(G3), .b(G326), .O(G402) );
nand2 gate82( .a(G7), .b(G326), .O(G403) );

  xor2  gate1667(.a(G329), .b(G11), .O(gate83inter0));
  nand2 gate1668(.a(gate83inter0), .b(s_160), .O(gate83inter1));
  and2  gate1669(.a(G329), .b(G11), .O(gate83inter2));
  inv1  gate1670(.a(s_160), .O(gate83inter3));
  inv1  gate1671(.a(s_161), .O(gate83inter4));
  nand2 gate1672(.a(gate83inter4), .b(gate83inter3), .O(gate83inter5));
  nor2  gate1673(.a(gate83inter5), .b(gate83inter2), .O(gate83inter6));
  inv1  gate1674(.a(G11), .O(gate83inter7));
  inv1  gate1675(.a(G329), .O(gate83inter8));
  nand2 gate1676(.a(gate83inter8), .b(gate83inter7), .O(gate83inter9));
  nand2 gate1677(.a(s_161), .b(gate83inter3), .O(gate83inter10));
  nor2  gate1678(.a(gate83inter10), .b(gate83inter9), .O(gate83inter11));
  nor2  gate1679(.a(gate83inter11), .b(gate83inter6), .O(gate83inter12));
  nand2 gate1680(.a(gate83inter12), .b(gate83inter1), .O(G404));
nand2 gate84( .a(G15), .b(G329), .O(G405) );
nand2 gate85( .a(G4), .b(G332), .O(G406) );

  xor2  gate1009(.a(G332), .b(G8), .O(gate86inter0));
  nand2 gate1010(.a(gate86inter0), .b(s_66), .O(gate86inter1));
  and2  gate1011(.a(G332), .b(G8), .O(gate86inter2));
  inv1  gate1012(.a(s_66), .O(gate86inter3));
  inv1  gate1013(.a(s_67), .O(gate86inter4));
  nand2 gate1014(.a(gate86inter4), .b(gate86inter3), .O(gate86inter5));
  nor2  gate1015(.a(gate86inter5), .b(gate86inter2), .O(gate86inter6));
  inv1  gate1016(.a(G8), .O(gate86inter7));
  inv1  gate1017(.a(G332), .O(gate86inter8));
  nand2 gate1018(.a(gate86inter8), .b(gate86inter7), .O(gate86inter9));
  nand2 gate1019(.a(s_67), .b(gate86inter3), .O(gate86inter10));
  nor2  gate1020(.a(gate86inter10), .b(gate86inter9), .O(gate86inter11));
  nor2  gate1021(.a(gate86inter11), .b(gate86inter6), .O(gate86inter12));
  nand2 gate1022(.a(gate86inter12), .b(gate86inter1), .O(G407));

  xor2  gate1695(.a(G335), .b(G12), .O(gate87inter0));
  nand2 gate1696(.a(gate87inter0), .b(s_164), .O(gate87inter1));
  and2  gate1697(.a(G335), .b(G12), .O(gate87inter2));
  inv1  gate1698(.a(s_164), .O(gate87inter3));
  inv1  gate1699(.a(s_165), .O(gate87inter4));
  nand2 gate1700(.a(gate87inter4), .b(gate87inter3), .O(gate87inter5));
  nor2  gate1701(.a(gate87inter5), .b(gate87inter2), .O(gate87inter6));
  inv1  gate1702(.a(G12), .O(gate87inter7));
  inv1  gate1703(.a(G335), .O(gate87inter8));
  nand2 gate1704(.a(gate87inter8), .b(gate87inter7), .O(gate87inter9));
  nand2 gate1705(.a(s_165), .b(gate87inter3), .O(gate87inter10));
  nor2  gate1706(.a(gate87inter10), .b(gate87inter9), .O(gate87inter11));
  nor2  gate1707(.a(gate87inter11), .b(gate87inter6), .O(gate87inter12));
  nand2 gate1708(.a(gate87inter12), .b(gate87inter1), .O(G408));
nand2 gate88( .a(G16), .b(G335), .O(G409) );
nand2 gate89( .a(G17), .b(G338), .O(G410) );
nand2 gate90( .a(G21), .b(G338), .O(G411) );
nand2 gate91( .a(G25), .b(G341), .O(G412) );
nand2 gate92( .a(G29), .b(G341), .O(G413) );
nand2 gate93( .a(G18), .b(G344), .O(G414) );

  xor2  gate1415(.a(G344), .b(G22), .O(gate94inter0));
  nand2 gate1416(.a(gate94inter0), .b(s_124), .O(gate94inter1));
  and2  gate1417(.a(G344), .b(G22), .O(gate94inter2));
  inv1  gate1418(.a(s_124), .O(gate94inter3));
  inv1  gate1419(.a(s_125), .O(gate94inter4));
  nand2 gate1420(.a(gate94inter4), .b(gate94inter3), .O(gate94inter5));
  nor2  gate1421(.a(gate94inter5), .b(gate94inter2), .O(gate94inter6));
  inv1  gate1422(.a(G22), .O(gate94inter7));
  inv1  gate1423(.a(G344), .O(gate94inter8));
  nand2 gate1424(.a(gate94inter8), .b(gate94inter7), .O(gate94inter9));
  nand2 gate1425(.a(s_125), .b(gate94inter3), .O(gate94inter10));
  nor2  gate1426(.a(gate94inter10), .b(gate94inter9), .O(gate94inter11));
  nor2  gate1427(.a(gate94inter11), .b(gate94inter6), .O(gate94inter12));
  nand2 gate1428(.a(gate94inter12), .b(gate94inter1), .O(G415));
nand2 gate95( .a(G26), .b(G347), .O(G416) );
nand2 gate96( .a(G30), .b(G347), .O(G417) );
nand2 gate97( .a(G19), .b(G350), .O(G418) );
nand2 gate98( .a(G23), .b(G350), .O(G419) );
nand2 gate99( .a(G27), .b(G353), .O(G420) );
nand2 gate100( .a(G31), .b(G353), .O(G421) );
nand2 gate101( .a(G20), .b(G356), .O(G422) );
nand2 gate102( .a(G24), .b(G356), .O(G423) );
nand2 gate103( .a(G28), .b(G359), .O(G424) );
nand2 gate104( .a(G32), .b(G359), .O(G425) );
nand2 gate105( .a(G362), .b(G363), .O(G426) );

  xor2  gate1877(.a(G365), .b(G364), .O(gate106inter0));
  nand2 gate1878(.a(gate106inter0), .b(s_190), .O(gate106inter1));
  and2  gate1879(.a(G365), .b(G364), .O(gate106inter2));
  inv1  gate1880(.a(s_190), .O(gate106inter3));
  inv1  gate1881(.a(s_191), .O(gate106inter4));
  nand2 gate1882(.a(gate106inter4), .b(gate106inter3), .O(gate106inter5));
  nor2  gate1883(.a(gate106inter5), .b(gate106inter2), .O(gate106inter6));
  inv1  gate1884(.a(G364), .O(gate106inter7));
  inv1  gate1885(.a(G365), .O(gate106inter8));
  nand2 gate1886(.a(gate106inter8), .b(gate106inter7), .O(gate106inter9));
  nand2 gate1887(.a(s_191), .b(gate106inter3), .O(gate106inter10));
  nor2  gate1888(.a(gate106inter10), .b(gate106inter9), .O(gate106inter11));
  nor2  gate1889(.a(gate106inter11), .b(gate106inter6), .O(gate106inter12));
  nand2 gate1890(.a(gate106inter12), .b(gate106inter1), .O(G429));
nand2 gate107( .a(G366), .b(G367), .O(G432) );
nand2 gate108( .a(G368), .b(G369), .O(G435) );

  xor2  gate1037(.a(G371), .b(G370), .O(gate109inter0));
  nand2 gate1038(.a(gate109inter0), .b(s_70), .O(gate109inter1));
  and2  gate1039(.a(G371), .b(G370), .O(gate109inter2));
  inv1  gate1040(.a(s_70), .O(gate109inter3));
  inv1  gate1041(.a(s_71), .O(gate109inter4));
  nand2 gate1042(.a(gate109inter4), .b(gate109inter3), .O(gate109inter5));
  nor2  gate1043(.a(gate109inter5), .b(gate109inter2), .O(gate109inter6));
  inv1  gate1044(.a(G370), .O(gate109inter7));
  inv1  gate1045(.a(G371), .O(gate109inter8));
  nand2 gate1046(.a(gate109inter8), .b(gate109inter7), .O(gate109inter9));
  nand2 gate1047(.a(s_71), .b(gate109inter3), .O(gate109inter10));
  nor2  gate1048(.a(gate109inter10), .b(gate109inter9), .O(gate109inter11));
  nor2  gate1049(.a(gate109inter11), .b(gate109inter6), .O(gate109inter12));
  nand2 gate1050(.a(gate109inter12), .b(gate109inter1), .O(G438));

  xor2  gate1135(.a(G373), .b(G372), .O(gate110inter0));
  nand2 gate1136(.a(gate110inter0), .b(s_84), .O(gate110inter1));
  and2  gate1137(.a(G373), .b(G372), .O(gate110inter2));
  inv1  gate1138(.a(s_84), .O(gate110inter3));
  inv1  gate1139(.a(s_85), .O(gate110inter4));
  nand2 gate1140(.a(gate110inter4), .b(gate110inter3), .O(gate110inter5));
  nor2  gate1141(.a(gate110inter5), .b(gate110inter2), .O(gate110inter6));
  inv1  gate1142(.a(G372), .O(gate110inter7));
  inv1  gate1143(.a(G373), .O(gate110inter8));
  nand2 gate1144(.a(gate110inter8), .b(gate110inter7), .O(gate110inter9));
  nand2 gate1145(.a(s_85), .b(gate110inter3), .O(gate110inter10));
  nor2  gate1146(.a(gate110inter10), .b(gate110inter9), .O(gate110inter11));
  nor2  gate1147(.a(gate110inter11), .b(gate110inter6), .O(gate110inter12));
  nand2 gate1148(.a(gate110inter12), .b(gate110inter1), .O(G441));

  xor2  gate939(.a(G375), .b(G374), .O(gate111inter0));
  nand2 gate940(.a(gate111inter0), .b(s_56), .O(gate111inter1));
  and2  gate941(.a(G375), .b(G374), .O(gate111inter2));
  inv1  gate942(.a(s_56), .O(gate111inter3));
  inv1  gate943(.a(s_57), .O(gate111inter4));
  nand2 gate944(.a(gate111inter4), .b(gate111inter3), .O(gate111inter5));
  nor2  gate945(.a(gate111inter5), .b(gate111inter2), .O(gate111inter6));
  inv1  gate946(.a(G374), .O(gate111inter7));
  inv1  gate947(.a(G375), .O(gate111inter8));
  nand2 gate948(.a(gate111inter8), .b(gate111inter7), .O(gate111inter9));
  nand2 gate949(.a(s_57), .b(gate111inter3), .O(gate111inter10));
  nor2  gate950(.a(gate111inter10), .b(gate111inter9), .O(gate111inter11));
  nor2  gate951(.a(gate111inter11), .b(gate111inter6), .O(gate111inter12));
  nand2 gate952(.a(gate111inter12), .b(gate111inter1), .O(G444));
nand2 gate112( .a(G376), .b(G377), .O(G447) );
nand2 gate113( .a(G378), .b(G379), .O(G450) );
nand2 gate114( .a(G380), .b(G381), .O(G453) );
nand2 gate115( .a(G382), .b(G383), .O(G456) );
nand2 gate116( .a(G384), .b(G385), .O(G459) );
nand2 gate117( .a(G386), .b(G387), .O(G462) );
nand2 gate118( .a(G388), .b(G389), .O(G465) );

  xor2  gate2059(.a(G391), .b(G390), .O(gate119inter0));
  nand2 gate2060(.a(gate119inter0), .b(s_216), .O(gate119inter1));
  and2  gate2061(.a(G391), .b(G390), .O(gate119inter2));
  inv1  gate2062(.a(s_216), .O(gate119inter3));
  inv1  gate2063(.a(s_217), .O(gate119inter4));
  nand2 gate2064(.a(gate119inter4), .b(gate119inter3), .O(gate119inter5));
  nor2  gate2065(.a(gate119inter5), .b(gate119inter2), .O(gate119inter6));
  inv1  gate2066(.a(G390), .O(gate119inter7));
  inv1  gate2067(.a(G391), .O(gate119inter8));
  nand2 gate2068(.a(gate119inter8), .b(gate119inter7), .O(gate119inter9));
  nand2 gate2069(.a(s_217), .b(gate119inter3), .O(gate119inter10));
  nor2  gate2070(.a(gate119inter10), .b(gate119inter9), .O(gate119inter11));
  nor2  gate2071(.a(gate119inter11), .b(gate119inter6), .O(gate119inter12));
  nand2 gate2072(.a(gate119inter12), .b(gate119inter1), .O(G468));
nand2 gate120( .a(G392), .b(G393), .O(G471) );

  xor2  gate673(.a(G395), .b(G394), .O(gate121inter0));
  nand2 gate674(.a(gate121inter0), .b(s_18), .O(gate121inter1));
  and2  gate675(.a(G395), .b(G394), .O(gate121inter2));
  inv1  gate676(.a(s_18), .O(gate121inter3));
  inv1  gate677(.a(s_19), .O(gate121inter4));
  nand2 gate678(.a(gate121inter4), .b(gate121inter3), .O(gate121inter5));
  nor2  gate679(.a(gate121inter5), .b(gate121inter2), .O(gate121inter6));
  inv1  gate680(.a(G394), .O(gate121inter7));
  inv1  gate681(.a(G395), .O(gate121inter8));
  nand2 gate682(.a(gate121inter8), .b(gate121inter7), .O(gate121inter9));
  nand2 gate683(.a(s_19), .b(gate121inter3), .O(gate121inter10));
  nor2  gate684(.a(gate121inter10), .b(gate121inter9), .O(gate121inter11));
  nor2  gate685(.a(gate121inter11), .b(gate121inter6), .O(gate121inter12));
  nand2 gate686(.a(gate121inter12), .b(gate121inter1), .O(G474));

  xor2  gate1247(.a(G397), .b(G396), .O(gate122inter0));
  nand2 gate1248(.a(gate122inter0), .b(s_100), .O(gate122inter1));
  and2  gate1249(.a(G397), .b(G396), .O(gate122inter2));
  inv1  gate1250(.a(s_100), .O(gate122inter3));
  inv1  gate1251(.a(s_101), .O(gate122inter4));
  nand2 gate1252(.a(gate122inter4), .b(gate122inter3), .O(gate122inter5));
  nor2  gate1253(.a(gate122inter5), .b(gate122inter2), .O(gate122inter6));
  inv1  gate1254(.a(G396), .O(gate122inter7));
  inv1  gate1255(.a(G397), .O(gate122inter8));
  nand2 gate1256(.a(gate122inter8), .b(gate122inter7), .O(gate122inter9));
  nand2 gate1257(.a(s_101), .b(gate122inter3), .O(gate122inter10));
  nor2  gate1258(.a(gate122inter10), .b(gate122inter9), .O(gate122inter11));
  nor2  gate1259(.a(gate122inter11), .b(gate122inter6), .O(gate122inter12));
  nand2 gate1260(.a(gate122inter12), .b(gate122inter1), .O(G477));
nand2 gate123( .a(G398), .b(G399), .O(G480) );
nand2 gate124( .a(G400), .b(G401), .O(G483) );
nand2 gate125( .a(G402), .b(G403), .O(G486) );

  xor2  gate659(.a(G405), .b(G404), .O(gate126inter0));
  nand2 gate660(.a(gate126inter0), .b(s_16), .O(gate126inter1));
  and2  gate661(.a(G405), .b(G404), .O(gate126inter2));
  inv1  gate662(.a(s_16), .O(gate126inter3));
  inv1  gate663(.a(s_17), .O(gate126inter4));
  nand2 gate664(.a(gate126inter4), .b(gate126inter3), .O(gate126inter5));
  nor2  gate665(.a(gate126inter5), .b(gate126inter2), .O(gate126inter6));
  inv1  gate666(.a(G404), .O(gate126inter7));
  inv1  gate667(.a(G405), .O(gate126inter8));
  nand2 gate668(.a(gate126inter8), .b(gate126inter7), .O(gate126inter9));
  nand2 gate669(.a(s_17), .b(gate126inter3), .O(gate126inter10));
  nor2  gate670(.a(gate126inter10), .b(gate126inter9), .O(gate126inter11));
  nor2  gate671(.a(gate126inter11), .b(gate126inter6), .O(gate126inter12));
  nand2 gate672(.a(gate126inter12), .b(gate126inter1), .O(G489));

  xor2  gate2409(.a(G407), .b(G406), .O(gate127inter0));
  nand2 gate2410(.a(gate127inter0), .b(s_266), .O(gate127inter1));
  and2  gate2411(.a(G407), .b(G406), .O(gate127inter2));
  inv1  gate2412(.a(s_266), .O(gate127inter3));
  inv1  gate2413(.a(s_267), .O(gate127inter4));
  nand2 gate2414(.a(gate127inter4), .b(gate127inter3), .O(gate127inter5));
  nor2  gate2415(.a(gate127inter5), .b(gate127inter2), .O(gate127inter6));
  inv1  gate2416(.a(G406), .O(gate127inter7));
  inv1  gate2417(.a(G407), .O(gate127inter8));
  nand2 gate2418(.a(gate127inter8), .b(gate127inter7), .O(gate127inter9));
  nand2 gate2419(.a(s_267), .b(gate127inter3), .O(gate127inter10));
  nor2  gate2420(.a(gate127inter10), .b(gate127inter9), .O(gate127inter11));
  nor2  gate2421(.a(gate127inter11), .b(gate127inter6), .O(gate127inter12));
  nand2 gate2422(.a(gate127inter12), .b(gate127inter1), .O(G492));
nand2 gate128( .a(G408), .b(G409), .O(G495) );
nand2 gate129( .a(G410), .b(G411), .O(G498) );
nand2 gate130( .a(G412), .b(G413), .O(G501) );

  xor2  gate2045(.a(G415), .b(G414), .O(gate131inter0));
  nand2 gate2046(.a(gate131inter0), .b(s_214), .O(gate131inter1));
  and2  gate2047(.a(G415), .b(G414), .O(gate131inter2));
  inv1  gate2048(.a(s_214), .O(gate131inter3));
  inv1  gate2049(.a(s_215), .O(gate131inter4));
  nand2 gate2050(.a(gate131inter4), .b(gate131inter3), .O(gate131inter5));
  nor2  gate2051(.a(gate131inter5), .b(gate131inter2), .O(gate131inter6));
  inv1  gate2052(.a(G414), .O(gate131inter7));
  inv1  gate2053(.a(G415), .O(gate131inter8));
  nand2 gate2054(.a(gate131inter8), .b(gate131inter7), .O(gate131inter9));
  nand2 gate2055(.a(s_215), .b(gate131inter3), .O(gate131inter10));
  nor2  gate2056(.a(gate131inter10), .b(gate131inter9), .O(gate131inter11));
  nor2  gate2057(.a(gate131inter11), .b(gate131inter6), .O(gate131inter12));
  nand2 gate2058(.a(gate131inter12), .b(gate131inter1), .O(G504));
nand2 gate132( .a(G416), .b(G417), .O(G507) );
nand2 gate133( .a(G418), .b(G419), .O(G510) );
nand2 gate134( .a(G420), .b(G421), .O(G513) );
nand2 gate135( .a(G422), .b(G423), .O(G516) );
nand2 gate136( .a(G424), .b(G425), .O(G519) );

  xor2  gate1681(.a(G429), .b(G426), .O(gate137inter0));
  nand2 gate1682(.a(gate137inter0), .b(s_162), .O(gate137inter1));
  and2  gate1683(.a(G429), .b(G426), .O(gate137inter2));
  inv1  gate1684(.a(s_162), .O(gate137inter3));
  inv1  gate1685(.a(s_163), .O(gate137inter4));
  nand2 gate1686(.a(gate137inter4), .b(gate137inter3), .O(gate137inter5));
  nor2  gate1687(.a(gate137inter5), .b(gate137inter2), .O(gate137inter6));
  inv1  gate1688(.a(G426), .O(gate137inter7));
  inv1  gate1689(.a(G429), .O(gate137inter8));
  nand2 gate1690(.a(gate137inter8), .b(gate137inter7), .O(gate137inter9));
  nand2 gate1691(.a(s_163), .b(gate137inter3), .O(gate137inter10));
  nor2  gate1692(.a(gate137inter10), .b(gate137inter9), .O(gate137inter11));
  nor2  gate1693(.a(gate137inter11), .b(gate137inter6), .O(gate137inter12));
  nand2 gate1694(.a(gate137inter12), .b(gate137inter1), .O(G522));

  xor2  gate1051(.a(G435), .b(G432), .O(gate138inter0));
  nand2 gate1052(.a(gate138inter0), .b(s_72), .O(gate138inter1));
  and2  gate1053(.a(G435), .b(G432), .O(gate138inter2));
  inv1  gate1054(.a(s_72), .O(gate138inter3));
  inv1  gate1055(.a(s_73), .O(gate138inter4));
  nand2 gate1056(.a(gate138inter4), .b(gate138inter3), .O(gate138inter5));
  nor2  gate1057(.a(gate138inter5), .b(gate138inter2), .O(gate138inter6));
  inv1  gate1058(.a(G432), .O(gate138inter7));
  inv1  gate1059(.a(G435), .O(gate138inter8));
  nand2 gate1060(.a(gate138inter8), .b(gate138inter7), .O(gate138inter9));
  nand2 gate1061(.a(s_73), .b(gate138inter3), .O(gate138inter10));
  nor2  gate1062(.a(gate138inter10), .b(gate138inter9), .O(gate138inter11));
  nor2  gate1063(.a(gate138inter11), .b(gate138inter6), .O(gate138inter12));
  nand2 gate1064(.a(gate138inter12), .b(gate138inter1), .O(G525));
nand2 gate139( .a(G438), .b(G441), .O(G528) );
nand2 gate140( .a(G444), .b(G447), .O(G531) );

  xor2  gate631(.a(G453), .b(G450), .O(gate141inter0));
  nand2 gate632(.a(gate141inter0), .b(s_12), .O(gate141inter1));
  and2  gate633(.a(G453), .b(G450), .O(gate141inter2));
  inv1  gate634(.a(s_12), .O(gate141inter3));
  inv1  gate635(.a(s_13), .O(gate141inter4));
  nand2 gate636(.a(gate141inter4), .b(gate141inter3), .O(gate141inter5));
  nor2  gate637(.a(gate141inter5), .b(gate141inter2), .O(gate141inter6));
  inv1  gate638(.a(G450), .O(gate141inter7));
  inv1  gate639(.a(G453), .O(gate141inter8));
  nand2 gate640(.a(gate141inter8), .b(gate141inter7), .O(gate141inter9));
  nand2 gate641(.a(s_13), .b(gate141inter3), .O(gate141inter10));
  nor2  gate642(.a(gate141inter10), .b(gate141inter9), .O(gate141inter11));
  nor2  gate643(.a(gate141inter11), .b(gate141inter6), .O(gate141inter12));
  nand2 gate644(.a(gate141inter12), .b(gate141inter1), .O(G534));

  xor2  gate1429(.a(G459), .b(G456), .O(gate142inter0));
  nand2 gate1430(.a(gate142inter0), .b(s_126), .O(gate142inter1));
  and2  gate1431(.a(G459), .b(G456), .O(gate142inter2));
  inv1  gate1432(.a(s_126), .O(gate142inter3));
  inv1  gate1433(.a(s_127), .O(gate142inter4));
  nand2 gate1434(.a(gate142inter4), .b(gate142inter3), .O(gate142inter5));
  nor2  gate1435(.a(gate142inter5), .b(gate142inter2), .O(gate142inter6));
  inv1  gate1436(.a(G456), .O(gate142inter7));
  inv1  gate1437(.a(G459), .O(gate142inter8));
  nand2 gate1438(.a(gate142inter8), .b(gate142inter7), .O(gate142inter9));
  nand2 gate1439(.a(s_127), .b(gate142inter3), .O(gate142inter10));
  nor2  gate1440(.a(gate142inter10), .b(gate142inter9), .O(gate142inter11));
  nor2  gate1441(.a(gate142inter11), .b(gate142inter6), .O(gate142inter12));
  nand2 gate1442(.a(gate142inter12), .b(gate142inter1), .O(G537));

  xor2  gate897(.a(G465), .b(G462), .O(gate143inter0));
  nand2 gate898(.a(gate143inter0), .b(s_50), .O(gate143inter1));
  and2  gate899(.a(G465), .b(G462), .O(gate143inter2));
  inv1  gate900(.a(s_50), .O(gate143inter3));
  inv1  gate901(.a(s_51), .O(gate143inter4));
  nand2 gate902(.a(gate143inter4), .b(gate143inter3), .O(gate143inter5));
  nor2  gate903(.a(gate143inter5), .b(gate143inter2), .O(gate143inter6));
  inv1  gate904(.a(G462), .O(gate143inter7));
  inv1  gate905(.a(G465), .O(gate143inter8));
  nand2 gate906(.a(gate143inter8), .b(gate143inter7), .O(gate143inter9));
  nand2 gate907(.a(s_51), .b(gate143inter3), .O(gate143inter10));
  nor2  gate908(.a(gate143inter10), .b(gate143inter9), .O(gate143inter11));
  nor2  gate909(.a(gate143inter11), .b(gate143inter6), .O(gate143inter12));
  nand2 gate910(.a(gate143inter12), .b(gate143inter1), .O(G540));

  xor2  gate1527(.a(G471), .b(G468), .O(gate144inter0));
  nand2 gate1528(.a(gate144inter0), .b(s_140), .O(gate144inter1));
  and2  gate1529(.a(G471), .b(G468), .O(gate144inter2));
  inv1  gate1530(.a(s_140), .O(gate144inter3));
  inv1  gate1531(.a(s_141), .O(gate144inter4));
  nand2 gate1532(.a(gate144inter4), .b(gate144inter3), .O(gate144inter5));
  nor2  gate1533(.a(gate144inter5), .b(gate144inter2), .O(gate144inter6));
  inv1  gate1534(.a(G468), .O(gate144inter7));
  inv1  gate1535(.a(G471), .O(gate144inter8));
  nand2 gate1536(.a(gate144inter8), .b(gate144inter7), .O(gate144inter9));
  nand2 gate1537(.a(s_141), .b(gate144inter3), .O(gate144inter10));
  nor2  gate1538(.a(gate144inter10), .b(gate144inter9), .O(gate144inter11));
  nor2  gate1539(.a(gate144inter11), .b(gate144inter6), .O(gate144inter12));
  nand2 gate1540(.a(gate144inter12), .b(gate144inter1), .O(G543));
nand2 gate145( .a(G474), .b(G477), .O(G546) );

  xor2  gate2311(.a(G483), .b(G480), .O(gate146inter0));
  nand2 gate2312(.a(gate146inter0), .b(s_252), .O(gate146inter1));
  and2  gate2313(.a(G483), .b(G480), .O(gate146inter2));
  inv1  gate2314(.a(s_252), .O(gate146inter3));
  inv1  gate2315(.a(s_253), .O(gate146inter4));
  nand2 gate2316(.a(gate146inter4), .b(gate146inter3), .O(gate146inter5));
  nor2  gate2317(.a(gate146inter5), .b(gate146inter2), .O(gate146inter6));
  inv1  gate2318(.a(G480), .O(gate146inter7));
  inv1  gate2319(.a(G483), .O(gate146inter8));
  nand2 gate2320(.a(gate146inter8), .b(gate146inter7), .O(gate146inter9));
  nand2 gate2321(.a(s_253), .b(gate146inter3), .O(gate146inter10));
  nor2  gate2322(.a(gate146inter10), .b(gate146inter9), .O(gate146inter11));
  nor2  gate2323(.a(gate146inter11), .b(gate146inter6), .O(gate146inter12));
  nand2 gate2324(.a(gate146inter12), .b(gate146inter1), .O(G549));
nand2 gate147( .a(G486), .b(G489), .O(G552) );
nand2 gate148( .a(G492), .b(G495), .O(G555) );
nand2 gate149( .a(G498), .b(G501), .O(G558) );

  xor2  gate2325(.a(G507), .b(G504), .O(gate150inter0));
  nand2 gate2326(.a(gate150inter0), .b(s_254), .O(gate150inter1));
  and2  gate2327(.a(G507), .b(G504), .O(gate150inter2));
  inv1  gate2328(.a(s_254), .O(gate150inter3));
  inv1  gate2329(.a(s_255), .O(gate150inter4));
  nand2 gate2330(.a(gate150inter4), .b(gate150inter3), .O(gate150inter5));
  nor2  gate2331(.a(gate150inter5), .b(gate150inter2), .O(gate150inter6));
  inv1  gate2332(.a(G504), .O(gate150inter7));
  inv1  gate2333(.a(G507), .O(gate150inter8));
  nand2 gate2334(.a(gate150inter8), .b(gate150inter7), .O(gate150inter9));
  nand2 gate2335(.a(s_255), .b(gate150inter3), .O(gate150inter10));
  nor2  gate2336(.a(gate150inter10), .b(gate150inter9), .O(gate150inter11));
  nor2  gate2337(.a(gate150inter11), .b(gate150inter6), .O(gate150inter12));
  nand2 gate2338(.a(gate150inter12), .b(gate150inter1), .O(G561));
nand2 gate151( .a(G510), .b(G513), .O(G564) );
nand2 gate152( .a(G516), .b(G519), .O(G567) );

  xor2  gate1079(.a(G522), .b(G426), .O(gate153inter0));
  nand2 gate1080(.a(gate153inter0), .b(s_76), .O(gate153inter1));
  and2  gate1081(.a(G522), .b(G426), .O(gate153inter2));
  inv1  gate1082(.a(s_76), .O(gate153inter3));
  inv1  gate1083(.a(s_77), .O(gate153inter4));
  nand2 gate1084(.a(gate153inter4), .b(gate153inter3), .O(gate153inter5));
  nor2  gate1085(.a(gate153inter5), .b(gate153inter2), .O(gate153inter6));
  inv1  gate1086(.a(G426), .O(gate153inter7));
  inv1  gate1087(.a(G522), .O(gate153inter8));
  nand2 gate1088(.a(gate153inter8), .b(gate153inter7), .O(gate153inter9));
  nand2 gate1089(.a(s_77), .b(gate153inter3), .O(gate153inter10));
  nor2  gate1090(.a(gate153inter10), .b(gate153inter9), .O(gate153inter11));
  nor2  gate1091(.a(gate153inter11), .b(gate153inter6), .O(gate153inter12));
  nand2 gate1092(.a(gate153inter12), .b(gate153inter1), .O(G570));

  xor2  gate1737(.a(G522), .b(G429), .O(gate154inter0));
  nand2 gate1738(.a(gate154inter0), .b(s_170), .O(gate154inter1));
  and2  gate1739(.a(G522), .b(G429), .O(gate154inter2));
  inv1  gate1740(.a(s_170), .O(gate154inter3));
  inv1  gate1741(.a(s_171), .O(gate154inter4));
  nand2 gate1742(.a(gate154inter4), .b(gate154inter3), .O(gate154inter5));
  nor2  gate1743(.a(gate154inter5), .b(gate154inter2), .O(gate154inter6));
  inv1  gate1744(.a(G429), .O(gate154inter7));
  inv1  gate1745(.a(G522), .O(gate154inter8));
  nand2 gate1746(.a(gate154inter8), .b(gate154inter7), .O(gate154inter9));
  nand2 gate1747(.a(s_171), .b(gate154inter3), .O(gate154inter10));
  nor2  gate1748(.a(gate154inter10), .b(gate154inter9), .O(gate154inter11));
  nor2  gate1749(.a(gate154inter11), .b(gate154inter6), .O(gate154inter12));
  nand2 gate1750(.a(gate154inter12), .b(gate154inter1), .O(G571));
nand2 gate155( .a(G432), .b(G525), .O(G572) );
nand2 gate156( .a(G435), .b(G525), .O(G573) );
nand2 gate157( .a(G438), .b(G528), .O(G574) );
nand2 gate158( .a(G441), .b(G528), .O(G575) );

  xor2  gate1065(.a(G531), .b(G444), .O(gate159inter0));
  nand2 gate1066(.a(gate159inter0), .b(s_74), .O(gate159inter1));
  and2  gate1067(.a(G531), .b(G444), .O(gate159inter2));
  inv1  gate1068(.a(s_74), .O(gate159inter3));
  inv1  gate1069(.a(s_75), .O(gate159inter4));
  nand2 gate1070(.a(gate159inter4), .b(gate159inter3), .O(gate159inter5));
  nor2  gate1071(.a(gate159inter5), .b(gate159inter2), .O(gate159inter6));
  inv1  gate1072(.a(G444), .O(gate159inter7));
  inv1  gate1073(.a(G531), .O(gate159inter8));
  nand2 gate1074(.a(gate159inter8), .b(gate159inter7), .O(gate159inter9));
  nand2 gate1075(.a(s_75), .b(gate159inter3), .O(gate159inter10));
  nor2  gate1076(.a(gate159inter10), .b(gate159inter9), .O(gate159inter11));
  nor2  gate1077(.a(gate159inter11), .b(gate159inter6), .O(gate159inter12));
  nand2 gate1078(.a(gate159inter12), .b(gate159inter1), .O(G576));
nand2 gate160( .a(G447), .b(G531), .O(G577) );

  xor2  gate1373(.a(G534), .b(G450), .O(gate161inter0));
  nand2 gate1374(.a(gate161inter0), .b(s_118), .O(gate161inter1));
  and2  gate1375(.a(G534), .b(G450), .O(gate161inter2));
  inv1  gate1376(.a(s_118), .O(gate161inter3));
  inv1  gate1377(.a(s_119), .O(gate161inter4));
  nand2 gate1378(.a(gate161inter4), .b(gate161inter3), .O(gate161inter5));
  nor2  gate1379(.a(gate161inter5), .b(gate161inter2), .O(gate161inter6));
  inv1  gate1380(.a(G450), .O(gate161inter7));
  inv1  gate1381(.a(G534), .O(gate161inter8));
  nand2 gate1382(.a(gate161inter8), .b(gate161inter7), .O(gate161inter9));
  nand2 gate1383(.a(s_119), .b(gate161inter3), .O(gate161inter10));
  nor2  gate1384(.a(gate161inter10), .b(gate161inter9), .O(gate161inter11));
  nor2  gate1385(.a(gate161inter11), .b(gate161inter6), .O(gate161inter12));
  nand2 gate1386(.a(gate161inter12), .b(gate161inter1), .O(G578));
nand2 gate162( .a(G453), .b(G534), .O(G579) );
nand2 gate163( .a(G456), .b(G537), .O(G580) );

  xor2  gate1723(.a(G537), .b(G459), .O(gate164inter0));
  nand2 gate1724(.a(gate164inter0), .b(s_168), .O(gate164inter1));
  and2  gate1725(.a(G537), .b(G459), .O(gate164inter2));
  inv1  gate1726(.a(s_168), .O(gate164inter3));
  inv1  gate1727(.a(s_169), .O(gate164inter4));
  nand2 gate1728(.a(gate164inter4), .b(gate164inter3), .O(gate164inter5));
  nor2  gate1729(.a(gate164inter5), .b(gate164inter2), .O(gate164inter6));
  inv1  gate1730(.a(G459), .O(gate164inter7));
  inv1  gate1731(.a(G537), .O(gate164inter8));
  nand2 gate1732(.a(gate164inter8), .b(gate164inter7), .O(gate164inter9));
  nand2 gate1733(.a(s_169), .b(gate164inter3), .O(gate164inter10));
  nor2  gate1734(.a(gate164inter10), .b(gate164inter9), .O(gate164inter11));
  nor2  gate1735(.a(gate164inter11), .b(gate164inter6), .O(gate164inter12));
  nand2 gate1736(.a(gate164inter12), .b(gate164inter1), .O(G581));

  xor2  gate2115(.a(G540), .b(G462), .O(gate165inter0));
  nand2 gate2116(.a(gate165inter0), .b(s_224), .O(gate165inter1));
  and2  gate2117(.a(G540), .b(G462), .O(gate165inter2));
  inv1  gate2118(.a(s_224), .O(gate165inter3));
  inv1  gate2119(.a(s_225), .O(gate165inter4));
  nand2 gate2120(.a(gate165inter4), .b(gate165inter3), .O(gate165inter5));
  nor2  gate2121(.a(gate165inter5), .b(gate165inter2), .O(gate165inter6));
  inv1  gate2122(.a(G462), .O(gate165inter7));
  inv1  gate2123(.a(G540), .O(gate165inter8));
  nand2 gate2124(.a(gate165inter8), .b(gate165inter7), .O(gate165inter9));
  nand2 gate2125(.a(s_225), .b(gate165inter3), .O(gate165inter10));
  nor2  gate2126(.a(gate165inter10), .b(gate165inter9), .O(gate165inter11));
  nor2  gate2127(.a(gate165inter11), .b(gate165inter6), .O(gate165inter12));
  nand2 gate2128(.a(gate165inter12), .b(gate165inter1), .O(G582));
nand2 gate166( .a(G465), .b(G540), .O(G583) );
nand2 gate167( .a(G468), .b(G543), .O(G584) );

  xor2  gate1793(.a(G543), .b(G471), .O(gate168inter0));
  nand2 gate1794(.a(gate168inter0), .b(s_178), .O(gate168inter1));
  and2  gate1795(.a(G543), .b(G471), .O(gate168inter2));
  inv1  gate1796(.a(s_178), .O(gate168inter3));
  inv1  gate1797(.a(s_179), .O(gate168inter4));
  nand2 gate1798(.a(gate168inter4), .b(gate168inter3), .O(gate168inter5));
  nor2  gate1799(.a(gate168inter5), .b(gate168inter2), .O(gate168inter6));
  inv1  gate1800(.a(G471), .O(gate168inter7));
  inv1  gate1801(.a(G543), .O(gate168inter8));
  nand2 gate1802(.a(gate168inter8), .b(gate168inter7), .O(gate168inter9));
  nand2 gate1803(.a(s_179), .b(gate168inter3), .O(gate168inter10));
  nor2  gate1804(.a(gate168inter10), .b(gate168inter9), .O(gate168inter11));
  nor2  gate1805(.a(gate168inter11), .b(gate168inter6), .O(gate168inter12));
  nand2 gate1806(.a(gate168inter12), .b(gate168inter1), .O(G585));
nand2 gate169( .a(G474), .b(G546), .O(G586) );
nand2 gate170( .a(G477), .b(G546), .O(G587) );
nand2 gate171( .a(G480), .b(G549), .O(G588) );
nand2 gate172( .a(G483), .b(G549), .O(G589) );

  xor2  gate1233(.a(G552), .b(G486), .O(gate173inter0));
  nand2 gate1234(.a(gate173inter0), .b(s_98), .O(gate173inter1));
  and2  gate1235(.a(G552), .b(G486), .O(gate173inter2));
  inv1  gate1236(.a(s_98), .O(gate173inter3));
  inv1  gate1237(.a(s_99), .O(gate173inter4));
  nand2 gate1238(.a(gate173inter4), .b(gate173inter3), .O(gate173inter5));
  nor2  gate1239(.a(gate173inter5), .b(gate173inter2), .O(gate173inter6));
  inv1  gate1240(.a(G486), .O(gate173inter7));
  inv1  gate1241(.a(G552), .O(gate173inter8));
  nand2 gate1242(.a(gate173inter8), .b(gate173inter7), .O(gate173inter9));
  nand2 gate1243(.a(s_99), .b(gate173inter3), .O(gate173inter10));
  nor2  gate1244(.a(gate173inter10), .b(gate173inter9), .O(gate173inter11));
  nor2  gate1245(.a(gate173inter11), .b(gate173inter6), .O(gate173inter12));
  nand2 gate1246(.a(gate173inter12), .b(gate173inter1), .O(G590));
nand2 gate174( .a(G489), .b(G552), .O(G591) );

  xor2  gate1611(.a(G555), .b(G492), .O(gate175inter0));
  nand2 gate1612(.a(gate175inter0), .b(s_152), .O(gate175inter1));
  and2  gate1613(.a(G555), .b(G492), .O(gate175inter2));
  inv1  gate1614(.a(s_152), .O(gate175inter3));
  inv1  gate1615(.a(s_153), .O(gate175inter4));
  nand2 gate1616(.a(gate175inter4), .b(gate175inter3), .O(gate175inter5));
  nor2  gate1617(.a(gate175inter5), .b(gate175inter2), .O(gate175inter6));
  inv1  gate1618(.a(G492), .O(gate175inter7));
  inv1  gate1619(.a(G555), .O(gate175inter8));
  nand2 gate1620(.a(gate175inter8), .b(gate175inter7), .O(gate175inter9));
  nand2 gate1621(.a(s_153), .b(gate175inter3), .O(gate175inter10));
  nor2  gate1622(.a(gate175inter10), .b(gate175inter9), .O(gate175inter11));
  nor2  gate1623(.a(gate175inter11), .b(gate175inter6), .O(gate175inter12));
  nand2 gate1624(.a(gate175inter12), .b(gate175inter1), .O(G592));
nand2 gate176( .a(G495), .b(G555), .O(G593) );
nand2 gate177( .a(G498), .b(G558), .O(G594) );
nand2 gate178( .a(G501), .b(G558), .O(G595) );
nand2 gate179( .a(G504), .b(G561), .O(G596) );
nand2 gate180( .a(G507), .b(G561), .O(G597) );
nand2 gate181( .a(G510), .b(G564), .O(G598) );
nand2 gate182( .a(G513), .b(G564), .O(G599) );
nand2 gate183( .a(G516), .b(G567), .O(G600) );
nand2 gate184( .a(G519), .b(G567), .O(G601) );
nand2 gate185( .a(G570), .b(G571), .O(G602) );
nand2 gate186( .a(G572), .b(G573), .O(G607) );

  xor2  gate1583(.a(G575), .b(G574), .O(gate187inter0));
  nand2 gate1584(.a(gate187inter0), .b(s_148), .O(gate187inter1));
  and2  gate1585(.a(G575), .b(G574), .O(gate187inter2));
  inv1  gate1586(.a(s_148), .O(gate187inter3));
  inv1  gate1587(.a(s_149), .O(gate187inter4));
  nand2 gate1588(.a(gate187inter4), .b(gate187inter3), .O(gate187inter5));
  nor2  gate1589(.a(gate187inter5), .b(gate187inter2), .O(gate187inter6));
  inv1  gate1590(.a(G574), .O(gate187inter7));
  inv1  gate1591(.a(G575), .O(gate187inter8));
  nand2 gate1592(.a(gate187inter8), .b(gate187inter7), .O(gate187inter9));
  nand2 gate1593(.a(s_149), .b(gate187inter3), .O(gate187inter10));
  nor2  gate1594(.a(gate187inter10), .b(gate187inter9), .O(gate187inter11));
  nor2  gate1595(.a(gate187inter11), .b(gate187inter6), .O(gate187inter12));
  nand2 gate1596(.a(gate187inter12), .b(gate187inter1), .O(G612));
nand2 gate188( .a(G576), .b(G577), .O(G617) );

  xor2  gate1933(.a(G579), .b(G578), .O(gate189inter0));
  nand2 gate1934(.a(gate189inter0), .b(s_198), .O(gate189inter1));
  and2  gate1935(.a(G579), .b(G578), .O(gate189inter2));
  inv1  gate1936(.a(s_198), .O(gate189inter3));
  inv1  gate1937(.a(s_199), .O(gate189inter4));
  nand2 gate1938(.a(gate189inter4), .b(gate189inter3), .O(gate189inter5));
  nor2  gate1939(.a(gate189inter5), .b(gate189inter2), .O(gate189inter6));
  inv1  gate1940(.a(G578), .O(gate189inter7));
  inv1  gate1941(.a(G579), .O(gate189inter8));
  nand2 gate1942(.a(gate189inter8), .b(gate189inter7), .O(gate189inter9));
  nand2 gate1943(.a(s_199), .b(gate189inter3), .O(gate189inter10));
  nor2  gate1944(.a(gate189inter10), .b(gate189inter9), .O(gate189inter11));
  nor2  gate1945(.a(gate189inter11), .b(gate189inter6), .O(gate189inter12));
  nand2 gate1946(.a(gate189inter12), .b(gate189inter1), .O(G622));

  xor2  gate1499(.a(G581), .b(G580), .O(gate190inter0));
  nand2 gate1500(.a(gate190inter0), .b(s_136), .O(gate190inter1));
  and2  gate1501(.a(G581), .b(G580), .O(gate190inter2));
  inv1  gate1502(.a(s_136), .O(gate190inter3));
  inv1  gate1503(.a(s_137), .O(gate190inter4));
  nand2 gate1504(.a(gate190inter4), .b(gate190inter3), .O(gate190inter5));
  nor2  gate1505(.a(gate190inter5), .b(gate190inter2), .O(gate190inter6));
  inv1  gate1506(.a(G580), .O(gate190inter7));
  inv1  gate1507(.a(G581), .O(gate190inter8));
  nand2 gate1508(.a(gate190inter8), .b(gate190inter7), .O(gate190inter9));
  nand2 gate1509(.a(s_137), .b(gate190inter3), .O(gate190inter10));
  nor2  gate1510(.a(gate190inter10), .b(gate190inter9), .O(gate190inter11));
  nor2  gate1511(.a(gate190inter11), .b(gate190inter6), .O(gate190inter12));
  nand2 gate1512(.a(gate190inter12), .b(gate190inter1), .O(G627));
nand2 gate191( .a(G582), .b(G583), .O(G632) );

  xor2  gate981(.a(G585), .b(G584), .O(gate192inter0));
  nand2 gate982(.a(gate192inter0), .b(s_62), .O(gate192inter1));
  and2  gate983(.a(G585), .b(G584), .O(gate192inter2));
  inv1  gate984(.a(s_62), .O(gate192inter3));
  inv1  gate985(.a(s_63), .O(gate192inter4));
  nand2 gate986(.a(gate192inter4), .b(gate192inter3), .O(gate192inter5));
  nor2  gate987(.a(gate192inter5), .b(gate192inter2), .O(gate192inter6));
  inv1  gate988(.a(G584), .O(gate192inter7));
  inv1  gate989(.a(G585), .O(gate192inter8));
  nand2 gate990(.a(gate192inter8), .b(gate192inter7), .O(gate192inter9));
  nand2 gate991(.a(s_63), .b(gate192inter3), .O(gate192inter10));
  nor2  gate992(.a(gate192inter10), .b(gate192inter9), .O(gate192inter11));
  nor2  gate993(.a(gate192inter11), .b(gate192inter6), .O(gate192inter12));
  nand2 gate994(.a(gate192inter12), .b(gate192inter1), .O(G637));
nand2 gate193( .a(G586), .b(G587), .O(G642) );
nand2 gate194( .a(G588), .b(G589), .O(G645) );
nand2 gate195( .a(G590), .b(G591), .O(G648) );
nand2 gate196( .a(G592), .b(G593), .O(G651) );

  xor2  gate1303(.a(G595), .b(G594), .O(gate197inter0));
  nand2 gate1304(.a(gate197inter0), .b(s_108), .O(gate197inter1));
  and2  gate1305(.a(G595), .b(G594), .O(gate197inter2));
  inv1  gate1306(.a(s_108), .O(gate197inter3));
  inv1  gate1307(.a(s_109), .O(gate197inter4));
  nand2 gate1308(.a(gate197inter4), .b(gate197inter3), .O(gate197inter5));
  nor2  gate1309(.a(gate197inter5), .b(gate197inter2), .O(gate197inter6));
  inv1  gate1310(.a(G594), .O(gate197inter7));
  inv1  gate1311(.a(G595), .O(gate197inter8));
  nand2 gate1312(.a(gate197inter8), .b(gate197inter7), .O(gate197inter9));
  nand2 gate1313(.a(s_109), .b(gate197inter3), .O(gate197inter10));
  nor2  gate1314(.a(gate197inter10), .b(gate197inter9), .O(gate197inter11));
  nor2  gate1315(.a(gate197inter11), .b(gate197inter6), .O(gate197inter12));
  nand2 gate1316(.a(gate197inter12), .b(gate197inter1), .O(G654));
nand2 gate198( .a(G596), .b(G597), .O(G657) );
nand2 gate199( .a(G598), .b(G599), .O(G660) );

  xor2  gate1177(.a(G601), .b(G600), .O(gate200inter0));
  nand2 gate1178(.a(gate200inter0), .b(s_90), .O(gate200inter1));
  and2  gate1179(.a(G601), .b(G600), .O(gate200inter2));
  inv1  gate1180(.a(s_90), .O(gate200inter3));
  inv1  gate1181(.a(s_91), .O(gate200inter4));
  nand2 gate1182(.a(gate200inter4), .b(gate200inter3), .O(gate200inter5));
  nor2  gate1183(.a(gate200inter5), .b(gate200inter2), .O(gate200inter6));
  inv1  gate1184(.a(G600), .O(gate200inter7));
  inv1  gate1185(.a(G601), .O(gate200inter8));
  nand2 gate1186(.a(gate200inter8), .b(gate200inter7), .O(gate200inter9));
  nand2 gate1187(.a(s_91), .b(gate200inter3), .O(gate200inter10));
  nor2  gate1188(.a(gate200inter10), .b(gate200inter9), .O(gate200inter11));
  nor2  gate1189(.a(gate200inter11), .b(gate200inter6), .O(gate200inter12));
  nand2 gate1190(.a(gate200inter12), .b(gate200inter1), .O(G663));

  xor2  gate2087(.a(G607), .b(G602), .O(gate201inter0));
  nand2 gate2088(.a(gate201inter0), .b(s_220), .O(gate201inter1));
  and2  gate2089(.a(G607), .b(G602), .O(gate201inter2));
  inv1  gate2090(.a(s_220), .O(gate201inter3));
  inv1  gate2091(.a(s_221), .O(gate201inter4));
  nand2 gate2092(.a(gate201inter4), .b(gate201inter3), .O(gate201inter5));
  nor2  gate2093(.a(gate201inter5), .b(gate201inter2), .O(gate201inter6));
  inv1  gate2094(.a(G602), .O(gate201inter7));
  inv1  gate2095(.a(G607), .O(gate201inter8));
  nand2 gate2096(.a(gate201inter8), .b(gate201inter7), .O(gate201inter9));
  nand2 gate2097(.a(s_221), .b(gate201inter3), .O(gate201inter10));
  nor2  gate2098(.a(gate201inter10), .b(gate201inter9), .O(gate201inter11));
  nor2  gate2099(.a(gate201inter11), .b(gate201inter6), .O(gate201inter12));
  nand2 gate2100(.a(gate201inter12), .b(gate201inter1), .O(G666));
nand2 gate202( .a(G612), .b(G617), .O(G669) );
nand2 gate203( .a(G602), .b(G612), .O(G672) );

  xor2  gate1107(.a(G617), .b(G607), .O(gate204inter0));
  nand2 gate1108(.a(gate204inter0), .b(s_80), .O(gate204inter1));
  and2  gate1109(.a(G617), .b(G607), .O(gate204inter2));
  inv1  gate1110(.a(s_80), .O(gate204inter3));
  inv1  gate1111(.a(s_81), .O(gate204inter4));
  nand2 gate1112(.a(gate204inter4), .b(gate204inter3), .O(gate204inter5));
  nor2  gate1113(.a(gate204inter5), .b(gate204inter2), .O(gate204inter6));
  inv1  gate1114(.a(G607), .O(gate204inter7));
  inv1  gate1115(.a(G617), .O(gate204inter8));
  nand2 gate1116(.a(gate204inter8), .b(gate204inter7), .O(gate204inter9));
  nand2 gate1117(.a(s_81), .b(gate204inter3), .O(gate204inter10));
  nor2  gate1118(.a(gate204inter10), .b(gate204inter9), .O(gate204inter11));
  nor2  gate1119(.a(gate204inter11), .b(gate204inter6), .O(gate204inter12));
  nand2 gate1120(.a(gate204inter12), .b(gate204inter1), .O(G675));

  xor2  gate1835(.a(G627), .b(G622), .O(gate205inter0));
  nand2 gate1836(.a(gate205inter0), .b(s_184), .O(gate205inter1));
  and2  gate1837(.a(G627), .b(G622), .O(gate205inter2));
  inv1  gate1838(.a(s_184), .O(gate205inter3));
  inv1  gate1839(.a(s_185), .O(gate205inter4));
  nand2 gate1840(.a(gate205inter4), .b(gate205inter3), .O(gate205inter5));
  nor2  gate1841(.a(gate205inter5), .b(gate205inter2), .O(gate205inter6));
  inv1  gate1842(.a(G622), .O(gate205inter7));
  inv1  gate1843(.a(G627), .O(gate205inter8));
  nand2 gate1844(.a(gate205inter8), .b(gate205inter7), .O(gate205inter9));
  nand2 gate1845(.a(s_185), .b(gate205inter3), .O(gate205inter10));
  nor2  gate1846(.a(gate205inter10), .b(gate205inter9), .O(gate205inter11));
  nor2  gate1847(.a(gate205inter11), .b(gate205inter6), .O(gate205inter12));
  nand2 gate1848(.a(gate205inter12), .b(gate205inter1), .O(G678));
nand2 gate206( .a(G632), .b(G637), .O(G681) );
nand2 gate207( .a(G622), .b(G632), .O(G684) );
nand2 gate208( .a(G627), .b(G637), .O(G687) );

  xor2  gate589(.a(G666), .b(G602), .O(gate209inter0));
  nand2 gate590(.a(gate209inter0), .b(s_6), .O(gate209inter1));
  and2  gate591(.a(G666), .b(G602), .O(gate209inter2));
  inv1  gate592(.a(s_6), .O(gate209inter3));
  inv1  gate593(.a(s_7), .O(gate209inter4));
  nand2 gate594(.a(gate209inter4), .b(gate209inter3), .O(gate209inter5));
  nor2  gate595(.a(gate209inter5), .b(gate209inter2), .O(gate209inter6));
  inv1  gate596(.a(G602), .O(gate209inter7));
  inv1  gate597(.a(G666), .O(gate209inter8));
  nand2 gate598(.a(gate209inter8), .b(gate209inter7), .O(gate209inter9));
  nand2 gate599(.a(s_7), .b(gate209inter3), .O(gate209inter10));
  nor2  gate600(.a(gate209inter10), .b(gate209inter9), .O(gate209inter11));
  nor2  gate601(.a(gate209inter11), .b(gate209inter6), .O(gate209inter12));
  nand2 gate602(.a(gate209inter12), .b(gate209inter1), .O(G690));

  xor2  gate1331(.a(G666), .b(G607), .O(gate210inter0));
  nand2 gate1332(.a(gate210inter0), .b(s_112), .O(gate210inter1));
  and2  gate1333(.a(G666), .b(G607), .O(gate210inter2));
  inv1  gate1334(.a(s_112), .O(gate210inter3));
  inv1  gate1335(.a(s_113), .O(gate210inter4));
  nand2 gate1336(.a(gate210inter4), .b(gate210inter3), .O(gate210inter5));
  nor2  gate1337(.a(gate210inter5), .b(gate210inter2), .O(gate210inter6));
  inv1  gate1338(.a(G607), .O(gate210inter7));
  inv1  gate1339(.a(G666), .O(gate210inter8));
  nand2 gate1340(.a(gate210inter8), .b(gate210inter7), .O(gate210inter9));
  nand2 gate1341(.a(s_113), .b(gate210inter3), .O(gate210inter10));
  nor2  gate1342(.a(gate210inter10), .b(gate210inter9), .O(gate210inter11));
  nor2  gate1343(.a(gate210inter11), .b(gate210inter6), .O(gate210inter12));
  nand2 gate1344(.a(gate210inter12), .b(gate210inter1), .O(G691));

  xor2  gate995(.a(G669), .b(G612), .O(gate211inter0));
  nand2 gate996(.a(gate211inter0), .b(s_64), .O(gate211inter1));
  and2  gate997(.a(G669), .b(G612), .O(gate211inter2));
  inv1  gate998(.a(s_64), .O(gate211inter3));
  inv1  gate999(.a(s_65), .O(gate211inter4));
  nand2 gate1000(.a(gate211inter4), .b(gate211inter3), .O(gate211inter5));
  nor2  gate1001(.a(gate211inter5), .b(gate211inter2), .O(gate211inter6));
  inv1  gate1002(.a(G612), .O(gate211inter7));
  inv1  gate1003(.a(G669), .O(gate211inter8));
  nand2 gate1004(.a(gate211inter8), .b(gate211inter7), .O(gate211inter9));
  nand2 gate1005(.a(s_65), .b(gate211inter3), .O(gate211inter10));
  nor2  gate1006(.a(gate211inter10), .b(gate211inter9), .O(gate211inter11));
  nor2  gate1007(.a(gate211inter11), .b(gate211inter6), .O(gate211inter12));
  nand2 gate1008(.a(gate211inter12), .b(gate211inter1), .O(G692));

  xor2  gate1947(.a(G669), .b(G617), .O(gate212inter0));
  nand2 gate1948(.a(gate212inter0), .b(s_200), .O(gate212inter1));
  and2  gate1949(.a(G669), .b(G617), .O(gate212inter2));
  inv1  gate1950(.a(s_200), .O(gate212inter3));
  inv1  gate1951(.a(s_201), .O(gate212inter4));
  nand2 gate1952(.a(gate212inter4), .b(gate212inter3), .O(gate212inter5));
  nor2  gate1953(.a(gate212inter5), .b(gate212inter2), .O(gate212inter6));
  inv1  gate1954(.a(G617), .O(gate212inter7));
  inv1  gate1955(.a(G669), .O(gate212inter8));
  nand2 gate1956(.a(gate212inter8), .b(gate212inter7), .O(gate212inter9));
  nand2 gate1957(.a(s_201), .b(gate212inter3), .O(gate212inter10));
  nor2  gate1958(.a(gate212inter10), .b(gate212inter9), .O(gate212inter11));
  nor2  gate1959(.a(gate212inter11), .b(gate212inter6), .O(gate212inter12));
  nand2 gate1960(.a(gate212inter12), .b(gate212inter1), .O(G693));
nand2 gate213( .a(G602), .b(G672), .O(G694) );
nand2 gate214( .a(G612), .b(G672), .O(G695) );
nand2 gate215( .a(G607), .b(G675), .O(G696) );

  xor2  gate743(.a(G675), .b(G617), .O(gate216inter0));
  nand2 gate744(.a(gate216inter0), .b(s_28), .O(gate216inter1));
  and2  gate745(.a(G675), .b(G617), .O(gate216inter2));
  inv1  gate746(.a(s_28), .O(gate216inter3));
  inv1  gate747(.a(s_29), .O(gate216inter4));
  nand2 gate748(.a(gate216inter4), .b(gate216inter3), .O(gate216inter5));
  nor2  gate749(.a(gate216inter5), .b(gate216inter2), .O(gate216inter6));
  inv1  gate750(.a(G617), .O(gate216inter7));
  inv1  gate751(.a(G675), .O(gate216inter8));
  nand2 gate752(.a(gate216inter8), .b(gate216inter7), .O(gate216inter9));
  nand2 gate753(.a(s_29), .b(gate216inter3), .O(gate216inter10));
  nor2  gate754(.a(gate216inter10), .b(gate216inter9), .O(gate216inter11));
  nor2  gate755(.a(gate216inter11), .b(gate216inter6), .O(gate216inter12));
  nand2 gate756(.a(gate216inter12), .b(gate216inter1), .O(G697));

  xor2  gate575(.a(G678), .b(G622), .O(gate217inter0));
  nand2 gate576(.a(gate217inter0), .b(s_4), .O(gate217inter1));
  and2  gate577(.a(G678), .b(G622), .O(gate217inter2));
  inv1  gate578(.a(s_4), .O(gate217inter3));
  inv1  gate579(.a(s_5), .O(gate217inter4));
  nand2 gate580(.a(gate217inter4), .b(gate217inter3), .O(gate217inter5));
  nor2  gate581(.a(gate217inter5), .b(gate217inter2), .O(gate217inter6));
  inv1  gate582(.a(G622), .O(gate217inter7));
  inv1  gate583(.a(G678), .O(gate217inter8));
  nand2 gate584(.a(gate217inter8), .b(gate217inter7), .O(gate217inter9));
  nand2 gate585(.a(s_5), .b(gate217inter3), .O(gate217inter10));
  nor2  gate586(.a(gate217inter10), .b(gate217inter9), .O(gate217inter11));
  nor2  gate587(.a(gate217inter11), .b(gate217inter6), .O(gate217inter12));
  nand2 gate588(.a(gate217inter12), .b(gate217inter1), .O(G698));

  xor2  gate2423(.a(G678), .b(G627), .O(gate218inter0));
  nand2 gate2424(.a(gate218inter0), .b(s_268), .O(gate218inter1));
  and2  gate2425(.a(G678), .b(G627), .O(gate218inter2));
  inv1  gate2426(.a(s_268), .O(gate218inter3));
  inv1  gate2427(.a(s_269), .O(gate218inter4));
  nand2 gate2428(.a(gate218inter4), .b(gate218inter3), .O(gate218inter5));
  nor2  gate2429(.a(gate218inter5), .b(gate218inter2), .O(gate218inter6));
  inv1  gate2430(.a(G627), .O(gate218inter7));
  inv1  gate2431(.a(G678), .O(gate218inter8));
  nand2 gate2432(.a(gate218inter8), .b(gate218inter7), .O(gate218inter9));
  nand2 gate2433(.a(s_269), .b(gate218inter3), .O(gate218inter10));
  nor2  gate2434(.a(gate218inter10), .b(gate218inter9), .O(gate218inter11));
  nor2  gate2435(.a(gate218inter11), .b(gate218inter6), .O(gate218inter12));
  nand2 gate2436(.a(gate218inter12), .b(gate218inter1), .O(G699));

  xor2  gate1849(.a(G681), .b(G632), .O(gate219inter0));
  nand2 gate1850(.a(gate219inter0), .b(s_186), .O(gate219inter1));
  and2  gate1851(.a(G681), .b(G632), .O(gate219inter2));
  inv1  gate1852(.a(s_186), .O(gate219inter3));
  inv1  gate1853(.a(s_187), .O(gate219inter4));
  nand2 gate1854(.a(gate219inter4), .b(gate219inter3), .O(gate219inter5));
  nor2  gate1855(.a(gate219inter5), .b(gate219inter2), .O(gate219inter6));
  inv1  gate1856(.a(G632), .O(gate219inter7));
  inv1  gate1857(.a(G681), .O(gate219inter8));
  nand2 gate1858(.a(gate219inter8), .b(gate219inter7), .O(gate219inter9));
  nand2 gate1859(.a(s_187), .b(gate219inter3), .O(gate219inter10));
  nor2  gate1860(.a(gate219inter10), .b(gate219inter9), .O(gate219inter11));
  nor2  gate1861(.a(gate219inter11), .b(gate219inter6), .O(gate219inter12));
  nand2 gate1862(.a(gate219inter12), .b(gate219inter1), .O(G700));
nand2 gate220( .a(G637), .b(G681), .O(G701) );
nand2 gate221( .a(G622), .b(G684), .O(G702) );

  xor2  gate967(.a(G684), .b(G632), .O(gate222inter0));
  nand2 gate968(.a(gate222inter0), .b(s_60), .O(gate222inter1));
  and2  gate969(.a(G684), .b(G632), .O(gate222inter2));
  inv1  gate970(.a(s_60), .O(gate222inter3));
  inv1  gate971(.a(s_61), .O(gate222inter4));
  nand2 gate972(.a(gate222inter4), .b(gate222inter3), .O(gate222inter5));
  nor2  gate973(.a(gate222inter5), .b(gate222inter2), .O(gate222inter6));
  inv1  gate974(.a(G632), .O(gate222inter7));
  inv1  gate975(.a(G684), .O(gate222inter8));
  nand2 gate976(.a(gate222inter8), .b(gate222inter7), .O(gate222inter9));
  nand2 gate977(.a(s_61), .b(gate222inter3), .O(gate222inter10));
  nor2  gate978(.a(gate222inter10), .b(gate222inter9), .O(gate222inter11));
  nor2  gate979(.a(gate222inter11), .b(gate222inter6), .O(gate222inter12));
  nand2 gate980(.a(gate222inter12), .b(gate222inter1), .O(G703));
nand2 gate223( .a(G627), .b(G687), .O(G704) );
nand2 gate224( .a(G637), .b(G687), .O(G705) );
nand2 gate225( .a(G690), .b(G691), .O(G706) );
nand2 gate226( .a(G692), .b(G693), .O(G709) );
nand2 gate227( .a(G694), .b(G695), .O(G712) );
nand2 gate228( .a(G696), .b(G697), .O(G715) );
nand2 gate229( .a(G698), .b(G699), .O(G718) );
nand2 gate230( .a(G700), .b(G701), .O(G721) );

  xor2  gate953(.a(G703), .b(G702), .O(gate231inter0));
  nand2 gate954(.a(gate231inter0), .b(s_58), .O(gate231inter1));
  and2  gate955(.a(G703), .b(G702), .O(gate231inter2));
  inv1  gate956(.a(s_58), .O(gate231inter3));
  inv1  gate957(.a(s_59), .O(gate231inter4));
  nand2 gate958(.a(gate231inter4), .b(gate231inter3), .O(gate231inter5));
  nor2  gate959(.a(gate231inter5), .b(gate231inter2), .O(gate231inter6));
  inv1  gate960(.a(G702), .O(gate231inter7));
  inv1  gate961(.a(G703), .O(gate231inter8));
  nand2 gate962(.a(gate231inter8), .b(gate231inter7), .O(gate231inter9));
  nand2 gate963(.a(s_59), .b(gate231inter3), .O(gate231inter10));
  nor2  gate964(.a(gate231inter10), .b(gate231inter9), .O(gate231inter11));
  nor2  gate965(.a(gate231inter11), .b(gate231inter6), .O(gate231inter12));
  nand2 gate966(.a(gate231inter12), .b(gate231inter1), .O(G724));
nand2 gate232( .a(G704), .b(G705), .O(G727) );

  xor2  gate1653(.a(G718), .b(G242), .O(gate233inter0));
  nand2 gate1654(.a(gate233inter0), .b(s_158), .O(gate233inter1));
  and2  gate1655(.a(G718), .b(G242), .O(gate233inter2));
  inv1  gate1656(.a(s_158), .O(gate233inter3));
  inv1  gate1657(.a(s_159), .O(gate233inter4));
  nand2 gate1658(.a(gate233inter4), .b(gate233inter3), .O(gate233inter5));
  nor2  gate1659(.a(gate233inter5), .b(gate233inter2), .O(gate233inter6));
  inv1  gate1660(.a(G242), .O(gate233inter7));
  inv1  gate1661(.a(G718), .O(gate233inter8));
  nand2 gate1662(.a(gate233inter8), .b(gate233inter7), .O(gate233inter9));
  nand2 gate1663(.a(s_159), .b(gate233inter3), .O(gate233inter10));
  nor2  gate1664(.a(gate233inter10), .b(gate233inter9), .O(gate233inter11));
  nor2  gate1665(.a(gate233inter11), .b(gate233inter6), .O(gate233inter12));
  nand2 gate1666(.a(gate233inter12), .b(gate233inter1), .O(G730));

  xor2  gate1905(.a(G721), .b(G245), .O(gate234inter0));
  nand2 gate1906(.a(gate234inter0), .b(s_194), .O(gate234inter1));
  and2  gate1907(.a(G721), .b(G245), .O(gate234inter2));
  inv1  gate1908(.a(s_194), .O(gate234inter3));
  inv1  gate1909(.a(s_195), .O(gate234inter4));
  nand2 gate1910(.a(gate234inter4), .b(gate234inter3), .O(gate234inter5));
  nor2  gate1911(.a(gate234inter5), .b(gate234inter2), .O(gate234inter6));
  inv1  gate1912(.a(G245), .O(gate234inter7));
  inv1  gate1913(.a(G721), .O(gate234inter8));
  nand2 gate1914(.a(gate234inter8), .b(gate234inter7), .O(gate234inter9));
  nand2 gate1915(.a(s_195), .b(gate234inter3), .O(gate234inter10));
  nor2  gate1916(.a(gate234inter10), .b(gate234inter9), .O(gate234inter11));
  nor2  gate1917(.a(gate234inter11), .b(gate234inter6), .O(gate234inter12));
  nand2 gate1918(.a(gate234inter12), .b(gate234inter1), .O(G733));
nand2 gate235( .a(G248), .b(G724), .O(G736) );
nand2 gate236( .a(G251), .b(G727), .O(G739) );

  xor2  gate1401(.a(G706), .b(G254), .O(gate237inter0));
  nand2 gate1402(.a(gate237inter0), .b(s_122), .O(gate237inter1));
  and2  gate1403(.a(G706), .b(G254), .O(gate237inter2));
  inv1  gate1404(.a(s_122), .O(gate237inter3));
  inv1  gate1405(.a(s_123), .O(gate237inter4));
  nand2 gate1406(.a(gate237inter4), .b(gate237inter3), .O(gate237inter5));
  nor2  gate1407(.a(gate237inter5), .b(gate237inter2), .O(gate237inter6));
  inv1  gate1408(.a(G254), .O(gate237inter7));
  inv1  gate1409(.a(G706), .O(gate237inter8));
  nand2 gate1410(.a(gate237inter8), .b(gate237inter7), .O(gate237inter9));
  nand2 gate1411(.a(s_123), .b(gate237inter3), .O(gate237inter10));
  nor2  gate1412(.a(gate237inter10), .b(gate237inter9), .O(gate237inter11));
  nor2  gate1413(.a(gate237inter11), .b(gate237inter6), .O(gate237inter12));
  nand2 gate1414(.a(gate237inter12), .b(gate237inter1), .O(G742));

  xor2  gate2157(.a(G709), .b(G257), .O(gate238inter0));
  nand2 gate2158(.a(gate238inter0), .b(s_230), .O(gate238inter1));
  and2  gate2159(.a(G709), .b(G257), .O(gate238inter2));
  inv1  gate2160(.a(s_230), .O(gate238inter3));
  inv1  gate2161(.a(s_231), .O(gate238inter4));
  nand2 gate2162(.a(gate238inter4), .b(gate238inter3), .O(gate238inter5));
  nor2  gate2163(.a(gate238inter5), .b(gate238inter2), .O(gate238inter6));
  inv1  gate2164(.a(G257), .O(gate238inter7));
  inv1  gate2165(.a(G709), .O(gate238inter8));
  nand2 gate2166(.a(gate238inter8), .b(gate238inter7), .O(gate238inter9));
  nand2 gate2167(.a(s_231), .b(gate238inter3), .O(gate238inter10));
  nor2  gate2168(.a(gate238inter10), .b(gate238inter9), .O(gate238inter11));
  nor2  gate2169(.a(gate238inter11), .b(gate238inter6), .O(gate238inter12));
  nand2 gate2170(.a(gate238inter12), .b(gate238inter1), .O(G745));
nand2 gate239( .a(G260), .b(G712), .O(G748) );
nand2 gate240( .a(G263), .b(G715), .O(G751) );
nand2 gate241( .a(G242), .b(G730), .O(G754) );
nand2 gate242( .a(G718), .b(G730), .O(G755) );
nand2 gate243( .a(G245), .b(G733), .O(G756) );
nand2 gate244( .a(G721), .b(G733), .O(G757) );

  xor2  gate645(.a(G736), .b(G248), .O(gate245inter0));
  nand2 gate646(.a(gate245inter0), .b(s_14), .O(gate245inter1));
  and2  gate647(.a(G736), .b(G248), .O(gate245inter2));
  inv1  gate648(.a(s_14), .O(gate245inter3));
  inv1  gate649(.a(s_15), .O(gate245inter4));
  nand2 gate650(.a(gate245inter4), .b(gate245inter3), .O(gate245inter5));
  nor2  gate651(.a(gate245inter5), .b(gate245inter2), .O(gate245inter6));
  inv1  gate652(.a(G248), .O(gate245inter7));
  inv1  gate653(.a(G736), .O(gate245inter8));
  nand2 gate654(.a(gate245inter8), .b(gate245inter7), .O(gate245inter9));
  nand2 gate655(.a(s_15), .b(gate245inter3), .O(gate245inter10));
  nor2  gate656(.a(gate245inter10), .b(gate245inter9), .O(gate245inter11));
  nor2  gate657(.a(gate245inter11), .b(gate245inter6), .O(gate245inter12));
  nand2 gate658(.a(gate245inter12), .b(gate245inter1), .O(G758));

  xor2  gate2017(.a(G736), .b(G724), .O(gate246inter0));
  nand2 gate2018(.a(gate246inter0), .b(s_210), .O(gate246inter1));
  and2  gate2019(.a(G736), .b(G724), .O(gate246inter2));
  inv1  gate2020(.a(s_210), .O(gate246inter3));
  inv1  gate2021(.a(s_211), .O(gate246inter4));
  nand2 gate2022(.a(gate246inter4), .b(gate246inter3), .O(gate246inter5));
  nor2  gate2023(.a(gate246inter5), .b(gate246inter2), .O(gate246inter6));
  inv1  gate2024(.a(G724), .O(gate246inter7));
  inv1  gate2025(.a(G736), .O(gate246inter8));
  nand2 gate2026(.a(gate246inter8), .b(gate246inter7), .O(gate246inter9));
  nand2 gate2027(.a(s_211), .b(gate246inter3), .O(gate246inter10));
  nor2  gate2028(.a(gate246inter10), .b(gate246inter9), .O(gate246inter11));
  nor2  gate2029(.a(gate246inter11), .b(gate246inter6), .O(gate246inter12));
  nand2 gate2030(.a(gate246inter12), .b(gate246inter1), .O(G759));
nand2 gate247( .a(G251), .b(G739), .O(G760) );

  xor2  gate2297(.a(G739), .b(G727), .O(gate248inter0));
  nand2 gate2298(.a(gate248inter0), .b(s_250), .O(gate248inter1));
  and2  gate2299(.a(G739), .b(G727), .O(gate248inter2));
  inv1  gate2300(.a(s_250), .O(gate248inter3));
  inv1  gate2301(.a(s_251), .O(gate248inter4));
  nand2 gate2302(.a(gate248inter4), .b(gate248inter3), .O(gate248inter5));
  nor2  gate2303(.a(gate248inter5), .b(gate248inter2), .O(gate248inter6));
  inv1  gate2304(.a(G727), .O(gate248inter7));
  inv1  gate2305(.a(G739), .O(gate248inter8));
  nand2 gate2306(.a(gate248inter8), .b(gate248inter7), .O(gate248inter9));
  nand2 gate2307(.a(s_251), .b(gate248inter3), .O(gate248inter10));
  nor2  gate2308(.a(gate248inter10), .b(gate248inter9), .O(gate248inter11));
  nor2  gate2309(.a(gate248inter11), .b(gate248inter6), .O(gate248inter12));
  nand2 gate2310(.a(gate248inter12), .b(gate248inter1), .O(G761));
nand2 gate249( .a(G254), .b(G742), .O(G762) );
nand2 gate250( .a(G706), .b(G742), .O(G763) );
nand2 gate251( .a(G257), .b(G745), .O(G764) );

  xor2  gate1597(.a(G745), .b(G709), .O(gate252inter0));
  nand2 gate1598(.a(gate252inter0), .b(s_150), .O(gate252inter1));
  and2  gate1599(.a(G745), .b(G709), .O(gate252inter2));
  inv1  gate1600(.a(s_150), .O(gate252inter3));
  inv1  gate1601(.a(s_151), .O(gate252inter4));
  nand2 gate1602(.a(gate252inter4), .b(gate252inter3), .O(gate252inter5));
  nor2  gate1603(.a(gate252inter5), .b(gate252inter2), .O(gate252inter6));
  inv1  gate1604(.a(G709), .O(gate252inter7));
  inv1  gate1605(.a(G745), .O(gate252inter8));
  nand2 gate1606(.a(gate252inter8), .b(gate252inter7), .O(gate252inter9));
  nand2 gate1607(.a(s_151), .b(gate252inter3), .O(gate252inter10));
  nor2  gate1608(.a(gate252inter10), .b(gate252inter9), .O(gate252inter11));
  nor2  gate1609(.a(gate252inter11), .b(gate252inter6), .O(gate252inter12));
  nand2 gate1610(.a(gate252inter12), .b(gate252inter1), .O(G765));

  xor2  gate2101(.a(G748), .b(G260), .O(gate253inter0));
  nand2 gate2102(.a(gate253inter0), .b(s_222), .O(gate253inter1));
  and2  gate2103(.a(G748), .b(G260), .O(gate253inter2));
  inv1  gate2104(.a(s_222), .O(gate253inter3));
  inv1  gate2105(.a(s_223), .O(gate253inter4));
  nand2 gate2106(.a(gate253inter4), .b(gate253inter3), .O(gate253inter5));
  nor2  gate2107(.a(gate253inter5), .b(gate253inter2), .O(gate253inter6));
  inv1  gate2108(.a(G260), .O(gate253inter7));
  inv1  gate2109(.a(G748), .O(gate253inter8));
  nand2 gate2110(.a(gate253inter8), .b(gate253inter7), .O(gate253inter9));
  nand2 gate2111(.a(s_223), .b(gate253inter3), .O(gate253inter10));
  nor2  gate2112(.a(gate253inter10), .b(gate253inter9), .O(gate253inter11));
  nor2  gate2113(.a(gate253inter11), .b(gate253inter6), .O(gate253inter12));
  nand2 gate2114(.a(gate253inter12), .b(gate253inter1), .O(G766));

  xor2  gate1163(.a(G748), .b(G712), .O(gate254inter0));
  nand2 gate1164(.a(gate254inter0), .b(s_88), .O(gate254inter1));
  and2  gate1165(.a(G748), .b(G712), .O(gate254inter2));
  inv1  gate1166(.a(s_88), .O(gate254inter3));
  inv1  gate1167(.a(s_89), .O(gate254inter4));
  nand2 gate1168(.a(gate254inter4), .b(gate254inter3), .O(gate254inter5));
  nor2  gate1169(.a(gate254inter5), .b(gate254inter2), .O(gate254inter6));
  inv1  gate1170(.a(G712), .O(gate254inter7));
  inv1  gate1171(.a(G748), .O(gate254inter8));
  nand2 gate1172(.a(gate254inter8), .b(gate254inter7), .O(gate254inter9));
  nand2 gate1173(.a(s_89), .b(gate254inter3), .O(gate254inter10));
  nor2  gate1174(.a(gate254inter10), .b(gate254inter9), .O(gate254inter11));
  nor2  gate1175(.a(gate254inter11), .b(gate254inter6), .O(gate254inter12));
  nand2 gate1176(.a(gate254inter12), .b(gate254inter1), .O(G767));
nand2 gate255( .a(G263), .b(G751), .O(G768) );

  xor2  gate1975(.a(G751), .b(G715), .O(gate256inter0));
  nand2 gate1976(.a(gate256inter0), .b(s_204), .O(gate256inter1));
  and2  gate1977(.a(G751), .b(G715), .O(gate256inter2));
  inv1  gate1978(.a(s_204), .O(gate256inter3));
  inv1  gate1979(.a(s_205), .O(gate256inter4));
  nand2 gate1980(.a(gate256inter4), .b(gate256inter3), .O(gate256inter5));
  nor2  gate1981(.a(gate256inter5), .b(gate256inter2), .O(gate256inter6));
  inv1  gate1982(.a(G715), .O(gate256inter7));
  inv1  gate1983(.a(G751), .O(gate256inter8));
  nand2 gate1984(.a(gate256inter8), .b(gate256inter7), .O(gate256inter9));
  nand2 gate1985(.a(s_205), .b(gate256inter3), .O(gate256inter10));
  nor2  gate1986(.a(gate256inter10), .b(gate256inter9), .O(gate256inter11));
  nor2  gate1987(.a(gate256inter11), .b(gate256inter6), .O(gate256inter12));
  nand2 gate1988(.a(gate256inter12), .b(gate256inter1), .O(G769));
nand2 gate257( .a(G754), .b(G755), .O(G770) );

  xor2  gate2255(.a(G757), .b(G756), .O(gate258inter0));
  nand2 gate2256(.a(gate258inter0), .b(s_244), .O(gate258inter1));
  and2  gate2257(.a(G757), .b(G756), .O(gate258inter2));
  inv1  gate2258(.a(s_244), .O(gate258inter3));
  inv1  gate2259(.a(s_245), .O(gate258inter4));
  nand2 gate2260(.a(gate258inter4), .b(gate258inter3), .O(gate258inter5));
  nor2  gate2261(.a(gate258inter5), .b(gate258inter2), .O(gate258inter6));
  inv1  gate2262(.a(G756), .O(gate258inter7));
  inv1  gate2263(.a(G757), .O(gate258inter8));
  nand2 gate2264(.a(gate258inter8), .b(gate258inter7), .O(gate258inter9));
  nand2 gate2265(.a(s_245), .b(gate258inter3), .O(gate258inter10));
  nor2  gate2266(.a(gate258inter10), .b(gate258inter9), .O(gate258inter11));
  nor2  gate2267(.a(gate258inter11), .b(gate258inter6), .O(gate258inter12));
  nand2 gate2268(.a(gate258inter12), .b(gate258inter1), .O(G773));
nand2 gate259( .a(G758), .b(G759), .O(G776) );

  xor2  gate603(.a(G761), .b(G760), .O(gate260inter0));
  nand2 gate604(.a(gate260inter0), .b(s_8), .O(gate260inter1));
  and2  gate605(.a(G761), .b(G760), .O(gate260inter2));
  inv1  gate606(.a(s_8), .O(gate260inter3));
  inv1  gate607(.a(s_9), .O(gate260inter4));
  nand2 gate608(.a(gate260inter4), .b(gate260inter3), .O(gate260inter5));
  nor2  gate609(.a(gate260inter5), .b(gate260inter2), .O(gate260inter6));
  inv1  gate610(.a(G760), .O(gate260inter7));
  inv1  gate611(.a(G761), .O(gate260inter8));
  nand2 gate612(.a(gate260inter8), .b(gate260inter7), .O(gate260inter9));
  nand2 gate613(.a(s_9), .b(gate260inter3), .O(gate260inter10));
  nor2  gate614(.a(gate260inter10), .b(gate260inter9), .O(gate260inter11));
  nor2  gate615(.a(gate260inter11), .b(gate260inter6), .O(gate260inter12));
  nand2 gate616(.a(gate260inter12), .b(gate260inter1), .O(G779));
nand2 gate261( .a(G762), .b(G763), .O(G782) );

  xor2  gate2031(.a(G765), .b(G764), .O(gate262inter0));
  nand2 gate2032(.a(gate262inter0), .b(s_212), .O(gate262inter1));
  and2  gate2033(.a(G765), .b(G764), .O(gate262inter2));
  inv1  gate2034(.a(s_212), .O(gate262inter3));
  inv1  gate2035(.a(s_213), .O(gate262inter4));
  nand2 gate2036(.a(gate262inter4), .b(gate262inter3), .O(gate262inter5));
  nor2  gate2037(.a(gate262inter5), .b(gate262inter2), .O(gate262inter6));
  inv1  gate2038(.a(G764), .O(gate262inter7));
  inv1  gate2039(.a(G765), .O(gate262inter8));
  nand2 gate2040(.a(gate262inter8), .b(gate262inter7), .O(gate262inter9));
  nand2 gate2041(.a(s_213), .b(gate262inter3), .O(gate262inter10));
  nor2  gate2042(.a(gate262inter10), .b(gate262inter9), .O(gate262inter11));
  nor2  gate2043(.a(gate262inter11), .b(gate262inter6), .O(gate262inter12));
  nand2 gate2044(.a(gate262inter12), .b(gate262inter1), .O(G785));
nand2 gate263( .a(G766), .b(G767), .O(G788) );
nand2 gate264( .a(G768), .b(G769), .O(G791) );
nand2 gate265( .a(G642), .b(G770), .O(G794) );
nand2 gate266( .a(G645), .b(G773), .O(G797) );
nand2 gate267( .a(G648), .b(G776), .O(G800) );
nand2 gate268( .a(G651), .b(G779), .O(G803) );
nand2 gate269( .a(G654), .b(G782), .O(G806) );

  xor2  gate701(.a(G785), .b(G657), .O(gate270inter0));
  nand2 gate702(.a(gate270inter0), .b(s_22), .O(gate270inter1));
  and2  gate703(.a(G785), .b(G657), .O(gate270inter2));
  inv1  gate704(.a(s_22), .O(gate270inter3));
  inv1  gate705(.a(s_23), .O(gate270inter4));
  nand2 gate706(.a(gate270inter4), .b(gate270inter3), .O(gate270inter5));
  nor2  gate707(.a(gate270inter5), .b(gate270inter2), .O(gate270inter6));
  inv1  gate708(.a(G657), .O(gate270inter7));
  inv1  gate709(.a(G785), .O(gate270inter8));
  nand2 gate710(.a(gate270inter8), .b(gate270inter7), .O(gate270inter9));
  nand2 gate711(.a(s_23), .b(gate270inter3), .O(gate270inter10));
  nor2  gate712(.a(gate270inter10), .b(gate270inter9), .O(gate270inter11));
  nor2  gate713(.a(gate270inter11), .b(gate270inter6), .O(gate270inter12));
  nand2 gate714(.a(gate270inter12), .b(gate270inter1), .O(G809));
nand2 gate271( .a(G660), .b(G788), .O(G812) );
nand2 gate272( .a(G663), .b(G791), .O(G815) );
nand2 gate273( .a(G642), .b(G794), .O(G818) );
nand2 gate274( .a(G770), .b(G794), .O(G819) );
nand2 gate275( .a(G645), .b(G797), .O(G820) );
nand2 gate276( .a(G773), .b(G797), .O(G821) );
nand2 gate277( .a(G648), .b(G800), .O(G822) );
nand2 gate278( .a(G776), .b(G800), .O(G823) );
nand2 gate279( .a(G651), .b(G803), .O(G824) );
nand2 gate280( .a(G779), .b(G803), .O(G825) );
nand2 gate281( .a(G654), .b(G806), .O(G826) );
nand2 gate282( .a(G782), .b(G806), .O(G827) );
nand2 gate283( .a(G657), .b(G809), .O(G828) );
nand2 gate284( .a(G785), .b(G809), .O(G829) );
nand2 gate285( .a(G660), .b(G812), .O(G830) );
nand2 gate286( .a(G788), .b(G812), .O(G831) );
nand2 gate287( .a(G663), .b(G815), .O(G832) );
nand2 gate288( .a(G791), .b(G815), .O(G833) );

  xor2  gate757(.a(G819), .b(G818), .O(gate289inter0));
  nand2 gate758(.a(gate289inter0), .b(s_30), .O(gate289inter1));
  and2  gate759(.a(G819), .b(G818), .O(gate289inter2));
  inv1  gate760(.a(s_30), .O(gate289inter3));
  inv1  gate761(.a(s_31), .O(gate289inter4));
  nand2 gate762(.a(gate289inter4), .b(gate289inter3), .O(gate289inter5));
  nor2  gate763(.a(gate289inter5), .b(gate289inter2), .O(gate289inter6));
  inv1  gate764(.a(G818), .O(gate289inter7));
  inv1  gate765(.a(G819), .O(gate289inter8));
  nand2 gate766(.a(gate289inter8), .b(gate289inter7), .O(gate289inter9));
  nand2 gate767(.a(s_31), .b(gate289inter3), .O(gate289inter10));
  nor2  gate768(.a(gate289inter10), .b(gate289inter9), .O(gate289inter11));
  nor2  gate769(.a(gate289inter11), .b(gate289inter6), .O(gate289inter12));
  nand2 gate770(.a(gate289inter12), .b(gate289inter1), .O(G834));
nand2 gate290( .a(G820), .b(G821), .O(G847) );

  xor2  gate2171(.a(G823), .b(G822), .O(gate291inter0));
  nand2 gate2172(.a(gate291inter0), .b(s_232), .O(gate291inter1));
  and2  gate2173(.a(G823), .b(G822), .O(gate291inter2));
  inv1  gate2174(.a(s_232), .O(gate291inter3));
  inv1  gate2175(.a(s_233), .O(gate291inter4));
  nand2 gate2176(.a(gate291inter4), .b(gate291inter3), .O(gate291inter5));
  nor2  gate2177(.a(gate291inter5), .b(gate291inter2), .O(gate291inter6));
  inv1  gate2178(.a(G822), .O(gate291inter7));
  inv1  gate2179(.a(G823), .O(gate291inter8));
  nand2 gate2180(.a(gate291inter8), .b(gate291inter7), .O(gate291inter9));
  nand2 gate2181(.a(s_233), .b(gate291inter3), .O(gate291inter10));
  nor2  gate2182(.a(gate291inter10), .b(gate291inter9), .O(gate291inter11));
  nor2  gate2183(.a(gate291inter11), .b(gate291inter6), .O(gate291inter12));
  nand2 gate2184(.a(gate291inter12), .b(gate291inter1), .O(G860));
nand2 gate292( .a(G824), .b(G825), .O(G873) );
nand2 gate293( .a(G828), .b(G829), .O(G886) );

  xor2  gate2353(.a(G833), .b(G832), .O(gate294inter0));
  nand2 gate2354(.a(gate294inter0), .b(s_258), .O(gate294inter1));
  and2  gate2355(.a(G833), .b(G832), .O(gate294inter2));
  inv1  gate2356(.a(s_258), .O(gate294inter3));
  inv1  gate2357(.a(s_259), .O(gate294inter4));
  nand2 gate2358(.a(gate294inter4), .b(gate294inter3), .O(gate294inter5));
  nor2  gate2359(.a(gate294inter5), .b(gate294inter2), .O(gate294inter6));
  inv1  gate2360(.a(G832), .O(gate294inter7));
  inv1  gate2361(.a(G833), .O(gate294inter8));
  nand2 gate2362(.a(gate294inter8), .b(gate294inter7), .O(gate294inter9));
  nand2 gate2363(.a(s_259), .b(gate294inter3), .O(gate294inter10));
  nor2  gate2364(.a(gate294inter10), .b(gate294inter9), .O(gate294inter11));
  nor2  gate2365(.a(gate294inter11), .b(gate294inter6), .O(gate294inter12));
  nand2 gate2366(.a(gate294inter12), .b(gate294inter1), .O(G899));
nand2 gate295( .a(G830), .b(G831), .O(G912) );
nand2 gate296( .a(G826), .b(G827), .O(G925) );
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );
nand2 gate387( .a(G1), .b(G1036), .O(G1132) );

  xor2  gate1387(.a(G1039), .b(G2), .O(gate388inter0));
  nand2 gate1388(.a(gate388inter0), .b(s_120), .O(gate388inter1));
  and2  gate1389(.a(G1039), .b(G2), .O(gate388inter2));
  inv1  gate1390(.a(s_120), .O(gate388inter3));
  inv1  gate1391(.a(s_121), .O(gate388inter4));
  nand2 gate1392(.a(gate388inter4), .b(gate388inter3), .O(gate388inter5));
  nor2  gate1393(.a(gate388inter5), .b(gate388inter2), .O(gate388inter6));
  inv1  gate1394(.a(G2), .O(gate388inter7));
  inv1  gate1395(.a(G1039), .O(gate388inter8));
  nand2 gate1396(.a(gate388inter8), .b(gate388inter7), .O(gate388inter9));
  nand2 gate1397(.a(s_121), .b(gate388inter3), .O(gate388inter10));
  nor2  gate1398(.a(gate388inter10), .b(gate388inter9), .O(gate388inter11));
  nor2  gate1399(.a(gate388inter11), .b(gate388inter6), .O(gate388inter12));
  nand2 gate1400(.a(gate388inter12), .b(gate388inter1), .O(G1135));

  xor2  gate1779(.a(G1042), .b(G3), .O(gate389inter0));
  nand2 gate1780(.a(gate389inter0), .b(s_176), .O(gate389inter1));
  and2  gate1781(.a(G1042), .b(G3), .O(gate389inter2));
  inv1  gate1782(.a(s_176), .O(gate389inter3));
  inv1  gate1783(.a(s_177), .O(gate389inter4));
  nand2 gate1784(.a(gate389inter4), .b(gate389inter3), .O(gate389inter5));
  nor2  gate1785(.a(gate389inter5), .b(gate389inter2), .O(gate389inter6));
  inv1  gate1786(.a(G3), .O(gate389inter7));
  inv1  gate1787(.a(G1042), .O(gate389inter8));
  nand2 gate1788(.a(gate389inter8), .b(gate389inter7), .O(gate389inter9));
  nand2 gate1789(.a(s_177), .b(gate389inter3), .O(gate389inter10));
  nor2  gate1790(.a(gate389inter10), .b(gate389inter9), .O(gate389inter11));
  nor2  gate1791(.a(gate389inter11), .b(gate389inter6), .O(gate389inter12));
  nand2 gate1792(.a(gate389inter12), .b(gate389inter1), .O(G1138));

  xor2  gate687(.a(G1045), .b(G4), .O(gate390inter0));
  nand2 gate688(.a(gate390inter0), .b(s_20), .O(gate390inter1));
  and2  gate689(.a(G1045), .b(G4), .O(gate390inter2));
  inv1  gate690(.a(s_20), .O(gate390inter3));
  inv1  gate691(.a(s_21), .O(gate390inter4));
  nand2 gate692(.a(gate390inter4), .b(gate390inter3), .O(gate390inter5));
  nor2  gate693(.a(gate390inter5), .b(gate390inter2), .O(gate390inter6));
  inv1  gate694(.a(G4), .O(gate390inter7));
  inv1  gate695(.a(G1045), .O(gate390inter8));
  nand2 gate696(.a(gate390inter8), .b(gate390inter7), .O(gate390inter9));
  nand2 gate697(.a(s_21), .b(gate390inter3), .O(gate390inter10));
  nor2  gate698(.a(gate390inter10), .b(gate390inter9), .O(gate390inter11));
  nor2  gate699(.a(gate390inter11), .b(gate390inter6), .O(gate390inter12));
  nand2 gate700(.a(gate390inter12), .b(gate390inter1), .O(G1141));

  xor2  gate2437(.a(G1048), .b(G5), .O(gate391inter0));
  nand2 gate2438(.a(gate391inter0), .b(s_270), .O(gate391inter1));
  and2  gate2439(.a(G1048), .b(G5), .O(gate391inter2));
  inv1  gate2440(.a(s_270), .O(gate391inter3));
  inv1  gate2441(.a(s_271), .O(gate391inter4));
  nand2 gate2442(.a(gate391inter4), .b(gate391inter3), .O(gate391inter5));
  nor2  gate2443(.a(gate391inter5), .b(gate391inter2), .O(gate391inter6));
  inv1  gate2444(.a(G5), .O(gate391inter7));
  inv1  gate2445(.a(G1048), .O(gate391inter8));
  nand2 gate2446(.a(gate391inter8), .b(gate391inter7), .O(gate391inter9));
  nand2 gate2447(.a(s_271), .b(gate391inter3), .O(gate391inter10));
  nor2  gate2448(.a(gate391inter10), .b(gate391inter9), .O(gate391inter11));
  nor2  gate2449(.a(gate391inter11), .b(gate391inter6), .O(gate391inter12));
  nand2 gate2450(.a(gate391inter12), .b(gate391inter1), .O(G1144));
nand2 gate392( .a(G6), .b(G1051), .O(G1147) );
nand2 gate393( .a(G7), .b(G1054), .O(G1150) );
nand2 gate394( .a(G8), .b(G1057), .O(G1153) );

  xor2  gate1821(.a(G1060), .b(G9), .O(gate395inter0));
  nand2 gate1822(.a(gate395inter0), .b(s_182), .O(gate395inter1));
  and2  gate1823(.a(G1060), .b(G9), .O(gate395inter2));
  inv1  gate1824(.a(s_182), .O(gate395inter3));
  inv1  gate1825(.a(s_183), .O(gate395inter4));
  nand2 gate1826(.a(gate395inter4), .b(gate395inter3), .O(gate395inter5));
  nor2  gate1827(.a(gate395inter5), .b(gate395inter2), .O(gate395inter6));
  inv1  gate1828(.a(G9), .O(gate395inter7));
  inv1  gate1829(.a(G1060), .O(gate395inter8));
  nand2 gate1830(.a(gate395inter8), .b(gate395inter7), .O(gate395inter9));
  nand2 gate1831(.a(s_183), .b(gate395inter3), .O(gate395inter10));
  nor2  gate1832(.a(gate395inter10), .b(gate395inter9), .O(gate395inter11));
  nor2  gate1833(.a(gate395inter11), .b(gate395inter6), .O(gate395inter12));
  nand2 gate1834(.a(gate395inter12), .b(gate395inter1), .O(G1156));
nand2 gate396( .a(G10), .b(G1063), .O(G1159) );
nand2 gate397( .a(G11), .b(G1066), .O(G1162) );
nand2 gate398( .a(G12), .b(G1069), .O(G1165) );
nand2 gate399( .a(G13), .b(G1072), .O(G1168) );
nand2 gate400( .a(G14), .b(G1075), .O(G1171) );

  xor2  gate2395(.a(G1078), .b(G15), .O(gate401inter0));
  nand2 gate2396(.a(gate401inter0), .b(s_264), .O(gate401inter1));
  and2  gate2397(.a(G1078), .b(G15), .O(gate401inter2));
  inv1  gate2398(.a(s_264), .O(gate401inter3));
  inv1  gate2399(.a(s_265), .O(gate401inter4));
  nand2 gate2400(.a(gate401inter4), .b(gate401inter3), .O(gate401inter5));
  nor2  gate2401(.a(gate401inter5), .b(gate401inter2), .O(gate401inter6));
  inv1  gate2402(.a(G15), .O(gate401inter7));
  inv1  gate2403(.a(G1078), .O(gate401inter8));
  nand2 gate2404(.a(gate401inter8), .b(gate401inter7), .O(gate401inter9));
  nand2 gate2405(.a(s_265), .b(gate401inter3), .O(gate401inter10));
  nor2  gate2406(.a(gate401inter10), .b(gate401inter9), .O(gate401inter11));
  nor2  gate2407(.a(gate401inter11), .b(gate401inter6), .O(gate401inter12));
  nand2 gate2408(.a(gate401inter12), .b(gate401inter1), .O(G1174));
nand2 gate402( .a(G16), .b(G1081), .O(G1177) );

  xor2  gate1625(.a(G1084), .b(G17), .O(gate403inter0));
  nand2 gate1626(.a(gate403inter0), .b(s_154), .O(gate403inter1));
  and2  gate1627(.a(G1084), .b(G17), .O(gate403inter2));
  inv1  gate1628(.a(s_154), .O(gate403inter3));
  inv1  gate1629(.a(s_155), .O(gate403inter4));
  nand2 gate1630(.a(gate403inter4), .b(gate403inter3), .O(gate403inter5));
  nor2  gate1631(.a(gate403inter5), .b(gate403inter2), .O(gate403inter6));
  inv1  gate1632(.a(G17), .O(gate403inter7));
  inv1  gate1633(.a(G1084), .O(gate403inter8));
  nand2 gate1634(.a(gate403inter8), .b(gate403inter7), .O(gate403inter9));
  nand2 gate1635(.a(s_155), .b(gate403inter3), .O(gate403inter10));
  nor2  gate1636(.a(gate403inter10), .b(gate403inter9), .O(gate403inter11));
  nor2  gate1637(.a(gate403inter11), .b(gate403inter6), .O(gate403inter12));
  nand2 gate1638(.a(gate403inter12), .b(gate403inter1), .O(G1180));

  xor2  gate2367(.a(G1087), .b(G18), .O(gate404inter0));
  nand2 gate2368(.a(gate404inter0), .b(s_260), .O(gate404inter1));
  and2  gate2369(.a(G1087), .b(G18), .O(gate404inter2));
  inv1  gate2370(.a(s_260), .O(gate404inter3));
  inv1  gate2371(.a(s_261), .O(gate404inter4));
  nand2 gate2372(.a(gate404inter4), .b(gate404inter3), .O(gate404inter5));
  nor2  gate2373(.a(gate404inter5), .b(gate404inter2), .O(gate404inter6));
  inv1  gate2374(.a(G18), .O(gate404inter7));
  inv1  gate2375(.a(G1087), .O(gate404inter8));
  nand2 gate2376(.a(gate404inter8), .b(gate404inter7), .O(gate404inter9));
  nand2 gate2377(.a(s_261), .b(gate404inter3), .O(gate404inter10));
  nor2  gate2378(.a(gate404inter10), .b(gate404inter9), .O(gate404inter11));
  nor2  gate2379(.a(gate404inter11), .b(gate404inter6), .O(gate404inter12));
  nand2 gate2380(.a(gate404inter12), .b(gate404inter1), .O(G1183));
nand2 gate405( .a(G19), .b(G1090), .O(G1186) );
nand2 gate406( .a(G20), .b(G1093), .O(G1189) );

  xor2  gate2213(.a(G1096), .b(G21), .O(gate407inter0));
  nand2 gate2214(.a(gate407inter0), .b(s_238), .O(gate407inter1));
  and2  gate2215(.a(G1096), .b(G21), .O(gate407inter2));
  inv1  gate2216(.a(s_238), .O(gate407inter3));
  inv1  gate2217(.a(s_239), .O(gate407inter4));
  nand2 gate2218(.a(gate407inter4), .b(gate407inter3), .O(gate407inter5));
  nor2  gate2219(.a(gate407inter5), .b(gate407inter2), .O(gate407inter6));
  inv1  gate2220(.a(G21), .O(gate407inter7));
  inv1  gate2221(.a(G1096), .O(gate407inter8));
  nand2 gate2222(.a(gate407inter8), .b(gate407inter7), .O(gate407inter9));
  nand2 gate2223(.a(s_239), .b(gate407inter3), .O(gate407inter10));
  nor2  gate2224(.a(gate407inter10), .b(gate407inter9), .O(gate407inter11));
  nor2  gate2225(.a(gate407inter11), .b(gate407inter6), .O(gate407inter12));
  nand2 gate2226(.a(gate407inter12), .b(gate407inter1), .O(G1192));
nand2 gate408( .a(G22), .b(G1099), .O(G1195) );
nand2 gate409( .a(G23), .b(G1102), .O(G1198) );
nand2 gate410( .a(G24), .b(G1105), .O(G1201) );
nand2 gate411( .a(G25), .b(G1108), .O(G1204) );
nand2 gate412( .a(G26), .b(G1111), .O(G1207) );
nand2 gate413( .a(G27), .b(G1114), .O(G1210) );

  xor2  gate1443(.a(G1117), .b(G28), .O(gate414inter0));
  nand2 gate1444(.a(gate414inter0), .b(s_128), .O(gate414inter1));
  and2  gate1445(.a(G1117), .b(G28), .O(gate414inter2));
  inv1  gate1446(.a(s_128), .O(gate414inter3));
  inv1  gate1447(.a(s_129), .O(gate414inter4));
  nand2 gate1448(.a(gate414inter4), .b(gate414inter3), .O(gate414inter5));
  nor2  gate1449(.a(gate414inter5), .b(gate414inter2), .O(gate414inter6));
  inv1  gate1450(.a(G28), .O(gate414inter7));
  inv1  gate1451(.a(G1117), .O(gate414inter8));
  nand2 gate1452(.a(gate414inter8), .b(gate414inter7), .O(gate414inter9));
  nand2 gate1453(.a(s_129), .b(gate414inter3), .O(gate414inter10));
  nor2  gate1454(.a(gate414inter10), .b(gate414inter9), .O(gate414inter11));
  nor2  gate1455(.a(gate414inter11), .b(gate414inter6), .O(gate414inter12));
  nand2 gate1456(.a(gate414inter12), .b(gate414inter1), .O(G1213));
nand2 gate415( .a(G29), .b(G1120), .O(G1216) );
nand2 gate416( .a(G30), .b(G1123), .O(G1219) );
nand2 gate417( .a(G31), .b(G1126), .O(G1222) );
nand2 gate418( .a(G32), .b(G1129), .O(G1225) );
nand2 gate419( .a(G1), .b(G1132), .O(G1228) );
nand2 gate420( .a(G1036), .b(G1132), .O(G1229) );

  xor2  gate2199(.a(G1135), .b(G2), .O(gate421inter0));
  nand2 gate2200(.a(gate421inter0), .b(s_236), .O(gate421inter1));
  and2  gate2201(.a(G1135), .b(G2), .O(gate421inter2));
  inv1  gate2202(.a(s_236), .O(gate421inter3));
  inv1  gate2203(.a(s_237), .O(gate421inter4));
  nand2 gate2204(.a(gate421inter4), .b(gate421inter3), .O(gate421inter5));
  nor2  gate2205(.a(gate421inter5), .b(gate421inter2), .O(gate421inter6));
  inv1  gate2206(.a(G2), .O(gate421inter7));
  inv1  gate2207(.a(G1135), .O(gate421inter8));
  nand2 gate2208(.a(gate421inter8), .b(gate421inter7), .O(gate421inter9));
  nand2 gate2209(.a(s_237), .b(gate421inter3), .O(gate421inter10));
  nor2  gate2210(.a(gate421inter10), .b(gate421inter9), .O(gate421inter11));
  nor2  gate2211(.a(gate421inter11), .b(gate421inter6), .O(gate421inter12));
  nand2 gate2212(.a(gate421inter12), .b(gate421inter1), .O(G1230));
nand2 gate422( .a(G1039), .b(G1135), .O(G1231) );
nand2 gate423( .a(G3), .b(G1138), .O(G1232) );
nand2 gate424( .a(G1042), .b(G1138), .O(G1233) );
nand2 gate425( .a(G4), .b(G1141), .O(G1234) );

  xor2  gate2227(.a(G1141), .b(G1045), .O(gate426inter0));
  nand2 gate2228(.a(gate426inter0), .b(s_240), .O(gate426inter1));
  and2  gate2229(.a(G1141), .b(G1045), .O(gate426inter2));
  inv1  gate2230(.a(s_240), .O(gate426inter3));
  inv1  gate2231(.a(s_241), .O(gate426inter4));
  nand2 gate2232(.a(gate426inter4), .b(gate426inter3), .O(gate426inter5));
  nor2  gate2233(.a(gate426inter5), .b(gate426inter2), .O(gate426inter6));
  inv1  gate2234(.a(G1045), .O(gate426inter7));
  inv1  gate2235(.a(G1141), .O(gate426inter8));
  nand2 gate2236(.a(gate426inter8), .b(gate426inter7), .O(gate426inter9));
  nand2 gate2237(.a(s_241), .b(gate426inter3), .O(gate426inter10));
  nor2  gate2238(.a(gate426inter10), .b(gate426inter9), .O(gate426inter11));
  nor2  gate2239(.a(gate426inter11), .b(gate426inter6), .O(gate426inter12));
  nand2 gate2240(.a(gate426inter12), .b(gate426inter1), .O(G1235));
nand2 gate427( .a(G5), .b(G1144), .O(G1236) );

  xor2  gate883(.a(G1144), .b(G1048), .O(gate428inter0));
  nand2 gate884(.a(gate428inter0), .b(s_48), .O(gate428inter1));
  and2  gate885(.a(G1144), .b(G1048), .O(gate428inter2));
  inv1  gate886(.a(s_48), .O(gate428inter3));
  inv1  gate887(.a(s_49), .O(gate428inter4));
  nand2 gate888(.a(gate428inter4), .b(gate428inter3), .O(gate428inter5));
  nor2  gate889(.a(gate428inter5), .b(gate428inter2), .O(gate428inter6));
  inv1  gate890(.a(G1048), .O(gate428inter7));
  inv1  gate891(.a(G1144), .O(gate428inter8));
  nand2 gate892(.a(gate428inter8), .b(gate428inter7), .O(gate428inter9));
  nand2 gate893(.a(s_49), .b(gate428inter3), .O(gate428inter10));
  nor2  gate894(.a(gate428inter10), .b(gate428inter9), .O(gate428inter11));
  nor2  gate895(.a(gate428inter11), .b(gate428inter6), .O(gate428inter12));
  nand2 gate896(.a(gate428inter12), .b(gate428inter1), .O(G1237));
nand2 gate429( .a(G6), .b(G1147), .O(G1238) );
nand2 gate430( .a(G1051), .b(G1147), .O(G1239) );
nand2 gate431( .a(G7), .b(G1150), .O(G1240) );

  xor2  gate1457(.a(G1150), .b(G1054), .O(gate432inter0));
  nand2 gate1458(.a(gate432inter0), .b(s_130), .O(gate432inter1));
  and2  gate1459(.a(G1150), .b(G1054), .O(gate432inter2));
  inv1  gate1460(.a(s_130), .O(gate432inter3));
  inv1  gate1461(.a(s_131), .O(gate432inter4));
  nand2 gate1462(.a(gate432inter4), .b(gate432inter3), .O(gate432inter5));
  nor2  gate1463(.a(gate432inter5), .b(gate432inter2), .O(gate432inter6));
  inv1  gate1464(.a(G1054), .O(gate432inter7));
  inv1  gate1465(.a(G1150), .O(gate432inter8));
  nand2 gate1466(.a(gate432inter8), .b(gate432inter7), .O(gate432inter9));
  nand2 gate1467(.a(s_131), .b(gate432inter3), .O(gate432inter10));
  nor2  gate1468(.a(gate432inter10), .b(gate432inter9), .O(gate432inter11));
  nor2  gate1469(.a(gate432inter11), .b(gate432inter6), .O(gate432inter12));
  nand2 gate1470(.a(gate432inter12), .b(gate432inter1), .O(G1241));
nand2 gate433( .a(G8), .b(G1153), .O(G1242) );

  xor2  gate1289(.a(G1153), .b(G1057), .O(gate434inter0));
  nand2 gate1290(.a(gate434inter0), .b(s_106), .O(gate434inter1));
  and2  gate1291(.a(G1153), .b(G1057), .O(gate434inter2));
  inv1  gate1292(.a(s_106), .O(gate434inter3));
  inv1  gate1293(.a(s_107), .O(gate434inter4));
  nand2 gate1294(.a(gate434inter4), .b(gate434inter3), .O(gate434inter5));
  nor2  gate1295(.a(gate434inter5), .b(gate434inter2), .O(gate434inter6));
  inv1  gate1296(.a(G1057), .O(gate434inter7));
  inv1  gate1297(.a(G1153), .O(gate434inter8));
  nand2 gate1298(.a(gate434inter8), .b(gate434inter7), .O(gate434inter9));
  nand2 gate1299(.a(s_107), .b(gate434inter3), .O(gate434inter10));
  nor2  gate1300(.a(gate434inter10), .b(gate434inter9), .O(gate434inter11));
  nor2  gate1301(.a(gate434inter11), .b(gate434inter6), .O(gate434inter12));
  nand2 gate1302(.a(gate434inter12), .b(gate434inter1), .O(G1243));

  xor2  gate1149(.a(G1156), .b(G9), .O(gate435inter0));
  nand2 gate1150(.a(gate435inter0), .b(s_86), .O(gate435inter1));
  and2  gate1151(.a(G1156), .b(G9), .O(gate435inter2));
  inv1  gate1152(.a(s_86), .O(gate435inter3));
  inv1  gate1153(.a(s_87), .O(gate435inter4));
  nand2 gate1154(.a(gate435inter4), .b(gate435inter3), .O(gate435inter5));
  nor2  gate1155(.a(gate435inter5), .b(gate435inter2), .O(gate435inter6));
  inv1  gate1156(.a(G9), .O(gate435inter7));
  inv1  gate1157(.a(G1156), .O(gate435inter8));
  nand2 gate1158(.a(gate435inter8), .b(gate435inter7), .O(gate435inter9));
  nand2 gate1159(.a(s_87), .b(gate435inter3), .O(gate435inter10));
  nor2  gate1160(.a(gate435inter10), .b(gate435inter9), .O(gate435inter11));
  nor2  gate1161(.a(gate435inter11), .b(gate435inter6), .O(gate435inter12));
  nand2 gate1162(.a(gate435inter12), .b(gate435inter1), .O(G1244));

  xor2  gate1555(.a(G1156), .b(G1060), .O(gate436inter0));
  nand2 gate1556(.a(gate436inter0), .b(s_144), .O(gate436inter1));
  and2  gate1557(.a(G1156), .b(G1060), .O(gate436inter2));
  inv1  gate1558(.a(s_144), .O(gate436inter3));
  inv1  gate1559(.a(s_145), .O(gate436inter4));
  nand2 gate1560(.a(gate436inter4), .b(gate436inter3), .O(gate436inter5));
  nor2  gate1561(.a(gate436inter5), .b(gate436inter2), .O(gate436inter6));
  inv1  gate1562(.a(G1060), .O(gate436inter7));
  inv1  gate1563(.a(G1156), .O(gate436inter8));
  nand2 gate1564(.a(gate436inter8), .b(gate436inter7), .O(gate436inter9));
  nand2 gate1565(.a(s_145), .b(gate436inter3), .O(gate436inter10));
  nor2  gate1566(.a(gate436inter10), .b(gate436inter9), .O(gate436inter11));
  nor2  gate1567(.a(gate436inter11), .b(gate436inter6), .O(gate436inter12));
  nand2 gate1568(.a(gate436inter12), .b(gate436inter1), .O(G1245));
nand2 gate437( .a(G10), .b(G1159), .O(G1246) );
nand2 gate438( .a(G1063), .b(G1159), .O(G1247) );

  xor2  gate1765(.a(G1162), .b(G11), .O(gate439inter0));
  nand2 gate1766(.a(gate439inter0), .b(s_174), .O(gate439inter1));
  and2  gate1767(.a(G1162), .b(G11), .O(gate439inter2));
  inv1  gate1768(.a(s_174), .O(gate439inter3));
  inv1  gate1769(.a(s_175), .O(gate439inter4));
  nand2 gate1770(.a(gate439inter4), .b(gate439inter3), .O(gate439inter5));
  nor2  gate1771(.a(gate439inter5), .b(gate439inter2), .O(gate439inter6));
  inv1  gate1772(.a(G11), .O(gate439inter7));
  inv1  gate1773(.a(G1162), .O(gate439inter8));
  nand2 gate1774(.a(gate439inter8), .b(gate439inter7), .O(gate439inter9));
  nand2 gate1775(.a(s_175), .b(gate439inter3), .O(gate439inter10));
  nor2  gate1776(.a(gate439inter10), .b(gate439inter9), .O(gate439inter11));
  nor2  gate1777(.a(gate439inter11), .b(gate439inter6), .O(gate439inter12));
  nand2 gate1778(.a(gate439inter12), .b(gate439inter1), .O(G1248));

  xor2  gate1863(.a(G1162), .b(G1066), .O(gate440inter0));
  nand2 gate1864(.a(gate440inter0), .b(s_188), .O(gate440inter1));
  and2  gate1865(.a(G1162), .b(G1066), .O(gate440inter2));
  inv1  gate1866(.a(s_188), .O(gate440inter3));
  inv1  gate1867(.a(s_189), .O(gate440inter4));
  nand2 gate1868(.a(gate440inter4), .b(gate440inter3), .O(gate440inter5));
  nor2  gate1869(.a(gate440inter5), .b(gate440inter2), .O(gate440inter6));
  inv1  gate1870(.a(G1066), .O(gate440inter7));
  inv1  gate1871(.a(G1162), .O(gate440inter8));
  nand2 gate1872(.a(gate440inter8), .b(gate440inter7), .O(gate440inter9));
  nand2 gate1873(.a(s_189), .b(gate440inter3), .O(gate440inter10));
  nor2  gate1874(.a(gate440inter10), .b(gate440inter9), .O(gate440inter11));
  nor2  gate1875(.a(gate440inter11), .b(gate440inter6), .O(gate440inter12));
  nand2 gate1876(.a(gate440inter12), .b(gate440inter1), .O(G1249));
nand2 gate441( .a(G12), .b(G1165), .O(G1250) );
nand2 gate442( .a(G1069), .b(G1165), .O(G1251) );
nand2 gate443( .a(G13), .b(G1168), .O(G1252) );
nand2 gate444( .a(G1072), .b(G1168), .O(G1253) );

  xor2  gate1541(.a(G1171), .b(G14), .O(gate445inter0));
  nand2 gate1542(.a(gate445inter0), .b(s_142), .O(gate445inter1));
  and2  gate1543(.a(G1171), .b(G14), .O(gate445inter2));
  inv1  gate1544(.a(s_142), .O(gate445inter3));
  inv1  gate1545(.a(s_143), .O(gate445inter4));
  nand2 gate1546(.a(gate445inter4), .b(gate445inter3), .O(gate445inter5));
  nor2  gate1547(.a(gate445inter5), .b(gate445inter2), .O(gate445inter6));
  inv1  gate1548(.a(G14), .O(gate445inter7));
  inv1  gate1549(.a(G1171), .O(gate445inter8));
  nand2 gate1550(.a(gate445inter8), .b(gate445inter7), .O(gate445inter9));
  nand2 gate1551(.a(s_143), .b(gate445inter3), .O(gate445inter10));
  nor2  gate1552(.a(gate445inter10), .b(gate445inter9), .O(gate445inter11));
  nor2  gate1553(.a(gate445inter11), .b(gate445inter6), .O(gate445inter12));
  nand2 gate1554(.a(gate445inter12), .b(gate445inter1), .O(G1254));
nand2 gate446( .a(G1075), .b(G1171), .O(G1255) );
nand2 gate447( .a(G15), .b(G1174), .O(G1256) );
nand2 gate448( .a(G1078), .b(G1174), .O(G1257) );
nand2 gate449( .a(G16), .b(G1177), .O(G1258) );
nand2 gate450( .a(G1081), .b(G1177), .O(G1259) );
nand2 gate451( .a(G17), .b(G1180), .O(G1260) );
nand2 gate452( .a(G1084), .b(G1180), .O(G1261) );

  xor2  gate2283(.a(G1183), .b(G18), .O(gate453inter0));
  nand2 gate2284(.a(gate453inter0), .b(s_248), .O(gate453inter1));
  and2  gate2285(.a(G1183), .b(G18), .O(gate453inter2));
  inv1  gate2286(.a(s_248), .O(gate453inter3));
  inv1  gate2287(.a(s_249), .O(gate453inter4));
  nand2 gate2288(.a(gate453inter4), .b(gate453inter3), .O(gate453inter5));
  nor2  gate2289(.a(gate453inter5), .b(gate453inter2), .O(gate453inter6));
  inv1  gate2290(.a(G18), .O(gate453inter7));
  inv1  gate2291(.a(G1183), .O(gate453inter8));
  nand2 gate2292(.a(gate453inter8), .b(gate453inter7), .O(gate453inter9));
  nand2 gate2293(.a(s_249), .b(gate453inter3), .O(gate453inter10));
  nor2  gate2294(.a(gate453inter10), .b(gate453inter9), .O(gate453inter11));
  nor2  gate2295(.a(gate453inter11), .b(gate453inter6), .O(gate453inter12));
  nand2 gate2296(.a(gate453inter12), .b(gate453inter1), .O(G1262));

  xor2  gate547(.a(G1183), .b(G1087), .O(gate454inter0));
  nand2 gate548(.a(gate454inter0), .b(s_0), .O(gate454inter1));
  and2  gate549(.a(G1183), .b(G1087), .O(gate454inter2));
  inv1  gate550(.a(s_0), .O(gate454inter3));
  inv1  gate551(.a(s_1), .O(gate454inter4));
  nand2 gate552(.a(gate454inter4), .b(gate454inter3), .O(gate454inter5));
  nor2  gate553(.a(gate454inter5), .b(gate454inter2), .O(gate454inter6));
  inv1  gate554(.a(G1087), .O(gate454inter7));
  inv1  gate555(.a(G1183), .O(gate454inter8));
  nand2 gate556(.a(gate454inter8), .b(gate454inter7), .O(gate454inter9));
  nand2 gate557(.a(s_1), .b(gate454inter3), .O(gate454inter10));
  nor2  gate558(.a(gate454inter10), .b(gate454inter9), .O(gate454inter11));
  nor2  gate559(.a(gate454inter11), .b(gate454inter6), .O(gate454inter12));
  nand2 gate560(.a(gate454inter12), .b(gate454inter1), .O(G1263));
nand2 gate455( .a(G19), .b(G1186), .O(G1264) );
nand2 gate456( .a(G1090), .b(G1186), .O(G1265) );
nand2 gate457( .a(G20), .b(G1189), .O(G1266) );
nand2 gate458( .a(G1093), .b(G1189), .O(G1267) );

  xor2  gate1961(.a(G1192), .b(G21), .O(gate459inter0));
  nand2 gate1962(.a(gate459inter0), .b(s_202), .O(gate459inter1));
  and2  gate1963(.a(G1192), .b(G21), .O(gate459inter2));
  inv1  gate1964(.a(s_202), .O(gate459inter3));
  inv1  gate1965(.a(s_203), .O(gate459inter4));
  nand2 gate1966(.a(gate459inter4), .b(gate459inter3), .O(gate459inter5));
  nor2  gate1967(.a(gate459inter5), .b(gate459inter2), .O(gate459inter6));
  inv1  gate1968(.a(G21), .O(gate459inter7));
  inv1  gate1969(.a(G1192), .O(gate459inter8));
  nand2 gate1970(.a(gate459inter8), .b(gate459inter7), .O(gate459inter9));
  nand2 gate1971(.a(s_203), .b(gate459inter3), .O(gate459inter10));
  nor2  gate1972(.a(gate459inter10), .b(gate459inter9), .O(gate459inter11));
  nor2  gate1973(.a(gate459inter11), .b(gate459inter6), .O(gate459inter12));
  nand2 gate1974(.a(gate459inter12), .b(gate459inter1), .O(G1268));
nand2 gate460( .a(G1096), .b(G1192), .O(G1269) );
nand2 gate461( .a(G22), .b(G1195), .O(G1270) );
nand2 gate462( .a(G1099), .b(G1195), .O(G1271) );

  xor2  gate1471(.a(G1198), .b(G23), .O(gate463inter0));
  nand2 gate1472(.a(gate463inter0), .b(s_132), .O(gate463inter1));
  and2  gate1473(.a(G1198), .b(G23), .O(gate463inter2));
  inv1  gate1474(.a(s_132), .O(gate463inter3));
  inv1  gate1475(.a(s_133), .O(gate463inter4));
  nand2 gate1476(.a(gate463inter4), .b(gate463inter3), .O(gate463inter5));
  nor2  gate1477(.a(gate463inter5), .b(gate463inter2), .O(gate463inter6));
  inv1  gate1478(.a(G23), .O(gate463inter7));
  inv1  gate1479(.a(G1198), .O(gate463inter8));
  nand2 gate1480(.a(gate463inter8), .b(gate463inter7), .O(gate463inter9));
  nand2 gate1481(.a(s_133), .b(gate463inter3), .O(gate463inter10));
  nor2  gate1482(.a(gate463inter10), .b(gate463inter9), .O(gate463inter11));
  nor2  gate1483(.a(gate463inter11), .b(gate463inter6), .O(gate463inter12));
  nand2 gate1484(.a(gate463inter12), .b(gate463inter1), .O(G1272));
nand2 gate464( .a(G1102), .b(G1198), .O(G1273) );

  xor2  gate715(.a(G1201), .b(G24), .O(gate465inter0));
  nand2 gate716(.a(gate465inter0), .b(s_24), .O(gate465inter1));
  and2  gate717(.a(G1201), .b(G24), .O(gate465inter2));
  inv1  gate718(.a(s_24), .O(gate465inter3));
  inv1  gate719(.a(s_25), .O(gate465inter4));
  nand2 gate720(.a(gate465inter4), .b(gate465inter3), .O(gate465inter5));
  nor2  gate721(.a(gate465inter5), .b(gate465inter2), .O(gate465inter6));
  inv1  gate722(.a(G24), .O(gate465inter7));
  inv1  gate723(.a(G1201), .O(gate465inter8));
  nand2 gate724(.a(gate465inter8), .b(gate465inter7), .O(gate465inter9));
  nand2 gate725(.a(s_25), .b(gate465inter3), .O(gate465inter10));
  nor2  gate726(.a(gate465inter10), .b(gate465inter9), .O(gate465inter11));
  nor2  gate727(.a(gate465inter11), .b(gate465inter6), .O(gate465inter12));
  nand2 gate728(.a(gate465inter12), .b(gate465inter1), .O(G1274));
nand2 gate466( .a(G1105), .b(G1201), .O(G1275) );

  xor2  gate785(.a(G1204), .b(G25), .O(gate467inter0));
  nand2 gate786(.a(gate467inter0), .b(s_34), .O(gate467inter1));
  and2  gate787(.a(G1204), .b(G25), .O(gate467inter2));
  inv1  gate788(.a(s_34), .O(gate467inter3));
  inv1  gate789(.a(s_35), .O(gate467inter4));
  nand2 gate790(.a(gate467inter4), .b(gate467inter3), .O(gate467inter5));
  nor2  gate791(.a(gate467inter5), .b(gate467inter2), .O(gate467inter6));
  inv1  gate792(.a(G25), .O(gate467inter7));
  inv1  gate793(.a(G1204), .O(gate467inter8));
  nand2 gate794(.a(gate467inter8), .b(gate467inter7), .O(gate467inter9));
  nand2 gate795(.a(s_35), .b(gate467inter3), .O(gate467inter10));
  nor2  gate796(.a(gate467inter10), .b(gate467inter9), .O(gate467inter11));
  nor2  gate797(.a(gate467inter11), .b(gate467inter6), .O(gate467inter12));
  nand2 gate798(.a(gate467inter12), .b(gate467inter1), .O(G1276));

  xor2  gate911(.a(G1204), .b(G1108), .O(gate468inter0));
  nand2 gate912(.a(gate468inter0), .b(s_52), .O(gate468inter1));
  and2  gate913(.a(G1204), .b(G1108), .O(gate468inter2));
  inv1  gate914(.a(s_52), .O(gate468inter3));
  inv1  gate915(.a(s_53), .O(gate468inter4));
  nand2 gate916(.a(gate468inter4), .b(gate468inter3), .O(gate468inter5));
  nor2  gate917(.a(gate468inter5), .b(gate468inter2), .O(gate468inter6));
  inv1  gate918(.a(G1108), .O(gate468inter7));
  inv1  gate919(.a(G1204), .O(gate468inter8));
  nand2 gate920(.a(gate468inter8), .b(gate468inter7), .O(gate468inter9));
  nand2 gate921(.a(s_53), .b(gate468inter3), .O(gate468inter10));
  nor2  gate922(.a(gate468inter10), .b(gate468inter9), .O(gate468inter11));
  nor2  gate923(.a(gate468inter11), .b(gate468inter6), .O(gate468inter12));
  nand2 gate924(.a(gate468inter12), .b(gate468inter1), .O(G1277));
nand2 gate469( .a(G26), .b(G1207), .O(G1278) );
nand2 gate470( .a(G1111), .b(G1207), .O(G1279) );
nand2 gate471( .a(G27), .b(G1210), .O(G1280) );

  xor2  gate2339(.a(G1210), .b(G1114), .O(gate472inter0));
  nand2 gate2340(.a(gate472inter0), .b(s_256), .O(gate472inter1));
  and2  gate2341(.a(G1210), .b(G1114), .O(gate472inter2));
  inv1  gate2342(.a(s_256), .O(gate472inter3));
  inv1  gate2343(.a(s_257), .O(gate472inter4));
  nand2 gate2344(.a(gate472inter4), .b(gate472inter3), .O(gate472inter5));
  nor2  gate2345(.a(gate472inter5), .b(gate472inter2), .O(gate472inter6));
  inv1  gate2346(.a(G1114), .O(gate472inter7));
  inv1  gate2347(.a(G1210), .O(gate472inter8));
  nand2 gate2348(.a(gate472inter8), .b(gate472inter7), .O(gate472inter9));
  nand2 gate2349(.a(s_257), .b(gate472inter3), .O(gate472inter10));
  nor2  gate2350(.a(gate472inter10), .b(gate472inter9), .O(gate472inter11));
  nor2  gate2351(.a(gate472inter11), .b(gate472inter6), .O(gate472inter12));
  nand2 gate2352(.a(gate472inter12), .b(gate472inter1), .O(G1281));
nand2 gate473( .a(G28), .b(G1213), .O(G1282) );
nand2 gate474( .a(G1117), .b(G1213), .O(G1283) );
nand2 gate475( .a(G29), .b(G1216), .O(G1284) );
nand2 gate476( .a(G1120), .b(G1216), .O(G1285) );

  xor2  gate1513(.a(G1219), .b(G30), .O(gate477inter0));
  nand2 gate1514(.a(gate477inter0), .b(s_138), .O(gate477inter1));
  and2  gate1515(.a(G1219), .b(G30), .O(gate477inter2));
  inv1  gate1516(.a(s_138), .O(gate477inter3));
  inv1  gate1517(.a(s_139), .O(gate477inter4));
  nand2 gate1518(.a(gate477inter4), .b(gate477inter3), .O(gate477inter5));
  nor2  gate1519(.a(gate477inter5), .b(gate477inter2), .O(gate477inter6));
  inv1  gate1520(.a(G30), .O(gate477inter7));
  inv1  gate1521(.a(G1219), .O(gate477inter8));
  nand2 gate1522(.a(gate477inter8), .b(gate477inter7), .O(gate477inter9));
  nand2 gate1523(.a(s_139), .b(gate477inter3), .O(gate477inter10));
  nor2  gate1524(.a(gate477inter10), .b(gate477inter9), .O(gate477inter11));
  nor2  gate1525(.a(gate477inter11), .b(gate477inter6), .O(gate477inter12));
  nand2 gate1526(.a(gate477inter12), .b(gate477inter1), .O(G1286));
nand2 gate478( .a(G1123), .b(G1219), .O(G1287) );
nand2 gate479( .a(G31), .b(G1222), .O(G1288) );
nand2 gate480( .a(G1126), .b(G1222), .O(G1289) );
nand2 gate481( .a(G32), .b(G1225), .O(G1290) );

  xor2  gate1261(.a(G1225), .b(G1129), .O(gate482inter0));
  nand2 gate1262(.a(gate482inter0), .b(s_102), .O(gate482inter1));
  and2  gate1263(.a(G1225), .b(G1129), .O(gate482inter2));
  inv1  gate1264(.a(s_102), .O(gate482inter3));
  inv1  gate1265(.a(s_103), .O(gate482inter4));
  nand2 gate1266(.a(gate482inter4), .b(gate482inter3), .O(gate482inter5));
  nor2  gate1267(.a(gate482inter5), .b(gate482inter2), .O(gate482inter6));
  inv1  gate1268(.a(G1129), .O(gate482inter7));
  inv1  gate1269(.a(G1225), .O(gate482inter8));
  nand2 gate1270(.a(gate482inter8), .b(gate482inter7), .O(gate482inter9));
  nand2 gate1271(.a(s_103), .b(gate482inter3), .O(gate482inter10));
  nor2  gate1272(.a(gate482inter10), .b(gate482inter9), .O(gate482inter11));
  nor2  gate1273(.a(gate482inter11), .b(gate482inter6), .O(gate482inter12));
  nand2 gate1274(.a(gate482inter12), .b(gate482inter1), .O(G1291));

  xor2  gate925(.a(G1229), .b(G1228), .O(gate483inter0));
  nand2 gate926(.a(gate483inter0), .b(s_54), .O(gate483inter1));
  and2  gate927(.a(G1229), .b(G1228), .O(gate483inter2));
  inv1  gate928(.a(s_54), .O(gate483inter3));
  inv1  gate929(.a(s_55), .O(gate483inter4));
  nand2 gate930(.a(gate483inter4), .b(gate483inter3), .O(gate483inter5));
  nor2  gate931(.a(gate483inter5), .b(gate483inter2), .O(gate483inter6));
  inv1  gate932(.a(G1228), .O(gate483inter7));
  inv1  gate933(.a(G1229), .O(gate483inter8));
  nand2 gate934(.a(gate483inter8), .b(gate483inter7), .O(gate483inter9));
  nand2 gate935(.a(s_55), .b(gate483inter3), .O(gate483inter10));
  nor2  gate936(.a(gate483inter10), .b(gate483inter9), .O(gate483inter11));
  nor2  gate937(.a(gate483inter11), .b(gate483inter6), .O(gate483inter12));
  nand2 gate938(.a(gate483inter12), .b(gate483inter1), .O(G1292));
nand2 gate484( .a(G1230), .b(G1231), .O(G1293) );
nand2 gate485( .a(G1232), .b(G1233), .O(G1294) );
nand2 gate486( .a(G1234), .b(G1235), .O(G1295) );

  xor2  gate1751(.a(G1237), .b(G1236), .O(gate487inter0));
  nand2 gate1752(.a(gate487inter0), .b(s_172), .O(gate487inter1));
  and2  gate1753(.a(G1237), .b(G1236), .O(gate487inter2));
  inv1  gate1754(.a(s_172), .O(gate487inter3));
  inv1  gate1755(.a(s_173), .O(gate487inter4));
  nand2 gate1756(.a(gate487inter4), .b(gate487inter3), .O(gate487inter5));
  nor2  gate1757(.a(gate487inter5), .b(gate487inter2), .O(gate487inter6));
  inv1  gate1758(.a(G1236), .O(gate487inter7));
  inv1  gate1759(.a(G1237), .O(gate487inter8));
  nand2 gate1760(.a(gate487inter8), .b(gate487inter7), .O(gate487inter9));
  nand2 gate1761(.a(s_173), .b(gate487inter3), .O(gate487inter10));
  nor2  gate1762(.a(gate487inter10), .b(gate487inter9), .O(gate487inter11));
  nor2  gate1763(.a(gate487inter11), .b(gate487inter6), .O(gate487inter12));
  nand2 gate1764(.a(gate487inter12), .b(gate487inter1), .O(G1296));
nand2 gate488( .a(G1238), .b(G1239), .O(G1297) );
nand2 gate489( .a(G1240), .b(G1241), .O(G1298) );
nand2 gate490( .a(G1242), .b(G1243), .O(G1299) );

  xor2  gate1219(.a(G1245), .b(G1244), .O(gate491inter0));
  nand2 gate1220(.a(gate491inter0), .b(s_96), .O(gate491inter1));
  and2  gate1221(.a(G1245), .b(G1244), .O(gate491inter2));
  inv1  gate1222(.a(s_96), .O(gate491inter3));
  inv1  gate1223(.a(s_97), .O(gate491inter4));
  nand2 gate1224(.a(gate491inter4), .b(gate491inter3), .O(gate491inter5));
  nor2  gate1225(.a(gate491inter5), .b(gate491inter2), .O(gate491inter6));
  inv1  gate1226(.a(G1244), .O(gate491inter7));
  inv1  gate1227(.a(G1245), .O(gate491inter8));
  nand2 gate1228(.a(gate491inter8), .b(gate491inter7), .O(gate491inter9));
  nand2 gate1229(.a(s_97), .b(gate491inter3), .O(gate491inter10));
  nor2  gate1230(.a(gate491inter10), .b(gate491inter9), .O(gate491inter11));
  nor2  gate1231(.a(gate491inter11), .b(gate491inter6), .O(gate491inter12));
  nand2 gate1232(.a(gate491inter12), .b(gate491inter1), .O(G1300));

  xor2  gate841(.a(G1247), .b(G1246), .O(gate492inter0));
  nand2 gate842(.a(gate492inter0), .b(s_42), .O(gate492inter1));
  and2  gate843(.a(G1247), .b(G1246), .O(gate492inter2));
  inv1  gate844(.a(s_42), .O(gate492inter3));
  inv1  gate845(.a(s_43), .O(gate492inter4));
  nand2 gate846(.a(gate492inter4), .b(gate492inter3), .O(gate492inter5));
  nor2  gate847(.a(gate492inter5), .b(gate492inter2), .O(gate492inter6));
  inv1  gate848(.a(G1246), .O(gate492inter7));
  inv1  gate849(.a(G1247), .O(gate492inter8));
  nand2 gate850(.a(gate492inter8), .b(gate492inter7), .O(gate492inter9));
  nand2 gate851(.a(s_43), .b(gate492inter3), .O(gate492inter10));
  nor2  gate852(.a(gate492inter10), .b(gate492inter9), .O(gate492inter11));
  nor2  gate853(.a(gate492inter11), .b(gate492inter6), .O(gate492inter12));
  nand2 gate854(.a(gate492inter12), .b(gate492inter1), .O(G1301));

  xor2  gate2269(.a(G1249), .b(G1248), .O(gate493inter0));
  nand2 gate2270(.a(gate493inter0), .b(s_246), .O(gate493inter1));
  and2  gate2271(.a(G1249), .b(G1248), .O(gate493inter2));
  inv1  gate2272(.a(s_246), .O(gate493inter3));
  inv1  gate2273(.a(s_247), .O(gate493inter4));
  nand2 gate2274(.a(gate493inter4), .b(gate493inter3), .O(gate493inter5));
  nor2  gate2275(.a(gate493inter5), .b(gate493inter2), .O(gate493inter6));
  inv1  gate2276(.a(G1248), .O(gate493inter7));
  inv1  gate2277(.a(G1249), .O(gate493inter8));
  nand2 gate2278(.a(gate493inter8), .b(gate493inter7), .O(gate493inter9));
  nand2 gate2279(.a(s_247), .b(gate493inter3), .O(gate493inter10));
  nor2  gate2280(.a(gate493inter10), .b(gate493inter9), .O(gate493inter11));
  nor2  gate2281(.a(gate493inter11), .b(gate493inter6), .O(gate493inter12));
  nand2 gate2282(.a(gate493inter12), .b(gate493inter1), .O(G1302));

  xor2  gate1807(.a(G1251), .b(G1250), .O(gate494inter0));
  nand2 gate1808(.a(gate494inter0), .b(s_180), .O(gate494inter1));
  and2  gate1809(.a(G1251), .b(G1250), .O(gate494inter2));
  inv1  gate1810(.a(s_180), .O(gate494inter3));
  inv1  gate1811(.a(s_181), .O(gate494inter4));
  nand2 gate1812(.a(gate494inter4), .b(gate494inter3), .O(gate494inter5));
  nor2  gate1813(.a(gate494inter5), .b(gate494inter2), .O(gate494inter6));
  inv1  gate1814(.a(G1250), .O(gate494inter7));
  inv1  gate1815(.a(G1251), .O(gate494inter8));
  nand2 gate1816(.a(gate494inter8), .b(gate494inter7), .O(gate494inter9));
  nand2 gate1817(.a(s_181), .b(gate494inter3), .O(gate494inter10));
  nor2  gate1818(.a(gate494inter10), .b(gate494inter9), .O(gate494inter11));
  nor2  gate1819(.a(gate494inter11), .b(gate494inter6), .O(gate494inter12));
  nand2 gate1820(.a(gate494inter12), .b(gate494inter1), .O(G1303));
nand2 gate495( .a(G1252), .b(G1253), .O(G1304) );
nand2 gate496( .a(G1254), .b(G1255), .O(G1305) );
nand2 gate497( .a(G1256), .b(G1257), .O(G1306) );
nand2 gate498( .a(G1258), .b(G1259), .O(G1307) );
nand2 gate499( .a(G1260), .b(G1261), .O(G1308) );

  xor2  gate1891(.a(G1263), .b(G1262), .O(gate500inter0));
  nand2 gate1892(.a(gate500inter0), .b(s_192), .O(gate500inter1));
  and2  gate1893(.a(G1263), .b(G1262), .O(gate500inter2));
  inv1  gate1894(.a(s_192), .O(gate500inter3));
  inv1  gate1895(.a(s_193), .O(gate500inter4));
  nand2 gate1896(.a(gate500inter4), .b(gate500inter3), .O(gate500inter5));
  nor2  gate1897(.a(gate500inter5), .b(gate500inter2), .O(gate500inter6));
  inv1  gate1898(.a(G1262), .O(gate500inter7));
  inv1  gate1899(.a(G1263), .O(gate500inter8));
  nand2 gate1900(.a(gate500inter8), .b(gate500inter7), .O(gate500inter9));
  nand2 gate1901(.a(s_193), .b(gate500inter3), .O(gate500inter10));
  nor2  gate1902(.a(gate500inter10), .b(gate500inter9), .O(gate500inter11));
  nor2  gate1903(.a(gate500inter11), .b(gate500inter6), .O(gate500inter12));
  nand2 gate1904(.a(gate500inter12), .b(gate500inter1), .O(G1309));
nand2 gate501( .a(G1264), .b(G1265), .O(G1310) );
nand2 gate502( .a(G1266), .b(G1267), .O(G1311) );
nand2 gate503( .a(G1268), .b(G1269), .O(G1312) );
nand2 gate504( .a(G1270), .b(G1271), .O(G1313) );
nand2 gate505( .a(G1272), .b(G1273), .O(G1314) );
nand2 gate506( .a(G1274), .b(G1275), .O(G1315) );

  xor2  gate1989(.a(G1277), .b(G1276), .O(gate507inter0));
  nand2 gate1990(.a(gate507inter0), .b(s_206), .O(gate507inter1));
  and2  gate1991(.a(G1277), .b(G1276), .O(gate507inter2));
  inv1  gate1992(.a(s_206), .O(gate507inter3));
  inv1  gate1993(.a(s_207), .O(gate507inter4));
  nand2 gate1994(.a(gate507inter4), .b(gate507inter3), .O(gate507inter5));
  nor2  gate1995(.a(gate507inter5), .b(gate507inter2), .O(gate507inter6));
  inv1  gate1996(.a(G1276), .O(gate507inter7));
  inv1  gate1997(.a(G1277), .O(gate507inter8));
  nand2 gate1998(.a(gate507inter8), .b(gate507inter7), .O(gate507inter9));
  nand2 gate1999(.a(s_207), .b(gate507inter3), .O(gate507inter10));
  nor2  gate2000(.a(gate507inter10), .b(gate507inter9), .O(gate507inter11));
  nor2  gate2001(.a(gate507inter11), .b(gate507inter6), .O(gate507inter12));
  nand2 gate2002(.a(gate507inter12), .b(gate507inter1), .O(G1316));
nand2 gate508( .a(G1278), .b(G1279), .O(G1317) );
nand2 gate509( .a(G1280), .b(G1281), .O(G1318) );
nand2 gate510( .a(G1282), .b(G1283), .O(G1319) );

  xor2  gate1205(.a(G1285), .b(G1284), .O(gate511inter0));
  nand2 gate1206(.a(gate511inter0), .b(s_94), .O(gate511inter1));
  and2  gate1207(.a(G1285), .b(G1284), .O(gate511inter2));
  inv1  gate1208(.a(s_94), .O(gate511inter3));
  inv1  gate1209(.a(s_95), .O(gate511inter4));
  nand2 gate1210(.a(gate511inter4), .b(gate511inter3), .O(gate511inter5));
  nor2  gate1211(.a(gate511inter5), .b(gate511inter2), .O(gate511inter6));
  inv1  gate1212(.a(G1284), .O(gate511inter7));
  inv1  gate1213(.a(G1285), .O(gate511inter8));
  nand2 gate1214(.a(gate511inter8), .b(gate511inter7), .O(gate511inter9));
  nand2 gate1215(.a(s_95), .b(gate511inter3), .O(gate511inter10));
  nor2  gate1216(.a(gate511inter10), .b(gate511inter9), .O(gate511inter11));
  nor2  gate1217(.a(gate511inter11), .b(gate511inter6), .O(gate511inter12));
  nand2 gate1218(.a(gate511inter12), .b(gate511inter1), .O(G1320));

  xor2  gate1919(.a(G1287), .b(G1286), .O(gate512inter0));
  nand2 gate1920(.a(gate512inter0), .b(s_196), .O(gate512inter1));
  and2  gate1921(.a(G1287), .b(G1286), .O(gate512inter2));
  inv1  gate1922(.a(s_196), .O(gate512inter3));
  inv1  gate1923(.a(s_197), .O(gate512inter4));
  nand2 gate1924(.a(gate512inter4), .b(gate512inter3), .O(gate512inter5));
  nor2  gate1925(.a(gate512inter5), .b(gate512inter2), .O(gate512inter6));
  inv1  gate1926(.a(G1286), .O(gate512inter7));
  inv1  gate1927(.a(G1287), .O(gate512inter8));
  nand2 gate1928(.a(gate512inter8), .b(gate512inter7), .O(gate512inter9));
  nand2 gate1929(.a(s_197), .b(gate512inter3), .O(gate512inter10));
  nor2  gate1930(.a(gate512inter10), .b(gate512inter9), .O(gate512inter11));
  nor2  gate1931(.a(gate512inter11), .b(gate512inter6), .O(gate512inter12));
  nand2 gate1932(.a(gate512inter12), .b(gate512inter1), .O(G1321));

  xor2  gate1093(.a(G1289), .b(G1288), .O(gate513inter0));
  nand2 gate1094(.a(gate513inter0), .b(s_78), .O(gate513inter1));
  and2  gate1095(.a(G1289), .b(G1288), .O(gate513inter2));
  inv1  gate1096(.a(s_78), .O(gate513inter3));
  inv1  gate1097(.a(s_79), .O(gate513inter4));
  nand2 gate1098(.a(gate513inter4), .b(gate513inter3), .O(gate513inter5));
  nor2  gate1099(.a(gate513inter5), .b(gate513inter2), .O(gate513inter6));
  inv1  gate1100(.a(G1288), .O(gate513inter7));
  inv1  gate1101(.a(G1289), .O(gate513inter8));
  nand2 gate1102(.a(gate513inter8), .b(gate513inter7), .O(gate513inter9));
  nand2 gate1103(.a(s_79), .b(gate513inter3), .O(gate513inter10));
  nor2  gate1104(.a(gate513inter10), .b(gate513inter9), .O(gate513inter11));
  nor2  gate1105(.a(gate513inter11), .b(gate513inter6), .O(gate513inter12));
  nand2 gate1106(.a(gate513inter12), .b(gate513inter1), .O(G1322));

  xor2  gate1569(.a(G1291), .b(G1290), .O(gate514inter0));
  nand2 gate1570(.a(gate514inter0), .b(s_146), .O(gate514inter1));
  and2  gate1571(.a(G1291), .b(G1290), .O(gate514inter2));
  inv1  gate1572(.a(s_146), .O(gate514inter3));
  inv1  gate1573(.a(s_147), .O(gate514inter4));
  nand2 gate1574(.a(gate514inter4), .b(gate514inter3), .O(gate514inter5));
  nor2  gate1575(.a(gate514inter5), .b(gate514inter2), .O(gate514inter6));
  inv1  gate1576(.a(G1290), .O(gate514inter7));
  inv1  gate1577(.a(G1291), .O(gate514inter8));
  nand2 gate1578(.a(gate514inter8), .b(gate514inter7), .O(gate514inter9));
  nand2 gate1579(.a(s_147), .b(gate514inter3), .O(gate514inter10));
  nor2  gate1580(.a(gate514inter10), .b(gate514inter9), .O(gate514inter11));
  nor2  gate1581(.a(gate514inter11), .b(gate514inter6), .O(gate514inter12));
  nand2 gate1582(.a(gate514inter12), .b(gate514inter1), .O(G1323));
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule