module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);

input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;//RE__PI;

input s_0,s_1;//RE__ALLOW(00,01,10,11);
input s_2,s_3;//RE__ALLOW(00,01,10,11);
input s_4,s_5;//RE__ALLOW(00,01,10,11);
input s_6,s_7;//RE__ALLOW(00,01,10,11);
input s_8,s_9;//RE__ALLOW(00,01,10,11);
input s_10,s_11;//RE__ALLOW(00,01,10,11);
input s_12,s_13;//RE__ALLOW(00,01,10,11);
input s_14,s_15;//RE__ALLOW(00,01,10,11);
input s_16,s_17;//RE__ALLOW(00,01,10,11);
input s_18,s_19;//RE__ALLOW(00,01,10,11);
input s_20,s_21;//RE__ALLOW(00,01,10,11);
input s_22,s_23;//RE__ALLOW(00,01,10,11);
input s_24,s_25;//RE__ALLOW(00,01,10,11);
input s_26,s_27;//RE__ALLOW(00,01,10,11);
input s_28,s_29;//RE__ALLOW(00,01,10,11);
input s_30,s_31;//RE__ALLOW(00,01,10,11);
input s_32,s_33;//RE__ALLOW(00,01,10,11);
input s_34,s_35;//RE__ALLOW(00,01,10,11);
input s_36,s_37;//RE__ALLOW(00,01,10,11);
input s_38,s_39;//RE__ALLOW(00,01,10,11);
input s_40,s_41;//RE__ALLOW(00,01,10,11);
input s_42,s_43;//RE__ALLOW(00,01,10,11);
input s_44,s_45;//RE__ALLOW(00,01,10,11);
input s_46,s_47;//RE__ALLOW(00,01,10,11);
input s_48,s_49;//RE__ALLOW(00,01,10,11);
input s_50,s_51;//RE__ALLOW(00,01,10,11);
input s_52,s_53;//RE__ALLOW(00,01,10,11);
input s_54,s_55;//RE__ALLOW(00,01,10,11);
input s_56,s_57;//RE__ALLOW(00,01,10,11);
input s_58,s_59;//RE__ALLOW(00,01,10,11);
input s_60,s_61;//RE__ALLOW(00,01,10,11);
input s_62,s_63;//RE__ALLOW(00,01,10,11);
input s_64,s_65;//RE__ALLOW(00,01,10,11);
input s_66,s_67;//RE__ALLOW(00,01,10,11);
input s_68,s_69;//RE__ALLOW(00,01,10,11);
input s_70,s_71;//RE__ALLOW(00,01,10,11);
input s_72,s_73;//RE__ALLOW(00,01,10,11);
input s_74,s_75;//RE__ALLOW(00,01,10,11);
input s_76,s_77;//RE__ALLOW(00,01,10,11);
input s_78,s_79;//RE__ALLOW(00,01,10,11);
input s_80,s_81;//RE__ALLOW(00,01,10,11);
input s_82,s_83;//RE__ALLOW(00,01,10,11);
input s_84,s_85;//RE__ALLOW(00,01,10,11);
input s_86,s_87;//RE__ALLOW(00,01,10,11);
input s_88,s_89;//RE__ALLOW(00,01,10,11);
input s_90,s_91;//RE__ALLOW(00,01,10,11);
input s_92,s_93;//RE__ALLOW(00,01,10,11);
input s_94,s_95;//RE__ALLOW(00,01,10,11);
input s_96,s_97;//RE__ALLOW(00,01,10,11);
input s_98,s_99;//RE__ALLOW(00,01,10,11);
input s_100,s_101;//RE__ALLOW(00,01,10,11);
input s_102,s_103;//RE__ALLOW(00,01,10,11);
input s_104,s_105;//RE__ALLOW(00,01,10,11);
input s_106,s_107;//RE__ALLOW(00,01,10,11);
input s_108,s_109;//RE__ALLOW(00,01,10,11);
input s_110,s_111;//RE__ALLOW(00,01,10,11);
input s_112,s_113;//RE__ALLOW(00,01,10,11);
input s_114,s_115;//RE__ALLOW(00,01,10,11);
input s_116,s_117;//RE__ALLOW(00,01,10,11);
input s_118,s_119;//RE__ALLOW(00,01,10,11);
input s_120,s_121;//RE__ALLOW(00,01,10,11);
input s_122,s_123;//RE__ALLOW(00,01,10,11);
input s_124,s_125;//RE__ALLOW(00,01,10,11);
input s_126,s_127;//RE__ALLOW(00,01,10,11);
input s_128,s_129;//RE__ALLOW(00,01,10,11);
input s_130,s_131;//RE__ALLOW(00,01,10,11);
input s_132,s_133;//RE__ALLOW(00,01,10,11);
input s_134,s_135;//RE__ALLOW(00,01,10,11);
input s_136,s_137;//RE__ALLOW(00,01,10,11);
input s_138,s_139;//RE__ALLOW(00,01,10,11);
input s_140,s_141;//RE__ALLOW(00,01,10,11);
input s_142,s_143;//RE__ALLOW(00,01,10,11);
input s_144,s_145;//RE__ALLOW(00,01,10,11);
input s_146,s_147;//RE__ALLOW(00,01,10,11);
input s_148,s_149;//RE__ALLOW(00,01,10,11);
input s_150,s_151;//RE__ALLOW(00,01,10,11);
input s_152,s_153;//RE__ALLOW(00,01,10,11);
input s_154,s_155;//RE__ALLOW(00,01,10,11);
input s_156,s_157;//RE__ALLOW(00,01,10,11);
input s_158,s_159;//RE__ALLOW(00,01,10,11);
input s_160,s_161;//RE__ALLOW(00,01,10,11);
input s_162,s_163;//RE__ALLOW(00,01,10,11);
input s_164,s_165;//RE__ALLOW(00,01,10,11);
input s_166,s_167;//RE__ALLOW(00,01,10,11);
input s_168,s_169;//RE__ALLOW(00,01,10,11);
input s_170,s_171;//RE__ALLOW(00,01,10,11);
input s_172,s_173;//RE__ALLOW(00,01,10,11);
input s_174,s_175;//RE__ALLOW(00,01,10,11);
input s_176,s_177;//RE__ALLOW(00,01,10,11);
input s_178,s_179;//RE__ALLOW(00,01,10,11);
input s_180,s_181;//RE__ALLOW(00,01,10,11);
input s_182,s_183;//RE__ALLOW(00,01,10,11);
input s_184,s_185;//RE__ALLOW(00,01,10,11);
input s_186,s_187;//RE__ALLOW(00,01,10,11);
input s_188,s_189;//RE__ALLOW(00,01,10,11);
input s_190,s_191;//RE__ALLOW(00,01,10,11);
input s_192,s_193;//RE__ALLOW(00,01,10,11);
input s_194,s_195;//RE__ALLOW(00,01,10,11);
input s_196,s_197;//RE__ALLOW(00,01,10,11);
input s_198,s_199;//RE__ALLOW(00,01,10,11);
input s_200,s_201;//RE__ALLOW(00,01,10,11);
input s_202,s_203;//RE__ALLOW(00,01,10,11);
input s_204,s_205;//RE__ALLOW(00,01,10,11);
input s_206,s_207;//RE__ALLOW(00,01,10,11);
input s_208,s_209;//RE__ALLOW(00,01,10,11);
input s_210,s_211;//RE__ALLOW(00,01,10,11);
input s_212,s_213;//RE__ALLOW(00,01,10,11);
input s_214,s_215;//RE__ALLOW(00,01,10,11);
input s_216,s_217;//RE__ALLOW(00,01,10,11);
input s_218,s_219;//RE__ALLOW(00,01,10,11);
input s_220,s_221;//RE__ALLOW(00,01,10,11);
input s_222,s_223;//RE__ALLOW(00,01,10,11);
input s_224,s_225;//RE__ALLOW(00,01,10,11);
input s_226,s_227;//RE__ALLOW(00,01,10,11);
input s_228,s_229;//RE__ALLOW(00,01,10,11);
input s_230,s_231;//RE__ALLOW(00,01,10,11);
input s_232,s_233;//RE__ALLOW(00,01,10,11);
input s_234,s_235;//RE__ALLOW(00,01,10,11);
input s_236,s_237;//RE__ALLOW(00,01,10,11);
input s_238,s_239;//RE__ALLOW(00,01,10,11);
input s_240,s_241;//RE__ALLOW(00,01,10,11);
input s_242,s_243;//RE__ALLOW(00,01,10,11);
input s_244,s_245;//RE__ALLOW(00,01,10,11);
input s_246,s_247;//RE__ALLOW(00,01,10,11);
input s_248,s_249;//RE__ALLOW(00,01,10,11);
input s_250,s_251;//RE__ALLOW(00,01,10,11);
input s_252,s_253;//RE__ALLOW(00,01,10,11);
input s_254,s_255;//RE__ALLOW(00,01,10,11);
input s_256,s_257;//RE__ALLOW(00,01,10,11);
input s_258,s_259;//RE__ALLOW(00,01,10,11);
input s_260,s_261;//RE__ALLOW(00,01,10,11);
input s_262,s_263;//RE__ALLOW(00,01,10,11);
input s_264,s_265;//RE__ALLOW(00,01,10,11);
input s_266,s_267;//RE__ALLOW(00,01,10,11);
input s_268,s_269;//RE__ALLOW(00,01,10,11);
input s_270,s_271;//RE__ALLOW(00,01,10,11);
input s_272,s_273;//RE__ALLOW(00,01,10,11);
input s_274,s_275;//RE__ALLOW(00,01,10,11);
input s_276,s_277;//RE__ALLOW(00,01,10,11);
input s_278,s_279;//RE__ALLOW(00,01,10,11);
input s_280,s_281;//RE__ALLOW(00,01,10,11);
input s_282,s_283;//RE__ALLOW(00,01,10,11);
input s_284,s_285;//RE__ALLOW(00,01,10,11);
input s_286,s_287;//RE__ALLOW(00,01,10,11);
input s_288,s_289;//RE__ALLOW(00,01,10,11);
input s_290,s_291;//RE__ALLOW(00,01,10,11);
input s_292,s_293;//RE__ALLOW(00,01,10,11);
input s_294,s_295;//RE__ALLOW(00,01,10,11);
input s_296,s_297;//RE__ALLOW(00,01,10,11);
input s_298,s_299;//RE__ALLOW(00,01,10,11);
input s_300,s_301;//RE__ALLOW(00,01,10,11);
input s_302,s_303;//RE__ALLOW(00,01,10,11);
input s_304,s_305;//RE__ALLOW(00,01,10,11);
input s_306,s_307;//RE__ALLOW(00,01,10,11);
input s_308,s_309;//RE__ALLOW(00,01,10,11);
input s_310,s_311;//RE__ALLOW(00,01,10,11);
input s_312,s_313;//RE__ALLOW(00,01,10,11);
input s_314,s_315;//RE__ALLOW(00,01,10,11);
input s_316,s_317;//RE__ALLOW(00,01,10,11);
input s_318,s_319;//RE__ALLOW(00,01,10,11);
input s_320,s_321;//RE__ALLOW(00,01,10,11);
input s_322,s_323;//RE__ALLOW(00,01,10,11);
input s_324,s_325;//RE__ALLOW(00,01,10,11);
input s_326,s_327;//RE__ALLOW(00,01,10,11);
input s_328,s_329;//RE__ALLOW(00,01,10,11);
input s_330,s_331;//RE__ALLOW(00,01,10,11);
input s_332,s_333;//RE__ALLOW(00,01,10,11);
input s_334,s_335;//RE__ALLOW(00,01,10,11);
input s_336,s_337;//RE__ALLOW(00,01,10,11);
input s_338,s_339;//RE__ALLOW(00,01,10,11);
input s_340,s_341;//RE__ALLOW(00,01,10,11);
input s_342,s_343;//RE__ALLOW(00,01,10,11);
input s_344,s_345;//RE__ALLOW(00,01,10,11);
input s_346,s_347;//RE__ALLOW(00,01,10,11);
input s_348,s_349;//RE__ALLOW(00,01,10,11);
input s_350,s_351;//RE__ALLOW(00,01,10,11);
input s_352,s_353;//RE__ALLOW(00,01,10,11);
input s_354,s_355;//RE__ALLOW(00,01,10,11);
input s_356,s_357;//RE__ALLOW(00,01,10,11);
input s_358,s_359;//RE__ALLOW(00,01,10,11);
input s_360,s_361;//RE__ALLOW(00,01,10,11);
input s_362,s_363;//RE__ALLOW(00,01,10,11);
input s_364,s_365;//RE__ALLOW(00,01,10,11);
input s_366,s_367;//RE__ALLOW(00,01,10,11);
input s_368,s_369;//RE__ALLOW(00,01,10,11);
input s_370,s_371;//RE__ALLOW(00,01,10,11);
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;

  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate42inter0, gate42inter1, gate42inter2, gate42inter3, gate42inter4, gate42inter5, gate42inter6, gate42inter7, gate42inter8, gate42inter9, gate42inter10, gate42inter11, gate42inter12, gate63inter0, gate63inter1, gate63inter2, gate63inter3, gate63inter4, gate63inter5, gate63inter6, gate63inter7, gate63inter8, gate63inter9, gate63inter10, gate63inter11, gate63inter12, gate431inter0, gate431inter1, gate431inter2, gate431inter3, gate431inter4, gate431inter5, gate431inter6, gate431inter7, gate431inter8, gate431inter9, gate431inter10, gate431inter11, gate431inter12, gate82inter0, gate82inter1, gate82inter2, gate82inter3, gate82inter4, gate82inter5, gate82inter6, gate82inter7, gate82inter8, gate82inter9, gate82inter10, gate82inter11, gate82inter12, gate496inter0, gate496inter1, gate496inter2, gate496inter3, gate496inter4, gate496inter5, gate496inter6, gate496inter7, gate496inter8, gate496inter9, gate496inter10, gate496inter11, gate496inter12, gate232inter0, gate232inter1, gate232inter2, gate232inter3, gate232inter4, gate232inter5, gate232inter6, gate232inter7, gate232inter8, gate232inter9, gate232inter10, gate232inter11, gate232inter12, gate123inter0, gate123inter1, gate123inter2, gate123inter3, gate123inter4, gate123inter5, gate123inter6, gate123inter7, gate123inter8, gate123inter9, gate123inter10, gate123inter11, gate123inter12, gate421inter0, gate421inter1, gate421inter2, gate421inter3, gate421inter4, gate421inter5, gate421inter6, gate421inter7, gate421inter8, gate421inter9, gate421inter10, gate421inter11, gate421inter12, gate148inter0, gate148inter1, gate148inter2, gate148inter3, gate148inter4, gate148inter5, gate148inter6, gate148inter7, gate148inter8, gate148inter9, gate148inter10, gate148inter11, gate148inter12, gate71inter0, gate71inter1, gate71inter2, gate71inter3, gate71inter4, gate71inter5, gate71inter6, gate71inter7, gate71inter8, gate71inter9, gate71inter10, gate71inter11, gate71inter12, gate173inter0, gate173inter1, gate173inter2, gate173inter3, gate173inter4, gate173inter5, gate173inter6, gate173inter7, gate173inter8, gate173inter9, gate173inter10, gate173inter11, gate173inter12, gate198inter0, gate198inter1, gate198inter2, gate198inter3, gate198inter4, gate198inter5, gate198inter6, gate198inter7, gate198inter8, gate198inter9, gate198inter10, gate198inter11, gate198inter12, gate40inter0, gate40inter1, gate40inter2, gate40inter3, gate40inter4, gate40inter5, gate40inter6, gate40inter7, gate40inter8, gate40inter9, gate40inter10, gate40inter11, gate40inter12, gate462inter0, gate462inter1, gate462inter2, gate462inter3, gate462inter4, gate462inter5, gate462inter6, gate462inter7, gate462inter8, gate462inter9, gate462inter10, gate462inter11, gate462inter12, gate495inter0, gate495inter1, gate495inter2, gate495inter3, gate495inter4, gate495inter5, gate495inter6, gate495inter7, gate495inter8, gate495inter9, gate495inter10, gate495inter11, gate495inter12, gate60inter0, gate60inter1, gate60inter2, gate60inter3, gate60inter4, gate60inter5, gate60inter6, gate60inter7, gate60inter8, gate60inter9, gate60inter10, gate60inter11, gate60inter12, gate390inter0, gate390inter1, gate390inter2, gate390inter3, gate390inter4, gate390inter5, gate390inter6, gate390inter7, gate390inter8, gate390inter9, gate390inter10, gate390inter11, gate390inter12, gate168inter0, gate168inter1, gate168inter2, gate168inter3, gate168inter4, gate168inter5, gate168inter6, gate168inter7, gate168inter8, gate168inter9, gate168inter10, gate168inter11, gate168inter12, gate501inter0, gate501inter1, gate501inter2, gate501inter3, gate501inter4, gate501inter5, gate501inter6, gate501inter7, gate501inter8, gate501inter9, gate501inter10, gate501inter11, gate501inter12, gate25inter0, gate25inter1, gate25inter2, gate25inter3, gate25inter4, gate25inter5, gate25inter6, gate25inter7, gate25inter8, gate25inter9, gate25inter10, gate25inter11, gate25inter12, gate183inter0, gate183inter1, gate183inter2, gate183inter3, gate183inter4, gate183inter5, gate183inter6, gate183inter7, gate183inter8, gate183inter9, gate183inter10, gate183inter11, gate183inter12, gate442inter0, gate442inter1, gate442inter2, gate442inter3, gate442inter4, gate442inter5, gate442inter6, gate442inter7, gate442inter8, gate442inter9, gate442inter10, gate442inter11, gate442inter12, gate399inter0, gate399inter1, gate399inter2, gate399inter3, gate399inter4, gate399inter5, gate399inter6, gate399inter7, gate399inter8, gate399inter9, gate399inter10, gate399inter11, gate399inter12, gate37inter0, gate37inter1, gate37inter2, gate37inter3, gate37inter4, gate37inter5, gate37inter6, gate37inter7, gate37inter8, gate37inter9, gate37inter10, gate37inter11, gate37inter12, gate263inter0, gate263inter1, gate263inter2, gate263inter3, gate263inter4, gate263inter5, gate263inter6, gate263inter7, gate263inter8, gate263inter9, gate263inter10, gate263inter11, gate263inter12, gate427inter0, gate427inter1, gate427inter2, gate427inter3, gate427inter4, gate427inter5, gate427inter6, gate427inter7, gate427inter8, gate427inter9, gate427inter10, gate427inter11, gate427inter12, gate38inter0, gate38inter1, gate38inter2, gate38inter3, gate38inter4, gate38inter5, gate38inter6, gate38inter7, gate38inter8, gate38inter9, gate38inter10, gate38inter11, gate38inter12, gate67inter0, gate67inter1, gate67inter2, gate67inter3, gate67inter4, gate67inter5, gate67inter6, gate67inter7, gate67inter8, gate67inter9, gate67inter10, gate67inter11, gate67inter12, gate224inter0, gate224inter1, gate224inter2, gate224inter3, gate224inter4, gate224inter5, gate224inter6, gate224inter7, gate224inter8, gate224inter9, gate224inter10, gate224inter11, gate224inter12, gate169inter0, gate169inter1, gate169inter2, gate169inter3, gate169inter4, gate169inter5, gate169inter6, gate169inter7, gate169inter8, gate169inter9, gate169inter10, gate169inter11, gate169inter12, gate212inter0, gate212inter1, gate212inter2, gate212inter3, gate212inter4, gate212inter5, gate212inter6, gate212inter7, gate212inter8, gate212inter9, gate212inter10, gate212inter11, gate212inter12, gate61inter0, gate61inter1, gate61inter2, gate61inter3, gate61inter4, gate61inter5, gate61inter6, gate61inter7, gate61inter8, gate61inter9, gate61inter10, gate61inter11, gate61inter12, gate110inter0, gate110inter1, gate110inter2, gate110inter3, gate110inter4, gate110inter5, gate110inter6, gate110inter7, gate110inter8, gate110inter9, gate110inter10, gate110inter11, gate110inter12, gate398inter0, gate398inter1, gate398inter2, gate398inter3, gate398inter4, gate398inter5, gate398inter6, gate398inter7, gate398inter8, gate398inter9, gate398inter10, gate398inter11, gate398inter12, gate451inter0, gate451inter1, gate451inter2, gate451inter3, gate451inter4, gate451inter5, gate451inter6, gate451inter7, gate451inter8, gate451inter9, gate451inter10, gate451inter11, gate451inter12, gate121inter0, gate121inter1, gate121inter2, gate121inter3, gate121inter4, gate121inter5, gate121inter6, gate121inter7, gate121inter8, gate121inter9, gate121inter10, gate121inter11, gate121inter12, gate98inter0, gate98inter1, gate98inter2, gate98inter3, gate98inter4, gate98inter5, gate98inter6, gate98inter7, gate98inter8, gate98inter9, gate98inter10, gate98inter11, gate98inter12, gate195inter0, gate195inter1, gate195inter2, gate195inter3, gate195inter4, gate195inter5, gate195inter6, gate195inter7, gate195inter8, gate195inter9, gate195inter10, gate195inter11, gate195inter12, gate213inter0, gate213inter1, gate213inter2, gate213inter3, gate213inter4, gate213inter5, gate213inter6, gate213inter7, gate213inter8, gate213inter9, gate213inter10, gate213inter11, gate213inter12, gate471inter0, gate471inter1, gate471inter2, gate471inter3, gate471inter4, gate471inter5, gate471inter6, gate471inter7, gate471inter8, gate471inter9, gate471inter10, gate471inter11, gate471inter12, gate268inter0, gate268inter1, gate268inter2, gate268inter3, gate268inter4, gate268inter5, gate268inter6, gate268inter7, gate268inter8, gate268inter9, gate268inter10, gate268inter11, gate268inter12, gate153inter0, gate153inter1, gate153inter2, gate153inter3, gate153inter4, gate153inter5, gate153inter6, gate153inter7, gate153inter8, gate153inter9, gate153inter10, gate153inter11, gate153inter12, gate12inter0, gate12inter1, gate12inter2, gate12inter3, gate12inter4, gate12inter5, gate12inter6, gate12inter7, gate12inter8, gate12inter9, gate12inter10, gate12inter11, gate12inter12, gate190inter0, gate190inter1, gate190inter2, gate190inter3, gate190inter4, gate190inter5, gate190inter6, gate190inter7, gate190inter8, gate190inter9, gate190inter10, gate190inter11, gate190inter12, gate226inter0, gate226inter1, gate226inter2, gate226inter3, gate226inter4, gate226inter5, gate226inter6, gate226inter7, gate226inter8, gate226inter9, gate226inter10, gate226inter11, gate226inter12, gate251inter0, gate251inter1, gate251inter2, gate251inter3, gate251inter4, gate251inter5, gate251inter6, gate251inter7, gate251inter8, gate251inter9, gate251inter10, gate251inter11, gate251inter12, gate512inter0, gate512inter1, gate512inter2, gate512inter3, gate512inter4, gate512inter5, gate512inter6, gate512inter7, gate512inter8, gate512inter9, gate512inter10, gate512inter11, gate512inter12, gate191inter0, gate191inter1, gate191inter2, gate191inter3, gate191inter4, gate191inter5, gate191inter6, gate191inter7, gate191inter8, gate191inter9, gate191inter10, gate191inter11, gate191inter12, gate470inter0, gate470inter1, gate470inter2, gate470inter3, gate470inter4, gate470inter5, gate470inter6, gate470inter7, gate470inter8, gate470inter9, gate470inter10, gate470inter11, gate470inter12, gate211inter0, gate211inter1, gate211inter2, gate211inter3, gate211inter4, gate211inter5, gate211inter6, gate211inter7, gate211inter8, gate211inter9, gate211inter10, gate211inter11, gate211inter12, gate402inter0, gate402inter1, gate402inter2, gate402inter3, gate402inter4, gate402inter5, gate402inter6, gate402inter7, gate402inter8, gate402inter9, gate402inter10, gate402inter11, gate402inter12, gate138inter0, gate138inter1, gate138inter2, gate138inter3, gate138inter4, gate138inter5, gate138inter6, gate138inter7, gate138inter8, gate138inter9, gate138inter10, gate138inter11, gate138inter12, gate117inter0, gate117inter1, gate117inter2, gate117inter3, gate117inter4, gate117inter5, gate117inter6, gate117inter7, gate117inter8, gate117inter9, gate117inter10, gate117inter11, gate117inter12, gate84inter0, gate84inter1, gate84inter2, gate84inter3, gate84inter4, gate84inter5, gate84inter6, gate84inter7, gate84inter8, gate84inter9, gate84inter10, gate84inter11, gate84inter12, gate253inter0, gate253inter1, gate253inter2, gate253inter3, gate253inter4, gate253inter5, gate253inter6, gate253inter7, gate253inter8, gate253inter9, gate253inter10, gate253inter11, gate253inter12, gate237inter0, gate237inter1, gate237inter2, gate237inter3, gate237inter4, gate237inter5, gate237inter6, gate237inter7, gate237inter8, gate237inter9, gate237inter10, gate237inter11, gate237inter12, gate58inter0, gate58inter1, gate58inter2, gate58inter3, gate58inter4, gate58inter5, gate58inter6, gate58inter7, gate58inter8, gate58inter9, gate58inter10, gate58inter11, gate58inter12, gate438inter0, gate438inter1, gate438inter2, gate438inter3, gate438inter4, gate438inter5, gate438inter6, gate438inter7, gate438inter8, gate438inter9, gate438inter10, gate438inter11, gate438inter12, gate143inter0, gate143inter1, gate143inter2, gate143inter3, gate143inter4, gate143inter5, gate143inter6, gate143inter7, gate143inter8, gate143inter9, gate143inter10, gate143inter11, gate143inter12, gate228inter0, gate228inter1, gate228inter2, gate228inter3, gate228inter4, gate228inter5, gate228inter6, gate228inter7, gate228inter8, gate228inter9, gate228inter10, gate228inter11, gate228inter12, gate270inter0, gate270inter1, gate270inter2, gate270inter3, gate270inter4, gate270inter5, gate270inter6, gate270inter7, gate270inter8, gate270inter9, gate270inter10, gate270inter11, gate270inter12, gate467inter0, gate467inter1, gate467inter2, gate467inter3, gate467inter4, gate467inter5, gate467inter6, gate467inter7, gate467inter8, gate467inter9, gate467inter10, gate467inter11, gate467inter12, gate219inter0, gate219inter1, gate219inter2, gate219inter3, gate219inter4, gate219inter5, gate219inter6, gate219inter7, gate219inter8, gate219inter9, gate219inter10, gate219inter11, gate219inter12, gate85inter0, gate85inter1, gate85inter2, gate85inter3, gate85inter4, gate85inter5, gate85inter6, gate85inter7, gate85inter8, gate85inter9, gate85inter10, gate85inter11, gate85inter12, gate194inter0, gate194inter1, gate194inter2, gate194inter3, gate194inter4, gate194inter5, gate194inter6, gate194inter7, gate194inter8, gate194inter9, gate194inter10, gate194inter11, gate194inter12, gate205inter0, gate205inter1, gate205inter2, gate205inter3, gate205inter4, gate205inter5, gate205inter6, gate205inter7, gate205inter8, gate205inter9, gate205inter10, gate205inter11, gate205inter12, gate146inter0, gate146inter1, gate146inter2, gate146inter3, gate146inter4, gate146inter5, gate146inter6, gate146inter7, gate146inter8, gate146inter9, gate146inter10, gate146inter11, gate146inter12, gate408inter0, gate408inter1, gate408inter2, gate408inter3, gate408inter4, gate408inter5, gate408inter6, gate408inter7, gate408inter8, gate408inter9, gate408inter10, gate408inter11, gate408inter12, gate502inter0, gate502inter1, gate502inter2, gate502inter3, gate502inter4, gate502inter5, gate502inter6, gate502inter7, gate502inter8, gate502inter9, gate502inter10, gate502inter11, gate502inter12, gate104inter0, gate104inter1, gate104inter2, gate104inter3, gate104inter4, gate104inter5, gate104inter6, gate104inter7, gate104inter8, gate104inter9, gate104inter10, gate104inter11, gate104inter12, gate86inter0, gate86inter1, gate86inter2, gate86inter3, gate86inter4, gate86inter5, gate86inter6, gate86inter7, gate86inter8, gate86inter9, gate86inter10, gate86inter11, gate86inter12, gate83inter0, gate83inter1, gate83inter2, gate83inter3, gate83inter4, gate83inter5, gate83inter6, gate83inter7, gate83inter8, gate83inter9, gate83inter10, gate83inter11, gate83inter12, gate262inter0, gate262inter1, gate262inter2, gate262inter3, gate262inter4, gate262inter5, gate262inter6, gate262inter7, gate262inter8, gate262inter9, gate262inter10, gate262inter11, gate262inter12, gate436inter0, gate436inter1, gate436inter2, gate436inter3, gate436inter4, gate436inter5, gate436inter6, gate436inter7, gate436inter8, gate436inter9, gate436inter10, gate436inter11, gate436inter12, gate508inter0, gate508inter1, gate508inter2, gate508inter3, gate508inter4, gate508inter5, gate508inter6, gate508inter7, gate508inter8, gate508inter9, gate508inter10, gate508inter11, gate508inter12, gate53inter0, gate53inter1, gate53inter2, gate53inter3, gate53inter4, gate53inter5, gate53inter6, gate53inter7, gate53inter8, gate53inter9, gate53inter10, gate53inter11, gate53inter12, gate93inter0, gate93inter1, gate93inter2, gate93inter3, gate93inter4, gate93inter5, gate93inter6, gate93inter7, gate93inter8, gate93inter9, gate93inter10, gate93inter11, gate93inter12, gate435inter0, gate435inter1, gate435inter2, gate435inter3, gate435inter4, gate435inter5, gate435inter6, gate435inter7, gate435inter8, gate435inter9, gate435inter10, gate435inter11, gate435inter12, gate493inter0, gate493inter1, gate493inter2, gate493inter3, gate493inter4, gate493inter5, gate493inter6, gate493inter7, gate493inter8, gate493inter9, gate493inter10, gate493inter11, gate493inter12, gate434inter0, gate434inter1, gate434inter2, gate434inter3, gate434inter4, gate434inter5, gate434inter6, gate434inter7, gate434inter8, gate434inter9, gate434inter10, gate434inter11, gate434inter12, gate405inter0, gate405inter1, gate405inter2, gate405inter3, gate405inter4, gate405inter5, gate405inter6, gate405inter7, gate405inter8, gate405inter9, gate405inter10, gate405inter11, gate405inter12, gate422inter0, gate422inter1, gate422inter2, gate422inter3, gate422inter4, gate422inter5, gate422inter6, gate422inter7, gate422inter8, gate422inter9, gate422inter10, gate422inter11, gate422inter12, gate393inter0, gate393inter1, gate393inter2, gate393inter3, gate393inter4, gate393inter5, gate393inter6, gate393inter7, gate393inter8, gate393inter9, gate393inter10, gate393inter11, gate393inter12, gate466inter0, gate466inter1, gate466inter2, gate466inter3, gate466inter4, gate466inter5, gate466inter6, gate466inter7, gate466inter8, gate466inter9, gate466inter10, gate466inter11, gate466inter12, gate202inter0, gate202inter1, gate202inter2, gate202inter3, gate202inter4, gate202inter5, gate202inter6, gate202inter7, gate202inter8, gate202inter9, gate202inter10, gate202inter11, gate202inter12, gate469inter0, gate469inter1, gate469inter2, gate469inter3, gate469inter4, gate469inter5, gate469inter6, gate469inter7, gate469inter8, gate469inter9, gate469inter10, gate469inter11, gate469inter12, gate155inter0, gate155inter1, gate155inter2, gate155inter3, gate155inter4, gate155inter5, gate155inter6, gate155inter7, gate155inter8, gate155inter9, gate155inter10, gate155inter11, gate155inter12, gate214inter0, gate214inter1, gate214inter2, gate214inter3, gate214inter4, gate214inter5, gate214inter6, gate214inter7, gate214inter8, gate214inter9, gate214inter10, gate214inter11, gate214inter12, gate440inter0, gate440inter1, gate440inter2, gate440inter3, gate440inter4, gate440inter5, gate440inter6, gate440inter7, gate440inter8, gate440inter9, gate440inter10, gate440inter11, gate440inter12, gate229inter0, gate229inter1, gate229inter2, gate229inter3, gate229inter4, gate229inter5, gate229inter6, gate229inter7, gate229inter8, gate229inter9, gate229inter10, gate229inter11, gate229inter12, gate511inter0, gate511inter1, gate511inter2, gate511inter3, gate511inter4, gate511inter5, gate511inter6, gate511inter7, gate511inter8, gate511inter9, gate511inter10, gate511inter11, gate511inter12, gate166inter0, gate166inter1, gate166inter2, gate166inter3, gate166inter4, gate166inter5, gate166inter6, gate166inter7, gate166inter8, gate166inter9, gate166inter10, gate166inter11, gate166inter12, gate171inter0, gate171inter1, gate171inter2, gate171inter3, gate171inter4, gate171inter5, gate171inter6, gate171inter7, gate171inter8, gate171inter9, gate171inter10, gate171inter11, gate171inter12, gate285inter0, gate285inter1, gate285inter2, gate285inter3, gate285inter4, gate285inter5, gate285inter6, gate285inter7, gate285inter8, gate285inter9, gate285inter10, gate285inter11, gate285inter12, gate56inter0, gate56inter1, gate56inter2, gate56inter3, gate56inter4, gate56inter5, gate56inter6, gate56inter7, gate56inter8, gate56inter9, gate56inter10, gate56inter11, gate56inter12, gate417inter0, gate417inter1, gate417inter2, gate417inter3, gate417inter4, gate417inter5, gate417inter6, gate417inter7, gate417inter8, gate417inter9, gate417inter10, gate417inter11, gate417inter12, gate407inter0, gate407inter1, gate407inter2, gate407inter3, gate407inter4, gate407inter5, gate407inter6, gate407inter7, gate407inter8, gate407inter9, gate407inter10, gate407inter11, gate407inter12, gate473inter0, gate473inter1, gate473inter2, gate473inter3, gate473inter4, gate473inter5, gate473inter6, gate473inter7, gate473inter8, gate473inter9, gate473inter10, gate473inter11, gate473inter12, gate234inter0, gate234inter1, gate234inter2, gate234inter3, gate234inter4, gate234inter5, gate234inter6, gate234inter7, gate234inter8, gate234inter9, gate234inter10, gate234inter11, gate234inter12, gate208inter0, gate208inter1, gate208inter2, gate208inter3, gate208inter4, gate208inter5, gate208inter6, gate208inter7, gate208inter8, gate208inter9, gate208inter10, gate208inter11, gate208inter12, gate132inter0, gate132inter1, gate132inter2, gate132inter3, gate132inter4, gate132inter5, gate132inter6, gate132inter7, gate132inter8, gate132inter9, gate132inter10, gate132inter11, gate132inter12, gate57inter0, gate57inter1, gate57inter2, gate57inter3, gate57inter4, gate57inter5, gate57inter6, gate57inter7, gate57inter8, gate57inter9, gate57inter10, gate57inter11, gate57inter12, gate43inter0, gate43inter1, gate43inter2, gate43inter3, gate43inter4, gate43inter5, gate43inter6, gate43inter7, gate43inter8, gate43inter9, gate43inter10, gate43inter11, gate43inter12, gate281inter0, gate281inter1, gate281inter2, gate281inter3, gate281inter4, gate281inter5, gate281inter6, gate281inter7, gate281inter8, gate281inter9, gate281inter10, gate281inter11, gate281inter12, gate31inter0, gate31inter1, gate31inter2, gate31inter3, gate31inter4, gate31inter5, gate31inter6, gate31inter7, gate31inter8, gate31inter9, gate31inter10, gate31inter11, gate31inter12, gate282inter0, gate282inter1, gate282inter2, gate282inter3, gate282inter4, gate282inter5, gate282inter6, gate282inter7, gate282inter8, gate282inter9, gate282inter10, gate282inter11, gate282inter12, gate464inter0, gate464inter1, gate464inter2, gate464inter3, gate464inter4, gate464inter5, gate464inter6, gate464inter7, gate464inter8, gate464inter9, gate464inter10, gate464inter11, gate464inter12, gate114inter0, gate114inter1, gate114inter2, gate114inter3, gate114inter4, gate114inter5, gate114inter6, gate114inter7, gate114inter8, gate114inter9, gate114inter10, gate114inter11, gate114inter12, gate139inter0, gate139inter1, gate139inter2, gate139inter3, gate139inter4, gate139inter5, gate139inter6, gate139inter7, gate139inter8, gate139inter9, gate139inter10, gate139inter11, gate139inter12, gate32inter0, gate32inter1, gate32inter2, gate32inter3, gate32inter4, gate32inter5, gate32inter6, gate32inter7, gate32inter8, gate32inter9, gate32inter10, gate32inter11, gate32inter12, gate465inter0, gate465inter1, gate465inter2, gate465inter3, gate465inter4, gate465inter5, gate465inter6, gate465inter7, gate465inter8, gate465inter9, gate465inter10, gate465inter11, gate465inter12, gate147inter0, gate147inter1, gate147inter2, gate147inter3, gate147inter4, gate147inter5, gate147inter6, gate147inter7, gate147inter8, gate147inter9, gate147inter10, gate147inter11, gate147inter12, gate106inter0, gate106inter1, gate106inter2, gate106inter3, gate106inter4, gate106inter5, gate106inter6, gate106inter7, gate106inter8, gate106inter9, gate106inter10, gate106inter11, gate106inter12, gate478inter0, gate478inter1, gate478inter2, gate478inter3, gate478inter4, gate478inter5, gate478inter6, gate478inter7, gate478inter8, gate478inter9, gate478inter10, gate478inter11, gate478inter12, gate432inter0, gate432inter1, gate432inter2, gate432inter3, gate432inter4, gate432inter5, gate432inter6, gate432inter7, gate432inter8, gate432inter9, gate432inter10, gate432inter11, gate432inter12, gate418inter0, gate418inter1, gate418inter2, gate418inter3, gate418inter4, gate418inter5, gate418inter6, gate418inter7, gate418inter8, gate418inter9, gate418inter10, gate418inter11, gate418inter12, gate136inter0, gate136inter1, gate136inter2, gate136inter3, gate136inter4, gate136inter5, gate136inter6, gate136inter7, gate136inter8, gate136inter9, gate136inter10, gate136inter11, gate136inter12, gate188inter0, gate188inter1, gate188inter2, gate188inter3, gate188inter4, gate188inter5, gate188inter6, gate188inter7, gate188inter8, gate188inter9, gate188inter10, gate188inter11, gate188inter12, gate280inter0, gate280inter1, gate280inter2, gate280inter3, gate280inter4, gate280inter5, gate280inter6, gate280inter7, gate280inter8, gate280inter9, gate280inter10, gate280inter11, gate280inter12, gate33inter0, gate33inter1, gate33inter2, gate33inter3, gate33inter4, gate33inter5, gate33inter6, gate33inter7, gate33inter8, gate33inter9, gate33inter10, gate33inter11, gate33inter12, gate187inter0, gate187inter1, gate187inter2, gate187inter3, gate187inter4, gate187inter5, gate187inter6, gate187inter7, gate187inter8, gate187inter9, gate187inter10, gate187inter11, gate187inter12, gate403inter0, gate403inter1, gate403inter2, gate403inter3, gate403inter4, gate403inter5, gate403inter6, gate403inter7, gate403inter8, gate403inter9, gate403inter10, gate403inter11, gate403inter12, gate509inter0, gate509inter1, gate509inter2, gate509inter3, gate509inter4, gate509inter5, gate509inter6, gate509inter7, gate509inter8, gate509inter9, gate509inter10, gate509inter11, gate509inter12, gate91inter0, gate91inter1, gate91inter2, gate91inter3, gate91inter4, gate91inter5, gate91inter6, gate91inter7, gate91inter8, gate91inter9, gate91inter10, gate91inter11, gate91inter12, gate154inter0, gate154inter1, gate154inter2, gate154inter3, gate154inter4, gate154inter5, gate154inter6, gate154inter7, gate154inter8, gate154inter9, gate154inter10, gate154inter11, gate154inter12, gate102inter0, gate102inter1, gate102inter2, gate102inter3, gate102inter4, gate102inter5, gate102inter6, gate102inter7, gate102inter8, gate102inter9, gate102inter10, gate102inter11, gate102inter12, gate170inter0, gate170inter1, gate170inter2, gate170inter3, gate170inter4, gate170inter5, gate170inter6, gate170inter7, gate170inter8, gate170inter9, gate170inter10, gate170inter11, gate170inter12, gate201inter0, gate201inter1, gate201inter2, gate201inter3, gate201inter4, gate201inter5, gate201inter6, gate201inter7, gate201inter8, gate201inter9, gate201inter10, gate201inter11, gate201inter12, gate233inter0, gate233inter1, gate233inter2, gate233inter3, gate233inter4, gate233inter5, gate233inter6, gate233inter7, gate233inter8, gate233inter9, gate233inter10, gate233inter11, gate233inter12, gate97inter0, gate97inter1, gate97inter2, gate97inter3, gate97inter4, gate97inter5, gate97inter6, gate97inter7, gate97inter8, gate97inter9, gate97inter10, gate97inter11, gate97inter12, gate193inter0, gate193inter1, gate193inter2, gate193inter3, gate193inter4, gate193inter5, gate193inter6, gate193inter7, gate193inter8, gate193inter9, gate193inter10, gate193inter11, gate193inter12, gate130inter0, gate130inter1, gate130inter2, gate130inter3, gate130inter4, gate130inter5, gate130inter6, gate130inter7, gate130inter8, gate130inter9, gate130inter10, gate130inter11, gate130inter12, gate283inter0, gate283inter1, gate283inter2, gate283inter3, gate283inter4, gate283inter5, gate283inter6, gate283inter7, gate283inter8, gate283inter9, gate283inter10, gate283inter11, gate283inter12, gate209inter0, gate209inter1, gate209inter2, gate209inter3, gate209inter4, gate209inter5, gate209inter6, gate209inter7, gate209inter8, gate209inter9, gate209inter10, gate209inter11, gate209inter12, gate9inter0, gate9inter1, gate9inter2, gate9inter3, gate9inter4, gate9inter5, gate9inter6, gate9inter7, gate9inter8, gate9inter9, gate9inter10, gate9inter11, gate9inter12, gate265inter0, gate265inter1, gate265inter2, gate265inter3, gate265inter4, gate265inter5, gate265inter6, gate265inter7, gate265inter8, gate265inter9, gate265inter10, gate265inter11, gate265inter12, gate161inter0, gate161inter1, gate161inter2, gate161inter3, gate161inter4, gate161inter5, gate161inter6, gate161inter7, gate161inter8, gate161inter9, gate161inter10, gate161inter11, gate161inter12, gate150inter0, gate150inter1, gate150inter2, gate150inter3, gate150inter4, gate150inter5, gate150inter6, gate150inter7, gate150inter8, gate150inter9, gate150inter10, gate150inter11, gate150inter12, gate45inter0, gate45inter1, gate45inter2, gate45inter3, gate45inter4, gate45inter5, gate45inter6, gate45inter7, gate45inter8, gate45inter9, gate45inter10, gate45inter11, gate45inter12, gate291inter0, gate291inter1, gate291inter2, gate291inter3, gate291inter4, gate291inter5, gate291inter6, gate291inter7, gate291inter8, gate291inter9, gate291inter10, gate291inter11, gate291inter12, gate425inter0, gate425inter1, gate425inter2, gate425inter3, gate425inter4, gate425inter5, gate425inter6, gate425inter7, gate425inter8, gate425inter9, gate425inter10, gate425inter11, gate425inter12, gate95inter0, gate95inter1, gate95inter2, gate95inter3, gate95inter4, gate95inter5, gate95inter6, gate95inter7, gate95inter8, gate95inter9, gate95inter10, gate95inter11, gate95inter12, gate199inter0, gate199inter1, gate199inter2, gate199inter3, gate199inter4, gate199inter5, gate199inter6, gate199inter7, gate199inter8, gate199inter9, gate199inter10, gate199inter11, gate199inter12, gate475inter0, gate475inter1, gate475inter2, gate475inter3, gate475inter4, gate475inter5, gate475inter6, gate475inter7, gate475inter8, gate475inter9, gate475inter10, gate475inter11, gate475inter12, gate222inter0, gate222inter1, gate222inter2, gate222inter3, gate222inter4, gate222inter5, gate222inter6, gate222inter7, gate222inter8, gate222inter9, gate222inter10, gate222inter11, gate222inter12, gate141inter0, gate141inter1, gate141inter2, gate141inter3, gate141inter4, gate141inter5, gate141inter6, gate141inter7, gate141inter8, gate141inter9, gate141inter10, gate141inter11, gate141inter12, gate133inter0, gate133inter1, gate133inter2, gate133inter3, gate133inter4, gate133inter5, gate133inter6, gate133inter7, gate133inter8, gate133inter9, gate133inter10, gate133inter11, gate133inter12, gate266inter0, gate266inter1, gate266inter2, gate266inter3, gate266inter4, gate266inter5, gate266inter6, gate266inter7, gate266inter8, gate266inter9, gate266inter10, gate266inter11, gate266inter12, gate157inter0, gate157inter1, gate157inter2, gate157inter3, gate157inter4, gate157inter5, gate157inter6, gate157inter7, gate157inter8, gate157inter9, gate157inter10, gate157inter11, gate157inter12, gate483inter0, gate483inter1, gate483inter2, gate483inter3, gate483inter4, gate483inter5, gate483inter6, gate483inter7, gate483inter8, gate483inter9, gate483inter10, gate483inter11, gate483inter12, gate499inter0, gate499inter1, gate499inter2, gate499inter3, gate499inter4, gate499inter5, gate499inter6, gate499inter7, gate499inter8, gate499inter9, gate499inter10, gate499inter11, gate499inter12, gate78inter0, gate78inter1, gate78inter2, gate78inter3, gate78inter4, gate78inter5, gate78inter6, gate78inter7, gate78inter8, gate78inter9, gate78inter10, gate78inter11, gate78inter12, gate39inter0, gate39inter1, gate39inter2, gate39inter3, gate39inter4, gate39inter5, gate39inter6, gate39inter7, gate39inter8, gate39inter9, gate39inter10, gate39inter11, gate39inter12, gate127inter0, gate127inter1, gate127inter2, gate127inter3, gate127inter4, gate127inter5, gate127inter6, gate127inter7, gate127inter8, gate127inter9, gate127inter10, gate127inter11, gate127inter12, gate491inter0, gate491inter1, gate491inter2, gate491inter3, gate491inter4, gate491inter5, gate491inter6, gate491inter7, gate491inter8, gate491inter9, gate491inter10, gate491inter11, gate491inter12, gate250inter0, gate250inter1, gate250inter2, gate250inter3, gate250inter4, gate250inter5, gate250inter6, gate250inter7, gate250inter8, gate250inter9, gate250inter10, gate250inter11, gate250inter12, gate387inter0, gate387inter1, gate387inter2, gate387inter3, gate387inter4, gate387inter5, gate387inter6, gate387inter7, gate387inter8, gate387inter9, gate387inter10, gate387inter11, gate387inter12, gate29inter0, gate29inter1, gate29inter2, gate29inter3, gate29inter4, gate29inter5, gate29inter6, gate29inter7, gate29inter8, gate29inter9, gate29inter10, gate29inter11, gate29inter12, gate419inter0, gate419inter1, gate419inter2, gate419inter3, gate419inter4, gate419inter5, gate419inter6, gate419inter7, gate419inter8, gate419inter9, gate419inter10, gate419inter11, gate419inter12, gate474inter0, gate474inter1, gate474inter2, gate474inter3, gate474inter4, gate474inter5, gate474inter6, gate474inter7, gate474inter8, gate474inter9, gate474inter10, gate474inter11, gate474inter12, gate30inter0, gate30inter1, gate30inter2, gate30inter3, gate30inter4, gate30inter5, gate30inter6, gate30inter7, gate30inter8, gate30inter9, gate30inter10, gate30inter11, gate30inter12, gate55inter0, gate55inter1, gate55inter2, gate55inter3, gate55inter4, gate55inter5, gate55inter6, gate55inter7, gate55inter8, gate55inter9, gate55inter10, gate55inter11, gate55inter12, gate489inter0, gate489inter1, gate489inter2, gate489inter3, gate489inter4, gate489inter5, gate489inter6, gate489inter7, gate489inter8, gate489inter9, gate489inter10, gate489inter11, gate489inter12, gate433inter0, gate433inter1, gate433inter2, gate433inter3, gate433inter4, gate433inter5, gate433inter6, gate433inter7, gate433inter8, gate433inter9, gate433inter10, gate433inter11, gate433inter12, gate248inter0, gate248inter1, gate248inter2, gate248inter3, gate248inter4, gate248inter5, gate248inter6, gate248inter7, gate248inter8, gate248inter9, gate248inter10, gate248inter11, gate248inter12, gate238inter0, gate238inter1, gate238inter2, gate238inter3, gate238inter4, gate238inter5, gate238inter6, gate238inter7, gate238inter8, gate238inter9, gate238inter10, gate238inter11, gate238inter12, gate51inter0, gate51inter1, gate51inter2, gate51inter3, gate51inter4, gate51inter5, gate51inter6, gate51inter7, gate51inter8, gate51inter9, gate51inter10, gate51inter11, gate51inter12, gate92inter0, gate92inter1, gate92inter2, gate92inter3, gate92inter4, gate92inter5, gate92inter6, gate92inter7, gate92inter8, gate92inter9, gate92inter10, gate92inter11, gate92inter12, gate392inter0, gate392inter1, gate392inter2, gate392inter3, gate392inter4, gate392inter5, gate392inter6, gate392inter7, gate392inter8, gate392inter9, gate392inter10, gate392inter11, gate392inter12, gate255inter0, gate255inter1, gate255inter2, gate255inter3, gate255inter4, gate255inter5, gate255inter6, gate255inter7, gate255inter8, gate255inter9, gate255inter10, gate255inter11, gate255inter12, gate461inter0, gate461inter1, gate461inter2, gate461inter3, gate461inter4, gate461inter5, gate461inter6, gate461inter7, gate461inter8, gate461inter9, gate461inter10, gate461inter11, gate461inter12, gate64inter0, gate64inter1, gate64inter2, gate64inter3, gate64inter4, gate64inter5, gate64inter6, gate64inter7, gate64inter8, gate64inter9, gate64inter10, gate64inter11, gate64inter12, gate413inter0, gate413inter1, gate413inter2, gate413inter3, gate413inter4, gate413inter5, gate413inter6, gate413inter7, gate413inter8, gate413inter9, gate413inter10, gate413inter11, gate413inter12, gate49inter0, gate49inter1, gate49inter2, gate49inter3, gate49inter4, gate49inter5, gate49inter6, gate49inter7, gate49inter8, gate49inter9, gate49inter10, gate49inter11, gate49inter12, gate244inter0, gate244inter1, gate244inter2, gate244inter3, gate244inter4, gate244inter5, gate244inter6, gate244inter7, gate244inter8, gate244inter9, gate244inter10, gate244inter11, gate244inter12, gate295inter0, gate295inter1, gate295inter2, gate295inter3, gate295inter4, gate295inter5, gate295inter6, gate295inter7, gate295inter8, gate295inter9, gate295inter10, gate295inter11, gate295inter12, gate100inter0, gate100inter1, gate100inter2, gate100inter3, gate100inter4, gate100inter5, gate100inter6, gate100inter7, gate100inter8, gate100inter9, gate100inter10, gate100inter11, gate100inter12, gate10inter0, gate10inter1, gate10inter2, gate10inter3, gate10inter4, gate10inter5, gate10inter6, gate10inter7, gate10inter8, gate10inter9, gate10inter10, gate10inter11, gate10inter12, gate134inter0, gate134inter1, gate134inter2, gate134inter3, gate134inter4, gate134inter5, gate134inter6, gate134inter7, gate134inter8, gate134inter9, gate134inter10, gate134inter11, gate134inter12, gate429inter0, gate429inter1, gate429inter2, gate429inter3, gate429inter4, gate429inter5, gate429inter6, gate429inter7, gate429inter8, gate429inter9, gate429inter10, gate429inter11, gate429inter12, gate388inter0, gate388inter1, gate388inter2, gate388inter3, gate388inter4, gate388inter5, gate388inter6, gate388inter7, gate388inter8, gate388inter9, gate388inter10, gate388inter11, gate388inter12, gate167inter0, gate167inter1, gate167inter2, gate167inter3, gate167inter4, gate167inter5, gate167inter6, gate167inter7, gate167inter8, gate167inter9, gate167inter10, gate167inter11, gate167inter12, gate485inter0, gate485inter1, gate485inter2, gate485inter3, gate485inter4, gate485inter5, gate485inter6, gate485inter7, gate485inter8, gate485inter9, gate485inter10, gate485inter11, gate485inter12, gate176inter0, gate176inter1, gate176inter2, gate176inter3, gate176inter4, gate176inter5, gate176inter6, gate176inter7, gate176inter8, gate176inter9, gate176inter10, gate176inter11, gate176inter12, gate290inter0, gate290inter1, gate290inter2, gate290inter3, gate290inter4, gate290inter5, gate290inter6, gate290inter7, gate290inter8, gate290inter9, gate290inter10, gate290inter11, gate290inter12, gate175inter0, gate175inter1, gate175inter2, gate175inter3, gate175inter4, gate175inter5, gate175inter6, gate175inter7, gate175inter8, gate175inter9, gate175inter10, gate175inter11, gate175inter12;



and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );

  xor2  gate2423(.a(G2), .b(G1), .O(gate9inter0));
  nand2 gate2424(.a(gate9inter0), .b(s_268), .O(gate9inter1));
  and2  gate2425(.a(G2), .b(G1), .O(gate9inter2));
  inv1  gate2426(.a(s_268), .O(gate9inter3));
  inv1  gate2427(.a(s_269), .O(gate9inter4));
  nand2 gate2428(.a(gate9inter4), .b(gate9inter3), .O(gate9inter5));
  nor2  gate2429(.a(gate9inter5), .b(gate9inter2), .O(gate9inter6));
  inv1  gate2430(.a(G1), .O(gate9inter7));
  inv1  gate2431(.a(G2), .O(gate9inter8));
  nand2 gate2432(.a(gate9inter8), .b(gate9inter7), .O(gate9inter9));
  nand2 gate2433(.a(s_269), .b(gate9inter3), .O(gate9inter10));
  nor2  gate2434(.a(gate9inter10), .b(gate9inter9), .O(gate9inter11));
  nor2  gate2435(.a(gate9inter11), .b(gate9inter6), .O(gate9inter12));
  nand2 gate2436(.a(gate9inter12), .b(gate9inter1), .O(G266));

  xor2  gate3025(.a(G4), .b(G3), .O(gate10inter0));
  nand2 gate3026(.a(gate10inter0), .b(s_354), .O(gate10inter1));
  and2  gate3027(.a(G4), .b(G3), .O(gate10inter2));
  inv1  gate3028(.a(s_354), .O(gate10inter3));
  inv1  gate3029(.a(s_355), .O(gate10inter4));
  nand2 gate3030(.a(gate10inter4), .b(gate10inter3), .O(gate10inter5));
  nor2  gate3031(.a(gate10inter5), .b(gate10inter2), .O(gate10inter6));
  inv1  gate3032(.a(G3), .O(gate10inter7));
  inv1  gate3033(.a(G4), .O(gate10inter8));
  nand2 gate3034(.a(gate10inter8), .b(gate10inter7), .O(gate10inter9));
  nand2 gate3035(.a(s_355), .b(gate10inter3), .O(gate10inter10));
  nor2  gate3036(.a(gate10inter10), .b(gate10inter9), .O(gate10inter11));
  nor2  gate3037(.a(gate10inter11), .b(gate10inter6), .O(gate10inter12));
  nand2 gate3038(.a(gate10inter12), .b(gate10inter1), .O(G269));
nand2 gate11( .a(G5), .b(G6), .O(G272) );

  xor2  gate1135(.a(G8), .b(G7), .O(gate12inter0));
  nand2 gate1136(.a(gate12inter0), .b(s_84), .O(gate12inter1));
  and2  gate1137(.a(G8), .b(G7), .O(gate12inter2));
  inv1  gate1138(.a(s_84), .O(gate12inter3));
  inv1  gate1139(.a(s_85), .O(gate12inter4));
  nand2 gate1140(.a(gate12inter4), .b(gate12inter3), .O(gate12inter5));
  nor2  gate1141(.a(gate12inter5), .b(gate12inter2), .O(gate12inter6));
  inv1  gate1142(.a(G7), .O(gate12inter7));
  inv1  gate1143(.a(G8), .O(gate12inter8));
  nand2 gate1144(.a(gate12inter8), .b(gate12inter7), .O(gate12inter9));
  nand2 gate1145(.a(s_85), .b(gate12inter3), .O(gate12inter10));
  nor2  gate1146(.a(gate12inter10), .b(gate12inter9), .O(gate12inter11));
  nor2  gate1147(.a(gate12inter11), .b(gate12inter6), .O(gate12inter12));
  nand2 gate1148(.a(gate12inter12), .b(gate12inter1), .O(G275));
nand2 gate13( .a(G9), .b(G10), .O(G278) );
nand2 gate14( .a(G11), .b(G12), .O(G281) );
nand2 gate15( .a(G13), .b(G14), .O(G284) );
nand2 gate16( .a(G15), .b(G16), .O(G287) );
nand2 gate17( .a(G17), .b(G18), .O(G290) );
nand2 gate18( .a(G19), .b(G20), .O(G293) );
nand2 gate19( .a(G21), .b(G22), .O(G296) );
nand2 gate20( .a(G23), .b(G24), .O(G299) );
nand2 gate21( .a(G25), .b(G26), .O(G302) );
nand2 gate22( .a(G27), .b(G28), .O(G305) );
nand2 gate23( .a(G29), .b(G30), .O(G308) );
nand2 gate24( .a(G31), .b(G32), .O(G311) );

  xor2  gate813(.a(G5), .b(G1), .O(gate25inter0));
  nand2 gate814(.a(gate25inter0), .b(s_38), .O(gate25inter1));
  and2  gate815(.a(G5), .b(G1), .O(gate25inter2));
  inv1  gate816(.a(s_38), .O(gate25inter3));
  inv1  gate817(.a(s_39), .O(gate25inter4));
  nand2 gate818(.a(gate25inter4), .b(gate25inter3), .O(gate25inter5));
  nor2  gate819(.a(gate25inter5), .b(gate25inter2), .O(gate25inter6));
  inv1  gate820(.a(G1), .O(gate25inter7));
  inv1  gate821(.a(G5), .O(gate25inter8));
  nand2 gate822(.a(gate25inter8), .b(gate25inter7), .O(gate25inter9));
  nand2 gate823(.a(s_39), .b(gate25inter3), .O(gate25inter10));
  nor2  gate824(.a(gate25inter10), .b(gate25inter9), .O(gate25inter11));
  nor2  gate825(.a(gate25inter11), .b(gate25inter6), .O(gate25inter12));
  nand2 gate826(.a(gate25inter12), .b(gate25inter1), .O(G314));
nand2 gate26( .a(G9), .b(G13), .O(G317) );
nand2 gate27( .a(G2), .b(G6), .O(G320) );
nand2 gate28( .a(G10), .b(G14), .O(G323) );

  xor2  gate2745(.a(G7), .b(G3), .O(gate29inter0));
  nand2 gate2746(.a(gate29inter0), .b(s_314), .O(gate29inter1));
  and2  gate2747(.a(G7), .b(G3), .O(gate29inter2));
  inv1  gate2748(.a(s_314), .O(gate29inter3));
  inv1  gate2749(.a(s_315), .O(gate29inter4));
  nand2 gate2750(.a(gate29inter4), .b(gate29inter3), .O(gate29inter5));
  nor2  gate2751(.a(gate29inter5), .b(gate29inter2), .O(gate29inter6));
  inv1  gate2752(.a(G3), .O(gate29inter7));
  inv1  gate2753(.a(G7), .O(gate29inter8));
  nand2 gate2754(.a(gate29inter8), .b(gate29inter7), .O(gate29inter9));
  nand2 gate2755(.a(s_315), .b(gate29inter3), .O(gate29inter10));
  nor2  gate2756(.a(gate29inter10), .b(gate29inter9), .O(gate29inter11));
  nor2  gate2757(.a(gate29inter11), .b(gate29inter6), .O(gate29inter12));
  nand2 gate2758(.a(gate29inter12), .b(gate29inter1), .O(G326));

  xor2  gate2787(.a(G15), .b(G11), .O(gate30inter0));
  nand2 gate2788(.a(gate30inter0), .b(s_320), .O(gate30inter1));
  and2  gate2789(.a(G15), .b(G11), .O(gate30inter2));
  inv1  gate2790(.a(s_320), .O(gate30inter3));
  inv1  gate2791(.a(s_321), .O(gate30inter4));
  nand2 gate2792(.a(gate30inter4), .b(gate30inter3), .O(gate30inter5));
  nor2  gate2793(.a(gate30inter5), .b(gate30inter2), .O(gate30inter6));
  inv1  gate2794(.a(G11), .O(gate30inter7));
  inv1  gate2795(.a(G15), .O(gate30inter8));
  nand2 gate2796(.a(gate30inter8), .b(gate30inter7), .O(gate30inter9));
  nand2 gate2797(.a(s_321), .b(gate30inter3), .O(gate30inter10));
  nor2  gate2798(.a(gate30inter10), .b(gate30inter9), .O(gate30inter11));
  nor2  gate2799(.a(gate30inter11), .b(gate30inter6), .O(gate30inter12));
  nand2 gate2800(.a(gate30inter12), .b(gate30inter1), .O(G329));

  xor2  gate2003(.a(G8), .b(G4), .O(gate31inter0));
  nand2 gate2004(.a(gate31inter0), .b(s_208), .O(gate31inter1));
  and2  gate2005(.a(G8), .b(G4), .O(gate31inter2));
  inv1  gate2006(.a(s_208), .O(gate31inter3));
  inv1  gate2007(.a(s_209), .O(gate31inter4));
  nand2 gate2008(.a(gate31inter4), .b(gate31inter3), .O(gate31inter5));
  nor2  gate2009(.a(gate31inter5), .b(gate31inter2), .O(gate31inter6));
  inv1  gate2010(.a(G4), .O(gate31inter7));
  inv1  gate2011(.a(G8), .O(gate31inter8));
  nand2 gate2012(.a(gate31inter8), .b(gate31inter7), .O(gate31inter9));
  nand2 gate2013(.a(s_209), .b(gate31inter3), .O(gate31inter10));
  nor2  gate2014(.a(gate31inter10), .b(gate31inter9), .O(gate31inter11));
  nor2  gate2015(.a(gate31inter11), .b(gate31inter6), .O(gate31inter12));
  nand2 gate2016(.a(gate31inter12), .b(gate31inter1), .O(G332));

  xor2  gate2073(.a(G16), .b(G12), .O(gate32inter0));
  nand2 gate2074(.a(gate32inter0), .b(s_218), .O(gate32inter1));
  and2  gate2075(.a(G16), .b(G12), .O(gate32inter2));
  inv1  gate2076(.a(s_218), .O(gate32inter3));
  inv1  gate2077(.a(s_219), .O(gate32inter4));
  nand2 gate2078(.a(gate32inter4), .b(gate32inter3), .O(gate32inter5));
  nor2  gate2079(.a(gate32inter5), .b(gate32inter2), .O(gate32inter6));
  inv1  gate2080(.a(G12), .O(gate32inter7));
  inv1  gate2081(.a(G16), .O(gate32inter8));
  nand2 gate2082(.a(gate32inter8), .b(gate32inter7), .O(gate32inter9));
  nand2 gate2083(.a(s_219), .b(gate32inter3), .O(gate32inter10));
  nor2  gate2084(.a(gate32inter10), .b(gate32inter9), .O(gate32inter11));
  nor2  gate2085(.a(gate32inter11), .b(gate32inter6), .O(gate32inter12));
  nand2 gate2086(.a(gate32inter12), .b(gate32inter1), .O(G335));

  xor2  gate2213(.a(G21), .b(G17), .O(gate33inter0));
  nand2 gate2214(.a(gate33inter0), .b(s_238), .O(gate33inter1));
  and2  gate2215(.a(G21), .b(G17), .O(gate33inter2));
  inv1  gate2216(.a(s_238), .O(gate33inter3));
  inv1  gate2217(.a(s_239), .O(gate33inter4));
  nand2 gate2218(.a(gate33inter4), .b(gate33inter3), .O(gate33inter5));
  nor2  gate2219(.a(gate33inter5), .b(gate33inter2), .O(gate33inter6));
  inv1  gate2220(.a(G17), .O(gate33inter7));
  inv1  gate2221(.a(G21), .O(gate33inter8));
  nand2 gate2222(.a(gate33inter8), .b(gate33inter7), .O(gate33inter9));
  nand2 gate2223(.a(s_239), .b(gate33inter3), .O(gate33inter10));
  nor2  gate2224(.a(gate33inter10), .b(gate33inter9), .O(gate33inter11));
  nor2  gate2225(.a(gate33inter11), .b(gate33inter6), .O(gate33inter12));
  nand2 gate2226(.a(gate33inter12), .b(gate33inter1), .O(G338));
nand2 gate34( .a(G25), .b(G29), .O(G341) );
nand2 gate35( .a(G18), .b(G22), .O(G344) );
nand2 gate36( .a(G26), .b(G30), .O(G347) );

  xor2  gate869(.a(G23), .b(G19), .O(gate37inter0));
  nand2 gate870(.a(gate37inter0), .b(s_46), .O(gate37inter1));
  and2  gate871(.a(G23), .b(G19), .O(gate37inter2));
  inv1  gate872(.a(s_46), .O(gate37inter3));
  inv1  gate873(.a(s_47), .O(gate37inter4));
  nand2 gate874(.a(gate37inter4), .b(gate37inter3), .O(gate37inter5));
  nor2  gate875(.a(gate37inter5), .b(gate37inter2), .O(gate37inter6));
  inv1  gate876(.a(G19), .O(gate37inter7));
  inv1  gate877(.a(G23), .O(gate37inter8));
  nand2 gate878(.a(gate37inter8), .b(gate37inter7), .O(gate37inter9));
  nand2 gate879(.a(s_47), .b(gate37inter3), .O(gate37inter10));
  nor2  gate880(.a(gate37inter10), .b(gate37inter9), .O(gate37inter11));
  nor2  gate881(.a(gate37inter11), .b(gate37inter6), .O(gate37inter12));
  nand2 gate882(.a(gate37inter12), .b(gate37inter1), .O(G350));

  xor2  gate911(.a(G31), .b(G27), .O(gate38inter0));
  nand2 gate912(.a(gate38inter0), .b(s_52), .O(gate38inter1));
  and2  gate913(.a(G31), .b(G27), .O(gate38inter2));
  inv1  gate914(.a(s_52), .O(gate38inter3));
  inv1  gate915(.a(s_53), .O(gate38inter4));
  nand2 gate916(.a(gate38inter4), .b(gate38inter3), .O(gate38inter5));
  nor2  gate917(.a(gate38inter5), .b(gate38inter2), .O(gate38inter6));
  inv1  gate918(.a(G27), .O(gate38inter7));
  inv1  gate919(.a(G31), .O(gate38inter8));
  nand2 gate920(.a(gate38inter8), .b(gate38inter7), .O(gate38inter9));
  nand2 gate921(.a(s_53), .b(gate38inter3), .O(gate38inter10));
  nor2  gate922(.a(gate38inter10), .b(gate38inter9), .O(gate38inter11));
  nor2  gate923(.a(gate38inter11), .b(gate38inter6), .O(gate38inter12));
  nand2 gate924(.a(gate38inter12), .b(gate38inter1), .O(G353));

  xor2  gate2675(.a(G24), .b(G20), .O(gate39inter0));
  nand2 gate2676(.a(gate39inter0), .b(s_304), .O(gate39inter1));
  and2  gate2677(.a(G24), .b(G20), .O(gate39inter2));
  inv1  gate2678(.a(s_304), .O(gate39inter3));
  inv1  gate2679(.a(s_305), .O(gate39inter4));
  nand2 gate2680(.a(gate39inter4), .b(gate39inter3), .O(gate39inter5));
  nor2  gate2681(.a(gate39inter5), .b(gate39inter2), .O(gate39inter6));
  inv1  gate2682(.a(G20), .O(gate39inter7));
  inv1  gate2683(.a(G24), .O(gate39inter8));
  nand2 gate2684(.a(gate39inter8), .b(gate39inter7), .O(gate39inter9));
  nand2 gate2685(.a(s_305), .b(gate39inter3), .O(gate39inter10));
  nor2  gate2686(.a(gate39inter10), .b(gate39inter9), .O(gate39inter11));
  nor2  gate2687(.a(gate39inter11), .b(gate39inter6), .O(gate39inter12));
  nand2 gate2688(.a(gate39inter12), .b(gate39inter1), .O(G356));

  xor2  gate715(.a(G32), .b(G28), .O(gate40inter0));
  nand2 gate716(.a(gate40inter0), .b(s_24), .O(gate40inter1));
  and2  gate717(.a(G32), .b(G28), .O(gate40inter2));
  inv1  gate718(.a(s_24), .O(gate40inter3));
  inv1  gate719(.a(s_25), .O(gate40inter4));
  nand2 gate720(.a(gate40inter4), .b(gate40inter3), .O(gate40inter5));
  nor2  gate721(.a(gate40inter5), .b(gate40inter2), .O(gate40inter6));
  inv1  gate722(.a(G28), .O(gate40inter7));
  inv1  gate723(.a(G32), .O(gate40inter8));
  nand2 gate724(.a(gate40inter8), .b(gate40inter7), .O(gate40inter9));
  nand2 gate725(.a(s_25), .b(gate40inter3), .O(gate40inter10));
  nor2  gate726(.a(gate40inter10), .b(gate40inter9), .O(gate40inter11));
  nor2  gate727(.a(gate40inter11), .b(gate40inter6), .O(gate40inter12));
  nand2 gate728(.a(gate40inter12), .b(gate40inter1), .O(G359));
nand2 gate41( .a(G1), .b(G266), .O(G362) );

  xor2  gate547(.a(G266), .b(G2), .O(gate42inter0));
  nand2 gate548(.a(gate42inter0), .b(s_0), .O(gate42inter1));
  and2  gate549(.a(G266), .b(G2), .O(gate42inter2));
  inv1  gate550(.a(s_0), .O(gate42inter3));
  inv1  gate551(.a(s_1), .O(gate42inter4));
  nand2 gate552(.a(gate42inter4), .b(gate42inter3), .O(gate42inter5));
  nor2  gate553(.a(gate42inter5), .b(gate42inter2), .O(gate42inter6));
  inv1  gate554(.a(G2), .O(gate42inter7));
  inv1  gate555(.a(G266), .O(gate42inter8));
  nand2 gate556(.a(gate42inter8), .b(gate42inter7), .O(gate42inter9));
  nand2 gate557(.a(s_1), .b(gate42inter3), .O(gate42inter10));
  nor2  gate558(.a(gate42inter10), .b(gate42inter9), .O(gate42inter11));
  nor2  gate559(.a(gate42inter11), .b(gate42inter6), .O(gate42inter12));
  nand2 gate560(.a(gate42inter12), .b(gate42inter1), .O(G363));

  xor2  gate1975(.a(G269), .b(G3), .O(gate43inter0));
  nand2 gate1976(.a(gate43inter0), .b(s_204), .O(gate43inter1));
  and2  gate1977(.a(G269), .b(G3), .O(gate43inter2));
  inv1  gate1978(.a(s_204), .O(gate43inter3));
  inv1  gate1979(.a(s_205), .O(gate43inter4));
  nand2 gate1980(.a(gate43inter4), .b(gate43inter3), .O(gate43inter5));
  nor2  gate1981(.a(gate43inter5), .b(gate43inter2), .O(gate43inter6));
  inv1  gate1982(.a(G3), .O(gate43inter7));
  inv1  gate1983(.a(G269), .O(gate43inter8));
  nand2 gate1984(.a(gate43inter8), .b(gate43inter7), .O(gate43inter9));
  nand2 gate1985(.a(s_205), .b(gate43inter3), .O(gate43inter10));
  nor2  gate1986(.a(gate43inter10), .b(gate43inter9), .O(gate43inter11));
  nor2  gate1987(.a(gate43inter11), .b(gate43inter6), .O(gate43inter12));
  nand2 gate1988(.a(gate43inter12), .b(gate43inter1), .O(G364));
nand2 gate44( .a(G4), .b(G269), .O(G365) );

  xor2  gate2479(.a(G272), .b(G5), .O(gate45inter0));
  nand2 gate2480(.a(gate45inter0), .b(s_276), .O(gate45inter1));
  and2  gate2481(.a(G272), .b(G5), .O(gate45inter2));
  inv1  gate2482(.a(s_276), .O(gate45inter3));
  inv1  gate2483(.a(s_277), .O(gate45inter4));
  nand2 gate2484(.a(gate45inter4), .b(gate45inter3), .O(gate45inter5));
  nor2  gate2485(.a(gate45inter5), .b(gate45inter2), .O(gate45inter6));
  inv1  gate2486(.a(G5), .O(gate45inter7));
  inv1  gate2487(.a(G272), .O(gate45inter8));
  nand2 gate2488(.a(gate45inter8), .b(gate45inter7), .O(gate45inter9));
  nand2 gate2489(.a(s_277), .b(gate45inter3), .O(gate45inter10));
  nor2  gate2490(.a(gate45inter10), .b(gate45inter9), .O(gate45inter11));
  nor2  gate2491(.a(gate45inter11), .b(gate45inter6), .O(gate45inter12));
  nand2 gate2492(.a(gate45inter12), .b(gate45inter1), .O(G366));
nand2 gate46( .a(G6), .b(G272), .O(G367) );
nand2 gate47( .a(G7), .b(G275), .O(G368) );
nand2 gate48( .a(G8), .b(G275), .O(G369) );

  xor2  gate2969(.a(G278), .b(G9), .O(gate49inter0));
  nand2 gate2970(.a(gate49inter0), .b(s_346), .O(gate49inter1));
  and2  gate2971(.a(G278), .b(G9), .O(gate49inter2));
  inv1  gate2972(.a(s_346), .O(gate49inter3));
  inv1  gate2973(.a(s_347), .O(gate49inter4));
  nand2 gate2974(.a(gate49inter4), .b(gate49inter3), .O(gate49inter5));
  nor2  gate2975(.a(gate49inter5), .b(gate49inter2), .O(gate49inter6));
  inv1  gate2976(.a(G9), .O(gate49inter7));
  inv1  gate2977(.a(G278), .O(gate49inter8));
  nand2 gate2978(.a(gate49inter8), .b(gate49inter7), .O(gate49inter9));
  nand2 gate2979(.a(s_347), .b(gate49inter3), .O(gate49inter10));
  nor2  gate2980(.a(gate49inter10), .b(gate49inter9), .O(gate49inter11));
  nor2  gate2981(.a(gate49inter11), .b(gate49inter6), .O(gate49inter12));
  nand2 gate2982(.a(gate49inter12), .b(gate49inter1), .O(G370));
nand2 gate50( .a(G10), .b(G278), .O(G371) );

  xor2  gate2871(.a(G281), .b(G11), .O(gate51inter0));
  nand2 gate2872(.a(gate51inter0), .b(s_332), .O(gate51inter1));
  and2  gate2873(.a(G281), .b(G11), .O(gate51inter2));
  inv1  gate2874(.a(s_332), .O(gate51inter3));
  inv1  gate2875(.a(s_333), .O(gate51inter4));
  nand2 gate2876(.a(gate51inter4), .b(gate51inter3), .O(gate51inter5));
  nor2  gate2877(.a(gate51inter5), .b(gate51inter2), .O(gate51inter6));
  inv1  gate2878(.a(G11), .O(gate51inter7));
  inv1  gate2879(.a(G281), .O(gate51inter8));
  nand2 gate2880(.a(gate51inter8), .b(gate51inter7), .O(gate51inter9));
  nand2 gate2881(.a(s_333), .b(gate51inter3), .O(gate51inter10));
  nor2  gate2882(.a(gate51inter10), .b(gate51inter9), .O(gate51inter11));
  nor2  gate2883(.a(gate51inter11), .b(gate51inter6), .O(gate51inter12));
  nand2 gate2884(.a(gate51inter12), .b(gate51inter1), .O(G372));
nand2 gate52( .a(G12), .b(G281), .O(G373) );

  xor2  gate1597(.a(G284), .b(G13), .O(gate53inter0));
  nand2 gate1598(.a(gate53inter0), .b(s_150), .O(gate53inter1));
  and2  gate1599(.a(G284), .b(G13), .O(gate53inter2));
  inv1  gate1600(.a(s_150), .O(gate53inter3));
  inv1  gate1601(.a(s_151), .O(gate53inter4));
  nand2 gate1602(.a(gate53inter4), .b(gate53inter3), .O(gate53inter5));
  nor2  gate1603(.a(gate53inter5), .b(gate53inter2), .O(gate53inter6));
  inv1  gate1604(.a(G13), .O(gate53inter7));
  inv1  gate1605(.a(G284), .O(gate53inter8));
  nand2 gate1606(.a(gate53inter8), .b(gate53inter7), .O(gate53inter9));
  nand2 gate1607(.a(s_151), .b(gate53inter3), .O(gate53inter10));
  nor2  gate1608(.a(gate53inter10), .b(gate53inter9), .O(gate53inter11));
  nor2  gate1609(.a(gate53inter11), .b(gate53inter6), .O(gate53inter12));
  nand2 gate1610(.a(gate53inter12), .b(gate53inter1), .O(G374));
nand2 gate54( .a(G14), .b(G284), .O(G375) );

  xor2  gate2801(.a(G287), .b(G15), .O(gate55inter0));
  nand2 gate2802(.a(gate55inter0), .b(s_322), .O(gate55inter1));
  and2  gate2803(.a(G287), .b(G15), .O(gate55inter2));
  inv1  gate2804(.a(s_322), .O(gate55inter3));
  inv1  gate2805(.a(s_323), .O(gate55inter4));
  nand2 gate2806(.a(gate55inter4), .b(gate55inter3), .O(gate55inter5));
  nor2  gate2807(.a(gate55inter5), .b(gate55inter2), .O(gate55inter6));
  inv1  gate2808(.a(G15), .O(gate55inter7));
  inv1  gate2809(.a(G287), .O(gate55inter8));
  nand2 gate2810(.a(gate55inter8), .b(gate55inter7), .O(gate55inter9));
  nand2 gate2811(.a(s_323), .b(gate55inter3), .O(gate55inter10));
  nor2  gate2812(.a(gate55inter10), .b(gate55inter9), .O(gate55inter11));
  nor2  gate2813(.a(gate55inter11), .b(gate55inter6), .O(gate55inter12));
  nand2 gate2814(.a(gate55inter12), .b(gate55inter1), .O(G376));

  xor2  gate1863(.a(G287), .b(G16), .O(gate56inter0));
  nand2 gate1864(.a(gate56inter0), .b(s_188), .O(gate56inter1));
  and2  gate1865(.a(G287), .b(G16), .O(gate56inter2));
  inv1  gate1866(.a(s_188), .O(gate56inter3));
  inv1  gate1867(.a(s_189), .O(gate56inter4));
  nand2 gate1868(.a(gate56inter4), .b(gate56inter3), .O(gate56inter5));
  nor2  gate1869(.a(gate56inter5), .b(gate56inter2), .O(gate56inter6));
  inv1  gate1870(.a(G16), .O(gate56inter7));
  inv1  gate1871(.a(G287), .O(gate56inter8));
  nand2 gate1872(.a(gate56inter8), .b(gate56inter7), .O(gate56inter9));
  nand2 gate1873(.a(s_189), .b(gate56inter3), .O(gate56inter10));
  nor2  gate1874(.a(gate56inter10), .b(gate56inter9), .O(gate56inter11));
  nor2  gate1875(.a(gate56inter11), .b(gate56inter6), .O(gate56inter12));
  nand2 gate1876(.a(gate56inter12), .b(gate56inter1), .O(G377));

  xor2  gate1961(.a(G290), .b(G17), .O(gate57inter0));
  nand2 gate1962(.a(gate57inter0), .b(s_202), .O(gate57inter1));
  and2  gate1963(.a(G290), .b(G17), .O(gate57inter2));
  inv1  gate1964(.a(s_202), .O(gate57inter3));
  inv1  gate1965(.a(s_203), .O(gate57inter4));
  nand2 gate1966(.a(gate57inter4), .b(gate57inter3), .O(gate57inter5));
  nor2  gate1967(.a(gate57inter5), .b(gate57inter2), .O(gate57inter6));
  inv1  gate1968(.a(G17), .O(gate57inter7));
  inv1  gate1969(.a(G290), .O(gate57inter8));
  nand2 gate1970(.a(gate57inter8), .b(gate57inter7), .O(gate57inter9));
  nand2 gate1971(.a(s_203), .b(gate57inter3), .O(gate57inter10));
  nor2  gate1972(.a(gate57inter10), .b(gate57inter9), .O(gate57inter11));
  nor2  gate1973(.a(gate57inter11), .b(gate57inter6), .O(gate57inter12));
  nand2 gate1974(.a(gate57inter12), .b(gate57inter1), .O(G378));

  xor2  gate1331(.a(G290), .b(G18), .O(gate58inter0));
  nand2 gate1332(.a(gate58inter0), .b(s_112), .O(gate58inter1));
  and2  gate1333(.a(G290), .b(G18), .O(gate58inter2));
  inv1  gate1334(.a(s_112), .O(gate58inter3));
  inv1  gate1335(.a(s_113), .O(gate58inter4));
  nand2 gate1336(.a(gate58inter4), .b(gate58inter3), .O(gate58inter5));
  nor2  gate1337(.a(gate58inter5), .b(gate58inter2), .O(gate58inter6));
  inv1  gate1338(.a(G18), .O(gate58inter7));
  inv1  gate1339(.a(G290), .O(gate58inter8));
  nand2 gate1340(.a(gate58inter8), .b(gate58inter7), .O(gate58inter9));
  nand2 gate1341(.a(s_113), .b(gate58inter3), .O(gate58inter10));
  nor2  gate1342(.a(gate58inter10), .b(gate58inter9), .O(gate58inter11));
  nor2  gate1343(.a(gate58inter11), .b(gate58inter6), .O(gate58inter12));
  nand2 gate1344(.a(gate58inter12), .b(gate58inter1), .O(G379));
nand2 gate59( .a(G19), .b(G293), .O(G380) );

  xor2  gate757(.a(G293), .b(G20), .O(gate60inter0));
  nand2 gate758(.a(gate60inter0), .b(s_30), .O(gate60inter1));
  and2  gate759(.a(G293), .b(G20), .O(gate60inter2));
  inv1  gate760(.a(s_30), .O(gate60inter3));
  inv1  gate761(.a(s_31), .O(gate60inter4));
  nand2 gate762(.a(gate60inter4), .b(gate60inter3), .O(gate60inter5));
  nor2  gate763(.a(gate60inter5), .b(gate60inter2), .O(gate60inter6));
  inv1  gate764(.a(G20), .O(gate60inter7));
  inv1  gate765(.a(G293), .O(gate60inter8));
  nand2 gate766(.a(gate60inter8), .b(gate60inter7), .O(gate60inter9));
  nand2 gate767(.a(s_31), .b(gate60inter3), .O(gate60inter10));
  nor2  gate768(.a(gate60inter10), .b(gate60inter9), .O(gate60inter11));
  nor2  gate769(.a(gate60inter11), .b(gate60inter6), .O(gate60inter12));
  nand2 gate770(.a(gate60inter12), .b(gate60inter1), .O(G381));

  xor2  gate981(.a(G296), .b(G21), .O(gate61inter0));
  nand2 gate982(.a(gate61inter0), .b(s_62), .O(gate61inter1));
  and2  gate983(.a(G296), .b(G21), .O(gate61inter2));
  inv1  gate984(.a(s_62), .O(gate61inter3));
  inv1  gate985(.a(s_63), .O(gate61inter4));
  nand2 gate986(.a(gate61inter4), .b(gate61inter3), .O(gate61inter5));
  nor2  gate987(.a(gate61inter5), .b(gate61inter2), .O(gate61inter6));
  inv1  gate988(.a(G21), .O(gate61inter7));
  inv1  gate989(.a(G296), .O(gate61inter8));
  nand2 gate990(.a(gate61inter8), .b(gate61inter7), .O(gate61inter9));
  nand2 gate991(.a(s_63), .b(gate61inter3), .O(gate61inter10));
  nor2  gate992(.a(gate61inter10), .b(gate61inter9), .O(gate61inter11));
  nor2  gate993(.a(gate61inter11), .b(gate61inter6), .O(gate61inter12));
  nand2 gate994(.a(gate61inter12), .b(gate61inter1), .O(G382));
nand2 gate62( .a(G22), .b(G296), .O(G383) );

  xor2  gate561(.a(G299), .b(G23), .O(gate63inter0));
  nand2 gate562(.a(gate63inter0), .b(s_2), .O(gate63inter1));
  and2  gate563(.a(G299), .b(G23), .O(gate63inter2));
  inv1  gate564(.a(s_2), .O(gate63inter3));
  inv1  gate565(.a(s_3), .O(gate63inter4));
  nand2 gate566(.a(gate63inter4), .b(gate63inter3), .O(gate63inter5));
  nor2  gate567(.a(gate63inter5), .b(gate63inter2), .O(gate63inter6));
  inv1  gate568(.a(G23), .O(gate63inter7));
  inv1  gate569(.a(G299), .O(gate63inter8));
  nand2 gate570(.a(gate63inter8), .b(gate63inter7), .O(gate63inter9));
  nand2 gate571(.a(s_3), .b(gate63inter3), .O(gate63inter10));
  nor2  gate572(.a(gate63inter10), .b(gate63inter9), .O(gate63inter11));
  nor2  gate573(.a(gate63inter11), .b(gate63inter6), .O(gate63inter12));
  nand2 gate574(.a(gate63inter12), .b(gate63inter1), .O(G384));

  xor2  gate2941(.a(G299), .b(G24), .O(gate64inter0));
  nand2 gate2942(.a(gate64inter0), .b(s_342), .O(gate64inter1));
  and2  gate2943(.a(G299), .b(G24), .O(gate64inter2));
  inv1  gate2944(.a(s_342), .O(gate64inter3));
  inv1  gate2945(.a(s_343), .O(gate64inter4));
  nand2 gate2946(.a(gate64inter4), .b(gate64inter3), .O(gate64inter5));
  nor2  gate2947(.a(gate64inter5), .b(gate64inter2), .O(gate64inter6));
  inv1  gate2948(.a(G24), .O(gate64inter7));
  inv1  gate2949(.a(G299), .O(gate64inter8));
  nand2 gate2950(.a(gate64inter8), .b(gate64inter7), .O(gate64inter9));
  nand2 gate2951(.a(s_343), .b(gate64inter3), .O(gate64inter10));
  nor2  gate2952(.a(gate64inter10), .b(gate64inter9), .O(gate64inter11));
  nor2  gate2953(.a(gate64inter11), .b(gate64inter6), .O(gate64inter12));
  nand2 gate2954(.a(gate64inter12), .b(gate64inter1), .O(G385));
nand2 gate65( .a(G25), .b(G302), .O(G386) );
nand2 gate66( .a(G26), .b(G302), .O(G387) );

  xor2  gate925(.a(G305), .b(G27), .O(gate67inter0));
  nand2 gate926(.a(gate67inter0), .b(s_54), .O(gate67inter1));
  and2  gate927(.a(G305), .b(G27), .O(gate67inter2));
  inv1  gate928(.a(s_54), .O(gate67inter3));
  inv1  gate929(.a(s_55), .O(gate67inter4));
  nand2 gate930(.a(gate67inter4), .b(gate67inter3), .O(gate67inter5));
  nor2  gate931(.a(gate67inter5), .b(gate67inter2), .O(gate67inter6));
  inv1  gate932(.a(G27), .O(gate67inter7));
  inv1  gate933(.a(G305), .O(gate67inter8));
  nand2 gate934(.a(gate67inter8), .b(gate67inter7), .O(gate67inter9));
  nand2 gate935(.a(s_55), .b(gate67inter3), .O(gate67inter10));
  nor2  gate936(.a(gate67inter10), .b(gate67inter9), .O(gate67inter11));
  nor2  gate937(.a(gate67inter11), .b(gate67inter6), .O(gate67inter12));
  nand2 gate938(.a(gate67inter12), .b(gate67inter1), .O(G388));
nand2 gate68( .a(G28), .b(G305), .O(G389) );
nand2 gate69( .a(G29), .b(G308), .O(G390) );
nand2 gate70( .a(G30), .b(G308), .O(G391) );

  xor2  gate673(.a(G311), .b(G31), .O(gate71inter0));
  nand2 gate674(.a(gate71inter0), .b(s_18), .O(gate71inter1));
  and2  gate675(.a(G311), .b(G31), .O(gate71inter2));
  inv1  gate676(.a(s_18), .O(gate71inter3));
  inv1  gate677(.a(s_19), .O(gate71inter4));
  nand2 gate678(.a(gate71inter4), .b(gate71inter3), .O(gate71inter5));
  nor2  gate679(.a(gate71inter5), .b(gate71inter2), .O(gate71inter6));
  inv1  gate680(.a(G31), .O(gate71inter7));
  inv1  gate681(.a(G311), .O(gate71inter8));
  nand2 gate682(.a(gate71inter8), .b(gate71inter7), .O(gate71inter9));
  nand2 gate683(.a(s_19), .b(gate71inter3), .O(gate71inter10));
  nor2  gate684(.a(gate71inter10), .b(gate71inter9), .O(gate71inter11));
  nor2  gate685(.a(gate71inter11), .b(gate71inter6), .O(gate71inter12));
  nand2 gate686(.a(gate71inter12), .b(gate71inter1), .O(G392));
nand2 gate72( .a(G32), .b(G311), .O(G393) );
nand2 gate73( .a(G1), .b(G314), .O(G394) );
nand2 gate74( .a(G5), .b(G314), .O(G395) );
nand2 gate75( .a(G9), .b(G317), .O(G396) );
nand2 gate76( .a(G13), .b(G317), .O(G397) );
nand2 gate77( .a(G2), .b(G320), .O(G398) );

  xor2  gate2661(.a(G320), .b(G6), .O(gate78inter0));
  nand2 gate2662(.a(gate78inter0), .b(s_302), .O(gate78inter1));
  and2  gate2663(.a(G320), .b(G6), .O(gate78inter2));
  inv1  gate2664(.a(s_302), .O(gate78inter3));
  inv1  gate2665(.a(s_303), .O(gate78inter4));
  nand2 gate2666(.a(gate78inter4), .b(gate78inter3), .O(gate78inter5));
  nor2  gate2667(.a(gate78inter5), .b(gate78inter2), .O(gate78inter6));
  inv1  gate2668(.a(G6), .O(gate78inter7));
  inv1  gate2669(.a(G320), .O(gate78inter8));
  nand2 gate2670(.a(gate78inter8), .b(gate78inter7), .O(gate78inter9));
  nand2 gate2671(.a(s_303), .b(gate78inter3), .O(gate78inter10));
  nor2  gate2672(.a(gate78inter10), .b(gate78inter9), .O(gate78inter11));
  nor2  gate2673(.a(gate78inter11), .b(gate78inter6), .O(gate78inter12));
  nand2 gate2674(.a(gate78inter12), .b(gate78inter1), .O(G399));
nand2 gate79( .a(G10), .b(G323), .O(G400) );
nand2 gate80( .a(G14), .b(G323), .O(G401) );
nand2 gate81( .a(G3), .b(G326), .O(G402) );

  xor2  gate589(.a(G326), .b(G7), .O(gate82inter0));
  nand2 gate590(.a(gate82inter0), .b(s_6), .O(gate82inter1));
  and2  gate591(.a(G326), .b(G7), .O(gate82inter2));
  inv1  gate592(.a(s_6), .O(gate82inter3));
  inv1  gate593(.a(s_7), .O(gate82inter4));
  nand2 gate594(.a(gate82inter4), .b(gate82inter3), .O(gate82inter5));
  nor2  gate595(.a(gate82inter5), .b(gate82inter2), .O(gate82inter6));
  inv1  gate596(.a(G7), .O(gate82inter7));
  inv1  gate597(.a(G326), .O(gate82inter8));
  nand2 gate598(.a(gate82inter8), .b(gate82inter7), .O(gate82inter9));
  nand2 gate599(.a(s_7), .b(gate82inter3), .O(gate82inter10));
  nor2  gate600(.a(gate82inter10), .b(gate82inter9), .O(gate82inter11));
  nor2  gate601(.a(gate82inter11), .b(gate82inter6), .O(gate82inter12));
  nand2 gate602(.a(gate82inter12), .b(gate82inter1), .O(G403));

  xor2  gate1541(.a(G329), .b(G11), .O(gate83inter0));
  nand2 gate1542(.a(gate83inter0), .b(s_142), .O(gate83inter1));
  and2  gate1543(.a(G329), .b(G11), .O(gate83inter2));
  inv1  gate1544(.a(s_142), .O(gate83inter3));
  inv1  gate1545(.a(s_143), .O(gate83inter4));
  nand2 gate1546(.a(gate83inter4), .b(gate83inter3), .O(gate83inter5));
  nor2  gate1547(.a(gate83inter5), .b(gate83inter2), .O(gate83inter6));
  inv1  gate1548(.a(G11), .O(gate83inter7));
  inv1  gate1549(.a(G329), .O(gate83inter8));
  nand2 gate1550(.a(gate83inter8), .b(gate83inter7), .O(gate83inter9));
  nand2 gate1551(.a(s_143), .b(gate83inter3), .O(gate83inter10));
  nor2  gate1552(.a(gate83inter10), .b(gate83inter9), .O(gate83inter11));
  nor2  gate1553(.a(gate83inter11), .b(gate83inter6), .O(gate83inter12));
  nand2 gate1554(.a(gate83inter12), .b(gate83inter1), .O(G404));

  xor2  gate1289(.a(G329), .b(G15), .O(gate84inter0));
  nand2 gate1290(.a(gate84inter0), .b(s_106), .O(gate84inter1));
  and2  gate1291(.a(G329), .b(G15), .O(gate84inter2));
  inv1  gate1292(.a(s_106), .O(gate84inter3));
  inv1  gate1293(.a(s_107), .O(gate84inter4));
  nand2 gate1294(.a(gate84inter4), .b(gate84inter3), .O(gate84inter5));
  nor2  gate1295(.a(gate84inter5), .b(gate84inter2), .O(gate84inter6));
  inv1  gate1296(.a(G15), .O(gate84inter7));
  inv1  gate1297(.a(G329), .O(gate84inter8));
  nand2 gate1298(.a(gate84inter8), .b(gate84inter7), .O(gate84inter9));
  nand2 gate1299(.a(s_107), .b(gate84inter3), .O(gate84inter10));
  nor2  gate1300(.a(gate84inter10), .b(gate84inter9), .O(gate84inter11));
  nor2  gate1301(.a(gate84inter11), .b(gate84inter6), .O(gate84inter12));
  nand2 gate1302(.a(gate84inter12), .b(gate84inter1), .O(G405));

  xor2  gate1429(.a(G332), .b(G4), .O(gate85inter0));
  nand2 gate1430(.a(gate85inter0), .b(s_126), .O(gate85inter1));
  and2  gate1431(.a(G332), .b(G4), .O(gate85inter2));
  inv1  gate1432(.a(s_126), .O(gate85inter3));
  inv1  gate1433(.a(s_127), .O(gate85inter4));
  nand2 gate1434(.a(gate85inter4), .b(gate85inter3), .O(gate85inter5));
  nor2  gate1435(.a(gate85inter5), .b(gate85inter2), .O(gate85inter6));
  inv1  gate1436(.a(G4), .O(gate85inter7));
  inv1  gate1437(.a(G332), .O(gate85inter8));
  nand2 gate1438(.a(gate85inter8), .b(gate85inter7), .O(gate85inter9));
  nand2 gate1439(.a(s_127), .b(gate85inter3), .O(gate85inter10));
  nor2  gate1440(.a(gate85inter10), .b(gate85inter9), .O(gate85inter11));
  nor2  gate1441(.a(gate85inter11), .b(gate85inter6), .O(gate85inter12));
  nand2 gate1442(.a(gate85inter12), .b(gate85inter1), .O(G406));

  xor2  gate1527(.a(G332), .b(G8), .O(gate86inter0));
  nand2 gate1528(.a(gate86inter0), .b(s_140), .O(gate86inter1));
  and2  gate1529(.a(G332), .b(G8), .O(gate86inter2));
  inv1  gate1530(.a(s_140), .O(gate86inter3));
  inv1  gate1531(.a(s_141), .O(gate86inter4));
  nand2 gate1532(.a(gate86inter4), .b(gate86inter3), .O(gate86inter5));
  nor2  gate1533(.a(gate86inter5), .b(gate86inter2), .O(gate86inter6));
  inv1  gate1534(.a(G8), .O(gate86inter7));
  inv1  gate1535(.a(G332), .O(gate86inter8));
  nand2 gate1536(.a(gate86inter8), .b(gate86inter7), .O(gate86inter9));
  nand2 gate1537(.a(s_141), .b(gate86inter3), .O(gate86inter10));
  nor2  gate1538(.a(gate86inter10), .b(gate86inter9), .O(gate86inter11));
  nor2  gate1539(.a(gate86inter11), .b(gate86inter6), .O(gate86inter12));
  nand2 gate1540(.a(gate86inter12), .b(gate86inter1), .O(G407));
nand2 gate87( .a(G12), .b(G335), .O(G408) );
nand2 gate88( .a(G16), .b(G335), .O(G409) );
nand2 gate89( .a(G17), .b(G338), .O(G410) );
nand2 gate90( .a(G21), .b(G338), .O(G411) );

  xor2  gate2269(.a(G341), .b(G25), .O(gate91inter0));
  nand2 gate2270(.a(gate91inter0), .b(s_246), .O(gate91inter1));
  and2  gate2271(.a(G341), .b(G25), .O(gate91inter2));
  inv1  gate2272(.a(s_246), .O(gate91inter3));
  inv1  gate2273(.a(s_247), .O(gate91inter4));
  nand2 gate2274(.a(gate91inter4), .b(gate91inter3), .O(gate91inter5));
  nor2  gate2275(.a(gate91inter5), .b(gate91inter2), .O(gate91inter6));
  inv1  gate2276(.a(G25), .O(gate91inter7));
  inv1  gate2277(.a(G341), .O(gate91inter8));
  nand2 gate2278(.a(gate91inter8), .b(gate91inter7), .O(gate91inter9));
  nand2 gate2279(.a(s_247), .b(gate91inter3), .O(gate91inter10));
  nor2  gate2280(.a(gate91inter10), .b(gate91inter9), .O(gate91inter11));
  nor2  gate2281(.a(gate91inter11), .b(gate91inter6), .O(gate91inter12));
  nand2 gate2282(.a(gate91inter12), .b(gate91inter1), .O(G412));

  xor2  gate2885(.a(G341), .b(G29), .O(gate92inter0));
  nand2 gate2886(.a(gate92inter0), .b(s_334), .O(gate92inter1));
  and2  gate2887(.a(G341), .b(G29), .O(gate92inter2));
  inv1  gate2888(.a(s_334), .O(gate92inter3));
  inv1  gate2889(.a(s_335), .O(gate92inter4));
  nand2 gate2890(.a(gate92inter4), .b(gate92inter3), .O(gate92inter5));
  nor2  gate2891(.a(gate92inter5), .b(gate92inter2), .O(gate92inter6));
  inv1  gate2892(.a(G29), .O(gate92inter7));
  inv1  gate2893(.a(G341), .O(gate92inter8));
  nand2 gate2894(.a(gate92inter8), .b(gate92inter7), .O(gate92inter9));
  nand2 gate2895(.a(s_335), .b(gate92inter3), .O(gate92inter10));
  nor2  gate2896(.a(gate92inter10), .b(gate92inter9), .O(gate92inter11));
  nor2  gate2897(.a(gate92inter11), .b(gate92inter6), .O(gate92inter12));
  nand2 gate2898(.a(gate92inter12), .b(gate92inter1), .O(G413));

  xor2  gate1611(.a(G344), .b(G18), .O(gate93inter0));
  nand2 gate1612(.a(gate93inter0), .b(s_152), .O(gate93inter1));
  and2  gate1613(.a(G344), .b(G18), .O(gate93inter2));
  inv1  gate1614(.a(s_152), .O(gate93inter3));
  inv1  gate1615(.a(s_153), .O(gate93inter4));
  nand2 gate1616(.a(gate93inter4), .b(gate93inter3), .O(gate93inter5));
  nor2  gate1617(.a(gate93inter5), .b(gate93inter2), .O(gate93inter6));
  inv1  gate1618(.a(G18), .O(gate93inter7));
  inv1  gate1619(.a(G344), .O(gate93inter8));
  nand2 gate1620(.a(gate93inter8), .b(gate93inter7), .O(gate93inter9));
  nand2 gate1621(.a(s_153), .b(gate93inter3), .O(gate93inter10));
  nor2  gate1622(.a(gate93inter10), .b(gate93inter9), .O(gate93inter11));
  nor2  gate1623(.a(gate93inter11), .b(gate93inter6), .O(gate93inter12));
  nand2 gate1624(.a(gate93inter12), .b(gate93inter1), .O(G414));
nand2 gate94( .a(G22), .b(G344), .O(G415) );

  xor2  gate2521(.a(G347), .b(G26), .O(gate95inter0));
  nand2 gate2522(.a(gate95inter0), .b(s_282), .O(gate95inter1));
  and2  gate2523(.a(G347), .b(G26), .O(gate95inter2));
  inv1  gate2524(.a(s_282), .O(gate95inter3));
  inv1  gate2525(.a(s_283), .O(gate95inter4));
  nand2 gate2526(.a(gate95inter4), .b(gate95inter3), .O(gate95inter5));
  nor2  gate2527(.a(gate95inter5), .b(gate95inter2), .O(gate95inter6));
  inv1  gate2528(.a(G26), .O(gate95inter7));
  inv1  gate2529(.a(G347), .O(gate95inter8));
  nand2 gate2530(.a(gate95inter8), .b(gate95inter7), .O(gate95inter9));
  nand2 gate2531(.a(s_283), .b(gate95inter3), .O(gate95inter10));
  nor2  gate2532(.a(gate95inter10), .b(gate95inter9), .O(gate95inter11));
  nor2  gate2533(.a(gate95inter11), .b(gate95inter6), .O(gate95inter12));
  nand2 gate2534(.a(gate95inter12), .b(gate95inter1), .O(G416));
nand2 gate96( .a(G30), .b(G347), .O(G417) );

  xor2  gate2353(.a(G350), .b(G19), .O(gate97inter0));
  nand2 gate2354(.a(gate97inter0), .b(s_258), .O(gate97inter1));
  and2  gate2355(.a(G350), .b(G19), .O(gate97inter2));
  inv1  gate2356(.a(s_258), .O(gate97inter3));
  inv1  gate2357(.a(s_259), .O(gate97inter4));
  nand2 gate2358(.a(gate97inter4), .b(gate97inter3), .O(gate97inter5));
  nor2  gate2359(.a(gate97inter5), .b(gate97inter2), .O(gate97inter6));
  inv1  gate2360(.a(G19), .O(gate97inter7));
  inv1  gate2361(.a(G350), .O(gate97inter8));
  nand2 gate2362(.a(gate97inter8), .b(gate97inter7), .O(gate97inter9));
  nand2 gate2363(.a(s_259), .b(gate97inter3), .O(gate97inter10));
  nor2  gate2364(.a(gate97inter10), .b(gate97inter9), .O(gate97inter11));
  nor2  gate2365(.a(gate97inter11), .b(gate97inter6), .O(gate97inter12));
  nand2 gate2366(.a(gate97inter12), .b(gate97inter1), .O(G418));

  xor2  gate1051(.a(G350), .b(G23), .O(gate98inter0));
  nand2 gate1052(.a(gate98inter0), .b(s_72), .O(gate98inter1));
  and2  gate1053(.a(G350), .b(G23), .O(gate98inter2));
  inv1  gate1054(.a(s_72), .O(gate98inter3));
  inv1  gate1055(.a(s_73), .O(gate98inter4));
  nand2 gate1056(.a(gate98inter4), .b(gate98inter3), .O(gate98inter5));
  nor2  gate1057(.a(gate98inter5), .b(gate98inter2), .O(gate98inter6));
  inv1  gate1058(.a(G23), .O(gate98inter7));
  inv1  gate1059(.a(G350), .O(gate98inter8));
  nand2 gate1060(.a(gate98inter8), .b(gate98inter7), .O(gate98inter9));
  nand2 gate1061(.a(s_73), .b(gate98inter3), .O(gate98inter10));
  nor2  gate1062(.a(gate98inter10), .b(gate98inter9), .O(gate98inter11));
  nor2  gate1063(.a(gate98inter11), .b(gate98inter6), .O(gate98inter12));
  nand2 gate1064(.a(gate98inter12), .b(gate98inter1), .O(G419));
nand2 gate99( .a(G27), .b(G353), .O(G420) );

  xor2  gate3011(.a(G353), .b(G31), .O(gate100inter0));
  nand2 gate3012(.a(gate100inter0), .b(s_352), .O(gate100inter1));
  and2  gate3013(.a(G353), .b(G31), .O(gate100inter2));
  inv1  gate3014(.a(s_352), .O(gate100inter3));
  inv1  gate3015(.a(s_353), .O(gate100inter4));
  nand2 gate3016(.a(gate100inter4), .b(gate100inter3), .O(gate100inter5));
  nor2  gate3017(.a(gate100inter5), .b(gate100inter2), .O(gate100inter6));
  inv1  gate3018(.a(G31), .O(gate100inter7));
  inv1  gate3019(.a(G353), .O(gate100inter8));
  nand2 gate3020(.a(gate100inter8), .b(gate100inter7), .O(gate100inter9));
  nand2 gate3021(.a(s_353), .b(gate100inter3), .O(gate100inter10));
  nor2  gate3022(.a(gate100inter10), .b(gate100inter9), .O(gate100inter11));
  nor2  gate3023(.a(gate100inter11), .b(gate100inter6), .O(gate100inter12));
  nand2 gate3024(.a(gate100inter12), .b(gate100inter1), .O(G421));
nand2 gate101( .a(G20), .b(G356), .O(G422) );

  xor2  gate2297(.a(G356), .b(G24), .O(gate102inter0));
  nand2 gate2298(.a(gate102inter0), .b(s_250), .O(gate102inter1));
  and2  gate2299(.a(G356), .b(G24), .O(gate102inter2));
  inv1  gate2300(.a(s_250), .O(gate102inter3));
  inv1  gate2301(.a(s_251), .O(gate102inter4));
  nand2 gate2302(.a(gate102inter4), .b(gate102inter3), .O(gate102inter5));
  nor2  gate2303(.a(gate102inter5), .b(gate102inter2), .O(gate102inter6));
  inv1  gate2304(.a(G24), .O(gate102inter7));
  inv1  gate2305(.a(G356), .O(gate102inter8));
  nand2 gate2306(.a(gate102inter8), .b(gate102inter7), .O(gate102inter9));
  nand2 gate2307(.a(s_251), .b(gate102inter3), .O(gate102inter10));
  nor2  gate2308(.a(gate102inter10), .b(gate102inter9), .O(gate102inter11));
  nor2  gate2309(.a(gate102inter11), .b(gate102inter6), .O(gate102inter12));
  nand2 gate2310(.a(gate102inter12), .b(gate102inter1), .O(G423));
nand2 gate103( .a(G28), .b(G359), .O(G424) );

  xor2  gate1513(.a(G359), .b(G32), .O(gate104inter0));
  nand2 gate1514(.a(gate104inter0), .b(s_138), .O(gate104inter1));
  and2  gate1515(.a(G359), .b(G32), .O(gate104inter2));
  inv1  gate1516(.a(s_138), .O(gate104inter3));
  inv1  gate1517(.a(s_139), .O(gate104inter4));
  nand2 gate1518(.a(gate104inter4), .b(gate104inter3), .O(gate104inter5));
  nor2  gate1519(.a(gate104inter5), .b(gate104inter2), .O(gate104inter6));
  inv1  gate1520(.a(G32), .O(gate104inter7));
  inv1  gate1521(.a(G359), .O(gate104inter8));
  nand2 gate1522(.a(gate104inter8), .b(gate104inter7), .O(gate104inter9));
  nand2 gate1523(.a(s_139), .b(gate104inter3), .O(gate104inter10));
  nor2  gate1524(.a(gate104inter10), .b(gate104inter9), .O(gate104inter11));
  nor2  gate1525(.a(gate104inter11), .b(gate104inter6), .O(gate104inter12));
  nand2 gate1526(.a(gate104inter12), .b(gate104inter1), .O(G425));
nand2 gate105( .a(G362), .b(G363), .O(G426) );

  xor2  gate2115(.a(G365), .b(G364), .O(gate106inter0));
  nand2 gate2116(.a(gate106inter0), .b(s_224), .O(gate106inter1));
  and2  gate2117(.a(G365), .b(G364), .O(gate106inter2));
  inv1  gate2118(.a(s_224), .O(gate106inter3));
  inv1  gate2119(.a(s_225), .O(gate106inter4));
  nand2 gate2120(.a(gate106inter4), .b(gate106inter3), .O(gate106inter5));
  nor2  gate2121(.a(gate106inter5), .b(gate106inter2), .O(gate106inter6));
  inv1  gate2122(.a(G364), .O(gate106inter7));
  inv1  gate2123(.a(G365), .O(gate106inter8));
  nand2 gate2124(.a(gate106inter8), .b(gate106inter7), .O(gate106inter9));
  nand2 gate2125(.a(s_225), .b(gate106inter3), .O(gate106inter10));
  nor2  gate2126(.a(gate106inter10), .b(gate106inter9), .O(gate106inter11));
  nor2  gate2127(.a(gate106inter11), .b(gate106inter6), .O(gate106inter12));
  nand2 gate2128(.a(gate106inter12), .b(gate106inter1), .O(G429));
nand2 gate107( .a(G366), .b(G367), .O(G432) );
nand2 gate108( .a(G368), .b(G369), .O(G435) );
nand2 gate109( .a(G370), .b(G371), .O(G438) );

  xor2  gate995(.a(G373), .b(G372), .O(gate110inter0));
  nand2 gate996(.a(gate110inter0), .b(s_64), .O(gate110inter1));
  and2  gate997(.a(G373), .b(G372), .O(gate110inter2));
  inv1  gate998(.a(s_64), .O(gate110inter3));
  inv1  gate999(.a(s_65), .O(gate110inter4));
  nand2 gate1000(.a(gate110inter4), .b(gate110inter3), .O(gate110inter5));
  nor2  gate1001(.a(gate110inter5), .b(gate110inter2), .O(gate110inter6));
  inv1  gate1002(.a(G372), .O(gate110inter7));
  inv1  gate1003(.a(G373), .O(gate110inter8));
  nand2 gate1004(.a(gate110inter8), .b(gate110inter7), .O(gate110inter9));
  nand2 gate1005(.a(s_65), .b(gate110inter3), .O(gate110inter10));
  nor2  gate1006(.a(gate110inter10), .b(gate110inter9), .O(gate110inter11));
  nor2  gate1007(.a(gate110inter11), .b(gate110inter6), .O(gate110inter12));
  nand2 gate1008(.a(gate110inter12), .b(gate110inter1), .O(G441));
nand2 gate111( .a(G374), .b(G375), .O(G444) );
nand2 gate112( .a(G376), .b(G377), .O(G447) );
nand2 gate113( .a(G378), .b(G379), .O(G450) );

  xor2  gate2045(.a(G381), .b(G380), .O(gate114inter0));
  nand2 gate2046(.a(gate114inter0), .b(s_214), .O(gate114inter1));
  and2  gate2047(.a(G381), .b(G380), .O(gate114inter2));
  inv1  gate2048(.a(s_214), .O(gate114inter3));
  inv1  gate2049(.a(s_215), .O(gate114inter4));
  nand2 gate2050(.a(gate114inter4), .b(gate114inter3), .O(gate114inter5));
  nor2  gate2051(.a(gate114inter5), .b(gate114inter2), .O(gate114inter6));
  inv1  gate2052(.a(G380), .O(gate114inter7));
  inv1  gate2053(.a(G381), .O(gate114inter8));
  nand2 gate2054(.a(gate114inter8), .b(gate114inter7), .O(gate114inter9));
  nand2 gate2055(.a(s_215), .b(gate114inter3), .O(gate114inter10));
  nor2  gate2056(.a(gate114inter10), .b(gate114inter9), .O(gate114inter11));
  nor2  gate2057(.a(gate114inter11), .b(gate114inter6), .O(gate114inter12));
  nand2 gate2058(.a(gate114inter12), .b(gate114inter1), .O(G453));
nand2 gate115( .a(G382), .b(G383), .O(G456) );
nand2 gate116( .a(G384), .b(G385), .O(G459) );

  xor2  gate1275(.a(G387), .b(G386), .O(gate117inter0));
  nand2 gate1276(.a(gate117inter0), .b(s_104), .O(gate117inter1));
  and2  gate1277(.a(G387), .b(G386), .O(gate117inter2));
  inv1  gate1278(.a(s_104), .O(gate117inter3));
  inv1  gate1279(.a(s_105), .O(gate117inter4));
  nand2 gate1280(.a(gate117inter4), .b(gate117inter3), .O(gate117inter5));
  nor2  gate1281(.a(gate117inter5), .b(gate117inter2), .O(gate117inter6));
  inv1  gate1282(.a(G386), .O(gate117inter7));
  inv1  gate1283(.a(G387), .O(gate117inter8));
  nand2 gate1284(.a(gate117inter8), .b(gate117inter7), .O(gate117inter9));
  nand2 gate1285(.a(s_105), .b(gate117inter3), .O(gate117inter10));
  nor2  gate1286(.a(gate117inter10), .b(gate117inter9), .O(gate117inter11));
  nor2  gate1287(.a(gate117inter11), .b(gate117inter6), .O(gate117inter12));
  nand2 gate1288(.a(gate117inter12), .b(gate117inter1), .O(G462));
nand2 gate118( .a(G388), .b(G389), .O(G465) );
nand2 gate119( .a(G390), .b(G391), .O(G468) );
nand2 gate120( .a(G392), .b(G393), .O(G471) );

  xor2  gate1037(.a(G395), .b(G394), .O(gate121inter0));
  nand2 gate1038(.a(gate121inter0), .b(s_70), .O(gate121inter1));
  and2  gate1039(.a(G395), .b(G394), .O(gate121inter2));
  inv1  gate1040(.a(s_70), .O(gate121inter3));
  inv1  gate1041(.a(s_71), .O(gate121inter4));
  nand2 gate1042(.a(gate121inter4), .b(gate121inter3), .O(gate121inter5));
  nor2  gate1043(.a(gate121inter5), .b(gate121inter2), .O(gate121inter6));
  inv1  gate1044(.a(G394), .O(gate121inter7));
  inv1  gate1045(.a(G395), .O(gate121inter8));
  nand2 gate1046(.a(gate121inter8), .b(gate121inter7), .O(gate121inter9));
  nand2 gate1047(.a(s_71), .b(gate121inter3), .O(gate121inter10));
  nor2  gate1048(.a(gate121inter10), .b(gate121inter9), .O(gate121inter11));
  nor2  gate1049(.a(gate121inter11), .b(gate121inter6), .O(gate121inter12));
  nand2 gate1050(.a(gate121inter12), .b(gate121inter1), .O(G474));
nand2 gate122( .a(G396), .b(G397), .O(G477) );

  xor2  gate631(.a(G399), .b(G398), .O(gate123inter0));
  nand2 gate632(.a(gate123inter0), .b(s_12), .O(gate123inter1));
  and2  gate633(.a(G399), .b(G398), .O(gate123inter2));
  inv1  gate634(.a(s_12), .O(gate123inter3));
  inv1  gate635(.a(s_13), .O(gate123inter4));
  nand2 gate636(.a(gate123inter4), .b(gate123inter3), .O(gate123inter5));
  nor2  gate637(.a(gate123inter5), .b(gate123inter2), .O(gate123inter6));
  inv1  gate638(.a(G398), .O(gate123inter7));
  inv1  gate639(.a(G399), .O(gate123inter8));
  nand2 gate640(.a(gate123inter8), .b(gate123inter7), .O(gate123inter9));
  nand2 gate641(.a(s_13), .b(gate123inter3), .O(gate123inter10));
  nor2  gate642(.a(gate123inter10), .b(gate123inter9), .O(gate123inter11));
  nor2  gate643(.a(gate123inter11), .b(gate123inter6), .O(gate123inter12));
  nand2 gate644(.a(gate123inter12), .b(gate123inter1), .O(G480));
nand2 gate124( .a(G400), .b(G401), .O(G483) );
nand2 gate125( .a(G402), .b(G403), .O(G486) );
nand2 gate126( .a(G404), .b(G405), .O(G489) );

  xor2  gate2689(.a(G407), .b(G406), .O(gate127inter0));
  nand2 gate2690(.a(gate127inter0), .b(s_306), .O(gate127inter1));
  and2  gate2691(.a(G407), .b(G406), .O(gate127inter2));
  inv1  gate2692(.a(s_306), .O(gate127inter3));
  inv1  gate2693(.a(s_307), .O(gate127inter4));
  nand2 gate2694(.a(gate127inter4), .b(gate127inter3), .O(gate127inter5));
  nor2  gate2695(.a(gate127inter5), .b(gate127inter2), .O(gate127inter6));
  inv1  gate2696(.a(G406), .O(gate127inter7));
  inv1  gate2697(.a(G407), .O(gate127inter8));
  nand2 gate2698(.a(gate127inter8), .b(gate127inter7), .O(gate127inter9));
  nand2 gate2699(.a(s_307), .b(gate127inter3), .O(gate127inter10));
  nor2  gate2700(.a(gate127inter10), .b(gate127inter9), .O(gate127inter11));
  nor2  gate2701(.a(gate127inter11), .b(gate127inter6), .O(gate127inter12));
  nand2 gate2702(.a(gate127inter12), .b(gate127inter1), .O(G492));
nand2 gate128( .a(G408), .b(G409), .O(G495) );
nand2 gate129( .a(G410), .b(G411), .O(G498) );

  xor2  gate2381(.a(G413), .b(G412), .O(gate130inter0));
  nand2 gate2382(.a(gate130inter0), .b(s_262), .O(gate130inter1));
  and2  gate2383(.a(G413), .b(G412), .O(gate130inter2));
  inv1  gate2384(.a(s_262), .O(gate130inter3));
  inv1  gate2385(.a(s_263), .O(gate130inter4));
  nand2 gate2386(.a(gate130inter4), .b(gate130inter3), .O(gate130inter5));
  nor2  gate2387(.a(gate130inter5), .b(gate130inter2), .O(gate130inter6));
  inv1  gate2388(.a(G412), .O(gate130inter7));
  inv1  gate2389(.a(G413), .O(gate130inter8));
  nand2 gate2390(.a(gate130inter8), .b(gate130inter7), .O(gate130inter9));
  nand2 gate2391(.a(s_263), .b(gate130inter3), .O(gate130inter10));
  nor2  gate2392(.a(gate130inter10), .b(gate130inter9), .O(gate130inter11));
  nor2  gate2393(.a(gate130inter11), .b(gate130inter6), .O(gate130inter12));
  nand2 gate2394(.a(gate130inter12), .b(gate130inter1), .O(G501));
nand2 gate131( .a(G414), .b(G415), .O(G504) );

  xor2  gate1947(.a(G417), .b(G416), .O(gate132inter0));
  nand2 gate1948(.a(gate132inter0), .b(s_200), .O(gate132inter1));
  and2  gate1949(.a(G417), .b(G416), .O(gate132inter2));
  inv1  gate1950(.a(s_200), .O(gate132inter3));
  inv1  gate1951(.a(s_201), .O(gate132inter4));
  nand2 gate1952(.a(gate132inter4), .b(gate132inter3), .O(gate132inter5));
  nor2  gate1953(.a(gate132inter5), .b(gate132inter2), .O(gate132inter6));
  inv1  gate1954(.a(G416), .O(gate132inter7));
  inv1  gate1955(.a(G417), .O(gate132inter8));
  nand2 gate1956(.a(gate132inter8), .b(gate132inter7), .O(gate132inter9));
  nand2 gate1957(.a(s_201), .b(gate132inter3), .O(gate132inter10));
  nor2  gate1958(.a(gate132inter10), .b(gate132inter9), .O(gate132inter11));
  nor2  gate1959(.a(gate132inter11), .b(gate132inter6), .O(gate132inter12));
  nand2 gate1960(.a(gate132inter12), .b(gate132inter1), .O(G507));

  xor2  gate2591(.a(G419), .b(G418), .O(gate133inter0));
  nand2 gate2592(.a(gate133inter0), .b(s_292), .O(gate133inter1));
  and2  gate2593(.a(G419), .b(G418), .O(gate133inter2));
  inv1  gate2594(.a(s_292), .O(gate133inter3));
  inv1  gate2595(.a(s_293), .O(gate133inter4));
  nand2 gate2596(.a(gate133inter4), .b(gate133inter3), .O(gate133inter5));
  nor2  gate2597(.a(gate133inter5), .b(gate133inter2), .O(gate133inter6));
  inv1  gate2598(.a(G418), .O(gate133inter7));
  inv1  gate2599(.a(G419), .O(gate133inter8));
  nand2 gate2600(.a(gate133inter8), .b(gate133inter7), .O(gate133inter9));
  nand2 gate2601(.a(s_293), .b(gate133inter3), .O(gate133inter10));
  nor2  gate2602(.a(gate133inter10), .b(gate133inter9), .O(gate133inter11));
  nor2  gate2603(.a(gate133inter11), .b(gate133inter6), .O(gate133inter12));
  nand2 gate2604(.a(gate133inter12), .b(gate133inter1), .O(G510));

  xor2  gate3039(.a(G421), .b(G420), .O(gate134inter0));
  nand2 gate3040(.a(gate134inter0), .b(s_356), .O(gate134inter1));
  and2  gate3041(.a(G421), .b(G420), .O(gate134inter2));
  inv1  gate3042(.a(s_356), .O(gate134inter3));
  inv1  gate3043(.a(s_357), .O(gate134inter4));
  nand2 gate3044(.a(gate134inter4), .b(gate134inter3), .O(gate134inter5));
  nor2  gate3045(.a(gate134inter5), .b(gate134inter2), .O(gate134inter6));
  inv1  gate3046(.a(G420), .O(gate134inter7));
  inv1  gate3047(.a(G421), .O(gate134inter8));
  nand2 gate3048(.a(gate134inter8), .b(gate134inter7), .O(gate134inter9));
  nand2 gate3049(.a(s_357), .b(gate134inter3), .O(gate134inter10));
  nor2  gate3050(.a(gate134inter10), .b(gate134inter9), .O(gate134inter11));
  nor2  gate3051(.a(gate134inter11), .b(gate134inter6), .O(gate134inter12));
  nand2 gate3052(.a(gate134inter12), .b(gate134inter1), .O(G513));
nand2 gate135( .a(G422), .b(G423), .O(G516) );

  xor2  gate2171(.a(G425), .b(G424), .O(gate136inter0));
  nand2 gate2172(.a(gate136inter0), .b(s_232), .O(gate136inter1));
  and2  gate2173(.a(G425), .b(G424), .O(gate136inter2));
  inv1  gate2174(.a(s_232), .O(gate136inter3));
  inv1  gate2175(.a(s_233), .O(gate136inter4));
  nand2 gate2176(.a(gate136inter4), .b(gate136inter3), .O(gate136inter5));
  nor2  gate2177(.a(gate136inter5), .b(gate136inter2), .O(gate136inter6));
  inv1  gate2178(.a(G424), .O(gate136inter7));
  inv1  gate2179(.a(G425), .O(gate136inter8));
  nand2 gate2180(.a(gate136inter8), .b(gate136inter7), .O(gate136inter9));
  nand2 gate2181(.a(s_233), .b(gate136inter3), .O(gate136inter10));
  nor2  gate2182(.a(gate136inter10), .b(gate136inter9), .O(gate136inter11));
  nor2  gate2183(.a(gate136inter11), .b(gate136inter6), .O(gate136inter12));
  nand2 gate2184(.a(gate136inter12), .b(gate136inter1), .O(G519));
nand2 gate137( .a(G426), .b(G429), .O(G522) );

  xor2  gate1261(.a(G435), .b(G432), .O(gate138inter0));
  nand2 gate1262(.a(gate138inter0), .b(s_102), .O(gate138inter1));
  and2  gate1263(.a(G435), .b(G432), .O(gate138inter2));
  inv1  gate1264(.a(s_102), .O(gate138inter3));
  inv1  gate1265(.a(s_103), .O(gate138inter4));
  nand2 gate1266(.a(gate138inter4), .b(gate138inter3), .O(gate138inter5));
  nor2  gate1267(.a(gate138inter5), .b(gate138inter2), .O(gate138inter6));
  inv1  gate1268(.a(G432), .O(gate138inter7));
  inv1  gate1269(.a(G435), .O(gate138inter8));
  nand2 gate1270(.a(gate138inter8), .b(gate138inter7), .O(gate138inter9));
  nand2 gate1271(.a(s_103), .b(gate138inter3), .O(gate138inter10));
  nor2  gate1272(.a(gate138inter10), .b(gate138inter9), .O(gate138inter11));
  nor2  gate1273(.a(gate138inter11), .b(gate138inter6), .O(gate138inter12));
  nand2 gate1274(.a(gate138inter12), .b(gate138inter1), .O(G525));

  xor2  gate2059(.a(G441), .b(G438), .O(gate139inter0));
  nand2 gate2060(.a(gate139inter0), .b(s_216), .O(gate139inter1));
  and2  gate2061(.a(G441), .b(G438), .O(gate139inter2));
  inv1  gate2062(.a(s_216), .O(gate139inter3));
  inv1  gate2063(.a(s_217), .O(gate139inter4));
  nand2 gate2064(.a(gate139inter4), .b(gate139inter3), .O(gate139inter5));
  nor2  gate2065(.a(gate139inter5), .b(gate139inter2), .O(gate139inter6));
  inv1  gate2066(.a(G438), .O(gate139inter7));
  inv1  gate2067(.a(G441), .O(gate139inter8));
  nand2 gate2068(.a(gate139inter8), .b(gate139inter7), .O(gate139inter9));
  nand2 gate2069(.a(s_217), .b(gate139inter3), .O(gate139inter10));
  nor2  gate2070(.a(gate139inter10), .b(gate139inter9), .O(gate139inter11));
  nor2  gate2071(.a(gate139inter11), .b(gate139inter6), .O(gate139inter12));
  nand2 gate2072(.a(gate139inter12), .b(gate139inter1), .O(G528));
nand2 gate140( .a(G444), .b(G447), .O(G531) );

  xor2  gate2577(.a(G453), .b(G450), .O(gate141inter0));
  nand2 gate2578(.a(gate141inter0), .b(s_290), .O(gate141inter1));
  and2  gate2579(.a(G453), .b(G450), .O(gate141inter2));
  inv1  gate2580(.a(s_290), .O(gate141inter3));
  inv1  gate2581(.a(s_291), .O(gate141inter4));
  nand2 gate2582(.a(gate141inter4), .b(gate141inter3), .O(gate141inter5));
  nor2  gate2583(.a(gate141inter5), .b(gate141inter2), .O(gate141inter6));
  inv1  gate2584(.a(G450), .O(gate141inter7));
  inv1  gate2585(.a(G453), .O(gate141inter8));
  nand2 gate2586(.a(gate141inter8), .b(gate141inter7), .O(gate141inter9));
  nand2 gate2587(.a(s_291), .b(gate141inter3), .O(gate141inter10));
  nor2  gate2588(.a(gate141inter10), .b(gate141inter9), .O(gate141inter11));
  nor2  gate2589(.a(gate141inter11), .b(gate141inter6), .O(gate141inter12));
  nand2 gate2590(.a(gate141inter12), .b(gate141inter1), .O(G534));
nand2 gate142( .a(G456), .b(G459), .O(G537) );

  xor2  gate1359(.a(G465), .b(G462), .O(gate143inter0));
  nand2 gate1360(.a(gate143inter0), .b(s_116), .O(gate143inter1));
  and2  gate1361(.a(G465), .b(G462), .O(gate143inter2));
  inv1  gate1362(.a(s_116), .O(gate143inter3));
  inv1  gate1363(.a(s_117), .O(gate143inter4));
  nand2 gate1364(.a(gate143inter4), .b(gate143inter3), .O(gate143inter5));
  nor2  gate1365(.a(gate143inter5), .b(gate143inter2), .O(gate143inter6));
  inv1  gate1366(.a(G462), .O(gate143inter7));
  inv1  gate1367(.a(G465), .O(gate143inter8));
  nand2 gate1368(.a(gate143inter8), .b(gate143inter7), .O(gate143inter9));
  nand2 gate1369(.a(s_117), .b(gate143inter3), .O(gate143inter10));
  nor2  gate1370(.a(gate143inter10), .b(gate143inter9), .O(gate143inter11));
  nor2  gate1371(.a(gate143inter11), .b(gate143inter6), .O(gate143inter12));
  nand2 gate1372(.a(gate143inter12), .b(gate143inter1), .O(G540));
nand2 gate144( .a(G468), .b(G471), .O(G543) );
nand2 gate145( .a(G474), .b(G477), .O(G546) );

  xor2  gate1471(.a(G483), .b(G480), .O(gate146inter0));
  nand2 gate1472(.a(gate146inter0), .b(s_132), .O(gate146inter1));
  and2  gate1473(.a(G483), .b(G480), .O(gate146inter2));
  inv1  gate1474(.a(s_132), .O(gate146inter3));
  inv1  gate1475(.a(s_133), .O(gate146inter4));
  nand2 gate1476(.a(gate146inter4), .b(gate146inter3), .O(gate146inter5));
  nor2  gate1477(.a(gate146inter5), .b(gate146inter2), .O(gate146inter6));
  inv1  gate1478(.a(G480), .O(gate146inter7));
  inv1  gate1479(.a(G483), .O(gate146inter8));
  nand2 gate1480(.a(gate146inter8), .b(gate146inter7), .O(gate146inter9));
  nand2 gate1481(.a(s_133), .b(gate146inter3), .O(gate146inter10));
  nor2  gate1482(.a(gate146inter10), .b(gate146inter9), .O(gate146inter11));
  nor2  gate1483(.a(gate146inter11), .b(gate146inter6), .O(gate146inter12));
  nand2 gate1484(.a(gate146inter12), .b(gate146inter1), .O(G549));

  xor2  gate2101(.a(G489), .b(G486), .O(gate147inter0));
  nand2 gate2102(.a(gate147inter0), .b(s_222), .O(gate147inter1));
  and2  gate2103(.a(G489), .b(G486), .O(gate147inter2));
  inv1  gate2104(.a(s_222), .O(gate147inter3));
  inv1  gate2105(.a(s_223), .O(gate147inter4));
  nand2 gate2106(.a(gate147inter4), .b(gate147inter3), .O(gate147inter5));
  nor2  gate2107(.a(gate147inter5), .b(gate147inter2), .O(gate147inter6));
  inv1  gate2108(.a(G486), .O(gate147inter7));
  inv1  gate2109(.a(G489), .O(gate147inter8));
  nand2 gate2110(.a(gate147inter8), .b(gate147inter7), .O(gate147inter9));
  nand2 gate2111(.a(s_223), .b(gate147inter3), .O(gate147inter10));
  nor2  gate2112(.a(gate147inter10), .b(gate147inter9), .O(gate147inter11));
  nor2  gate2113(.a(gate147inter11), .b(gate147inter6), .O(gate147inter12));
  nand2 gate2114(.a(gate147inter12), .b(gate147inter1), .O(G552));

  xor2  gate659(.a(G495), .b(G492), .O(gate148inter0));
  nand2 gate660(.a(gate148inter0), .b(s_16), .O(gate148inter1));
  and2  gate661(.a(G495), .b(G492), .O(gate148inter2));
  inv1  gate662(.a(s_16), .O(gate148inter3));
  inv1  gate663(.a(s_17), .O(gate148inter4));
  nand2 gate664(.a(gate148inter4), .b(gate148inter3), .O(gate148inter5));
  nor2  gate665(.a(gate148inter5), .b(gate148inter2), .O(gate148inter6));
  inv1  gate666(.a(G492), .O(gate148inter7));
  inv1  gate667(.a(G495), .O(gate148inter8));
  nand2 gate668(.a(gate148inter8), .b(gate148inter7), .O(gate148inter9));
  nand2 gate669(.a(s_17), .b(gate148inter3), .O(gate148inter10));
  nor2  gate670(.a(gate148inter10), .b(gate148inter9), .O(gate148inter11));
  nor2  gate671(.a(gate148inter11), .b(gate148inter6), .O(gate148inter12));
  nand2 gate672(.a(gate148inter12), .b(gate148inter1), .O(G555));
nand2 gate149( .a(G498), .b(G501), .O(G558) );

  xor2  gate2465(.a(G507), .b(G504), .O(gate150inter0));
  nand2 gate2466(.a(gate150inter0), .b(s_274), .O(gate150inter1));
  and2  gate2467(.a(G507), .b(G504), .O(gate150inter2));
  inv1  gate2468(.a(s_274), .O(gate150inter3));
  inv1  gate2469(.a(s_275), .O(gate150inter4));
  nand2 gate2470(.a(gate150inter4), .b(gate150inter3), .O(gate150inter5));
  nor2  gate2471(.a(gate150inter5), .b(gate150inter2), .O(gate150inter6));
  inv1  gate2472(.a(G504), .O(gate150inter7));
  inv1  gate2473(.a(G507), .O(gate150inter8));
  nand2 gate2474(.a(gate150inter8), .b(gate150inter7), .O(gate150inter9));
  nand2 gate2475(.a(s_275), .b(gate150inter3), .O(gate150inter10));
  nor2  gate2476(.a(gate150inter10), .b(gate150inter9), .O(gate150inter11));
  nor2  gate2477(.a(gate150inter11), .b(gate150inter6), .O(gate150inter12));
  nand2 gate2478(.a(gate150inter12), .b(gate150inter1), .O(G561));
nand2 gate151( .a(G510), .b(G513), .O(G564) );
nand2 gate152( .a(G516), .b(G519), .O(G567) );

  xor2  gate1121(.a(G522), .b(G426), .O(gate153inter0));
  nand2 gate1122(.a(gate153inter0), .b(s_82), .O(gate153inter1));
  and2  gate1123(.a(G522), .b(G426), .O(gate153inter2));
  inv1  gate1124(.a(s_82), .O(gate153inter3));
  inv1  gate1125(.a(s_83), .O(gate153inter4));
  nand2 gate1126(.a(gate153inter4), .b(gate153inter3), .O(gate153inter5));
  nor2  gate1127(.a(gate153inter5), .b(gate153inter2), .O(gate153inter6));
  inv1  gate1128(.a(G426), .O(gate153inter7));
  inv1  gate1129(.a(G522), .O(gate153inter8));
  nand2 gate1130(.a(gate153inter8), .b(gate153inter7), .O(gate153inter9));
  nand2 gate1131(.a(s_83), .b(gate153inter3), .O(gate153inter10));
  nor2  gate1132(.a(gate153inter10), .b(gate153inter9), .O(gate153inter11));
  nor2  gate1133(.a(gate153inter11), .b(gate153inter6), .O(gate153inter12));
  nand2 gate1134(.a(gate153inter12), .b(gate153inter1), .O(G570));

  xor2  gate2283(.a(G522), .b(G429), .O(gate154inter0));
  nand2 gate2284(.a(gate154inter0), .b(s_248), .O(gate154inter1));
  and2  gate2285(.a(G522), .b(G429), .O(gate154inter2));
  inv1  gate2286(.a(s_248), .O(gate154inter3));
  inv1  gate2287(.a(s_249), .O(gate154inter4));
  nand2 gate2288(.a(gate154inter4), .b(gate154inter3), .O(gate154inter5));
  nor2  gate2289(.a(gate154inter5), .b(gate154inter2), .O(gate154inter6));
  inv1  gate2290(.a(G429), .O(gate154inter7));
  inv1  gate2291(.a(G522), .O(gate154inter8));
  nand2 gate2292(.a(gate154inter8), .b(gate154inter7), .O(gate154inter9));
  nand2 gate2293(.a(s_249), .b(gate154inter3), .O(gate154inter10));
  nor2  gate2294(.a(gate154inter10), .b(gate154inter9), .O(gate154inter11));
  nor2  gate2295(.a(gate154inter11), .b(gate154inter6), .O(gate154inter12));
  nand2 gate2296(.a(gate154inter12), .b(gate154inter1), .O(G571));

  xor2  gate1751(.a(G525), .b(G432), .O(gate155inter0));
  nand2 gate1752(.a(gate155inter0), .b(s_172), .O(gate155inter1));
  and2  gate1753(.a(G525), .b(G432), .O(gate155inter2));
  inv1  gate1754(.a(s_172), .O(gate155inter3));
  inv1  gate1755(.a(s_173), .O(gate155inter4));
  nand2 gate1756(.a(gate155inter4), .b(gate155inter3), .O(gate155inter5));
  nor2  gate1757(.a(gate155inter5), .b(gate155inter2), .O(gate155inter6));
  inv1  gate1758(.a(G432), .O(gate155inter7));
  inv1  gate1759(.a(G525), .O(gate155inter8));
  nand2 gate1760(.a(gate155inter8), .b(gate155inter7), .O(gate155inter9));
  nand2 gate1761(.a(s_173), .b(gate155inter3), .O(gate155inter10));
  nor2  gate1762(.a(gate155inter10), .b(gate155inter9), .O(gate155inter11));
  nor2  gate1763(.a(gate155inter11), .b(gate155inter6), .O(gate155inter12));
  nand2 gate1764(.a(gate155inter12), .b(gate155inter1), .O(G572));
nand2 gate156( .a(G435), .b(G525), .O(G573) );

  xor2  gate2619(.a(G528), .b(G438), .O(gate157inter0));
  nand2 gate2620(.a(gate157inter0), .b(s_296), .O(gate157inter1));
  and2  gate2621(.a(G528), .b(G438), .O(gate157inter2));
  inv1  gate2622(.a(s_296), .O(gate157inter3));
  inv1  gate2623(.a(s_297), .O(gate157inter4));
  nand2 gate2624(.a(gate157inter4), .b(gate157inter3), .O(gate157inter5));
  nor2  gate2625(.a(gate157inter5), .b(gate157inter2), .O(gate157inter6));
  inv1  gate2626(.a(G438), .O(gate157inter7));
  inv1  gate2627(.a(G528), .O(gate157inter8));
  nand2 gate2628(.a(gate157inter8), .b(gate157inter7), .O(gate157inter9));
  nand2 gate2629(.a(s_297), .b(gate157inter3), .O(gate157inter10));
  nor2  gate2630(.a(gate157inter10), .b(gate157inter9), .O(gate157inter11));
  nor2  gate2631(.a(gate157inter11), .b(gate157inter6), .O(gate157inter12));
  nand2 gate2632(.a(gate157inter12), .b(gate157inter1), .O(G574));
nand2 gate158( .a(G441), .b(G528), .O(G575) );
nand2 gate159( .a(G444), .b(G531), .O(G576) );
nand2 gate160( .a(G447), .b(G531), .O(G577) );

  xor2  gate2451(.a(G534), .b(G450), .O(gate161inter0));
  nand2 gate2452(.a(gate161inter0), .b(s_272), .O(gate161inter1));
  and2  gate2453(.a(G534), .b(G450), .O(gate161inter2));
  inv1  gate2454(.a(s_272), .O(gate161inter3));
  inv1  gate2455(.a(s_273), .O(gate161inter4));
  nand2 gate2456(.a(gate161inter4), .b(gate161inter3), .O(gate161inter5));
  nor2  gate2457(.a(gate161inter5), .b(gate161inter2), .O(gate161inter6));
  inv1  gate2458(.a(G450), .O(gate161inter7));
  inv1  gate2459(.a(G534), .O(gate161inter8));
  nand2 gate2460(.a(gate161inter8), .b(gate161inter7), .O(gate161inter9));
  nand2 gate2461(.a(s_273), .b(gate161inter3), .O(gate161inter10));
  nor2  gate2462(.a(gate161inter10), .b(gate161inter9), .O(gate161inter11));
  nor2  gate2463(.a(gate161inter11), .b(gate161inter6), .O(gate161inter12));
  nand2 gate2464(.a(gate161inter12), .b(gate161inter1), .O(G578));
nand2 gate162( .a(G453), .b(G534), .O(G579) );
nand2 gate163( .a(G456), .b(G537), .O(G580) );
nand2 gate164( .a(G459), .b(G537), .O(G581) );
nand2 gate165( .a(G462), .b(G540), .O(G582) );

  xor2  gate1821(.a(G540), .b(G465), .O(gate166inter0));
  nand2 gate1822(.a(gate166inter0), .b(s_182), .O(gate166inter1));
  and2  gate1823(.a(G540), .b(G465), .O(gate166inter2));
  inv1  gate1824(.a(s_182), .O(gate166inter3));
  inv1  gate1825(.a(s_183), .O(gate166inter4));
  nand2 gate1826(.a(gate166inter4), .b(gate166inter3), .O(gate166inter5));
  nor2  gate1827(.a(gate166inter5), .b(gate166inter2), .O(gate166inter6));
  inv1  gate1828(.a(G465), .O(gate166inter7));
  inv1  gate1829(.a(G540), .O(gate166inter8));
  nand2 gate1830(.a(gate166inter8), .b(gate166inter7), .O(gate166inter9));
  nand2 gate1831(.a(s_183), .b(gate166inter3), .O(gate166inter10));
  nor2  gate1832(.a(gate166inter10), .b(gate166inter9), .O(gate166inter11));
  nor2  gate1833(.a(gate166inter11), .b(gate166inter6), .O(gate166inter12));
  nand2 gate1834(.a(gate166inter12), .b(gate166inter1), .O(G583));

  xor2  gate3081(.a(G543), .b(G468), .O(gate167inter0));
  nand2 gate3082(.a(gate167inter0), .b(s_362), .O(gate167inter1));
  and2  gate3083(.a(G543), .b(G468), .O(gate167inter2));
  inv1  gate3084(.a(s_362), .O(gate167inter3));
  inv1  gate3085(.a(s_363), .O(gate167inter4));
  nand2 gate3086(.a(gate167inter4), .b(gate167inter3), .O(gate167inter5));
  nor2  gate3087(.a(gate167inter5), .b(gate167inter2), .O(gate167inter6));
  inv1  gate3088(.a(G468), .O(gate167inter7));
  inv1  gate3089(.a(G543), .O(gate167inter8));
  nand2 gate3090(.a(gate167inter8), .b(gate167inter7), .O(gate167inter9));
  nand2 gate3091(.a(s_363), .b(gate167inter3), .O(gate167inter10));
  nor2  gate3092(.a(gate167inter10), .b(gate167inter9), .O(gate167inter11));
  nor2  gate3093(.a(gate167inter11), .b(gate167inter6), .O(gate167inter12));
  nand2 gate3094(.a(gate167inter12), .b(gate167inter1), .O(G584));

  xor2  gate785(.a(G543), .b(G471), .O(gate168inter0));
  nand2 gate786(.a(gate168inter0), .b(s_34), .O(gate168inter1));
  and2  gate787(.a(G543), .b(G471), .O(gate168inter2));
  inv1  gate788(.a(s_34), .O(gate168inter3));
  inv1  gate789(.a(s_35), .O(gate168inter4));
  nand2 gate790(.a(gate168inter4), .b(gate168inter3), .O(gate168inter5));
  nor2  gate791(.a(gate168inter5), .b(gate168inter2), .O(gate168inter6));
  inv1  gate792(.a(G471), .O(gate168inter7));
  inv1  gate793(.a(G543), .O(gate168inter8));
  nand2 gate794(.a(gate168inter8), .b(gate168inter7), .O(gate168inter9));
  nand2 gate795(.a(s_35), .b(gate168inter3), .O(gate168inter10));
  nor2  gate796(.a(gate168inter10), .b(gate168inter9), .O(gate168inter11));
  nor2  gate797(.a(gate168inter11), .b(gate168inter6), .O(gate168inter12));
  nand2 gate798(.a(gate168inter12), .b(gate168inter1), .O(G585));

  xor2  gate953(.a(G546), .b(G474), .O(gate169inter0));
  nand2 gate954(.a(gate169inter0), .b(s_58), .O(gate169inter1));
  and2  gate955(.a(G546), .b(G474), .O(gate169inter2));
  inv1  gate956(.a(s_58), .O(gate169inter3));
  inv1  gate957(.a(s_59), .O(gate169inter4));
  nand2 gate958(.a(gate169inter4), .b(gate169inter3), .O(gate169inter5));
  nor2  gate959(.a(gate169inter5), .b(gate169inter2), .O(gate169inter6));
  inv1  gate960(.a(G474), .O(gate169inter7));
  inv1  gate961(.a(G546), .O(gate169inter8));
  nand2 gate962(.a(gate169inter8), .b(gate169inter7), .O(gate169inter9));
  nand2 gate963(.a(s_59), .b(gate169inter3), .O(gate169inter10));
  nor2  gate964(.a(gate169inter10), .b(gate169inter9), .O(gate169inter11));
  nor2  gate965(.a(gate169inter11), .b(gate169inter6), .O(gate169inter12));
  nand2 gate966(.a(gate169inter12), .b(gate169inter1), .O(G586));

  xor2  gate2311(.a(G546), .b(G477), .O(gate170inter0));
  nand2 gate2312(.a(gate170inter0), .b(s_252), .O(gate170inter1));
  and2  gate2313(.a(G546), .b(G477), .O(gate170inter2));
  inv1  gate2314(.a(s_252), .O(gate170inter3));
  inv1  gate2315(.a(s_253), .O(gate170inter4));
  nand2 gate2316(.a(gate170inter4), .b(gate170inter3), .O(gate170inter5));
  nor2  gate2317(.a(gate170inter5), .b(gate170inter2), .O(gate170inter6));
  inv1  gate2318(.a(G477), .O(gate170inter7));
  inv1  gate2319(.a(G546), .O(gate170inter8));
  nand2 gate2320(.a(gate170inter8), .b(gate170inter7), .O(gate170inter9));
  nand2 gate2321(.a(s_253), .b(gate170inter3), .O(gate170inter10));
  nor2  gate2322(.a(gate170inter10), .b(gate170inter9), .O(gate170inter11));
  nor2  gate2323(.a(gate170inter11), .b(gate170inter6), .O(gate170inter12));
  nand2 gate2324(.a(gate170inter12), .b(gate170inter1), .O(G587));

  xor2  gate1835(.a(G549), .b(G480), .O(gate171inter0));
  nand2 gate1836(.a(gate171inter0), .b(s_184), .O(gate171inter1));
  and2  gate1837(.a(G549), .b(G480), .O(gate171inter2));
  inv1  gate1838(.a(s_184), .O(gate171inter3));
  inv1  gate1839(.a(s_185), .O(gate171inter4));
  nand2 gate1840(.a(gate171inter4), .b(gate171inter3), .O(gate171inter5));
  nor2  gate1841(.a(gate171inter5), .b(gate171inter2), .O(gate171inter6));
  inv1  gate1842(.a(G480), .O(gate171inter7));
  inv1  gate1843(.a(G549), .O(gate171inter8));
  nand2 gate1844(.a(gate171inter8), .b(gate171inter7), .O(gate171inter9));
  nand2 gate1845(.a(s_185), .b(gate171inter3), .O(gate171inter10));
  nor2  gate1846(.a(gate171inter10), .b(gate171inter9), .O(gate171inter11));
  nor2  gate1847(.a(gate171inter11), .b(gate171inter6), .O(gate171inter12));
  nand2 gate1848(.a(gate171inter12), .b(gate171inter1), .O(G588));
nand2 gate172( .a(G483), .b(G549), .O(G589) );

  xor2  gate687(.a(G552), .b(G486), .O(gate173inter0));
  nand2 gate688(.a(gate173inter0), .b(s_20), .O(gate173inter1));
  and2  gate689(.a(G552), .b(G486), .O(gate173inter2));
  inv1  gate690(.a(s_20), .O(gate173inter3));
  inv1  gate691(.a(s_21), .O(gate173inter4));
  nand2 gate692(.a(gate173inter4), .b(gate173inter3), .O(gate173inter5));
  nor2  gate693(.a(gate173inter5), .b(gate173inter2), .O(gate173inter6));
  inv1  gate694(.a(G486), .O(gate173inter7));
  inv1  gate695(.a(G552), .O(gate173inter8));
  nand2 gate696(.a(gate173inter8), .b(gate173inter7), .O(gate173inter9));
  nand2 gate697(.a(s_21), .b(gate173inter3), .O(gate173inter10));
  nor2  gate698(.a(gate173inter10), .b(gate173inter9), .O(gate173inter11));
  nor2  gate699(.a(gate173inter11), .b(gate173inter6), .O(gate173inter12));
  nand2 gate700(.a(gate173inter12), .b(gate173inter1), .O(G590));
nand2 gate174( .a(G489), .b(G552), .O(G591) );

  xor2  gate3137(.a(G555), .b(G492), .O(gate175inter0));
  nand2 gate3138(.a(gate175inter0), .b(s_370), .O(gate175inter1));
  and2  gate3139(.a(G555), .b(G492), .O(gate175inter2));
  inv1  gate3140(.a(s_370), .O(gate175inter3));
  inv1  gate3141(.a(s_371), .O(gate175inter4));
  nand2 gate3142(.a(gate175inter4), .b(gate175inter3), .O(gate175inter5));
  nor2  gate3143(.a(gate175inter5), .b(gate175inter2), .O(gate175inter6));
  inv1  gate3144(.a(G492), .O(gate175inter7));
  inv1  gate3145(.a(G555), .O(gate175inter8));
  nand2 gate3146(.a(gate175inter8), .b(gate175inter7), .O(gate175inter9));
  nand2 gate3147(.a(s_371), .b(gate175inter3), .O(gate175inter10));
  nor2  gate3148(.a(gate175inter10), .b(gate175inter9), .O(gate175inter11));
  nor2  gate3149(.a(gate175inter11), .b(gate175inter6), .O(gate175inter12));
  nand2 gate3150(.a(gate175inter12), .b(gate175inter1), .O(G592));

  xor2  gate3109(.a(G555), .b(G495), .O(gate176inter0));
  nand2 gate3110(.a(gate176inter0), .b(s_366), .O(gate176inter1));
  and2  gate3111(.a(G555), .b(G495), .O(gate176inter2));
  inv1  gate3112(.a(s_366), .O(gate176inter3));
  inv1  gate3113(.a(s_367), .O(gate176inter4));
  nand2 gate3114(.a(gate176inter4), .b(gate176inter3), .O(gate176inter5));
  nor2  gate3115(.a(gate176inter5), .b(gate176inter2), .O(gate176inter6));
  inv1  gate3116(.a(G495), .O(gate176inter7));
  inv1  gate3117(.a(G555), .O(gate176inter8));
  nand2 gate3118(.a(gate176inter8), .b(gate176inter7), .O(gate176inter9));
  nand2 gate3119(.a(s_367), .b(gate176inter3), .O(gate176inter10));
  nor2  gate3120(.a(gate176inter10), .b(gate176inter9), .O(gate176inter11));
  nor2  gate3121(.a(gate176inter11), .b(gate176inter6), .O(gate176inter12));
  nand2 gate3122(.a(gate176inter12), .b(gate176inter1), .O(G593));
nand2 gate177( .a(G498), .b(G558), .O(G594) );
nand2 gate178( .a(G501), .b(G558), .O(G595) );
nand2 gate179( .a(G504), .b(G561), .O(G596) );
nand2 gate180( .a(G507), .b(G561), .O(G597) );
nand2 gate181( .a(G510), .b(G564), .O(G598) );
nand2 gate182( .a(G513), .b(G564), .O(G599) );

  xor2  gate827(.a(G567), .b(G516), .O(gate183inter0));
  nand2 gate828(.a(gate183inter0), .b(s_40), .O(gate183inter1));
  and2  gate829(.a(G567), .b(G516), .O(gate183inter2));
  inv1  gate830(.a(s_40), .O(gate183inter3));
  inv1  gate831(.a(s_41), .O(gate183inter4));
  nand2 gate832(.a(gate183inter4), .b(gate183inter3), .O(gate183inter5));
  nor2  gate833(.a(gate183inter5), .b(gate183inter2), .O(gate183inter6));
  inv1  gate834(.a(G516), .O(gate183inter7));
  inv1  gate835(.a(G567), .O(gate183inter8));
  nand2 gate836(.a(gate183inter8), .b(gate183inter7), .O(gate183inter9));
  nand2 gate837(.a(s_41), .b(gate183inter3), .O(gate183inter10));
  nor2  gate838(.a(gate183inter10), .b(gate183inter9), .O(gate183inter11));
  nor2  gate839(.a(gate183inter11), .b(gate183inter6), .O(gate183inter12));
  nand2 gate840(.a(gate183inter12), .b(gate183inter1), .O(G600));
nand2 gate184( .a(G519), .b(G567), .O(G601) );
nand2 gate185( .a(G570), .b(G571), .O(G602) );
nand2 gate186( .a(G572), .b(G573), .O(G607) );

  xor2  gate2227(.a(G575), .b(G574), .O(gate187inter0));
  nand2 gate2228(.a(gate187inter0), .b(s_240), .O(gate187inter1));
  and2  gate2229(.a(G575), .b(G574), .O(gate187inter2));
  inv1  gate2230(.a(s_240), .O(gate187inter3));
  inv1  gate2231(.a(s_241), .O(gate187inter4));
  nand2 gate2232(.a(gate187inter4), .b(gate187inter3), .O(gate187inter5));
  nor2  gate2233(.a(gate187inter5), .b(gate187inter2), .O(gate187inter6));
  inv1  gate2234(.a(G574), .O(gate187inter7));
  inv1  gate2235(.a(G575), .O(gate187inter8));
  nand2 gate2236(.a(gate187inter8), .b(gate187inter7), .O(gate187inter9));
  nand2 gate2237(.a(s_241), .b(gate187inter3), .O(gate187inter10));
  nor2  gate2238(.a(gate187inter10), .b(gate187inter9), .O(gate187inter11));
  nor2  gate2239(.a(gate187inter11), .b(gate187inter6), .O(gate187inter12));
  nand2 gate2240(.a(gate187inter12), .b(gate187inter1), .O(G612));

  xor2  gate2185(.a(G577), .b(G576), .O(gate188inter0));
  nand2 gate2186(.a(gate188inter0), .b(s_234), .O(gate188inter1));
  and2  gate2187(.a(G577), .b(G576), .O(gate188inter2));
  inv1  gate2188(.a(s_234), .O(gate188inter3));
  inv1  gate2189(.a(s_235), .O(gate188inter4));
  nand2 gate2190(.a(gate188inter4), .b(gate188inter3), .O(gate188inter5));
  nor2  gate2191(.a(gate188inter5), .b(gate188inter2), .O(gate188inter6));
  inv1  gate2192(.a(G576), .O(gate188inter7));
  inv1  gate2193(.a(G577), .O(gate188inter8));
  nand2 gate2194(.a(gate188inter8), .b(gate188inter7), .O(gate188inter9));
  nand2 gate2195(.a(s_235), .b(gate188inter3), .O(gate188inter10));
  nor2  gate2196(.a(gate188inter10), .b(gate188inter9), .O(gate188inter11));
  nor2  gate2197(.a(gate188inter11), .b(gate188inter6), .O(gate188inter12));
  nand2 gate2198(.a(gate188inter12), .b(gate188inter1), .O(G617));
nand2 gate189( .a(G578), .b(G579), .O(G622) );

  xor2  gate1149(.a(G581), .b(G580), .O(gate190inter0));
  nand2 gate1150(.a(gate190inter0), .b(s_86), .O(gate190inter1));
  and2  gate1151(.a(G581), .b(G580), .O(gate190inter2));
  inv1  gate1152(.a(s_86), .O(gate190inter3));
  inv1  gate1153(.a(s_87), .O(gate190inter4));
  nand2 gate1154(.a(gate190inter4), .b(gate190inter3), .O(gate190inter5));
  nor2  gate1155(.a(gate190inter5), .b(gate190inter2), .O(gate190inter6));
  inv1  gate1156(.a(G580), .O(gate190inter7));
  inv1  gate1157(.a(G581), .O(gate190inter8));
  nand2 gate1158(.a(gate190inter8), .b(gate190inter7), .O(gate190inter9));
  nand2 gate1159(.a(s_87), .b(gate190inter3), .O(gate190inter10));
  nor2  gate1160(.a(gate190inter10), .b(gate190inter9), .O(gate190inter11));
  nor2  gate1161(.a(gate190inter11), .b(gate190inter6), .O(gate190inter12));
  nand2 gate1162(.a(gate190inter12), .b(gate190inter1), .O(G627));

  xor2  gate1205(.a(G583), .b(G582), .O(gate191inter0));
  nand2 gate1206(.a(gate191inter0), .b(s_94), .O(gate191inter1));
  and2  gate1207(.a(G583), .b(G582), .O(gate191inter2));
  inv1  gate1208(.a(s_94), .O(gate191inter3));
  inv1  gate1209(.a(s_95), .O(gate191inter4));
  nand2 gate1210(.a(gate191inter4), .b(gate191inter3), .O(gate191inter5));
  nor2  gate1211(.a(gate191inter5), .b(gate191inter2), .O(gate191inter6));
  inv1  gate1212(.a(G582), .O(gate191inter7));
  inv1  gate1213(.a(G583), .O(gate191inter8));
  nand2 gate1214(.a(gate191inter8), .b(gate191inter7), .O(gate191inter9));
  nand2 gate1215(.a(s_95), .b(gate191inter3), .O(gate191inter10));
  nor2  gate1216(.a(gate191inter10), .b(gate191inter9), .O(gate191inter11));
  nor2  gate1217(.a(gate191inter11), .b(gate191inter6), .O(gate191inter12));
  nand2 gate1218(.a(gate191inter12), .b(gate191inter1), .O(G632));
nand2 gate192( .a(G584), .b(G585), .O(G637) );

  xor2  gate2367(.a(G587), .b(G586), .O(gate193inter0));
  nand2 gate2368(.a(gate193inter0), .b(s_260), .O(gate193inter1));
  and2  gate2369(.a(G587), .b(G586), .O(gate193inter2));
  inv1  gate2370(.a(s_260), .O(gate193inter3));
  inv1  gate2371(.a(s_261), .O(gate193inter4));
  nand2 gate2372(.a(gate193inter4), .b(gate193inter3), .O(gate193inter5));
  nor2  gate2373(.a(gate193inter5), .b(gate193inter2), .O(gate193inter6));
  inv1  gate2374(.a(G586), .O(gate193inter7));
  inv1  gate2375(.a(G587), .O(gate193inter8));
  nand2 gate2376(.a(gate193inter8), .b(gate193inter7), .O(gate193inter9));
  nand2 gate2377(.a(s_261), .b(gate193inter3), .O(gate193inter10));
  nor2  gate2378(.a(gate193inter10), .b(gate193inter9), .O(gate193inter11));
  nor2  gate2379(.a(gate193inter11), .b(gate193inter6), .O(gate193inter12));
  nand2 gate2380(.a(gate193inter12), .b(gate193inter1), .O(G642));

  xor2  gate1443(.a(G589), .b(G588), .O(gate194inter0));
  nand2 gate1444(.a(gate194inter0), .b(s_128), .O(gate194inter1));
  and2  gate1445(.a(G589), .b(G588), .O(gate194inter2));
  inv1  gate1446(.a(s_128), .O(gate194inter3));
  inv1  gate1447(.a(s_129), .O(gate194inter4));
  nand2 gate1448(.a(gate194inter4), .b(gate194inter3), .O(gate194inter5));
  nor2  gate1449(.a(gate194inter5), .b(gate194inter2), .O(gate194inter6));
  inv1  gate1450(.a(G588), .O(gate194inter7));
  inv1  gate1451(.a(G589), .O(gate194inter8));
  nand2 gate1452(.a(gate194inter8), .b(gate194inter7), .O(gate194inter9));
  nand2 gate1453(.a(s_129), .b(gate194inter3), .O(gate194inter10));
  nor2  gate1454(.a(gate194inter10), .b(gate194inter9), .O(gate194inter11));
  nor2  gate1455(.a(gate194inter11), .b(gate194inter6), .O(gate194inter12));
  nand2 gate1456(.a(gate194inter12), .b(gate194inter1), .O(G645));

  xor2  gate1065(.a(G591), .b(G590), .O(gate195inter0));
  nand2 gate1066(.a(gate195inter0), .b(s_74), .O(gate195inter1));
  and2  gate1067(.a(G591), .b(G590), .O(gate195inter2));
  inv1  gate1068(.a(s_74), .O(gate195inter3));
  inv1  gate1069(.a(s_75), .O(gate195inter4));
  nand2 gate1070(.a(gate195inter4), .b(gate195inter3), .O(gate195inter5));
  nor2  gate1071(.a(gate195inter5), .b(gate195inter2), .O(gate195inter6));
  inv1  gate1072(.a(G590), .O(gate195inter7));
  inv1  gate1073(.a(G591), .O(gate195inter8));
  nand2 gate1074(.a(gate195inter8), .b(gate195inter7), .O(gate195inter9));
  nand2 gate1075(.a(s_75), .b(gate195inter3), .O(gate195inter10));
  nor2  gate1076(.a(gate195inter10), .b(gate195inter9), .O(gate195inter11));
  nor2  gate1077(.a(gate195inter11), .b(gate195inter6), .O(gate195inter12));
  nand2 gate1078(.a(gate195inter12), .b(gate195inter1), .O(G648));
nand2 gate196( .a(G592), .b(G593), .O(G651) );
nand2 gate197( .a(G594), .b(G595), .O(G654) );

  xor2  gate701(.a(G597), .b(G596), .O(gate198inter0));
  nand2 gate702(.a(gate198inter0), .b(s_22), .O(gate198inter1));
  and2  gate703(.a(G597), .b(G596), .O(gate198inter2));
  inv1  gate704(.a(s_22), .O(gate198inter3));
  inv1  gate705(.a(s_23), .O(gate198inter4));
  nand2 gate706(.a(gate198inter4), .b(gate198inter3), .O(gate198inter5));
  nor2  gate707(.a(gate198inter5), .b(gate198inter2), .O(gate198inter6));
  inv1  gate708(.a(G596), .O(gate198inter7));
  inv1  gate709(.a(G597), .O(gate198inter8));
  nand2 gate710(.a(gate198inter8), .b(gate198inter7), .O(gate198inter9));
  nand2 gate711(.a(s_23), .b(gate198inter3), .O(gate198inter10));
  nor2  gate712(.a(gate198inter10), .b(gate198inter9), .O(gate198inter11));
  nor2  gate713(.a(gate198inter11), .b(gate198inter6), .O(gate198inter12));
  nand2 gate714(.a(gate198inter12), .b(gate198inter1), .O(G657));

  xor2  gate2535(.a(G599), .b(G598), .O(gate199inter0));
  nand2 gate2536(.a(gate199inter0), .b(s_284), .O(gate199inter1));
  and2  gate2537(.a(G599), .b(G598), .O(gate199inter2));
  inv1  gate2538(.a(s_284), .O(gate199inter3));
  inv1  gate2539(.a(s_285), .O(gate199inter4));
  nand2 gate2540(.a(gate199inter4), .b(gate199inter3), .O(gate199inter5));
  nor2  gate2541(.a(gate199inter5), .b(gate199inter2), .O(gate199inter6));
  inv1  gate2542(.a(G598), .O(gate199inter7));
  inv1  gate2543(.a(G599), .O(gate199inter8));
  nand2 gate2544(.a(gate199inter8), .b(gate199inter7), .O(gate199inter9));
  nand2 gate2545(.a(s_285), .b(gate199inter3), .O(gate199inter10));
  nor2  gate2546(.a(gate199inter10), .b(gate199inter9), .O(gate199inter11));
  nor2  gate2547(.a(gate199inter11), .b(gate199inter6), .O(gate199inter12));
  nand2 gate2548(.a(gate199inter12), .b(gate199inter1), .O(G660));
nand2 gate200( .a(G600), .b(G601), .O(G663) );

  xor2  gate2325(.a(G607), .b(G602), .O(gate201inter0));
  nand2 gate2326(.a(gate201inter0), .b(s_254), .O(gate201inter1));
  and2  gate2327(.a(G607), .b(G602), .O(gate201inter2));
  inv1  gate2328(.a(s_254), .O(gate201inter3));
  inv1  gate2329(.a(s_255), .O(gate201inter4));
  nand2 gate2330(.a(gate201inter4), .b(gate201inter3), .O(gate201inter5));
  nor2  gate2331(.a(gate201inter5), .b(gate201inter2), .O(gate201inter6));
  inv1  gate2332(.a(G602), .O(gate201inter7));
  inv1  gate2333(.a(G607), .O(gate201inter8));
  nand2 gate2334(.a(gate201inter8), .b(gate201inter7), .O(gate201inter9));
  nand2 gate2335(.a(s_255), .b(gate201inter3), .O(gate201inter10));
  nor2  gate2336(.a(gate201inter10), .b(gate201inter9), .O(gate201inter11));
  nor2  gate2337(.a(gate201inter11), .b(gate201inter6), .O(gate201inter12));
  nand2 gate2338(.a(gate201inter12), .b(gate201inter1), .O(G666));

  xor2  gate1723(.a(G617), .b(G612), .O(gate202inter0));
  nand2 gate1724(.a(gate202inter0), .b(s_168), .O(gate202inter1));
  and2  gate1725(.a(G617), .b(G612), .O(gate202inter2));
  inv1  gate1726(.a(s_168), .O(gate202inter3));
  inv1  gate1727(.a(s_169), .O(gate202inter4));
  nand2 gate1728(.a(gate202inter4), .b(gate202inter3), .O(gate202inter5));
  nor2  gate1729(.a(gate202inter5), .b(gate202inter2), .O(gate202inter6));
  inv1  gate1730(.a(G612), .O(gate202inter7));
  inv1  gate1731(.a(G617), .O(gate202inter8));
  nand2 gate1732(.a(gate202inter8), .b(gate202inter7), .O(gate202inter9));
  nand2 gate1733(.a(s_169), .b(gate202inter3), .O(gate202inter10));
  nor2  gate1734(.a(gate202inter10), .b(gate202inter9), .O(gate202inter11));
  nor2  gate1735(.a(gate202inter11), .b(gate202inter6), .O(gate202inter12));
  nand2 gate1736(.a(gate202inter12), .b(gate202inter1), .O(G669));
nand2 gate203( .a(G602), .b(G612), .O(G672) );
nand2 gate204( .a(G607), .b(G617), .O(G675) );

  xor2  gate1457(.a(G627), .b(G622), .O(gate205inter0));
  nand2 gate1458(.a(gate205inter0), .b(s_130), .O(gate205inter1));
  and2  gate1459(.a(G627), .b(G622), .O(gate205inter2));
  inv1  gate1460(.a(s_130), .O(gate205inter3));
  inv1  gate1461(.a(s_131), .O(gate205inter4));
  nand2 gate1462(.a(gate205inter4), .b(gate205inter3), .O(gate205inter5));
  nor2  gate1463(.a(gate205inter5), .b(gate205inter2), .O(gate205inter6));
  inv1  gate1464(.a(G622), .O(gate205inter7));
  inv1  gate1465(.a(G627), .O(gate205inter8));
  nand2 gate1466(.a(gate205inter8), .b(gate205inter7), .O(gate205inter9));
  nand2 gate1467(.a(s_131), .b(gate205inter3), .O(gate205inter10));
  nor2  gate1468(.a(gate205inter10), .b(gate205inter9), .O(gate205inter11));
  nor2  gate1469(.a(gate205inter11), .b(gate205inter6), .O(gate205inter12));
  nand2 gate1470(.a(gate205inter12), .b(gate205inter1), .O(G678));
nand2 gate206( .a(G632), .b(G637), .O(G681) );
nand2 gate207( .a(G622), .b(G632), .O(G684) );

  xor2  gate1933(.a(G637), .b(G627), .O(gate208inter0));
  nand2 gate1934(.a(gate208inter0), .b(s_198), .O(gate208inter1));
  and2  gate1935(.a(G637), .b(G627), .O(gate208inter2));
  inv1  gate1936(.a(s_198), .O(gate208inter3));
  inv1  gate1937(.a(s_199), .O(gate208inter4));
  nand2 gate1938(.a(gate208inter4), .b(gate208inter3), .O(gate208inter5));
  nor2  gate1939(.a(gate208inter5), .b(gate208inter2), .O(gate208inter6));
  inv1  gate1940(.a(G627), .O(gate208inter7));
  inv1  gate1941(.a(G637), .O(gate208inter8));
  nand2 gate1942(.a(gate208inter8), .b(gate208inter7), .O(gate208inter9));
  nand2 gate1943(.a(s_199), .b(gate208inter3), .O(gate208inter10));
  nor2  gate1944(.a(gate208inter10), .b(gate208inter9), .O(gate208inter11));
  nor2  gate1945(.a(gate208inter11), .b(gate208inter6), .O(gate208inter12));
  nand2 gate1946(.a(gate208inter12), .b(gate208inter1), .O(G687));

  xor2  gate2409(.a(G666), .b(G602), .O(gate209inter0));
  nand2 gate2410(.a(gate209inter0), .b(s_266), .O(gate209inter1));
  and2  gate2411(.a(G666), .b(G602), .O(gate209inter2));
  inv1  gate2412(.a(s_266), .O(gate209inter3));
  inv1  gate2413(.a(s_267), .O(gate209inter4));
  nand2 gate2414(.a(gate209inter4), .b(gate209inter3), .O(gate209inter5));
  nor2  gate2415(.a(gate209inter5), .b(gate209inter2), .O(gate209inter6));
  inv1  gate2416(.a(G602), .O(gate209inter7));
  inv1  gate2417(.a(G666), .O(gate209inter8));
  nand2 gate2418(.a(gate209inter8), .b(gate209inter7), .O(gate209inter9));
  nand2 gate2419(.a(s_267), .b(gate209inter3), .O(gate209inter10));
  nor2  gate2420(.a(gate209inter10), .b(gate209inter9), .O(gate209inter11));
  nor2  gate2421(.a(gate209inter11), .b(gate209inter6), .O(gate209inter12));
  nand2 gate2422(.a(gate209inter12), .b(gate209inter1), .O(G690));
nand2 gate210( .a(G607), .b(G666), .O(G691) );

  xor2  gate1233(.a(G669), .b(G612), .O(gate211inter0));
  nand2 gate1234(.a(gate211inter0), .b(s_98), .O(gate211inter1));
  and2  gate1235(.a(G669), .b(G612), .O(gate211inter2));
  inv1  gate1236(.a(s_98), .O(gate211inter3));
  inv1  gate1237(.a(s_99), .O(gate211inter4));
  nand2 gate1238(.a(gate211inter4), .b(gate211inter3), .O(gate211inter5));
  nor2  gate1239(.a(gate211inter5), .b(gate211inter2), .O(gate211inter6));
  inv1  gate1240(.a(G612), .O(gate211inter7));
  inv1  gate1241(.a(G669), .O(gate211inter8));
  nand2 gate1242(.a(gate211inter8), .b(gate211inter7), .O(gate211inter9));
  nand2 gate1243(.a(s_99), .b(gate211inter3), .O(gate211inter10));
  nor2  gate1244(.a(gate211inter10), .b(gate211inter9), .O(gate211inter11));
  nor2  gate1245(.a(gate211inter11), .b(gate211inter6), .O(gate211inter12));
  nand2 gate1246(.a(gate211inter12), .b(gate211inter1), .O(G692));

  xor2  gate967(.a(G669), .b(G617), .O(gate212inter0));
  nand2 gate968(.a(gate212inter0), .b(s_60), .O(gate212inter1));
  and2  gate969(.a(G669), .b(G617), .O(gate212inter2));
  inv1  gate970(.a(s_60), .O(gate212inter3));
  inv1  gate971(.a(s_61), .O(gate212inter4));
  nand2 gate972(.a(gate212inter4), .b(gate212inter3), .O(gate212inter5));
  nor2  gate973(.a(gate212inter5), .b(gate212inter2), .O(gate212inter6));
  inv1  gate974(.a(G617), .O(gate212inter7));
  inv1  gate975(.a(G669), .O(gate212inter8));
  nand2 gate976(.a(gate212inter8), .b(gate212inter7), .O(gate212inter9));
  nand2 gate977(.a(s_61), .b(gate212inter3), .O(gate212inter10));
  nor2  gate978(.a(gate212inter10), .b(gate212inter9), .O(gate212inter11));
  nor2  gate979(.a(gate212inter11), .b(gate212inter6), .O(gate212inter12));
  nand2 gate980(.a(gate212inter12), .b(gate212inter1), .O(G693));

  xor2  gate1079(.a(G672), .b(G602), .O(gate213inter0));
  nand2 gate1080(.a(gate213inter0), .b(s_76), .O(gate213inter1));
  and2  gate1081(.a(G672), .b(G602), .O(gate213inter2));
  inv1  gate1082(.a(s_76), .O(gate213inter3));
  inv1  gate1083(.a(s_77), .O(gate213inter4));
  nand2 gate1084(.a(gate213inter4), .b(gate213inter3), .O(gate213inter5));
  nor2  gate1085(.a(gate213inter5), .b(gate213inter2), .O(gate213inter6));
  inv1  gate1086(.a(G602), .O(gate213inter7));
  inv1  gate1087(.a(G672), .O(gate213inter8));
  nand2 gate1088(.a(gate213inter8), .b(gate213inter7), .O(gate213inter9));
  nand2 gate1089(.a(s_77), .b(gate213inter3), .O(gate213inter10));
  nor2  gate1090(.a(gate213inter10), .b(gate213inter9), .O(gate213inter11));
  nor2  gate1091(.a(gate213inter11), .b(gate213inter6), .O(gate213inter12));
  nand2 gate1092(.a(gate213inter12), .b(gate213inter1), .O(G694));

  xor2  gate1765(.a(G672), .b(G612), .O(gate214inter0));
  nand2 gate1766(.a(gate214inter0), .b(s_174), .O(gate214inter1));
  and2  gate1767(.a(G672), .b(G612), .O(gate214inter2));
  inv1  gate1768(.a(s_174), .O(gate214inter3));
  inv1  gate1769(.a(s_175), .O(gate214inter4));
  nand2 gate1770(.a(gate214inter4), .b(gate214inter3), .O(gate214inter5));
  nor2  gate1771(.a(gate214inter5), .b(gate214inter2), .O(gate214inter6));
  inv1  gate1772(.a(G612), .O(gate214inter7));
  inv1  gate1773(.a(G672), .O(gate214inter8));
  nand2 gate1774(.a(gate214inter8), .b(gate214inter7), .O(gate214inter9));
  nand2 gate1775(.a(s_175), .b(gate214inter3), .O(gate214inter10));
  nor2  gate1776(.a(gate214inter10), .b(gate214inter9), .O(gate214inter11));
  nor2  gate1777(.a(gate214inter11), .b(gate214inter6), .O(gate214inter12));
  nand2 gate1778(.a(gate214inter12), .b(gate214inter1), .O(G695));
nand2 gate215( .a(G607), .b(G675), .O(G696) );
nand2 gate216( .a(G617), .b(G675), .O(G697) );
nand2 gate217( .a(G622), .b(G678), .O(G698) );
nand2 gate218( .a(G627), .b(G678), .O(G699) );

  xor2  gate1415(.a(G681), .b(G632), .O(gate219inter0));
  nand2 gate1416(.a(gate219inter0), .b(s_124), .O(gate219inter1));
  and2  gate1417(.a(G681), .b(G632), .O(gate219inter2));
  inv1  gate1418(.a(s_124), .O(gate219inter3));
  inv1  gate1419(.a(s_125), .O(gate219inter4));
  nand2 gate1420(.a(gate219inter4), .b(gate219inter3), .O(gate219inter5));
  nor2  gate1421(.a(gate219inter5), .b(gate219inter2), .O(gate219inter6));
  inv1  gate1422(.a(G632), .O(gate219inter7));
  inv1  gate1423(.a(G681), .O(gate219inter8));
  nand2 gate1424(.a(gate219inter8), .b(gate219inter7), .O(gate219inter9));
  nand2 gate1425(.a(s_125), .b(gate219inter3), .O(gate219inter10));
  nor2  gate1426(.a(gate219inter10), .b(gate219inter9), .O(gate219inter11));
  nor2  gate1427(.a(gate219inter11), .b(gate219inter6), .O(gate219inter12));
  nand2 gate1428(.a(gate219inter12), .b(gate219inter1), .O(G700));
nand2 gate220( .a(G637), .b(G681), .O(G701) );
nand2 gate221( .a(G622), .b(G684), .O(G702) );

  xor2  gate2563(.a(G684), .b(G632), .O(gate222inter0));
  nand2 gate2564(.a(gate222inter0), .b(s_288), .O(gate222inter1));
  and2  gate2565(.a(G684), .b(G632), .O(gate222inter2));
  inv1  gate2566(.a(s_288), .O(gate222inter3));
  inv1  gate2567(.a(s_289), .O(gate222inter4));
  nand2 gate2568(.a(gate222inter4), .b(gate222inter3), .O(gate222inter5));
  nor2  gate2569(.a(gate222inter5), .b(gate222inter2), .O(gate222inter6));
  inv1  gate2570(.a(G632), .O(gate222inter7));
  inv1  gate2571(.a(G684), .O(gate222inter8));
  nand2 gate2572(.a(gate222inter8), .b(gate222inter7), .O(gate222inter9));
  nand2 gate2573(.a(s_289), .b(gate222inter3), .O(gate222inter10));
  nor2  gate2574(.a(gate222inter10), .b(gate222inter9), .O(gate222inter11));
  nor2  gate2575(.a(gate222inter11), .b(gate222inter6), .O(gate222inter12));
  nand2 gate2576(.a(gate222inter12), .b(gate222inter1), .O(G703));
nand2 gate223( .a(G627), .b(G687), .O(G704) );

  xor2  gate939(.a(G687), .b(G637), .O(gate224inter0));
  nand2 gate940(.a(gate224inter0), .b(s_56), .O(gate224inter1));
  and2  gate941(.a(G687), .b(G637), .O(gate224inter2));
  inv1  gate942(.a(s_56), .O(gate224inter3));
  inv1  gate943(.a(s_57), .O(gate224inter4));
  nand2 gate944(.a(gate224inter4), .b(gate224inter3), .O(gate224inter5));
  nor2  gate945(.a(gate224inter5), .b(gate224inter2), .O(gate224inter6));
  inv1  gate946(.a(G637), .O(gate224inter7));
  inv1  gate947(.a(G687), .O(gate224inter8));
  nand2 gate948(.a(gate224inter8), .b(gate224inter7), .O(gate224inter9));
  nand2 gate949(.a(s_57), .b(gate224inter3), .O(gate224inter10));
  nor2  gate950(.a(gate224inter10), .b(gate224inter9), .O(gate224inter11));
  nor2  gate951(.a(gate224inter11), .b(gate224inter6), .O(gate224inter12));
  nand2 gate952(.a(gate224inter12), .b(gate224inter1), .O(G705));
nand2 gate225( .a(G690), .b(G691), .O(G706) );

  xor2  gate1163(.a(G693), .b(G692), .O(gate226inter0));
  nand2 gate1164(.a(gate226inter0), .b(s_88), .O(gate226inter1));
  and2  gate1165(.a(G693), .b(G692), .O(gate226inter2));
  inv1  gate1166(.a(s_88), .O(gate226inter3));
  inv1  gate1167(.a(s_89), .O(gate226inter4));
  nand2 gate1168(.a(gate226inter4), .b(gate226inter3), .O(gate226inter5));
  nor2  gate1169(.a(gate226inter5), .b(gate226inter2), .O(gate226inter6));
  inv1  gate1170(.a(G692), .O(gate226inter7));
  inv1  gate1171(.a(G693), .O(gate226inter8));
  nand2 gate1172(.a(gate226inter8), .b(gate226inter7), .O(gate226inter9));
  nand2 gate1173(.a(s_89), .b(gate226inter3), .O(gate226inter10));
  nor2  gate1174(.a(gate226inter10), .b(gate226inter9), .O(gate226inter11));
  nor2  gate1175(.a(gate226inter11), .b(gate226inter6), .O(gate226inter12));
  nand2 gate1176(.a(gate226inter12), .b(gate226inter1), .O(G709));
nand2 gate227( .a(G694), .b(G695), .O(G712) );

  xor2  gate1373(.a(G697), .b(G696), .O(gate228inter0));
  nand2 gate1374(.a(gate228inter0), .b(s_118), .O(gate228inter1));
  and2  gate1375(.a(G697), .b(G696), .O(gate228inter2));
  inv1  gate1376(.a(s_118), .O(gate228inter3));
  inv1  gate1377(.a(s_119), .O(gate228inter4));
  nand2 gate1378(.a(gate228inter4), .b(gate228inter3), .O(gate228inter5));
  nor2  gate1379(.a(gate228inter5), .b(gate228inter2), .O(gate228inter6));
  inv1  gate1380(.a(G696), .O(gate228inter7));
  inv1  gate1381(.a(G697), .O(gate228inter8));
  nand2 gate1382(.a(gate228inter8), .b(gate228inter7), .O(gate228inter9));
  nand2 gate1383(.a(s_119), .b(gate228inter3), .O(gate228inter10));
  nor2  gate1384(.a(gate228inter10), .b(gate228inter9), .O(gate228inter11));
  nor2  gate1385(.a(gate228inter11), .b(gate228inter6), .O(gate228inter12));
  nand2 gate1386(.a(gate228inter12), .b(gate228inter1), .O(G715));

  xor2  gate1793(.a(G699), .b(G698), .O(gate229inter0));
  nand2 gate1794(.a(gate229inter0), .b(s_178), .O(gate229inter1));
  and2  gate1795(.a(G699), .b(G698), .O(gate229inter2));
  inv1  gate1796(.a(s_178), .O(gate229inter3));
  inv1  gate1797(.a(s_179), .O(gate229inter4));
  nand2 gate1798(.a(gate229inter4), .b(gate229inter3), .O(gate229inter5));
  nor2  gate1799(.a(gate229inter5), .b(gate229inter2), .O(gate229inter6));
  inv1  gate1800(.a(G698), .O(gate229inter7));
  inv1  gate1801(.a(G699), .O(gate229inter8));
  nand2 gate1802(.a(gate229inter8), .b(gate229inter7), .O(gate229inter9));
  nand2 gate1803(.a(s_179), .b(gate229inter3), .O(gate229inter10));
  nor2  gate1804(.a(gate229inter10), .b(gate229inter9), .O(gate229inter11));
  nor2  gate1805(.a(gate229inter11), .b(gate229inter6), .O(gate229inter12));
  nand2 gate1806(.a(gate229inter12), .b(gate229inter1), .O(G718));
nand2 gate230( .a(G700), .b(G701), .O(G721) );
nand2 gate231( .a(G702), .b(G703), .O(G724) );

  xor2  gate617(.a(G705), .b(G704), .O(gate232inter0));
  nand2 gate618(.a(gate232inter0), .b(s_10), .O(gate232inter1));
  and2  gate619(.a(G705), .b(G704), .O(gate232inter2));
  inv1  gate620(.a(s_10), .O(gate232inter3));
  inv1  gate621(.a(s_11), .O(gate232inter4));
  nand2 gate622(.a(gate232inter4), .b(gate232inter3), .O(gate232inter5));
  nor2  gate623(.a(gate232inter5), .b(gate232inter2), .O(gate232inter6));
  inv1  gate624(.a(G704), .O(gate232inter7));
  inv1  gate625(.a(G705), .O(gate232inter8));
  nand2 gate626(.a(gate232inter8), .b(gate232inter7), .O(gate232inter9));
  nand2 gate627(.a(s_11), .b(gate232inter3), .O(gate232inter10));
  nor2  gate628(.a(gate232inter10), .b(gate232inter9), .O(gate232inter11));
  nor2  gate629(.a(gate232inter11), .b(gate232inter6), .O(gate232inter12));
  nand2 gate630(.a(gate232inter12), .b(gate232inter1), .O(G727));

  xor2  gate2339(.a(G718), .b(G242), .O(gate233inter0));
  nand2 gate2340(.a(gate233inter0), .b(s_256), .O(gate233inter1));
  and2  gate2341(.a(G718), .b(G242), .O(gate233inter2));
  inv1  gate2342(.a(s_256), .O(gate233inter3));
  inv1  gate2343(.a(s_257), .O(gate233inter4));
  nand2 gate2344(.a(gate233inter4), .b(gate233inter3), .O(gate233inter5));
  nor2  gate2345(.a(gate233inter5), .b(gate233inter2), .O(gate233inter6));
  inv1  gate2346(.a(G242), .O(gate233inter7));
  inv1  gate2347(.a(G718), .O(gate233inter8));
  nand2 gate2348(.a(gate233inter8), .b(gate233inter7), .O(gate233inter9));
  nand2 gate2349(.a(s_257), .b(gate233inter3), .O(gate233inter10));
  nor2  gate2350(.a(gate233inter10), .b(gate233inter9), .O(gate233inter11));
  nor2  gate2351(.a(gate233inter11), .b(gate233inter6), .O(gate233inter12));
  nand2 gate2352(.a(gate233inter12), .b(gate233inter1), .O(G730));

  xor2  gate1919(.a(G721), .b(G245), .O(gate234inter0));
  nand2 gate1920(.a(gate234inter0), .b(s_196), .O(gate234inter1));
  and2  gate1921(.a(G721), .b(G245), .O(gate234inter2));
  inv1  gate1922(.a(s_196), .O(gate234inter3));
  inv1  gate1923(.a(s_197), .O(gate234inter4));
  nand2 gate1924(.a(gate234inter4), .b(gate234inter3), .O(gate234inter5));
  nor2  gate1925(.a(gate234inter5), .b(gate234inter2), .O(gate234inter6));
  inv1  gate1926(.a(G245), .O(gate234inter7));
  inv1  gate1927(.a(G721), .O(gate234inter8));
  nand2 gate1928(.a(gate234inter8), .b(gate234inter7), .O(gate234inter9));
  nand2 gate1929(.a(s_197), .b(gate234inter3), .O(gate234inter10));
  nor2  gate1930(.a(gate234inter10), .b(gate234inter9), .O(gate234inter11));
  nor2  gate1931(.a(gate234inter11), .b(gate234inter6), .O(gate234inter12));
  nand2 gate1932(.a(gate234inter12), .b(gate234inter1), .O(G733));
nand2 gate235( .a(G248), .b(G724), .O(G736) );
nand2 gate236( .a(G251), .b(G727), .O(G739) );

  xor2  gate1317(.a(G706), .b(G254), .O(gate237inter0));
  nand2 gate1318(.a(gate237inter0), .b(s_110), .O(gate237inter1));
  and2  gate1319(.a(G706), .b(G254), .O(gate237inter2));
  inv1  gate1320(.a(s_110), .O(gate237inter3));
  inv1  gate1321(.a(s_111), .O(gate237inter4));
  nand2 gate1322(.a(gate237inter4), .b(gate237inter3), .O(gate237inter5));
  nor2  gate1323(.a(gate237inter5), .b(gate237inter2), .O(gate237inter6));
  inv1  gate1324(.a(G254), .O(gate237inter7));
  inv1  gate1325(.a(G706), .O(gate237inter8));
  nand2 gate1326(.a(gate237inter8), .b(gate237inter7), .O(gate237inter9));
  nand2 gate1327(.a(s_111), .b(gate237inter3), .O(gate237inter10));
  nor2  gate1328(.a(gate237inter10), .b(gate237inter9), .O(gate237inter11));
  nor2  gate1329(.a(gate237inter11), .b(gate237inter6), .O(gate237inter12));
  nand2 gate1330(.a(gate237inter12), .b(gate237inter1), .O(G742));

  xor2  gate2857(.a(G709), .b(G257), .O(gate238inter0));
  nand2 gate2858(.a(gate238inter0), .b(s_330), .O(gate238inter1));
  and2  gate2859(.a(G709), .b(G257), .O(gate238inter2));
  inv1  gate2860(.a(s_330), .O(gate238inter3));
  inv1  gate2861(.a(s_331), .O(gate238inter4));
  nand2 gate2862(.a(gate238inter4), .b(gate238inter3), .O(gate238inter5));
  nor2  gate2863(.a(gate238inter5), .b(gate238inter2), .O(gate238inter6));
  inv1  gate2864(.a(G257), .O(gate238inter7));
  inv1  gate2865(.a(G709), .O(gate238inter8));
  nand2 gate2866(.a(gate238inter8), .b(gate238inter7), .O(gate238inter9));
  nand2 gate2867(.a(s_331), .b(gate238inter3), .O(gate238inter10));
  nor2  gate2868(.a(gate238inter10), .b(gate238inter9), .O(gate238inter11));
  nor2  gate2869(.a(gate238inter11), .b(gate238inter6), .O(gate238inter12));
  nand2 gate2870(.a(gate238inter12), .b(gate238inter1), .O(G745));
nand2 gate239( .a(G260), .b(G712), .O(G748) );
nand2 gate240( .a(G263), .b(G715), .O(G751) );
nand2 gate241( .a(G242), .b(G730), .O(G754) );
nand2 gate242( .a(G718), .b(G730), .O(G755) );
nand2 gate243( .a(G245), .b(G733), .O(G756) );

  xor2  gate2983(.a(G733), .b(G721), .O(gate244inter0));
  nand2 gate2984(.a(gate244inter0), .b(s_348), .O(gate244inter1));
  and2  gate2985(.a(G733), .b(G721), .O(gate244inter2));
  inv1  gate2986(.a(s_348), .O(gate244inter3));
  inv1  gate2987(.a(s_349), .O(gate244inter4));
  nand2 gate2988(.a(gate244inter4), .b(gate244inter3), .O(gate244inter5));
  nor2  gate2989(.a(gate244inter5), .b(gate244inter2), .O(gate244inter6));
  inv1  gate2990(.a(G721), .O(gate244inter7));
  inv1  gate2991(.a(G733), .O(gate244inter8));
  nand2 gate2992(.a(gate244inter8), .b(gate244inter7), .O(gate244inter9));
  nand2 gate2993(.a(s_349), .b(gate244inter3), .O(gate244inter10));
  nor2  gate2994(.a(gate244inter10), .b(gate244inter9), .O(gate244inter11));
  nor2  gate2995(.a(gate244inter11), .b(gate244inter6), .O(gate244inter12));
  nand2 gate2996(.a(gate244inter12), .b(gate244inter1), .O(G757));
nand2 gate245( .a(G248), .b(G736), .O(G758) );
nand2 gate246( .a(G724), .b(G736), .O(G759) );
nand2 gate247( .a(G251), .b(G739), .O(G760) );

  xor2  gate2843(.a(G739), .b(G727), .O(gate248inter0));
  nand2 gate2844(.a(gate248inter0), .b(s_328), .O(gate248inter1));
  and2  gate2845(.a(G739), .b(G727), .O(gate248inter2));
  inv1  gate2846(.a(s_328), .O(gate248inter3));
  inv1  gate2847(.a(s_329), .O(gate248inter4));
  nand2 gate2848(.a(gate248inter4), .b(gate248inter3), .O(gate248inter5));
  nor2  gate2849(.a(gate248inter5), .b(gate248inter2), .O(gate248inter6));
  inv1  gate2850(.a(G727), .O(gate248inter7));
  inv1  gate2851(.a(G739), .O(gate248inter8));
  nand2 gate2852(.a(gate248inter8), .b(gate248inter7), .O(gate248inter9));
  nand2 gate2853(.a(s_329), .b(gate248inter3), .O(gate248inter10));
  nor2  gate2854(.a(gate248inter10), .b(gate248inter9), .O(gate248inter11));
  nor2  gate2855(.a(gate248inter11), .b(gate248inter6), .O(gate248inter12));
  nand2 gate2856(.a(gate248inter12), .b(gate248inter1), .O(G761));
nand2 gate249( .a(G254), .b(G742), .O(G762) );

  xor2  gate2717(.a(G742), .b(G706), .O(gate250inter0));
  nand2 gate2718(.a(gate250inter0), .b(s_310), .O(gate250inter1));
  and2  gate2719(.a(G742), .b(G706), .O(gate250inter2));
  inv1  gate2720(.a(s_310), .O(gate250inter3));
  inv1  gate2721(.a(s_311), .O(gate250inter4));
  nand2 gate2722(.a(gate250inter4), .b(gate250inter3), .O(gate250inter5));
  nor2  gate2723(.a(gate250inter5), .b(gate250inter2), .O(gate250inter6));
  inv1  gate2724(.a(G706), .O(gate250inter7));
  inv1  gate2725(.a(G742), .O(gate250inter8));
  nand2 gate2726(.a(gate250inter8), .b(gate250inter7), .O(gate250inter9));
  nand2 gate2727(.a(s_311), .b(gate250inter3), .O(gate250inter10));
  nor2  gate2728(.a(gate250inter10), .b(gate250inter9), .O(gate250inter11));
  nor2  gate2729(.a(gate250inter11), .b(gate250inter6), .O(gate250inter12));
  nand2 gate2730(.a(gate250inter12), .b(gate250inter1), .O(G763));

  xor2  gate1177(.a(G745), .b(G257), .O(gate251inter0));
  nand2 gate1178(.a(gate251inter0), .b(s_90), .O(gate251inter1));
  and2  gate1179(.a(G745), .b(G257), .O(gate251inter2));
  inv1  gate1180(.a(s_90), .O(gate251inter3));
  inv1  gate1181(.a(s_91), .O(gate251inter4));
  nand2 gate1182(.a(gate251inter4), .b(gate251inter3), .O(gate251inter5));
  nor2  gate1183(.a(gate251inter5), .b(gate251inter2), .O(gate251inter6));
  inv1  gate1184(.a(G257), .O(gate251inter7));
  inv1  gate1185(.a(G745), .O(gate251inter8));
  nand2 gate1186(.a(gate251inter8), .b(gate251inter7), .O(gate251inter9));
  nand2 gate1187(.a(s_91), .b(gate251inter3), .O(gate251inter10));
  nor2  gate1188(.a(gate251inter10), .b(gate251inter9), .O(gate251inter11));
  nor2  gate1189(.a(gate251inter11), .b(gate251inter6), .O(gate251inter12));
  nand2 gate1190(.a(gate251inter12), .b(gate251inter1), .O(G764));
nand2 gate252( .a(G709), .b(G745), .O(G765) );

  xor2  gate1303(.a(G748), .b(G260), .O(gate253inter0));
  nand2 gate1304(.a(gate253inter0), .b(s_108), .O(gate253inter1));
  and2  gate1305(.a(G748), .b(G260), .O(gate253inter2));
  inv1  gate1306(.a(s_108), .O(gate253inter3));
  inv1  gate1307(.a(s_109), .O(gate253inter4));
  nand2 gate1308(.a(gate253inter4), .b(gate253inter3), .O(gate253inter5));
  nor2  gate1309(.a(gate253inter5), .b(gate253inter2), .O(gate253inter6));
  inv1  gate1310(.a(G260), .O(gate253inter7));
  inv1  gate1311(.a(G748), .O(gate253inter8));
  nand2 gate1312(.a(gate253inter8), .b(gate253inter7), .O(gate253inter9));
  nand2 gate1313(.a(s_109), .b(gate253inter3), .O(gate253inter10));
  nor2  gate1314(.a(gate253inter10), .b(gate253inter9), .O(gate253inter11));
  nor2  gate1315(.a(gate253inter11), .b(gate253inter6), .O(gate253inter12));
  nand2 gate1316(.a(gate253inter12), .b(gate253inter1), .O(G766));
nand2 gate254( .a(G712), .b(G748), .O(G767) );

  xor2  gate2913(.a(G751), .b(G263), .O(gate255inter0));
  nand2 gate2914(.a(gate255inter0), .b(s_338), .O(gate255inter1));
  and2  gate2915(.a(G751), .b(G263), .O(gate255inter2));
  inv1  gate2916(.a(s_338), .O(gate255inter3));
  inv1  gate2917(.a(s_339), .O(gate255inter4));
  nand2 gate2918(.a(gate255inter4), .b(gate255inter3), .O(gate255inter5));
  nor2  gate2919(.a(gate255inter5), .b(gate255inter2), .O(gate255inter6));
  inv1  gate2920(.a(G263), .O(gate255inter7));
  inv1  gate2921(.a(G751), .O(gate255inter8));
  nand2 gate2922(.a(gate255inter8), .b(gate255inter7), .O(gate255inter9));
  nand2 gate2923(.a(s_339), .b(gate255inter3), .O(gate255inter10));
  nor2  gate2924(.a(gate255inter10), .b(gate255inter9), .O(gate255inter11));
  nor2  gate2925(.a(gate255inter11), .b(gate255inter6), .O(gate255inter12));
  nand2 gate2926(.a(gate255inter12), .b(gate255inter1), .O(G768));
nand2 gate256( .a(G715), .b(G751), .O(G769) );
nand2 gate257( .a(G754), .b(G755), .O(G770) );
nand2 gate258( .a(G756), .b(G757), .O(G773) );
nand2 gate259( .a(G758), .b(G759), .O(G776) );
nand2 gate260( .a(G760), .b(G761), .O(G779) );
nand2 gate261( .a(G762), .b(G763), .O(G782) );

  xor2  gate1555(.a(G765), .b(G764), .O(gate262inter0));
  nand2 gate1556(.a(gate262inter0), .b(s_144), .O(gate262inter1));
  and2  gate1557(.a(G765), .b(G764), .O(gate262inter2));
  inv1  gate1558(.a(s_144), .O(gate262inter3));
  inv1  gate1559(.a(s_145), .O(gate262inter4));
  nand2 gate1560(.a(gate262inter4), .b(gate262inter3), .O(gate262inter5));
  nor2  gate1561(.a(gate262inter5), .b(gate262inter2), .O(gate262inter6));
  inv1  gate1562(.a(G764), .O(gate262inter7));
  inv1  gate1563(.a(G765), .O(gate262inter8));
  nand2 gate1564(.a(gate262inter8), .b(gate262inter7), .O(gate262inter9));
  nand2 gate1565(.a(s_145), .b(gate262inter3), .O(gate262inter10));
  nor2  gate1566(.a(gate262inter10), .b(gate262inter9), .O(gate262inter11));
  nor2  gate1567(.a(gate262inter11), .b(gate262inter6), .O(gate262inter12));
  nand2 gate1568(.a(gate262inter12), .b(gate262inter1), .O(G785));

  xor2  gate883(.a(G767), .b(G766), .O(gate263inter0));
  nand2 gate884(.a(gate263inter0), .b(s_48), .O(gate263inter1));
  and2  gate885(.a(G767), .b(G766), .O(gate263inter2));
  inv1  gate886(.a(s_48), .O(gate263inter3));
  inv1  gate887(.a(s_49), .O(gate263inter4));
  nand2 gate888(.a(gate263inter4), .b(gate263inter3), .O(gate263inter5));
  nor2  gate889(.a(gate263inter5), .b(gate263inter2), .O(gate263inter6));
  inv1  gate890(.a(G766), .O(gate263inter7));
  inv1  gate891(.a(G767), .O(gate263inter8));
  nand2 gate892(.a(gate263inter8), .b(gate263inter7), .O(gate263inter9));
  nand2 gate893(.a(s_49), .b(gate263inter3), .O(gate263inter10));
  nor2  gate894(.a(gate263inter10), .b(gate263inter9), .O(gate263inter11));
  nor2  gate895(.a(gate263inter11), .b(gate263inter6), .O(gate263inter12));
  nand2 gate896(.a(gate263inter12), .b(gate263inter1), .O(G788));
nand2 gate264( .a(G768), .b(G769), .O(G791) );

  xor2  gate2437(.a(G770), .b(G642), .O(gate265inter0));
  nand2 gate2438(.a(gate265inter0), .b(s_270), .O(gate265inter1));
  and2  gate2439(.a(G770), .b(G642), .O(gate265inter2));
  inv1  gate2440(.a(s_270), .O(gate265inter3));
  inv1  gate2441(.a(s_271), .O(gate265inter4));
  nand2 gate2442(.a(gate265inter4), .b(gate265inter3), .O(gate265inter5));
  nor2  gate2443(.a(gate265inter5), .b(gate265inter2), .O(gate265inter6));
  inv1  gate2444(.a(G642), .O(gate265inter7));
  inv1  gate2445(.a(G770), .O(gate265inter8));
  nand2 gate2446(.a(gate265inter8), .b(gate265inter7), .O(gate265inter9));
  nand2 gate2447(.a(s_271), .b(gate265inter3), .O(gate265inter10));
  nor2  gate2448(.a(gate265inter10), .b(gate265inter9), .O(gate265inter11));
  nor2  gate2449(.a(gate265inter11), .b(gate265inter6), .O(gate265inter12));
  nand2 gate2450(.a(gate265inter12), .b(gate265inter1), .O(G794));

  xor2  gate2605(.a(G773), .b(G645), .O(gate266inter0));
  nand2 gate2606(.a(gate266inter0), .b(s_294), .O(gate266inter1));
  and2  gate2607(.a(G773), .b(G645), .O(gate266inter2));
  inv1  gate2608(.a(s_294), .O(gate266inter3));
  inv1  gate2609(.a(s_295), .O(gate266inter4));
  nand2 gate2610(.a(gate266inter4), .b(gate266inter3), .O(gate266inter5));
  nor2  gate2611(.a(gate266inter5), .b(gate266inter2), .O(gate266inter6));
  inv1  gate2612(.a(G645), .O(gate266inter7));
  inv1  gate2613(.a(G773), .O(gate266inter8));
  nand2 gate2614(.a(gate266inter8), .b(gate266inter7), .O(gate266inter9));
  nand2 gate2615(.a(s_295), .b(gate266inter3), .O(gate266inter10));
  nor2  gate2616(.a(gate266inter10), .b(gate266inter9), .O(gate266inter11));
  nor2  gate2617(.a(gate266inter11), .b(gate266inter6), .O(gate266inter12));
  nand2 gate2618(.a(gate266inter12), .b(gate266inter1), .O(G797));
nand2 gate267( .a(G648), .b(G776), .O(G800) );

  xor2  gate1107(.a(G779), .b(G651), .O(gate268inter0));
  nand2 gate1108(.a(gate268inter0), .b(s_80), .O(gate268inter1));
  and2  gate1109(.a(G779), .b(G651), .O(gate268inter2));
  inv1  gate1110(.a(s_80), .O(gate268inter3));
  inv1  gate1111(.a(s_81), .O(gate268inter4));
  nand2 gate1112(.a(gate268inter4), .b(gate268inter3), .O(gate268inter5));
  nor2  gate1113(.a(gate268inter5), .b(gate268inter2), .O(gate268inter6));
  inv1  gate1114(.a(G651), .O(gate268inter7));
  inv1  gate1115(.a(G779), .O(gate268inter8));
  nand2 gate1116(.a(gate268inter8), .b(gate268inter7), .O(gate268inter9));
  nand2 gate1117(.a(s_81), .b(gate268inter3), .O(gate268inter10));
  nor2  gate1118(.a(gate268inter10), .b(gate268inter9), .O(gate268inter11));
  nor2  gate1119(.a(gate268inter11), .b(gate268inter6), .O(gate268inter12));
  nand2 gate1120(.a(gate268inter12), .b(gate268inter1), .O(G803));
nand2 gate269( .a(G654), .b(G782), .O(G806) );

  xor2  gate1387(.a(G785), .b(G657), .O(gate270inter0));
  nand2 gate1388(.a(gate270inter0), .b(s_120), .O(gate270inter1));
  and2  gate1389(.a(G785), .b(G657), .O(gate270inter2));
  inv1  gate1390(.a(s_120), .O(gate270inter3));
  inv1  gate1391(.a(s_121), .O(gate270inter4));
  nand2 gate1392(.a(gate270inter4), .b(gate270inter3), .O(gate270inter5));
  nor2  gate1393(.a(gate270inter5), .b(gate270inter2), .O(gate270inter6));
  inv1  gate1394(.a(G657), .O(gate270inter7));
  inv1  gate1395(.a(G785), .O(gate270inter8));
  nand2 gate1396(.a(gate270inter8), .b(gate270inter7), .O(gate270inter9));
  nand2 gate1397(.a(s_121), .b(gate270inter3), .O(gate270inter10));
  nor2  gate1398(.a(gate270inter10), .b(gate270inter9), .O(gate270inter11));
  nor2  gate1399(.a(gate270inter11), .b(gate270inter6), .O(gate270inter12));
  nand2 gate1400(.a(gate270inter12), .b(gate270inter1), .O(G809));
nand2 gate271( .a(G660), .b(G788), .O(G812) );
nand2 gate272( .a(G663), .b(G791), .O(G815) );
nand2 gate273( .a(G642), .b(G794), .O(G818) );
nand2 gate274( .a(G770), .b(G794), .O(G819) );
nand2 gate275( .a(G645), .b(G797), .O(G820) );
nand2 gate276( .a(G773), .b(G797), .O(G821) );
nand2 gate277( .a(G648), .b(G800), .O(G822) );
nand2 gate278( .a(G776), .b(G800), .O(G823) );
nand2 gate279( .a(G651), .b(G803), .O(G824) );

  xor2  gate2199(.a(G803), .b(G779), .O(gate280inter0));
  nand2 gate2200(.a(gate280inter0), .b(s_236), .O(gate280inter1));
  and2  gate2201(.a(G803), .b(G779), .O(gate280inter2));
  inv1  gate2202(.a(s_236), .O(gate280inter3));
  inv1  gate2203(.a(s_237), .O(gate280inter4));
  nand2 gate2204(.a(gate280inter4), .b(gate280inter3), .O(gate280inter5));
  nor2  gate2205(.a(gate280inter5), .b(gate280inter2), .O(gate280inter6));
  inv1  gate2206(.a(G779), .O(gate280inter7));
  inv1  gate2207(.a(G803), .O(gate280inter8));
  nand2 gate2208(.a(gate280inter8), .b(gate280inter7), .O(gate280inter9));
  nand2 gate2209(.a(s_237), .b(gate280inter3), .O(gate280inter10));
  nor2  gate2210(.a(gate280inter10), .b(gate280inter9), .O(gate280inter11));
  nor2  gate2211(.a(gate280inter11), .b(gate280inter6), .O(gate280inter12));
  nand2 gate2212(.a(gate280inter12), .b(gate280inter1), .O(G825));

  xor2  gate1989(.a(G806), .b(G654), .O(gate281inter0));
  nand2 gate1990(.a(gate281inter0), .b(s_206), .O(gate281inter1));
  and2  gate1991(.a(G806), .b(G654), .O(gate281inter2));
  inv1  gate1992(.a(s_206), .O(gate281inter3));
  inv1  gate1993(.a(s_207), .O(gate281inter4));
  nand2 gate1994(.a(gate281inter4), .b(gate281inter3), .O(gate281inter5));
  nor2  gate1995(.a(gate281inter5), .b(gate281inter2), .O(gate281inter6));
  inv1  gate1996(.a(G654), .O(gate281inter7));
  inv1  gate1997(.a(G806), .O(gate281inter8));
  nand2 gate1998(.a(gate281inter8), .b(gate281inter7), .O(gate281inter9));
  nand2 gate1999(.a(s_207), .b(gate281inter3), .O(gate281inter10));
  nor2  gate2000(.a(gate281inter10), .b(gate281inter9), .O(gate281inter11));
  nor2  gate2001(.a(gate281inter11), .b(gate281inter6), .O(gate281inter12));
  nand2 gate2002(.a(gate281inter12), .b(gate281inter1), .O(G826));

  xor2  gate2017(.a(G806), .b(G782), .O(gate282inter0));
  nand2 gate2018(.a(gate282inter0), .b(s_210), .O(gate282inter1));
  and2  gate2019(.a(G806), .b(G782), .O(gate282inter2));
  inv1  gate2020(.a(s_210), .O(gate282inter3));
  inv1  gate2021(.a(s_211), .O(gate282inter4));
  nand2 gate2022(.a(gate282inter4), .b(gate282inter3), .O(gate282inter5));
  nor2  gate2023(.a(gate282inter5), .b(gate282inter2), .O(gate282inter6));
  inv1  gate2024(.a(G782), .O(gate282inter7));
  inv1  gate2025(.a(G806), .O(gate282inter8));
  nand2 gate2026(.a(gate282inter8), .b(gate282inter7), .O(gate282inter9));
  nand2 gate2027(.a(s_211), .b(gate282inter3), .O(gate282inter10));
  nor2  gate2028(.a(gate282inter10), .b(gate282inter9), .O(gate282inter11));
  nor2  gate2029(.a(gate282inter11), .b(gate282inter6), .O(gate282inter12));
  nand2 gate2030(.a(gate282inter12), .b(gate282inter1), .O(G827));

  xor2  gate2395(.a(G809), .b(G657), .O(gate283inter0));
  nand2 gate2396(.a(gate283inter0), .b(s_264), .O(gate283inter1));
  and2  gate2397(.a(G809), .b(G657), .O(gate283inter2));
  inv1  gate2398(.a(s_264), .O(gate283inter3));
  inv1  gate2399(.a(s_265), .O(gate283inter4));
  nand2 gate2400(.a(gate283inter4), .b(gate283inter3), .O(gate283inter5));
  nor2  gate2401(.a(gate283inter5), .b(gate283inter2), .O(gate283inter6));
  inv1  gate2402(.a(G657), .O(gate283inter7));
  inv1  gate2403(.a(G809), .O(gate283inter8));
  nand2 gate2404(.a(gate283inter8), .b(gate283inter7), .O(gate283inter9));
  nand2 gate2405(.a(s_265), .b(gate283inter3), .O(gate283inter10));
  nor2  gate2406(.a(gate283inter10), .b(gate283inter9), .O(gate283inter11));
  nor2  gate2407(.a(gate283inter11), .b(gate283inter6), .O(gate283inter12));
  nand2 gate2408(.a(gate283inter12), .b(gate283inter1), .O(G828));
nand2 gate284( .a(G785), .b(G809), .O(G829) );

  xor2  gate1849(.a(G812), .b(G660), .O(gate285inter0));
  nand2 gate1850(.a(gate285inter0), .b(s_186), .O(gate285inter1));
  and2  gate1851(.a(G812), .b(G660), .O(gate285inter2));
  inv1  gate1852(.a(s_186), .O(gate285inter3));
  inv1  gate1853(.a(s_187), .O(gate285inter4));
  nand2 gate1854(.a(gate285inter4), .b(gate285inter3), .O(gate285inter5));
  nor2  gate1855(.a(gate285inter5), .b(gate285inter2), .O(gate285inter6));
  inv1  gate1856(.a(G660), .O(gate285inter7));
  inv1  gate1857(.a(G812), .O(gate285inter8));
  nand2 gate1858(.a(gate285inter8), .b(gate285inter7), .O(gate285inter9));
  nand2 gate1859(.a(s_187), .b(gate285inter3), .O(gate285inter10));
  nor2  gate1860(.a(gate285inter10), .b(gate285inter9), .O(gate285inter11));
  nor2  gate1861(.a(gate285inter11), .b(gate285inter6), .O(gate285inter12));
  nand2 gate1862(.a(gate285inter12), .b(gate285inter1), .O(G830));
nand2 gate286( .a(G788), .b(G812), .O(G831) );
nand2 gate287( .a(G663), .b(G815), .O(G832) );
nand2 gate288( .a(G791), .b(G815), .O(G833) );
nand2 gate289( .a(G818), .b(G819), .O(G834) );

  xor2  gate3123(.a(G821), .b(G820), .O(gate290inter0));
  nand2 gate3124(.a(gate290inter0), .b(s_368), .O(gate290inter1));
  and2  gate3125(.a(G821), .b(G820), .O(gate290inter2));
  inv1  gate3126(.a(s_368), .O(gate290inter3));
  inv1  gate3127(.a(s_369), .O(gate290inter4));
  nand2 gate3128(.a(gate290inter4), .b(gate290inter3), .O(gate290inter5));
  nor2  gate3129(.a(gate290inter5), .b(gate290inter2), .O(gate290inter6));
  inv1  gate3130(.a(G820), .O(gate290inter7));
  inv1  gate3131(.a(G821), .O(gate290inter8));
  nand2 gate3132(.a(gate290inter8), .b(gate290inter7), .O(gate290inter9));
  nand2 gate3133(.a(s_369), .b(gate290inter3), .O(gate290inter10));
  nor2  gate3134(.a(gate290inter10), .b(gate290inter9), .O(gate290inter11));
  nor2  gate3135(.a(gate290inter11), .b(gate290inter6), .O(gate290inter12));
  nand2 gate3136(.a(gate290inter12), .b(gate290inter1), .O(G847));

  xor2  gate2493(.a(G823), .b(G822), .O(gate291inter0));
  nand2 gate2494(.a(gate291inter0), .b(s_278), .O(gate291inter1));
  and2  gate2495(.a(G823), .b(G822), .O(gate291inter2));
  inv1  gate2496(.a(s_278), .O(gate291inter3));
  inv1  gate2497(.a(s_279), .O(gate291inter4));
  nand2 gate2498(.a(gate291inter4), .b(gate291inter3), .O(gate291inter5));
  nor2  gate2499(.a(gate291inter5), .b(gate291inter2), .O(gate291inter6));
  inv1  gate2500(.a(G822), .O(gate291inter7));
  inv1  gate2501(.a(G823), .O(gate291inter8));
  nand2 gate2502(.a(gate291inter8), .b(gate291inter7), .O(gate291inter9));
  nand2 gate2503(.a(s_279), .b(gate291inter3), .O(gate291inter10));
  nor2  gate2504(.a(gate291inter10), .b(gate291inter9), .O(gate291inter11));
  nor2  gate2505(.a(gate291inter11), .b(gate291inter6), .O(gate291inter12));
  nand2 gate2506(.a(gate291inter12), .b(gate291inter1), .O(G860));
nand2 gate292( .a(G824), .b(G825), .O(G873) );
nand2 gate293( .a(G828), .b(G829), .O(G886) );
nand2 gate294( .a(G832), .b(G833), .O(G899) );

  xor2  gate2997(.a(G831), .b(G830), .O(gate295inter0));
  nand2 gate2998(.a(gate295inter0), .b(s_350), .O(gate295inter1));
  and2  gate2999(.a(G831), .b(G830), .O(gate295inter2));
  inv1  gate3000(.a(s_350), .O(gate295inter3));
  inv1  gate3001(.a(s_351), .O(gate295inter4));
  nand2 gate3002(.a(gate295inter4), .b(gate295inter3), .O(gate295inter5));
  nor2  gate3003(.a(gate295inter5), .b(gate295inter2), .O(gate295inter6));
  inv1  gate3004(.a(G830), .O(gate295inter7));
  inv1  gate3005(.a(G831), .O(gate295inter8));
  nand2 gate3006(.a(gate295inter8), .b(gate295inter7), .O(gate295inter9));
  nand2 gate3007(.a(s_351), .b(gate295inter3), .O(gate295inter10));
  nor2  gate3008(.a(gate295inter10), .b(gate295inter9), .O(gate295inter11));
  nor2  gate3009(.a(gate295inter11), .b(gate295inter6), .O(gate295inter12));
  nand2 gate3010(.a(gate295inter12), .b(gate295inter1), .O(G912));
nand2 gate296( .a(G826), .b(G827), .O(G925) );
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );

  xor2  gate2731(.a(G1036), .b(G1), .O(gate387inter0));
  nand2 gate2732(.a(gate387inter0), .b(s_312), .O(gate387inter1));
  and2  gate2733(.a(G1036), .b(G1), .O(gate387inter2));
  inv1  gate2734(.a(s_312), .O(gate387inter3));
  inv1  gate2735(.a(s_313), .O(gate387inter4));
  nand2 gate2736(.a(gate387inter4), .b(gate387inter3), .O(gate387inter5));
  nor2  gate2737(.a(gate387inter5), .b(gate387inter2), .O(gate387inter6));
  inv1  gate2738(.a(G1), .O(gate387inter7));
  inv1  gate2739(.a(G1036), .O(gate387inter8));
  nand2 gate2740(.a(gate387inter8), .b(gate387inter7), .O(gate387inter9));
  nand2 gate2741(.a(s_313), .b(gate387inter3), .O(gate387inter10));
  nor2  gate2742(.a(gate387inter10), .b(gate387inter9), .O(gate387inter11));
  nor2  gate2743(.a(gate387inter11), .b(gate387inter6), .O(gate387inter12));
  nand2 gate2744(.a(gate387inter12), .b(gate387inter1), .O(G1132));

  xor2  gate3067(.a(G1039), .b(G2), .O(gate388inter0));
  nand2 gate3068(.a(gate388inter0), .b(s_360), .O(gate388inter1));
  and2  gate3069(.a(G1039), .b(G2), .O(gate388inter2));
  inv1  gate3070(.a(s_360), .O(gate388inter3));
  inv1  gate3071(.a(s_361), .O(gate388inter4));
  nand2 gate3072(.a(gate388inter4), .b(gate388inter3), .O(gate388inter5));
  nor2  gate3073(.a(gate388inter5), .b(gate388inter2), .O(gate388inter6));
  inv1  gate3074(.a(G2), .O(gate388inter7));
  inv1  gate3075(.a(G1039), .O(gate388inter8));
  nand2 gate3076(.a(gate388inter8), .b(gate388inter7), .O(gate388inter9));
  nand2 gate3077(.a(s_361), .b(gate388inter3), .O(gate388inter10));
  nor2  gate3078(.a(gate388inter10), .b(gate388inter9), .O(gate388inter11));
  nor2  gate3079(.a(gate388inter11), .b(gate388inter6), .O(gate388inter12));
  nand2 gate3080(.a(gate388inter12), .b(gate388inter1), .O(G1135));
nand2 gate389( .a(G3), .b(G1042), .O(G1138) );

  xor2  gate771(.a(G1045), .b(G4), .O(gate390inter0));
  nand2 gate772(.a(gate390inter0), .b(s_32), .O(gate390inter1));
  and2  gate773(.a(G1045), .b(G4), .O(gate390inter2));
  inv1  gate774(.a(s_32), .O(gate390inter3));
  inv1  gate775(.a(s_33), .O(gate390inter4));
  nand2 gate776(.a(gate390inter4), .b(gate390inter3), .O(gate390inter5));
  nor2  gate777(.a(gate390inter5), .b(gate390inter2), .O(gate390inter6));
  inv1  gate778(.a(G4), .O(gate390inter7));
  inv1  gate779(.a(G1045), .O(gate390inter8));
  nand2 gate780(.a(gate390inter8), .b(gate390inter7), .O(gate390inter9));
  nand2 gate781(.a(s_33), .b(gate390inter3), .O(gate390inter10));
  nor2  gate782(.a(gate390inter10), .b(gate390inter9), .O(gate390inter11));
  nor2  gate783(.a(gate390inter11), .b(gate390inter6), .O(gate390inter12));
  nand2 gate784(.a(gate390inter12), .b(gate390inter1), .O(G1141));
nand2 gate391( .a(G5), .b(G1048), .O(G1144) );

  xor2  gate2899(.a(G1051), .b(G6), .O(gate392inter0));
  nand2 gate2900(.a(gate392inter0), .b(s_336), .O(gate392inter1));
  and2  gate2901(.a(G1051), .b(G6), .O(gate392inter2));
  inv1  gate2902(.a(s_336), .O(gate392inter3));
  inv1  gate2903(.a(s_337), .O(gate392inter4));
  nand2 gate2904(.a(gate392inter4), .b(gate392inter3), .O(gate392inter5));
  nor2  gate2905(.a(gate392inter5), .b(gate392inter2), .O(gate392inter6));
  inv1  gate2906(.a(G6), .O(gate392inter7));
  inv1  gate2907(.a(G1051), .O(gate392inter8));
  nand2 gate2908(.a(gate392inter8), .b(gate392inter7), .O(gate392inter9));
  nand2 gate2909(.a(s_337), .b(gate392inter3), .O(gate392inter10));
  nor2  gate2910(.a(gate392inter10), .b(gate392inter9), .O(gate392inter11));
  nor2  gate2911(.a(gate392inter11), .b(gate392inter6), .O(gate392inter12));
  nand2 gate2912(.a(gate392inter12), .b(gate392inter1), .O(G1147));

  xor2  gate1695(.a(G1054), .b(G7), .O(gate393inter0));
  nand2 gate1696(.a(gate393inter0), .b(s_164), .O(gate393inter1));
  and2  gate1697(.a(G1054), .b(G7), .O(gate393inter2));
  inv1  gate1698(.a(s_164), .O(gate393inter3));
  inv1  gate1699(.a(s_165), .O(gate393inter4));
  nand2 gate1700(.a(gate393inter4), .b(gate393inter3), .O(gate393inter5));
  nor2  gate1701(.a(gate393inter5), .b(gate393inter2), .O(gate393inter6));
  inv1  gate1702(.a(G7), .O(gate393inter7));
  inv1  gate1703(.a(G1054), .O(gate393inter8));
  nand2 gate1704(.a(gate393inter8), .b(gate393inter7), .O(gate393inter9));
  nand2 gate1705(.a(s_165), .b(gate393inter3), .O(gate393inter10));
  nor2  gate1706(.a(gate393inter10), .b(gate393inter9), .O(gate393inter11));
  nor2  gate1707(.a(gate393inter11), .b(gate393inter6), .O(gate393inter12));
  nand2 gate1708(.a(gate393inter12), .b(gate393inter1), .O(G1150));
nand2 gate394( .a(G8), .b(G1057), .O(G1153) );
nand2 gate395( .a(G9), .b(G1060), .O(G1156) );
nand2 gate396( .a(G10), .b(G1063), .O(G1159) );
nand2 gate397( .a(G11), .b(G1066), .O(G1162) );

  xor2  gate1009(.a(G1069), .b(G12), .O(gate398inter0));
  nand2 gate1010(.a(gate398inter0), .b(s_66), .O(gate398inter1));
  and2  gate1011(.a(G1069), .b(G12), .O(gate398inter2));
  inv1  gate1012(.a(s_66), .O(gate398inter3));
  inv1  gate1013(.a(s_67), .O(gate398inter4));
  nand2 gate1014(.a(gate398inter4), .b(gate398inter3), .O(gate398inter5));
  nor2  gate1015(.a(gate398inter5), .b(gate398inter2), .O(gate398inter6));
  inv1  gate1016(.a(G12), .O(gate398inter7));
  inv1  gate1017(.a(G1069), .O(gate398inter8));
  nand2 gate1018(.a(gate398inter8), .b(gate398inter7), .O(gate398inter9));
  nand2 gate1019(.a(s_67), .b(gate398inter3), .O(gate398inter10));
  nor2  gate1020(.a(gate398inter10), .b(gate398inter9), .O(gate398inter11));
  nor2  gate1021(.a(gate398inter11), .b(gate398inter6), .O(gate398inter12));
  nand2 gate1022(.a(gate398inter12), .b(gate398inter1), .O(G1165));

  xor2  gate855(.a(G1072), .b(G13), .O(gate399inter0));
  nand2 gate856(.a(gate399inter0), .b(s_44), .O(gate399inter1));
  and2  gate857(.a(G1072), .b(G13), .O(gate399inter2));
  inv1  gate858(.a(s_44), .O(gate399inter3));
  inv1  gate859(.a(s_45), .O(gate399inter4));
  nand2 gate860(.a(gate399inter4), .b(gate399inter3), .O(gate399inter5));
  nor2  gate861(.a(gate399inter5), .b(gate399inter2), .O(gate399inter6));
  inv1  gate862(.a(G13), .O(gate399inter7));
  inv1  gate863(.a(G1072), .O(gate399inter8));
  nand2 gate864(.a(gate399inter8), .b(gate399inter7), .O(gate399inter9));
  nand2 gate865(.a(s_45), .b(gate399inter3), .O(gate399inter10));
  nor2  gate866(.a(gate399inter10), .b(gate399inter9), .O(gate399inter11));
  nor2  gate867(.a(gate399inter11), .b(gate399inter6), .O(gate399inter12));
  nand2 gate868(.a(gate399inter12), .b(gate399inter1), .O(G1168));
nand2 gate400( .a(G14), .b(G1075), .O(G1171) );
nand2 gate401( .a(G15), .b(G1078), .O(G1174) );

  xor2  gate1247(.a(G1081), .b(G16), .O(gate402inter0));
  nand2 gate1248(.a(gate402inter0), .b(s_100), .O(gate402inter1));
  and2  gate1249(.a(G1081), .b(G16), .O(gate402inter2));
  inv1  gate1250(.a(s_100), .O(gate402inter3));
  inv1  gate1251(.a(s_101), .O(gate402inter4));
  nand2 gate1252(.a(gate402inter4), .b(gate402inter3), .O(gate402inter5));
  nor2  gate1253(.a(gate402inter5), .b(gate402inter2), .O(gate402inter6));
  inv1  gate1254(.a(G16), .O(gate402inter7));
  inv1  gate1255(.a(G1081), .O(gate402inter8));
  nand2 gate1256(.a(gate402inter8), .b(gate402inter7), .O(gate402inter9));
  nand2 gate1257(.a(s_101), .b(gate402inter3), .O(gate402inter10));
  nor2  gate1258(.a(gate402inter10), .b(gate402inter9), .O(gate402inter11));
  nor2  gate1259(.a(gate402inter11), .b(gate402inter6), .O(gate402inter12));
  nand2 gate1260(.a(gate402inter12), .b(gate402inter1), .O(G1177));

  xor2  gate2241(.a(G1084), .b(G17), .O(gate403inter0));
  nand2 gate2242(.a(gate403inter0), .b(s_242), .O(gate403inter1));
  and2  gate2243(.a(G1084), .b(G17), .O(gate403inter2));
  inv1  gate2244(.a(s_242), .O(gate403inter3));
  inv1  gate2245(.a(s_243), .O(gate403inter4));
  nand2 gate2246(.a(gate403inter4), .b(gate403inter3), .O(gate403inter5));
  nor2  gate2247(.a(gate403inter5), .b(gate403inter2), .O(gate403inter6));
  inv1  gate2248(.a(G17), .O(gate403inter7));
  inv1  gate2249(.a(G1084), .O(gate403inter8));
  nand2 gate2250(.a(gate403inter8), .b(gate403inter7), .O(gate403inter9));
  nand2 gate2251(.a(s_243), .b(gate403inter3), .O(gate403inter10));
  nor2  gate2252(.a(gate403inter10), .b(gate403inter9), .O(gate403inter11));
  nor2  gate2253(.a(gate403inter11), .b(gate403inter6), .O(gate403inter12));
  nand2 gate2254(.a(gate403inter12), .b(gate403inter1), .O(G1180));
nand2 gate404( .a(G18), .b(G1087), .O(G1183) );

  xor2  gate1667(.a(G1090), .b(G19), .O(gate405inter0));
  nand2 gate1668(.a(gate405inter0), .b(s_160), .O(gate405inter1));
  and2  gate1669(.a(G1090), .b(G19), .O(gate405inter2));
  inv1  gate1670(.a(s_160), .O(gate405inter3));
  inv1  gate1671(.a(s_161), .O(gate405inter4));
  nand2 gate1672(.a(gate405inter4), .b(gate405inter3), .O(gate405inter5));
  nor2  gate1673(.a(gate405inter5), .b(gate405inter2), .O(gate405inter6));
  inv1  gate1674(.a(G19), .O(gate405inter7));
  inv1  gate1675(.a(G1090), .O(gate405inter8));
  nand2 gate1676(.a(gate405inter8), .b(gate405inter7), .O(gate405inter9));
  nand2 gate1677(.a(s_161), .b(gate405inter3), .O(gate405inter10));
  nor2  gate1678(.a(gate405inter10), .b(gate405inter9), .O(gate405inter11));
  nor2  gate1679(.a(gate405inter11), .b(gate405inter6), .O(gate405inter12));
  nand2 gate1680(.a(gate405inter12), .b(gate405inter1), .O(G1186));
nand2 gate406( .a(G20), .b(G1093), .O(G1189) );

  xor2  gate1891(.a(G1096), .b(G21), .O(gate407inter0));
  nand2 gate1892(.a(gate407inter0), .b(s_192), .O(gate407inter1));
  and2  gate1893(.a(G1096), .b(G21), .O(gate407inter2));
  inv1  gate1894(.a(s_192), .O(gate407inter3));
  inv1  gate1895(.a(s_193), .O(gate407inter4));
  nand2 gate1896(.a(gate407inter4), .b(gate407inter3), .O(gate407inter5));
  nor2  gate1897(.a(gate407inter5), .b(gate407inter2), .O(gate407inter6));
  inv1  gate1898(.a(G21), .O(gate407inter7));
  inv1  gate1899(.a(G1096), .O(gate407inter8));
  nand2 gate1900(.a(gate407inter8), .b(gate407inter7), .O(gate407inter9));
  nand2 gate1901(.a(s_193), .b(gate407inter3), .O(gate407inter10));
  nor2  gate1902(.a(gate407inter10), .b(gate407inter9), .O(gate407inter11));
  nor2  gate1903(.a(gate407inter11), .b(gate407inter6), .O(gate407inter12));
  nand2 gate1904(.a(gate407inter12), .b(gate407inter1), .O(G1192));

  xor2  gate1485(.a(G1099), .b(G22), .O(gate408inter0));
  nand2 gate1486(.a(gate408inter0), .b(s_134), .O(gate408inter1));
  and2  gate1487(.a(G1099), .b(G22), .O(gate408inter2));
  inv1  gate1488(.a(s_134), .O(gate408inter3));
  inv1  gate1489(.a(s_135), .O(gate408inter4));
  nand2 gate1490(.a(gate408inter4), .b(gate408inter3), .O(gate408inter5));
  nor2  gate1491(.a(gate408inter5), .b(gate408inter2), .O(gate408inter6));
  inv1  gate1492(.a(G22), .O(gate408inter7));
  inv1  gate1493(.a(G1099), .O(gate408inter8));
  nand2 gate1494(.a(gate408inter8), .b(gate408inter7), .O(gate408inter9));
  nand2 gate1495(.a(s_135), .b(gate408inter3), .O(gate408inter10));
  nor2  gate1496(.a(gate408inter10), .b(gate408inter9), .O(gate408inter11));
  nor2  gate1497(.a(gate408inter11), .b(gate408inter6), .O(gate408inter12));
  nand2 gate1498(.a(gate408inter12), .b(gate408inter1), .O(G1195));
nand2 gate409( .a(G23), .b(G1102), .O(G1198) );
nand2 gate410( .a(G24), .b(G1105), .O(G1201) );
nand2 gate411( .a(G25), .b(G1108), .O(G1204) );
nand2 gate412( .a(G26), .b(G1111), .O(G1207) );

  xor2  gate2955(.a(G1114), .b(G27), .O(gate413inter0));
  nand2 gate2956(.a(gate413inter0), .b(s_344), .O(gate413inter1));
  and2  gate2957(.a(G1114), .b(G27), .O(gate413inter2));
  inv1  gate2958(.a(s_344), .O(gate413inter3));
  inv1  gate2959(.a(s_345), .O(gate413inter4));
  nand2 gate2960(.a(gate413inter4), .b(gate413inter3), .O(gate413inter5));
  nor2  gate2961(.a(gate413inter5), .b(gate413inter2), .O(gate413inter6));
  inv1  gate2962(.a(G27), .O(gate413inter7));
  inv1  gate2963(.a(G1114), .O(gate413inter8));
  nand2 gate2964(.a(gate413inter8), .b(gate413inter7), .O(gate413inter9));
  nand2 gate2965(.a(s_345), .b(gate413inter3), .O(gate413inter10));
  nor2  gate2966(.a(gate413inter10), .b(gate413inter9), .O(gate413inter11));
  nor2  gate2967(.a(gate413inter11), .b(gate413inter6), .O(gate413inter12));
  nand2 gate2968(.a(gate413inter12), .b(gate413inter1), .O(G1210));
nand2 gate414( .a(G28), .b(G1117), .O(G1213) );
nand2 gate415( .a(G29), .b(G1120), .O(G1216) );
nand2 gate416( .a(G30), .b(G1123), .O(G1219) );

  xor2  gate1877(.a(G1126), .b(G31), .O(gate417inter0));
  nand2 gate1878(.a(gate417inter0), .b(s_190), .O(gate417inter1));
  and2  gate1879(.a(G1126), .b(G31), .O(gate417inter2));
  inv1  gate1880(.a(s_190), .O(gate417inter3));
  inv1  gate1881(.a(s_191), .O(gate417inter4));
  nand2 gate1882(.a(gate417inter4), .b(gate417inter3), .O(gate417inter5));
  nor2  gate1883(.a(gate417inter5), .b(gate417inter2), .O(gate417inter6));
  inv1  gate1884(.a(G31), .O(gate417inter7));
  inv1  gate1885(.a(G1126), .O(gate417inter8));
  nand2 gate1886(.a(gate417inter8), .b(gate417inter7), .O(gate417inter9));
  nand2 gate1887(.a(s_191), .b(gate417inter3), .O(gate417inter10));
  nor2  gate1888(.a(gate417inter10), .b(gate417inter9), .O(gate417inter11));
  nor2  gate1889(.a(gate417inter11), .b(gate417inter6), .O(gate417inter12));
  nand2 gate1890(.a(gate417inter12), .b(gate417inter1), .O(G1222));

  xor2  gate2157(.a(G1129), .b(G32), .O(gate418inter0));
  nand2 gate2158(.a(gate418inter0), .b(s_230), .O(gate418inter1));
  and2  gate2159(.a(G1129), .b(G32), .O(gate418inter2));
  inv1  gate2160(.a(s_230), .O(gate418inter3));
  inv1  gate2161(.a(s_231), .O(gate418inter4));
  nand2 gate2162(.a(gate418inter4), .b(gate418inter3), .O(gate418inter5));
  nor2  gate2163(.a(gate418inter5), .b(gate418inter2), .O(gate418inter6));
  inv1  gate2164(.a(G32), .O(gate418inter7));
  inv1  gate2165(.a(G1129), .O(gate418inter8));
  nand2 gate2166(.a(gate418inter8), .b(gate418inter7), .O(gate418inter9));
  nand2 gate2167(.a(s_231), .b(gate418inter3), .O(gate418inter10));
  nor2  gate2168(.a(gate418inter10), .b(gate418inter9), .O(gate418inter11));
  nor2  gate2169(.a(gate418inter11), .b(gate418inter6), .O(gate418inter12));
  nand2 gate2170(.a(gate418inter12), .b(gate418inter1), .O(G1225));

  xor2  gate2759(.a(G1132), .b(G1), .O(gate419inter0));
  nand2 gate2760(.a(gate419inter0), .b(s_316), .O(gate419inter1));
  and2  gate2761(.a(G1132), .b(G1), .O(gate419inter2));
  inv1  gate2762(.a(s_316), .O(gate419inter3));
  inv1  gate2763(.a(s_317), .O(gate419inter4));
  nand2 gate2764(.a(gate419inter4), .b(gate419inter3), .O(gate419inter5));
  nor2  gate2765(.a(gate419inter5), .b(gate419inter2), .O(gate419inter6));
  inv1  gate2766(.a(G1), .O(gate419inter7));
  inv1  gate2767(.a(G1132), .O(gate419inter8));
  nand2 gate2768(.a(gate419inter8), .b(gate419inter7), .O(gate419inter9));
  nand2 gate2769(.a(s_317), .b(gate419inter3), .O(gate419inter10));
  nor2  gate2770(.a(gate419inter10), .b(gate419inter9), .O(gate419inter11));
  nor2  gate2771(.a(gate419inter11), .b(gate419inter6), .O(gate419inter12));
  nand2 gate2772(.a(gate419inter12), .b(gate419inter1), .O(G1228));
nand2 gate420( .a(G1036), .b(G1132), .O(G1229) );

  xor2  gate645(.a(G1135), .b(G2), .O(gate421inter0));
  nand2 gate646(.a(gate421inter0), .b(s_14), .O(gate421inter1));
  and2  gate647(.a(G1135), .b(G2), .O(gate421inter2));
  inv1  gate648(.a(s_14), .O(gate421inter3));
  inv1  gate649(.a(s_15), .O(gate421inter4));
  nand2 gate650(.a(gate421inter4), .b(gate421inter3), .O(gate421inter5));
  nor2  gate651(.a(gate421inter5), .b(gate421inter2), .O(gate421inter6));
  inv1  gate652(.a(G2), .O(gate421inter7));
  inv1  gate653(.a(G1135), .O(gate421inter8));
  nand2 gate654(.a(gate421inter8), .b(gate421inter7), .O(gate421inter9));
  nand2 gate655(.a(s_15), .b(gate421inter3), .O(gate421inter10));
  nor2  gate656(.a(gate421inter10), .b(gate421inter9), .O(gate421inter11));
  nor2  gate657(.a(gate421inter11), .b(gate421inter6), .O(gate421inter12));
  nand2 gate658(.a(gate421inter12), .b(gate421inter1), .O(G1230));

  xor2  gate1681(.a(G1135), .b(G1039), .O(gate422inter0));
  nand2 gate1682(.a(gate422inter0), .b(s_162), .O(gate422inter1));
  and2  gate1683(.a(G1135), .b(G1039), .O(gate422inter2));
  inv1  gate1684(.a(s_162), .O(gate422inter3));
  inv1  gate1685(.a(s_163), .O(gate422inter4));
  nand2 gate1686(.a(gate422inter4), .b(gate422inter3), .O(gate422inter5));
  nor2  gate1687(.a(gate422inter5), .b(gate422inter2), .O(gate422inter6));
  inv1  gate1688(.a(G1039), .O(gate422inter7));
  inv1  gate1689(.a(G1135), .O(gate422inter8));
  nand2 gate1690(.a(gate422inter8), .b(gate422inter7), .O(gate422inter9));
  nand2 gate1691(.a(s_163), .b(gate422inter3), .O(gate422inter10));
  nor2  gate1692(.a(gate422inter10), .b(gate422inter9), .O(gate422inter11));
  nor2  gate1693(.a(gate422inter11), .b(gate422inter6), .O(gate422inter12));
  nand2 gate1694(.a(gate422inter12), .b(gate422inter1), .O(G1231));
nand2 gate423( .a(G3), .b(G1138), .O(G1232) );
nand2 gate424( .a(G1042), .b(G1138), .O(G1233) );

  xor2  gate2507(.a(G1141), .b(G4), .O(gate425inter0));
  nand2 gate2508(.a(gate425inter0), .b(s_280), .O(gate425inter1));
  and2  gate2509(.a(G1141), .b(G4), .O(gate425inter2));
  inv1  gate2510(.a(s_280), .O(gate425inter3));
  inv1  gate2511(.a(s_281), .O(gate425inter4));
  nand2 gate2512(.a(gate425inter4), .b(gate425inter3), .O(gate425inter5));
  nor2  gate2513(.a(gate425inter5), .b(gate425inter2), .O(gate425inter6));
  inv1  gate2514(.a(G4), .O(gate425inter7));
  inv1  gate2515(.a(G1141), .O(gate425inter8));
  nand2 gate2516(.a(gate425inter8), .b(gate425inter7), .O(gate425inter9));
  nand2 gate2517(.a(s_281), .b(gate425inter3), .O(gate425inter10));
  nor2  gate2518(.a(gate425inter10), .b(gate425inter9), .O(gate425inter11));
  nor2  gate2519(.a(gate425inter11), .b(gate425inter6), .O(gate425inter12));
  nand2 gate2520(.a(gate425inter12), .b(gate425inter1), .O(G1234));
nand2 gate426( .a(G1045), .b(G1141), .O(G1235) );

  xor2  gate897(.a(G1144), .b(G5), .O(gate427inter0));
  nand2 gate898(.a(gate427inter0), .b(s_50), .O(gate427inter1));
  and2  gate899(.a(G1144), .b(G5), .O(gate427inter2));
  inv1  gate900(.a(s_50), .O(gate427inter3));
  inv1  gate901(.a(s_51), .O(gate427inter4));
  nand2 gate902(.a(gate427inter4), .b(gate427inter3), .O(gate427inter5));
  nor2  gate903(.a(gate427inter5), .b(gate427inter2), .O(gate427inter6));
  inv1  gate904(.a(G5), .O(gate427inter7));
  inv1  gate905(.a(G1144), .O(gate427inter8));
  nand2 gate906(.a(gate427inter8), .b(gate427inter7), .O(gate427inter9));
  nand2 gate907(.a(s_51), .b(gate427inter3), .O(gate427inter10));
  nor2  gate908(.a(gate427inter10), .b(gate427inter9), .O(gate427inter11));
  nor2  gate909(.a(gate427inter11), .b(gate427inter6), .O(gate427inter12));
  nand2 gate910(.a(gate427inter12), .b(gate427inter1), .O(G1236));
nand2 gate428( .a(G1048), .b(G1144), .O(G1237) );

  xor2  gate3053(.a(G1147), .b(G6), .O(gate429inter0));
  nand2 gate3054(.a(gate429inter0), .b(s_358), .O(gate429inter1));
  and2  gate3055(.a(G1147), .b(G6), .O(gate429inter2));
  inv1  gate3056(.a(s_358), .O(gate429inter3));
  inv1  gate3057(.a(s_359), .O(gate429inter4));
  nand2 gate3058(.a(gate429inter4), .b(gate429inter3), .O(gate429inter5));
  nor2  gate3059(.a(gate429inter5), .b(gate429inter2), .O(gate429inter6));
  inv1  gate3060(.a(G6), .O(gate429inter7));
  inv1  gate3061(.a(G1147), .O(gate429inter8));
  nand2 gate3062(.a(gate429inter8), .b(gate429inter7), .O(gate429inter9));
  nand2 gate3063(.a(s_359), .b(gate429inter3), .O(gate429inter10));
  nor2  gate3064(.a(gate429inter10), .b(gate429inter9), .O(gate429inter11));
  nor2  gate3065(.a(gate429inter11), .b(gate429inter6), .O(gate429inter12));
  nand2 gate3066(.a(gate429inter12), .b(gate429inter1), .O(G1238));
nand2 gate430( .a(G1051), .b(G1147), .O(G1239) );

  xor2  gate575(.a(G1150), .b(G7), .O(gate431inter0));
  nand2 gate576(.a(gate431inter0), .b(s_4), .O(gate431inter1));
  and2  gate577(.a(G1150), .b(G7), .O(gate431inter2));
  inv1  gate578(.a(s_4), .O(gate431inter3));
  inv1  gate579(.a(s_5), .O(gate431inter4));
  nand2 gate580(.a(gate431inter4), .b(gate431inter3), .O(gate431inter5));
  nor2  gate581(.a(gate431inter5), .b(gate431inter2), .O(gate431inter6));
  inv1  gate582(.a(G7), .O(gate431inter7));
  inv1  gate583(.a(G1150), .O(gate431inter8));
  nand2 gate584(.a(gate431inter8), .b(gate431inter7), .O(gate431inter9));
  nand2 gate585(.a(s_5), .b(gate431inter3), .O(gate431inter10));
  nor2  gate586(.a(gate431inter10), .b(gate431inter9), .O(gate431inter11));
  nor2  gate587(.a(gate431inter11), .b(gate431inter6), .O(gate431inter12));
  nand2 gate588(.a(gate431inter12), .b(gate431inter1), .O(G1240));

  xor2  gate2143(.a(G1150), .b(G1054), .O(gate432inter0));
  nand2 gate2144(.a(gate432inter0), .b(s_228), .O(gate432inter1));
  and2  gate2145(.a(G1150), .b(G1054), .O(gate432inter2));
  inv1  gate2146(.a(s_228), .O(gate432inter3));
  inv1  gate2147(.a(s_229), .O(gate432inter4));
  nand2 gate2148(.a(gate432inter4), .b(gate432inter3), .O(gate432inter5));
  nor2  gate2149(.a(gate432inter5), .b(gate432inter2), .O(gate432inter6));
  inv1  gate2150(.a(G1054), .O(gate432inter7));
  inv1  gate2151(.a(G1150), .O(gate432inter8));
  nand2 gate2152(.a(gate432inter8), .b(gate432inter7), .O(gate432inter9));
  nand2 gate2153(.a(s_229), .b(gate432inter3), .O(gate432inter10));
  nor2  gate2154(.a(gate432inter10), .b(gate432inter9), .O(gate432inter11));
  nor2  gate2155(.a(gate432inter11), .b(gate432inter6), .O(gate432inter12));
  nand2 gate2156(.a(gate432inter12), .b(gate432inter1), .O(G1241));

  xor2  gate2829(.a(G1153), .b(G8), .O(gate433inter0));
  nand2 gate2830(.a(gate433inter0), .b(s_326), .O(gate433inter1));
  and2  gate2831(.a(G1153), .b(G8), .O(gate433inter2));
  inv1  gate2832(.a(s_326), .O(gate433inter3));
  inv1  gate2833(.a(s_327), .O(gate433inter4));
  nand2 gate2834(.a(gate433inter4), .b(gate433inter3), .O(gate433inter5));
  nor2  gate2835(.a(gate433inter5), .b(gate433inter2), .O(gate433inter6));
  inv1  gate2836(.a(G8), .O(gate433inter7));
  inv1  gate2837(.a(G1153), .O(gate433inter8));
  nand2 gate2838(.a(gate433inter8), .b(gate433inter7), .O(gate433inter9));
  nand2 gate2839(.a(s_327), .b(gate433inter3), .O(gate433inter10));
  nor2  gate2840(.a(gate433inter10), .b(gate433inter9), .O(gate433inter11));
  nor2  gate2841(.a(gate433inter11), .b(gate433inter6), .O(gate433inter12));
  nand2 gate2842(.a(gate433inter12), .b(gate433inter1), .O(G1242));

  xor2  gate1653(.a(G1153), .b(G1057), .O(gate434inter0));
  nand2 gate1654(.a(gate434inter0), .b(s_158), .O(gate434inter1));
  and2  gate1655(.a(G1153), .b(G1057), .O(gate434inter2));
  inv1  gate1656(.a(s_158), .O(gate434inter3));
  inv1  gate1657(.a(s_159), .O(gate434inter4));
  nand2 gate1658(.a(gate434inter4), .b(gate434inter3), .O(gate434inter5));
  nor2  gate1659(.a(gate434inter5), .b(gate434inter2), .O(gate434inter6));
  inv1  gate1660(.a(G1057), .O(gate434inter7));
  inv1  gate1661(.a(G1153), .O(gate434inter8));
  nand2 gate1662(.a(gate434inter8), .b(gate434inter7), .O(gate434inter9));
  nand2 gate1663(.a(s_159), .b(gate434inter3), .O(gate434inter10));
  nor2  gate1664(.a(gate434inter10), .b(gate434inter9), .O(gate434inter11));
  nor2  gate1665(.a(gate434inter11), .b(gate434inter6), .O(gate434inter12));
  nand2 gate1666(.a(gate434inter12), .b(gate434inter1), .O(G1243));

  xor2  gate1625(.a(G1156), .b(G9), .O(gate435inter0));
  nand2 gate1626(.a(gate435inter0), .b(s_154), .O(gate435inter1));
  and2  gate1627(.a(G1156), .b(G9), .O(gate435inter2));
  inv1  gate1628(.a(s_154), .O(gate435inter3));
  inv1  gate1629(.a(s_155), .O(gate435inter4));
  nand2 gate1630(.a(gate435inter4), .b(gate435inter3), .O(gate435inter5));
  nor2  gate1631(.a(gate435inter5), .b(gate435inter2), .O(gate435inter6));
  inv1  gate1632(.a(G9), .O(gate435inter7));
  inv1  gate1633(.a(G1156), .O(gate435inter8));
  nand2 gate1634(.a(gate435inter8), .b(gate435inter7), .O(gate435inter9));
  nand2 gate1635(.a(s_155), .b(gate435inter3), .O(gate435inter10));
  nor2  gate1636(.a(gate435inter10), .b(gate435inter9), .O(gate435inter11));
  nor2  gate1637(.a(gate435inter11), .b(gate435inter6), .O(gate435inter12));
  nand2 gate1638(.a(gate435inter12), .b(gate435inter1), .O(G1244));

  xor2  gate1569(.a(G1156), .b(G1060), .O(gate436inter0));
  nand2 gate1570(.a(gate436inter0), .b(s_146), .O(gate436inter1));
  and2  gate1571(.a(G1156), .b(G1060), .O(gate436inter2));
  inv1  gate1572(.a(s_146), .O(gate436inter3));
  inv1  gate1573(.a(s_147), .O(gate436inter4));
  nand2 gate1574(.a(gate436inter4), .b(gate436inter3), .O(gate436inter5));
  nor2  gate1575(.a(gate436inter5), .b(gate436inter2), .O(gate436inter6));
  inv1  gate1576(.a(G1060), .O(gate436inter7));
  inv1  gate1577(.a(G1156), .O(gate436inter8));
  nand2 gate1578(.a(gate436inter8), .b(gate436inter7), .O(gate436inter9));
  nand2 gate1579(.a(s_147), .b(gate436inter3), .O(gate436inter10));
  nor2  gate1580(.a(gate436inter10), .b(gate436inter9), .O(gate436inter11));
  nor2  gate1581(.a(gate436inter11), .b(gate436inter6), .O(gate436inter12));
  nand2 gate1582(.a(gate436inter12), .b(gate436inter1), .O(G1245));
nand2 gate437( .a(G10), .b(G1159), .O(G1246) );

  xor2  gate1345(.a(G1159), .b(G1063), .O(gate438inter0));
  nand2 gate1346(.a(gate438inter0), .b(s_114), .O(gate438inter1));
  and2  gate1347(.a(G1159), .b(G1063), .O(gate438inter2));
  inv1  gate1348(.a(s_114), .O(gate438inter3));
  inv1  gate1349(.a(s_115), .O(gate438inter4));
  nand2 gate1350(.a(gate438inter4), .b(gate438inter3), .O(gate438inter5));
  nor2  gate1351(.a(gate438inter5), .b(gate438inter2), .O(gate438inter6));
  inv1  gate1352(.a(G1063), .O(gate438inter7));
  inv1  gate1353(.a(G1159), .O(gate438inter8));
  nand2 gate1354(.a(gate438inter8), .b(gate438inter7), .O(gate438inter9));
  nand2 gate1355(.a(s_115), .b(gate438inter3), .O(gate438inter10));
  nor2  gate1356(.a(gate438inter10), .b(gate438inter9), .O(gate438inter11));
  nor2  gate1357(.a(gate438inter11), .b(gate438inter6), .O(gate438inter12));
  nand2 gate1358(.a(gate438inter12), .b(gate438inter1), .O(G1247));
nand2 gate439( .a(G11), .b(G1162), .O(G1248) );

  xor2  gate1779(.a(G1162), .b(G1066), .O(gate440inter0));
  nand2 gate1780(.a(gate440inter0), .b(s_176), .O(gate440inter1));
  and2  gate1781(.a(G1162), .b(G1066), .O(gate440inter2));
  inv1  gate1782(.a(s_176), .O(gate440inter3));
  inv1  gate1783(.a(s_177), .O(gate440inter4));
  nand2 gate1784(.a(gate440inter4), .b(gate440inter3), .O(gate440inter5));
  nor2  gate1785(.a(gate440inter5), .b(gate440inter2), .O(gate440inter6));
  inv1  gate1786(.a(G1066), .O(gate440inter7));
  inv1  gate1787(.a(G1162), .O(gate440inter8));
  nand2 gate1788(.a(gate440inter8), .b(gate440inter7), .O(gate440inter9));
  nand2 gate1789(.a(s_177), .b(gate440inter3), .O(gate440inter10));
  nor2  gate1790(.a(gate440inter10), .b(gate440inter9), .O(gate440inter11));
  nor2  gate1791(.a(gate440inter11), .b(gate440inter6), .O(gate440inter12));
  nand2 gate1792(.a(gate440inter12), .b(gate440inter1), .O(G1249));
nand2 gate441( .a(G12), .b(G1165), .O(G1250) );

  xor2  gate841(.a(G1165), .b(G1069), .O(gate442inter0));
  nand2 gate842(.a(gate442inter0), .b(s_42), .O(gate442inter1));
  and2  gate843(.a(G1165), .b(G1069), .O(gate442inter2));
  inv1  gate844(.a(s_42), .O(gate442inter3));
  inv1  gate845(.a(s_43), .O(gate442inter4));
  nand2 gate846(.a(gate442inter4), .b(gate442inter3), .O(gate442inter5));
  nor2  gate847(.a(gate442inter5), .b(gate442inter2), .O(gate442inter6));
  inv1  gate848(.a(G1069), .O(gate442inter7));
  inv1  gate849(.a(G1165), .O(gate442inter8));
  nand2 gate850(.a(gate442inter8), .b(gate442inter7), .O(gate442inter9));
  nand2 gate851(.a(s_43), .b(gate442inter3), .O(gate442inter10));
  nor2  gate852(.a(gate442inter10), .b(gate442inter9), .O(gate442inter11));
  nor2  gate853(.a(gate442inter11), .b(gate442inter6), .O(gate442inter12));
  nand2 gate854(.a(gate442inter12), .b(gate442inter1), .O(G1251));
nand2 gate443( .a(G13), .b(G1168), .O(G1252) );
nand2 gate444( .a(G1072), .b(G1168), .O(G1253) );
nand2 gate445( .a(G14), .b(G1171), .O(G1254) );
nand2 gate446( .a(G1075), .b(G1171), .O(G1255) );
nand2 gate447( .a(G15), .b(G1174), .O(G1256) );
nand2 gate448( .a(G1078), .b(G1174), .O(G1257) );
nand2 gate449( .a(G16), .b(G1177), .O(G1258) );
nand2 gate450( .a(G1081), .b(G1177), .O(G1259) );

  xor2  gate1023(.a(G1180), .b(G17), .O(gate451inter0));
  nand2 gate1024(.a(gate451inter0), .b(s_68), .O(gate451inter1));
  and2  gate1025(.a(G1180), .b(G17), .O(gate451inter2));
  inv1  gate1026(.a(s_68), .O(gate451inter3));
  inv1  gate1027(.a(s_69), .O(gate451inter4));
  nand2 gate1028(.a(gate451inter4), .b(gate451inter3), .O(gate451inter5));
  nor2  gate1029(.a(gate451inter5), .b(gate451inter2), .O(gate451inter6));
  inv1  gate1030(.a(G17), .O(gate451inter7));
  inv1  gate1031(.a(G1180), .O(gate451inter8));
  nand2 gate1032(.a(gate451inter8), .b(gate451inter7), .O(gate451inter9));
  nand2 gate1033(.a(s_69), .b(gate451inter3), .O(gate451inter10));
  nor2  gate1034(.a(gate451inter10), .b(gate451inter9), .O(gate451inter11));
  nor2  gate1035(.a(gate451inter11), .b(gate451inter6), .O(gate451inter12));
  nand2 gate1036(.a(gate451inter12), .b(gate451inter1), .O(G1260));
nand2 gate452( .a(G1084), .b(G1180), .O(G1261) );
nand2 gate453( .a(G18), .b(G1183), .O(G1262) );
nand2 gate454( .a(G1087), .b(G1183), .O(G1263) );
nand2 gate455( .a(G19), .b(G1186), .O(G1264) );
nand2 gate456( .a(G1090), .b(G1186), .O(G1265) );
nand2 gate457( .a(G20), .b(G1189), .O(G1266) );
nand2 gate458( .a(G1093), .b(G1189), .O(G1267) );
nand2 gate459( .a(G21), .b(G1192), .O(G1268) );
nand2 gate460( .a(G1096), .b(G1192), .O(G1269) );

  xor2  gate2927(.a(G1195), .b(G22), .O(gate461inter0));
  nand2 gate2928(.a(gate461inter0), .b(s_340), .O(gate461inter1));
  and2  gate2929(.a(G1195), .b(G22), .O(gate461inter2));
  inv1  gate2930(.a(s_340), .O(gate461inter3));
  inv1  gate2931(.a(s_341), .O(gate461inter4));
  nand2 gate2932(.a(gate461inter4), .b(gate461inter3), .O(gate461inter5));
  nor2  gate2933(.a(gate461inter5), .b(gate461inter2), .O(gate461inter6));
  inv1  gate2934(.a(G22), .O(gate461inter7));
  inv1  gate2935(.a(G1195), .O(gate461inter8));
  nand2 gate2936(.a(gate461inter8), .b(gate461inter7), .O(gate461inter9));
  nand2 gate2937(.a(s_341), .b(gate461inter3), .O(gate461inter10));
  nor2  gate2938(.a(gate461inter10), .b(gate461inter9), .O(gate461inter11));
  nor2  gate2939(.a(gate461inter11), .b(gate461inter6), .O(gate461inter12));
  nand2 gate2940(.a(gate461inter12), .b(gate461inter1), .O(G1270));

  xor2  gate729(.a(G1195), .b(G1099), .O(gate462inter0));
  nand2 gate730(.a(gate462inter0), .b(s_26), .O(gate462inter1));
  and2  gate731(.a(G1195), .b(G1099), .O(gate462inter2));
  inv1  gate732(.a(s_26), .O(gate462inter3));
  inv1  gate733(.a(s_27), .O(gate462inter4));
  nand2 gate734(.a(gate462inter4), .b(gate462inter3), .O(gate462inter5));
  nor2  gate735(.a(gate462inter5), .b(gate462inter2), .O(gate462inter6));
  inv1  gate736(.a(G1099), .O(gate462inter7));
  inv1  gate737(.a(G1195), .O(gate462inter8));
  nand2 gate738(.a(gate462inter8), .b(gate462inter7), .O(gate462inter9));
  nand2 gate739(.a(s_27), .b(gate462inter3), .O(gate462inter10));
  nor2  gate740(.a(gate462inter10), .b(gate462inter9), .O(gate462inter11));
  nor2  gate741(.a(gate462inter11), .b(gate462inter6), .O(gate462inter12));
  nand2 gate742(.a(gate462inter12), .b(gate462inter1), .O(G1271));
nand2 gate463( .a(G23), .b(G1198), .O(G1272) );

  xor2  gate2031(.a(G1198), .b(G1102), .O(gate464inter0));
  nand2 gate2032(.a(gate464inter0), .b(s_212), .O(gate464inter1));
  and2  gate2033(.a(G1198), .b(G1102), .O(gate464inter2));
  inv1  gate2034(.a(s_212), .O(gate464inter3));
  inv1  gate2035(.a(s_213), .O(gate464inter4));
  nand2 gate2036(.a(gate464inter4), .b(gate464inter3), .O(gate464inter5));
  nor2  gate2037(.a(gate464inter5), .b(gate464inter2), .O(gate464inter6));
  inv1  gate2038(.a(G1102), .O(gate464inter7));
  inv1  gate2039(.a(G1198), .O(gate464inter8));
  nand2 gate2040(.a(gate464inter8), .b(gate464inter7), .O(gate464inter9));
  nand2 gate2041(.a(s_213), .b(gate464inter3), .O(gate464inter10));
  nor2  gate2042(.a(gate464inter10), .b(gate464inter9), .O(gate464inter11));
  nor2  gate2043(.a(gate464inter11), .b(gate464inter6), .O(gate464inter12));
  nand2 gate2044(.a(gate464inter12), .b(gate464inter1), .O(G1273));

  xor2  gate2087(.a(G1201), .b(G24), .O(gate465inter0));
  nand2 gate2088(.a(gate465inter0), .b(s_220), .O(gate465inter1));
  and2  gate2089(.a(G1201), .b(G24), .O(gate465inter2));
  inv1  gate2090(.a(s_220), .O(gate465inter3));
  inv1  gate2091(.a(s_221), .O(gate465inter4));
  nand2 gate2092(.a(gate465inter4), .b(gate465inter3), .O(gate465inter5));
  nor2  gate2093(.a(gate465inter5), .b(gate465inter2), .O(gate465inter6));
  inv1  gate2094(.a(G24), .O(gate465inter7));
  inv1  gate2095(.a(G1201), .O(gate465inter8));
  nand2 gate2096(.a(gate465inter8), .b(gate465inter7), .O(gate465inter9));
  nand2 gate2097(.a(s_221), .b(gate465inter3), .O(gate465inter10));
  nor2  gate2098(.a(gate465inter10), .b(gate465inter9), .O(gate465inter11));
  nor2  gate2099(.a(gate465inter11), .b(gate465inter6), .O(gate465inter12));
  nand2 gate2100(.a(gate465inter12), .b(gate465inter1), .O(G1274));

  xor2  gate1709(.a(G1201), .b(G1105), .O(gate466inter0));
  nand2 gate1710(.a(gate466inter0), .b(s_166), .O(gate466inter1));
  and2  gate1711(.a(G1201), .b(G1105), .O(gate466inter2));
  inv1  gate1712(.a(s_166), .O(gate466inter3));
  inv1  gate1713(.a(s_167), .O(gate466inter4));
  nand2 gate1714(.a(gate466inter4), .b(gate466inter3), .O(gate466inter5));
  nor2  gate1715(.a(gate466inter5), .b(gate466inter2), .O(gate466inter6));
  inv1  gate1716(.a(G1105), .O(gate466inter7));
  inv1  gate1717(.a(G1201), .O(gate466inter8));
  nand2 gate1718(.a(gate466inter8), .b(gate466inter7), .O(gate466inter9));
  nand2 gate1719(.a(s_167), .b(gate466inter3), .O(gate466inter10));
  nor2  gate1720(.a(gate466inter10), .b(gate466inter9), .O(gate466inter11));
  nor2  gate1721(.a(gate466inter11), .b(gate466inter6), .O(gate466inter12));
  nand2 gate1722(.a(gate466inter12), .b(gate466inter1), .O(G1275));

  xor2  gate1401(.a(G1204), .b(G25), .O(gate467inter0));
  nand2 gate1402(.a(gate467inter0), .b(s_122), .O(gate467inter1));
  and2  gate1403(.a(G1204), .b(G25), .O(gate467inter2));
  inv1  gate1404(.a(s_122), .O(gate467inter3));
  inv1  gate1405(.a(s_123), .O(gate467inter4));
  nand2 gate1406(.a(gate467inter4), .b(gate467inter3), .O(gate467inter5));
  nor2  gate1407(.a(gate467inter5), .b(gate467inter2), .O(gate467inter6));
  inv1  gate1408(.a(G25), .O(gate467inter7));
  inv1  gate1409(.a(G1204), .O(gate467inter8));
  nand2 gate1410(.a(gate467inter8), .b(gate467inter7), .O(gate467inter9));
  nand2 gate1411(.a(s_123), .b(gate467inter3), .O(gate467inter10));
  nor2  gate1412(.a(gate467inter10), .b(gate467inter9), .O(gate467inter11));
  nor2  gate1413(.a(gate467inter11), .b(gate467inter6), .O(gate467inter12));
  nand2 gate1414(.a(gate467inter12), .b(gate467inter1), .O(G1276));
nand2 gate468( .a(G1108), .b(G1204), .O(G1277) );

  xor2  gate1737(.a(G1207), .b(G26), .O(gate469inter0));
  nand2 gate1738(.a(gate469inter0), .b(s_170), .O(gate469inter1));
  and2  gate1739(.a(G1207), .b(G26), .O(gate469inter2));
  inv1  gate1740(.a(s_170), .O(gate469inter3));
  inv1  gate1741(.a(s_171), .O(gate469inter4));
  nand2 gate1742(.a(gate469inter4), .b(gate469inter3), .O(gate469inter5));
  nor2  gate1743(.a(gate469inter5), .b(gate469inter2), .O(gate469inter6));
  inv1  gate1744(.a(G26), .O(gate469inter7));
  inv1  gate1745(.a(G1207), .O(gate469inter8));
  nand2 gate1746(.a(gate469inter8), .b(gate469inter7), .O(gate469inter9));
  nand2 gate1747(.a(s_171), .b(gate469inter3), .O(gate469inter10));
  nor2  gate1748(.a(gate469inter10), .b(gate469inter9), .O(gate469inter11));
  nor2  gate1749(.a(gate469inter11), .b(gate469inter6), .O(gate469inter12));
  nand2 gate1750(.a(gate469inter12), .b(gate469inter1), .O(G1278));

  xor2  gate1219(.a(G1207), .b(G1111), .O(gate470inter0));
  nand2 gate1220(.a(gate470inter0), .b(s_96), .O(gate470inter1));
  and2  gate1221(.a(G1207), .b(G1111), .O(gate470inter2));
  inv1  gate1222(.a(s_96), .O(gate470inter3));
  inv1  gate1223(.a(s_97), .O(gate470inter4));
  nand2 gate1224(.a(gate470inter4), .b(gate470inter3), .O(gate470inter5));
  nor2  gate1225(.a(gate470inter5), .b(gate470inter2), .O(gate470inter6));
  inv1  gate1226(.a(G1111), .O(gate470inter7));
  inv1  gate1227(.a(G1207), .O(gate470inter8));
  nand2 gate1228(.a(gate470inter8), .b(gate470inter7), .O(gate470inter9));
  nand2 gate1229(.a(s_97), .b(gate470inter3), .O(gate470inter10));
  nor2  gate1230(.a(gate470inter10), .b(gate470inter9), .O(gate470inter11));
  nor2  gate1231(.a(gate470inter11), .b(gate470inter6), .O(gate470inter12));
  nand2 gate1232(.a(gate470inter12), .b(gate470inter1), .O(G1279));

  xor2  gate1093(.a(G1210), .b(G27), .O(gate471inter0));
  nand2 gate1094(.a(gate471inter0), .b(s_78), .O(gate471inter1));
  and2  gate1095(.a(G1210), .b(G27), .O(gate471inter2));
  inv1  gate1096(.a(s_78), .O(gate471inter3));
  inv1  gate1097(.a(s_79), .O(gate471inter4));
  nand2 gate1098(.a(gate471inter4), .b(gate471inter3), .O(gate471inter5));
  nor2  gate1099(.a(gate471inter5), .b(gate471inter2), .O(gate471inter6));
  inv1  gate1100(.a(G27), .O(gate471inter7));
  inv1  gate1101(.a(G1210), .O(gate471inter8));
  nand2 gate1102(.a(gate471inter8), .b(gate471inter7), .O(gate471inter9));
  nand2 gate1103(.a(s_79), .b(gate471inter3), .O(gate471inter10));
  nor2  gate1104(.a(gate471inter10), .b(gate471inter9), .O(gate471inter11));
  nor2  gate1105(.a(gate471inter11), .b(gate471inter6), .O(gate471inter12));
  nand2 gate1106(.a(gate471inter12), .b(gate471inter1), .O(G1280));
nand2 gate472( .a(G1114), .b(G1210), .O(G1281) );

  xor2  gate1905(.a(G1213), .b(G28), .O(gate473inter0));
  nand2 gate1906(.a(gate473inter0), .b(s_194), .O(gate473inter1));
  and2  gate1907(.a(G1213), .b(G28), .O(gate473inter2));
  inv1  gate1908(.a(s_194), .O(gate473inter3));
  inv1  gate1909(.a(s_195), .O(gate473inter4));
  nand2 gate1910(.a(gate473inter4), .b(gate473inter3), .O(gate473inter5));
  nor2  gate1911(.a(gate473inter5), .b(gate473inter2), .O(gate473inter6));
  inv1  gate1912(.a(G28), .O(gate473inter7));
  inv1  gate1913(.a(G1213), .O(gate473inter8));
  nand2 gate1914(.a(gate473inter8), .b(gate473inter7), .O(gate473inter9));
  nand2 gate1915(.a(s_195), .b(gate473inter3), .O(gate473inter10));
  nor2  gate1916(.a(gate473inter10), .b(gate473inter9), .O(gate473inter11));
  nor2  gate1917(.a(gate473inter11), .b(gate473inter6), .O(gate473inter12));
  nand2 gate1918(.a(gate473inter12), .b(gate473inter1), .O(G1282));

  xor2  gate2773(.a(G1213), .b(G1117), .O(gate474inter0));
  nand2 gate2774(.a(gate474inter0), .b(s_318), .O(gate474inter1));
  and2  gate2775(.a(G1213), .b(G1117), .O(gate474inter2));
  inv1  gate2776(.a(s_318), .O(gate474inter3));
  inv1  gate2777(.a(s_319), .O(gate474inter4));
  nand2 gate2778(.a(gate474inter4), .b(gate474inter3), .O(gate474inter5));
  nor2  gate2779(.a(gate474inter5), .b(gate474inter2), .O(gate474inter6));
  inv1  gate2780(.a(G1117), .O(gate474inter7));
  inv1  gate2781(.a(G1213), .O(gate474inter8));
  nand2 gate2782(.a(gate474inter8), .b(gate474inter7), .O(gate474inter9));
  nand2 gate2783(.a(s_319), .b(gate474inter3), .O(gate474inter10));
  nor2  gate2784(.a(gate474inter10), .b(gate474inter9), .O(gate474inter11));
  nor2  gate2785(.a(gate474inter11), .b(gate474inter6), .O(gate474inter12));
  nand2 gate2786(.a(gate474inter12), .b(gate474inter1), .O(G1283));

  xor2  gate2549(.a(G1216), .b(G29), .O(gate475inter0));
  nand2 gate2550(.a(gate475inter0), .b(s_286), .O(gate475inter1));
  and2  gate2551(.a(G1216), .b(G29), .O(gate475inter2));
  inv1  gate2552(.a(s_286), .O(gate475inter3));
  inv1  gate2553(.a(s_287), .O(gate475inter4));
  nand2 gate2554(.a(gate475inter4), .b(gate475inter3), .O(gate475inter5));
  nor2  gate2555(.a(gate475inter5), .b(gate475inter2), .O(gate475inter6));
  inv1  gate2556(.a(G29), .O(gate475inter7));
  inv1  gate2557(.a(G1216), .O(gate475inter8));
  nand2 gate2558(.a(gate475inter8), .b(gate475inter7), .O(gate475inter9));
  nand2 gate2559(.a(s_287), .b(gate475inter3), .O(gate475inter10));
  nor2  gate2560(.a(gate475inter10), .b(gate475inter9), .O(gate475inter11));
  nor2  gate2561(.a(gate475inter11), .b(gate475inter6), .O(gate475inter12));
  nand2 gate2562(.a(gate475inter12), .b(gate475inter1), .O(G1284));
nand2 gate476( .a(G1120), .b(G1216), .O(G1285) );
nand2 gate477( .a(G30), .b(G1219), .O(G1286) );

  xor2  gate2129(.a(G1219), .b(G1123), .O(gate478inter0));
  nand2 gate2130(.a(gate478inter0), .b(s_226), .O(gate478inter1));
  and2  gate2131(.a(G1219), .b(G1123), .O(gate478inter2));
  inv1  gate2132(.a(s_226), .O(gate478inter3));
  inv1  gate2133(.a(s_227), .O(gate478inter4));
  nand2 gate2134(.a(gate478inter4), .b(gate478inter3), .O(gate478inter5));
  nor2  gate2135(.a(gate478inter5), .b(gate478inter2), .O(gate478inter6));
  inv1  gate2136(.a(G1123), .O(gate478inter7));
  inv1  gate2137(.a(G1219), .O(gate478inter8));
  nand2 gate2138(.a(gate478inter8), .b(gate478inter7), .O(gate478inter9));
  nand2 gate2139(.a(s_227), .b(gate478inter3), .O(gate478inter10));
  nor2  gate2140(.a(gate478inter10), .b(gate478inter9), .O(gate478inter11));
  nor2  gate2141(.a(gate478inter11), .b(gate478inter6), .O(gate478inter12));
  nand2 gate2142(.a(gate478inter12), .b(gate478inter1), .O(G1287));
nand2 gate479( .a(G31), .b(G1222), .O(G1288) );
nand2 gate480( .a(G1126), .b(G1222), .O(G1289) );
nand2 gate481( .a(G32), .b(G1225), .O(G1290) );
nand2 gate482( .a(G1129), .b(G1225), .O(G1291) );

  xor2  gate2633(.a(G1229), .b(G1228), .O(gate483inter0));
  nand2 gate2634(.a(gate483inter0), .b(s_298), .O(gate483inter1));
  and2  gate2635(.a(G1229), .b(G1228), .O(gate483inter2));
  inv1  gate2636(.a(s_298), .O(gate483inter3));
  inv1  gate2637(.a(s_299), .O(gate483inter4));
  nand2 gate2638(.a(gate483inter4), .b(gate483inter3), .O(gate483inter5));
  nor2  gate2639(.a(gate483inter5), .b(gate483inter2), .O(gate483inter6));
  inv1  gate2640(.a(G1228), .O(gate483inter7));
  inv1  gate2641(.a(G1229), .O(gate483inter8));
  nand2 gate2642(.a(gate483inter8), .b(gate483inter7), .O(gate483inter9));
  nand2 gate2643(.a(s_299), .b(gate483inter3), .O(gate483inter10));
  nor2  gate2644(.a(gate483inter10), .b(gate483inter9), .O(gate483inter11));
  nor2  gate2645(.a(gate483inter11), .b(gate483inter6), .O(gate483inter12));
  nand2 gate2646(.a(gate483inter12), .b(gate483inter1), .O(G1292));
nand2 gate484( .a(G1230), .b(G1231), .O(G1293) );

  xor2  gate3095(.a(G1233), .b(G1232), .O(gate485inter0));
  nand2 gate3096(.a(gate485inter0), .b(s_364), .O(gate485inter1));
  and2  gate3097(.a(G1233), .b(G1232), .O(gate485inter2));
  inv1  gate3098(.a(s_364), .O(gate485inter3));
  inv1  gate3099(.a(s_365), .O(gate485inter4));
  nand2 gate3100(.a(gate485inter4), .b(gate485inter3), .O(gate485inter5));
  nor2  gate3101(.a(gate485inter5), .b(gate485inter2), .O(gate485inter6));
  inv1  gate3102(.a(G1232), .O(gate485inter7));
  inv1  gate3103(.a(G1233), .O(gate485inter8));
  nand2 gate3104(.a(gate485inter8), .b(gate485inter7), .O(gate485inter9));
  nand2 gate3105(.a(s_365), .b(gate485inter3), .O(gate485inter10));
  nor2  gate3106(.a(gate485inter10), .b(gate485inter9), .O(gate485inter11));
  nor2  gate3107(.a(gate485inter11), .b(gate485inter6), .O(gate485inter12));
  nand2 gate3108(.a(gate485inter12), .b(gate485inter1), .O(G1294));
nand2 gate486( .a(G1234), .b(G1235), .O(G1295) );
nand2 gate487( .a(G1236), .b(G1237), .O(G1296) );
nand2 gate488( .a(G1238), .b(G1239), .O(G1297) );

  xor2  gate2815(.a(G1241), .b(G1240), .O(gate489inter0));
  nand2 gate2816(.a(gate489inter0), .b(s_324), .O(gate489inter1));
  and2  gate2817(.a(G1241), .b(G1240), .O(gate489inter2));
  inv1  gate2818(.a(s_324), .O(gate489inter3));
  inv1  gate2819(.a(s_325), .O(gate489inter4));
  nand2 gate2820(.a(gate489inter4), .b(gate489inter3), .O(gate489inter5));
  nor2  gate2821(.a(gate489inter5), .b(gate489inter2), .O(gate489inter6));
  inv1  gate2822(.a(G1240), .O(gate489inter7));
  inv1  gate2823(.a(G1241), .O(gate489inter8));
  nand2 gate2824(.a(gate489inter8), .b(gate489inter7), .O(gate489inter9));
  nand2 gate2825(.a(s_325), .b(gate489inter3), .O(gate489inter10));
  nor2  gate2826(.a(gate489inter10), .b(gate489inter9), .O(gate489inter11));
  nor2  gate2827(.a(gate489inter11), .b(gate489inter6), .O(gate489inter12));
  nand2 gate2828(.a(gate489inter12), .b(gate489inter1), .O(G1298));
nand2 gate490( .a(G1242), .b(G1243), .O(G1299) );

  xor2  gate2703(.a(G1245), .b(G1244), .O(gate491inter0));
  nand2 gate2704(.a(gate491inter0), .b(s_308), .O(gate491inter1));
  and2  gate2705(.a(G1245), .b(G1244), .O(gate491inter2));
  inv1  gate2706(.a(s_308), .O(gate491inter3));
  inv1  gate2707(.a(s_309), .O(gate491inter4));
  nand2 gate2708(.a(gate491inter4), .b(gate491inter3), .O(gate491inter5));
  nor2  gate2709(.a(gate491inter5), .b(gate491inter2), .O(gate491inter6));
  inv1  gate2710(.a(G1244), .O(gate491inter7));
  inv1  gate2711(.a(G1245), .O(gate491inter8));
  nand2 gate2712(.a(gate491inter8), .b(gate491inter7), .O(gate491inter9));
  nand2 gate2713(.a(s_309), .b(gate491inter3), .O(gate491inter10));
  nor2  gate2714(.a(gate491inter10), .b(gate491inter9), .O(gate491inter11));
  nor2  gate2715(.a(gate491inter11), .b(gate491inter6), .O(gate491inter12));
  nand2 gate2716(.a(gate491inter12), .b(gate491inter1), .O(G1300));
nand2 gate492( .a(G1246), .b(G1247), .O(G1301) );

  xor2  gate1639(.a(G1249), .b(G1248), .O(gate493inter0));
  nand2 gate1640(.a(gate493inter0), .b(s_156), .O(gate493inter1));
  and2  gate1641(.a(G1249), .b(G1248), .O(gate493inter2));
  inv1  gate1642(.a(s_156), .O(gate493inter3));
  inv1  gate1643(.a(s_157), .O(gate493inter4));
  nand2 gate1644(.a(gate493inter4), .b(gate493inter3), .O(gate493inter5));
  nor2  gate1645(.a(gate493inter5), .b(gate493inter2), .O(gate493inter6));
  inv1  gate1646(.a(G1248), .O(gate493inter7));
  inv1  gate1647(.a(G1249), .O(gate493inter8));
  nand2 gate1648(.a(gate493inter8), .b(gate493inter7), .O(gate493inter9));
  nand2 gate1649(.a(s_157), .b(gate493inter3), .O(gate493inter10));
  nor2  gate1650(.a(gate493inter10), .b(gate493inter9), .O(gate493inter11));
  nor2  gate1651(.a(gate493inter11), .b(gate493inter6), .O(gate493inter12));
  nand2 gate1652(.a(gate493inter12), .b(gate493inter1), .O(G1302));
nand2 gate494( .a(G1250), .b(G1251), .O(G1303) );

  xor2  gate743(.a(G1253), .b(G1252), .O(gate495inter0));
  nand2 gate744(.a(gate495inter0), .b(s_28), .O(gate495inter1));
  and2  gate745(.a(G1253), .b(G1252), .O(gate495inter2));
  inv1  gate746(.a(s_28), .O(gate495inter3));
  inv1  gate747(.a(s_29), .O(gate495inter4));
  nand2 gate748(.a(gate495inter4), .b(gate495inter3), .O(gate495inter5));
  nor2  gate749(.a(gate495inter5), .b(gate495inter2), .O(gate495inter6));
  inv1  gate750(.a(G1252), .O(gate495inter7));
  inv1  gate751(.a(G1253), .O(gate495inter8));
  nand2 gate752(.a(gate495inter8), .b(gate495inter7), .O(gate495inter9));
  nand2 gate753(.a(s_29), .b(gate495inter3), .O(gate495inter10));
  nor2  gate754(.a(gate495inter10), .b(gate495inter9), .O(gate495inter11));
  nor2  gate755(.a(gate495inter11), .b(gate495inter6), .O(gate495inter12));
  nand2 gate756(.a(gate495inter12), .b(gate495inter1), .O(G1304));

  xor2  gate603(.a(G1255), .b(G1254), .O(gate496inter0));
  nand2 gate604(.a(gate496inter0), .b(s_8), .O(gate496inter1));
  and2  gate605(.a(G1255), .b(G1254), .O(gate496inter2));
  inv1  gate606(.a(s_8), .O(gate496inter3));
  inv1  gate607(.a(s_9), .O(gate496inter4));
  nand2 gate608(.a(gate496inter4), .b(gate496inter3), .O(gate496inter5));
  nor2  gate609(.a(gate496inter5), .b(gate496inter2), .O(gate496inter6));
  inv1  gate610(.a(G1254), .O(gate496inter7));
  inv1  gate611(.a(G1255), .O(gate496inter8));
  nand2 gate612(.a(gate496inter8), .b(gate496inter7), .O(gate496inter9));
  nand2 gate613(.a(s_9), .b(gate496inter3), .O(gate496inter10));
  nor2  gate614(.a(gate496inter10), .b(gate496inter9), .O(gate496inter11));
  nor2  gate615(.a(gate496inter11), .b(gate496inter6), .O(gate496inter12));
  nand2 gate616(.a(gate496inter12), .b(gate496inter1), .O(G1305));
nand2 gate497( .a(G1256), .b(G1257), .O(G1306) );
nand2 gate498( .a(G1258), .b(G1259), .O(G1307) );

  xor2  gate2647(.a(G1261), .b(G1260), .O(gate499inter0));
  nand2 gate2648(.a(gate499inter0), .b(s_300), .O(gate499inter1));
  and2  gate2649(.a(G1261), .b(G1260), .O(gate499inter2));
  inv1  gate2650(.a(s_300), .O(gate499inter3));
  inv1  gate2651(.a(s_301), .O(gate499inter4));
  nand2 gate2652(.a(gate499inter4), .b(gate499inter3), .O(gate499inter5));
  nor2  gate2653(.a(gate499inter5), .b(gate499inter2), .O(gate499inter6));
  inv1  gate2654(.a(G1260), .O(gate499inter7));
  inv1  gate2655(.a(G1261), .O(gate499inter8));
  nand2 gate2656(.a(gate499inter8), .b(gate499inter7), .O(gate499inter9));
  nand2 gate2657(.a(s_301), .b(gate499inter3), .O(gate499inter10));
  nor2  gate2658(.a(gate499inter10), .b(gate499inter9), .O(gate499inter11));
  nor2  gate2659(.a(gate499inter11), .b(gate499inter6), .O(gate499inter12));
  nand2 gate2660(.a(gate499inter12), .b(gate499inter1), .O(G1308));
nand2 gate500( .a(G1262), .b(G1263), .O(G1309) );

  xor2  gate799(.a(G1265), .b(G1264), .O(gate501inter0));
  nand2 gate800(.a(gate501inter0), .b(s_36), .O(gate501inter1));
  and2  gate801(.a(G1265), .b(G1264), .O(gate501inter2));
  inv1  gate802(.a(s_36), .O(gate501inter3));
  inv1  gate803(.a(s_37), .O(gate501inter4));
  nand2 gate804(.a(gate501inter4), .b(gate501inter3), .O(gate501inter5));
  nor2  gate805(.a(gate501inter5), .b(gate501inter2), .O(gate501inter6));
  inv1  gate806(.a(G1264), .O(gate501inter7));
  inv1  gate807(.a(G1265), .O(gate501inter8));
  nand2 gate808(.a(gate501inter8), .b(gate501inter7), .O(gate501inter9));
  nand2 gate809(.a(s_37), .b(gate501inter3), .O(gate501inter10));
  nor2  gate810(.a(gate501inter10), .b(gate501inter9), .O(gate501inter11));
  nor2  gate811(.a(gate501inter11), .b(gate501inter6), .O(gate501inter12));
  nand2 gate812(.a(gate501inter12), .b(gate501inter1), .O(G1310));

  xor2  gate1499(.a(G1267), .b(G1266), .O(gate502inter0));
  nand2 gate1500(.a(gate502inter0), .b(s_136), .O(gate502inter1));
  and2  gate1501(.a(G1267), .b(G1266), .O(gate502inter2));
  inv1  gate1502(.a(s_136), .O(gate502inter3));
  inv1  gate1503(.a(s_137), .O(gate502inter4));
  nand2 gate1504(.a(gate502inter4), .b(gate502inter3), .O(gate502inter5));
  nor2  gate1505(.a(gate502inter5), .b(gate502inter2), .O(gate502inter6));
  inv1  gate1506(.a(G1266), .O(gate502inter7));
  inv1  gate1507(.a(G1267), .O(gate502inter8));
  nand2 gate1508(.a(gate502inter8), .b(gate502inter7), .O(gate502inter9));
  nand2 gate1509(.a(s_137), .b(gate502inter3), .O(gate502inter10));
  nor2  gate1510(.a(gate502inter10), .b(gate502inter9), .O(gate502inter11));
  nor2  gate1511(.a(gate502inter11), .b(gate502inter6), .O(gate502inter12));
  nand2 gate1512(.a(gate502inter12), .b(gate502inter1), .O(G1311));
nand2 gate503( .a(G1268), .b(G1269), .O(G1312) );
nand2 gate504( .a(G1270), .b(G1271), .O(G1313) );
nand2 gate505( .a(G1272), .b(G1273), .O(G1314) );
nand2 gate506( .a(G1274), .b(G1275), .O(G1315) );
nand2 gate507( .a(G1276), .b(G1277), .O(G1316) );

  xor2  gate1583(.a(G1279), .b(G1278), .O(gate508inter0));
  nand2 gate1584(.a(gate508inter0), .b(s_148), .O(gate508inter1));
  and2  gate1585(.a(G1279), .b(G1278), .O(gate508inter2));
  inv1  gate1586(.a(s_148), .O(gate508inter3));
  inv1  gate1587(.a(s_149), .O(gate508inter4));
  nand2 gate1588(.a(gate508inter4), .b(gate508inter3), .O(gate508inter5));
  nor2  gate1589(.a(gate508inter5), .b(gate508inter2), .O(gate508inter6));
  inv1  gate1590(.a(G1278), .O(gate508inter7));
  inv1  gate1591(.a(G1279), .O(gate508inter8));
  nand2 gate1592(.a(gate508inter8), .b(gate508inter7), .O(gate508inter9));
  nand2 gate1593(.a(s_149), .b(gate508inter3), .O(gate508inter10));
  nor2  gate1594(.a(gate508inter10), .b(gate508inter9), .O(gate508inter11));
  nor2  gate1595(.a(gate508inter11), .b(gate508inter6), .O(gate508inter12));
  nand2 gate1596(.a(gate508inter12), .b(gate508inter1), .O(G1317));

  xor2  gate2255(.a(G1281), .b(G1280), .O(gate509inter0));
  nand2 gate2256(.a(gate509inter0), .b(s_244), .O(gate509inter1));
  and2  gate2257(.a(G1281), .b(G1280), .O(gate509inter2));
  inv1  gate2258(.a(s_244), .O(gate509inter3));
  inv1  gate2259(.a(s_245), .O(gate509inter4));
  nand2 gate2260(.a(gate509inter4), .b(gate509inter3), .O(gate509inter5));
  nor2  gate2261(.a(gate509inter5), .b(gate509inter2), .O(gate509inter6));
  inv1  gate2262(.a(G1280), .O(gate509inter7));
  inv1  gate2263(.a(G1281), .O(gate509inter8));
  nand2 gate2264(.a(gate509inter8), .b(gate509inter7), .O(gate509inter9));
  nand2 gate2265(.a(s_245), .b(gate509inter3), .O(gate509inter10));
  nor2  gate2266(.a(gate509inter10), .b(gate509inter9), .O(gate509inter11));
  nor2  gate2267(.a(gate509inter11), .b(gate509inter6), .O(gate509inter12));
  nand2 gate2268(.a(gate509inter12), .b(gate509inter1), .O(G1318));
nand2 gate510( .a(G1282), .b(G1283), .O(G1319) );

  xor2  gate1807(.a(G1285), .b(G1284), .O(gate511inter0));
  nand2 gate1808(.a(gate511inter0), .b(s_180), .O(gate511inter1));
  and2  gate1809(.a(G1285), .b(G1284), .O(gate511inter2));
  inv1  gate1810(.a(s_180), .O(gate511inter3));
  inv1  gate1811(.a(s_181), .O(gate511inter4));
  nand2 gate1812(.a(gate511inter4), .b(gate511inter3), .O(gate511inter5));
  nor2  gate1813(.a(gate511inter5), .b(gate511inter2), .O(gate511inter6));
  inv1  gate1814(.a(G1284), .O(gate511inter7));
  inv1  gate1815(.a(G1285), .O(gate511inter8));
  nand2 gate1816(.a(gate511inter8), .b(gate511inter7), .O(gate511inter9));
  nand2 gate1817(.a(s_181), .b(gate511inter3), .O(gate511inter10));
  nor2  gate1818(.a(gate511inter10), .b(gate511inter9), .O(gate511inter11));
  nor2  gate1819(.a(gate511inter11), .b(gate511inter6), .O(gate511inter12));
  nand2 gate1820(.a(gate511inter12), .b(gate511inter1), .O(G1320));

  xor2  gate1191(.a(G1287), .b(G1286), .O(gate512inter0));
  nand2 gate1192(.a(gate512inter0), .b(s_92), .O(gate512inter1));
  and2  gate1193(.a(G1287), .b(G1286), .O(gate512inter2));
  inv1  gate1194(.a(s_92), .O(gate512inter3));
  inv1  gate1195(.a(s_93), .O(gate512inter4));
  nand2 gate1196(.a(gate512inter4), .b(gate512inter3), .O(gate512inter5));
  nor2  gate1197(.a(gate512inter5), .b(gate512inter2), .O(gate512inter6));
  inv1  gate1198(.a(G1286), .O(gate512inter7));
  inv1  gate1199(.a(G1287), .O(gate512inter8));
  nand2 gate1200(.a(gate512inter8), .b(gate512inter7), .O(gate512inter9));
  nand2 gate1201(.a(s_93), .b(gate512inter3), .O(gate512inter10));
  nor2  gate1202(.a(gate512inter10), .b(gate512inter9), .O(gate512inter11));
  nor2  gate1203(.a(gate512inter11), .b(gate512inter6), .O(gate512inter12));
  nand2 gate1204(.a(gate512inter12), .b(gate512inter1), .O(G1321));
nand2 gate513( .a(G1288), .b(G1289), .O(G1322) );
nand2 gate514( .a(G1290), .b(G1291), .O(G1323) );
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule