module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);

input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;//RE__PI;

input s_0,s_1;//RE__ALLOW(00,01,10,11);
input s_2,s_3;//RE__ALLOW(00,01,10,11);
input s_4,s_5;//RE__ALLOW(00,01,10,11);
input s_6,s_7;//RE__ALLOW(00,01,10,11);
input s_8,s_9;//RE__ALLOW(00,01,10,11);
input s_10,s_11;//RE__ALLOW(00,01,10,11);
input s_12,s_13;//RE__ALLOW(00,01,10,11);
input s_14,s_15;//RE__ALLOW(00,01,10,11);
input s_16,s_17;//RE__ALLOW(00,01,10,11);
input s_18,s_19;//RE__ALLOW(00,01,10,11);
input s_20,s_21;//RE__ALLOW(00,01,10,11);
input s_22,s_23;//RE__ALLOW(00,01,10,11);
input s_24,s_25;//RE__ALLOW(00,01,10,11);
input s_26,s_27;//RE__ALLOW(00,01,10,11);
input s_28,s_29;//RE__ALLOW(00,01,10,11);
input s_30,s_31;//RE__ALLOW(00,01,10,11);
input s_32,s_33;//RE__ALLOW(00,01,10,11);
input s_34,s_35;//RE__ALLOW(00,01,10,11);
input s_36,s_37;//RE__ALLOW(00,01,10,11);
input s_38,s_39;//RE__ALLOW(00,01,10,11);
input s_40,s_41;//RE__ALLOW(00,01,10,11);
input s_42,s_43;//RE__ALLOW(00,01,10,11);
input s_44,s_45;//RE__ALLOW(00,01,10,11);
input s_46,s_47;//RE__ALLOW(00,01,10,11);
input s_48,s_49;//RE__ALLOW(00,01,10,11);
input s_50,s_51;//RE__ALLOW(00,01,10,11);
input s_52,s_53;//RE__ALLOW(00,01,10,11);
input s_54,s_55;//RE__ALLOW(00,01,10,11);
input s_56,s_57;//RE__ALLOW(00,01,10,11);
input s_58,s_59;//RE__ALLOW(00,01,10,11);
input s_60,s_61;//RE__ALLOW(00,01,10,11);
input s_62,s_63;//RE__ALLOW(00,01,10,11);
input s_64,s_65;//RE__ALLOW(00,01,10,11);
input s_66,s_67;//RE__ALLOW(00,01,10,11);
input s_68,s_69;//RE__ALLOW(00,01,10,11);
input s_70,s_71;//RE__ALLOW(00,01,10,11);
input s_72,s_73;//RE__ALLOW(00,01,10,11);
input s_74,s_75;//RE__ALLOW(00,01,10,11);
input s_76,s_77;//RE__ALLOW(00,01,10,11);
input s_78,s_79;//RE__ALLOW(00,01,10,11);
input s_80,s_81;//RE__ALLOW(00,01,10,11);
input s_82,s_83;//RE__ALLOW(00,01,10,11);
input s_84,s_85;//RE__ALLOW(00,01,10,11);
input s_86,s_87;//RE__ALLOW(00,01,10,11);
input s_88,s_89;//RE__ALLOW(00,01,10,11);
input s_90,s_91;//RE__ALLOW(00,01,10,11);
input s_92,s_93;//RE__ALLOW(00,01,10,11);
input s_94,s_95;//RE__ALLOW(00,01,10,11);
input s_96,s_97;//RE__ALLOW(00,01,10,11);
input s_98,s_99;//RE__ALLOW(00,01,10,11);
input s_100,s_101;//RE__ALLOW(00,01,10,11);
input s_102,s_103;//RE__ALLOW(00,01,10,11);
input s_104,s_105;//RE__ALLOW(00,01,10,11);
input s_106,s_107;//RE__ALLOW(00,01,10,11);
input s_108,s_109;//RE__ALLOW(00,01,10,11);
input s_110,s_111;//RE__ALLOW(00,01,10,11);
input s_112,s_113;//RE__ALLOW(00,01,10,11);
input s_114,s_115;//RE__ALLOW(00,01,10,11);
input s_116,s_117;//RE__ALLOW(00,01,10,11);
input s_118,s_119;//RE__ALLOW(00,01,10,11);
input s_120,s_121;//RE__ALLOW(00,01,10,11);
input s_122,s_123;//RE__ALLOW(00,01,10,11);
input s_124,s_125;//RE__ALLOW(00,01,10,11);
input s_126,s_127;//RE__ALLOW(00,01,10,11);
input s_128,s_129;//RE__ALLOW(00,01,10,11);
input s_130,s_131;//RE__ALLOW(00,01,10,11);
input s_132,s_133;//RE__ALLOW(00,01,10,11);
input s_134,s_135;//RE__ALLOW(00,01,10,11);
input s_136,s_137;//RE__ALLOW(00,01,10,11);
input s_138,s_139;//RE__ALLOW(00,01,10,11);
input s_140,s_141;//RE__ALLOW(00,01,10,11);
input s_142,s_143;//RE__ALLOW(00,01,10,11);
input s_144,s_145;//RE__ALLOW(00,01,10,11);
input s_146,s_147;//RE__ALLOW(00,01,10,11);
input s_148,s_149;//RE__ALLOW(00,01,10,11);
input s_150,s_151;//RE__ALLOW(00,01,10,11);
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;

  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate263inter0, gate263inter1, gate263inter2, gate263inter3, gate263inter4, gate263inter5, gate263inter6, gate263inter7, gate263inter8, gate263inter9, gate263inter10, gate263inter11, gate263inter12, gate120inter0, gate120inter1, gate120inter2, gate120inter3, gate120inter4, gate120inter5, gate120inter6, gate120inter7, gate120inter8, gate120inter9, gate120inter10, gate120inter11, gate120inter12, gate407inter0, gate407inter1, gate407inter2, gate407inter3, gate407inter4, gate407inter5, gate407inter6, gate407inter7, gate407inter8, gate407inter9, gate407inter10, gate407inter11, gate407inter12, gate462inter0, gate462inter1, gate462inter2, gate462inter3, gate462inter4, gate462inter5, gate462inter6, gate462inter7, gate462inter8, gate462inter9, gate462inter10, gate462inter11, gate462inter12, gate148inter0, gate148inter1, gate148inter2, gate148inter3, gate148inter4, gate148inter5, gate148inter6, gate148inter7, gate148inter8, gate148inter9, gate148inter10, gate148inter11, gate148inter12, gate193inter0, gate193inter1, gate193inter2, gate193inter3, gate193inter4, gate193inter5, gate193inter6, gate193inter7, gate193inter8, gate193inter9, gate193inter10, gate193inter11, gate193inter12, gate15inter0, gate15inter1, gate15inter2, gate15inter3, gate15inter4, gate15inter5, gate15inter6, gate15inter7, gate15inter8, gate15inter9, gate15inter10, gate15inter11, gate15inter12, gate216inter0, gate216inter1, gate216inter2, gate216inter3, gate216inter4, gate216inter5, gate216inter6, gate216inter7, gate216inter8, gate216inter9, gate216inter10, gate216inter11, gate216inter12, gate276inter0, gate276inter1, gate276inter2, gate276inter3, gate276inter4, gate276inter5, gate276inter6, gate276inter7, gate276inter8, gate276inter9, gate276inter10, gate276inter11, gate276inter12, gate153inter0, gate153inter1, gate153inter2, gate153inter3, gate153inter4, gate153inter5, gate153inter6, gate153inter7, gate153inter8, gate153inter9, gate153inter10, gate153inter11, gate153inter12, gate192inter0, gate192inter1, gate192inter2, gate192inter3, gate192inter4, gate192inter5, gate192inter6, gate192inter7, gate192inter8, gate192inter9, gate192inter10, gate192inter11, gate192inter12, gate170inter0, gate170inter1, gate170inter2, gate170inter3, gate170inter4, gate170inter5, gate170inter6, gate170inter7, gate170inter8, gate170inter9, gate170inter10, gate170inter11, gate170inter12, gate160inter0, gate160inter1, gate160inter2, gate160inter3, gate160inter4, gate160inter5, gate160inter6, gate160inter7, gate160inter8, gate160inter9, gate160inter10, gate160inter11, gate160inter12, gate214inter0, gate214inter1, gate214inter2, gate214inter3, gate214inter4, gate214inter5, gate214inter6, gate214inter7, gate214inter8, gate214inter9, gate214inter10, gate214inter11, gate214inter12, gate471inter0, gate471inter1, gate471inter2, gate471inter3, gate471inter4, gate471inter5, gate471inter6, gate471inter7, gate471inter8, gate471inter9, gate471inter10, gate471inter11, gate471inter12, gate122inter0, gate122inter1, gate122inter2, gate122inter3, gate122inter4, gate122inter5, gate122inter6, gate122inter7, gate122inter8, gate122inter9, gate122inter10, gate122inter11, gate122inter12, gate428inter0, gate428inter1, gate428inter2, gate428inter3, gate428inter4, gate428inter5, gate428inter6, gate428inter7, gate428inter8, gate428inter9, gate428inter10, gate428inter11, gate428inter12, gate212inter0, gate212inter1, gate212inter2, gate212inter3, gate212inter4, gate212inter5, gate212inter6, gate212inter7, gate212inter8, gate212inter9, gate212inter10, gate212inter11, gate212inter12, gate436inter0, gate436inter1, gate436inter2, gate436inter3, gate436inter4, gate436inter5, gate436inter6, gate436inter7, gate436inter8, gate436inter9, gate436inter10, gate436inter11, gate436inter12, gate467inter0, gate467inter1, gate467inter2, gate467inter3, gate467inter4, gate467inter5, gate467inter6, gate467inter7, gate467inter8, gate467inter9, gate467inter10, gate467inter11, gate467inter12, gate11inter0, gate11inter1, gate11inter2, gate11inter3, gate11inter4, gate11inter5, gate11inter6, gate11inter7, gate11inter8, gate11inter9, gate11inter10, gate11inter11, gate11inter12, gate81inter0, gate81inter1, gate81inter2, gate81inter3, gate81inter4, gate81inter5, gate81inter6, gate81inter7, gate81inter8, gate81inter9, gate81inter10, gate81inter11, gate81inter12, gate247inter0, gate247inter1, gate247inter2, gate247inter3, gate247inter4, gate247inter5, gate247inter6, gate247inter7, gate247inter8, gate247inter9, gate247inter10, gate247inter11, gate247inter12, gate387inter0, gate387inter1, gate387inter2, gate387inter3, gate387inter4, gate387inter5, gate387inter6, gate387inter7, gate387inter8, gate387inter9, gate387inter10, gate387inter11, gate387inter12, gate432inter0, gate432inter1, gate432inter2, gate432inter3, gate432inter4, gate432inter5, gate432inter6, gate432inter7, gate432inter8, gate432inter9, gate432inter10, gate432inter11, gate432inter12, gate45inter0, gate45inter1, gate45inter2, gate45inter3, gate45inter4, gate45inter5, gate45inter6, gate45inter7, gate45inter8, gate45inter9, gate45inter10, gate45inter11, gate45inter12, gate269inter0, gate269inter1, gate269inter2, gate269inter3, gate269inter4, gate269inter5, gate269inter6, gate269inter7, gate269inter8, gate269inter9, gate269inter10, gate269inter11, gate269inter12, gate272inter0, gate272inter1, gate272inter2, gate272inter3, gate272inter4, gate272inter5, gate272inter6, gate272inter7, gate272inter8, gate272inter9, gate272inter10, gate272inter11, gate272inter12, gate415inter0, gate415inter1, gate415inter2, gate415inter3, gate415inter4, gate415inter5, gate415inter6, gate415inter7, gate415inter8, gate415inter9, gate415inter10, gate415inter11, gate415inter12, gate90inter0, gate90inter1, gate90inter2, gate90inter3, gate90inter4, gate90inter5, gate90inter6, gate90inter7, gate90inter8, gate90inter9, gate90inter10, gate90inter11, gate90inter12, gate491inter0, gate491inter1, gate491inter2, gate491inter3, gate491inter4, gate491inter5, gate491inter6, gate491inter7, gate491inter8, gate491inter9, gate491inter10, gate491inter11, gate491inter12, gate164inter0, gate164inter1, gate164inter2, gate164inter3, gate164inter4, gate164inter5, gate164inter6, gate164inter7, gate164inter8, gate164inter9, gate164inter10, gate164inter11, gate164inter12, gate433inter0, gate433inter1, gate433inter2, gate433inter3, gate433inter4, gate433inter5, gate433inter6, gate433inter7, gate433inter8, gate433inter9, gate433inter10, gate433inter11, gate433inter12, gate435inter0, gate435inter1, gate435inter2, gate435inter3, gate435inter4, gate435inter5, gate435inter6, gate435inter7, gate435inter8, gate435inter9, gate435inter10, gate435inter11, gate435inter12, gate31inter0, gate31inter1, gate31inter2, gate31inter3, gate31inter4, gate31inter5, gate31inter6, gate31inter7, gate31inter8, gate31inter9, gate31inter10, gate31inter11, gate31inter12, gate217inter0, gate217inter1, gate217inter2, gate217inter3, gate217inter4, gate217inter5, gate217inter6, gate217inter7, gate217inter8, gate217inter9, gate217inter10, gate217inter11, gate217inter12, gate190inter0, gate190inter1, gate190inter2, gate190inter3, gate190inter4, gate190inter5, gate190inter6, gate190inter7, gate190inter8, gate190inter9, gate190inter10, gate190inter11, gate190inter12, gate444inter0, gate444inter1, gate444inter2, gate444inter3, gate444inter4, gate444inter5, gate444inter6, gate444inter7, gate444inter8, gate444inter9, gate444inter10, gate444inter11, gate444inter12, gate264inter0, gate264inter1, gate264inter2, gate264inter3, gate264inter4, gate264inter5, gate264inter6, gate264inter7, gate264inter8, gate264inter9, gate264inter10, gate264inter11, gate264inter12, gate75inter0, gate75inter1, gate75inter2, gate75inter3, gate75inter4, gate75inter5, gate75inter6, gate75inter7, gate75inter8, gate75inter9, gate75inter10, gate75inter11, gate75inter12, gate14inter0, gate14inter1, gate14inter2, gate14inter3, gate14inter4, gate14inter5, gate14inter6, gate14inter7, gate14inter8, gate14inter9, gate14inter10, gate14inter11, gate14inter12, gate97inter0, gate97inter1, gate97inter2, gate97inter3, gate97inter4, gate97inter5, gate97inter6, gate97inter7, gate97inter8, gate97inter9, gate97inter10, gate97inter11, gate97inter12, gate104inter0, gate104inter1, gate104inter2, gate104inter3, gate104inter4, gate104inter5, gate104inter6, gate104inter7, gate104inter8, gate104inter9, gate104inter10, gate104inter11, gate104inter12, gate218inter0, gate218inter1, gate218inter2, gate218inter3, gate218inter4, gate218inter5, gate218inter6, gate218inter7, gate218inter8, gate218inter9, gate218inter10, gate218inter11, gate218inter12, gate416inter0, gate416inter1, gate416inter2, gate416inter3, gate416inter4, gate416inter5, gate416inter6, gate416inter7, gate416inter8, gate416inter9, gate416inter10, gate416inter11, gate416inter12, gate497inter0, gate497inter1, gate497inter2, gate497inter3, gate497inter4, gate497inter5, gate497inter6, gate497inter7, gate497inter8, gate497inter9, gate497inter10, gate497inter11, gate497inter12, gate191inter0, gate191inter1, gate191inter2, gate191inter3, gate191inter4, gate191inter5, gate191inter6, gate191inter7, gate191inter8, gate191inter9, gate191inter10, gate191inter11, gate191inter12, gate201inter0, gate201inter1, gate201inter2, gate201inter3, gate201inter4, gate201inter5, gate201inter6, gate201inter7, gate201inter8, gate201inter9, gate201inter10, gate201inter11, gate201inter12, gate211inter0, gate211inter1, gate211inter2, gate211inter3, gate211inter4, gate211inter5, gate211inter6, gate211inter7, gate211inter8, gate211inter9, gate211inter10, gate211inter11, gate211inter12, gate95inter0, gate95inter1, gate95inter2, gate95inter3, gate95inter4, gate95inter5, gate95inter6, gate95inter7, gate95inter8, gate95inter9, gate95inter10, gate95inter11, gate95inter12, gate96inter0, gate96inter1, gate96inter2, gate96inter3, gate96inter4, gate96inter5, gate96inter6, gate96inter7, gate96inter8, gate96inter9, gate96inter10, gate96inter11, gate96inter12, gate226inter0, gate226inter1, gate226inter2, gate226inter3, gate226inter4, gate226inter5, gate226inter6, gate226inter7, gate226inter8, gate226inter9, gate226inter10, gate226inter11, gate226inter12, gate388inter0, gate388inter1, gate388inter2, gate388inter3, gate388inter4, gate388inter5, gate388inter6, gate388inter7, gate388inter8, gate388inter9, gate388inter10, gate388inter11, gate388inter12, gate271inter0, gate271inter1, gate271inter2, gate271inter3, gate271inter4, gate271inter5, gate271inter6, gate271inter7, gate271inter8, gate271inter9, gate271inter10, gate271inter11, gate271inter12, gate157inter0, gate157inter1, gate157inter2, gate157inter3, gate157inter4, gate157inter5, gate157inter6, gate157inter7, gate157inter8, gate157inter9, gate157inter10, gate157inter11, gate157inter12, gate468inter0, gate468inter1, gate468inter2, gate468inter3, gate468inter4, gate468inter5, gate468inter6, gate468inter7, gate468inter8, gate468inter9, gate468inter10, gate468inter11, gate468inter12, gate125inter0, gate125inter1, gate125inter2, gate125inter3, gate125inter4, gate125inter5, gate125inter6, gate125inter7, gate125inter8, gate125inter9, gate125inter10, gate125inter11, gate125inter12, gate184inter0, gate184inter1, gate184inter2, gate184inter3, gate184inter4, gate184inter5, gate184inter6, gate184inter7, gate184inter8, gate184inter9, gate184inter10, gate184inter11, gate184inter12, gate228inter0, gate228inter1, gate228inter2, gate228inter3, gate228inter4, gate228inter5, gate228inter6, gate228inter7, gate228inter8, gate228inter9, gate228inter10, gate228inter11, gate228inter12, gate277inter0, gate277inter1, gate277inter2, gate277inter3, gate277inter4, gate277inter5, gate277inter6, gate277inter7, gate277inter8, gate277inter9, gate277inter10, gate277inter11, gate277inter12, gate20inter0, gate20inter1, gate20inter2, gate20inter3, gate20inter4, gate20inter5, gate20inter6, gate20inter7, gate20inter8, gate20inter9, gate20inter10, gate20inter11, gate20inter12, gate250inter0, gate250inter1, gate250inter2, gate250inter3, gate250inter4, gate250inter5, gate250inter6, gate250inter7, gate250inter8, gate250inter9, gate250inter10, gate250inter11, gate250inter12, gate254inter0, gate254inter1, gate254inter2, gate254inter3, gate254inter4, gate254inter5, gate254inter6, gate254inter7, gate254inter8, gate254inter9, gate254inter10, gate254inter11, gate254inter12, gate38inter0, gate38inter1, gate38inter2, gate38inter3, gate38inter4, gate38inter5, gate38inter6, gate38inter7, gate38inter8, gate38inter9, gate38inter10, gate38inter11, gate38inter12, gate46inter0, gate46inter1, gate46inter2, gate46inter3, gate46inter4, gate46inter5, gate46inter6, gate46inter7, gate46inter8, gate46inter9, gate46inter10, gate46inter11, gate46inter12, gate73inter0, gate73inter1, gate73inter2, gate73inter3, gate73inter4, gate73inter5, gate73inter6, gate73inter7, gate73inter8, gate73inter9, gate73inter10, gate73inter11, gate73inter12, gate10inter0, gate10inter1, gate10inter2, gate10inter3, gate10inter4, gate10inter5, gate10inter6, gate10inter7, gate10inter8, gate10inter9, gate10inter10, gate10inter11, gate10inter12, gate427inter0, gate427inter1, gate427inter2, gate427inter3, gate427inter4, gate427inter5, gate427inter6, gate427inter7, gate427inter8, gate427inter9, gate427inter10, gate427inter11, gate427inter12, gate431inter0, gate431inter1, gate431inter2, gate431inter3, gate431inter4, gate431inter5, gate431inter6, gate431inter7, gate431inter8, gate431inter9, gate431inter10, gate431inter11, gate431inter12, gate107inter0, gate107inter1, gate107inter2, gate107inter3, gate107inter4, gate107inter5, gate107inter6, gate107inter7, gate107inter8, gate107inter9, gate107inter10, gate107inter11, gate107inter12, gate140inter0, gate140inter1, gate140inter2, gate140inter3, gate140inter4, gate140inter5, gate140inter6, gate140inter7, gate140inter8, gate140inter9, gate140inter10, gate140inter11, gate140inter12, gate482inter0, gate482inter1, gate482inter2, gate482inter3, gate482inter4, gate482inter5, gate482inter6, gate482inter7, gate482inter8, gate482inter9, gate482inter10, gate482inter11, gate482inter12, gate93inter0, gate93inter1, gate93inter2, gate93inter3, gate93inter4, gate93inter5, gate93inter6, gate93inter7, gate93inter8, gate93inter9, gate93inter10, gate93inter11, gate93inter12, gate83inter0, gate83inter1, gate83inter2, gate83inter3, gate83inter4, gate83inter5, gate83inter6, gate83inter7, gate83inter8, gate83inter9, gate83inter10, gate83inter11, gate83inter12, gate279inter0, gate279inter1, gate279inter2, gate279inter3, gate279inter4, gate279inter5, gate279inter6, gate279inter7, gate279inter8, gate279inter9, gate279inter10, gate279inter11, gate279inter12, gate403inter0, gate403inter1, gate403inter2, gate403inter3, gate403inter4, gate403inter5, gate403inter6, gate403inter7, gate403inter8, gate403inter9, gate403inter10, gate403inter11, gate403inter12;



and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );
nand2 gate9( .a(G1), .b(G2), .O(G266) );

  xor2  gate1471(.a(G4), .b(G3), .O(gate10inter0));
  nand2 gate1472(.a(gate10inter0), .b(s_132), .O(gate10inter1));
  and2  gate1473(.a(G4), .b(G3), .O(gate10inter2));
  inv1  gate1474(.a(s_132), .O(gate10inter3));
  inv1  gate1475(.a(s_133), .O(gate10inter4));
  nand2 gate1476(.a(gate10inter4), .b(gate10inter3), .O(gate10inter5));
  nor2  gate1477(.a(gate10inter5), .b(gate10inter2), .O(gate10inter6));
  inv1  gate1478(.a(G3), .O(gate10inter7));
  inv1  gate1479(.a(G4), .O(gate10inter8));
  nand2 gate1480(.a(gate10inter8), .b(gate10inter7), .O(gate10inter9));
  nand2 gate1481(.a(s_133), .b(gate10inter3), .O(gate10inter10));
  nor2  gate1482(.a(gate10inter10), .b(gate10inter9), .O(gate10inter11));
  nor2  gate1483(.a(gate10inter11), .b(gate10inter6), .O(gate10inter12));
  nand2 gate1484(.a(gate10inter12), .b(gate10inter1), .O(G269));

  xor2  gate827(.a(G6), .b(G5), .O(gate11inter0));
  nand2 gate828(.a(gate11inter0), .b(s_40), .O(gate11inter1));
  and2  gate829(.a(G6), .b(G5), .O(gate11inter2));
  inv1  gate830(.a(s_40), .O(gate11inter3));
  inv1  gate831(.a(s_41), .O(gate11inter4));
  nand2 gate832(.a(gate11inter4), .b(gate11inter3), .O(gate11inter5));
  nor2  gate833(.a(gate11inter5), .b(gate11inter2), .O(gate11inter6));
  inv1  gate834(.a(G5), .O(gate11inter7));
  inv1  gate835(.a(G6), .O(gate11inter8));
  nand2 gate836(.a(gate11inter8), .b(gate11inter7), .O(gate11inter9));
  nand2 gate837(.a(s_41), .b(gate11inter3), .O(gate11inter10));
  nor2  gate838(.a(gate11inter10), .b(gate11inter9), .O(gate11inter11));
  nor2  gate839(.a(gate11inter11), .b(gate11inter6), .O(gate11inter12));
  nand2 gate840(.a(gate11inter12), .b(gate11inter1), .O(G272));
nand2 gate12( .a(G7), .b(G8), .O(G275) );
nand2 gate13( .a(G9), .b(G10), .O(G278) );

  xor2  gate1107(.a(G12), .b(G11), .O(gate14inter0));
  nand2 gate1108(.a(gate14inter0), .b(s_80), .O(gate14inter1));
  and2  gate1109(.a(G12), .b(G11), .O(gate14inter2));
  inv1  gate1110(.a(s_80), .O(gate14inter3));
  inv1  gate1111(.a(s_81), .O(gate14inter4));
  nand2 gate1112(.a(gate14inter4), .b(gate14inter3), .O(gate14inter5));
  nor2  gate1113(.a(gate14inter5), .b(gate14inter2), .O(gate14inter6));
  inv1  gate1114(.a(G11), .O(gate14inter7));
  inv1  gate1115(.a(G12), .O(gate14inter8));
  nand2 gate1116(.a(gate14inter8), .b(gate14inter7), .O(gate14inter9));
  nand2 gate1117(.a(s_81), .b(gate14inter3), .O(gate14inter10));
  nor2  gate1118(.a(gate14inter10), .b(gate14inter9), .O(gate14inter11));
  nor2  gate1119(.a(gate14inter11), .b(gate14inter6), .O(gate14inter12));
  nand2 gate1120(.a(gate14inter12), .b(gate14inter1), .O(G281));

  xor2  gate631(.a(G14), .b(G13), .O(gate15inter0));
  nand2 gate632(.a(gate15inter0), .b(s_12), .O(gate15inter1));
  and2  gate633(.a(G14), .b(G13), .O(gate15inter2));
  inv1  gate634(.a(s_12), .O(gate15inter3));
  inv1  gate635(.a(s_13), .O(gate15inter4));
  nand2 gate636(.a(gate15inter4), .b(gate15inter3), .O(gate15inter5));
  nor2  gate637(.a(gate15inter5), .b(gate15inter2), .O(gate15inter6));
  inv1  gate638(.a(G13), .O(gate15inter7));
  inv1  gate639(.a(G14), .O(gate15inter8));
  nand2 gate640(.a(gate15inter8), .b(gate15inter7), .O(gate15inter9));
  nand2 gate641(.a(s_13), .b(gate15inter3), .O(gate15inter10));
  nor2  gate642(.a(gate15inter10), .b(gate15inter9), .O(gate15inter11));
  nor2  gate643(.a(gate15inter11), .b(gate15inter6), .O(gate15inter12));
  nand2 gate644(.a(gate15inter12), .b(gate15inter1), .O(G284));
nand2 gate16( .a(G15), .b(G16), .O(G287) );
nand2 gate17( .a(G17), .b(G18), .O(G290) );
nand2 gate18( .a(G19), .b(G20), .O(G293) );
nand2 gate19( .a(G21), .b(G22), .O(G296) );

  xor2  gate1387(.a(G24), .b(G23), .O(gate20inter0));
  nand2 gate1388(.a(gate20inter0), .b(s_120), .O(gate20inter1));
  and2  gate1389(.a(G24), .b(G23), .O(gate20inter2));
  inv1  gate1390(.a(s_120), .O(gate20inter3));
  inv1  gate1391(.a(s_121), .O(gate20inter4));
  nand2 gate1392(.a(gate20inter4), .b(gate20inter3), .O(gate20inter5));
  nor2  gate1393(.a(gate20inter5), .b(gate20inter2), .O(gate20inter6));
  inv1  gate1394(.a(G23), .O(gate20inter7));
  inv1  gate1395(.a(G24), .O(gate20inter8));
  nand2 gate1396(.a(gate20inter8), .b(gate20inter7), .O(gate20inter9));
  nand2 gate1397(.a(s_121), .b(gate20inter3), .O(gate20inter10));
  nor2  gate1398(.a(gate20inter10), .b(gate20inter9), .O(gate20inter11));
  nor2  gate1399(.a(gate20inter11), .b(gate20inter6), .O(gate20inter12));
  nand2 gate1400(.a(gate20inter12), .b(gate20inter1), .O(G299));
nand2 gate21( .a(G25), .b(G26), .O(G302) );
nand2 gate22( .a(G27), .b(G28), .O(G305) );
nand2 gate23( .a(G29), .b(G30), .O(G308) );
nand2 gate24( .a(G31), .b(G32), .O(G311) );
nand2 gate25( .a(G1), .b(G5), .O(G314) );
nand2 gate26( .a(G9), .b(G13), .O(G317) );
nand2 gate27( .a(G2), .b(G6), .O(G320) );
nand2 gate28( .a(G10), .b(G14), .O(G323) );
nand2 gate29( .a(G3), .b(G7), .O(G326) );
nand2 gate30( .a(G11), .b(G15), .O(G329) );

  xor2  gate1023(.a(G8), .b(G4), .O(gate31inter0));
  nand2 gate1024(.a(gate31inter0), .b(s_68), .O(gate31inter1));
  and2  gate1025(.a(G8), .b(G4), .O(gate31inter2));
  inv1  gate1026(.a(s_68), .O(gate31inter3));
  inv1  gate1027(.a(s_69), .O(gate31inter4));
  nand2 gate1028(.a(gate31inter4), .b(gate31inter3), .O(gate31inter5));
  nor2  gate1029(.a(gate31inter5), .b(gate31inter2), .O(gate31inter6));
  inv1  gate1030(.a(G4), .O(gate31inter7));
  inv1  gate1031(.a(G8), .O(gate31inter8));
  nand2 gate1032(.a(gate31inter8), .b(gate31inter7), .O(gate31inter9));
  nand2 gate1033(.a(s_69), .b(gate31inter3), .O(gate31inter10));
  nor2  gate1034(.a(gate31inter10), .b(gate31inter9), .O(gate31inter11));
  nor2  gate1035(.a(gate31inter11), .b(gate31inter6), .O(gate31inter12));
  nand2 gate1036(.a(gate31inter12), .b(gate31inter1), .O(G332));
nand2 gate32( .a(G12), .b(G16), .O(G335) );
nand2 gate33( .a(G17), .b(G21), .O(G338) );
nand2 gate34( .a(G25), .b(G29), .O(G341) );
nand2 gate35( .a(G18), .b(G22), .O(G344) );
nand2 gate36( .a(G26), .b(G30), .O(G347) );
nand2 gate37( .a(G19), .b(G23), .O(G350) );

  xor2  gate1429(.a(G31), .b(G27), .O(gate38inter0));
  nand2 gate1430(.a(gate38inter0), .b(s_126), .O(gate38inter1));
  and2  gate1431(.a(G31), .b(G27), .O(gate38inter2));
  inv1  gate1432(.a(s_126), .O(gate38inter3));
  inv1  gate1433(.a(s_127), .O(gate38inter4));
  nand2 gate1434(.a(gate38inter4), .b(gate38inter3), .O(gate38inter5));
  nor2  gate1435(.a(gate38inter5), .b(gate38inter2), .O(gate38inter6));
  inv1  gate1436(.a(G27), .O(gate38inter7));
  inv1  gate1437(.a(G31), .O(gate38inter8));
  nand2 gate1438(.a(gate38inter8), .b(gate38inter7), .O(gate38inter9));
  nand2 gate1439(.a(s_127), .b(gate38inter3), .O(gate38inter10));
  nor2  gate1440(.a(gate38inter10), .b(gate38inter9), .O(gate38inter11));
  nor2  gate1441(.a(gate38inter11), .b(gate38inter6), .O(gate38inter12));
  nand2 gate1442(.a(gate38inter12), .b(gate38inter1), .O(G353));
nand2 gate39( .a(G20), .b(G24), .O(G356) );
nand2 gate40( .a(G28), .b(G32), .O(G359) );
nand2 gate41( .a(G1), .b(G266), .O(G362) );
nand2 gate42( .a(G2), .b(G266), .O(G363) );
nand2 gate43( .a(G3), .b(G269), .O(G364) );
nand2 gate44( .a(G4), .b(G269), .O(G365) );

  xor2  gate897(.a(G272), .b(G5), .O(gate45inter0));
  nand2 gate898(.a(gate45inter0), .b(s_50), .O(gate45inter1));
  and2  gate899(.a(G272), .b(G5), .O(gate45inter2));
  inv1  gate900(.a(s_50), .O(gate45inter3));
  inv1  gate901(.a(s_51), .O(gate45inter4));
  nand2 gate902(.a(gate45inter4), .b(gate45inter3), .O(gate45inter5));
  nor2  gate903(.a(gate45inter5), .b(gate45inter2), .O(gate45inter6));
  inv1  gate904(.a(G5), .O(gate45inter7));
  inv1  gate905(.a(G272), .O(gate45inter8));
  nand2 gate906(.a(gate45inter8), .b(gate45inter7), .O(gate45inter9));
  nand2 gate907(.a(s_51), .b(gate45inter3), .O(gate45inter10));
  nor2  gate908(.a(gate45inter10), .b(gate45inter9), .O(gate45inter11));
  nor2  gate909(.a(gate45inter11), .b(gate45inter6), .O(gate45inter12));
  nand2 gate910(.a(gate45inter12), .b(gate45inter1), .O(G366));

  xor2  gate1443(.a(G272), .b(G6), .O(gate46inter0));
  nand2 gate1444(.a(gate46inter0), .b(s_128), .O(gate46inter1));
  and2  gate1445(.a(G272), .b(G6), .O(gate46inter2));
  inv1  gate1446(.a(s_128), .O(gate46inter3));
  inv1  gate1447(.a(s_129), .O(gate46inter4));
  nand2 gate1448(.a(gate46inter4), .b(gate46inter3), .O(gate46inter5));
  nor2  gate1449(.a(gate46inter5), .b(gate46inter2), .O(gate46inter6));
  inv1  gate1450(.a(G6), .O(gate46inter7));
  inv1  gate1451(.a(G272), .O(gate46inter8));
  nand2 gate1452(.a(gate46inter8), .b(gate46inter7), .O(gate46inter9));
  nand2 gate1453(.a(s_129), .b(gate46inter3), .O(gate46inter10));
  nor2  gate1454(.a(gate46inter10), .b(gate46inter9), .O(gate46inter11));
  nor2  gate1455(.a(gate46inter11), .b(gate46inter6), .O(gate46inter12));
  nand2 gate1456(.a(gate46inter12), .b(gate46inter1), .O(G367));
nand2 gate47( .a(G7), .b(G275), .O(G368) );
nand2 gate48( .a(G8), .b(G275), .O(G369) );
nand2 gate49( .a(G9), .b(G278), .O(G370) );
nand2 gate50( .a(G10), .b(G278), .O(G371) );
nand2 gate51( .a(G11), .b(G281), .O(G372) );
nand2 gate52( .a(G12), .b(G281), .O(G373) );
nand2 gate53( .a(G13), .b(G284), .O(G374) );
nand2 gate54( .a(G14), .b(G284), .O(G375) );
nand2 gate55( .a(G15), .b(G287), .O(G376) );
nand2 gate56( .a(G16), .b(G287), .O(G377) );
nand2 gate57( .a(G17), .b(G290), .O(G378) );
nand2 gate58( .a(G18), .b(G290), .O(G379) );
nand2 gate59( .a(G19), .b(G293), .O(G380) );
nand2 gate60( .a(G20), .b(G293), .O(G381) );
nand2 gate61( .a(G21), .b(G296), .O(G382) );
nand2 gate62( .a(G22), .b(G296), .O(G383) );
nand2 gate63( .a(G23), .b(G299), .O(G384) );
nand2 gate64( .a(G24), .b(G299), .O(G385) );
nand2 gate65( .a(G25), .b(G302), .O(G386) );
nand2 gate66( .a(G26), .b(G302), .O(G387) );
nand2 gate67( .a(G27), .b(G305), .O(G388) );
nand2 gate68( .a(G28), .b(G305), .O(G389) );
nand2 gate69( .a(G29), .b(G308), .O(G390) );
nand2 gate70( .a(G30), .b(G308), .O(G391) );
nand2 gate71( .a(G31), .b(G311), .O(G392) );
nand2 gate72( .a(G32), .b(G311), .O(G393) );

  xor2  gate1457(.a(G314), .b(G1), .O(gate73inter0));
  nand2 gate1458(.a(gate73inter0), .b(s_130), .O(gate73inter1));
  and2  gate1459(.a(G314), .b(G1), .O(gate73inter2));
  inv1  gate1460(.a(s_130), .O(gate73inter3));
  inv1  gate1461(.a(s_131), .O(gate73inter4));
  nand2 gate1462(.a(gate73inter4), .b(gate73inter3), .O(gate73inter5));
  nor2  gate1463(.a(gate73inter5), .b(gate73inter2), .O(gate73inter6));
  inv1  gate1464(.a(G1), .O(gate73inter7));
  inv1  gate1465(.a(G314), .O(gate73inter8));
  nand2 gate1466(.a(gate73inter8), .b(gate73inter7), .O(gate73inter9));
  nand2 gate1467(.a(s_131), .b(gate73inter3), .O(gate73inter10));
  nor2  gate1468(.a(gate73inter10), .b(gate73inter9), .O(gate73inter11));
  nor2  gate1469(.a(gate73inter11), .b(gate73inter6), .O(gate73inter12));
  nand2 gate1470(.a(gate73inter12), .b(gate73inter1), .O(G394));
nand2 gate74( .a(G5), .b(G314), .O(G395) );

  xor2  gate1093(.a(G317), .b(G9), .O(gate75inter0));
  nand2 gate1094(.a(gate75inter0), .b(s_78), .O(gate75inter1));
  and2  gate1095(.a(G317), .b(G9), .O(gate75inter2));
  inv1  gate1096(.a(s_78), .O(gate75inter3));
  inv1  gate1097(.a(s_79), .O(gate75inter4));
  nand2 gate1098(.a(gate75inter4), .b(gate75inter3), .O(gate75inter5));
  nor2  gate1099(.a(gate75inter5), .b(gate75inter2), .O(gate75inter6));
  inv1  gate1100(.a(G9), .O(gate75inter7));
  inv1  gate1101(.a(G317), .O(gate75inter8));
  nand2 gate1102(.a(gate75inter8), .b(gate75inter7), .O(gate75inter9));
  nand2 gate1103(.a(s_79), .b(gate75inter3), .O(gate75inter10));
  nor2  gate1104(.a(gate75inter10), .b(gate75inter9), .O(gate75inter11));
  nor2  gate1105(.a(gate75inter11), .b(gate75inter6), .O(gate75inter12));
  nand2 gate1106(.a(gate75inter12), .b(gate75inter1), .O(G396));
nand2 gate76( .a(G13), .b(G317), .O(G397) );
nand2 gate77( .a(G2), .b(G320), .O(G398) );
nand2 gate78( .a(G6), .b(G320), .O(G399) );
nand2 gate79( .a(G10), .b(G323), .O(G400) );
nand2 gate80( .a(G14), .b(G323), .O(G401) );

  xor2  gate841(.a(G326), .b(G3), .O(gate81inter0));
  nand2 gate842(.a(gate81inter0), .b(s_42), .O(gate81inter1));
  and2  gate843(.a(G326), .b(G3), .O(gate81inter2));
  inv1  gate844(.a(s_42), .O(gate81inter3));
  inv1  gate845(.a(s_43), .O(gate81inter4));
  nand2 gate846(.a(gate81inter4), .b(gate81inter3), .O(gate81inter5));
  nor2  gate847(.a(gate81inter5), .b(gate81inter2), .O(gate81inter6));
  inv1  gate848(.a(G3), .O(gate81inter7));
  inv1  gate849(.a(G326), .O(gate81inter8));
  nand2 gate850(.a(gate81inter8), .b(gate81inter7), .O(gate81inter9));
  nand2 gate851(.a(s_43), .b(gate81inter3), .O(gate81inter10));
  nor2  gate852(.a(gate81inter10), .b(gate81inter9), .O(gate81inter11));
  nor2  gate853(.a(gate81inter11), .b(gate81inter6), .O(gate81inter12));
  nand2 gate854(.a(gate81inter12), .b(gate81inter1), .O(G402));
nand2 gate82( .a(G7), .b(G326), .O(G403) );

  xor2  gate1569(.a(G329), .b(G11), .O(gate83inter0));
  nand2 gate1570(.a(gate83inter0), .b(s_146), .O(gate83inter1));
  and2  gate1571(.a(G329), .b(G11), .O(gate83inter2));
  inv1  gate1572(.a(s_146), .O(gate83inter3));
  inv1  gate1573(.a(s_147), .O(gate83inter4));
  nand2 gate1574(.a(gate83inter4), .b(gate83inter3), .O(gate83inter5));
  nor2  gate1575(.a(gate83inter5), .b(gate83inter2), .O(gate83inter6));
  inv1  gate1576(.a(G11), .O(gate83inter7));
  inv1  gate1577(.a(G329), .O(gate83inter8));
  nand2 gate1578(.a(gate83inter8), .b(gate83inter7), .O(gate83inter9));
  nand2 gate1579(.a(s_147), .b(gate83inter3), .O(gate83inter10));
  nor2  gate1580(.a(gate83inter10), .b(gate83inter9), .O(gate83inter11));
  nor2  gate1581(.a(gate83inter11), .b(gate83inter6), .O(gate83inter12));
  nand2 gate1582(.a(gate83inter12), .b(gate83inter1), .O(G404));
nand2 gate84( .a(G15), .b(G329), .O(G405) );
nand2 gate85( .a(G4), .b(G332), .O(G406) );
nand2 gate86( .a(G8), .b(G332), .O(G407) );
nand2 gate87( .a(G12), .b(G335), .O(G408) );
nand2 gate88( .a(G16), .b(G335), .O(G409) );
nand2 gate89( .a(G17), .b(G338), .O(G410) );

  xor2  gate953(.a(G338), .b(G21), .O(gate90inter0));
  nand2 gate954(.a(gate90inter0), .b(s_58), .O(gate90inter1));
  and2  gate955(.a(G338), .b(G21), .O(gate90inter2));
  inv1  gate956(.a(s_58), .O(gate90inter3));
  inv1  gate957(.a(s_59), .O(gate90inter4));
  nand2 gate958(.a(gate90inter4), .b(gate90inter3), .O(gate90inter5));
  nor2  gate959(.a(gate90inter5), .b(gate90inter2), .O(gate90inter6));
  inv1  gate960(.a(G21), .O(gate90inter7));
  inv1  gate961(.a(G338), .O(gate90inter8));
  nand2 gate962(.a(gate90inter8), .b(gate90inter7), .O(gate90inter9));
  nand2 gate963(.a(s_59), .b(gate90inter3), .O(gate90inter10));
  nor2  gate964(.a(gate90inter10), .b(gate90inter9), .O(gate90inter11));
  nor2  gate965(.a(gate90inter11), .b(gate90inter6), .O(gate90inter12));
  nand2 gate966(.a(gate90inter12), .b(gate90inter1), .O(G411));
nand2 gate91( .a(G25), .b(G341), .O(G412) );
nand2 gate92( .a(G29), .b(G341), .O(G413) );

  xor2  gate1555(.a(G344), .b(G18), .O(gate93inter0));
  nand2 gate1556(.a(gate93inter0), .b(s_144), .O(gate93inter1));
  and2  gate1557(.a(G344), .b(G18), .O(gate93inter2));
  inv1  gate1558(.a(s_144), .O(gate93inter3));
  inv1  gate1559(.a(s_145), .O(gate93inter4));
  nand2 gate1560(.a(gate93inter4), .b(gate93inter3), .O(gate93inter5));
  nor2  gate1561(.a(gate93inter5), .b(gate93inter2), .O(gate93inter6));
  inv1  gate1562(.a(G18), .O(gate93inter7));
  inv1  gate1563(.a(G344), .O(gate93inter8));
  nand2 gate1564(.a(gate93inter8), .b(gate93inter7), .O(gate93inter9));
  nand2 gate1565(.a(s_145), .b(gate93inter3), .O(gate93inter10));
  nor2  gate1566(.a(gate93inter10), .b(gate93inter9), .O(gate93inter11));
  nor2  gate1567(.a(gate93inter11), .b(gate93inter6), .O(gate93inter12));
  nand2 gate1568(.a(gate93inter12), .b(gate93inter1), .O(G414));
nand2 gate94( .a(G22), .b(G344), .O(G415) );

  xor2  gate1233(.a(G347), .b(G26), .O(gate95inter0));
  nand2 gate1234(.a(gate95inter0), .b(s_98), .O(gate95inter1));
  and2  gate1235(.a(G347), .b(G26), .O(gate95inter2));
  inv1  gate1236(.a(s_98), .O(gate95inter3));
  inv1  gate1237(.a(s_99), .O(gate95inter4));
  nand2 gate1238(.a(gate95inter4), .b(gate95inter3), .O(gate95inter5));
  nor2  gate1239(.a(gate95inter5), .b(gate95inter2), .O(gate95inter6));
  inv1  gate1240(.a(G26), .O(gate95inter7));
  inv1  gate1241(.a(G347), .O(gate95inter8));
  nand2 gate1242(.a(gate95inter8), .b(gate95inter7), .O(gate95inter9));
  nand2 gate1243(.a(s_99), .b(gate95inter3), .O(gate95inter10));
  nor2  gate1244(.a(gate95inter10), .b(gate95inter9), .O(gate95inter11));
  nor2  gate1245(.a(gate95inter11), .b(gate95inter6), .O(gate95inter12));
  nand2 gate1246(.a(gate95inter12), .b(gate95inter1), .O(G416));

  xor2  gate1247(.a(G347), .b(G30), .O(gate96inter0));
  nand2 gate1248(.a(gate96inter0), .b(s_100), .O(gate96inter1));
  and2  gate1249(.a(G347), .b(G30), .O(gate96inter2));
  inv1  gate1250(.a(s_100), .O(gate96inter3));
  inv1  gate1251(.a(s_101), .O(gate96inter4));
  nand2 gate1252(.a(gate96inter4), .b(gate96inter3), .O(gate96inter5));
  nor2  gate1253(.a(gate96inter5), .b(gate96inter2), .O(gate96inter6));
  inv1  gate1254(.a(G30), .O(gate96inter7));
  inv1  gate1255(.a(G347), .O(gate96inter8));
  nand2 gate1256(.a(gate96inter8), .b(gate96inter7), .O(gate96inter9));
  nand2 gate1257(.a(s_101), .b(gate96inter3), .O(gate96inter10));
  nor2  gate1258(.a(gate96inter10), .b(gate96inter9), .O(gate96inter11));
  nor2  gate1259(.a(gate96inter11), .b(gate96inter6), .O(gate96inter12));
  nand2 gate1260(.a(gate96inter12), .b(gate96inter1), .O(G417));

  xor2  gate1121(.a(G350), .b(G19), .O(gate97inter0));
  nand2 gate1122(.a(gate97inter0), .b(s_82), .O(gate97inter1));
  and2  gate1123(.a(G350), .b(G19), .O(gate97inter2));
  inv1  gate1124(.a(s_82), .O(gate97inter3));
  inv1  gate1125(.a(s_83), .O(gate97inter4));
  nand2 gate1126(.a(gate97inter4), .b(gate97inter3), .O(gate97inter5));
  nor2  gate1127(.a(gate97inter5), .b(gate97inter2), .O(gate97inter6));
  inv1  gate1128(.a(G19), .O(gate97inter7));
  inv1  gate1129(.a(G350), .O(gate97inter8));
  nand2 gate1130(.a(gate97inter8), .b(gate97inter7), .O(gate97inter9));
  nand2 gate1131(.a(s_83), .b(gate97inter3), .O(gate97inter10));
  nor2  gate1132(.a(gate97inter10), .b(gate97inter9), .O(gate97inter11));
  nor2  gate1133(.a(gate97inter11), .b(gate97inter6), .O(gate97inter12));
  nand2 gate1134(.a(gate97inter12), .b(gate97inter1), .O(G418));
nand2 gate98( .a(G23), .b(G350), .O(G419) );
nand2 gate99( .a(G27), .b(G353), .O(G420) );
nand2 gate100( .a(G31), .b(G353), .O(G421) );
nand2 gate101( .a(G20), .b(G356), .O(G422) );
nand2 gate102( .a(G24), .b(G356), .O(G423) );
nand2 gate103( .a(G28), .b(G359), .O(G424) );

  xor2  gate1135(.a(G359), .b(G32), .O(gate104inter0));
  nand2 gate1136(.a(gate104inter0), .b(s_84), .O(gate104inter1));
  and2  gate1137(.a(G359), .b(G32), .O(gate104inter2));
  inv1  gate1138(.a(s_84), .O(gate104inter3));
  inv1  gate1139(.a(s_85), .O(gate104inter4));
  nand2 gate1140(.a(gate104inter4), .b(gate104inter3), .O(gate104inter5));
  nor2  gate1141(.a(gate104inter5), .b(gate104inter2), .O(gate104inter6));
  inv1  gate1142(.a(G32), .O(gate104inter7));
  inv1  gate1143(.a(G359), .O(gate104inter8));
  nand2 gate1144(.a(gate104inter8), .b(gate104inter7), .O(gate104inter9));
  nand2 gate1145(.a(s_85), .b(gate104inter3), .O(gate104inter10));
  nor2  gate1146(.a(gate104inter10), .b(gate104inter9), .O(gate104inter11));
  nor2  gate1147(.a(gate104inter11), .b(gate104inter6), .O(gate104inter12));
  nand2 gate1148(.a(gate104inter12), .b(gate104inter1), .O(G425));
nand2 gate105( .a(G362), .b(G363), .O(G426) );
nand2 gate106( .a(G364), .b(G365), .O(G429) );

  xor2  gate1513(.a(G367), .b(G366), .O(gate107inter0));
  nand2 gate1514(.a(gate107inter0), .b(s_138), .O(gate107inter1));
  and2  gate1515(.a(G367), .b(G366), .O(gate107inter2));
  inv1  gate1516(.a(s_138), .O(gate107inter3));
  inv1  gate1517(.a(s_139), .O(gate107inter4));
  nand2 gate1518(.a(gate107inter4), .b(gate107inter3), .O(gate107inter5));
  nor2  gate1519(.a(gate107inter5), .b(gate107inter2), .O(gate107inter6));
  inv1  gate1520(.a(G366), .O(gate107inter7));
  inv1  gate1521(.a(G367), .O(gate107inter8));
  nand2 gate1522(.a(gate107inter8), .b(gate107inter7), .O(gate107inter9));
  nand2 gate1523(.a(s_139), .b(gate107inter3), .O(gate107inter10));
  nor2  gate1524(.a(gate107inter10), .b(gate107inter9), .O(gate107inter11));
  nor2  gate1525(.a(gate107inter11), .b(gate107inter6), .O(gate107inter12));
  nand2 gate1526(.a(gate107inter12), .b(gate107inter1), .O(G432));
nand2 gate108( .a(G368), .b(G369), .O(G435) );
nand2 gate109( .a(G370), .b(G371), .O(G438) );
nand2 gate110( .a(G372), .b(G373), .O(G441) );
nand2 gate111( .a(G374), .b(G375), .O(G444) );
nand2 gate112( .a(G376), .b(G377), .O(G447) );
nand2 gate113( .a(G378), .b(G379), .O(G450) );
nand2 gate114( .a(G380), .b(G381), .O(G453) );
nand2 gate115( .a(G382), .b(G383), .O(G456) );
nand2 gate116( .a(G384), .b(G385), .O(G459) );
nand2 gate117( .a(G386), .b(G387), .O(G462) );
nand2 gate118( .a(G388), .b(G389), .O(G465) );
nand2 gate119( .a(G390), .b(G391), .O(G468) );

  xor2  gate561(.a(G393), .b(G392), .O(gate120inter0));
  nand2 gate562(.a(gate120inter0), .b(s_2), .O(gate120inter1));
  and2  gate563(.a(G393), .b(G392), .O(gate120inter2));
  inv1  gate564(.a(s_2), .O(gate120inter3));
  inv1  gate565(.a(s_3), .O(gate120inter4));
  nand2 gate566(.a(gate120inter4), .b(gate120inter3), .O(gate120inter5));
  nor2  gate567(.a(gate120inter5), .b(gate120inter2), .O(gate120inter6));
  inv1  gate568(.a(G392), .O(gate120inter7));
  inv1  gate569(.a(G393), .O(gate120inter8));
  nand2 gate570(.a(gate120inter8), .b(gate120inter7), .O(gate120inter9));
  nand2 gate571(.a(s_3), .b(gate120inter3), .O(gate120inter10));
  nor2  gate572(.a(gate120inter10), .b(gate120inter9), .O(gate120inter11));
  nor2  gate573(.a(gate120inter11), .b(gate120inter6), .O(gate120inter12));
  nand2 gate574(.a(gate120inter12), .b(gate120inter1), .O(G471));
nand2 gate121( .a(G394), .b(G395), .O(G474) );

  xor2  gate757(.a(G397), .b(G396), .O(gate122inter0));
  nand2 gate758(.a(gate122inter0), .b(s_30), .O(gate122inter1));
  and2  gate759(.a(G397), .b(G396), .O(gate122inter2));
  inv1  gate760(.a(s_30), .O(gate122inter3));
  inv1  gate761(.a(s_31), .O(gate122inter4));
  nand2 gate762(.a(gate122inter4), .b(gate122inter3), .O(gate122inter5));
  nor2  gate763(.a(gate122inter5), .b(gate122inter2), .O(gate122inter6));
  inv1  gate764(.a(G396), .O(gate122inter7));
  inv1  gate765(.a(G397), .O(gate122inter8));
  nand2 gate766(.a(gate122inter8), .b(gate122inter7), .O(gate122inter9));
  nand2 gate767(.a(s_31), .b(gate122inter3), .O(gate122inter10));
  nor2  gate768(.a(gate122inter10), .b(gate122inter9), .O(gate122inter11));
  nor2  gate769(.a(gate122inter11), .b(gate122inter6), .O(gate122inter12));
  nand2 gate770(.a(gate122inter12), .b(gate122inter1), .O(G477));
nand2 gate123( .a(G398), .b(G399), .O(G480) );
nand2 gate124( .a(G400), .b(G401), .O(G483) );

  xor2  gate1331(.a(G403), .b(G402), .O(gate125inter0));
  nand2 gate1332(.a(gate125inter0), .b(s_112), .O(gate125inter1));
  and2  gate1333(.a(G403), .b(G402), .O(gate125inter2));
  inv1  gate1334(.a(s_112), .O(gate125inter3));
  inv1  gate1335(.a(s_113), .O(gate125inter4));
  nand2 gate1336(.a(gate125inter4), .b(gate125inter3), .O(gate125inter5));
  nor2  gate1337(.a(gate125inter5), .b(gate125inter2), .O(gate125inter6));
  inv1  gate1338(.a(G402), .O(gate125inter7));
  inv1  gate1339(.a(G403), .O(gate125inter8));
  nand2 gate1340(.a(gate125inter8), .b(gate125inter7), .O(gate125inter9));
  nand2 gate1341(.a(s_113), .b(gate125inter3), .O(gate125inter10));
  nor2  gate1342(.a(gate125inter10), .b(gate125inter9), .O(gate125inter11));
  nor2  gate1343(.a(gate125inter11), .b(gate125inter6), .O(gate125inter12));
  nand2 gate1344(.a(gate125inter12), .b(gate125inter1), .O(G486));
nand2 gate126( .a(G404), .b(G405), .O(G489) );
nand2 gate127( .a(G406), .b(G407), .O(G492) );
nand2 gate128( .a(G408), .b(G409), .O(G495) );
nand2 gate129( .a(G410), .b(G411), .O(G498) );
nand2 gate130( .a(G412), .b(G413), .O(G501) );
nand2 gate131( .a(G414), .b(G415), .O(G504) );
nand2 gate132( .a(G416), .b(G417), .O(G507) );
nand2 gate133( .a(G418), .b(G419), .O(G510) );
nand2 gate134( .a(G420), .b(G421), .O(G513) );
nand2 gate135( .a(G422), .b(G423), .O(G516) );
nand2 gate136( .a(G424), .b(G425), .O(G519) );
nand2 gate137( .a(G426), .b(G429), .O(G522) );
nand2 gate138( .a(G432), .b(G435), .O(G525) );
nand2 gate139( .a(G438), .b(G441), .O(G528) );

  xor2  gate1527(.a(G447), .b(G444), .O(gate140inter0));
  nand2 gate1528(.a(gate140inter0), .b(s_140), .O(gate140inter1));
  and2  gate1529(.a(G447), .b(G444), .O(gate140inter2));
  inv1  gate1530(.a(s_140), .O(gate140inter3));
  inv1  gate1531(.a(s_141), .O(gate140inter4));
  nand2 gate1532(.a(gate140inter4), .b(gate140inter3), .O(gate140inter5));
  nor2  gate1533(.a(gate140inter5), .b(gate140inter2), .O(gate140inter6));
  inv1  gate1534(.a(G444), .O(gate140inter7));
  inv1  gate1535(.a(G447), .O(gate140inter8));
  nand2 gate1536(.a(gate140inter8), .b(gate140inter7), .O(gate140inter9));
  nand2 gate1537(.a(s_141), .b(gate140inter3), .O(gate140inter10));
  nor2  gate1538(.a(gate140inter10), .b(gate140inter9), .O(gate140inter11));
  nor2  gate1539(.a(gate140inter11), .b(gate140inter6), .O(gate140inter12));
  nand2 gate1540(.a(gate140inter12), .b(gate140inter1), .O(G531));
nand2 gate141( .a(G450), .b(G453), .O(G534) );
nand2 gate142( .a(G456), .b(G459), .O(G537) );
nand2 gate143( .a(G462), .b(G465), .O(G540) );
nand2 gate144( .a(G468), .b(G471), .O(G543) );
nand2 gate145( .a(G474), .b(G477), .O(G546) );
nand2 gate146( .a(G480), .b(G483), .O(G549) );
nand2 gate147( .a(G486), .b(G489), .O(G552) );

  xor2  gate603(.a(G495), .b(G492), .O(gate148inter0));
  nand2 gate604(.a(gate148inter0), .b(s_8), .O(gate148inter1));
  and2  gate605(.a(G495), .b(G492), .O(gate148inter2));
  inv1  gate606(.a(s_8), .O(gate148inter3));
  inv1  gate607(.a(s_9), .O(gate148inter4));
  nand2 gate608(.a(gate148inter4), .b(gate148inter3), .O(gate148inter5));
  nor2  gate609(.a(gate148inter5), .b(gate148inter2), .O(gate148inter6));
  inv1  gate610(.a(G492), .O(gate148inter7));
  inv1  gate611(.a(G495), .O(gate148inter8));
  nand2 gate612(.a(gate148inter8), .b(gate148inter7), .O(gate148inter9));
  nand2 gate613(.a(s_9), .b(gate148inter3), .O(gate148inter10));
  nor2  gate614(.a(gate148inter10), .b(gate148inter9), .O(gate148inter11));
  nor2  gate615(.a(gate148inter11), .b(gate148inter6), .O(gate148inter12));
  nand2 gate616(.a(gate148inter12), .b(gate148inter1), .O(G555));
nand2 gate149( .a(G498), .b(G501), .O(G558) );
nand2 gate150( .a(G504), .b(G507), .O(G561) );
nand2 gate151( .a(G510), .b(G513), .O(G564) );
nand2 gate152( .a(G516), .b(G519), .O(G567) );

  xor2  gate673(.a(G522), .b(G426), .O(gate153inter0));
  nand2 gate674(.a(gate153inter0), .b(s_18), .O(gate153inter1));
  and2  gate675(.a(G522), .b(G426), .O(gate153inter2));
  inv1  gate676(.a(s_18), .O(gate153inter3));
  inv1  gate677(.a(s_19), .O(gate153inter4));
  nand2 gate678(.a(gate153inter4), .b(gate153inter3), .O(gate153inter5));
  nor2  gate679(.a(gate153inter5), .b(gate153inter2), .O(gate153inter6));
  inv1  gate680(.a(G426), .O(gate153inter7));
  inv1  gate681(.a(G522), .O(gate153inter8));
  nand2 gate682(.a(gate153inter8), .b(gate153inter7), .O(gate153inter9));
  nand2 gate683(.a(s_19), .b(gate153inter3), .O(gate153inter10));
  nor2  gate684(.a(gate153inter10), .b(gate153inter9), .O(gate153inter11));
  nor2  gate685(.a(gate153inter11), .b(gate153inter6), .O(gate153inter12));
  nand2 gate686(.a(gate153inter12), .b(gate153inter1), .O(G570));
nand2 gate154( .a(G429), .b(G522), .O(G571) );
nand2 gate155( .a(G432), .b(G525), .O(G572) );
nand2 gate156( .a(G435), .b(G525), .O(G573) );

  xor2  gate1303(.a(G528), .b(G438), .O(gate157inter0));
  nand2 gate1304(.a(gate157inter0), .b(s_108), .O(gate157inter1));
  and2  gate1305(.a(G528), .b(G438), .O(gate157inter2));
  inv1  gate1306(.a(s_108), .O(gate157inter3));
  inv1  gate1307(.a(s_109), .O(gate157inter4));
  nand2 gate1308(.a(gate157inter4), .b(gate157inter3), .O(gate157inter5));
  nor2  gate1309(.a(gate157inter5), .b(gate157inter2), .O(gate157inter6));
  inv1  gate1310(.a(G438), .O(gate157inter7));
  inv1  gate1311(.a(G528), .O(gate157inter8));
  nand2 gate1312(.a(gate157inter8), .b(gate157inter7), .O(gate157inter9));
  nand2 gate1313(.a(s_109), .b(gate157inter3), .O(gate157inter10));
  nor2  gate1314(.a(gate157inter10), .b(gate157inter9), .O(gate157inter11));
  nor2  gate1315(.a(gate157inter11), .b(gate157inter6), .O(gate157inter12));
  nand2 gate1316(.a(gate157inter12), .b(gate157inter1), .O(G574));
nand2 gate158( .a(G441), .b(G528), .O(G575) );
nand2 gate159( .a(G444), .b(G531), .O(G576) );

  xor2  gate715(.a(G531), .b(G447), .O(gate160inter0));
  nand2 gate716(.a(gate160inter0), .b(s_24), .O(gate160inter1));
  and2  gate717(.a(G531), .b(G447), .O(gate160inter2));
  inv1  gate718(.a(s_24), .O(gate160inter3));
  inv1  gate719(.a(s_25), .O(gate160inter4));
  nand2 gate720(.a(gate160inter4), .b(gate160inter3), .O(gate160inter5));
  nor2  gate721(.a(gate160inter5), .b(gate160inter2), .O(gate160inter6));
  inv1  gate722(.a(G447), .O(gate160inter7));
  inv1  gate723(.a(G531), .O(gate160inter8));
  nand2 gate724(.a(gate160inter8), .b(gate160inter7), .O(gate160inter9));
  nand2 gate725(.a(s_25), .b(gate160inter3), .O(gate160inter10));
  nor2  gate726(.a(gate160inter10), .b(gate160inter9), .O(gate160inter11));
  nor2  gate727(.a(gate160inter11), .b(gate160inter6), .O(gate160inter12));
  nand2 gate728(.a(gate160inter12), .b(gate160inter1), .O(G577));
nand2 gate161( .a(G450), .b(G534), .O(G578) );
nand2 gate162( .a(G453), .b(G534), .O(G579) );
nand2 gate163( .a(G456), .b(G537), .O(G580) );

  xor2  gate981(.a(G537), .b(G459), .O(gate164inter0));
  nand2 gate982(.a(gate164inter0), .b(s_62), .O(gate164inter1));
  and2  gate983(.a(G537), .b(G459), .O(gate164inter2));
  inv1  gate984(.a(s_62), .O(gate164inter3));
  inv1  gate985(.a(s_63), .O(gate164inter4));
  nand2 gate986(.a(gate164inter4), .b(gate164inter3), .O(gate164inter5));
  nor2  gate987(.a(gate164inter5), .b(gate164inter2), .O(gate164inter6));
  inv1  gate988(.a(G459), .O(gate164inter7));
  inv1  gate989(.a(G537), .O(gate164inter8));
  nand2 gate990(.a(gate164inter8), .b(gate164inter7), .O(gate164inter9));
  nand2 gate991(.a(s_63), .b(gate164inter3), .O(gate164inter10));
  nor2  gate992(.a(gate164inter10), .b(gate164inter9), .O(gate164inter11));
  nor2  gate993(.a(gate164inter11), .b(gate164inter6), .O(gate164inter12));
  nand2 gate994(.a(gate164inter12), .b(gate164inter1), .O(G581));
nand2 gate165( .a(G462), .b(G540), .O(G582) );
nand2 gate166( .a(G465), .b(G540), .O(G583) );
nand2 gate167( .a(G468), .b(G543), .O(G584) );
nand2 gate168( .a(G471), .b(G543), .O(G585) );
nand2 gate169( .a(G474), .b(G546), .O(G586) );

  xor2  gate701(.a(G546), .b(G477), .O(gate170inter0));
  nand2 gate702(.a(gate170inter0), .b(s_22), .O(gate170inter1));
  and2  gate703(.a(G546), .b(G477), .O(gate170inter2));
  inv1  gate704(.a(s_22), .O(gate170inter3));
  inv1  gate705(.a(s_23), .O(gate170inter4));
  nand2 gate706(.a(gate170inter4), .b(gate170inter3), .O(gate170inter5));
  nor2  gate707(.a(gate170inter5), .b(gate170inter2), .O(gate170inter6));
  inv1  gate708(.a(G477), .O(gate170inter7));
  inv1  gate709(.a(G546), .O(gate170inter8));
  nand2 gate710(.a(gate170inter8), .b(gate170inter7), .O(gate170inter9));
  nand2 gate711(.a(s_23), .b(gate170inter3), .O(gate170inter10));
  nor2  gate712(.a(gate170inter10), .b(gate170inter9), .O(gate170inter11));
  nor2  gate713(.a(gate170inter11), .b(gate170inter6), .O(gate170inter12));
  nand2 gate714(.a(gate170inter12), .b(gate170inter1), .O(G587));
nand2 gate171( .a(G480), .b(G549), .O(G588) );
nand2 gate172( .a(G483), .b(G549), .O(G589) );
nand2 gate173( .a(G486), .b(G552), .O(G590) );
nand2 gate174( .a(G489), .b(G552), .O(G591) );
nand2 gate175( .a(G492), .b(G555), .O(G592) );
nand2 gate176( .a(G495), .b(G555), .O(G593) );
nand2 gate177( .a(G498), .b(G558), .O(G594) );
nand2 gate178( .a(G501), .b(G558), .O(G595) );
nand2 gate179( .a(G504), .b(G561), .O(G596) );
nand2 gate180( .a(G507), .b(G561), .O(G597) );
nand2 gate181( .a(G510), .b(G564), .O(G598) );
nand2 gate182( .a(G513), .b(G564), .O(G599) );
nand2 gate183( .a(G516), .b(G567), .O(G600) );

  xor2  gate1345(.a(G567), .b(G519), .O(gate184inter0));
  nand2 gate1346(.a(gate184inter0), .b(s_114), .O(gate184inter1));
  and2  gate1347(.a(G567), .b(G519), .O(gate184inter2));
  inv1  gate1348(.a(s_114), .O(gate184inter3));
  inv1  gate1349(.a(s_115), .O(gate184inter4));
  nand2 gate1350(.a(gate184inter4), .b(gate184inter3), .O(gate184inter5));
  nor2  gate1351(.a(gate184inter5), .b(gate184inter2), .O(gate184inter6));
  inv1  gate1352(.a(G519), .O(gate184inter7));
  inv1  gate1353(.a(G567), .O(gate184inter8));
  nand2 gate1354(.a(gate184inter8), .b(gate184inter7), .O(gate184inter9));
  nand2 gate1355(.a(s_115), .b(gate184inter3), .O(gate184inter10));
  nor2  gate1356(.a(gate184inter10), .b(gate184inter9), .O(gate184inter11));
  nor2  gate1357(.a(gate184inter11), .b(gate184inter6), .O(gate184inter12));
  nand2 gate1358(.a(gate184inter12), .b(gate184inter1), .O(G601));
nand2 gate185( .a(G570), .b(G571), .O(G602) );
nand2 gate186( .a(G572), .b(G573), .O(G607) );
nand2 gate187( .a(G574), .b(G575), .O(G612) );
nand2 gate188( .a(G576), .b(G577), .O(G617) );
nand2 gate189( .a(G578), .b(G579), .O(G622) );

  xor2  gate1051(.a(G581), .b(G580), .O(gate190inter0));
  nand2 gate1052(.a(gate190inter0), .b(s_72), .O(gate190inter1));
  and2  gate1053(.a(G581), .b(G580), .O(gate190inter2));
  inv1  gate1054(.a(s_72), .O(gate190inter3));
  inv1  gate1055(.a(s_73), .O(gate190inter4));
  nand2 gate1056(.a(gate190inter4), .b(gate190inter3), .O(gate190inter5));
  nor2  gate1057(.a(gate190inter5), .b(gate190inter2), .O(gate190inter6));
  inv1  gate1058(.a(G580), .O(gate190inter7));
  inv1  gate1059(.a(G581), .O(gate190inter8));
  nand2 gate1060(.a(gate190inter8), .b(gate190inter7), .O(gate190inter9));
  nand2 gate1061(.a(s_73), .b(gate190inter3), .O(gate190inter10));
  nor2  gate1062(.a(gate190inter10), .b(gate190inter9), .O(gate190inter11));
  nor2  gate1063(.a(gate190inter11), .b(gate190inter6), .O(gate190inter12));
  nand2 gate1064(.a(gate190inter12), .b(gate190inter1), .O(G627));

  xor2  gate1191(.a(G583), .b(G582), .O(gate191inter0));
  nand2 gate1192(.a(gate191inter0), .b(s_92), .O(gate191inter1));
  and2  gate1193(.a(G583), .b(G582), .O(gate191inter2));
  inv1  gate1194(.a(s_92), .O(gate191inter3));
  inv1  gate1195(.a(s_93), .O(gate191inter4));
  nand2 gate1196(.a(gate191inter4), .b(gate191inter3), .O(gate191inter5));
  nor2  gate1197(.a(gate191inter5), .b(gate191inter2), .O(gate191inter6));
  inv1  gate1198(.a(G582), .O(gate191inter7));
  inv1  gate1199(.a(G583), .O(gate191inter8));
  nand2 gate1200(.a(gate191inter8), .b(gate191inter7), .O(gate191inter9));
  nand2 gate1201(.a(s_93), .b(gate191inter3), .O(gate191inter10));
  nor2  gate1202(.a(gate191inter10), .b(gate191inter9), .O(gate191inter11));
  nor2  gate1203(.a(gate191inter11), .b(gate191inter6), .O(gate191inter12));
  nand2 gate1204(.a(gate191inter12), .b(gate191inter1), .O(G632));

  xor2  gate687(.a(G585), .b(G584), .O(gate192inter0));
  nand2 gate688(.a(gate192inter0), .b(s_20), .O(gate192inter1));
  and2  gate689(.a(G585), .b(G584), .O(gate192inter2));
  inv1  gate690(.a(s_20), .O(gate192inter3));
  inv1  gate691(.a(s_21), .O(gate192inter4));
  nand2 gate692(.a(gate192inter4), .b(gate192inter3), .O(gate192inter5));
  nor2  gate693(.a(gate192inter5), .b(gate192inter2), .O(gate192inter6));
  inv1  gate694(.a(G584), .O(gate192inter7));
  inv1  gate695(.a(G585), .O(gate192inter8));
  nand2 gate696(.a(gate192inter8), .b(gate192inter7), .O(gate192inter9));
  nand2 gate697(.a(s_21), .b(gate192inter3), .O(gate192inter10));
  nor2  gate698(.a(gate192inter10), .b(gate192inter9), .O(gate192inter11));
  nor2  gate699(.a(gate192inter11), .b(gate192inter6), .O(gate192inter12));
  nand2 gate700(.a(gate192inter12), .b(gate192inter1), .O(G637));

  xor2  gate617(.a(G587), .b(G586), .O(gate193inter0));
  nand2 gate618(.a(gate193inter0), .b(s_10), .O(gate193inter1));
  and2  gate619(.a(G587), .b(G586), .O(gate193inter2));
  inv1  gate620(.a(s_10), .O(gate193inter3));
  inv1  gate621(.a(s_11), .O(gate193inter4));
  nand2 gate622(.a(gate193inter4), .b(gate193inter3), .O(gate193inter5));
  nor2  gate623(.a(gate193inter5), .b(gate193inter2), .O(gate193inter6));
  inv1  gate624(.a(G586), .O(gate193inter7));
  inv1  gate625(.a(G587), .O(gate193inter8));
  nand2 gate626(.a(gate193inter8), .b(gate193inter7), .O(gate193inter9));
  nand2 gate627(.a(s_11), .b(gate193inter3), .O(gate193inter10));
  nor2  gate628(.a(gate193inter10), .b(gate193inter9), .O(gate193inter11));
  nor2  gate629(.a(gate193inter11), .b(gate193inter6), .O(gate193inter12));
  nand2 gate630(.a(gate193inter12), .b(gate193inter1), .O(G642));
nand2 gate194( .a(G588), .b(G589), .O(G645) );
nand2 gate195( .a(G590), .b(G591), .O(G648) );
nand2 gate196( .a(G592), .b(G593), .O(G651) );
nand2 gate197( .a(G594), .b(G595), .O(G654) );
nand2 gate198( .a(G596), .b(G597), .O(G657) );
nand2 gate199( .a(G598), .b(G599), .O(G660) );
nand2 gate200( .a(G600), .b(G601), .O(G663) );

  xor2  gate1205(.a(G607), .b(G602), .O(gate201inter0));
  nand2 gate1206(.a(gate201inter0), .b(s_94), .O(gate201inter1));
  and2  gate1207(.a(G607), .b(G602), .O(gate201inter2));
  inv1  gate1208(.a(s_94), .O(gate201inter3));
  inv1  gate1209(.a(s_95), .O(gate201inter4));
  nand2 gate1210(.a(gate201inter4), .b(gate201inter3), .O(gate201inter5));
  nor2  gate1211(.a(gate201inter5), .b(gate201inter2), .O(gate201inter6));
  inv1  gate1212(.a(G602), .O(gate201inter7));
  inv1  gate1213(.a(G607), .O(gate201inter8));
  nand2 gate1214(.a(gate201inter8), .b(gate201inter7), .O(gate201inter9));
  nand2 gate1215(.a(s_95), .b(gate201inter3), .O(gate201inter10));
  nor2  gate1216(.a(gate201inter10), .b(gate201inter9), .O(gate201inter11));
  nor2  gate1217(.a(gate201inter11), .b(gate201inter6), .O(gate201inter12));
  nand2 gate1218(.a(gate201inter12), .b(gate201inter1), .O(G666));
nand2 gate202( .a(G612), .b(G617), .O(G669) );
nand2 gate203( .a(G602), .b(G612), .O(G672) );
nand2 gate204( .a(G607), .b(G617), .O(G675) );
nand2 gate205( .a(G622), .b(G627), .O(G678) );
nand2 gate206( .a(G632), .b(G637), .O(G681) );
nand2 gate207( .a(G622), .b(G632), .O(G684) );
nand2 gate208( .a(G627), .b(G637), .O(G687) );
nand2 gate209( .a(G602), .b(G666), .O(G690) );
nand2 gate210( .a(G607), .b(G666), .O(G691) );

  xor2  gate1219(.a(G669), .b(G612), .O(gate211inter0));
  nand2 gate1220(.a(gate211inter0), .b(s_96), .O(gate211inter1));
  and2  gate1221(.a(G669), .b(G612), .O(gate211inter2));
  inv1  gate1222(.a(s_96), .O(gate211inter3));
  inv1  gate1223(.a(s_97), .O(gate211inter4));
  nand2 gate1224(.a(gate211inter4), .b(gate211inter3), .O(gate211inter5));
  nor2  gate1225(.a(gate211inter5), .b(gate211inter2), .O(gate211inter6));
  inv1  gate1226(.a(G612), .O(gate211inter7));
  inv1  gate1227(.a(G669), .O(gate211inter8));
  nand2 gate1228(.a(gate211inter8), .b(gate211inter7), .O(gate211inter9));
  nand2 gate1229(.a(s_97), .b(gate211inter3), .O(gate211inter10));
  nor2  gate1230(.a(gate211inter10), .b(gate211inter9), .O(gate211inter11));
  nor2  gate1231(.a(gate211inter11), .b(gate211inter6), .O(gate211inter12));
  nand2 gate1232(.a(gate211inter12), .b(gate211inter1), .O(G692));

  xor2  gate785(.a(G669), .b(G617), .O(gate212inter0));
  nand2 gate786(.a(gate212inter0), .b(s_34), .O(gate212inter1));
  and2  gate787(.a(G669), .b(G617), .O(gate212inter2));
  inv1  gate788(.a(s_34), .O(gate212inter3));
  inv1  gate789(.a(s_35), .O(gate212inter4));
  nand2 gate790(.a(gate212inter4), .b(gate212inter3), .O(gate212inter5));
  nor2  gate791(.a(gate212inter5), .b(gate212inter2), .O(gate212inter6));
  inv1  gate792(.a(G617), .O(gate212inter7));
  inv1  gate793(.a(G669), .O(gate212inter8));
  nand2 gate794(.a(gate212inter8), .b(gate212inter7), .O(gate212inter9));
  nand2 gate795(.a(s_35), .b(gate212inter3), .O(gate212inter10));
  nor2  gate796(.a(gate212inter10), .b(gate212inter9), .O(gate212inter11));
  nor2  gate797(.a(gate212inter11), .b(gate212inter6), .O(gate212inter12));
  nand2 gate798(.a(gate212inter12), .b(gate212inter1), .O(G693));
nand2 gate213( .a(G602), .b(G672), .O(G694) );

  xor2  gate729(.a(G672), .b(G612), .O(gate214inter0));
  nand2 gate730(.a(gate214inter0), .b(s_26), .O(gate214inter1));
  and2  gate731(.a(G672), .b(G612), .O(gate214inter2));
  inv1  gate732(.a(s_26), .O(gate214inter3));
  inv1  gate733(.a(s_27), .O(gate214inter4));
  nand2 gate734(.a(gate214inter4), .b(gate214inter3), .O(gate214inter5));
  nor2  gate735(.a(gate214inter5), .b(gate214inter2), .O(gate214inter6));
  inv1  gate736(.a(G612), .O(gate214inter7));
  inv1  gate737(.a(G672), .O(gate214inter8));
  nand2 gate738(.a(gate214inter8), .b(gate214inter7), .O(gate214inter9));
  nand2 gate739(.a(s_27), .b(gate214inter3), .O(gate214inter10));
  nor2  gate740(.a(gate214inter10), .b(gate214inter9), .O(gate214inter11));
  nor2  gate741(.a(gate214inter11), .b(gate214inter6), .O(gate214inter12));
  nand2 gate742(.a(gate214inter12), .b(gate214inter1), .O(G695));
nand2 gate215( .a(G607), .b(G675), .O(G696) );

  xor2  gate645(.a(G675), .b(G617), .O(gate216inter0));
  nand2 gate646(.a(gate216inter0), .b(s_14), .O(gate216inter1));
  and2  gate647(.a(G675), .b(G617), .O(gate216inter2));
  inv1  gate648(.a(s_14), .O(gate216inter3));
  inv1  gate649(.a(s_15), .O(gate216inter4));
  nand2 gate650(.a(gate216inter4), .b(gate216inter3), .O(gate216inter5));
  nor2  gate651(.a(gate216inter5), .b(gate216inter2), .O(gate216inter6));
  inv1  gate652(.a(G617), .O(gate216inter7));
  inv1  gate653(.a(G675), .O(gate216inter8));
  nand2 gate654(.a(gate216inter8), .b(gate216inter7), .O(gate216inter9));
  nand2 gate655(.a(s_15), .b(gate216inter3), .O(gate216inter10));
  nor2  gate656(.a(gate216inter10), .b(gate216inter9), .O(gate216inter11));
  nor2  gate657(.a(gate216inter11), .b(gate216inter6), .O(gate216inter12));
  nand2 gate658(.a(gate216inter12), .b(gate216inter1), .O(G697));

  xor2  gate1037(.a(G678), .b(G622), .O(gate217inter0));
  nand2 gate1038(.a(gate217inter0), .b(s_70), .O(gate217inter1));
  and2  gate1039(.a(G678), .b(G622), .O(gate217inter2));
  inv1  gate1040(.a(s_70), .O(gate217inter3));
  inv1  gate1041(.a(s_71), .O(gate217inter4));
  nand2 gate1042(.a(gate217inter4), .b(gate217inter3), .O(gate217inter5));
  nor2  gate1043(.a(gate217inter5), .b(gate217inter2), .O(gate217inter6));
  inv1  gate1044(.a(G622), .O(gate217inter7));
  inv1  gate1045(.a(G678), .O(gate217inter8));
  nand2 gate1046(.a(gate217inter8), .b(gate217inter7), .O(gate217inter9));
  nand2 gate1047(.a(s_71), .b(gate217inter3), .O(gate217inter10));
  nor2  gate1048(.a(gate217inter10), .b(gate217inter9), .O(gate217inter11));
  nor2  gate1049(.a(gate217inter11), .b(gate217inter6), .O(gate217inter12));
  nand2 gate1050(.a(gate217inter12), .b(gate217inter1), .O(G698));

  xor2  gate1149(.a(G678), .b(G627), .O(gate218inter0));
  nand2 gate1150(.a(gate218inter0), .b(s_86), .O(gate218inter1));
  and2  gate1151(.a(G678), .b(G627), .O(gate218inter2));
  inv1  gate1152(.a(s_86), .O(gate218inter3));
  inv1  gate1153(.a(s_87), .O(gate218inter4));
  nand2 gate1154(.a(gate218inter4), .b(gate218inter3), .O(gate218inter5));
  nor2  gate1155(.a(gate218inter5), .b(gate218inter2), .O(gate218inter6));
  inv1  gate1156(.a(G627), .O(gate218inter7));
  inv1  gate1157(.a(G678), .O(gate218inter8));
  nand2 gate1158(.a(gate218inter8), .b(gate218inter7), .O(gate218inter9));
  nand2 gate1159(.a(s_87), .b(gate218inter3), .O(gate218inter10));
  nor2  gate1160(.a(gate218inter10), .b(gate218inter9), .O(gate218inter11));
  nor2  gate1161(.a(gate218inter11), .b(gate218inter6), .O(gate218inter12));
  nand2 gate1162(.a(gate218inter12), .b(gate218inter1), .O(G699));
nand2 gate219( .a(G632), .b(G681), .O(G700) );
nand2 gate220( .a(G637), .b(G681), .O(G701) );
nand2 gate221( .a(G622), .b(G684), .O(G702) );
nand2 gate222( .a(G632), .b(G684), .O(G703) );
nand2 gate223( .a(G627), .b(G687), .O(G704) );
nand2 gate224( .a(G637), .b(G687), .O(G705) );
nand2 gate225( .a(G690), .b(G691), .O(G706) );

  xor2  gate1261(.a(G693), .b(G692), .O(gate226inter0));
  nand2 gate1262(.a(gate226inter0), .b(s_102), .O(gate226inter1));
  and2  gate1263(.a(G693), .b(G692), .O(gate226inter2));
  inv1  gate1264(.a(s_102), .O(gate226inter3));
  inv1  gate1265(.a(s_103), .O(gate226inter4));
  nand2 gate1266(.a(gate226inter4), .b(gate226inter3), .O(gate226inter5));
  nor2  gate1267(.a(gate226inter5), .b(gate226inter2), .O(gate226inter6));
  inv1  gate1268(.a(G692), .O(gate226inter7));
  inv1  gate1269(.a(G693), .O(gate226inter8));
  nand2 gate1270(.a(gate226inter8), .b(gate226inter7), .O(gate226inter9));
  nand2 gate1271(.a(s_103), .b(gate226inter3), .O(gate226inter10));
  nor2  gate1272(.a(gate226inter10), .b(gate226inter9), .O(gate226inter11));
  nor2  gate1273(.a(gate226inter11), .b(gate226inter6), .O(gate226inter12));
  nand2 gate1274(.a(gate226inter12), .b(gate226inter1), .O(G709));
nand2 gate227( .a(G694), .b(G695), .O(G712) );

  xor2  gate1359(.a(G697), .b(G696), .O(gate228inter0));
  nand2 gate1360(.a(gate228inter0), .b(s_116), .O(gate228inter1));
  and2  gate1361(.a(G697), .b(G696), .O(gate228inter2));
  inv1  gate1362(.a(s_116), .O(gate228inter3));
  inv1  gate1363(.a(s_117), .O(gate228inter4));
  nand2 gate1364(.a(gate228inter4), .b(gate228inter3), .O(gate228inter5));
  nor2  gate1365(.a(gate228inter5), .b(gate228inter2), .O(gate228inter6));
  inv1  gate1366(.a(G696), .O(gate228inter7));
  inv1  gate1367(.a(G697), .O(gate228inter8));
  nand2 gate1368(.a(gate228inter8), .b(gate228inter7), .O(gate228inter9));
  nand2 gate1369(.a(s_117), .b(gate228inter3), .O(gate228inter10));
  nor2  gate1370(.a(gate228inter10), .b(gate228inter9), .O(gate228inter11));
  nor2  gate1371(.a(gate228inter11), .b(gate228inter6), .O(gate228inter12));
  nand2 gate1372(.a(gate228inter12), .b(gate228inter1), .O(G715));
nand2 gate229( .a(G698), .b(G699), .O(G718) );
nand2 gate230( .a(G700), .b(G701), .O(G721) );
nand2 gate231( .a(G702), .b(G703), .O(G724) );
nand2 gate232( .a(G704), .b(G705), .O(G727) );
nand2 gate233( .a(G242), .b(G718), .O(G730) );
nand2 gate234( .a(G245), .b(G721), .O(G733) );
nand2 gate235( .a(G248), .b(G724), .O(G736) );
nand2 gate236( .a(G251), .b(G727), .O(G739) );
nand2 gate237( .a(G254), .b(G706), .O(G742) );
nand2 gate238( .a(G257), .b(G709), .O(G745) );
nand2 gate239( .a(G260), .b(G712), .O(G748) );
nand2 gate240( .a(G263), .b(G715), .O(G751) );
nand2 gate241( .a(G242), .b(G730), .O(G754) );
nand2 gate242( .a(G718), .b(G730), .O(G755) );
nand2 gate243( .a(G245), .b(G733), .O(G756) );
nand2 gate244( .a(G721), .b(G733), .O(G757) );
nand2 gate245( .a(G248), .b(G736), .O(G758) );
nand2 gate246( .a(G724), .b(G736), .O(G759) );

  xor2  gate855(.a(G739), .b(G251), .O(gate247inter0));
  nand2 gate856(.a(gate247inter0), .b(s_44), .O(gate247inter1));
  and2  gate857(.a(G739), .b(G251), .O(gate247inter2));
  inv1  gate858(.a(s_44), .O(gate247inter3));
  inv1  gate859(.a(s_45), .O(gate247inter4));
  nand2 gate860(.a(gate247inter4), .b(gate247inter3), .O(gate247inter5));
  nor2  gate861(.a(gate247inter5), .b(gate247inter2), .O(gate247inter6));
  inv1  gate862(.a(G251), .O(gate247inter7));
  inv1  gate863(.a(G739), .O(gate247inter8));
  nand2 gate864(.a(gate247inter8), .b(gate247inter7), .O(gate247inter9));
  nand2 gate865(.a(s_45), .b(gate247inter3), .O(gate247inter10));
  nor2  gate866(.a(gate247inter10), .b(gate247inter9), .O(gate247inter11));
  nor2  gate867(.a(gate247inter11), .b(gate247inter6), .O(gate247inter12));
  nand2 gate868(.a(gate247inter12), .b(gate247inter1), .O(G760));
nand2 gate248( .a(G727), .b(G739), .O(G761) );
nand2 gate249( .a(G254), .b(G742), .O(G762) );

  xor2  gate1401(.a(G742), .b(G706), .O(gate250inter0));
  nand2 gate1402(.a(gate250inter0), .b(s_122), .O(gate250inter1));
  and2  gate1403(.a(G742), .b(G706), .O(gate250inter2));
  inv1  gate1404(.a(s_122), .O(gate250inter3));
  inv1  gate1405(.a(s_123), .O(gate250inter4));
  nand2 gate1406(.a(gate250inter4), .b(gate250inter3), .O(gate250inter5));
  nor2  gate1407(.a(gate250inter5), .b(gate250inter2), .O(gate250inter6));
  inv1  gate1408(.a(G706), .O(gate250inter7));
  inv1  gate1409(.a(G742), .O(gate250inter8));
  nand2 gate1410(.a(gate250inter8), .b(gate250inter7), .O(gate250inter9));
  nand2 gate1411(.a(s_123), .b(gate250inter3), .O(gate250inter10));
  nor2  gate1412(.a(gate250inter10), .b(gate250inter9), .O(gate250inter11));
  nor2  gate1413(.a(gate250inter11), .b(gate250inter6), .O(gate250inter12));
  nand2 gate1414(.a(gate250inter12), .b(gate250inter1), .O(G763));
nand2 gate251( .a(G257), .b(G745), .O(G764) );
nand2 gate252( .a(G709), .b(G745), .O(G765) );
nand2 gate253( .a(G260), .b(G748), .O(G766) );

  xor2  gate1415(.a(G748), .b(G712), .O(gate254inter0));
  nand2 gate1416(.a(gate254inter0), .b(s_124), .O(gate254inter1));
  and2  gate1417(.a(G748), .b(G712), .O(gate254inter2));
  inv1  gate1418(.a(s_124), .O(gate254inter3));
  inv1  gate1419(.a(s_125), .O(gate254inter4));
  nand2 gate1420(.a(gate254inter4), .b(gate254inter3), .O(gate254inter5));
  nor2  gate1421(.a(gate254inter5), .b(gate254inter2), .O(gate254inter6));
  inv1  gate1422(.a(G712), .O(gate254inter7));
  inv1  gate1423(.a(G748), .O(gate254inter8));
  nand2 gate1424(.a(gate254inter8), .b(gate254inter7), .O(gate254inter9));
  nand2 gate1425(.a(s_125), .b(gate254inter3), .O(gate254inter10));
  nor2  gate1426(.a(gate254inter10), .b(gate254inter9), .O(gate254inter11));
  nor2  gate1427(.a(gate254inter11), .b(gate254inter6), .O(gate254inter12));
  nand2 gate1428(.a(gate254inter12), .b(gate254inter1), .O(G767));
nand2 gate255( .a(G263), .b(G751), .O(G768) );
nand2 gate256( .a(G715), .b(G751), .O(G769) );
nand2 gate257( .a(G754), .b(G755), .O(G770) );
nand2 gate258( .a(G756), .b(G757), .O(G773) );
nand2 gate259( .a(G758), .b(G759), .O(G776) );
nand2 gate260( .a(G760), .b(G761), .O(G779) );
nand2 gate261( .a(G762), .b(G763), .O(G782) );
nand2 gate262( .a(G764), .b(G765), .O(G785) );

  xor2  gate547(.a(G767), .b(G766), .O(gate263inter0));
  nand2 gate548(.a(gate263inter0), .b(s_0), .O(gate263inter1));
  and2  gate549(.a(G767), .b(G766), .O(gate263inter2));
  inv1  gate550(.a(s_0), .O(gate263inter3));
  inv1  gate551(.a(s_1), .O(gate263inter4));
  nand2 gate552(.a(gate263inter4), .b(gate263inter3), .O(gate263inter5));
  nor2  gate553(.a(gate263inter5), .b(gate263inter2), .O(gate263inter6));
  inv1  gate554(.a(G766), .O(gate263inter7));
  inv1  gate555(.a(G767), .O(gate263inter8));
  nand2 gate556(.a(gate263inter8), .b(gate263inter7), .O(gate263inter9));
  nand2 gate557(.a(s_1), .b(gate263inter3), .O(gate263inter10));
  nor2  gate558(.a(gate263inter10), .b(gate263inter9), .O(gate263inter11));
  nor2  gate559(.a(gate263inter11), .b(gate263inter6), .O(gate263inter12));
  nand2 gate560(.a(gate263inter12), .b(gate263inter1), .O(G788));

  xor2  gate1079(.a(G769), .b(G768), .O(gate264inter0));
  nand2 gate1080(.a(gate264inter0), .b(s_76), .O(gate264inter1));
  and2  gate1081(.a(G769), .b(G768), .O(gate264inter2));
  inv1  gate1082(.a(s_76), .O(gate264inter3));
  inv1  gate1083(.a(s_77), .O(gate264inter4));
  nand2 gate1084(.a(gate264inter4), .b(gate264inter3), .O(gate264inter5));
  nor2  gate1085(.a(gate264inter5), .b(gate264inter2), .O(gate264inter6));
  inv1  gate1086(.a(G768), .O(gate264inter7));
  inv1  gate1087(.a(G769), .O(gate264inter8));
  nand2 gate1088(.a(gate264inter8), .b(gate264inter7), .O(gate264inter9));
  nand2 gate1089(.a(s_77), .b(gate264inter3), .O(gate264inter10));
  nor2  gate1090(.a(gate264inter10), .b(gate264inter9), .O(gate264inter11));
  nor2  gate1091(.a(gate264inter11), .b(gate264inter6), .O(gate264inter12));
  nand2 gate1092(.a(gate264inter12), .b(gate264inter1), .O(G791));
nand2 gate265( .a(G642), .b(G770), .O(G794) );
nand2 gate266( .a(G645), .b(G773), .O(G797) );
nand2 gate267( .a(G648), .b(G776), .O(G800) );
nand2 gate268( .a(G651), .b(G779), .O(G803) );

  xor2  gate911(.a(G782), .b(G654), .O(gate269inter0));
  nand2 gate912(.a(gate269inter0), .b(s_52), .O(gate269inter1));
  and2  gate913(.a(G782), .b(G654), .O(gate269inter2));
  inv1  gate914(.a(s_52), .O(gate269inter3));
  inv1  gate915(.a(s_53), .O(gate269inter4));
  nand2 gate916(.a(gate269inter4), .b(gate269inter3), .O(gate269inter5));
  nor2  gate917(.a(gate269inter5), .b(gate269inter2), .O(gate269inter6));
  inv1  gate918(.a(G654), .O(gate269inter7));
  inv1  gate919(.a(G782), .O(gate269inter8));
  nand2 gate920(.a(gate269inter8), .b(gate269inter7), .O(gate269inter9));
  nand2 gate921(.a(s_53), .b(gate269inter3), .O(gate269inter10));
  nor2  gate922(.a(gate269inter10), .b(gate269inter9), .O(gate269inter11));
  nor2  gate923(.a(gate269inter11), .b(gate269inter6), .O(gate269inter12));
  nand2 gate924(.a(gate269inter12), .b(gate269inter1), .O(G806));
nand2 gate270( .a(G657), .b(G785), .O(G809) );

  xor2  gate1289(.a(G788), .b(G660), .O(gate271inter0));
  nand2 gate1290(.a(gate271inter0), .b(s_106), .O(gate271inter1));
  and2  gate1291(.a(G788), .b(G660), .O(gate271inter2));
  inv1  gate1292(.a(s_106), .O(gate271inter3));
  inv1  gate1293(.a(s_107), .O(gate271inter4));
  nand2 gate1294(.a(gate271inter4), .b(gate271inter3), .O(gate271inter5));
  nor2  gate1295(.a(gate271inter5), .b(gate271inter2), .O(gate271inter6));
  inv1  gate1296(.a(G660), .O(gate271inter7));
  inv1  gate1297(.a(G788), .O(gate271inter8));
  nand2 gate1298(.a(gate271inter8), .b(gate271inter7), .O(gate271inter9));
  nand2 gate1299(.a(s_107), .b(gate271inter3), .O(gate271inter10));
  nor2  gate1300(.a(gate271inter10), .b(gate271inter9), .O(gate271inter11));
  nor2  gate1301(.a(gate271inter11), .b(gate271inter6), .O(gate271inter12));
  nand2 gate1302(.a(gate271inter12), .b(gate271inter1), .O(G812));

  xor2  gate925(.a(G791), .b(G663), .O(gate272inter0));
  nand2 gate926(.a(gate272inter0), .b(s_54), .O(gate272inter1));
  and2  gate927(.a(G791), .b(G663), .O(gate272inter2));
  inv1  gate928(.a(s_54), .O(gate272inter3));
  inv1  gate929(.a(s_55), .O(gate272inter4));
  nand2 gate930(.a(gate272inter4), .b(gate272inter3), .O(gate272inter5));
  nor2  gate931(.a(gate272inter5), .b(gate272inter2), .O(gate272inter6));
  inv1  gate932(.a(G663), .O(gate272inter7));
  inv1  gate933(.a(G791), .O(gate272inter8));
  nand2 gate934(.a(gate272inter8), .b(gate272inter7), .O(gate272inter9));
  nand2 gate935(.a(s_55), .b(gate272inter3), .O(gate272inter10));
  nor2  gate936(.a(gate272inter10), .b(gate272inter9), .O(gate272inter11));
  nor2  gate937(.a(gate272inter11), .b(gate272inter6), .O(gate272inter12));
  nand2 gate938(.a(gate272inter12), .b(gate272inter1), .O(G815));
nand2 gate273( .a(G642), .b(G794), .O(G818) );
nand2 gate274( .a(G770), .b(G794), .O(G819) );
nand2 gate275( .a(G645), .b(G797), .O(G820) );

  xor2  gate659(.a(G797), .b(G773), .O(gate276inter0));
  nand2 gate660(.a(gate276inter0), .b(s_16), .O(gate276inter1));
  and2  gate661(.a(G797), .b(G773), .O(gate276inter2));
  inv1  gate662(.a(s_16), .O(gate276inter3));
  inv1  gate663(.a(s_17), .O(gate276inter4));
  nand2 gate664(.a(gate276inter4), .b(gate276inter3), .O(gate276inter5));
  nor2  gate665(.a(gate276inter5), .b(gate276inter2), .O(gate276inter6));
  inv1  gate666(.a(G773), .O(gate276inter7));
  inv1  gate667(.a(G797), .O(gate276inter8));
  nand2 gate668(.a(gate276inter8), .b(gate276inter7), .O(gate276inter9));
  nand2 gate669(.a(s_17), .b(gate276inter3), .O(gate276inter10));
  nor2  gate670(.a(gate276inter10), .b(gate276inter9), .O(gate276inter11));
  nor2  gate671(.a(gate276inter11), .b(gate276inter6), .O(gate276inter12));
  nand2 gate672(.a(gate276inter12), .b(gate276inter1), .O(G821));

  xor2  gate1373(.a(G800), .b(G648), .O(gate277inter0));
  nand2 gate1374(.a(gate277inter0), .b(s_118), .O(gate277inter1));
  and2  gate1375(.a(G800), .b(G648), .O(gate277inter2));
  inv1  gate1376(.a(s_118), .O(gate277inter3));
  inv1  gate1377(.a(s_119), .O(gate277inter4));
  nand2 gate1378(.a(gate277inter4), .b(gate277inter3), .O(gate277inter5));
  nor2  gate1379(.a(gate277inter5), .b(gate277inter2), .O(gate277inter6));
  inv1  gate1380(.a(G648), .O(gate277inter7));
  inv1  gate1381(.a(G800), .O(gate277inter8));
  nand2 gate1382(.a(gate277inter8), .b(gate277inter7), .O(gate277inter9));
  nand2 gate1383(.a(s_119), .b(gate277inter3), .O(gate277inter10));
  nor2  gate1384(.a(gate277inter10), .b(gate277inter9), .O(gate277inter11));
  nor2  gate1385(.a(gate277inter11), .b(gate277inter6), .O(gate277inter12));
  nand2 gate1386(.a(gate277inter12), .b(gate277inter1), .O(G822));
nand2 gate278( .a(G776), .b(G800), .O(G823) );

  xor2  gate1583(.a(G803), .b(G651), .O(gate279inter0));
  nand2 gate1584(.a(gate279inter0), .b(s_148), .O(gate279inter1));
  and2  gate1585(.a(G803), .b(G651), .O(gate279inter2));
  inv1  gate1586(.a(s_148), .O(gate279inter3));
  inv1  gate1587(.a(s_149), .O(gate279inter4));
  nand2 gate1588(.a(gate279inter4), .b(gate279inter3), .O(gate279inter5));
  nor2  gate1589(.a(gate279inter5), .b(gate279inter2), .O(gate279inter6));
  inv1  gate1590(.a(G651), .O(gate279inter7));
  inv1  gate1591(.a(G803), .O(gate279inter8));
  nand2 gate1592(.a(gate279inter8), .b(gate279inter7), .O(gate279inter9));
  nand2 gate1593(.a(s_149), .b(gate279inter3), .O(gate279inter10));
  nor2  gate1594(.a(gate279inter10), .b(gate279inter9), .O(gate279inter11));
  nor2  gate1595(.a(gate279inter11), .b(gate279inter6), .O(gate279inter12));
  nand2 gate1596(.a(gate279inter12), .b(gate279inter1), .O(G824));
nand2 gate280( .a(G779), .b(G803), .O(G825) );
nand2 gate281( .a(G654), .b(G806), .O(G826) );
nand2 gate282( .a(G782), .b(G806), .O(G827) );
nand2 gate283( .a(G657), .b(G809), .O(G828) );
nand2 gate284( .a(G785), .b(G809), .O(G829) );
nand2 gate285( .a(G660), .b(G812), .O(G830) );
nand2 gate286( .a(G788), .b(G812), .O(G831) );
nand2 gate287( .a(G663), .b(G815), .O(G832) );
nand2 gate288( .a(G791), .b(G815), .O(G833) );
nand2 gate289( .a(G818), .b(G819), .O(G834) );
nand2 gate290( .a(G820), .b(G821), .O(G847) );
nand2 gate291( .a(G822), .b(G823), .O(G860) );
nand2 gate292( .a(G824), .b(G825), .O(G873) );
nand2 gate293( .a(G828), .b(G829), .O(G886) );
nand2 gate294( .a(G832), .b(G833), .O(G899) );
nand2 gate295( .a(G830), .b(G831), .O(G912) );
nand2 gate296( .a(G826), .b(G827), .O(G925) );
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );

  xor2  gate869(.a(G1036), .b(G1), .O(gate387inter0));
  nand2 gate870(.a(gate387inter0), .b(s_46), .O(gate387inter1));
  and2  gate871(.a(G1036), .b(G1), .O(gate387inter2));
  inv1  gate872(.a(s_46), .O(gate387inter3));
  inv1  gate873(.a(s_47), .O(gate387inter4));
  nand2 gate874(.a(gate387inter4), .b(gate387inter3), .O(gate387inter5));
  nor2  gate875(.a(gate387inter5), .b(gate387inter2), .O(gate387inter6));
  inv1  gate876(.a(G1), .O(gate387inter7));
  inv1  gate877(.a(G1036), .O(gate387inter8));
  nand2 gate878(.a(gate387inter8), .b(gate387inter7), .O(gate387inter9));
  nand2 gate879(.a(s_47), .b(gate387inter3), .O(gate387inter10));
  nor2  gate880(.a(gate387inter10), .b(gate387inter9), .O(gate387inter11));
  nor2  gate881(.a(gate387inter11), .b(gate387inter6), .O(gate387inter12));
  nand2 gate882(.a(gate387inter12), .b(gate387inter1), .O(G1132));

  xor2  gate1275(.a(G1039), .b(G2), .O(gate388inter0));
  nand2 gate1276(.a(gate388inter0), .b(s_104), .O(gate388inter1));
  and2  gate1277(.a(G1039), .b(G2), .O(gate388inter2));
  inv1  gate1278(.a(s_104), .O(gate388inter3));
  inv1  gate1279(.a(s_105), .O(gate388inter4));
  nand2 gate1280(.a(gate388inter4), .b(gate388inter3), .O(gate388inter5));
  nor2  gate1281(.a(gate388inter5), .b(gate388inter2), .O(gate388inter6));
  inv1  gate1282(.a(G2), .O(gate388inter7));
  inv1  gate1283(.a(G1039), .O(gate388inter8));
  nand2 gate1284(.a(gate388inter8), .b(gate388inter7), .O(gate388inter9));
  nand2 gate1285(.a(s_105), .b(gate388inter3), .O(gate388inter10));
  nor2  gate1286(.a(gate388inter10), .b(gate388inter9), .O(gate388inter11));
  nor2  gate1287(.a(gate388inter11), .b(gate388inter6), .O(gate388inter12));
  nand2 gate1288(.a(gate388inter12), .b(gate388inter1), .O(G1135));
nand2 gate389( .a(G3), .b(G1042), .O(G1138) );
nand2 gate390( .a(G4), .b(G1045), .O(G1141) );
nand2 gate391( .a(G5), .b(G1048), .O(G1144) );
nand2 gate392( .a(G6), .b(G1051), .O(G1147) );
nand2 gate393( .a(G7), .b(G1054), .O(G1150) );
nand2 gate394( .a(G8), .b(G1057), .O(G1153) );
nand2 gate395( .a(G9), .b(G1060), .O(G1156) );
nand2 gate396( .a(G10), .b(G1063), .O(G1159) );
nand2 gate397( .a(G11), .b(G1066), .O(G1162) );
nand2 gate398( .a(G12), .b(G1069), .O(G1165) );
nand2 gate399( .a(G13), .b(G1072), .O(G1168) );
nand2 gate400( .a(G14), .b(G1075), .O(G1171) );
nand2 gate401( .a(G15), .b(G1078), .O(G1174) );
nand2 gate402( .a(G16), .b(G1081), .O(G1177) );

  xor2  gate1597(.a(G1084), .b(G17), .O(gate403inter0));
  nand2 gate1598(.a(gate403inter0), .b(s_150), .O(gate403inter1));
  and2  gate1599(.a(G1084), .b(G17), .O(gate403inter2));
  inv1  gate1600(.a(s_150), .O(gate403inter3));
  inv1  gate1601(.a(s_151), .O(gate403inter4));
  nand2 gate1602(.a(gate403inter4), .b(gate403inter3), .O(gate403inter5));
  nor2  gate1603(.a(gate403inter5), .b(gate403inter2), .O(gate403inter6));
  inv1  gate1604(.a(G17), .O(gate403inter7));
  inv1  gate1605(.a(G1084), .O(gate403inter8));
  nand2 gate1606(.a(gate403inter8), .b(gate403inter7), .O(gate403inter9));
  nand2 gate1607(.a(s_151), .b(gate403inter3), .O(gate403inter10));
  nor2  gate1608(.a(gate403inter10), .b(gate403inter9), .O(gate403inter11));
  nor2  gate1609(.a(gate403inter11), .b(gate403inter6), .O(gate403inter12));
  nand2 gate1610(.a(gate403inter12), .b(gate403inter1), .O(G1180));
nand2 gate404( .a(G18), .b(G1087), .O(G1183) );
nand2 gate405( .a(G19), .b(G1090), .O(G1186) );
nand2 gate406( .a(G20), .b(G1093), .O(G1189) );

  xor2  gate575(.a(G1096), .b(G21), .O(gate407inter0));
  nand2 gate576(.a(gate407inter0), .b(s_4), .O(gate407inter1));
  and2  gate577(.a(G1096), .b(G21), .O(gate407inter2));
  inv1  gate578(.a(s_4), .O(gate407inter3));
  inv1  gate579(.a(s_5), .O(gate407inter4));
  nand2 gate580(.a(gate407inter4), .b(gate407inter3), .O(gate407inter5));
  nor2  gate581(.a(gate407inter5), .b(gate407inter2), .O(gate407inter6));
  inv1  gate582(.a(G21), .O(gate407inter7));
  inv1  gate583(.a(G1096), .O(gate407inter8));
  nand2 gate584(.a(gate407inter8), .b(gate407inter7), .O(gate407inter9));
  nand2 gate585(.a(s_5), .b(gate407inter3), .O(gate407inter10));
  nor2  gate586(.a(gate407inter10), .b(gate407inter9), .O(gate407inter11));
  nor2  gate587(.a(gate407inter11), .b(gate407inter6), .O(gate407inter12));
  nand2 gate588(.a(gate407inter12), .b(gate407inter1), .O(G1192));
nand2 gate408( .a(G22), .b(G1099), .O(G1195) );
nand2 gate409( .a(G23), .b(G1102), .O(G1198) );
nand2 gate410( .a(G24), .b(G1105), .O(G1201) );
nand2 gate411( .a(G25), .b(G1108), .O(G1204) );
nand2 gate412( .a(G26), .b(G1111), .O(G1207) );
nand2 gate413( .a(G27), .b(G1114), .O(G1210) );
nand2 gate414( .a(G28), .b(G1117), .O(G1213) );

  xor2  gate939(.a(G1120), .b(G29), .O(gate415inter0));
  nand2 gate940(.a(gate415inter0), .b(s_56), .O(gate415inter1));
  and2  gate941(.a(G1120), .b(G29), .O(gate415inter2));
  inv1  gate942(.a(s_56), .O(gate415inter3));
  inv1  gate943(.a(s_57), .O(gate415inter4));
  nand2 gate944(.a(gate415inter4), .b(gate415inter3), .O(gate415inter5));
  nor2  gate945(.a(gate415inter5), .b(gate415inter2), .O(gate415inter6));
  inv1  gate946(.a(G29), .O(gate415inter7));
  inv1  gate947(.a(G1120), .O(gate415inter8));
  nand2 gate948(.a(gate415inter8), .b(gate415inter7), .O(gate415inter9));
  nand2 gate949(.a(s_57), .b(gate415inter3), .O(gate415inter10));
  nor2  gate950(.a(gate415inter10), .b(gate415inter9), .O(gate415inter11));
  nor2  gate951(.a(gate415inter11), .b(gate415inter6), .O(gate415inter12));
  nand2 gate952(.a(gate415inter12), .b(gate415inter1), .O(G1216));

  xor2  gate1163(.a(G1123), .b(G30), .O(gate416inter0));
  nand2 gate1164(.a(gate416inter0), .b(s_88), .O(gate416inter1));
  and2  gate1165(.a(G1123), .b(G30), .O(gate416inter2));
  inv1  gate1166(.a(s_88), .O(gate416inter3));
  inv1  gate1167(.a(s_89), .O(gate416inter4));
  nand2 gate1168(.a(gate416inter4), .b(gate416inter3), .O(gate416inter5));
  nor2  gate1169(.a(gate416inter5), .b(gate416inter2), .O(gate416inter6));
  inv1  gate1170(.a(G30), .O(gate416inter7));
  inv1  gate1171(.a(G1123), .O(gate416inter8));
  nand2 gate1172(.a(gate416inter8), .b(gate416inter7), .O(gate416inter9));
  nand2 gate1173(.a(s_89), .b(gate416inter3), .O(gate416inter10));
  nor2  gate1174(.a(gate416inter10), .b(gate416inter9), .O(gate416inter11));
  nor2  gate1175(.a(gate416inter11), .b(gate416inter6), .O(gate416inter12));
  nand2 gate1176(.a(gate416inter12), .b(gate416inter1), .O(G1219));
nand2 gate417( .a(G31), .b(G1126), .O(G1222) );
nand2 gate418( .a(G32), .b(G1129), .O(G1225) );
nand2 gate419( .a(G1), .b(G1132), .O(G1228) );
nand2 gate420( .a(G1036), .b(G1132), .O(G1229) );
nand2 gate421( .a(G2), .b(G1135), .O(G1230) );
nand2 gate422( .a(G1039), .b(G1135), .O(G1231) );
nand2 gate423( .a(G3), .b(G1138), .O(G1232) );
nand2 gate424( .a(G1042), .b(G1138), .O(G1233) );
nand2 gate425( .a(G4), .b(G1141), .O(G1234) );
nand2 gate426( .a(G1045), .b(G1141), .O(G1235) );

  xor2  gate1485(.a(G1144), .b(G5), .O(gate427inter0));
  nand2 gate1486(.a(gate427inter0), .b(s_134), .O(gate427inter1));
  and2  gate1487(.a(G1144), .b(G5), .O(gate427inter2));
  inv1  gate1488(.a(s_134), .O(gate427inter3));
  inv1  gate1489(.a(s_135), .O(gate427inter4));
  nand2 gate1490(.a(gate427inter4), .b(gate427inter3), .O(gate427inter5));
  nor2  gate1491(.a(gate427inter5), .b(gate427inter2), .O(gate427inter6));
  inv1  gate1492(.a(G5), .O(gate427inter7));
  inv1  gate1493(.a(G1144), .O(gate427inter8));
  nand2 gate1494(.a(gate427inter8), .b(gate427inter7), .O(gate427inter9));
  nand2 gate1495(.a(s_135), .b(gate427inter3), .O(gate427inter10));
  nor2  gate1496(.a(gate427inter10), .b(gate427inter9), .O(gate427inter11));
  nor2  gate1497(.a(gate427inter11), .b(gate427inter6), .O(gate427inter12));
  nand2 gate1498(.a(gate427inter12), .b(gate427inter1), .O(G1236));

  xor2  gate771(.a(G1144), .b(G1048), .O(gate428inter0));
  nand2 gate772(.a(gate428inter0), .b(s_32), .O(gate428inter1));
  and2  gate773(.a(G1144), .b(G1048), .O(gate428inter2));
  inv1  gate774(.a(s_32), .O(gate428inter3));
  inv1  gate775(.a(s_33), .O(gate428inter4));
  nand2 gate776(.a(gate428inter4), .b(gate428inter3), .O(gate428inter5));
  nor2  gate777(.a(gate428inter5), .b(gate428inter2), .O(gate428inter6));
  inv1  gate778(.a(G1048), .O(gate428inter7));
  inv1  gate779(.a(G1144), .O(gate428inter8));
  nand2 gate780(.a(gate428inter8), .b(gate428inter7), .O(gate428inter9));
  nand2 gate781(.a(s_33), .b(gate428inter3), .O(gate428inter10));
  nor2  gate782(.a(gate428inter10), .b(gate428inter9), .O(gate428inter11));
  nor2  gate783(.a(gate428inter11), .b(gate428inter6), .O(gate428inter12));
  nand2 gate784(.a(gate428inter12), .b(gate428inter1), .O(G1237));
nand2 gate429( .a(G6), .b(G1147), .O(G1238) );
nand2 gate430( .a(G1051), .b(G1147), .O(G1239) );

  xor2  gate1499(.a(G1150), .b(G7), .O(gate431inter0));
  nand2 gate1500(.a(gate431inter0), .b(s_136), .O(gate431inter1));
  and2  gate1501(.a(G1150), .b(G7), .O(gate431inter2));
  inv1  gate1502(.a(s_136), .O(gate431inter3));
  inv1  gate1503(.a(s_137), .O(gate431inter4));
  nand2 gate1504(.a(gate431inter4), .b(gate431inter3), .O(gate431inter5));
  nor2  gate1505(.a(gate431inter5), .b(gate431inter2), .O(gate431inter6));
  inv1  gate1506(.a(G7), .O(gate431inter7));
  inv1  gate1507(.a(G1150), .O(gate431inter8));
  nand2 gate1508(.a(gate431inter8), .b(gate431inter7), .O(gate431inter9));
  nand2 gate1509(.a(s_137), .b(gate431inter3), .O(gate431inter10));
  nor2  gate1510(.a(gate431inter10), .b(gate431inter9), .O(gate431inter11));
  nor2  gate1511(.a(gate431inter11), .b(gate431inter6), .O(gate431inter12));
  nand2 gate1512(.a(gate431inter12), .b(gate431inter1), .O(G1240));

  xor2  gate883(.a(G1150), .b(G1054), .O(gate432inter0));
  nand2 gate884(.a(gate432inter0), .b(s_48), .O(gate432inter1));
  and2  gate885(.a(G1150), .b(G1054), .O(gate432inter2));
  inv1  gate886(.a(s_48), .O(gate432inter3));
  inv1  gate887(.a(s_49), .O(gate432inter4));
  nand2 gate888(.a(gate432inter4), .b(gate432inter3), .O(gate432inter5));
  nor2  gate889(.a(gate432inter5), .b(gate432inter2), .O(gate432inter6));
  inv1  gate890(.a(G1054), .O(gate432inter7));
  inv1  gate891(.a(G1150), .O(gate432inter8));
  nand2 gate892(.a(gate432inter8), .b(gate432inter7), .O(gate432inter9));
  nand2 gate893(.a(s_49), .b(gate432inter3), .O(gate432inter10));
  nor2  gate894(.a(gate432inter10), .b(gate432inter9), .O(gate432inter11));
  nor2  gate895(.a(gate432inter11), .b(gate432inter6), .O(gate432inter12));
  nand2 gate896(.a(gate432inter12), .b(gate432inter1), .O(G1241));

  xor2  gate995(.a(G1153), .b(G8), .O(gate433inter0));
  nand2 gate996(.a(gate433inter0), .b(s_64), .O(gate433inter1));
  and2  gate997(.a(G1153), .b(G8), .O(gate433inter2));
  inv1  gate998(.a(s_64), .O(gate433inter3));
  inv1  gate999(.a(s_65), .O(gate433inter4));
  nand2 gate1000(.a(gate433inter4), .b(gate433inter3), .O(gate433inter5));
  nor2  gate1001(.a(gate433inter5), .b(gate433inter2), .O(gate433inter6));
  inv1  gate1002(.a(G8), .O(gate433inter7));
  inv1  gate1003(.a(G1153), .O(gate433inter8));
  nand2 gate1004(.a(gate433inter8), .b(gate433inter7), .O(gate433inter9));
  nand2 gate1005(.a(s_65), .b(gate433inter3), .O(gate433inter10));
  nor2  gate1006(.a(gate433inter10), .b(gate433inter9), .O(gate433inter11));
  nor2  gate1007(.a(gate433inter11), .b(gate433inter6), .O(gate433inter12));
  nand2 gate1008(.a(gate433inter12), .b(gate433inter1), .O(G1242));
nand2 gate434( .a(G1057), .b(G1153), .O(G1243) );

  xor2  gate1009(.a(G1156), .b(G9), .O(gate435inter0));
  nand2 gate1010(.a(gate435inter0), .b(s_66), .O(gate435inter1));
  and2  gate1011(.a(G1156), .b(G9), .O(gate435inter2));
  inv1  gate1012(.a(s_66), .O(gate435inter3));
  inv1  gate1013(.a(s_67), .O(gate435inter4));
  nand2 gate1014(.a(gate435inter4), .b(gate435inter3), .O(gate435inter5));
  nor2  gate1015(.a(gate435inter5), .b(gate435inter2), .O(gate435inter6));
  inv1  gate1016(.a(G9), .O(gate435inter7));
  inv1  gate1017(.a(G1156), .O(gate435inter8));
  nand2 gate1018(.a(gate435inter8), .b(gate435inter7), .O(gate435inter9));
  nand2 gate1019(.a(s_67), .b(gate435inter3), .O(gate435inter10));
  nor2  gate1020(.a(gate435inter10), .b(gate435inter9), .O(gate435inter11));
  nor2  gate1021(.a(gate435inter11), .b(gate435inter6), .O(gate435inter12));
  nand2 gate1022(.a(gate435inter12), .b(gate435inter1), .O(G1244));

  xor2  gate799(.a(G1156), .b(G1060), .O(gate436inter0));
  nand2 gate800(.a(gate436inter0), .b(s_36), .O(gate436inter1));
  and2  gate801(.a(G1156), .b(G1060), .O(gate436inter2));
  inv1  gate802(.a(s_36), .O(gate436inter3));
  inv1  gate803(.a(s_37), .O(gate436inter4));
  nand2 gate804(.a(gate436inter4), .b(gate436inter3), .O(gate436inter5));
  nor2  gate805(.a(gate436inter5), .b(gate436inter2), .O(gate436inter6));
  inv1  gate806(.a(G1060), .O(gate436inter7));
  inv1  gate807(.a(G1156), .O(gate436inter8));
  nand2 gate808(.a(gate436inter8), .b(gate436inter7), .O(gate436inter9));
  nand2 gate809(.a(s_37), .b(gate436inter3), .O(gate436inter10));
  nor2  gate810(.a(gate436inter10), .b(gate436inter9), .O(gate436inter11));
  nor2  gate811(.a(gate436inter11), .b(gate436inter6), .O(gate436inter12));
  nand2 gate812(.a(gate436inter12), .b(gate436inter1), .O(G1245));
nand2 gate437( .a(G10), .b(G1159), .O(G1246) );
nand2 gate438( .a(G1063), .b(G1159), .O(G1247) );
nand2 gate439( .a(G11), .b(G1162), .O(G1248) );
nand2 gate440( .a(G1066), .b(G1162), .O(G1249) );
nand2 gate441( .a(G12), .b(G1165), .O(G1250) );
nand2 gate442( .a(G1069), .b(G1165), .O(G1251) );
nand2 gate443( .a(G13), .b(G1168), .O(G1252) );

  xor2  gate1065(.a(G1168), .b(G1072), .O(gate444inter0));
  nand2 gate1066(.a(gate444inter0), .b(s_74), .O(gate444inter1));
  and2  gate1067(.a(G1168), .b(G1072), .O(gate444inter2));
  inv1  gate1068(.a(s_74), .O(gate444inter3));
  inv1  gate1069(.a(s_75), .O(gate444inter4));
  nand2 gate1070(.a(gate444inter4), .b(gate444inter3), .O(gate444inter5));
  nor2  gate1071(.a(gate444inter5), .b(gate444inter2), .O(gate444inter6));
  inv1  gate1072(.a(G1072), .O(gate444inter7));
  inv1  gate1073(.a(G1168), .O(gate444inter8));
  nand2 gate1074(.a(gate444inter8), .b(gate444inter7), .O(gate444inter9));
  nand2 gate1075(.a(s_75), .b(gate444inter3), .O(gate444inter10));
  nor2  gate1076(.a(gate444inter10), .b(gate444inter9), .O(gate444inter11));
  nor2  gate1077(.a(gate444inter11), .b(gate444inter6), .O(gate444inter12));
  nand2 gate1078(.a(gate444inter12), .b(gate444inter1), .O(G1253));
nand2 gate445( .a(G14), .b(G1171), .O(G1254) );
nand2 gate446( .a(G1075), .b(G1171), .O(G1255) );
nand2 gate447( .a(G15), .b(G1174), .O(G1256) );
nand2 gate448( .a(G1078), .b(G1174), .O(G1257) );
nand2 gate449( .a(G16), .b(G1177), .O(G1258) );
nand2 gate450( .a(G1081), .b(G1177), .O(G1259) );
nand2 gate451( .a(G17), .b(G1180), .O(G1260) );
nand2 gate452( .a(G1084), .b(G1180), .O(G1261) );
nand2 gate453( .a(G18), .b(G1183), .O(G1262) );
nand2 gate454( .a(G1087), .b(G1183), .O(G1263) );
nand2 gate455( .a(G19), .b(G1186), .O(G1264) );
nand2 gate456( .a(G1090), .b(G1186), .O(G1265) );
nand2 gate457( .a(G20), .b(G1189), .O(G1266) );
nand2 gate458( .a(G1093), .b(G1189), .O(G1267) );
nand2 gate459( .a(G21), .b(G1192), .O(G1268) );
nand2 gate460( .a(G1096), .b(G1192), .O(G1269) );
nand2 gate461( .a(G22), .b(G1195), .O(G1270) );

  xor2  gate589(.a(G1195), .b(G1099), .O(gate462inter0));
  nand2 gate590(.a(gate462inter0), .b(s_6), .O(gate462inter1));
  and2  gate591(.a(G1195), .b(G1099), .O(gate462inter2));
  inv1  gate592(.a(s_6), .O(gate462inter3));
  inv1  gate593(.a(s_7), .O(gate462inter4));
  nand2 gate594(.a(gate462inter4), .b(gate462inter3), .O(gate462inter5));
  nor2  gate595(.a(gate462inter5), .b(gate462inter2), .O(gate462inter6));
  inv1  gate596(.a(G1099), .O(gate462inter7));
  inv1  gate597(.a(G1195), .O(gate462inter8));
  nand2 gate598(.a(gate462inter8), .b(gate462inter7), .O(gate462inter9));
  nand2 gate599(.a(s_7), .b(gate462inter3), .O(gate462inter10));
  nor2  gate600(.a(gate462inter10), .b(gate462inter9), .O(gate462inter11));
  nor2  gate601(.a(gate462inter11), .b(gate462inter6), .O(gate462inter12));
  nand2 gate602(.a(gate462inter12), .b(gate462inter1), .O(G1271));
nand2 gate463( .a(G23), .b(G1198), .O(G1272) );
nand2 gate464( .a(G1102), .b(G1198), .O(G1273) );
nand2 gate465( .a(G24), .b(G1201), .O(G1274) );
nand2 gate466( .a(G1105), .b(G1201), .O(G1275) );

  xor2  gate813(.a(G1204), .b(G25), .O(gate467inter0));
  nand2 gate814(.a(gate467inter0), .b(s_38), .O(gate467inter1));
  and2  gate815(.a(G1204), .b(G25), .O(gate467inter2));
  inv1  gate816(.a(s_38), .O(gate467inter3));
  inv1  gate817(.a(s_39), .O(gate467inter4));
  nand2 gate818(.a(gate467inter4), .b(gate467inter3), .O(gate467inter5));
  nor2  gate819(.a(gate467inter5), .b(gate467inter2), .O(gate467inter6));
  inv1  gate820(.a(G25), .O(gate467inter7));
  inv1  gate821(.a(G1204), .O(gate467inter8));
  nand2 gate822(.a(gate467inter8), .b(gate467inter7), .O(gate467inter9));
  nand2 gate823(.a(s_39), .b(gate467inter3), .O(gate467inter10));
  nor2  gate824(.a(gate467inter10), .b(gate467inter9), .O(gate467inter11));
  nor2  gate825(.a(gate467inter11), .b(gate467inter6), .O(gate467inter12));
  nand2 gate826(.a(gate467inter12), .b(gate467inter1), .O(G1276));

  xor2  gate1317(.a(G1204), .b(G1108), .O(gate468inter0));
  nand2 gate1318(.a(gate468inter0), .b(s_110), .O(gate468inter1));
  and2  gate1319(.a(G1204), .b(G1108), .O(gate468inter2));
  inv1  gate1320(.a(s_110), .O(gate468inter3));
  inv1  gate1321(.a(s_111), .O(gate468inter4));
  nand2 gate1322(.a(gate468inter4), .b(gate468inter3), .O(gate468inter5));
  nor2  gate1323(.a(gate468inter5), .b(gate468inter2), .O(gate468inter6));
  inv1  gate1324(.a(G1108), .O(gate468inter7));
  inv1  gate1325(.a(G1204), .O(gate468inter8));
  nand2 gate1326(.a(gate468inter8), .b(gate468inter7), .O(gate468inter9));
  nand2 gate1327(.a(s_111), .b(gate468inter3), .O(gate468inter10));
  nor2  gate1328(.a(gate468inter10), .b(gate468inter9), .O(gate468inter11));
  nor2  gate1329(.a(gate468inter11), .b(gate468inter6), .O(gate468inter12));
  nand2 gate1330(.a(gate468inter12), .b(gate468inter1), .O(G1277));
nand2 gate469( .a(G26), .b(G1207), .O(G1278) );
nand2 gate470( .a(G1111), .b(G1207), .O(G1279) );

  xor2  gate743(.a(G1210), .b(G27), .O(gate471inter0));
  nand2 gate744(.a(gate471inter0), .b(s_28), .O(gate471inter1));
  and2  gate745(.a(G1210), .b(G27), .O(gate471inter2));
  inv1  gate746(.a(s_28), .O(gate471inter3));
  inv1  gate747(.a(s_29), .O(gate471inter4));
  nand2 gate748(.a(gate471inter4), .b(gate471inter3), .O(gate471inter5));
  nor2  gate749(.a(gate471inter5), .b(gate471inter2), .O(gate471inter6));
  inv1  gate750(.a(G27), .O(gate471inter7));
  inv1  gate751(.a(G1210), .O(gate471inter8));
  nand2 gate752(.a(gate471inter8), .b(gate471inter7), .O(gate471inter9));
  nand2 gate753(.a(s_29), .b(gate471inter3), .O(gate471inter10));
  nor2  gate754(.a(gate471inter10), .b(gate471inter9), .O(gate471inter11));
  nor2  gate755(.a(gate471inter11), .b(gate471inter6), .O(gate471inter12));
  nand2 gate756(.a(gate471inter12), .b(gate471inter1), .O(G1280));
nand2 gate472( .a(G1114), .b(G1210), .O(G1281) );
nand2 gate473( .a(G28), .b(G1213), .O(G1282) );
nand2 gate474( .a(G1117), .b(G1213), .O(G1283) );
nand2 gate475( .a(G29), .b(G1216), .O(G1284) );
nand2 gate476( .a(G1120), .b(G1216), .O(G1285) );
nand2 gate477( .a(G30), .b(G1219), .O(G1286) );
nand2 gate478( .a(G1123), .b(G1219), .O(G1287) );
nand2 gate479( .a(G31), .b(G1222), .O(G1288) );
nand2 gate480( .a(G1126), .b(G1222), .O(G1289) );
nand2 gate481( .a(G32), .b(G1225), .O(G1290) );

  xor2  gate1541(.a(G1225), .b(G1129), .O(gate482inter0));
  nand2 gate1542(.a(gate482inter0), .b(s_142), .O(gate482inter1));
  and2  gate1543(.a(G1225), .b(G1129), .O(gate482inter2));
  inv1  gate1544(.a(s_142), .O(gate482inter3));
  inv1  gate1545(.a(s_143), .O(gate482inter4));
  nand2 gate1546(.a(gate482inter4), .b(gate482inter3), .O(gate482inter5));
  nor2  gate1547(.a(gate482inter5), .b(gate482inter2), .O(gate482inter6));
  inv1  gate1548(.a(G1129), .O(gate482inter7));
  inv1  gate1549(.a(G1225), .O(gate482inter8));
  nand2 gate1550(.a(gate482inter8), .b(gate482inter7), .O(gate482inter9));
  nand2 gate1551(.a(s_143), .b(gate482inter3), .O(gate482inter10));
  nor2  gate1552(.a(gate482inter10), .b(gate482inter9), .O(gate482inter11));
  nor2  gate1553(.a(gate482inter11), .b(gate482inter6), .O(gate482inter12));
  nand2 gate1554(.a(gate482inter12), .b(gate482inter1), .O(G1291));
nand2 gate483( .a(G1228), .b(G1229), .O(G1292) );
nand2 gate484( .a(G1230), .b(G1231), .O(G1293) );
nand2 gate485( .a(G1232), .b(G1233), .O(G1294) );
nand2 gate486( .a(G1234), .b(G1235), .O(G1295) );
nand2 gate487( .a(G1236), .b(G1237), .O(G1296) );
nand2 gate488( .a(G1238), .b(G1239), .O(G1297) );
nand2 gate489( .a(G1240), .b(G1241), .O(G1298) );
nand2 gate490( .a(G1242), .b(G1243), .O(G1299) );

  xor2  gate967(.a(G1245), .b(G1244), .O(gate491inter0));
  nand2 gate968(.a(gate491inter0), .b(s_60), .O(gate491inter1));
  and2  gate969(.a(G1245), .b(G1244), .O(gate491inter2));
  inv1  gate970(.a(s_60), .O(gate491inter3));
  inv1  gate971(.a(s_61), .O(gate491inter4));
  nand2 gate972(.a(gate491inter4), .b(gate491inter3), .O(gate491inter5));
  nor2  gate973(.a(gate491inter5), .b(gate491inter2), .O(gate491inter6));
  inv1  gate974(.a(G1244), .O(gate491inter7));
  inv1  gate975(.a(G1245), .O(gate491inter8));
  nand2 gate976(.a(gate491inter8), .b(gate491inter7), .O(gate491inter9));
  nand2 gate977(.a(s_61), .b(gate491inter3), .O(gate491inter10));
  nor2  gate978(.a(gate491inter10), .b(gate491inter9), .O(gate491inter11));
  nor2  gate979(.a(gate491inter11), .b(gate491inter6), .O(gate491inter12));
  nand2 gate980(.a(gate491inter12), .b(gate491inter1), .O(G1300));
nand2 gate492( .a(G1246), .b(G1247), .O(G1301) );
nand2 gate493( .a(G1248), .b(G1249), .O(G1302) );
nand2 gate494( .a(G1250), .b(G1251), .O(G1303) );
nand2 gate495( .a(G1252), .b(G1253), .O(G1304) );
nand2 gate496( .a(G1254), .b(G1255), .O(G1305) );

  xor2  gate1177(.a(G1257), .b(G1256), .O(gate497inter0));
  nand2 gate1178(.a(gate497inter0), .b(s_90), .O(gate497inter1));
  and2  gate1179(.a(G1257), .b(G1256), .O(gate497inter2));
  inv1  gate1180(.a(s_90), .O(gate497inter3));
  inv1  gate1181(.a(s_91), .O(gate497inter4));
  nand2 gate1182(.a(gate497inter4), .b(gate497inter3), .O(gate497inter5));
  nor2  gate1183(.a(gate497inter5), .b(gate497inter2), .O(gate497inter6));
  inv1  gate1184(.a(G1256), .O(gate497inter7));
  inv1  gate1185(.a(G1257), .O(gate497inter8));
  nand2 gate1186(.a(gate497inter8), .b(gate497inter7), .O(gate497inter9));
  nand2 gate1187(.a(s_91), .b(gate497inter3), .O(gate497inter10));
  nor2  gate1188(.a(gate497inter10), .b(gate497inter9), .O(gate497inter11));
  nor2  gate1189(.a(gate497inter11), .b(gate497inter6), .O(gate497inter12));
  nand2 gate1190(.a(gate497inter12), .b(gate497inter1), .O(G1306));
nand2 gate498( .a(G1258), .b(G1259), .O(G1307) );
nand2 gate499( .a(G1260), .b(G1261), .O(G1308) );
nand2 gate500( .a(G1262), .b(G1263), .O(G1309) );
nand2 gate501( .a(G1264), .b(G1265), .O(G1310) );
nand2 gate502( .a(G1266), .b(G1267), .O(G1311) );
nand2 gate503( .a(G1268), .b(G1269), .O(G1312) );
nand2 gate504( .a(G1270), .b(G1271), .O(G1313) );
nand2 gate505( .a(G1272), .b(G1273), .O(G1314) );
nand2 gate506( .a(G1274), .b(G1275), .O(G1315) );
nand2 gate507( .a(G1276), .b(G1277), .O(G1316) );
nand2 gate508( .a(G1278), .b(G1279), .O(G1317) );
nand2 gate509( .a(G1280), .b(G1281), .O(G1318) );
nand2 gate510( .a(G1282), .b(G1283), .O(G1319) );
nand2 gate511( .a(G1284), .b(G1285), .O(G1320) );
nand2 gate512( .a(G1286), .b(G1287), .O(G1321) );
nand2 gate513( .a(G1288), .b(G1289), .O(G1322) );
nand2 gate514( .a(G1290), .b(G1291), .O(G1323) );
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule