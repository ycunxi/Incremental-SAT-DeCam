module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);

input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;//RE__PI;

input s_0,s_1;//RE__ALLOW(00,01,10,11);
input s_2,s_3;//RE__ALLOW(00,01,10,11);
input s_4,s_5;//RE__ALLOW(00,01,10,11);
input s_6,s_7;//RE__ALLOW(00,01,10,11);
input s_8,s_9;//RE__ALLOW(00,01,10,11);
input s_10,s_11;//RE__ALLOW(00,01,10,11);
input s_12,s_13;//RE__ALLOW(00,01,10,11);
input s_14,s_15;//RE__ALLOW(00,01,10,11);
input s_16,s_17;//RE__ALLOW(00,01,10,11);
input s_18,s_19;//RE__ALLOW(00,01,10,11);
input s_20,s_21;//RE__ALLOW(00,01,10,11);
input s_22,s_23;//RE__ALLOW(00,01,10,11);
input s_24,s_25;//RE__ALLOW(00,01,10,11);
input s_26,s_27;//RE__ALLOW(00,01,10,11);
input s_28,s_29;//RE__ALLOW(00,01,10,11);
input s_30,s_31;//RE__ALLOW(00,01,10,11);
input s_32,s_33;//RE__ALLOW(00,01,10,11);
input s_34,s_35;//RE__ALLOW(00,01,10,11);
input s_36,s_37;//RE__ALLOW(00,01,10,11);
input s_38,s_39;//RE__ALLOW(00,01,10,11);
input s_40,s_41;//RE__ALLOW(00,01,10,11);
input s_42,s_43;//RE__ALLOW(00,01,10,11);
input s_44,s_45;//RE__ALLOW(00,01,10,11);
input s_46,s_47;//RE__ALLOW(00,01,10,11);
input s_48,s_49;//RE__ALLOW(00,01,10,11);
input s_50,s_51;//RE__ALLOW(00,01,10,11);
input s_52,s_53;//RE__ALLOW(00,01,10,11);
input s_54,s_55;//RE__ALLOW(00,01,10,11);
input s_56,s_57;//RE__ALLOW(00,01,10,11);
input s_58,s_59;//RE__ALLOW(00,01,10,11);
input s_60,s_61;//RE__ALLOW(00,01,10,11);
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;

  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate275inter0, gate275inter1, gate275inter2, gate275inter3, gate275inter4, gate275inter5, gate275inter6, gate275inter7, gate275inter8, gate275inter9, gate275inter10, gate275inter11, gate275inter12, gate153inter0, gate153inter1, gate153inter2, gate153inter3, gate153inter4, gate153inter5, gate153inter6, gate153inter7, gate153inter8, gate153inter9, gate153inter10, gate153inter11, gate153inter12, gate112inter0, gate112inter1, gate112inter2, gate112inter3, gate112inter4, gate112inter5, gate112inter6, gate112inter7, gate112inter8, gate112inter9, gate112inter10, gate112inter11, gate112inter12, gate254inter0, gate254inter1, gate254inter2, gate254inter3, gate254inter4, gate254inter5, gate254inter6, gate254inter7, gate254inter8, gate254inter9, gate254inter10, gate254inter11, gate254inter12, gate183inter0, gate183inter1, gate183inter2, gate183inter3, gate183inter4, gate183inter5, gate183inter6, gate183inter7, gate183inter8, gate183inter9, gate183inter10, gate183inter11, gate183inter12, gate221inter0, gate221inter1, gate221inter2, gate221inter3, gate221inter4, gate221inter5, gate221inter6, gate221inter7, gate221inter8, gate221inter9, gate221inter10, gate221inter11, gate221inter12, gate390inter0, gate390inter1, gate390inter2, gate390inter3, gate390inter4, gate390inter5, gate390inter6, gate390inter7, gate390inter8, gate390inter9, gate390inter10, gate390inter11, gate390inter12, gate234inter0, gate234inter1, gate234inter2, gate234inter3, gate234inter4, gate234inter5, gate234inter6, gate234inter7, gate234inter8, gate234inter9, gate234inter10, gate234inter11, gate234inter12, gate276inter0, gate276inter1, gate276inter2, gate276inter3, gate276inter4, gate276inter5, gate276inter6, gate276inter7, gate276inter8, gate276inter9, gate276inter10, gate276inter11, gate276inter12, gate106inter0, gate106inter1, gate106inter2, gate106inter3, gate106inter4, gate106inter5, gate106inter6, gate106inter7, gate106inter8, gate106inter9, gate106inter10, gate106inter11, gate106inter12, gate483inter0, gate483inter1, gate483inter2, gate483inter3, gate483inter4, gate483inter5, gate483inter6, gate483inter7, gate483inter8, gate483inter9, gate483inter10, gate483inter11, gate483inter12, gate43inter0, gate43inter1, gate43inter2, gate43inter3, gate43inter4, gate43inter5, gate43inter6, gate43inter7, gate43inter8, gate43inter9, gate43inter10, gate43inter11, gate43inter12, gate28inter0, gate28inter1, gate28inter2, gate28inter3, gate28inter4, gate28inter5, gate28inter6, gate28inter7, gate28inter8, gate28inter9, gate28inter10, gate28inter11, gate28inter12, gate44inter0, gate44inter1, gate44inter2, gate44inter3, gate44inter4, gate44inter5, gate44inter6, gate44inter7, gate44inter8, gate44inter9, gate44inter10, gate44inter11, gate44inter12, gate115inter0, gate115inter1, gate115inter2, gate115inter3, gate115inter4, gate115inter5, gate115inter6, gate115inter7, gate115inter8, gate115inter9, gate115inter10, gate115inter11, gate115inter12, gate397inter0, gate397inter1, gate397inter2, gate397inter3, gate397inter4, gate397inter5, gate397inter6, gate397inter7, gate397inter8, gate397inter9, gate397inter10, gate397inter11, gate397inter12, gate124inter0, gate124inter1, gate124inter2, gate124inter3, gate124inter4, gate124inter5, gate124inter6, gate124inter7, gate124inter8, gate124inter9, gate124inter10, gate124inter11, gate124inter12, gate468inter0, gate468inter1, gate468inter2, gate468inter3, gate468inter4, gate468inter5, gate468inter6, gate468inter7, gate468inter8, gate468inter9, gate468inter10, gate468inter11, gate468inter12, gate161inter0, gate161inter1, gate161inter2, gate161inter3, gate161inter4, gate161inter5, gate161inter6, gate161inter7, gate161inter8, gate161inter9, gate161inter10, gate161inter11, gate161inter12, gate431inter0, gate431inter1, gate431inter2, gate431inter3, gate431inter4, gate431inter5, gate431inter6, gate431inter7, gate431inter8, gate431inter9, gate431inter10, gate431inter11, gate431inter12, gate496inter0, gate496inter1, gate496inter2, gate496inter3, gate496inter4, gate496inter5, gate496inter6, gate496inter7, gate496inter8, gate496inter9, gate496inter10, gate496inter11, gate496inter12, gate205inter0, gate205inter1, gate205inter2, gate205inter3, gate205inter4, gate205inter5, gate205inter6, gate205inter7, gate205inter8, gate205inter9, gate205inter10, gate205inter11, gate205inter12, gate31inter0, gate31inter1, gate31inter2, gate31inter3, gate31inter4, gate31inter5, gate31inter6, gate31inter7, gate31inter8, gate31inter9, gate31inter10, gate31inter11, gate31inter12, gate186inter0, gate186inter1, gate186inter2, gate186inter3, gate186inter4, gate186inter5, gate186inter6, gate186inter7, gate186inter8, gate186inter9, gate186inter10, gate186inter11, gate186inter12, gate238inter0, gate238inter1, gate238inter2, gate238inter3, gate238inter4, gate238inter5, gate238inter6, gate238inter7, gate238inter8, gate238inter9, gate238inter10, gate238inter11, gate238inter12, gate295inter0, gate295inter1, gate295inter2, gate295inter3, gate295inter4, gate295inter5, gate295inter6, gate295inter7, gate295inter8, gate295inter9, gate295inter10, gate295inter11, gate295inter12, gate190inter0, gate190inter1, gate190inter2, gate190inter3, gate190inter4, gate190inter5, gate190inter6, gate190inter7, gate190inter8, gate190inter9, gate190inter10, gate190inter11, gate190inter12, gate457inter0, gate457inter1, gate457inter2, gate457inter3, gate457inter4, gate457inter5, gate457inter6, gate457inter7, gate457inter8, gate457inter9, gate457inter10, gate457inter11, gate457inter12, gate179inter0, gate179inter1, gate179inter2, gate179inter3, gate179inter4, gate179inter5, gate179inter6, gate179inter7, gate179inter8, gate179inter9, gate179inter10, gate179inter11, gate179inter12, gate480inter0, gate480inter1, gate480inter2, gate480inter3, gate480inter4, gate480inter5, gate480inter6, gate480inter7, gate480inter8, gate480inter9, gate480inter10, gate480inter11, gate480inter12, gate281inter0, gate281inter1, gate281inter2, gate281inter3, gate281inter4, gate281inter5, gate281inter6, gate281inter7, gate281inter8, gate281inter9, gate281inter10, gate281inter11, gate281inter12;



and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );
nand2 gate9( .a(G1), .b(G2), .O(G266) );
nand2 gate10( .a(G3), .b(G4), .O(G269) );
nand2 gate11( .a(G5), .b(G6), .O(G272) );
nand2 gate12( .a(G7), .b(G8), .O(G275) );
nand2 gate13( .a(G9), .b(G10), .O(G278) );
nand2 gate14( .a(G11), .b(G12), .O(G281) );
nand2 gate15( .a(G13), .b(G14), .O(G284) );
nand2 gate16( .a(G15), .b(G16), .O(G287) );
nand2 gate17( .a(G17), .b(G18), .O(G290) );
nand2 gate18( .a(G19), .b(G20), .O(G293) );
nand2 gate19( .a(G21), .b(G22), .O(G296) );
nand2 gate20( .a(G23), .b(G24), .O(G299) );
nand2 gate21( .a(G25), .b(G26), .O(G302) );
nand2 gate22( .a(G27), .b(G28), .O(G305) );
nand2 gate23( .a(G29), .b(G30), .O(G308) );
nand2 gate24( .a(G31), .b(G32), .O(G311) );
nand2 gate25( .a(G1), .b(G5), .O(G314) );
nand2 gate26( .a(G9), .b(G13), .O(G317) );
nand2 gate27( .a(G2), .b(G6), .O(G320) );

  xor2  gate715(.a(G14), .b(G10), .O(gate28inter0));
  nand2 gate716(.a(gate28inter0), .b(s_24), .O(gate28inter1));
  and2  gate717(.a(G14), .b(G10), .O(gate28inter2));
  inv1  gate718(.a(s_24), .O(gate28inter3));
  inv1  gate719(.a(s_25), .O(gate28inter4));
  nand2 gate720(.a(gate28inter4), .b(gate28inter3), .O(gate28inter5));
  nor2  gate721(.a(gate28inter5), .b(gate28inter2), .O(gate28inter6));
  inv1  gate722(.a(G10), .O(gate28inter7));
  inv1  gate723(.a(G14), .O(gate28inter8));
  nand2 gate724(.a(gate28inter8), .b(gate28inter7), .O(gate28inter9));
  nand2 gate725(.a(s_25), .b(gate28inter3), .O(gate28inter10));
  nor2  gate726(.a(gate28inter10), .b(gate28inter9), .O(gate28inter11));
  nor2  gate727(.a(gate28inter11), .b(gate28inter6), .O(gate28inter12));
  nand2 gate728(.a(gate28inter12), .b(gate28inter1), .O(G323));
nand2 gate29( .a(G3), .b(G7), .O(G326) );
nand2 gate30( .a(G11), .b(G15), .O(G329) );

  xor2  gate855(.a(G8), .b(G4), .O(gate31inter0));
  nand2 gate856(.a(gate31inter0), .b(s_44), .O(gate31inter1));
  and2  gate857(.a(G8), .b(G4), .O(gate31inter2));
  inv1  gate858(.a(s_44), .O(gate31inter3));
  inv1  gate859(.a(s_45), .O(gate31inter4));
  nand2 gate860(.a(gate31inter4), .b(gate31inter3), .O(gate31inter5));
  nor2  gate861(.a(gate31inter5), .b(gate31inter2), .O(gate31inter6));
  inv1  gate862(.a(G4), .O(gate31inter7));
  inv1  gate863(.a(G8), .O(gate31inter8));
  nand2 gate864(.a(gate31inter8), .b(gate31inter7), .O(gate31inter9));
  nand2 gate865(.a(s_45), .b(gate31inter3), .O(gate31inter10));
  nor2  gate866(.a(gate31inter10), .b(gate31inter9), .O(gate31inter11));
  nor2  gate867(.a(gate31inter11), .b(gate31inter6), .O(gate31inter12));
  nand2 gate868(.a(gate31inter12), .b(gate31inter1), .O(G332));
nand2 gate32( .a(G12), .b(G16), .O(G335) );
nand2 gate33( .a(G17), .b(G21), .O(G338) );
nand2 gate34( .a(G25), .b(G29), .O(G341) );
nand2 gate35( .a(G18), .b(G22), .O(G344) );
nand2 gate36( .a(G26), .b(G30), .O(G347) );
nand2 gate37( .a(G19), .b(G23), .O(G350) );
nand2 gate38( .a(G27), .b(G31), .O(G353) );
nand2 gate39( .a(G20), .b(G24), .O(G356) );
nand2 gate40( .a(G28), .b(G32), .O(G359) );
nand2 gate41( .a(G1), .b(G266), .O(G362) );
nand2 gate42( .a(G2), .b(G266), .O(G363) );

  xor2  gate701(.a(G269), .b(G3), .O(gate43inter0));
  nand2 gate702(.a(gate43inter0), .b(s_22), .O(gate43inter1));
  and2  gate703(.a(G269), .b(G3), .O(gate43inter2));
  inv1  gate704(.a(s_22), .O(gate43inter3));
  inv1  gate705(.a(s_23), .O(gate43inter4));
  nand2 gate706(.a(gate43inter4), .b(gate43inter3), .O(gate43inter5));
  nor2  gate707(.a(gate43inter5), .b(gate43inter2), .O(gate43inter6));
  inv1  gate708(.a(G3), .O(gate43inter7));
  inv1  gate709(.a(G269), .O(gate43inter8));
  nand2 gate710(.a(gate43inter8), .b(gate43inter7), .O(gate43inter9));
  nand2 gate711(.a(s_23), .b(gate43inter3), .O(gate43inter10));
  nor2  gate712(.a(gate43inter10), .b(gate43inter9), .O(gate43inter11));
  nor2  gate713(.a(gate43inter11), .b(gate43inter6), .O(gate43inter12));
  nand2 gate714(.a(gate43inter12), .b(gate43inter1), .O(G364));

  xor2  gate729(.a(G269), .b(G4), .O(gate44inter0));
  nand2 gate730(.a(gate44inter0), .b(s_26), .O(gate44inter1));
  and2  gate731(.a(G269), .b(G4), .O(gate44inter2));
  inv1  gate732(.a(s_26), .O(gate44inter3));
  inv1  gate733(.a(s_27), .O(gate44inter4));
  nand2 gate734(.a(gate44inter4), .b(gate44inter3), .O(gate44inter5));
  nor2  gate735(.a(gate44inter5), .b(gate44inter2), .O(gate44inter6));
  inv1  gate736(.a(G4), .O(gate44inter7));
  inv1  gate737(.a(G269), .O(gate44inter8));
  nand2 gate738(.a(gate44inter8), .b(gate44inter7), .O(gate44inter9));
  nand2 gate739(.a(s_27), .b(gate44inter3), .O(gate44inter10));
  nor2  gate740(.a(gate44inter10), .b(gate44inter9), .O(gate44inter11));
  nor2  gate741(.a(gate44inter11), .b(gate44inter6), .O(gate44inter12));
  nand2 gate742(.a(gate44inter12), .b(gate44inter1), .O(G365));
nand2 gate45( .a(G5), .b(G272), .O(G366) );
nand2 gate46( .a(G6), .b(G272), .O(G367) );
nand2 gate47( .a(G7), .b(G275), .O(G368) );
nand2 gate48( .a(G8), .b(G275), .O(G369) );
nand2 gate49( .a(G9), .b(G278), .O(G370) );
nand2 gate50( .a(G10), .b(G278), .O(G371) );
nand2 gate51( .a(G11), .b(G281), .O(G372) );
nand2 gate52( .a(G12), .b(G281), .O(G373) );
nand2 gate53( .a(G13), .b(G284), .O(G374) );
nand2 gate54( .a(G14), .b(G284), .O(G375) );
nand2 gate55( .a(G15), .b(G287), .O(G376) );
nand2 gate56( .a(G16), .b(G287), .O(G377) );
nand2 gate57( .a(G17), .b(G290), .O(G378) );
nand2 gate58( .a(G18), .b(G290), .O(G379) );
nand2 gate59( .a(G19), .b(G293), .O(G380) );
nand2 gate60( .a(G20), .b(G293), .O(G381) );
nand2 gate61( .a(G21), .b(G296), .O(G382) );
nand2 gate62( .a(G22), .b(G296), .O(G383) );
nand2 gate63( .a(G23), .b(G299), .O(G384) );
nand2 gate64( .a(G24), .b(G299), .O(G385) );
nand2 gate65( .a(G25), .b(G302), .O(G386) );
nand2 gate66( .a(G26), .b(G302), .O(G387) );
nand2 gate67( .a(G27), .b(G305), .O(G388) );
nand2 gate68( .a(G28), .b(G305), .O(G389) );
nand2 gate69( .a(G29), .b(G308), .O(G390) );
nand2 gate70( .a(G30), .b(G308), .O(G391) );
nand2 gate71( .a(G31), .b(G311), .O(G392) );
nand2 gate72( .a(G32), .b(G311), .O(G393) );
nand2 gate73( .a(G1), .b(G314), .O(G394) );
nand2 gate74( .a(G5), .b(G314), .O(G395) );
nand2 gate75( .a(G9), .b(G317), .O(G396) );
nand2 gate76( .a(G13), .b(G317), .O(G397) );
nand2 gate77( .a(G2), .b(G320), .O(G398) );
nand2 gate78( .a(G6), .b(G320), .O(G399) );
nand2 gate79( .a(G10), .b(G323), .O(G400) );
nand2 gate80( .a(G14), .b(G323), .O(G401) );
nand2 gate81( .a(G3), .b(G326), .O(G402) );
nand2 gate82( .a(G7), .b(G326), .O(G403) );
nand2 gate83( .a(G11), .b(G329), .O(G404) );
nand2 gate84( .a(G15), .b(G329), .O(G405) );
nand2 gate85( .a(G4), .b(G332), .O(G406) );
nand2 gate86( .a(G8), .b(G332), .O(G407) );
nand2 gate87( .a(G12), .b(G335), .O(G408) );
nand2 gate88( .a(G16), .b(G335), .O(G409) );
nand2 gate89( .a(G17), .b(G338), .O(G410) );
nand2 gate90( .a(G21), .b(G338), .O(G411) );
nand2 gate91( .a(G25), .b(G341), .O(G412) );
nand2 gate92( .a(G29), .b(G341), .O(G413) );
nand2 gate93( .a(G18), .b(G344), .O(G414) );
nand2 gate94( .a(G22), .b(G344), .O(G415) );
nand2 gate95( .a(G26), .b(G347), .O(G416) );
nand2 gate96( .a(G30), .b(G347), .O(G417) );
nand2 gate97( .a(G19), .b(G350), .O(G418) );
nand2 gate98( .a(G23), .b(G350), .O(G419) );
nand2 gate99( .a(G27), .b(G353), .O(G420) );
nand2 gate100( .a(G31), .b(G353), .O(G421) );
nand2 gate101( .a(G20), .b(G356), .O(G422) );
nand2 gate102( .a(G24), .b(G356), .O(G423) );
nand2 gate103( .a(G28), .b(G359), .O(G424) );
nand2 gate104( .a(G32), .b(G359), .O(G425) );
nand2 gate105( .a(G362), .b(G363), .O(G426) );

  xor2  gate673(.a(G365), .b(G364), .O(gate106inter0));
  nand2 gate674(.a(gate106inter0), .b(s_18), .O(gate106inter1));
  and2  gate675(.a(G365), .b(G364), .O(gate106inter2));
  inv1  gate676(.a(s_18), .O(gate106inter3));
  inv1  gate677(.a(s_19), .O(gate106inter4));
  nand2 gate678(.a(gate106inter4), .b(gate106inter3), .O(gate106inter5));
  nor2  gate679(.a(gate106inter5), .b(gate106inter2), .O(gate106inter6));
  inv1  gate680(.a(G364), .O(gate106inter7));
  inv1  gate681(.a(G365), .O(gate106inter8));
  nand2 gate682(.a(gate106inter8), .b(gate106inter7), .O(gate106inter9));
  nand2 gate683(.a(s_19), .b(gate106inter3), .O(gate106inter10));
  nor2  gate684(.a(gate106inter10), .b(gate106inter9), .O(gate106inter11));
  nor2  gate685(.a(gate106inter11), .b(gate106inter6), .O(gate106inter12));
  nand2 gate686(.a(gate106inter12), .b(gate106inter1), .O(G429));
nand2 gate107( .a(G366), .b(G367), .O(G432) );
nand2 gate108( .a(G368), .b(G369), .O(G435) );
nand2 gate109( .a(G370), .b(G371), .O(G438) );
nand2 gate110( .a(G372), .b(G373), .O(G441) );
nand2 gate111( .a(G374), .b(G375), .O(G444) );

  xor2  gate575(.a(G377), .b(G376), .O(gate112inter0));
  nand2 gate576(.a(gate112inter0), .b(s_4), .O(gate112inter1));
  and2  gate577(.a(G377), .b(G376), .O(gate112inter2));
  inv1  gate578(.a(s_4), .O(gate112inter3));
  inv1  gate579(.a(s_5), .O(gate112inter4));
  nand2 gate580(.a(gate112inter4), .b(gate112inter3), .O(gate112inter5));
  nor2  gate581(.a(gate112inter5), .b(gate112inter2), .O(gate112inter6));
  inv1  gate582(.a(G376), .O(gate112inter7));
  inv1  gate583(.a(G377), .O(gate112inter8));
  nand2 gate584(.a(gate112inter8), .b(gate112inter7), .O(gate112inter9));
  nand2 gate585(.a(s_5), .b(gate112inter3), .O(gate112inter10));
  nor2  gate586(.a(gate112inter10), .b(gate112inter9), .O(gate112inter11));
  nor2  gate587(.a(gate112inter11), .b(gate112inter6), .O(gate112inter12));
  nand2 gate588(.a(gate112inter12), .b(gate112inter1), .O(G447));
nand2 gate113( .a(G378), .b(G379), .O(G450) );
nand2 gate114( .a(G380), .b(G381), .O(G453) );

  xor2  gate743(.a(G383), .b(G382), .O(gate115inter0));
  nand2 gate744(.a(gate115inter0), .b(s_28), .O(gate115inter1));
  and2  gate745(.a(G383), .b(G382), .O(gate115inter2));
  inv1  gate746(.a(s_28), .O(gate115inter3));
  inv1  gate747(.a(s_29), .O(gate115inter4));
  nand2 gate748(.a(gate115inter4), .b(gate115inter3), .O(gate115inter5));
  nor2  gate749(.a(gate115inter5), .b(gate115inter2), .O(gate115inter6));
  inv1  gate750(.a(G382), .O(gate115inter7));
  inv1  gate751(.a(G383), .O(gate115inter8));
  nand2 gate752(.a(gate115inter8), .b(gate115inter7), .O(gate115inter9));
  nand2 gate753(.a(s_29), .b(gate115inter3), .O(gate115inter10));
  nor2  gate754(.a(gate115inter10), .b(gate115inter9), .O(gate115inter11));
  nor2  gate755(.a(gate115inter11), .b(gate115inter6), .O(gate115inter12));
  nand2 gate756(.a(gate115inter12), .b(gate115inter1), .O(G456));
nand2 gate116( .a(G384), .b(G385), .O(G459) );
nand2 gate117( .a(G386), .b(G387), .O(G462) );
nand2 gate118( .a(G388), .b(G389), .O(G465) );
nand2 gate119( .a(G390), .b(G391), .O(G468) );
nand2 gate120( .a(G392), .b(G393), .O(G471) );
nand2 gate121( .a(G394), .b(G395), .O(G474) );
nand2 gate122( .a(G396), .b(G397), .O(G477) );
nand2 gate123( .a(G398), .b(G399), .O(G480) );

  xor2  gate771(.a(G401), .b(G400), .O(gate124inter0));
  nand2 gate772(.a(gate124inter0), .b(s_32), .O(gate124inter1));
  and2  gate773(.a(G401), .b(G400), .O(gate124inter2));
  inv1  gate774(.a(s_32), .O(gate124inter3));
  inv1  gate775(.a(s_33), .O(gate124inter4));
  nand2 gate776(.a(gate124inter4), .b(gate124inter3), .O(gate124inter5));
  nor2  gate777(.a(gate124inter5), .b(gate124inter2), .O(gate124inter6));
  inv1  gate778(.a(G400), .O(gate124inter7));
  inv1  gate779(.a(G401), .O(gate124inter8));
  nand2 gate780(.a(gate124inter8), .b(gate124inter7), .O(gate124inter9));
  nand2 gate781(.a(s_33), .b(gate124inter3), .O(gate124inter10));
  nor2  gate782(.a(gate124inter10), .b(gate124inter9), .O(gate124inter11));
  nor2  gate783(.a(gate124inter11), .b(gate124inter6), .O(gate124inter12));
  nand2 gate784(.a(gate124inter12), .b(gate124inter1), .O(G483));
nand2 gate125( .a(G402), .b(G403), .O(G486) );
nand2 gate126( .a(G404), .b(G405), .O(G489) );
nand2 gate127( .a(G406), .b(G407), .O(G492) );
nand2 gate128( .a(G408), .b(G409), .O(G495) );
nand2 gate129( .a(G410), .b(G411), .O(G498) );
nand2 gate130( .a(G412), .b(G413), .O(G501) );
nand2 gate131( .a(G414), .b(G415), .O(G504) );
nand2 gate132( .a(G416), .b(G417), .O(G507) );
nand2 gate133( .a(G418), .b(G419), .O(G510) );
nand2 gate134( .a(G420), .b(G421), .O(G513) );
nand2 gate135( .a(G422), .b(G423), .O(G516) );
nand2 gate136( .a(G424), .b(G425), .O(G519) );
nand2 gate137( .a(G426), .b(G429), .O(G522) );
nand2 gate138( .a(G432), .b(G435), .O(G525) );
nand2 gate139( .a(G438), .b(G441), .O(G528) );
nand2 gate140( .a(G444), .b(G447), .O(G531) );
nand2 gate141( .a(G450), .b(G453), .O(G534) );
nand2 gate142( .a(G456), .b(G459), .O(G537) );
nand2 gate143( .a(G462), .b(G465), .O(G540) );
nand2 gate144( .a(G468), .b(G471), .O(G543) );
nand2 gate145( .a(G474), .b(G477), .O(G546) );
nand2 gate146( .a(G480), .b(G483), .O(G549) );
nand2 gate147( .a(G486), .b(G489), .O(G552) );
nand2 gate148( .a(G492), .b(G495), .O(G555) );
nand2 gate149( .a(G498), .b(G501), .O(G558) );
nand2 gate150( .a(G504), .b(G507), .O(G561) );
nand2 gate151( .a(G510), .b(G513), .O(G564) );
nand2 gate152( .a(G516), .b(G519), .O(G567) );

  xor2  gate561(.a(G522), .b(G426), .O(gate153inter0));
  nand2 gate562(.a(gate153inter0), .b(s_2), .O(gate153inter1));
  and2  gate563(.a(G522), .b(G426), .O(gate153inter2));
  inv1  gate564(.a(s_2), .O(gate153inter3));
  inv1  gate565(.a(s_3), .O(gate153inter4));
  nand2 gate566(.a(gate153inter4), .b(gate153inter3), .O(gate153inter5));
  nor2  gate567(.a(gate153inter5), .b(gate153inter2), .O(gate153inter6));
  inv1  gate568(.a(G426), .O(gate153inter7));
  inv1  gate569(.a(G522), .O(gate153inter8));
  nand2 gate570(.a(gate153inter8), .b(gate153inter7), .O(gate153inter9));
  nand2 gate571(.a(s_3), .b(gate153inter3), .O(gate153inter10));
  nor2  gate572(.a(gate153inter10), .b(gate153inter9), .O(gate153inter11));
  nor2  gate573(.a(gate153inter11), .b(gate153inter6), .O(gate153inter12));
  nand2 gate574(.a(gate153inter12), .b(gate153inter1), .O(G570));
nand2 gate154( .a(G429), .b(G522), .O(G571) );
nand2 gate155( .a(G432), .b(G525), .O(G572) );
nand2 gate156( .a(G435), .b(G525), .O(G573) );
nand2 gate157( .a(G438), .b(G528), .O(G574) );
nand2 gate158( .a(G441), .b(G528), .O(G575) );
nand2 gate159( .a(G444), .b(G531), .O(G576) );
nand2 gate160( .a(G447), .b(G531), .O(G577) );

  xor2  gate799(.a(G534), .b(G450), .O(gate161inter0));
  nand2 gate800(.a(gate161inter0), .b(s_36), .O(gate161inter1));
  and2  gate801(.a(G534), .b(G450), .O(gate161inter2));
  inv1  gate802(.a(s_36), .O(gate161inter3));
  inv1  gate803(.a(s_37), .O(gate161inter4));
  nand2 gate804(.a(gate161inter4), .b(gate161inter3), .O(gate161inter5));
  nor2  gate805(.a(gate161inter5), .b(gate161inter2), .O(gate161inter6));
  inv1  gate806(.a(G450), .O(gate161inter7));
  inv1  gate807(.a(G534), .O(gate161inter8));
  nand2 gate808(.a(gate161inter8), .b(gate161inter7), .O(gate161inter9));
  nand2 gate809(.a(s_37), .b(gate161inter3), .O(gate161inter10));
  nor2  gate810(.a(gate161inter10), .b(gate161inter9), .O(gate161inter11));
  nor2  gate811(.a(gate161inter11), .b(gate161inter6), .O(gate161inter12));
  nand2 gate812(.a(gate161inter12), .b(gate161inter1), .O(G578));
nand2 gate162( .a(G453), .b(G534), .O(G579) );
nand2 gate163( .a(G456), .b(G537), .O(G580) );
nand2 gate164( .a(G459), .b(G537), .O(G581) );
nand2 gate165( .a(G462), .b(G540), .O(G582) );
nand2 gate166( .a(G465), .b(G540), .O(G583) );
nand2 gate167( .a(G468), .b(G543), .O(G584) );
nand2 gate168( .a(G471), .b(G543), .O(G585) );
nand2 gate169( .a(G474), .b(G546), .O(G586) );
nand2 gate170( .a(G477), .b(G546), .O(G587) );
nand2 gate171( .a(G480), .b(G549), .O(G588) );
nand2 gate172( .a(G483), .b(G549), .O(G589) );
nand2 gate173( .a(G486), .b(G552), .O(G590) );
nand2 gate174( .a(G489), .b(G552), .O(G591) );
nand2 gate175( .a(G492), .b(G555), .O(G592) );
nand2 gate176( .a(G495), .b(G555), .O(G593) );
nand2 gate177( .a(G498), .b(G558), .O(G594) );
nand2 gate178( .a(G501), .b(G558), .O(G595) );

  xor2  gate939(.a(G561), .b(G504), .O(gate179inter0));
  nand2 gate940(.a(gate179inter0), .b(s_56), .O(gate179inter1));
  and2  gate941(.a(G561), .b(G504), .O(gate179inter2));
  inv1  gate942(.a(s_56), .O(gate179inter3));
  inv1  gate943(.a(s_57), .O(gate179inter4));
  nand2 gate944(.a(gate179inter4), .b(gate179inter3), .O(gate179inter5));
  nor2  gate945(.a(gate179inter5), .b(gate179inter2), .O(gate179inter6));
  inv1  gate946(.a(G504), .O(gate179inter7));
  inv1  gate947(.a(G561), .O(gate179inter8));
  nand2 gate948(.a(gate179inter8), .b(gate179inter7), .O(gate179inter9));
  nand2 gate949(.a(s_57), .b(gate179inter3), .O(gate179inter10));
  nor2  gate950(.a(gate179inter10), .b(gate179inter9), .O(gate179inter11));
  nor2  gate951(.a(gate179inter11), .b(gate179inter6), .O(gate179inter12));
  nand2 gate952(.a(gate179inter12), .b(gate179inter1), .O(G596));
nand2 gate180( .a(G507), .b(G561), .O(G597) );
nand2 gate181( .a(G510), .b(G564), .O(G598) );
nand2 gate182( .a(G513), .b(G564), .O(G599) );

  xor2  gate603(.a(G567), .b(G516), .O(gate183inter0));
  nand2 gate604(.a(gate183inter0), .b(s_8), .O(gate183inter1));
  and2  gate605(.a(G567), .b(G516), .O(gate183inter2));
  inv1  gate606(.a(s_8), .O(gate183inter3));
  inv1  gate607(.a(s_9), .O(gate183inter4));
  nand2 gate608(.a(gate183inter4), .b(gate183inter3), .O(gate183inter5));
  nor2  gate609(.a(gate183inter5), .b(gate183inter2), .O(gate183inter6));
  inv1  gate610(.a(G516), .O(gate183inter7));
  inv1  gate611(.a(G567), .O(gate183inter8));
  nand2 gate612(.a(gate183inter8), .b(gate183inter7), .O(gate183inter9));
  nand2 gate613(.a(s_9), .b(gate183inter3), .O(gate183inter10));
  nor2  gate614(.a(gate183inter10), .b(gate183inter9), .O(gate183inter11));
  nor2  gate615(.a(gate183inter11), .b(gate183inter6), .O(gate183inter12));
  nand2 gate616(.a(gate183inter12), .b(gate183inter1), .O(G600));
nand2 gate184( .a(G519), .b(G567), .O(G601) );
nand2 gate185( .a(G570), .b(G571), .O(G602) );

  xor2  gate869(.a(G573), .b(G572), .O(gate186inter0));
  nand2 gate870(.a(gate186inter0), .b(s_46), .O(gate186inter1));
  and2  gate871(.a(G573), .b(G572), .O(gate186inter2));
  inv1  gate872(.a(s_46), .O(gate186inter3));
  inv1  gate873(.a(s_47), .O(gate186inter4));
  nand2 gate874(.a(gate186inter4), .b(gate186inter3), .O(gate186inter5));
  nor2  gate875(.a(gate186inter5), .b(gate186inter2), .O(gate186inter6));
  inv1  gate876(.a(G572), .O(gate186inter7));
  inv1  gate877(.a(G573), .O(gate186inter8));
  nand2 gate878(.a(gate186inter8), .b(gate186inter7), .O(gate186inter9));
  nand2 gate879(.a(s_47), .b(gate186inter3), .O(gate186inter10));
  nor2  gate880(.a(gate186inter10), .b(gate186inter9), .O(gate186inter11));
  nor2  gate881(.a(gate186inter11), .b(gate186inter6), .O(gate186inter12));
  nand2 gate882(.a(gate186inter12), .b(gate186inter1), .O(G607));
nand2 gate187( .a(G574), .b(G575), .O(G612) );
nand2 gate188( .a(G576), .b(G577), .O(G617) );
nand2 gate189( .a(G578), .b(G579), .O(G622) );

  xor2  gate911(.a(G581), .b(G580), .O(gate190inter0));
  nand2 gate912(.a(gate190inter0), .b(s_52), .O(gate190inter1));
  and2  gate913(.a(G581), .b(G580), .O(gate190inter2));
  inv1  gate914(.a(s_52), .O(gate190inter3));
  inv1  gate915(.a(s_53), .O(gate190inter4));
  nand2 gate916(.a(gate190inter4), .b(gate190inter3), .O(gate190inter5));
  nor2  gate917(.a(gate190inter5), .b(gate190inter2), .O(gate190inter6));
  inv1  gate918(.a(G580), .O(gate190inter7));
  inv1  gate919(.a(G581), .O(gate190inter8));
  nand2 gate920(.a(gate190inter8), .b(gate190inter7), .O(gate190inter9));
  nand2 gate921(.a(s_53), .b(gate190inter3), .O(gate190inter10));
  nor2  gate922(.a(gate190inter10), .b(gate190inter9), .O(gate190inter11));
  nor2  gate923(.a(gate190inter11), .b(gate190inter6), .O(gate190inter12));
  nand2 gate924(.a(gate190inter12), .b(gate190inter1), .O(G627));
nand2 gate191( .a(G582), .b(G583), .O(G632) );
nand2 gate192( .a(G584), .b(G585), .O(G637) );
nand2 gate193( .a(G586), .b(G587), .O(G642) );
nand2 gate194( .a(G588), .b(G589), .O(G645) );
nand2 gate195( .a(G590), .b(G591), .O(G648) );
nand2 gate196( .a(G592), .b(G593), .O(G651) );
nand2 gate197( .a(G594), .b(G595), .O(G654) );
nand2 gate198( .a(G596), .b(G597), .O(G657) );
nand2 gate199( .a(G598), .b(G599), .O(G660) );
nand2 gate200( .a(G600), .b(G601), .O(G663) );
nand2 gate201( .a(G602), .b(G607), .O(G666) );
nand2 gate202( .a(G612), .b(G617), .O(G669) );
nand2 gate203( .a(G602), .b(G612), .O(G672) );
nand2 gate204( .a(G607), .b(G617), .O(G675) );

  xor2  gate841(.a(G627), .b(G622), .O(gate205inter0));
  nand2 gate842(.a(gate205inter0), .b(s_42), .O(gate205inter1));
  and2  gate843(.a(G627), .b(G622), .O(gate205inter2));
  inv1  gate844(.a(s_42), .O(gate205inter3));
  inv1  gate845(.a(s_43), .O(gate205inter4));
  nand2 gate846(.a(gate205inter4), .b(gate205inter3), .O(gate205inter5));
  nor2  gate847(.a(gate205inter5), .b(gate205inter2), .O(gate205inter6));
  inv1  gate848(.a(G622), .O(gate205inter7));
  inv1  gate849(.a(G627), .O(gate205inter8));
  nand2 gate850(.a(gate205inter8), .b(gate205inter7), .O(gate205inter9));
  nand2 gate851(.a(s_43), .b(gate205inter3), .O(gate205inter10));
  nor2  gate852(.a(gate205inter10), .b(gate205inter9), .O(gate205inter11));
  nor2  gate853(.a(gate205inter11), .b(gate205inter6), .O(gate205inter12));
  nand2 gate854(.a(gate205inter12), .b(gate205inter1), .O(G678));
nand2 gate206( .a(G632), .b(G637), .O(G681) );
nand2 gate207( .a(G622), .b(G632), .O(G684) );
nand2 gate208( .a(G627), .b(G637), .O(G687) );
nand2 gate209( .a(G602), .b(G666), .O(G690) );
nand2 gate210( .a(G607), .b(G666), .O(G691) );
nand2 gate211( .a(G612), .b(G669), .O(G692) );
nand2 gate212( .a(G617), .b(G669), .O(G693) );
nand2 gate213( .a(G602), .b(G672), .O(G694) );
nand2 gate214( .a(G612), .b(G672), .O(G695) );
nand2 gate215( .a(G607), .b(G675), .O(G696) );
nand2 gate216( .a(G617), .b(G675), .O(G697) );
nand2 gate217( .a(G622), .b(G678), .O(G698) );
nand2 gate218( .a(G627), .b(G678), .O(G699) );
nand2 gate219( .a(G632), .b(G681), .O(G700) );
nand2 gate220( .a(G637), .b(G681), .O(G701) );

  xor2  gate617(.a(G684), .b(G622), .O(gate221inter0));
  nand2 gate618(.a(gate221inter0), .b(s_10), .O(gate221inter1));
  and2  gate619(.a(G684), .b(G622), .O(gate221inter2));
  inv1  gate620(.a(s_10), .O(gate221inter3));
  inv1  gate621(.a(s_11), .O(gate221inter4));
  nand2 gate622(.a(gate221inter4), .b(gate221inter3), .O(gate221inter5));
  nor2  gate623(.a(gate221inter5), .b(gate221inter2), .O(gate221inter6));
  inv1  gate624(.a(G622), .O(gate221inter7));
  inv1  gate625(.a(G684), .O(gate221inter8));
  nand2 gate626(.a(gate221inter8), .b(gate221inter7), .O(gate221inter9));
  nand2 gate627(.a(s_11), .b(gate221inter3), .O(gate221inter10));
  nor2  gate628(.a(gate221inter10), .b(gate221inter9), .O(gate221inter11));
  nor2  gate629(.a(gate221inter11), .b(gate221inter6), .O(gate221inter12));
  nand2 gate630(.a(gate221inter12), .b(gate221inter1), .O(G702));
nand2 gate222( .a(G632), .b(G684), .O(G703) );
nand2 gate223( .a(G627), .b(G687), .O(G704) );
nand2 gate224( .a(G637), .b(G687), .O(G705) );
nand2 gate225( .a(G690), .b(G691), .O(G706) );
nand2 gate226( .a(G692), .b(G693), .O(G709) );
nand2 gate227( .a(G694), .b(G695), .O(G712) );
nand2 gate228( .a(G696), .b(G697), .O(G715) );
nand2 gate229( .a(G698), .b(G699), .O(G718) );
nand2 gate230( .a(G700), .b(G701), .O(G721) );
nand2 gate231( .a(G702), .b(G703), .O(G724) );
nand2 gate232( .a(G704), .b(G705), .O(G727) );
nand2 gate233( .a(G242), .b(G718), .O(G730) );

  xor2  gate645(.a(G721), .b(G245), .O(gate234inter0));
  nand2 gate646(.a(gate234inter0), .b(s_14), .O(gate234inter1));
  and2  gate647(.a(G721), .b(G245), .O(gate234inter2));
  inv1  gate648(.a(s_14), .O(gate234inter3));
  inv1  gate649(.a(s_15), .O(gate234inter4));
  nand2 gate650(.a(gate234inter4), .b(gate234inter3), .O(gate234inter5));
  nor2  gate651(.a(gate234inter5), .b(gate234inter2), .O(gate234inter6));
  inv1  gate652(.a(G245), .O(gate234inter7));
  inv1  gate653(.a(G721), .O(gate234inter8));
  nand2 gate654(.a(gate234inter8), .b(gate234inter7), .O(gate234inter9));
  nand2 gate655(.a(s_15), .b(gate234inter3), .O(gate234inter10));
  nor2  gate656(.a(gate234inter10), .b(gate234inter9), .O(gate234inter11));
  nor2  gate657(.a(gate234inter11), .b(gate234inter6), .O(gate234inter12));
  nand2 gate658(.a(gate234inter12), .b(gate234inter1), .O(G733));
nand2 gate235( .a(G248), .b(G724), .O(G736) );
nand2 gate236( .a(G251), .b(G727), .O(G739) );
nand2 gate237( .a(G254), .b(G706), .O(G742) );

  xor2  gate883(.a(G709), .b(G257), .O(gate238inter0));
  nand2 gate884(.a(gate238inter0), .b(s_48), .O(gate238inter1));
  and2  gate885(.a(G709), .b(G257), .O(gate238inter2));
  inv1  gate886(.a(s_48), .O(gate238inter3));
  inv1  gate887(.a(s_49), .O(gate238inter4));
  nand2 gate888(.a(gate238inter4), .b(gate238inter3), .O(gate238inter5));
  nor2  gate889(.a(gate238inter5), .b(gate238inter2), .O(gate238inter6));
  inv1  gate890(.a(G257), .O(gate238inter7));
  inv1  gate891(.a(G709), .O(gate238inter8));
  nand2 gate892(.a(gate238inter8), .b(gate238inter7), .O(gate238inter9));
  nand2 gate893(.a(s_49), .b(gate238inter3), .O(gate238inter10));
  nor2  gate894(.a(gate238inter10), .b(gate238inter9), .O(gate238inter11));
  nor2  gate895(.a(gate238inter11), .b(gate238inter6), .O(gate238inter12));
  nand2 gate896(.a(gate238inter12), .b(gate238inter1), .O(G745));
nand2 gate239( .a(G260), .b(G712), .O(G748) );
nand2 gate240( .a(G263), .b(G715), .O(G751) );
nand2 gate241( .a(G242), .b(G730), .O(G754) );
nand2 gate242( .a(G718), .b(G730), .O(G755) );
nand2 gate243( .a(G245), .b(G733), .O(G756) );
nand2 gate244( .a(G721), .b(G733), .O(G757) );
nand2 gate245( .a(G248), .b(G736), .O(G758) );
nand2 gate246( .a(G724), .b(G736), .O(G759) );
nand2 gate247( .a(G251), .b(G739), .O(G760) );
nand2 gate248( .a(G727), .b(G739), .O(G761) );
nand2 gate249( .a(G254), .b(G742), .O(G762) );
nand2 gate250( .a(G706), .b(G742), .O(G763) );
nand2 gate251( .a(G257), .b(G745), .O(G764) );
nand2 gate252( .a(G709), .b(G745), .O(G765) );
nand2 gate253( .a(G260), .b(G748), .O(G766) );

  xor2  gate589(.a(G748), .b(G712), .O(gate254inter0));
  nand2 gate590(.a(gate254inter0), .b(s_6), .O(gate254inter1));
  and2  gate591(.a(G748), .b(G712), .O(gate254inter2));
  inv1  gate592(.a(s_6), .O(gate254inter3));
  inv1  gate593(.a(s_7), .O(gate254inter4));
  nand2 gate594(.a(gate254inter4), .b(gate254inter3), .O(gate254inter5));
  nor2  gate595(.a(gate254inter5), .b(gate254inter2), .O(gate254inter6));
  inv1  gate596(.a(G712), .O(gate254inter7));
  inv1  gate597(.a(G748), .O(gate254inter8));
  nand2 gate598(.a(gate254inter8), .b(gate254inter7), .O(gate254inter9));
  nand2 gate599(.a(s_7), .b(gate254inter3), .O(gate254inter10));
  nor2  gate600(.a(gate254inter10), .b(gate254inter9), .O(gate254inter11));
  nor2  gate601(.a(gate254inter11), .b(gate254inter6), .O(gate254inter12));
  nand2 gate602(.a(gate254inter12), .b(gate254inter1), .O(G767));
nand2 gate255( .a(G263), .b(G751), .O(G768) );
nand2 gate256( .a(G715), .b(G751), .O(G769) );
nand2 gate257( .a(G754), .b(G755), .O(G770) );
nand2 gate258( .a(G756), .b(G757), .O(G773) );
nand2 gate259( .a(G758), .b(G759), .O(G776) );
nand2 gate260( .a(G760), .b(G761), .O(G779) );
nand2 gate261( .a(G762), .b(G763), .O(G782) );
nand2 gate262( .a(G764), .b(G765), .O(G785) );
nand2 gate263( .a(G766), .b(G767), .O(G788) );
nand2 gate264( .a(G768), .b(G769), .O(G791) );
nand2 gate265( .a(G642), .b(G770), .O(G794) );
nand2 gate266( .a(G645), .b(G773), .O(G797) );
nand2 gate267( .a(G648), .b(G776), .O(G800) );
nand2 gate268( .a(G651), .b(G779), .O(G803) );
nand2 gate269( .a(G654), .b(G782), .O(G806) );
nand2 gate270( .a(G657), .b(G785), .O(G809) );
nand2 gate271( .a(G660), .b(G788), .O(G812) );
nand2 gate272( .a(G663), .b(G791), .O(G815) );
nand2 gate273( .a(G642), .b(G794), .O(G818) );
nand2 gate274( .a(G770), .b(G794), .O(G819) );

  xor2  gate547(.a(G797), .b(G645), .O(gate275inter0));
  nand2 gate548(.a(gate275inter0), .b(s_0), .O(gate275inter1));
  and2  gate549(.a(G797), .b(G645), .O(gate275inter2));
  inv1  gate550(.a(s_0), .O(gate275inter3));
  inv1  gate551(.a(s_1), .O(gate275inter4));
  nand2 gate552(.a(gate275inter4), .b(gate275inter3), .O(gate275inter5));
  nor2  gate553(.a(gate275inter5), .b(gate275inter2), .O(gate275inter6));
  inv1  gate554(.a(G645), .O(gate275inter7));
  inv1  gate555(.a(G797), .O(gate275inter8));
  nand2 gate556(.a(gate275inter8), .b(gate275inter7), .O(gate275inter9));
  nand2 gate557(.a(s_1), .b(gate275inter3), .O(gate275inter10));
  nor2  gate558(.a(gate275inter10), .b(gate275inter9), .O(gate275inter11));
  nor2  gate559(.a(gate275inter11), .b(gate275inter6), .O(gate275inter12));
  nand2 gate560(.a(gate275inter12), .b(gate275inter1), .O(G820));

  xor2  gate659(.a(G797), .b(G773), .O(gate276inter0));
  nand2 gate660(.a(gate276inter0), .b(s_16), .O(gate276inter1));
  and2  gate661(.a(G797), .b(G773), .O(gate276inter2));
  inv1  gate662(.a(s_16), .O(gate276inter3));
  inv1  gate663(.a(s_17), .O(gate276inter4));
  nand2 gate664(.a(gate276inter4), .b(gate276inter3), .O(gate276inter5));
  nor2  gate665(.a(gate276inter5), .b(gate276inter2), .O(gate276inter6));
  inv1  gate666(.a(G773), .O(gate276inter7));
  inv1  gate667(.a(G797), .O(gate276inter8));
  nand2 gate668(.a(gate276inter8), .b(gate276inter7), .O(gate276inter9));
  nand2 gate669(.a(s_17), .b(gate276inter3), .O(gate276inter10));
  nor2  gate670(.a(gate276inter10), .b(gate276inter9), .O(gate276inter11));
  nor2  gate671(.a(gate276inter11), .b(gate276inter6), .O(gate276inter12));
  nand2 gate672(.a(gate276inter12), .b(gate276inter1), .O(G821));
nand2 gate277( .a(G648), .b(G800), .O(G822) );
nand2 gate278( .a(G776), .b(G800), .O(G823) );
nand2 gate279( .a(G651), .b(G803), .O(G824) );
nand2 gate280( .a(G779), .b(G803), .O(G825) );

  xor2  gate967(.a(G806), .b(G654), .O(gate281inter0));
  nand2 gate968(.a(gate281inter0), .b(s_60), .O(gate281inter1));
  and2  gate969(.a(G806), .b(G654), .O(gate281inter2));
  inv1  gate970(.a(s_60), .O(gate281inter3));
  inv1  gate971(.a(s_61), .O(gate281inter4));
  nand2 gate972(.a(gate281inter4), .b(gate281inter3), .O(gate281inter5));
  nor2  gate973(.a(gate281inter5), .b(gate281inter2), .O(gate281inter6));
  inv1  gate974(.a(G654), .O(gate281inter7));
  inv1  gate975(.a(G806), .O(gate281inter8));
  nand2 gate976(.a(gate281inter8), .b(gate281inter7), .O(gate281inter9));
  nand2 gate977(.a(s_61), .b(gate281inter3), .O(gate281inter10));
  nor2  gate978(.a(gate281inter10), .b(gate281inter9), .O(gate281inter11));
  nor2  gate979(.a(gate281inter11), .b(gate281inter6), .O(gate281inter12));
  nand2 gate980(.a(gate281inter12), .b(gate281inter1), .O(G826));
nand2 gate282( .a(G782), .b(G806), .O(G827) );
nand2 gate283( .a(G657), .b(G809), .O(G828) );
nand2 gate284( .a(G785), .b(G809), .O(G829) );
nand2 gate285( .a(G660), .b(G812), .O(G830) );
nand2 gate286( .a(G788), .b(G812), .O(G831) );
nand2 gate287( .a(G663), .b(G815), .O(G832) );
nand2 gate288( .a(G791), .b(G815), .O(G833) );
nand2 gate289( .a(G818), .b(G819), .O(G834) );
nand2 gate290( .a(G820), .b(G821), .O(G847) );
nand2 gate291( .a(G822), .b(G823), .O(G860) );
nand2 gate292( .a(G824), .b(G825), .O(G873) );
nand2 gate293( .a(G828), .b(G829), .O(G886) );
nand2 gate294( .a(G832), .b(G833), .O(G899) );

  xor2  gate897(.a(G831), .b(G830), .O(gate295inter0));
  nand2 gate898(.a(gate295inter0), .b(s_50), .O(gate295inter1));
  and2  gate899(.a(G831), .b(G830), .O(gate295inter2));
  inv1  gate900(.a(s_50), .O(gate295inter3));
  inv1  gate901(.a(s_51), .O(gate295inter4));
  nand2 gate902(.a(gate295inter4), .b(gate295inter3), .O(gate295inter5));
  nor2  gate903(.a(gate295inter5), .b(gate295inter2), .O(gate295inter6));
  inv1  gate904(.a(G830), .O(gate295inter7));
  inv1  gate905(.a(G831), .O(gate295inter8));
  nand2 gate906(.a(gate295inter8), .b(gate295inter7), .O(gate295inter9));
  nand2 gate907(.a(s_51), .b(gate295inter3), .O(gate295inter10));
  nor2  gate908(.a(gate295inter10), .b(gate295inter9), .O(gate295inter11));
  nor2  gate909(.a(gate295inter11), .b(gate295inter6), .O(gate295inter12));
  nand2 gate910(.a(gate295inter12), .b(gate295inter1), .O(G912));
nand2 gate296( .a(G826), .b(G827), .O(G925) );
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );
nand2 gate387( .a(G1), .b(G1036), .O(G1132) );
nand2 gate388( .a(G2), .b(G1039), .O(G1135) );
nand2 gate389( .a(G3), .b(G1042), .O(G1138) );

  xor2  gate631(.a(G1045), .b(G4), .O(gate390inter0));
  nand2 gate632(.a(gate390inter0), .b(s_12), .O(gate390inter1));
  and2  gate633(.a(G1045), .b(G4), .O(gate390inter2));
  inv1  gate634(.a(s_12), .O(gate390inter3));
  inv1  gate635(.a(s_13), .O(gate390inter4));
  nand2 gate636(.a(gate390inter4), .b(gate390inter3), .O(gate390inter5));
  nor2  gate637(.a(gate390inter5), .b(gate390inter2), .O(gate390inter6));
  inv1  gate638(.a(G4), .O(gate390inter7));
  inv1  gate639(.a(G1045), .O(gate390inter8));
  nand2 gate640(.a(gate390inter8), .b(gate390inter7), .O(gate390inter9));
  nand2 gate641(.a(s_13), .b(gate390inter3), .O(gate390inter10));
  nor2  gate642(.a(gate390inter10), .b(gate390inter9), .O(gate390inter11));
  nor2  gate643(.a(gate390inter11), .b(gate390inter6), .O(gate390inter12));
  nand2 gate644(.a(gate390inter12), .b(gate390inter1), .O(G1141));
nand2 gate391( .a(G5), .b(G1048), .O(G1144) );
nand2 gate392( .a(G6), .b(G1051), .O(G1147) );
nand2 gate393( .a(G7), .b(G1054), .O(G1150) );
nand2 gate394( .a(G8), .b(G1057), .O(G1153) );
nand2 gate395( .a(G9), .b(G1060), .O(G1156) );
nand2 gate396( .a(G10), .b(G1063), .O(G1159) );

  xor2  gate757(.a(G1066), .b(G11), .O(gate397inter0));
  nand2 gate758(.a(gate397inter0), .b(s_30), .O(gate397inter1));
  and2  gate759(.a(G1066), .b(G11), .O(gate397inter2));
  inv1  gate760(.a(s_30), .O(gate397inter3));
  inv1  gate761(.a(s_31), .O(gate397inter4));
  nand2 gate762(.a(gate397inter4), .b(gate397inter3), .O(gate397inter5));
  nor2  gate763(.a(gate397inter5), .b(gate397inter2), .O(gate397inter6));
  inv1  gate764(.a(G11), .O(gate397inter7));
  inv1  gate765(.a(G1066), .O(gate397inter8));
  nand2 gate766(.a(gate397inter8), .b(gate397inter7), .O(gate397inter9));
  nand2 gate767(.a(s_31), .b(gate397inter3), .O(gate397inter10));
  nor2  gate768(.a(gate397inter10), .b(gate397inter9), .O(gate397inter11));
  nor2  gate769(.a(gate397inter11), .b(gate397inter6), .O(gate397inter12));
  nand2 gate770(.a(gate397inter12), .b(gate397inter1), .O(G1162));
nand2 gate398( .a(G12), .b(G1069), .O(G1165) );
nand2 gate399( .a(G13), .b(G1072), .O(G1168) );
nand2 gate400( .a(G14), .b(G1075), .O(G1171) );
nand2 gate401( .a(G15), .b(G1078), .O(G1174) );
nand2 gate402( .a(G16), .b(G1081), .O(G1177) );
nand2 gate403( .a(G17), .b(G1084), .O(G1180) );
nand2 gate404( .a(G18), .b(G1087), .O(G1183) );
nand2 gate405( .a(G19), .b(G1090), .O(G1186) );
nand2 gate406( .a(G20), .b(G1093), .O(G1189) );
nand2 gate407( .a(G21), .b(G1096), .O(G1192) );
nand2 gate408( .a(G22), .b(G1099), .O(G1195) );
nand2 gate409( .a(G23), .b(G1102), .O(G1198) );
nand2 gate410( .a(G24), .b(G1105), .O(G1201) );
nand2 gate411( .a(G25), .b(G1108), .O(G1204) );
nand2 gate412( .a(G26), .b(G1111), .O(G1207) );
nand2 gate413( .a(G27), .b(G1114), .O(G1210) );
nand2 gate414( .a(G28), .b(G1117), .O(G1213) );
nand2 gate415( .a(G29), .b(G1120), .O(G1216) );
nand2 gate416( .a(G30), .b(G1123), .O(G1219) );
nand2 gate417( .a(G31), .b(G1126), .O(G1222) );
nand2 gate418( .a(G32), .b(G1129), .O(G1225) );
nand2 gate419( .a(G1), .b(G1132), .O(G1228) );
nand2 gate420( .a(G1036), .b(G1132), .O(G1229) );
nand2 gate421( .a(G2), .b(G1135), .O(G1230) );
nand2 gate422( .a(G1039), .b(G1135), .O(G1231) );
nand2 gate423( .a(G3), .b(G1138), .O(G1232) );
nand2 gate424( .a(G1042), .b(G1138), .O(G1233) );
nand2 gate425( .a(G4), .b(G1141), .O(G1234) );
nand2 gate426( .a(G1045), .b(G1141), .O(G1235) );
nand2 gate427( .a(G5), .b(G1144), .O(G1236) );
nand2 gate428( .a(G1048), .b(G1144), .O(G1237) );
nand2 gate429( .a(G6), .b(G1147), .O(G1238) );
nand2 gate430( .a(G1051), .b(G1147), .O(G1239) );

  xor2  gate813(.a(G1150), .b(G7), .O(gate431inter0));
  nand2 gate814(.a(gate431inter0), .b(s_38), .O(gate431inter1));
  and2  gate815(.a(G1150), .b(G7), .O(gate431inter2));
  inv1  gate816(.a(s_38), .O(gate431inter3));
  inv1  gate817(.a(s_39), .O(gate431inter4));
  nand2 gate818(.a(gate431inter4), .b(gate431inter3), .O(gate431inter5));
  nor2  gate819(.a(gate431inter5), .b(gate431inter2), .O(gate431inter6));
  inv1  gate820(.a(G7), .O(gate431inter7));
  inv1  gate821(.a(G1150), .O(gate431inter8));
  nand2 gate822(.a(gate431inter8), .b(gate431inter7), .O(gate431inter9));
  nand2 gate823(.a(s_39), .b(gate431inter3), .O(gate431inter10));
  nor2  gate824(.a(gate431inter10), .b(gate431inter9), .O(gate431inter11));
  nor2  gate825(.a(gate431inter11), .b(gate431inter6), .O(gate431inter12));
  nand2 gate826(.a(gate431inter12), .b(gate431inter1), .O(G1240));
nand2 gate432( .a(G1054), .b(G1150), .O(G1241) );
nand2 gate433( .a(G8), .b(G1153), .O(G1242) );
nand2 gate434( .a(G1057), .b(G1153), .O(G1243) );
nand2 gate435( .a(G9), .b(G1156), .O(G1244) );
nand2 gate436( .a(G1060), .b(G1156), .O(G1245) );
nand2 gate437( .a(G10), .b(G1159), .O(G1246) );
nand2 gate438( .a(G1063), .b(G1159), .O(G1247) );
nand2 gate439( .a(G11), .b(G1162), .O(G1248) );
nand2 gate440( .a(G1066), .b(G1162), .O(G1249) );
nand2 gate441( .a(G12), .b(G1165), .O(G1250) );
nand2 gate442( .a(G1069), .b(G1165), .O(G1251) );
nand2 gate443( .a(G13), .b(G1168), .O(G1252) );
nand2 gate444( .a(G1072), .b(G1168), .O(G1253) );
nand2 gate445( .a(G14), .b(G1171), .O(G1254) );
nand2 gate446( .a(G1075), .b(G1171), .O(G1255) );
nand2 gate447( .a(G15), .b(G1174), .O(G1256) );
nand2 gate448( .a(G1078), .b(G1174), .O(G1257) );
nand2 gate449( .a(G16), .b(G1177), .O(G1258) );
nand2 gate450( .a(G1081), .b(G1177), .O(G1259) );
nand2 gate451( .a(G17), .b(G1180), .O(G1260) );
nand2 gate452( .a(G1084), .b(G1180), .O(G1261) );
nand2 gate453( .a(G18), .b(G1183), .O(G1262) );
nand2 gate454( .a(G1087), .b(G1183), .O(G1263) );
nand2 gate455( .a(G19), .b(G1186), .O(G1264) );
nand2 gate456( .a(G1090), .b(G1186), .O(G1265) );

  xor2  gate925(.a(G1189), .b(G20), .O(gate457inter0));
  nand2 gate926(.a(gate457inter0), .b(s_54), .O(gate457inter1));
  and2  gate927(.a(G1189), .b(G20), .O(gate457inter2));
  inv1  gate928(.a(s_54), .O(gate457inter3));
  inv1  gate929(.a(s_55), .O(gate457inter4));
  nand2 gate930(.a(gate457inter4), .b(gate457inter3), .O(gate457inter5));
  nor2  gate931(.a(gate457inter5), .b(gate457inter2), .O(gate457inter6));
  inv1  gate932(.a(G20), .O(gate457inter7));
  inv1  gate933(.a(G1189), .O(gate457inter8));
  nand2 gate934(.a(gate457inter8), .b(gate457inter7), .O(gate457inter9));
  nand2 gate935(.a(s_55), .b(gate457inter3), .O(gate457inter10));
  nor2  gate936(.a(gate457inter10), .b(gate457inter9), .O(gate457inter11));
  nor2  gate937(.a(gate457inter11), .b(gate457inter6), .O(gate457inter12));
  nand2 gate938(.a(gate457inter12), .b(gate457inter1), .O(G1266));
nand2 gate458( .a(G1093), .b(G1189), .O(G1267) );
nand2 gate459( .a(G21), .b(G1192), .O(G1268) );
nand2 gate460( .a(G1096), .b(G1192), .O(G1269) );
nand2 gate461( .a(G22), .b(G1195), .O(G1270) );
nand2 gate462( .a(G1099), .b(G1195), .O(G1271) );
nand2 gate463( .a(G23), .b(G1198), .O(G1272) );
nand2 gate464( .a(G1102), .b(G1198), .O(G1273) );
nand2 gate465( .a(G24), .b(G1201), .O(G1274) );
nand2 gate466( .a(G1105), .b(G1201), .O(G1275) );
nand2 gate467( .a(G25), .b(G1204), .O(G1276) );

  xor2  gate785(.a(G1204), .b(G1108), .O(gate468inter0));
  nand2 gate786(.a(gate468inter0), .b(s_34), .O(gate468inter1));
  and2  gate787(.a(G1204), .b(G1108), .O(gate468inter2));
  inv1  gate788(.a(s_34), .O(gate468inter3));
  inv1  gate789(.a(s_35), .O(gate468inter4));
  nand2 gate790(.a(gate468inter4), .b(gate468inter3), .O(gate468inter5));
  nor2  gate791(.a(gate468inter5), .b(gate468inter2), .O(gate468inter6));
  inv1  gate792(.a(G1108), .O(gate468inter7));
  inv1  gate793(.a(G1204), .O(gate468inter8));
  nand2 gate794(.a(gate468inter8), .b(gate468inter7), .O(gate468inter9));
  nand2 gate795(.a(s_35), .b(gate468inter3), .O(gate468inter10));
  nor2  gate796(.a(gate468inter10), .b(gate468inter9), .O(gate468inter11));
  nor2  gate797(.a(gate468inter11), .b(gate468inter6), .O(gate468inter12));
  nand2 gate798(.a(gate468inter12), .b(gate468inter1), .O(G1277));
nand2 gate469( .a(G26), .b(G1207), .O(G1278) );
nand2 gate470( .a(G1111), .b(G1207), .O(G1279) );
nand2 gate471( .a(G27), .b(G1210), .O(G1280) );
nand2 gate472( .a(G1114), .b(G1210), .O(G1281) );
nand2 gate473( .a(G28), .b(G1213), .O(G1282) );
nand2 gate474( .a(G1117), .b(G1213), .O(G1283) );
nand2 gate475( .a(G29), .b(G1216), .O(G1284) );
nand2 gate476( .a(G1120), .b(G1216), .O(G1285) );
nand2 gate477( .a(G30), .b(G1219), .O(G1286) );
nand2 gate478( .a(G1123), .b(G1219), .O(G1287) );
nand2 gate479( .a(G31), .b(G1222), .O(G1288) );

  xor2  gate953(.a(G1222), .b(G1126), .O(gate480inter0));
  nand2 gate954(.a(gate480inter0), .b(s_58), .O(gate480inter1));
  and2  gate955(.a(G1222), .b(G1126), .O(gate480inter2));
  inv1  gate956(.a(s_58), .O(gate480inter3));
  inv1  gate957(.a(s_59), .O(gate480inter4));
  nand2 gate958(.a(gate480inter4), .b(gate480inter3), .O(gate480inter5));
  nor2  gate959(.a(gate480inter5), .b(gate480inter2), .O(gate480inter6));
  inv1  gate960(.a(G1126), .O(gate480inter7));
  inv1  gate961(.a(G1222), .O(gate480inter8));
  nand2 gate962(.a(gate480inter8), .b(gate480inter7), .O(gate480inter9));
  nand2 gate963(.a(s_59), .b(gate480inter3), .O(gate480inter10));
  nor2  gate964(.a(gate480inter10), .b(gate480inter9), .O(gate480inter11));
  nor2  gate965(.a(gate480inter11), .b(gate480inter6), .O(gate480inter12));
  nand2 gate966(.a(gate480inter12), .b(gate480inter1), .O(G1289));
nand2 gate481( .a(G32), .b(G1225), .O(G1290) );
nand2 gate482( .a(G1129), .b(G1225), .O(G1291) );

  xor2  gate687(.a(G1229), .b(G1228), .O(gate483inter0));
  nand2 gate688(.a(gate483inter0), .b(s_20), .O(gate483inter1));
  and2  gate689(.a(G1229), .b(G1228), .O(gate483inter2));
  inv1  gate690(.a(s_20), .O(gate483inter3));
  inv1  gate691(.a(s_21), .O(gate483inter4));
  nand2 gate692(.a(gate483inter4), .b(gate483inter3), .O(gate483inter5));
  nor2  gate693(.a(gate483inter5), .b(gate483inter2), .O(gate483inter6));
  inv1  gate694(.a(G1228), .O(gate483inter7));
  inv1  gate695(.a(G1229), .O(gate483inter8));
  nand2 gate696(.a(gate483inter8), .b(gate483inter7), .O(gate483inter9));
  nand2 gate697(.a(s_21), .b(gate483inter3), .O(gate483inter10));
  nor2  gate698(.a(gate483inter10), .b(gate483inter9), .O(gate483inter11));
  nor2  gate699(.a(gate483inter11), .b(gate483inter6), .O(gate483inter12));
  nand2 gate700(.a(gate483inter12), .b(gate483inter1), .O(G1292));
nand2 gate484( .a(G1230), .b(G1231), .O(G1293) );
nand2 gate485( .a(G1232), .b(G1233), .O(G1294) );
nand2 gate486( .a(G1234), .b(G1235), .O(G1295) );
nand2 gate487( .a(G1236), .b(G1237), .O(G1296) );
nand2 gate488( .a(G1238), .b(G1239), .O(G1297) );
nand2 gate489( .a(G1240), .b(G1241), .O(G1298) );
nand2 gate490( .a(G1242), .b(G1243), .O(G1299) );
nand2 gate491( .a(G1244), .b(G1245), .O(G1300) );
nand2 gate492( .a(G1246), .b(G1247), .O(G1301) );
nand2 gate493( .a(G1248), .b(G1249), .O(G1302) );
nand2 gate494( .a(G1250), .b(G1251), .O(G1303) );
nand2 gate495( .a(G1252), .b(G1253), .O(G1304) );

  xor2  gate827(.a(G1255), .b(G1254), .O(gate496inter0));
  nand2 gate828(.a(gate496inter0), .b(s_40), .O(gate496inter1));
  and2  gate829(.a(G1255), .b(G1254), .O(gate496inter2));
  inv1  gate830(.a(s_40), .O(gate496inter3));
  inv1  gate831(.a(s_41), .O(gate496inter4));
  nand2 gate832(.a(gate496inter4), .b(gate496inter3), .O(gate496inter5));
  nor2  gate833(.a(gate496inter5), .b(gate496inter2), .O(gate496inter6));
  inv1  gate834(.a(G1254), .O(gate496inter7));
  inv1  gate835(.a(G1255), .O(gate496inter8));
  nand2 gate836(.a(gate496inter8), .b(gate496inter7), .O(gate496inter9));
  nand2 gate837(.a(s_41), .b(gate496inter3), .O(gate496inter10));
  nor2  gate838(.a(gate496inter10), .b(gate496inter9), .O(gate496inter11));
  nor2  gate839(.a(gate496inter11), .b(gate496inter6), .O(gate496inter12));
  nand2 gate840(.a(gate496inter12), .b(gate496inter1), .O(G1305));
nand2 gate497( .a(G1256), .b(G1257), .O(G1306) );
nand2 gate498( .a(G1258), .b(G1259), .O(G1307) );
nand2 gate499( .a(G1260), .b(G1261), .O(G1308) );
nand2 gate500( .a(G1262), .b(G1263), .O(G1309) );
nand2 gate501( .a(G1264), .b(G1265), .O(G1310) );
nand2 gate502( .a(G1266), .b(G1267), .O(G1311) );
nand2 gate503( .a(G1268), .b(G1269), .O(G1312) );
nand2 gate504( .a(G1270), .b(G1271), .O(G1313) );
nand2 gate505( .a(G1272), .b(G1273), .O(G1314) );
nand2 gate506( .a(G1274), .b(G1275), .O(G1315) );
nand2 gate507( .a(G1276), .b(G1277), .O(G1316) );
nand2 gate508( .a(G1278), .b(G1279), .O(G1317) );
nand2 gate509( .a(G1280), .b(G1281), .O(G1318) );
nand2 gate510( .a(G1282), .b(G1283), .O(G1319) );
nand2 gate511( .a(G1284), .b(G1285), .O(G1320) );
nand2 gate512( .a(G1286), .b(G1287), .O(G1321) );
nand2 gate513( .a(G1288), .b(G1289), .O(G1322) );
nand2 gate514( .a(G1290), .b(G1291), .O(G1323) );
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule