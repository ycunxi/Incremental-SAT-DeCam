module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);

input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;//RE__PI;

input s_0,s_1;//RE__ALLOW(00,01,10,11);
input s_2,s_3;//RE__ALLOW(00,01,10,11);
input s_4,s_5;//RE__ALLOW(00,01,10,11);
input s_6,s_7;//RE__ALLOW(00,01,10,11);
input s_8,s_9;//RE__ALLOW(00,01,10,11);
input s_10,s_11;//RE__ALLOW(00,01,10,11);
input s_12,s_13;//RE__ALLOW(00,01,10,11);
input s_14,s_15;//RE__ALLOW(00,01,10,11);
input s_16,s_17;//RE__ALLOW(00,01,10,11);
input s_18,s_19;//RE__ALLOW(00,01,10,11);
input s_20,s_21;//RE__ALLOW(00,01,10,11);
input s_22,s_23;//RE__ALLOW(00,01,10,11);
input s_24,s_25;//RE__ALLOW(00,01,10,11);
input s_26,s_27;//RE__ALLOW(00,01,10,11);
input s_28,s_29;//RE__ALLOW(00,01,10,11);
input s_30,s_31;//RE__ALLOW(00,01,10,11);
input s_32,s_33;//RE__ALLOW(00,01,10,11);
input s_34,s_35;//RE__ALLOW(00,01,10,11);
input s_36,s_37;//RE__ALLOW(00,01,10,11);
input s_38,s_39;//RE__ALLOW(00,01,10,11);
input s_40,s_41;//RE__ALLOW(00,01,10,11);
input s_42,s_43;//RE__ALLOW(00,01,10,11);
input s_44,s_45;//RE__ALLOW(00,01,10,11);
input s_46,s_47;//RE__ALLOW(00,01,10,11);
input s_48,s_49;//RE__ALLOW(00,01,10,11);
input s_50,s_51;//RE__ALLOW(00,01,10,11);
input s_52,s_53;//RE__ALLOW(00,01,10,11);
input s_54,s_55;//RE__ALLOW(00,01,10,11);
input s_56,s_57;//RE__ALLOW(00,01,10,11);
input s_58,s_59;//RE__ALLOW(00,01,10,11);
input s_60,s_61;//RE__ALLOW(00,01,10,11);
input s_62,s_63;//RE__ALLOW(00,01,10,11);
input s_64,s_65;//RE__ALLOW(00,01,10,11);
input s_66,s_67;//RE__ALLOW(00,01,10,11);
input s_68,s_69;//RE__ALLOW(00,01,10,11);
input s_70,s_71;//RE__ALLOW(00,01,10,11);
input s_72,s_73;//RE__ALLOW(00,01,10,11);
input s_74,s_75;//RE__ALLOW(00,01,10,11);
input s_76,s_77;//RE__ALLOW(00,01,10,11);
input s_78,s_79;//RE__ALLOW(00,01,10,11);
input s_80,s_81;//RE__ALLOW(00,01,10,11);
input s_82,s_83;//RE__ALLOW(00,01,10,11);
input s_84,s_85;//RE__ALLOW(00,01,10,11);
input s_86,s_87;//RE__ALLOW(00,01,10,11);
input s_88,s_89;//RE__ALLOW(00,01,10,11);
input s_90,s_91;//RE__ALLOW(00,01,10,11);
input s_92,s_93;//RE__ALLOW(00,01,10,11);
input s_94,s_95;//RE__ALLOW(00,01,10,11);
input s_96,s_97;//RE__ALLOW(00,01,10,11);
input s_98,s_99;//RE__ALLOW(00,01,10,11);
input s_100,s_101;//RE__ALLOW(00,01,10,11);
input s_102,s_103;//RE__ALLOW(00,01,10,11);
input s_104,s_105;//RE__ALLOW(00,01,10,11);
input s_106,s_107;//RE__ALLOW(00,01,10,11);
input s_108,s_109;//RE__ALLOW(00,01,10,11);
input s_110,s_111;//RE__ALLOW(00,01,10,11);
input s_112,s_113;//RE__ALLOW(00,01,10,11);
input s_114,s_115;//RE__ALLOW(00,01,10,11);
input s_116,s_117;//RE__ALLOW(00,01,10,11);
input s_118,s_119;//RE__ALLOW(00,01,10,11);
input s_120,s_121;//RE__ALLOW(00,01,10,11);
input s_122,s_123;//RE__ALLOW(00,01,10,11);
input s_124,s_125;//RE__ALLOW(00,01,10,11);
input s_126,s_127;//RE__ALLOW(00,01,10,11);
input s_128,s_129;//RE__ALLOW(00,01,10,11);
input s_130,s_131;//RE__ALLOW(00,01,10,11);
input s_132,s_133;//RE__ALLOW(00,01,10,11);
input s_134,s_135;//RE__ALLOW(00,01,10,11);
input s_136,s_137;//RE__ALLOW(00,01,10,11);
input s_138,s_139;//RE__ALLOW(00,01,10,11);
input s_140,s_141;//RE__ALLOW(00,01,10,11);
input s_142,s_143;//RE__ALLOW(00,01,10,11);
input s_144,s_145;//RE__ALLOW(00,01,10,11);
input s_146,s_147;//RE__ALLOW(00,01,10,11);
input s_148,s_149;//RE__ALLOW(00,01,10,11);
input s_150,s_151;//RE__ALLOW(00,01,10,11);
input s_152,s_153;//RE__ALLOW(00,01,10,11);
input s_154,s_155;//RE__ALLOW(00,01,10,11);
input s_156,s_157;//RE__ALLOW(00,01,10,11);
input s_158,s_159;//RE__ALLOW(00,01,10,11);
input s_160,s_161;//RE__ALLOW(00,01,10,11);
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;

  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate177inter0, gate177inter1, gate177inter2, gate177inter3, gate177inter4, gate177inter5, gate177inter6, gate177inter7, gate177inter8, gate177inter9, gate177inter10, gate177inter11, gate177inter12, gate157inter0, gate157inter1, gate157inter2, gate157inter3, gate157inter4, gate157inter5, gate157inter6, gate157inter7, gate157inter8, gate157inter9, gate157inter10, gate157inter11, gate157inter12, gate34inter0, gate34inter1, gate34inter2, gate34inter3, gate34inter4, gate34inter5, gate34inter6, gate34inter7, gate34inter8, gate34inter9, gate34inter10, gate34inter11, gate34inter12, gate136inter0, gate136inter1, gate136inter2, gate136inter3, gate136inter4, gate136inter5, gate136inter6, gate136inter7, gate136inter8, gate136inter9, gate136inter10, gate136inter11, gate136inter12, gate12inter0, gate12inter1, gate12inter2, gate12inter3, gate12inter4, gate12inter5, gate12inter6, gate12inter7, gate12inter8, gate12inter9, gate12inter10, gate12inter11, gate12inter12, gate233inter0, gate233inter1, gate233inter2, gate233inter3, gate233inter4, gate233inter5, gate233inter6, gate233inter7, gate233inter8, gate233inter9, gate233inter10, gate233inter11, gate233inter12, gate475inter0, gate475inter1, gate475inter2, gate475inter3, gate475inter4, gate475inter5, gate475inter6, gate475inter7, gate475inter8, gate475inter9, gate475inter10, gate475inter11, gate475inter12, gate147inter0, gate147inter1, gate147inter2, gate147inter3, gate147inter4, gate147inter5, gate147inter6, gate147inter7, gate147inter8, gate147inter9, gate147inter10, gate147inter11, gate147inter12, gate255inter0, gate255inter1, gate255inter2, gate255inter3, gate255inter4, gate255inter5, gate255inter6, gate255inter7, gate255inter8, gate255inter9, gate255inter10, gate255inter11, gate255inter12, gate240inter0, gate240inter1, gate240inter2, gate240inter3, gate240inter4, gate240inter5, gate240inter6, gate240inter7, gate240inter8, gate240inter9, gate240inter10, gate240inter11, gate240inter12, gate121inter0, gate121inter1, gate121inter2, gate121inter3, gate121inter4, gate121inter5, gate121inter6, gate121inter7, gate121inter8, gate121inter9, gate121inter10, gate121inter11, gate121inter12, gate22inter0, gate22inter1, gate22inter2, gate22inter3, gate22inter4, gate22inter5, gate22inter6, gate22inter7, gate22inter8, gate22inter9, gate22inter10, gate22inter11, gate22inter12, gate56inter0, gate56inter1, gate56inter2, gate56inter3, gate56inter4, gate56inter5, gate56inter6, gate56inter7, gate56inter8, gate56inter9, gate56inter10, gate56inter11, gate56inter12, gate252inter0, gate252inter1, gate252inter2, gate252inter3, gate252inter4, gate252inter5, gate252inter6, gate252inter7, gate252inter8, gate252inter9, gate252inter10, gate252inter11, gate252inter12, gate478inter0, gate478inter1, gate478inter2, gate478inter3, gate478inter4, gate478inter5, gate478inter6, gate478inter7, gate478inter8, gate478inter9, gate478inter10, gate478inter11, gate478inter12, gate286inter0, gate286inter1, gate286inter2, gate286inter3, gate286inter4, gate286inter5, gate286inter6, gate286inter7, gate286inter8, gate286inter9, gate286inter10, gate286inter11, gate286inter12, gate269inter0, gate269inter1, gate269inter2, gate269inter3, gate269inter4, gate269inter5, gate269inter6, gate269inter7, gate269inter8, gate269inter9, gate269inter10, gate269inter11, gate269inter12, gate245inter0, gate245inter1, gate245inter2, gate245inter3, gate245inter4, gate245inter5, gate245inter6, gate245inter7, gate245inter8, gate245inter9, gate245inter10, gate245inter11, gate245inter12, gate450inter0, gate450inter1, gate450inter2, gate450inter3, gate450inter4, gate450inter5, gate450inter6, gate450inter7, gate450inter8, gate450inter9, gate450inter10, gate450inter11, gate450inter12, gate44inter0, gate44inter1, gate44inter2, gate44inter3, gate44inter4, gate44inter5, gate44inter6, gate44inter7, gate44inter8, gate44inter9, gate44inter10, gate44inter11, gate44inter12, gate113inter0, gate113inter1, gate113inter2, gate113inter3, gate113inter4, gate113inter5, gate113inter6, gate113inter7, gate113inter8, gate113inter9, gate113inter10, gate113inter11, gate113inter12, gate123inter0, gate123inter1, gate123inter2, gate123inter3, gate123inter4, gate123inter5, gate123inter6, gate123inter7, gate123inter8, gate123inter9, gate123inter10, gate123inter11, gate123inter12, gate247inter0, gate247inter1, gate247inter2, gate247inter3, gate247inter4, gate247inter5, gate247inter6, gate247inter7, gate247inter8, gate247inter9, gate247inter10, gate247inter11, gate247inter12, gate173inter0, gate173inter1, gate173inter2, gate173inter3, gate173inter4, gate173inter5, gate173inter6, gate173inter7, gate173inter8, gate173inter9, gate173inter10, gate173inter11, gate173inter12, gate92inter0, gate92inter1, gate92inter2, gate92inter3, gate92inter4, gate92inter5, gate92inter6, gate92inter7, gate92inter8, gate92inter9, gate92inter10, gate92inter11, gate92inter12, gate161inter0, gate161inter1, gate161inter2, gate161inter3, gate161inter4, gate161inter5, gate161inter6, gate161inter7, gate161inter8, gate161inter9, gate161inter10, gate161inter11, gate161inter12, gate486inter0, gate486inter1, gate486inter2, gate486inter3, gate486inter4, gate486inter5, gate486inter6, gate486inter7, gate486inter8, gate486inter9, gate486inter10, gate486inter11, gate486inter12, gate29inter0, gate29inter1, gate29inter2, gate29inter3, gate29inter4, gate29inter5, gate29inter6, gate29inter7, gate29inter8, gate29inter9, gate29inter10, gate29inter11, gate29inter12, gate410inter0, gate410inter1, gate410inter2, gate410inter3, gate410inter4, gate410inter5, gate410inter6, gate410inter7, gate410inter8, gate410inter9, gate410inter10, gate410inter11, gate410inter12, gate15inter0, gate15inter1, gate15inter2, gate15inter3, gate15inter4, gate15inter5, gate15inter6, gate15inter7, gate15inter8, gate15inter9, gate15inter10, gate15inter11, gate15inter12, gate429inter0, gate429inter1, gate429inter2, gate429inter3, gate429inter4, gate429inter5, gate429inter6, gate429inter7, gate429inter8, gate429inter9, gate429inter10, gate429inter11, gate429inter12, gate224inter0, gate224inter1, gate224inter2, gate224inter3, gate224inter4, gate224inter5, gate224inter6, gate224inter7, gate224inter8, gate224inter9, gate224inter10, gate224inter11, gate224inter12, gate414inter0, gate414inter1, gate414inter2, gate414inter3, gate414inter4, gate414inter5, gate414inter6, gate414inter7, gate414inter8, gate414inter9, gate414inter10, gate414inter11, gate414inter12, gate417inter0, gate417inter1, gate417inter2, gate417inter3, gate417inter4, gate417inter5, gate417inter6, gate417inter7, gate417inter8, gate417inter9, gate417inter10, gate417inter11, gate417inter12, gate39inter0, gate39inter1, gate39inter2, gate39inter3, gate39inter4, gate39inter5, gate39inter6, gate39inter7, gate39inter8, gate39inter9, gate39inter10, gate39inter11, gate39inter12, gate205inter0, gate205inter1, gate205inter2, gate205inter3, gate205inter4, gate205inter5, gate205inter6, gate205inter7, gate205inter8, gate205inter9, gate205inter10, gate205inter11, gate205inter12, gate391inter0, gate391inter1, gate391inter2, gate391inter3, gate391inter4, gate391inter5, gate391inter6, gate391inter7, gate391inter8, gate391inter9, gate391inter10, gate391inter11, gate391inter12, gate285inter0, gate285inter1, gate285inter2, gate285inter3, gate285inter4, gate285inter5, gate285inter6, gate285inter7, gate285inter8, gate285inter9, gate285inter10, gate285inter11, gate285inter12, gate287inter0, gate287inter1, gate287inter2, gate287inter3, gate287inter4, gate287inter5, gate287inter6, gate287inter7, gate287inter8, gate287inter9, gate287inter10, gate287inter11, gate287inter12, gate149inter0, gate149inter1, gate149inter2, gate149inter3, gate149inter4, gate149inter5, gate149inter6, gate149inter7, gate149inter8, gate149inter9, gate149inter10, gate149inter11, gate149inter12, gate102inter0, gate102inter1, gate102inter2, gate102inter3, gate102inter4, gate102inter5, gate102inter6, gate102inter7, gate102inter8, gate102inter9, gate102inter10, gate102inter11, gate102inter12, gate49inter0, gate49inter1, gate49inter2, gate49inter3, gate49inter4, gate49inter5, gate49inter6, gate49inter7, gate49inter8, gate49inter9, gate49inter10, gate49inter11, gate49inter12, gate186inter0, gate186inter1, gate186inter2, gate186inter3, gate186inter4, gate186inter5, gate186inter6, gate186inter7, gate186inter8, gate186inter9, gate186inter10, gate186inter11, gate186inter12, gate132inter0, gate132inter1, gate132inter2, gate132inter3, gate132inter4, gate132inter5, gate132inter6, gate132inter7, gate132inter8, gate132inter9, gate132inter10, gate132inter11, gate132inter12, gate67inter0, gate67inter1, gate67inter2, gate67inter3, gate67inter4, gate67inter5, gate67inter6, gate67inter7, gate67inter8, gate67inter9, gate67inter10, gate67inter11, gate67inter12, gate387inter0, gate387inter1, gate387inter2, gate387inter3, gate387inter4, gate387inter5, gate387inter6, gate387inter7, gate387inter8, gate387inter9, gate387inter10, gate387inter11, gate387inter12, gate24inter0, gate24inter1, gate24inter2, gate24inter3, gate24inter4, gate24inter5, gate24inter6, gate24inter7, gate24inter8, gate24inter9, gate24inter10, gate24inter11, gate24inter12, gate260inter0, gate260inter1, gate260inter2, gate260inter3, gate260inter4, gate260inter5, gate260inter6, gate260inter7, gate260inter8, gate260inter9, gate260inter10, gate260inter11, gate260inter12, gate246inter0, gate246inter1, gate246inter2, gate246inter3, gate246inter4, gate246inter5, gate246inter6, gate246inter7, gate246inter8, gate246inter9, gate246inter10, gate246inter11, gate246inter12, gate272inter0, gate272inter1, gate272inter2, gate272inter3, gate272inter4, gate272inter5, gate272inter6, gate272inter7, gate272inter8, gate272inter9, gate272inter10, gate272inter11, gate272inter12, gate459inter0, gate459inter1, gate459inter2, gate459inter3, gate459inter4, gate459inter5, gate459inter6, gate459inter7, gate459inter8, gate459inter9, gate459inter10, gate459inter11, gate459inter12, gate251inter0, gate251inter1, gate251inter2, gate251inter3, gate251inter4, gate251inter5, gate251inter6, gate251inter7, gate251inter8, gate251inter9, gate251inter10, gate251inter11, gate251inter12, gate223inter0, gate223inter1, gate223inter2, gate223inter3, gate223inter4, gate223inter5, gate223inter6, gate223inter7, gate223inter8, gate223inter9, gate223inter10, gate223inter11, gate223inter12, gate166inter0, gate166inter1, gate166inter2, gate166inter3, gate166inter4, gate166inter5, gate166inter6, gate166inter7, gate166inter8, gate166inter9, gate166inter10, gate166inter11, gate166inter12, gate17inter0, gate17inter1, gate17inter2, gate17inter3, gate17inter4, gate17inter5, gate17inter6, gate17inter7, gate17inter8, gate17inter9, gate17inter10, gate17inter11, gate17inter12, gate174inter0, gate174inter1, gate174inter2, gate174inter3, gate174inter4, gate174inter5, gate174inter6, gate174inter7, gate174inter8, gate174inter9, gate174inter10, gate174inter11, gate174inter12, gate288inter0, gate288inter1, gate288inter2, gate288inter3, gate288inter4, gate288inter5, gate288inter6, gate288inter7, gate288inter8, gate288inter9, gate288inter10, gate288inter11, gate288inter12, gate207inter0, gate207inter1, gate207inter2, gate207inter3, gate207inter4, gate207inter5, gate207inter6, gate207inter7, gate207inter8, gate207inter9, gate207inter10, gate207inter11, gate207inter12, gate86inter0, gate86inter1, gate86inter2, gate86inter3, gate86inter4, gate86inter5, gate86inter6, gate86inter7, gate86inter8, gate86inter9, gate86inter10, gate86inter11, gate86inter12, gate219inter0, gate219inter1, gate219inter2, gate219inter3, gate219inter4, gate219inter5, gate219inter6, gate219inter7, gate219inter8, gate219inter9, gate219inter10, gate219inter11, gate219inter12, gate472inter0, gate472inter1, gate472inter2, gate472inter3, gate472inter4, gate472inter5, gate472inter6, gate472inter7, gate472inter8, gate472inter9, gate472inter10, gate472inter11, gate472inter12, gate468inter0, gate468inter1, gate468inter2, gate468inter3, gate468inter4, gate468inter5, gate468inter6, gate468inter7, gate468inter8, gate468inter9, gate468inter10, gate468inter11, gate468inter12, gate226inter0, gate226inter1, gate226inter2, gate226inter3, gate226inter4, gate226inter5, gate226inter6, gate226inter7, gate226inter8, gate226inter9, gate226inter10, gate226inter11, gate226inter12, gate418inter0, gate418inter1, gate418inter2, gate418inter3, gate418inter4, gate418inter5, gate418inter6, gate418inter7, gate418inter8, gate418inter9, gate418inter10, gate418inter11, gate418inter12, gate456inter0, gate456inter1, gate456inter2, gate456inter3, gate456inter4, gate456inter5, gate456inter6, gate456inter7, gate456inter8, gate456inter9, gate456inter10, gate456inter11, gate456inter12, gate402inter0, gate402inter1, gate402inter2, gate402inter3, gate402inter4, gate402inter5, gate402inter6, gate402inter7, gate402inter8, gate402inter9, gate402inter10, gate402inter11, gate402inter12, gate203inter0, gate203inter1, gate203inter2, gate203inter3, gate203inter4, gate203inter5, gate203inter6, gate203inter7, gate203inter8, gate203inter9, gate203inter10, gate203inter11, gate203inter12, gate432inter0, gate432inter1, gate432inter2, gate432inter3, gate432inter4, gate432inter5, gate432inter6, gate432inter7, gate432inter8, gate432inter9, gate432inter10, gate432inter11, gate432inter12, gate481inter0, gate481inter1, gate481inter2, gate481inter3, gate481inter4, gate481inter5, gate481inter6, gate481inter7, gate481inter8, gate481inter9, gate481inter10, gate481inter11, gate481inter12, gate488inter0, gate488inter1, gate488inter2, gate488inter3, gate488inter4, gate488inter5, gate488inter6, gate488inter7, gate488inter8, gate488inter9, gate488inter10, gate488inter11, gate488inter12, gate51inter0, gate51inter1, gate51inter2, gate51inter3, gate51inter4, gate51inter5, gate51inter6, gate51inter7, gate51inter8, gate51inter9, gate51inter10, gate51inter11, gate51inter12, gate124inter0, gate124inter1, gate124inter2, gate124inter3, gate124inter4, gate124inter5, gate124inter6, gate124inter7, gate124inter8, gate124inter9, gate124inter10, gate124inter11, gate124inter12, gate216inter0, gate216inter1, gate216inter2, gate216inter3, gate216inter4, gate216inter5, gate216inter6, gate216inter7, gate216inter8, gate216inter9, gate216inter10, gate216inter11, gate216inter12, gate407inter0, gate407inter1, gate407inter2, gate407inter3, gate407inter4, gate407inter5, gate407inter6, gate407inter7, gate407inter8, gate407inter9, gate407inter10, gate407inter11, gate407inter12, gate159inter0, gate159inter1, gate159inter2, gate159inter3, gate159inter4, gate159inter5, gate159inter6, gate159inter7, gate159inter8, gate159inter9, gate159inter10, gate159inter11, gate159inter12, gate279inter0, gate279inter1, gate279inter2, gate279inter3, gate279inter4, gate279inter5, gate279inter6, gate279inter7, gate279inter8, gate279inter9, gate279inter10, gate279inter11, gate279inter12, gate142inter0, gate142inter1, gate142inter2, gate142inter3, gate142inter4, gate142inter5, gate142inter6, gate142inter7, gate142inter8, gate142inter9, gate142inter10, gate142inter11, gate142inter12, gate93inter0, gate93inter1, gate93inter2, gate93inter3, gate93inter4, gate93inter5, gate93inter6, gate93inter7, gate93inter8, gate93inter9, gate93inter10, gate93inter11, gate93inter12, gate235inter0, gate235inter1, gate235inter2, gate235inter3, gate235inter4, gate235inter5, gate235inter6, gate235inter7, gate235inter8, gate235inter9, gate235inter10, gate235inter11, gate235inter12, gate507inter0, gate507inter1, gate507inter2, gate507inter3, gate507inter4, gate507inter5, gate507inter6, gate507inter7, gate507inter8, gate507inter9, gate507inter10, gate507inter11, gate507inter12, gate501inter0, gate501inter1, gate501inter2, gate501inter3, gate501inter4, gate501inter5, gate501inter6, gate501inter7, gate501inter8, gate501inter9, gate501inter10, gate501inter11, gate501inter12;



and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );
nand2 gate9( .a(G1), .b(G2), .O(G266) );
nand2 gate10( .a(G3), .b(G4), .O(G269) );
nand2 gate11( .a(G5), .b(G6), .O(G272) );

  xor2  gate603(.a(G8), .b(G7), .O(gate12inter0));
  nand2 gate604(.a(gate12inter0), .b(s_8), .O(gate12inter1));
  and2  gate605(.a(G8), .b(G7), .O(gate12inter2));
  inv1  gate606(.a(s_8), .O(gate12inter3));
  inv1  gate607(.a(s_9), .O(gate12inter4));
  nand2 gate608(.a(gate12inter4), .b(gate12inter3), .O(gate12inter5));
  nor2  gate609(.a(gate12inter5), .b(gate12inter2), .O(gate12inter6));
  inv1  gate610(.a(G7), .O(gate12inter7));
  inv1  gate611(.a(G8), .O(gate12inter8));
  nand2 gate612(.a(gate12inter8), .b(gate12inter7), .O(gate12inter9));
  nand2 gate613(.a(s_9), .b(gate12inter3), .O(gate12inter10));
  nor2  gate614(.a(gate12inter10), .b(gate12inter9), .O(gate12inter11));
  nor2  gate615(.a(gate12inter11), .b(gate12inter6), .O(gate12inter12));
  nand2 gate616(.a(gate12inter12), .b(gate12inter1), .O(G275));
nand2 gate13( .a(G9), .b(G10), .O(G278) );
nand2 gate14( .a(G11), .b(G12), .O(G281) );

  xor2  gate953(.a(G14), .b(G13), .O(gate15inter0));
  nand2 gate954(.a(gate15inter0), .b(s_58), .O(gate15inter1));
  and2  gate955(.a(G14), .b(G13), .O(gate15inter2));
  inv1  gate956(.a(s_58), .O(gate15inter3));
  inv1  gate957(.a(s_59), .O(gate15inter4));
  nand2 gate958(.a(gate15inter4), .b(gate15inter3), .O(gate15inter5));
  nor2  gate959(.a(gate15inter5), .b(gate15inter2), .O(gate15inter6));
  inv1  gate960(.a(G13), .O(gate15inter7));
  inv1  gate961(.a(G14), .O(gate15inter8));
  nand2 gate962(.a(gate15inter8), .b(gate15inter7), .O(gate15inter9));
  nand2 gate963(.a(s_59), .b(gate15inter3), .O(gate15inter10));
  nor2  gate964(.a(gate15inter10), .b(gate15inter9), .O(gate15inter11));
  nor2  gate965(.a(gate15inter11), .b(gate15inter6), .O(gate15inter12));
  nand2 gate966(.a(gate15inter12), .b(gate15inter1), .O(G284));
nand2 gate16( .a(G15), .b(G16), .O(G287) );

  xor2  gate1303(.a(G18), .b(G17), .O(gate17inter0));
  nand2 gate1304(.a(gate17inter0), .b(s_108), .O(gate17inter1));
  and2  gate1305(.a(G18), .b(G17), .O(gate17inter2));
  inv1  gate1306(.a(s_108), .O(gate17inter3));
  inv1  gate1307(.a(s_109), .O(gate17inter4));
  nand2 gate1308(.a(gate17inter4), .b(gate17inter3), .O(gate17inter5));
  nor2  gate1309(.a(gate17inter5), .b(gate17inter2), .O(gate17inter6));
  inv1  gate1310(.a(G17), .O(gate17inter7));
  inv1  gate1311(.a(G18), .O(gate17inter8));
  nand2 gate1312(.a(gate17inter8), .b(gate17inter7), .O(gate17inter9));
  nand2 gate1313(.a(s_109), .b(gate17inter3), .O(gate17inter10));
  nor2  gate1314(.a(gate17inter10), .b(gate17inter9), .O(gate17inter11));
  nor2  gate1315(.a(gate17inter11), .b(gate17inter6), .O(gate17inter12));
  nand2 gate1316(.a(gate17inter12), .b(gate17inter1), .O(G290));
nand2 gate18( .a(G19), .b(G20), .O(G293) );
nand2 gate19( .a(G21), .b(G22), .O(G296) );
nand2 gate20( .a(G23), .b(G24), .O(G299) );
nand2 gate21( .a(G25), .b(G26), .O(G302) );

  xor2  gate701(.a(G28), .b(G27), .O(gate22inter0));
  nand2 gate702(.a(gate22inter0), .b(s_22), .O(gate22inter1));
  and2  gate703(.a(G28), .b(G27), .O(gate22inter2));
  inv1  gate704(.a(s_22), .O(gate22inter3));
  inv1  gate705(.a(s_23), .O(gate22inter4));
  nand2 gate706(.a(gate22inter4), .b(gate22inter3), .O(gate22inter5));
  nor2  gate707(.a(gate22inter5), .b(gate22inter2), .O(gate22inter6));
  inv1  gate708(.a(G27), .O(gate22inter7));
  inv1  gate709(.a(G28), .O(gate22inter8));
  nand2 gate710(.a(gate22inter8), .b(gate22inter7), .O(gate22inter9));
  nand2 gate711(.a(s_23), .b(gate22inter3), .O(gate22inter10));
  nor2  gate712(.a(gate22inter10), .b(gate22inter9), .O(gate22inter11));
  nor2  gate713(.a(gate22inter11), .b(gate22inter6), .O(gate22inter12));
  nand2 gate714(.a(gate22inter12), .b(gate22inter1), .O(G305));
nand2 gate23( .a(G29), .b(G30), .O(G308) );

  xor2  gate1191(.a(G32), .b(G31), .O(gate24inter0));
  nand2 gate1192(.a(gate24inter0), .b(s_92), .O(gate24inter1));
  and2  gate1193(.a(G32), .b(G31), .O(gate24inter2));
  inv1  gate1194(.a(s_92), .O(gate24inter3));
  inv1  gate1195(.a(s_93), .O(gate24inter4));
  nand2 gate1196(.a(gate24inter4), .b(gate24inter3), .O(gate24inter5));
  nor2  gate1197(.a(gate24inter5), .b(gate24inter2), .O(gate24inter6));
  inv1  gate1198(.a(G31), .O(gate24inter7));
  inv1  gate1199(.a(G32), .O(gate24inter8));
  nand2 gate1200(.a(gate24inter8), .b(gate24inter7), .O(gate24inter9));
  nand2 gate1201(.a(s_93), .b(gate24inter3), .O(gate24inter10));
  nor2  gate1202(.a(gate24inter10), .b(gate24inter9), .O(gate24inter11));
  nor2  gate1203(.a(gate24inter11), .b(gate24inter6), .O(gate24inter12));
  nand2 gate1204(.a(gate24inter12), .b(gate24inter1), .O(G311));
nand2 gate25( .a(G1), .b(G5), .O(G314) );
nand2 gate26( .a(G9), .b(G13), .O(G317) );
nand2 gate27( .a(G2), .b(G6), .O(G320) );
nand2 gate28( .a(G10), .b(G14), .O(G323) );

  xor2  gate925(.a(G7), .b(G3), .O(gate29inter0));
  nand2 gate926(.a(gate29inter0), .b(s_54), .O(gate29inter1));
  and2  gate927(.a(G7), .b(G3), .O(gate29inter2));
  inv1  gate928(.a(s_54), .O(gate29inter3));
  inv1  gate929(.a(s_55), .O(gate29inter4));
  nand2 gate930(.a(gate29inter4), .b(gate29inter3), .O(gate29inter5));
  nor2  gate931(.a(gate29inter5), .b(gate29inter2), .O(gate29inter6));
  inv1  gate932(.a(G3), .O(gate29inter7));
  inv1  gate933(.a(G7), .O(gate29inter8));
  nand2 gate934(.a(gate29inter8), .b(gate29inter7), .O(gate29inter9));
  nand2 gate935(.a(s_55), .b(gate29inter3), .O(gate29inter10));
  nor2  gate936(.a(gate29inter10), .b(gate29inter9), .O(gate29inter11));
  nor2  gate937(.a(gate29inter11), .b(gate29inter6), .O(gate29inter12));
  nand2 gate938(.a(gate29inter12), .b(gate29inter1), .O(G326));
nand2 gate30( .a(G11), .b(G15), .O(G329) );
nand2 gate31( .a(G4), .b(G8), .O(G332) );
nand2 gate32( .a(G12), .b(G16), .O(G335) );
nand2 gate33( .a(G17), .b(G21), .O(G338) );

  xor2  gate575(.a(G29), .b(G25), .O(gate34inter0));
  nand2 gate576(.a(gate34inter0), .b(s_4), .O(gate34inter1));
  and2  gate577(.a(G29), .b(G25), .O(gate34inter2));
  inv1  gate578(.a(s_4), .O(gate34inter3));
  inv1  gate579(.a(s_5), .O(gate34inter4));
  nand2 gate580(.a(gate34inter4), .b(gate34inter3), .O(gate34inter5));
  nor2  gate581(.a(gate34inter5), .b(gate34inter2), .O(gate34inter6));
  inv1  gate582(.a(G25), .O(gate34inter7));
  inv1  gate583(.a(G29), .O(gate34inter8));
  nand2 gate584(.a(gate34inter8), .b(gate34inter7), .O(gate34inter9));
  nand2 gate585(.a(s_5), .b(gate34inter3), .O(gate34inter10));
  nor2  gate586(.a(gate34inter10), .b(gate34inter9), .O(gate34inter11));
  nor2  gate587(.a(gate34inter11), .b(gate34inter6), .O(gate34inter12));
  nand2 gate588(.a(gate34inter12), .b(gate34inter1), .O(G341));
nand2 gate35( .a(G18), .b(G22), .O(G344) );
nand2 gate36( .a(G26), .b(G30), .O(G347) );
nand2 gate37( .a(G19), .b(G23), .O(G350) );
nand2 gate38( .a(G27), .b(G31), .O(G353) );

  xor2  gate1023(.a(G24), .b(G20), .O(gate39inter0));
  nand2 gate1024(.a(gate39inter0), .b(s_68), .O(gate39inter1));
  and2  gate1025(.a(G24), .b(G20), .O(gate39inter2));
  inv1  gate1026(.a(s_68), .O(gate39inter3));
  inv1  gate1027(.a(s_69), .O(gate39inter4));
  nand2 gate1028(.a(gate39inter4), .b(gate39inter3), .O(gate39inter5));
  nor2  gate1029(.a(gate39inter5), .b(gate39inter2), .O(gate39inter6));
  inv1  gate1030(.a(G20), .O(gate39inter7));
  inv1  gate1031(.a(G24), .O(gate39inter8));
  nand2 gate1032(.a(gate39inter8), .b(gate39inter7), .O(gate39inter9));
  nand2 gate1033(.a(s_69), .b(gate39inter3), .O(gate39inter10));
  nor2  gate1034(.a(gate39inter10), .b(gate39inter9), .O(gate39inter11));
  nor2  gate1035(.a(gate39inter11), .b(gate39inter6), .O(gate39inter12));
  nand2 gate1036(.a(gate39inter12), .b(gate39inter1), .O(G356));
nand2 gate40( .a(G28), .b(G32), .O(G359) );
nand2 gate41( .a(G1), .b(G266), .O(G362) );
nand2 gate42( .a(G2), .b(G266), .O(G363) );
nand2 gate43( .a(G3), .b(G269), .O(G364) );

  xor2  gate813(.a(G269), .b(G4), .O(gate44inter0));
  nand2 gate814(.a(gate44inter0), .b(s_38), .O(gate44inter1));
  and2  gate815(.a(G269), .b(G4), .O(gate44inter2));
  inv1  gate816(.a(s_38), .O(gate44inter3));
  inv1  gate817(.a(s_39), .O(gate44inter4));
  nand2 gate818(.a(gate44inter4), .b(gate44inter3), .O(gate44inter5));
  nor2  gate819(.a(gate44inter5), .b(gate44inter2), .O(gate44inter6));
  inv1  gate820(.a(G4), .O(gate44inter7));
  inv1  gate821(.a(G269), .O(gate44inter8));
  nand2 gate822(.a(gate44inter8), .b(gate44inter7), .O(gate44inter9));
  nand2 gate823(.a(s_39), .b(gate44inter3), .O(gate44inter10));
  nor2  gate824(.a(gate44inter10), .b(gate44inter9), .O(gate44inter11));
  nor2  gate825(.a(gate44inter11), .b(gate44inter6), .O(gate44inter12));
  nand2 gate826(.a(gate44inter12), .b(gate44inter1), .O(G365));
nand2 gate45( .a(G5), .b(G272), .O(G366) );
nand2 gate46( .a(G6), .b(G272), .O(G367) );
nand2 gate47( .a(G7), .b(G275), .O(G368) );
nand2 gate48( .a(G8), .b(G275), .O(G369) );

  xor2  gate1121(.a(G278), .b(G9), .O(gate49inter0));
  nand2 gate1122(.a(gate49inter0), .b(s_82), .O(gate49inter1));
  and2  gate1123(.a(G278), .b(G9), .O(gate49inter2));
  inv1  gate1124(.a(s_82), .O(gate49inter3));
  inv1  gate1125(.a(s_83), .O(gate49inter4));
  nand2 gate1126(.a(gate49inter4), .b(gate49inter3), .O(gate49inter5));
  nor2  gate1127(.a(gate49inter5), .b(gate49inter2), .O(gate49inter6));
  inv1  gate1128(.a(G9), .O(gate49inter7));
  inv1  gate1129(.a(G278), .O(gate49inter8));
  nand2 gate1130(.a(gate49inter8), .b(gate49inter7), .O(gate49inter9));
  nand2 gate1131(.a(s_83), .b(gate49inter3), .O(gate49inter10));
  nor2  gate1132(.a(gate49inter10), .b(gate49inter9), .O(gate49inter11));
  nor2  gate1133(.a(gate49inter11), .b(gate49inter6), .O(gate49inter12));
  nand2 gate1134(.a(gate49inter12), .b(gate49inter1), .O(G370));
nand2 gate50( .a(G10), .b(G278), .O(G371) );

  xor2  gate1527(.a(G281), .b(G11), .O(gate51inter0));
  nand2 gate1528(.a(gate51inter0), .b(s_140), .O(gate51inter1));
  and2  gate1529(.a(G281), .b(G11), .O(gate51inter2));
  inv1  gate1530(.a(s_140), .O(gate51inter3));
  inv1  gate1531(.a(s_141), .O(gate51inter4));
  nand2 gate1532(.a(gate51inter4), .b(gate51inter3), .O(gate51inter5));
  nor2  gate1533(.a(gate51inter5), .b(gate51inter2), .O(gate51inter6));
  inv1  gate1534(.a(G11), .O(gate51inter7));
  inv1  gate1535(.a(G281), .O(gate51inter8));
  nand2 gate1536(.a(gate51inter8), .b(gate51inter7), .O(gate51inter9));
  nand2 gate1537(.a(s_141), .b(gate51inter3), .O(gate51inter10));
  nor2  gate1538(.a(gate51inter10), .b(gate51inter9), .O(gate51inter11));
  nor2  gate1539(.a(gate51inter11), .b(gate51inter6), .O(gate51inter12));
  nand2 gate1540(.a(gate51inter12), .b(gate51inter1), .O(G372));
nand2 gate52( .a(G12), .b(G281), .O(G373) );
nand2 gate53( .a(G13), .b(G284), .O(G374) );
nand2 gate54( .a(G14), .b(G284), .O(G375) );
nand2 gate55( .a(G15), .b(G287), .O(G376) );

  xor2  gate715(.a(G287), .b(G16), .O(gate56inter0));
  nand2 gate716(.a(gate56inter0), .b(s_24), .O(gate56inter1));
  and2  gate717(.a(G287), .b(G16), .O(gate56inter2));
  inv1  gate718(.a(s_24), .O(gate56inter3));
  inv1  gate719(.a(s_25), .O(gate56inter4));
  nand2 gate720(.a(gate56inter4), .b(gate56inter3), .O(gate56inter5));
  nor2  gate721(.a(gate56inter5), .b(gate56inter2), .O(gate56inter6));
  inv1  gate722(.a(G16), .O(gate56inter7));
  inv1  gate723(.a(G287), .O(gate56inter8));
  nand2 gate724(.a(gate56inter8), .b(gate56inter7), .O(gate56inter9));
  nand2 gate725(.a(s_25), .b(gate56inter3), .O(gate56inter10));
  nor2  gate726(.a(gate56inter10), .b(gate56inter9), .O(gate56inter11));
  nor2  gate727(.a(gate56inter11), .b(gate56inter6), .O(gate56inter12));
  nand2 gate728(.a(gate56inter12), .b(gate56inter1), .O(G377));
nand2 gate57( .a(G17), .b(G290), .O(G378) );
nand2 gate58( .a(G18), .b(G290), .O(G379) );
nand2 gate59( .a(G19), .b(G293), .O(G380) );
nand2 gate60( .a(G20), .b(G293), .O(G381) );
nand2 gate61( .a(G21), .b(G296), .O(G382) );
nand2 gate62( .a(G22), .b(G296), .O(G383) );
nand2 gate63( .a(G23), .b(G299), .O(G384) );
nand2 gate64( .a(G24), .b(G299), .O(G385) );
nand2 gate65( .a(G25), .b(G302), .O(G386) );
nand2 gate66( .a(G26), .b(G302), .O(G387) );

  xor2  gate1163(.a(G305), .b(G27), .O(gate67inter0));
  nand2 gate1164(.a(gate67inter0), .b(s_88), .O(gate67inter1));
  and2  gate1165(.a(G305), .b(G27), .O(gate67inter2));
  inv1  gate1166(.a(s_88), .O(gate67inter3));
  inv1  gate1167(.a(s_89), .O(gate67inter4));
  nand2 gate1168(.a(gate67inter4), .b(gate67inter3), .O(gate67inter5));
  nor2  gate1169(.a(gate67inter5), .b(gate67inter2), .O(gate67inter6));
  inv1  gate1170(.a(G27), .O(gate67inter7));
  inv1  gate1171(.a(G305), .O(gate67inter8));
  nand2 gate1172(.a(gate67inter8), .b(gate67inter7), .O(gate67inter9));
  nand2 gate1173(.a(s_89), .b(gate67inter3), .O(gate67inter10));
  nor2  gate1174(.a(gate67inter10), .b(gate67inter9), .O(gate67inter11));
  nor2  gate1175(.a(gate67inter11), .b(gate67inter6), .O(gate67inter12));
  nand2 gate1176(.a(gate67inter12), .b(gate67inter1), .O(G388));
nand2 gate68( .a(G28), .b(G305), .O(G389) );
nand2 gate69( .a(G29), .b(G308), .O(G390) );
nand2 gate70( .a(G30), .b(G308), .O(G391) );
nand2 gate71( .a(G31), .b(G311), .O(G392) );
nand2 gate72( .a(G32), .b(G311), .O(G393) );
nand2 gate73( .a(G1), .b(G314), .O(G394) );
nand2 gate74( .a(G5), .b(G314), .O(G395) );
nand2 gate75( .a(G9), .b(G317), .O(G396) );
nand2 gate76( .a(G13), .b(G317), .O(G397) );
nand2 gate77( .a(G2), .b(G320), .O(G398) );
nand2 gate78( .a(G6), .b(G320), .O(G399) );
nand2 gate79( .a(G10), .b(G323), .O(G400) );
nand2 gate80( .a(G14), .b(G323), .O(G401) );
nand2 gate81( .a(G3), .b(G326), .O(G402) );
nand2 gate82( .a(G7), .b(G326), .O(G403) );
nand2 gate83( .a(G11), .b(G329), .O(G404) );
nand2 gate84( .a(G15), .b(G329), .O(G405) );
nand2 gate85( .a(G4), .b(G332), .O(G406) );

  xor2  gate1359(.a(G332), .b(G8), .O(gate86inter0));
  nand2 gate1360(.a(gate86inter0), .b(s_116), .O(gate86inter1));
  and2  gate1361(.a(G332), .b(G8), .O(gate86inter2));
  inv1  gate1362(.a(s_116), .O(gate86inter3));
  inv1  gate1363(.a(s_117), .O(gate86inter4));
  nand2 gate1364(.a(gate86inter4), .b(gate86inter3), .O(gate86inter5));
  nor2  gate1365(.a(gate86inter5), .b(gate86inter2), .O(gate86inter6));
  inv1  gate1366(.a(G8), .O(gate86inter7));
  inv1  gate1367(.a(G332), .O(gate86inter8));
  nand2 gate1368(.a(gate86inter8), .b(gate86inter7), .O(gate86inter9));
  nand2 gate1369(.a(s_117), .b(gate86inter3), .O(gate86inter10));
  nor2  gate1370(.a(gate86inter10), .b(gate86inter9), .O(gate86inter11));
  nor2  gate1371(.a(gate86inter11), .b(gate86inter6), .O(gate86inter12));
  nand2 gate1372(.a(gate86inter12), .b(gate86inter1), .O(G407));
nand2 gate87( .a(G12), .b(G335), .O(G408) );
nand2 gate88( .a(G16), .b(G335), .O(G409) );
nand2 gate89( .a(G17), .b(G338), .O(G410) );
nand2 gate90( .a(G21), .b(G338), .O(G411) );
nand2 gate91( .a(G25), .b(G341), .O(G412) );

  xor2  gate883(.a(G341), .b(G29), .O(gate92inter0));
  nand2 gate884(.a(gate92inter0), .b(s_48), .O(gate92inter1));
  and2  gate885(.a(G341), .b(G29), .O(gate92inter2));
  inv1  gate886(.a(s_48), .O(gate92inter3));
  inv1  gate887(.a(s_49), .O(gate92inter4));
  nand2 gate888(.a(gate92inter4), .b(gate92inter3), .O(gate92inter5));
  nor2  gate889(.a(gate92inter5), .b(gate92inter2), .O(gate92inter6));
  inv1  gate890(.a(G29), .O(gate92inter7));
  inv1  gate891(.a(G341), .O(gate92inter8));
  nand2 gate892(.a(gate92inter8), .b(gate92inter7), .O(gate92inter9));
  nand2 gate893(.a(s_49), .b(gate92inter3), .O(gate92inter10));
  nor2  gate894(.a(gate92inter10), .b(gate92inter9), .O(gate92inter11));
  nor2  gate895(.a(gate92inter11), .b(gate92inter6), .O(gate92inter12));
  nand2 gate896(.a(gate92inter12), .b(gate92inter1), .O(G413));

  xor2  gate1625(.a(G344), .b(G18), .O(gate93inter0));
  nand2 gate1626(.a(gate93inter0), .b(s_154), .O(gate93inter1));
  and2  gate1627(.a(G344), .b(G18), .O(gate93inter2));
  inv1  gate1628(.a(s_154), .O(gate93inter3));
  inv1  gate1629(.a(s_155), .O(gate93inter4));
  nand2 gate1630(.a(gate93inter4), .b(gate93inter3), .O(gate93inter5));
  nor2  gate1631(.a(gate93inter5), .b(gate93inter2), .O(gate93inter6));
  inv1  gate1632(.a(G18), .O(gate93inter7));
  inv1  gate1633(.a(G344), .O(gate93inter8));
  nand2 gate1634(.a(gate93inter8), .b(gate93inter7), .O(gate93inter9));
  nand2 gate1635(.a(s_155), .b(gate93inter3), .O(gate93inter10));
  nor2  gate1636(.a(gate93inter10), .b(gate93inter9), .O(gate93inter11));
  nor2  gate1637(.a(gate93inter11), .b(gate93inter6), .O(gate93inter12));
  nand2 gate1638(.a(gate93inter12), .b(gate93inter1), .O(G414));
nand2 gate94( .a(G22), .b(G344), .O(G415) );
nand2 gate95( .a(G26), .b(G347), .O(G416) );
nand2 gate96( .a(G30), .b(G347), .O(G417) );
nand2 gate97( .a(G19), .b(G350), .O(G418) );
nand2 gate98( .a(G23), .b(G350), .O(G419) );
nand2 gate99( .a(G27), .b(G353), .O(G420) );
nand2 gate100( .a(G31), .b(G353), .O(G421) );
nand2 gate101( .a(G20), .b(G356), .O(G422) );

  xor2  gate1107(.a(G356), .b(G24), .O(gate102inter0));
  nand2 gate1108(.a(gate102inter0), .b(s_80), .O(gate102inter1));
  and2  gate1109(.a(G356), .b(G24), .O(gate102inter2));
  inv1  gate1110(.a(s_80), .O(gate102inter3));
  inv1  gate1111(.a(s_81), .O(gate102inter4));
  nand2 gate1112(.a(gate102inter4), .b(gate102inter3), .O(gate102inter5));
  nor2  gate1113(.a(gate102inter5), .b(gate102inter2), .O(gate102inter6));
  inv1  gate1114(.a(G24), .O(gate102inter7));
  inv1  gate1115(.a(G356), .O(gate102inter8));
  nand2 gate1116(.a(gate102inter8), .b(gate102inter7), .O(gate102inter9));
  nand2 gate1117(.a(s_81), .b(gate102inter3), .O(gate102inter10));
  nor2  gate1118(.a(gate102inter10), .b(gate102inter9), .O(gate102inter11));
  nor2  gate1119(.a(gate102inter11), .b(gate102inter6), .O(gate102inter12));
  nand2 gate1120(.a(gate102inter12), .b(gate102inter1), .O(G423));
nand2 gate103( .a(G28), .b(G359), .O(G424) );
nand2 gate104( .a(G32), .b(G359), .O(G425) );
nand2 gate105( .a(G362), .b(G363), .O(G426) );
nand2 gate106( .a(G364), .b(G365), .O(G429) );
nand2 gate107( .a(G366), .b(G367), .O(G432) );
nand2 gate108( .a(G368), .b(G369), .O(G435) );
nand2 gate109( .a(G370), .b(G371), .O(G438) );
nand2 gate110( .a(G372), .b(G373), .O(G441) );
nand2 gate111( .a(G374), .b(G375), .O(G444) );
nand2 gate112( .a(G376), .b(G377), .O(G447) );

  xor2  gate827(.a(G379), .b(G378), .O(gate113inter0));
  nand2 gate828(.a(gate113inter0), .b(s_40), .O(gate113inter1));
  and2  gate829(.a(G379), .b(G378), .O(gate113inter2));
  inv1  gate830(.a(s_40), .O(gate113inter3));
  inv1  gate831(.a(s_41), .O(gate113inter4));
  nand2 gate832(.a(gate113inter4), .b(gate113inter3), .O(gate113inter5));
  nor2  gate833(.a(gate113inter5), .b(gate113inter2), .O(gate113inter6));
  inv1  gate834(.a(G378), .O(gate113inter7));
  inv1  gate835(.a(G379), .O(gate113inter8));
  nand2 gate836(.a(gate113inter8), .b(gate113inter7), .O(gate113inter9));
  nand2 gate837(.a(s_41), .b(gate113inter3), .O(gate113inter10));
  nor2  gate838(.a(gate113inter10), .b(gate113inter9), .O(gate113inter11));
  nor2  gate839(.a(gate113inter11), .b(gate113inter6), .O(gate113inter12));
  nand2 gate840(.a(gate113inter12), .b(gate113inter1), .O(G450));
nand2 gate114( .a(G380), .b(G381), .O(G453) );
nand2 gate115( .a(G382), .b(G383), .O(G456) );
nand2 gate116( .a(G384), .b(G385), .O(G459) );
nand2 gate117( .a(G386), .b(G387), .O(G462) );
nand2 gate118( .a(G388), .b(G389), .O(G465) );
nand2 gate119( .a(G390), .b(G391), .O(G468) );
nand2 gate120( .a(G392), .b(G393), .O(G471) );

  xor2  gate687(.a(G395), .b(G394), .O(gate121inter0));
  nand2 gate688(.a(gate121inter0), .b(s_20), .O(gate121inter1));
  and2  gate689(.a(G395), .b(G394), .O(gate121inter2));
  inv1  gate690(.a(s_20), .O(gate121inter3));
  inv1  gate691(.a(s_21), .O(gate121inter4));
  nand2 gate692(.a(gate121inter4), .b(gate121inter3), .O(gate121inter5));
  nor2  gate693(.a(gate121inter5), .b(gate121inter2), .O(gate121inter6));
  inv1  gate694(.a(G394), .O(gate121inter7));
  inv1  gate695(.a(G395), .O(gate121inter8));
  nand2 gate696(.a(gate121inter8), .b(gate121inter7), .O(gate121inter9));
  nand2 gate697(.a(s_21), .b(gate121inter3), .O(gate121inter10));
  nor2  gate698(.a(gate121inter10), .b(gate121inter9), .O(gate121inter11));
  nor2  gate699(.a(gate121inter11), .b(gate121inter6), .O(gate121inter12));
  nand2 gate700(.a(gate121inter12), .b(gate121inter1), .O(G474));
nand2 gate122( .a(G396), .b(G397), .O(G477) );

  xor2  gate841(.a(G399), .b(G398), .O(gate123inter0));
  nand2 gate842(.a(gate123inter0), .b(s_42), .O(gate123inter1));
  and2  gate843(.a(G399), .b(G398), .O(gate123inter2));
  inv1  gate844(.a(s_42), .O(gate123inter3));
  inv1  gate845(.a(s_43), .O(gate123inter4));
  nand2 gate846(.a(gate123inter4), .b(gate123inter3), .O(gate123inter5));
  nor2  gate847(.a(gate123inter5), .b(gate123inter2), .O(gate123inter6));
  inv1  gate848(.a(G398), .O(gate123inter7));
  inv1  gate849(.a(G399), .O(gate123inter8));
  nand2 gate850(.a(gate123inter8), .b(gate123inter7), .O(gate123inter9));
  nand2 gate851(.a(s_43), .b(gate123inter3), .O(gate123inter10));
  nor2  gate852(.a(gate123inter10), .b(gate123inter9), .O(gate123inter11));
  nor2  gate853(.a(gate123inter11), .b(gate123inter6), .O(gate123inter12));
  nand2 gate854(.a(gate123inter12), .b(gate123inter1), .O(G480));

  xor2  gate1541(.a(G401), .b(G400), .O(gate124inter0));
  nand2 gate1542(.a(gate124inter0), .b(s_142), .O(gate124inter1));
  and2  gate1543(.a(G401), .b(G400), .O(gate124inter2));
  inv1  gate1544(.a(s_142), .O(gate124inter3));
  inv1  gate1545(.a(s_143), .O(gate124inter4));
  nand2 gate1546(.a(gate124inter4), .b(gate124inter3), .O(gate124inter5));
  nor2  gate1547(.a(gate124inter5), .b(gate124inter2), .O(gate124inter6));
  inv1  gate1548(.a(G400), .O(gate124inter7));
  inv1  gate1549(.a(G401), .O(gate124inter8));
  nand2 gate1550(.a(gate124inter8), .b(gate124inter7), .O(gate124inter9));
  nand2 gate1551(.a(s_143), .b(gate124inter3), .O(gate124inter10));
  nor2  gate1552(.a(gate124inter10), .b(gate124inter9), .O(gate124inter11));
  nor2  gate1553(.a(gate124inter11), .b(gate124inter6), .O(gate124inter12));
  nand2 gate1554(.a(gate124inter12), .b(gate124inter1), .O(G483));
nand2 gate125( .a(G402), .b(G403), .O(G486) );
nand2 gate126( .a(G404), .b(G405), .O(G489) );
nand2 gate127( .a(G406), .b(G407), .O(G492) );
nand2 gate128( .a(G408), .b(G409), .O(G495) );
nand2 gate129( .a(G410), .b(G411), .O(G498) );
nand2 gate130( .a(G412), .b(G413), .O(G501) );
nand2 gate131( .a(G414), .b(G415), .O(G504) );

  xor2  gate1149(.a(G417), .b(G416), .O(gate132inter0));
  nand2 gate1150(.a(gate132inter0), .b(s_86), .O(gate132inter1));
  and2  gate1151(.a(G417), .b(G416), .O(gate132inter2));
  inv1  gate1152(.a(s_86), .O(gate132inter3));
  inv1  gate1153(.a(s_87), .O(gate132inter4));
  nand2 gate1154(.a(gate132inter4), .b(gate132inter3), .O(gate132inter5));
  nor2  gate1155(.a(gate132inter5), .b(gate132inter2), .O(gate132inter6));
  inv1  gate1156(.a(G416), .O(gate132inter7));
  inv1  gate1157(.a(G417), .O(gate132inter8));
  nand2 gate1158(.a(gate132inter8), .b(gate132inter7), .O(gate132inter9));
  nand2 gate1159(.a(s_87), .b(gate132inter3), .O(gate132inter10));
  nor2  gate1160(.a(gate132inter10), .b(gate132inter9), .O(gate132inter11));
  nor2  gate1161(.a(gate132inter11), .b(gate132inter6), .O(gate132inter12));
  nand2 gate1162(.a(gate132inter12), .b(gate132inter1), .O(G507));
nand2 gate133( .a(G418), .b(G419), .O(G510) );
nand2 gate134( .a(G420), .b(G421), .O(G513) );
nand2 gate135( .a(G422), .b(G423), .O(G516) );

  xor2  gate589(.a(G425), .b(G424), .O(gate136inter0));
  nand2 gate590(.a(gate136inter0), .b(s_6), .O(gate136inter1));
  and2  gate591(.a(G425), .b(G424), .O(gate136inter2));
  inv1  gate592(.a(s_6), .O(gate136inter3));
  inv1  gate593(.a(s_7), .O(gate136inter4));
  nand2 gate594(.a(gate136inter4), .b(gate136inter3), .O(gate136inter5));
  nor2  gate595(.a(gate136inter5), .b(gate136inter2), .O(gate136inter6));
  inv1  gate596(.a(G424), .O(gate136inter7));
  inv1  gate597(.a(G425), .O(gate136inter8));
  nand2 gate598(.a(gate136inter8), .b(gate136inter7), .O(gate136inter9));
  nand2 gate599(.a(s_7), .b(gate136inter3), .O(gate136inter10));
  nor2  gate600(.a(gate136inter10), .b(gate136inter9), .O(gate136inter11));
  nor2  gate601(.a(gate136inter11), .b(gate136inter6), .O(gate136inter12));
  nand2 gate602(.a(gate136inter12), .b(gate136inter1), .O(G519));
nand2 gate137( .a(G426), .b(G429), .O(G522) );
nand2 gate138( .a(G432), .b(G435), .O(G525) );
nand2 gate139( .a(G438), .b(G441), .O(G528) );
nand2 gate140( .a(G444), .b(G447), .O(G531) );
nand2 gate141( .a(G450), .b(G453), .O(G534) );

  xor2  gate1611(.a(G459), .b(G456), .O(gate142inter0));
  nand2 gate1612(.a(gate142inter0), .b(s_152), .O(gate142inter1));
  and2  gate1613(.a(G459), .b(G456), .O(gate142inter2));
  inv1  gate1614(.a(s_152), .O(gate142inter3));
  inv1  gate1615(.a(s_153), .O(gate142inter4));
  nand2 gate1616(.a(gate142inter4), .b(gate142inter3), .O(gate142inter5));
  nor2  gate1617(.a(gate142inter5), .b(gate142inter2), .O(gate142inter6));
  inv1  gate1618(.a(G456), .O(gate142inter7));
  inv1  gate1619(.a(G459), .O(gate142inter8));
  nand2 gate1620(.a(gate142inter8), .b(gate142inter7), .O(gate142inter9));
  nand2 gate1621(.a(s_153), .b(gate142inter3), .O(gate142inter10));
  nor2  gate1622(.a(gate142inter10), .b(gate142inter9), .O(gate142inter11));
  nor2  gate1623(.a(gate142inter11), .b(gate142inter6), .O(gate142inter12));
  nand2 gate1624(.a(gate142inter12), .b(gate142inter1), .O(G537));
nand2 gate143( .a(G462), .b(G465), .O(G540) );
nand2 gate144( .a(G468), .b(G471), .O(G543) );
nand2 gate145( .a(G474), .b(G477), .O(G546) );
nand2 gate146( .a(G480), .b(G483), .O(G549) );

  xor2  gate645(.a(G489), .b(G486), .O(gate147inter0));
  nand2 gate646(.a(gate147inter0), .b(s_14), .O(gate147inter1));
  and2  gate647(.a(G489), .b(G486), .O(gate147inter2));
  inv1  gate648(.a(s_14), .O(gate147inter3));
  inv1  gate649(.a(s_15), .O(gate147inter4));
  nand2 gate650(.a(gate147inter4), .b(gate147inter3), .O(gate147inter5));
  nor2  gate651(.a(gate147inter5), .b(gate147inter2), .O(gate147inter6));
  inv1  gate652(.a(G486), .O(gate147inter7));
  inv1  gate653(.a(G489), .O(gate147inter8));
  nand2 gate654(.a(gate147inter8), .b(gate147inter7), .O(gate147inter9));
  nand2 gate655(.a(s_15), .b(gate147inter3), .O(gate147inter10));
  nor2  gate656(.a(gate147inter10), .b(gate147inter9), .O(gate147inter11));
  nor2  gate657(.a(gate147inter11), .b(gate147inter6), .O(gate147inter12));
  nand2 gate658(.a(gate147inter12), .b(gate147inter1), .O(G552));
nand2 gate148( .a(G492), .b(G495), .O(G555) );

  xor2  gate1093(.a(G501), .b(G498), .O(gate149inter0));
  nand2 gate1094(.a(gate149inter0), .b(s_78), .O(gate149inter1));
  and2  gate1095(.a(G501), .b(G498), .O(gate149inter2));
  inv1  gate1096(.a(s_78), .O(gate149inter3));
  inv1  gate1097(.a(s_79), .O(gate149inter4));
  nand2 gate1098(.a(gate149inter4), .b(gate149inter3), .O(gate149inter5));
  nor2  gate1099(.a(gate149inter5), .b(gate149inter2), .O(gate149inter6));
  inv1  gate1100(.a(G498), .O(gate149inter7));
  inv1  gate1101(.a(G501), .O(gate149inter8));
  nand2 gate1102(.a(gate149inter8), .b(gate149inter7), .O(gate149inter9));
  nand2 gate1103(.a(s_79), .b(gate149inter3), .O(gate149inter10));
  nor2  gate1104(.a(gate149inter10), .b(gate149inter9), .O(gate149inter11));
  nor2  gate1105(.a(gate149inter11), .b(gate149inter6), .O(gate149inter12));
  nand2 gate1106(.a(gate149inter12), .b(gate149inter1), .O(G558));
nand2 gate150( .a(G504), .b(G507), .O(G561) );
nand2 gate151( .a(G510), .b(G513), .O(G564) );
nand2 gate152( .a(G516), .b(G519), .O(G567) );
nand2 gate153( .a(G426), .b(G522), .O(G570) );
nand2 gate154( .a(G429), .b(G522), .O(G571) );
nand2 gate155( .a(G432), .b(G525), .O(G572) );
nand2 gate156( .a(G435), .b(G525), .O(G573) );

  xor2  gate561(.a(G528), .b(G438), .O(gate157inter0));
  nand2 gate562(.a(gate157inter0), .b(s_2), .O(gate157inter1));
  and2  gate563(.a(G528), .b(G438), .O(gate157inter2));
  inv1  gate564(.a(s_2), .O(gate157inter3));
  inv1  gate565(.a(s_3), .O(gate157inter4));
  nand2 gate566(.a(gate157inter4), .b(gate157inter3), .O(gate157inter5));
  nor2  gate567(.a(gate157inter5), .b(gate157inter2), .O(gate157inter6));
  inv1  gate568(.a(G438), .O(gate157inter7));
  inv1  gate569(.a(G528), .O(gate157inter8));
  nand2 gate570(.a(gate157inter8), .b(gate157inter7), .O(gate157inter9));
  nand2 gate571(.a(s_3), .b(gate157inter3), .O(gate157inter10));
  nor2  gate572(.a(gate157inter10), .b(gate157inter9), .O(gate157inter11));
  nor2  gate573(.a(gate157inter11), .b(gate157inter6), .O(gate157inter12));
  nand2 gate574(.a(gate157inter12), .b(gate157inter1), .O(G574));
nand2 gate158( .a(G441), .b(G528), .O(G575) );

  xor2  gate1583(.a(G531), .b(G444), .O(gate159inter0));
  nand2 gate1584(.a(gate159inter0), .b(s_148), .O(gate159inter1));
  and2  gate1585(.a(G531), .b(G444), .O(gate159inter2));
  inv1  gate1586(.a(s_148), .O(gate159inter3));
  inv1  gate1587(.a(s_149), .O(gate159inter4));
  nand2 gate1588(.a(gate159inter4), .b(gate159inter3), .O(gate159inter5));
  nor2  gate1589(.a(gate159inter5), .b(gate159inter2), .O(gate159inter6));
  inv1  gate1590(.a(G444), .O(gate159inter7));
  inv1  gate1591(.a(G531), .O(gate159inter8));
  nand2 gate1592(.a(gate159inter8), .b(gate159inter7), .O(gate159inter9));
  nand2 gate1593(.a(s_149), .b(gate159inter3), .O(gate159inter10));
  nor2  gate1594(.a(gate159inter10), .b(gate159inter9), .O(gate159inter11));
  nor2  gate1595(.a(gate159inter11), .b(gate159inter6), .O(gate159inter12));
  nand2 gate1596(.a(gate159inter12), .b(gate159inter1), .O(G576));
nand2 gate160( .a(G447), .b(G531), .O(G577) );

  xor2  gate897(.a(G534), .b(G450), .O(gate161inter0));
  nand2 gate898(.a(gate161inter0), .b(s_50), .O(gate161inter1));
  and2  gate899(.a(G534), .b(G450), .O(gate161inter2));
  inv1  gate900(.a(s_50), .O(gate161inter3));
  inv1  gate901(.a(s_51), .O(gate161inter4));
  nand2 gate902(.a(gate161inter4), .b(gate161inter3), .O(gate161inter5));
  nor2  gate903(.a(gate161inter5), .b(gate161inter2), .O(gate161inter6));
  inv1  gate904(.a(G450), .O(gate161inter7));
  inv1  gate905(.a(G534), .O(gate161inter8));
  nand2 gate906(.a(gate161inter8), .b(gate161inter7), .O(gate161inter9));
  nand2 gate907(.a(s_51), .b(gate161inter3), .O(gate161inter10));
  nor2  gate908(.a(gate161inter10), .b(gate161inter9), .O(gate161inter11));
  nor2  gate909(.a(gate161inter11), .b(gate161inter6), .O(gate161inter12));
  nand2 gate910(.a(gate161inter12), .b(gate161inter1), .O(G578));
nand2 gate162( .a(G453), .b(G534), .O(G579) );
nand2 gate163( .a(G456), .b(G537), .O(G580) );
nand2 gate164( .a(G459), .b(G537), .O(G581) );
nand2 gate165( .a(G462), .b(G540), .O(G582) );

  xor2  gate1289(.a(G540), .b(G465), .O(gate166inter0));
  nand2 gate1290(.a(gate166inter0), .b(s_106), .O(gate166inter1));
  and2  gate1291(.a(G540), .b(G465), .O(gate166inter2));
  inv1  gate1292(.a(s_106), .O(gate166inter3));
  inv1  gate1293(.a(s_107), .O(gate166inter4));
  nand2 gate1294(.a(gate166inter4), .b(gate166inter3), .O(gate166inter5));
  nor2  gate1295(.a(gate166inter5), .b(gate166inter2), .O(gate166inter6));
  inv1  gate1296(.a(G465), .O(gate166inter7));
  inv1  gate1297(.a(G540), .O(gate166inter8));
  nand2 gate1298(.a(gate166inter8), .b(gate166inter7), .O(gate166inter9));
  nand2 gate1299(.a(s_107), .b(gate166inter3), .O(gate166inter10));
  nor2  gate1300(.a(gate166inter10), .b(gate166inter9), .O(gate166inter11));
  nor2  gate1301(.a(gate166inter11), .b(gate166inter6), .O(gate166inter12));
  nand2 gate1302(.a(gate166inter12), .b(gate166inter1), .O(G583));
nand2 gate167( .a(G468), .b(G543), .O(G584) );
nand2 gate168( .a(G471), .b(G543), .O(G585) );
nand2 gate169( .a(G474), .b(G546), .O(G586) );
nand2 gate170( .a(G477), .b(G546), .O(G587) );
nand2 gate171( .a(G480), .b(G549), .O(G588) );
nand2 gate172( .a(G483), .b(G549), .O(G589) );

  xor2  gate869(.a(G552), .b(G486), .O(gate173inter0));
  nand2 gate870(.a(gate173inter0), .b(s_46), .O(gate173inter1));
  and2  gate871(.a(G552), .b(G486), .O(gate173inter2));
  inv1  gate872(.a(s_46), .O(gate173inter3));
  inv1  gate873(.a(s_47), .O(gate173inter4));
  nand2 gate874(.a(gate173inter4), .b(gate173inter3), .O(gate173inter5));
  nor2  gate875(.a(gate173inter5), .b(gate173inter2), .O(gate173inter6));
  inv1  gate876(.a(G486), .O(gate173inter7));
  inv1  gate877(.a(G552), .O(gate173inter8));
  nand2 gate878(.a(gate173inter8), .b(gate173inter7), .O(gate173inter9));
  nand2 gate879(.a(s_47), .b(gate173inter3), .O(gate173inter10));
  nor2  gate880(.a(gate173inter10), .b(gate173inter9), .O(gate173inter11));
  nor2  gate881(.a(gate173inter11), .b(gate173inter6), .O(gate173inter12));
  nand2 gate882(.a(gate173inter12), .b(gate173inter1), .O(G590));

  xor2  gate1317(.a(G552), .b(G489), .O(gate174inter0));
  nand2 gate1318(.a(gate174inter0), .b(s_110), .O(gate174inter1));
  and2  gate1319(.a(G552), .b(G489), .O(gate174inter2));
  inv1  gate1320(.a(s_110), .O(gate174inter3));
  inv1  gate1321(.a(s_111), .O(gate174inter4));
  nand2 gate1322(.a(gate174inter4), .b(gate174inter3), .O(gate174inter5));
  nor2  gate1323(.a(gate174inter5), .b(gate174inter2), .O(gate174inter6));
  inv1  gate1324(.a(G489), .O(gate174inter7));
  inv1  gate1325(.a(G552), .O(gate174inter8));
  nand2 gate1326(.a(gate174inter8), .b(gate174inter7), .O(gate174inter9));
  nand2 gate1327(.a(s_111), .b(gate174inter3), .O(gate174inter10));
  nor2  gate1328(.a(gate174inter10), .b(gate174inter9), .O(gate174inter11));
  nor2  gate1329(.a(gate174inter11), .b(gate174inter6), .O(gate174inter12));
  nand2 gate1330(.a(gate174inter12), .b(gate174inter1), .O(G591));
nand2 gate175( .a(G492), .b(G555), .O(G592) );
nand2 gate176( .a(G495), .b(G555), .O(G593) );

  xor2  gate547(.a(G558), .b(G498), .O(gate177inter0));
  nand2 gate548(.a(gate177inter0), .b(s_0), .O(gate177inter1));
  and2  gate549(.a(G558), .b(G498), .O(gate177inter2));
  inv1  gate550(.a(s_0), .O(gate177inter3));
  inv1  gate551(.a(s_1), .O(gate177inter4));
  nand2 gate552(.a(gate177inter4), .b(gate177inter3), .O(gate177inter5));
  nor2  gate553(.a(gate177inter5), .b(gate177inter2), .O(gate177inter6));
  inv1  gate554(.a(G498), .O(gate177inter7));
  inv1  gate555(.a(G558), .O(gate177inter8));
  nand2 gate556(.a(gate177inter8), .b(gate177inter7), .O(gate177inter9));
  nand2 gate557(.a(s_1), .b(gate177inter3), .O(gate177inter10));
  nor2  gate558(.a(gate177inter10), .b(gate177inter9), .O(gate177inter11));
  nor2  gate559(.a(gate177inter11), .b(gate177inter6), .O(gate177inter12));
  nand2 gate560(.a(gate177inter12), .b(gate177inter1), .O(G594));
nand2 gate178( .a(G501), .b(G558), .O(G595) );
nand2 gate179( .a(G504), .b(G561), .O(G596) );
nand2 gate180( .a(G507), .b(G561), .O(G597) );
nand2 gate181( .a(G510), .b(G564), .O(G598) );
nand2 gate182( .a(G513), .b(G564), .O(G599) );
nand2 gate183( .a(G516), .b(G567), .O(G600) );
nand2 gate184( .a(G519), .b(G567), .O(G601) );
nand2 gate185( .a(G570), .b(G571), .O(G602) );

  xor2  gate1135(.a(G573), .b(G572), .O(gate186inter0));
  nand2 gate1136(.a(gate186inter0), .b(s_84), .O(gate186inter1));
  and2  gate1137(.a(G573), .b(G572), .O(gate186inter2));
  inv1  gate1138(.a(s_84), .O(gate186inter3));
  inv1  gate1139(.a(s_85), .O(gate186inter4));
  nand2 gate1140(.a(gate186inter4), .b(gate186inter3), .O(gate186inter5));
  nor2  gate1141(.a(gate186inter5), .b(gate186inter2), .O(gate186inter6));
  inv1  gate1142(.a(G572), .O(gate186inter7));
  inv1  gate1143(.a(G573), .O(gate186inter8));
  nand2 gate1144(.a(gate186inter8), .b(gate186inter7), .O(gate186inter9));
  nand2 gate1145(.a(s_85), .b(gate186inter3), .O(gate186inter10));
  nor2  gate1146(.a(gate186inter10), .b(gate186inter9), .O(gate186inter11));
  nor2  gate1147(.a(gate186inter11), .b(gate186inter6), .O(gate186inter12));
  nand2 gate1148(.a(gate186inter12), .b(gate186inter1), .O(G607));
nand2 gate187( .a(G574), .b(G575), .O(G612) );
nand2 gate188( .a(G576), .b(G577), .O(G617) );
nand2 gate189( .a(G578), .b(G579), .O(G622) );
nand2 gate190( .a(G580), .b(G581), .O(G627) );
nand2 gate191( .a(G582), .b(G583), .O(G632) );
nand2 gate192( .a(G584), .b(G585), .O(G637) );
nand2 gate193( .a(G586), .b(G587), .O(G642) );
nand2 gate194( .a(G588), .b(G589), .O(G645) );
nand2 gate195( .a(G590), .b(G591), .O(G648) );
nand2 gate196( .a(G592), .b(G593), .O(G651) );
nand2 gate197( .a(G594), .b(G595), .O(G654) );
nand2 gate198( .a(G596), .b(G597), .O(G657) );
nand2 gate199( .a(G598), .b(G599), .O(G660) );
nand2 gate200( .a(G600), .b(G601), .O(G663) );
nand2 gate201( .a(G602), .b(G607), .O(G666) );
nand2 gate202( .a(G612), .b(G617), .O(G669) );

  xor2  gate1471(.a(G612), .b(G602), .O(gate203inter0));
  nand2 gate1472(.a(gate203inter0), .b(s_132), .O(gate203inter1));
  and2  gate1473(.a(G612), .b(G602), .O(gate203inter2));
  inv1  gate1474(.a(s_132), .O(gate203inter3));
  inv1  gate1475(.a(s_133), .O(gate203inter4));
  nand2 gate1476(.a(gate203inter4), .b(gate203inter3), .O(gate203inter5));
  nor2  gate1477(.a(gate203inter5), .b(gate203inter2), .O(gate203inter6));
  inv1  gate1478(.a(G602), .O(gate203inter7));
  inv1  gate1479(.a(G612), .O(gate203inter8));
  nand2 gate1480(.a(gate203inter8), .b(gate203inter7), .O(gate203inter9));
  nand2 gate1481(.a(s_133), .b(gate203inter3), .O(gate203inter10));
  nor2  gate1482(.a(gate203inter10), .b(gate203inter9), .O(gate203inter11));
  nor2  gate1483(.a(gate203inter11), .b(gate203inter6), .O(gate203inter12));
  nand2 gate1484(.a(gate203inter12), .b(gate203inter1), .O(G672));
nand2 gate204( .a(G607), .b(G617), .O(G675) );

  xor2  gate1037(.a(G627), .b(G622), .O(gate205inter0));
  nand2 gate1038(.a(gate205inter0), .b(s_70), .O(gate205inter1));
  and2  gate1039(.a(G627), .b(G622), .O(gate205inter2));
  inv1  gate1040(.a(s_70), .O(gate205inter3));
  inv1  gate1041(.a(s_71), .O(gate205inter4));
  nand2 gate1042(.a(gate205inter4), .b(gate205inter3), .O(gate205inter5));
  nor2  gate1043(.a(gate205inter5), .b(gate205inter2), .O(gate205inter6));
  inv1  gate1044(.a(G622), .O(gate205inter7));
  inv1  gate1045(.a(G627), .O(gate205inter8));
  nand2 gate1046(.a(gate205inter8), .b(gate205inter7), .O(gate205inter9));
  nand2 gate1047(.a(s_71), .b(gate205inter3), .O(gate205inter10));
  nor2  gate1048(.a(gate205inter10), .b(gate205inter9), .O(gate205inter11));
  nor2  gate1049(.a(gate205inter11), .b(gate205inter6), .O(gate205inter12));
  nand2 gate1050(.a(gate205inter12), .b(gate205inter1), .O(G678));
nand2 gate206( .a(G632), .b(G637), .O(G681) );

  xor2  gate1345(.a(G632), .b(G622), .O(gate207inter0));
  nand2 gate1346(.a(gate207inter0), .b(s_114), .O(gate207inter1));
  and2  gate1347(.a(G632), .b(G622), .O(gate207inter2));
  inv1  gate1348(.a(s_114), .O(gate207inter3));
  inv1  gate1349(.a(s_115), .O(gate207inter4));
  nand2 gate1350(.a(gate207inter4), .b(gate207inter3), .O(gate207inter5));
  nor2  gate1351(.a(gate207inter5), .b(gate207inter2), .O(gate207inter6));
  inv1  gate1352(.a(G622), .O(gate207inter7));
  inv1  gate1353(.a(G632), .O(gate207inter8));
  nand2 gate1354(.a(gate207inter8), .b(gate207inter7), .O(gate207inter9));
  nand2 gate1355(.a(s_115), .b(gate207inter3), .O(gate207inter10));
  nor2  gate1356(.a(gate207inter10), .b(gate207inter9), .O(gate207inter11));
  nor2  gate1357(.a(gate207inter11), .b(gate207inter6), .O(gate207inter12));
  nand2 gate1358(.a(gate207inter12), .b(gate207inter1), .O(G684));
nand2 gate208( .a(G627), .b(G637), .O(G687) );
nand2 gate209( .a(G602), .b(G666), .O(G690) );
nand2 gate210( .a(G607), .b(G666), .O(G691) );
nand2 gate211( .a(G612), .b(G669), .O(G692) );
nand2 gate212( .a(G617), .b(G669), .O(G693) );
nand2 gate213( .a(G602), .b(G672), .O(G694) );
nand2 gate214( .a(G612), .b(G672), .O(G695) );
nand2 gate215( .a(G607), .b(G675), .O(G696) );

  xor2  gate1555(.a(G675), .b(G617), .O(gate216inter0));
  nand2 gate1556(.a(gate216inter0), .b(s_144), .O(gate216inter1));
  and2  gate1557(.a(G675), .b(G617), .O(gate216inter2));
  inv1  gate1558(.a(s_144), .O(gate216inter3));
  inv1  gate1559(.a(s_145), .O(gate216inter4));
  nand2 gate1560(.a(gate216inter4), .b(gate216inter3), .O(gate216inter5));
  nor2  gate1561(.a(gate216inter5), .b(gate216inter2), .O(gate216inter6));
  inv1  gate1562(.a(G617), .O(gate216inter7));
  inv1  gate1563(.a(G675), .O(gate216inter8));
  nand2 gate1564(.a(gate216inter8), .b(gate216inter7), .O(gate216inter9));
  nand2 gate1565(.a(s_145), .b(gate216inter3), .O(gate216inter10));
  nor2  gate1566(.a(gate216inter10), .b(gate216inter9), .O(gate216inter11));
  nor2  gate1567(.a(gate216inter11), .b(gate216inter6), .O(gate216inter12));
  nand2 gate1568(.a(gate216inter12), .b(gate216inter1), .O(G697));
nand2 gate217( .a(G622), .b(G678), .O(G698) );
nand2 gate218( .a(G627), .b(G678), .O(G699) );

  xor2  gate1373(.a(G681), .b(G632), .O(gate219inter0));
  nand2 gate1374(.a(gate219inter0), .b(s_118), .O(gate219inter1));
  and2  gate1375(.a(G681), .b(G632), .O(gate219inter2));
  inv1  gate1376(.a(s_118), .O(gate219inter3));
  inv1  gate1377(.a(s_119), .O(gate219inter4));
  nand2 gate1378(.a(gate219inter4), .b(gate219inter3), .O(gate219inter5));
  nor2  gate1379(.a(gate219inter5), .b(gate219inter2), .O(gate219inter6));
  inv1  gate1380(.a(G632), .O(gate219inter7));
  inv1  gate1381(.a(G681), .O(gate219inter8));
  nand2 gate1382(.a(gate219inter8), .b(gate219inter7), .O(gate219inter9));
  nand2 gate1383(.a(s_119), .b(gate219inter3), .O(gate219inter10));
  nor2  gate1384(.a(gate219inter10), .b(gate219inter9), .O(gate219inter11));
  nor2  gate1385(.a(gate219inter11), .b(gate219inter6), .O(gate219inter12));
  nand2 gate1386(.a(gate219inter12), .b(gate219inter1), .O(G700));
nand2 gate220( .a(G637), .b(G681), .O(G701) );
nand2 gate221( .a(G622), .b(G684), .O(G702) );
nand2 gate222( .a(G632), .b(G684), .O(G703) );

  xor2  gate1275(.a(G687), .b(G627), .O(gate223inter0));
  nand2 gate1276(.a(gate223inter0), .b(s_104), .O(gate223inter1));
  and2  gate1277(.a(G687), .b(G627), .O(gate223inter2));
  inv1  gate1278(.a(s_104), .O(gate223inter3));
  inv1  gate1279(.a(s_105), .O(gate223inter4));
  nand2 gate1280(.a(gate223inter4), .b(gate223inter3), .O(gate223inter5));
  nor2  gate1281(.a(gate223inter5), .b(gate223inter2), .O(gate223inter6));
  inv1  gate1282(.a(G627), .O(gate223inter7));
  inv1  gate1283(.a(G687), .O(gate223inter8));
  nand2 gate1284(.a(gate223inter8), .b(gate223inter7), .O(gate223inter9));
  nand2 gate1285(.a(s_105), .b(gate223inter3), .O(gate223inter10));
  nor2  gate1286(.a(gate223inter10), .b(gate223inter9), .O(gate223inter11));
  nor2  gate1287(.a(gate223inter11), .b(gate223inter6), .O(gate223inter12));
  nand2 gate1288(.a(gate223inter12), .b(gate223inter1), .O(G704));

  xor2  gate981(.a(G687), .b(G637), .O(gate224inter0));
  nand2 gate982(.a(gate224inter0), .b(s_62), .O(gate224inter1));
  and2  gate983(.a(G687), .b(G637), .O(gate224inter2));
  inv1  gate984(.a(s_62), .O(gate224inter3));
  inv1  gate985(.a(s_63), .O(gate224inter4));
  nand2 gate986(.a(gate224inter4), .b(gate224inter3), .O(gate224inter5));
  nor2  gate987(.a(gate224inter5), .b(gate224inter2), .O(gate224inter6));
  inv1  gate988(.a(G637), .O(gate224inter7));
  inv1  gate989(.a(G687), .O(gate224inter8));
  nand2 gate990(.a(gate224inter8), .b(gate224inter7), .O(gate224inter9));
  nand2 gate991(.a(s_63), .b(gate224inter3), .O(gate224inter10));
  nor2  gate992(.a(gate224inter10), .b(gate224inter9), .O(gate224inter11));
  nor2  gate993(.a(gate224inter11), .b(gate224inter6), .O(gate224inter12));
  nand2 gate994(.a(gate224inter12), .b(gate224inter1), .O(G705));
nand2 gate225( .a(G690), .b(G691), .O(G706) );

  xor2  gate1415(.a(G693), .b(G692), .O(gate226inter0));
  nand2 gate1416(.a(gate226inter0), .b(s_124), .O(gate226inter1));
  and2  gate1417(.a(G693), .b(G692), .O(gate226inter2));
  inv1  gate1418(.a(s_124), .O(gate226inter3));
  inv1  gate1419(.a(s_125), .O(gate226inter4));
  nand2 gate1420(.a(gate226inter4), .b(gate226inter3), .O(gate226inter5));
  nor2  gate1421(.a(gate226inter5), .b(gate226inter2), .O(gate226inter6));
  inv1  gate1422(.a(G692), .O(gate226inter7));
  inv1  gate1423(.a(G693), .O(gate226inter8));
  nand2 gate1424(.a(gate226inter8), .b(gate226inter7), .O(gate226inter9));
  nand2 gate1425(.a(s_125), .b(gate226inter3), .O(gate226inter10));
  nor2  gate1426(.a(gate226inter10), .b(gate226inter9), .O(gate226inter11));
  nor2  gate1427(.a(gate226inter11), .b(gate226inter6), .O(gate226inter12));
  nand2 gate1428(.a(gate226inter12), .b(gate226inter1), .O(G709));
nand2 gate227( .a(G694), .b(G695), .O(G712) );
nand2 gate228( .a(G696), .b(G697), .O(G715) );
nand2 gate229( .a(G698), .b(G699), .O(G718) );
nand2 gate230( .a(G700), .b(G701), .O(G721) );
nand2 gate231( .a(G702), .b(G703), .O(G724) );
nand2 gate232( .a(G704), .b(G705), .O(G727) );

  xor2  gate617(.a(G718), .b(G242), .O(gate233inter0));
  nand2 gate618(.a(gate233inter0), .b(s_10), .O(gate233inter1));
  and2  gate619(.a(G718), .b(G242), .O(gate233inter2));
  inv1  gate620(.a(s_10), .O(gate233inter3));
  inv1  gate621(.a(s_11), .O(gate233inter4));
  nand2 gate622(.a(gate233inter4), .b(gate233inter3), .O(gate233inter5));
  nor2  gate623(.a(gate233inter5), .b(gate233inter2), .O(gate233inter6));
  inv1  gate624(.a(G242), .O(gate233inter7));
  inv1  gate625(.a(G718), .O(gate233inter8));
  nand2 gate626(.a(gate233inter8), .b(gate233inter7), .O(gate233inter9));
  nand2 gate627(.a(s_11), .b(gate233inter3), .O(gate233inter10));
  nor2  gate628(.a(gate233inter10), .b(gate233inter9), .O(gate233inter11));
  nor2  gate629(.a(gate233inter11), .b(gate233inter6), .O(gate233inter12));
  nand2 gate630(.a(gate233inter12), .b(gate233inter1), .O(G730));
nand2 gate234( .a(G245), .b(G721), .O(G733) );

  xor2  gate1639(.a(G724), .b(G248), .O(gate235inter0));
  nand2 gate1640(.a(gate235inter0), .b(s_156), .O(gate235inter1));
  and2  gate1641(.a(G724), .b(G248), .O(gate235inter2));
  inv1  gate1642(.a(s_156), .O(gate235inter3));
  inv1  gate1643(.a(s_157), .O(gate235inter4));
  nand2 gate1644(.a(gate235inter4), .b(gate235inter3), .O(gate235inter5));
  nor2  gate1645(.a(gate235inter5), .b(gate235inter2), .O(gate235inter6));
  inv1  gate1646(.a(G248), .O(gate235inter7));
  inv1  gate1647(.a(G724), .O(gate235inter8));
  nand2 gate1648(.a(gate235inter8), .b(gate235inter7), .O(gate235inter9));
  nand2 gate1649(.a(s_157), .b(gate235inter3), .O(gate235inter10));
  nor2  gate1650(.a(gate235inter10), .b(gate235inter9), .O(gate235inter11));
  nor2  gate1651(.a(gate235inter11), .b(gate235inter6), .O(gate235inter12));
  nand2 gate1652(.a(gate235inter12), .b(gate235inter1), .O(G736));
nand2 gate236( .a(G251), .b(G727), .O(G739) );
nand2 gate237( .a(G254), .b(G706), .O(G742) );
nand2 gate238( .a(G257), .b(G709), .O(G745) );
nand2 gate239( .a(G260), .b(G712), .O(G748) );

  xor2  gate673(.a(G715), .b(G263), .O(gate240inter0));
  nand2 gate674(.a(gate240inter0), .b(s_18), .O(gate240inter1));
  and2  gate675(.a(G715), .b(G263), .O(gate240inter2));
  inv1  gate676(.a(s_18), .O(gate240inter3));
  inv1  gate677(.a(s_19), .O(gate240inter4));
  nand2 gate678(.a(gate240inter4), .b(gate240inter3), .O(gate240inter5));
  nor2  gate679(.a(gate240inter5), .b(gate240inter2), .O(gate240inter6));
  inv1  gate680(.a(G263), .O(gate240inter7));
  inv1  gate681(.a(G715), .O(gate240inter8));
  nand2 gate682(.a(gate240inter8), .b(gate240inter7), .O(gate240inter9));
  nand2 gate683(.a(s_19), .b(gate240inter3), .O(gate240inter10));
  nor2  gate684(.a(gate240inter10), .b(gate240inter9), .O(gate240inter11));
  nor2  gate685(.a(gate240inter11), .b(gate240inter6), .O(gate240inter12));
  nand2 gate686(.a(gate240inter12), .b(gate240inter1), .O(G751));
nand2 gate241( .a(G242), .b(G730), .O(G754) );
nand2 gate242( .a(G718), .b(G730), .O(G755) );
nand2 gate243( .a(G245), .b(G733), .O(G756) );
nand2 gate244( .a(G721), .b(G733), .O(G757) );

  xor2  gate785(.a(G736), .b(G248), .O(gate245inter0));
  nand2 gate786(.a(gate245inter0), .b(s_34), .O(gate245inter1));
  and2  gate787(.a(G736), .b(G248), .O(gate245inter2));
  inv1  gate788(.a(s_34), .O(gate245inter3));
  inv1  gate789(.a(s_35), .O(gate245inter4));
  nand2 gate790(.a(gate245inter4), .b(gate245inter3), .O(gate245inter5));
  nor2  gate791(.a(gate245inter5), .b(gate245inter2), .O(gate245inter6));
  inv1  gate792(.a(G248), .O(gate245inter7));
  inv1  gate793(.a(G736), .O(gate245inter8));
  nand2 gate794(.a(gate245inter8), .b(gate245inter7), .O(gate245inter9));
  nand2 gate795(.a(s_35), .b(gate245inter3), .O(gate245inter10));
  nor2  gate796(.a(gate245inter10), .b(gate245inter9), .O(gate245inter11));
  nor2  gate797(.a(gate245inter11), .b(gate245inter6), .O(gate245inter12));
  nand2 gate798(.a(gate245inter12), .b(gate245inter1), .O(G758));

  xor2  gate1219(.a(G736), .b(G724), .O(gate246inter0));
  nand2 gate1220(.a(gate246inter0), .b(s_96), .O(gate246inter1));
  and2  gate1221(.a(G736), .b(G724), .O(gate246inter2));
  inv1  gate1222(.a(s_96), .O(gate246inter3));
  inv1  gate1223(.a(s_97), .O(gate246inter4));
  nand2 gate1224(.a(gate246inter4), .b(gate246inter3), .O(gate246inter5));
  nor2  gate1225(.a(gate246inter5), .b(gate246inter2), .O(gate246inter6));
  inv1  gate1226(.a(G724), .O(gate246inter7));
  inv1  gate1227(.a(G736), .O(gate246inter8));
  nand2 gate1228(.a(gate246inter8), .b(gate246inter7), .O(gate246inter9));
  nand2 gate1229(.a(s_97), .b(gate246inter3), .O(gate246inter10));
  nor2  gate1230(.a(gate246inter10), .b(gate246inter9), .O(gate246inter11));
  nor2  gate1231(.a(gate246inter11), .b(gate246inter6), .O(gate246inter12));
  nand2 gate1232(.a(gate246inter12), .b(gate246inter1), .O(G759));

  xor2  gate855(.a(G739), .b(G251), .O(gate247inter0));
  nand2 gate856(.a(gate247inter0), .b(s_44), .O(gate247inter1));
  and2  gate857(.a(G739), .b(G251), .O(gate247inter2));
  inv1  gate858(.a(s_44), .O(gate247inter3));
  inv1  gate859(.a(s_45), .O(gate247inter4));
  nand2 gate860(.a(gate247inter4), .b(gate247inter3), .O(gate247inter5));
  nor2  gate861(.a(gate247inter5), .b(gate247inter2), .O(gate247inter6));
  inv1  gate862(.a(G251), .O(gate247inter7));
  inv1  gate863(.a(G739), .O(gate247inter8));
  nand2 gate864(.a(gate247inter8), .b(gate247inter7), .O(gate247inter9));
  nand2 gate865(.a(s_45), .b(gate247inter3), .O(gate247inter10));
  nor2  gate866(.a(gate247inter10), .b(gate247inter9), .O(gate247inter11));
  nor2  gate867(.a(gate247inter11), .b(gate247inter6), .O(gate247inter12));
  nand2 gate868(.a(gate247inter12), .b(gate247inter1), .O(G760));
nand2 gate248( .a(G727), .b(G739), .O(G761) );
nand2 gate249( .a(G254), .b(G742), .O(G762) );
nand2 gate250( .a(G706), .b(G742), .O(G763) );

  xor2  gate1261(.a(G745), .b(G257), .O(gate251inter0));
  nand2 gate1262(.a(gate251inter0), .b(s_102), .O(gate251inter1));
  and2  gate1263(.a(G745), .b(G257), .O(gate251inter2));
  inv1  gate1264(.a(s_102), .O(gate251inter3));
  inv1  gate1265(.a(s_103), .O(gate251inter4));
  nand2 gate1266(.a(gate251inter4), .b(gate251inter3), .O(gate251inter5));
  nor2  gate1267(.a(gate251inter5), .b(gate251inter2), .O(gate251inter6));
  inv1  gate1268(.a(G257), .O(gate251inter7));
  inv1  gate1269(.a(G745), .O(gate251inter8));
  nand2 gate1270(.a(gate251inter8), .b(gate251inter7), .O(gate251inter9));
  nand2 gate1271(.a(s_103), .b(gate251inter3), .O(gate251inter10));
  nor2  gate1272(.a(gate251inter10), .b(gate251inter9), .O(gate251inter11));
  nor2  gate1273(.a(gate251inter11), .b(gate251inter6), .O(gate251inter12));
  nand2 gate1274(.a(gate251inter12), .b(gate251inter1), .O(G764));

  xor2  gate729(.a(G745), .b(G709), .O(gate252inter0));
  nand2 gate730(.a(gate252inter0), .b(s_26), .O(gate252inter1));
  and2  gate731(.a(G745), .b(G709), .O(gate252inter2));
  inv1  gate732(.a(s_26), .O(gate252inter3));
  inv1  gate733(.a(s_27), .O(gate252inter4));
  nand2 gate734(.a(gate252inter4), .b(gate252inter3), .O(gate252inter5));
  nor2  gate735(.a(gate252inter5), .b(gate252inter2), .O(gate252inter6));
  inv1  gate736(.a(G709), .O(gate252inter7));
  inv1  gate737(.a(G745), .O(gate252inter8));
  nand2 gate738(.a(gate252inter8), .b(gate252inter7), .O(gate252inter9));
  nand2 gate739(.a(s_27), .b(gate252inter3), .O(gate252inter10));
  nor2  gate740(.a(gate252inter10), .b(gate252inter9), .O(gate252inter11));
  nor2  gate741(.a(gate252inter11), .b(gate252inter6), .O(gate252inter12));
  nand2 gate742(.a(gate252inter12), .b(gate252inter1), .O(G765));
nand2 gate253( .a(G260), .b(G748), .O(G766) );
nand2 gate254( .a(G712), .b(G748), .O(G767) );

  xor2  gate659(.a(G751), .b(G263), .O(gate255inter0));
  nand2 gate660(.a(gate255inter0), .b(s_16), .O(gate255inter1));
  and2  gate661(.a(G751), .b(G263), .O(gate255inter2));
  inv1  gate662(.a(s_16), .O(gate255inter3));
  inv1  gate663(.a(s_17), .O(gate255inter4));
  nand2 gate664(.a(gate255inter4), .b(gate255inter3), .O(gate255inter5));
  nor2  gate665(.a(gate255inter5), .b(gate255inter2), .O(gate255inter6));
  inv1  gate666(.a(G263), .O(gate255inter7));
  inv1  gate667(.a(G751), .O(gate255inter8));
  nand2 gate668(.a(gate255inter8), .b(gate255inter7), .O(gate255inter9));
  nand2 gate669(.a(s_17), .b(gate255inter3), .O(gate255inter10));
  nor2  gate670(.a(gate255inter10), .b(gate255inter9), .O(gate255inter11));
  nor2  gate671(.a(gate255inter11), .b(gate255inter6), .O(gate255inter12));
  nand2 gate672(.a(gate255inter12), .b(gate255inter1), .O(G768));
nand2 gate256( .a(G715), .b(G751), .O(G769) );
nand2 gate257( .a(G754), .b(G755), .O(G770) );
nand2 gate258( .a(G756), .b(G757), .O(G773) );
nand2 gate259( .a(G758), .b(G759), .O(G776) );

  xor2  gate1205(.a(G761), .b(G760), .O(gate260inter0));
  nand2 gate1206(.a(gate260inter0), .b(s_94), .O(gate260inter1));
  and2  gate1207(.a(G761), .b(G760), .O(gate260inter2));
  inv1  gate1208(.a(s_94), .O(gate260inter3));
  inv1  gate1209(.a(s_95), .O(gate260inter4));
  nand2 gate1210(.a(gate260inter4), .b(gate260inter3), .O(gate260inter5));
  nor2  gate1211(.a(gate260inter5), .b(gate260inter2), .O(gate260inter6));
  inv1  gate1212(.a(G760), .O(gate260inter7));
  inv1  gate1213(.a(G761), .O(gate260inter8));
  nand2 gate1214(.a(gate260inter8), .b(gate260inter7), .O(gate260inter9));
  nand2 gate1215(.a(s_95), .b(gate260inter3), .O(gate260inter10));
  nor2  gate1216(.a(gate260inter10), .b(gate260inter9), .O(gate260inter11));
  nor2  gate1217(.a(gate260inter11), .b(gate260inter6), .O(gate260inter12));
  nand2 gate1218(.a(gate260inter12), .b(gate260inter1), .O(G779));
nand2 gate261( .a(G762), .b(G763), .O(G782) );
nand2 gate262( .a(G764), .b(G765), .O(G785) );
nand2 gate263( .a(G766), .b(G767), .O(G788) );
nand2 gate264( .a(G768), .b(G769), .O(G791) );
nand2 gate265( .a(G642), .b(G770), .O(G794) );
nand2 gate266( .a(G645), .b(G773), .O(G797) );
nand2 gate267( .a(G648), .b(G776), .O(G800) );
nand2 gate268( .a(G651), .b(G779), .O(G803) );

  xor2  gate771(.a(G782), .b(G654), .O(gate269inter0));
  nand2 gate772(.a(gate269inter0), .b(s_32), .O(gate269inter1));
  and2  gate773(.a(G782), .b(G654), .O(gate269inter2));
  inv1  gate774(.a(s_32), .O(gate269inter3));
  inv1  gate775(.a(s_33), .O(gate269inter4));
  nand2 gate776(.a(gate269inter4), .b(gate269inter3), .O(gate269inter5));
  nor2  gate777(.a(gate269inter5), .b(gate269inter2), .O(gate269inter6));
  inv1  gate778(.a(G654), .O(gate269inter7));
  inv1  gate779(.a(G782), .O(gate269inter8));
  nand2 gate780(.a(gate269inter8), .b(gate269inter7), .O(gate269inter9));
  nand2 gate781(.a(s_33), .b(gate269inter3), .O(gate269inter10));
  nor2  gate782(.a(gate269inter10), .b(gate269inter9), .O(gate269inter11));
  nor2  gate783(.a(gate269inter11), .b(gate269inter6), .O(gate269inter12));
  nand2 gate784(.a(gate269inter12), .b(gate269inter1), .O(G806));
nand2 gate270( .a(G657), .b(G785), .O(G809) );
nand2 gate271( .a(G660), .b(G788), .O(G812) );

  xor2  gate1233(.a(G791), .b(G663), .O(gate272inter0));
  nand2 gate1234(.a(gate272inter0), .b(s_98), .O(gate272inter1));
  and2  gate1235(.a(G791), .b(G663), .O(gate272inter2));
  inv1  gate1236(.a(s_98), .O(gate272inter3));
  inv1  gate1237(.a(s_99), .O(gate272inter4));
  nand2 gate1238(.a(gate272inter4), .b(gate272inter3), .O(gate272inter5));
  nor2  gate1239(.a(gate272inter5), .b(gate272inter2), .O(gate272inter6));
  inv1  gate1240(.a(G663), .O(gate272inter7));
  inv1  gate1241(.a(G791), .O(gate272inter8));
  nand2 gate1242(.a(gate272inter8), .b(gate272inter7), .O(gate272inter9));
  nand2 gate1243(.a(s_99), .b(gate272inter3), .O(gate272inter10));
  nor2  gate1244(.a(gate272inter10), .b(gate272inter9), .O(gate272inter11));
  nor2  gate1245(.a(gate272inter11), .b(gate272inter6), .O(gate272inter12));
  nand2 gate1246(.a(gate272inter12), .b(gate272inter1), .O(G815));
nand2 gate273( .a(G642), .b(G794), .O(G818) );
nand2 gate274( .a(G770), .b(G794), .O(G819) );
nand2 gate275( .a(G645), .b(G797), .O(G820) );
nand2 gate276( .a(G773), .b(G797), .O(G821) );
nand2 gate277( .a(G648), .b(G800), .O(G822) );
nand2 gate278( .a(G776), .b(G800), .O(G823) );

  xor2  gate1597(.a(G803), .b(G651), .O(gate279inter0));
  nand2 gate1598(.a(gate279inter0), .b(s_150), .O(gate279inter1));
  and2  gate1599(.a(G803), .b(G651), .O(gate279inter2));
  inv1  gate1600(.a(s_150), .O(gate279inter3));
  inv1  gate1601(.a(s_151), .O(gate279inter4));
  nand2 gate1602(.a(gate279inter4), .b(gate279inter3), .O(gate279inter5));
  nor2  gate1603(.a(gate279inter5), .b(gate279inter2), .O(gate279inter6));
  inv1  gate1604(.a(G651), .O(gate279inter7));
  inv1  gate1605(.a(G803), .O(gate279inter8));
  nand2 gate1606(.a(gate279inter8), .b(gate279inter7), .O(gate279inter9));
  nand2 gate1607(.a(s_151), .b(gate279inter3), .O(gate279inter10));
  nor2  gate1608(.a(gate279inter10), .b(gate279inter9), .O(gate279inter11));
  nor2  gate1609(.a(gate279inter11), .b(gate279inter6), .O(gate279inter12));
  nand2 gate1610(.a(gate279inter12), .b(gate279inter1), .O(G824));
nand2 gate280( .a(G779), .b(G803), .O(G825) );
nand2 gate281( .a(G654), .b(G806), .O(G826) );
nand2 gate282( .a(G782), .b(G806), .O(G827) );
nand2 gate283( .a(G657), .b(G809), .O(G828) );
nand2 gate284( .a(G785), .b(G809), .O(G829) );

  xor2  gate1065(.a(G812), .b(G660), .O(gate285inter0));
  nand2 gate1066(.a(gate285inter0), .b(s_74), .O(gate285inter1));
  and2  gate1067(.a(G812), .b(G660), .O(gate285inter2));
  inv1  gate1068(.a(s_74), .O(gate285inter3));
  inv1  gate1069(.a(s_75), .O(gate285inter4));
  nand2 gate1070(.a(gate285inter4), .b(gate285inter3), .O(gate285inter5));
  nor2  gate1071(.a(gate285inter5), .b(gate285inter2), .O(gate285inter6));
  inv1  gate1072(.a(G660), .O(gate285inter7));
  inv1  gate1073(.a(G812), .O(gate285inter8));
  nand2 gate1074(.a(gate285inter8), .b(gate285inter7), .O(gate285inter9));
  nand2 gate1075(.a(s_75), .b(gate285inter3), .O(gate285inter10));
  nor2  gate1076(.a(gate285inter10), .b(gate285inter9), .O(gate285inter11));
  nor2  gate1077(.a(gate285inter11), .b(gate285inter6), .O(gate285inter12));
  nand2 gate1078(.a(gate285inter12), .b(gate285inter1), .O(G830));

  xor2  gate757(.a(G812), .b(G788), .O(gate286inter0));
  nand2 gate758(.a(gate286inter0), .b(s_30), .O(gate286inter1));
  and2  gate759(.a(G812), .b(G788), .O(gate286inter2));
  inv1  gate760(.a(s_30), .O(gate286inter3));
  inv1  gate761(.a(s_31), .O(gate286inter4));
  nand2 gate762(.a(gate286inter4), .b(gate286inter3), .O(gate286inter5));
  nor2  gate763(.a(gate286inter5), .b(gate286inter2), .O(gate286inter6));
  inv1  gate764(.a(G788), .O(gate286inter7));
  inv1  gate765(.a(G812), .O(gate286inter8));
  nand2 gate766(.a(gate286inter8), .b(gate286inter7), .O(gate286inter9));
  nand2 gate767(.a(s_31), .b(gate286inter3), .O(gate286inter10));
  nor2  gate768(.a(gate286inter10), .b(gate286inter9), .O(gate286inter11));
  nor2  gate769(.a(gate286inter11), .b(gate286inter6), .O(gate286inter12));
  nand2 gate770(.a(gate286inter12), .b(gate286inter1), .O(G831));

  xor2  gate1079(.a(G815), .b(G663), .O(gate287inter0));
  nand2 gate1080(.a(gate287inter0), .b(s_76), .O(gate287inter1));
  and2  gate1081(.a(G815), .b(G663), .O(gate287inter2));
  inv1  gate1082(.a(s_76), .O(gate287inter3));
  inv1  gate1083(.a(s_77), .O(gate287inter4));
  nand2 gate1084(.a(gate287inter4), .b(gate287inter3), .O(gate287inter5));
  nor2  gate1085(.a(gate287inter5), .b(gate287inter2), .O(gate287inter6));
  inv1  gate1086(.a(G663), .O(gate287inter7));
  inv1  gate1087(.a(G815), .O(gate287inter8));
  nand2 gate1088(.a(gate287inter8), .b(gate287inter7), .O(gate287inter9));
  nand2 gate1089(.a(s_77), .b(gate287inter3), .O(gate287inter10));
  nor2  gate1090(.a(gate287inter10), .b(gate287inter9), .O(gate287inter11));
  nor2  gate1091(.a(gate287inter11), .b(gate287inter6), .O(gate287inter12));
  nand2 gate1092(.a(gate287inter12), .b(gate287inter1), .O(G832));

  xor2  gate1331(.a(G815), .b(G791), .O(gate288inter0));
  nand2 gate1332(.a(gate288inter0), .b(s_112), .O(gate288inter1));
  and2  gate1333(.a(G815), .b(G791), .O(gate288inter2));
  inv1  gate1334(.a(s_112), .O(gate288inter3));
  inv1  gate1335(.a(s_113), .O(gate288inter4));
  nand2 gate1336(.a(gate288inter4), .b(gate288inter3), .O(gate288inter5));
  nor2  gate1337(.a(gate288inter5), .b(gate288inter2), .O(gate288inter6));
  inv1  gate1338(.a(G791), .O(gate288inter7));
  inv1  gate1339(.a(G815), .O(gate288inter8));
  nand2 gate1340(.a(gate288inter8), .b(gate288inter7), .O(gate288inter9));
  nand2 gate1341(.a(s_113), .b(gate288inter3), .O(gate288inter10));
  nor2  gate1342(.a(gate288inter10), .b(gate288inter9), .O(gate288inter11));
  nor2  gate1343(.a(gate288inter11), .b(gate288inter6), .O(gate288inter12));
  nand2 gate1344(.a(gate288inter12), .b(gate288inter1), .O(G833));
nand2 gate289( .a(G818), .b(G819), .O(G834) );
nand2 gate290( .a(G820), .b(G821), .O(G847) );
nand2 gate291( .a(G822), .b(G823), .O(G860) );
nand2 gate292( .a(G824), .b(G825), .O(G873) );
nand2 gate293( .a(G828), .b(G829), .O(G886) );
nand2 gate294( .a(G832), .b(G833), .O(G899) );
nand2 gate295( .a(G830), .b(G831), .O(G912) );
nand2 gate296( .a(G826), .b(G827), .O(G925) );
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );

  xor2  gate1177(.a(G1036), .b(G1), .O(gate387inter0));
  nand2 gate1178(.a(gate387inter0), .b(s_90), .O(gate387inter1));
  and2  gate1179(.a(G1036), .b(G1), .O(gate387inter2));
  inv1  gate1180(.a(s_90), .O(gate387inter3));
  inv1  gate1181(.a(s_91), .O(gate387inter4));
  nand2 gate1182(.a(gate387inter4), .b(gate387inter3), .O(gate387inter5));
  nor2  gate1183(.a(gate387inter5), .b(gate387inter2), .O(gate387inter6));
  inv1  gate1184(.a(G1), .O(gate387inter7));
  inv1  gate1185(.a(G1036), .O(gate387inter8));
  nand2 gate1186(.a(gate387inter8), .b(gate387inter7), .O(gate387inter9));
  nand2 gate1187(.a(s_91), .b(gate387inter3), .O(gate387inter10));
  nor2  gate1188(.a(gate387inter10), .b(gate387inter9), .O(gate387inter11));
  nor2  gate1189(.a(gate387inter11), .b(gate387inter6), .O(gate387inter12));
  nand2 gate1190(.a(gate387inter12), .b(gate387inter1), .O(G1132));
nand2 gate388( .a(G2), .b(G1039), .O(G1135) );
nand2 gate389( .a(G3), .b(G1042), .O(G1138) );
nand2 gate390( .a(G4), .b(G1045), .O(G1141) );

  xor2  gate1051(.a(G1048), .b(G5), .O(gate391inter0));
  nand2 gate1052(.a(gate391inter0), .b(s_72), .O(gate391inter1));
  and2  gate1053(.a(G1048), .b(G5), .O(gate391inter2));
  inv1  gate1054(.a(s_72), .O(gate391inter3));
  inv1  gate1055(.a(s_73), .O(gate391inter4));
  nand2 gate1056(.a(gate391inter4), .b(gate391inter3), .O(gate391inter5));
  nor2  gate1057(.a(gate391inter5), .b(gate391inter2), .O(gate391inter6));
  inv1  gate1058(.a(G5), .O(gate391inter7));
  inv1  gate1059(.a(G1048), .O(gate391inter8));
  nand2 gate1060(.a(gate391inter8), .b(gate391inter7), .O(gate391inter9));
  nand2 gate1061(.a(s_73), .b(gate391inter3), .O(gate391inter10));
  nor2  gate1062(.a(gate391inter10), .b(gate391inter9), .O(gate391inter11));
  nor2  gate1063(.a(gate391inter11), .b(gate391inter6), .O(gate391inter12));
  nand2 gate1064(.a(gate391inter12), .b(gate391inter1), .O(G1144));
nand2 gate392( .a(G6), .b(G1051), .O(G1147) );
nand2 gate393( .a(G7), .b(G1054), .O(G1150) );
nand2 gate394( .a(G8), .b(G1057), .O(G1153) );
nand2 gate395( .a(G9), .b(G1060), .O(G1156) );
nand2 gate396( .a(G10), .b(G1063), .O(G1159) );
nand2 gate397( .a(G11), .b(G1066), .O(G1162) );
nand2 gate398( .a(G12), .b(G1069), .O(G1165) );
nand2 gate399( .a(G13), .b(G1072), .O(G1168) );
nand2 gate400( .a(G14), .b(G1075), .O(G1171) );
nand2 gate401( .a(G15), .b(G1078), .O(G1174) );

  xor2  gate1457(.a(G1081), .b(G16), .O(gate402inter0));
  nand2 gate1458(.a(gate402inter0), .b(s_130), .O(gate402inter1));
  and2  gate1459(.a(G1081), .b(G16), .O(gate402inter2));
  inv1  gate1460(.a(s_130), .O(gate402inter3));
  inv1  gate1461(.a(s_131), .O(gate402inter4));
  nand2 gate1462(.a(gate402inter4), .b(gate402inter3), .O(gate402inter5));
  nor2  gate1463(.a(gate402inter5), .b(gate402inter2), .O(gate402inter6));
  inv1  gate1464(.a(G16), .O(gate402inter7));
  inv1  gate1465(.a(G1081), .O(gate402inter8));
  nand2 gate1466(.a(gate402inter8), .b(gate402inter7), .O(gate402inter9));
  nand2 gate1467(.a(s_131), .b(gate402inter3), .O(gate402inter10));
  nor2  gate1468(.a(gate402inter10), .b(gate402inter9), .O(gate402inter11));
  nor2  gate1469(.a(gate402inter11), .b(gate402inter6), .O(gate402inter12));
  nand2 gate1470(.a(gate402inter12), .b(gate402inter1), .O(G1177));
nand2 gate403( .a(G17), .b(G1084), .O(G1180) );
nand2 gate404( .a(G18), .b(G1087), .O(G1183) );
nand2 gate405( .a(G19), .b(G1090), .O(G1186) );
nand2 gate406( .a(G20), .b(G1093), .O(G1189) );

  xor2  gate1569(.a(G1096), .b(G21), .O(gate407inter0));
  nand2 gate1570(.a(gate407inter0), .b(s_146), .O(gate407inter1));
  and2  gate1571(.a(G1096), .b(G21), .O(gate407inter2));
  inv1  gate1572(.a(s_146), .O(gate407inter3));
  inv1  gate1573(.a(s_147), .O(gate407inter4));
  nand2 gate1574(.a(gate407inter4), .b(gate407inter3), .O(gate407inter5));
  nor2  gate1575(.a(gate407inter5), .b(gate407inter2), .O(gate407inter6));
  inv1  gate1576(.a(G21), .O(gate407inter7));
  inv1  gate1577(.a(G1096), .O(gate407inter8));
  nand2 gate1578(.a(gate407inter8), .b(gate407inter7), .O(gate407inter9));
  nand2 gate1579(.a(s_147), .b(gate407inter3), .O(gate407inter10));
  nor2  gate1580(.a(gate407inter10), .b(gate407inter9), .O(gate407inter11));
  nor2  gate1581(.a(gate407inter11), .b(gate407inter6), .O(gate407inter12));
  nand2 gate1582(.a(gate407inter12), .b(gate407inter1), .O(G1192));
nand2 gate408( .a(G22), .b(G1099), .O(G1195) );
nand2 gate409( .a(G23), .b(G1102), .O(G1198) );

  xor2  gate939(.a(G1105), .b(G24), .O(gate410inter0));
  nand2 gate940(.a(gate410inter0), .b(s_56), .O(gate410inter1));
  and2  gate941(.a(G1105), .b(G24), .O(gate410inter2));
  inv1  gate942(.a(s_56), .O(gate410inter3));
  inv1  gate943(.a(s_57), .O(gate410inter4));
  nand2 gate944(.a(gate410inter4), .b(gate410inter3), .O(gate410inter5));
  nor2  gate945(.a(gate410inter5), .b(gate410inter2), .O(gate410inter6));
  inv1  gate946(.a(G24), .O(gate410inter7));
  inv1  gate947(.a(G1105), .O(gate410inter8));
  nand2 gate948(.a(gate410inter8), .b(gate410inter7), .O(gate410inter9));
  nand2 gate949(.a(s_57), .b(gate410inter3), .O(gate410inter10));
  nor2  gate950(.a(gate410inter10), .b(gate410inter9), .O(gate410inter11));
  nor2  gate951(.a(gate410inter11), .b(gate410inter6), .O(gate410inter12));
  nand2 gate952(.a(gate410inter12), .b(gate410inter1), .O(G1201));
nand2 gate411( .a(G25), .b(G1108), .O(G1204) );
nand2 gate412( .a(G26), .b(G1111), .O(G1207) );
nand2 gate413( .a(G27), .b(G1114), .O(G1210) );

  xor2  gate995(.a(G1117), .b(G28), .O(gate414inter0));
  nand2 gate996(.a(gate414inter0), .b(s_64), .O(gate414inter1));
  and2  gate997(.a(G1117), .b(G28), .O(gate414inter2));
  inv1  gate998(.a(s_64), .O(gate414inter3));
  inv1  gate999(.a(s_65), .O(gate414inter4));
  nand2 gate1000(.a(gate414inter4), .b(gate414inter3), .O(gate414inter5));
  nor2  gate1001(.a(gate414inter5), .b(gate414inter2), .O(gate414inter6));
  inv1  gate1002(.a(G28), .O(gate414inter7));
  inv1  gate1003(.a(G1117), .O(gate414inter8));
  nand2 gate1004(.a(gate414inter8), .b(gate414inter7), .O(gate414inter9));
  nand2 gate1005(.a(s_65), .b(gate414inter3), .O(gate414inter10));
  nor2  gate1006(.a(gate414inter10), .b(gate414inter9), .O(gate414inter11));
  nor2  gate1007(.a(gate414inter11), .b(gate414inter6), .O(gate414inter12));
  nand2 gate1008(.a(gate414inter12), .b(gate414inter1), .O(G1213));
nand2 gate415( .a(G29), .b(G1120), .O(G1216) );
nand2 gate416( .a(G30), .b(G1123), .O(G1219) );

  xor2  gate1009(.a(G1126), .b(G31), .O(gate417inter0));
  nand2 gate1010(.a(gate417inter0), .b(s_66), .O(gate417inter1));
  and2  gate1011(.a(G1126), .b(G31), .O(gate417inter2));
  inv1  gate1012(.a(s_66), .O(gate417inter3));
  inv1  gate1013(.a(s_67), .O(gate417inter4));
  nand2 gate1014(.a(gate417inter4), .b(gate417inter3), .O(gate417inter5));
  nor2  gate1015(.a(gate417inter5), .b(gate417inter2), .O(gate417inter6));
  inv1  gate1016(.a(G31), .O(gate417inter7));
  inv1  gate1017(.a(G1126), .O(gate417inter8));
  nand2 gate1018(.a(gate417inter8), .b(gate417inter7), .O(gate417inter9));
  nand2 gate1019(.a(s_67), .b(gate417inter3), .O(gate417inter10));
  nor2  gate1020(.a(gate417inter10), .b(gate417inter9), .O(gate417inter11));
  nor2  gate1021(.a(gate417inter11), .b(gate417inter6), .O(gate417inter12));
  nand2 gate1022(.a(gate417inter12), .b(gate417inter1), .O(G1222));

  xor2  gate1429(.a(G1129), .b(G32), .O(gate418inter0));
  nand2 gate1430(.a(gate418inter0), .b(s_126), .O(gate418inter1));
  and2  gate1431(.a(G1129), .b(G32), .O(gate418inter2));
  inv1  gate1432(.a(s_126), .O(gate418inter3));
  inv1  gate1433(.a(s_127), .O(gate418inter4));
  nand2 gate1434(.a(gate418inter4), .b(gate418inter3), .O(gate418inter5));
  nor2  gate1435(.a(gate418inter5), .b(gate418inter2), .O(gate418inter6));
  inv1  gate1436(.a(G32), .O(gate418inter7));
  inv1  gate1437(.a(G1129), .O(gate418inter8));
  nand2 gate1438(.a(gate418inter8), .b(gate418inter7), .O(gate418inter9));
  nand2 gate1439(.a(s_127), .b(gate418inter3), .O(gate418inter10));
  nor2  gate1440(.a(gate418inter10), .b(gate418inter9), .O(gate418inter11));
  nor2  gate1441(.a(gate418inter11), .b(gate418inter6), .O(gate418inter12));
  nand2 gate1442(.a(gate418inter12), .b(gate418inter1), .O(G1225));
nand2 gate419( .a(G1), .b(G1132), .O(G1228) );
nand2 gate420( .a(G1036), .b(G1132), .O(G1229) );
nand2 gate421( .a(G2), .b(G1135), .O(G1230) );
nand2 gate422( .a(G1039), .b(G1135), .O(G1231) );
nand2 gate423( .a(G3), .b(G1138), .O(G1232) );
nand2 gate424( .a(G1042), .b(G1138), .O(G1233) );
nand2 gate425( .a(G4), .b(G1141), .O(G1234) );
nand2 gate426( .a(G1045), .b(G1141), .O(G1235) );
nand2 gate427( .a(G5), .b(G1144), .O(G1236) );
nand2 gate428( .a(G1048), .b(G1144), .O(G1237) );

  xor2  gate967(.a(G1147), .b(G6), .O(gate429inter0));
  nand2 gate968(.a(gate429inter0), .b(s_60), .O(gate429inter1));
  and2  gate969(.a(G1147), .b(G6), .O(gate429inter2));
  inv1  gate970(.a(s_60), .O(gate429inter3));
  inv1  gate971(.a(s_61), .O(gate429inter4));
  nand2 gate972(.a(gate429inter4), .b(gate429inter3), .O(gate429inter5));
  nor2  gate973(.a(gate429inter5), .b(gate429inter2), .O(gate429inter6));
  inv1  gate974(.a(G6), .O(gate429inter7));
  inv1  gate975(.a(G1147), .O(gate429inter8));
  nand2 gate976(.a(gate429inter8), .b(gate429inter7), .O(gate429inter9));
  nand2 gate977(.a(s_61), .b(gate429inter3), .O(gate429inter10));
  nor2  gate978(.a(gate429inter10), .b(gate429inter9), .O(gate429inter11));
  nor2  gate979(.a(gate429inter11), .b(gate429inter6), .O(gate429inter12));
  nand2 gate980(.a(gate429inter12), .b(gate429inter1), .O(G1238));
nand2 gate430( .a(G1051), .b(G1147), .O(G1239) );
nand2 gate431( .a(G7), .b(G1150), .O(G1240) );

  xor2  gate1485(.a(G1150), .b(G1054), .O(gate432inter0));
  nand2 gate1486(.a(gate432inter0), .b(s_134), .O(gate432inter1));
  and2  gate1487(.a(G1150), .b(G1054), .O(gate432inter2));
  inv1  gate1488(.a(s_134), .O(gate432inter3));
  inv1  gate1489(.a(s_135), .O(gate432inter4));
  nand2 gate1490(.a(gate432inter4), .b(gate432inter3), .O(gate432inter5));
  nor2  gate1491(.a(gate432inter5), .b(gate432inter2), .O(gate432inter6));
  inv1  gate1492(.a(G1054), .O(gate432inter7));
  inv1  gate1493(.a(G1150), .O(gate432inter8));
  nand2 gate1494(.a(gate432inter8), .b(gate432inter7), .O(gate432inter9));
  nand2 gate1495(.a(s_135), .b(gate432inter3), .O(gate432inter10));
  nor2  gate1496(.a(gate432inter10), .b(gate432inter9), .O(gate432inter11));
  nor2  gate1497(.a(gate432inter11), .b(gate432inter6), .O(gate432inter12));
  nand2 gate1498(.a(gate432inter12), .b(gate432inter1), .O(G1241));
nand2 gate433( .a(G8), .b(G1153), .O(G1242) );
nand2 gate434( .a(G1057), .b(G1153), .O(G1243) );
nand2 gate435( .a(G9), .b(G1156), .O(G1244) );
nand2 gate436( .a(G1060), .b(G1156), .O(G1245) );
nand2 gate437( .a(G10), .b(G1159), .O(G1246) );
nand2 gate438( .a(G1063), .b(G1159), .O(G1247) );
nand2 gate439( .a(G11), .b(G1162), .O(G1248) );
nand2 gate440( .a(G1066), .b(G1162), .O(G1249) );
nand2 gate441( .a(G12), .b(G1165), .O(G1250) );
nand2 gate442( .a(G1069), .b(G1165), .O(G1251) );
nand2 gate443( .a(G13), .b(G1168), .O(G1252) );
nand2 gate444( .a(G1072), .b(G1168), .O(G1253) );
nand2 gate445( .a(G14), .b(G1171), .O(G1254) );
nand2 gate446( .a(G1075), .b(G1171), .O(G1255) );
nand2 gate447( .a(G15), .b(G1174), .O(G1256) );
nand2 gate448( .a(G1078), .b(G1174), .O(G1257) );
nand2 gate449( .a(G16), .b(G1177), .O(G1258) );

  xor2  gate799(.a(G1177), .b(G1081), .O(gate450inter0));
  nand2 gate800(.a(gate450inter0), .b(s_36), .O(gate450inter1));
  and2  gate801(.a(G1177), .b(G1081), .O(gate450inter2));
  inv1  gate802(.a(s_36), .O(gate450inter3));
  inv1  gate803(.a(s_37), .O(gate450inter4));
  nand2 gate804(.a(gate450inter4), .b(gate450inter3), .O(gate450inter5));
  nor2  gate805(.a(gate450inter5), .b(gate450inter2), .O(gate450inter6));
  inv1  gate806(.a(G1081), .O(gate450inter7));
  inv1  gate807(.a(G1177), .O(gate450inter8));
  nand2 gate808(.a(gate450inter8), .b(gate450inter7), .O(gate450inter9));
  nand2 gate809(.a(s_37), .b(gate450inter3), .O(gate450inter10));
  nor2  gate810(.a(gate450inter10), .b(gate450inter9), .O(gate450inter11));
  nor2  gate811(.a(gate450inter11), .b(gate450inter6), .O(gate450inter12));
  nand2 gate812(.a(gate450inter12), .b(gate450inter1), .O(G1259));
nand2 gate451( .a(G17), .b(G1180), .O(G1260) );
nand2 gate452( .a(G1084), .b(G1180), .O(G1261) );
nand2 gate453( .a(G18), .b(G1183), .O(G1262) );
nand2 gate454( .a(G1087), .b(G1183), .O(G1263) );
nand2 gate455( .a(G19), .b(G1186), .O(G1264) );

  xor2  gate1443(.a(G1186), .b(G1090), .O(gate456inter0));
  nand2 gate1444(.a(gate456inter0), .b(s_128), .O(gate456inter1));
  and2  gate1445(.a(G1186), .b(G1090), .O(gate456inter2));
  inv1  gate1446(.a(s_128), .O(gate456inter3));
  inv1  gate1447(.a(s_129), .O(gate456inter4));
  nand2 gate1448(.a(gate456inter4), .b(gate456inter3), .O(gate456inter5));
  nor2  gate1449(.a(gate456inter5), .b(gate456inter2), .O(gate456inter6));
  inv1  gate1450(.a(G1090), .O(gate456inter7));
  inv1  gate1451(.a(G1186), .O(gate456inter8));
  nand2 gate1452(.a(gate456inter8), .b(gate456inter7), .O(gate456inter9));
  nand2 gate1453(.a(s_129), .b(gate456inter3), .O(gate456inter10));
  nor2  gate1454(.a(gate456inter10), .b(gate456inter9), .O(gate456inter11));
  nor2  gate1455(.a(gate456inter11), .b(gate456inter6), .O(gate456inter12));
  nand2 gate1456(.a(gate456inter12), .b(gate456inter1), .O(G1265));
nand2 gate457( .a(G20), .b(G1189), .O(G1266) );
nand2 gate458( .a(G1093), .b(G1189), .O(G1267) );

  xor2  gate1247(.a(G1192), .b(G21), .O(gate459inter0));
  nand2 gate1248(.a(gate459inter0), .b(s_100), .O(gate459inter1));
  and2  gate1249(.a(G1192), .b(G21), .O(gate459inter2));
  inv1  gate1250(.a(s_100), .O(gate459inter3));
  inv1  gate1251(.a(s_101), .O(gate459inter4));
  nand2 gate1252(.a(gate459inter4), .b(gate459inter3), .O(gate459inter5));
  nor2  gate1253(.a(gate459inter5), .b(gate459inter2), .O(gate459inter6));
  inv1  gate1254(.a(G21), .O(gate459inter7));
  inv1  gate1255(.a(G1192), .O(gate459inter8));
  nand2 gate1256(.a(gate459inter8), .b(gate459inter7), .O(gate459inter9));
  nand2 gate1257(.a(s_101), .b(gate459inter3), .O(gate459inter10));
  nor2  gate1258(.a(gate459inter10), .b(gate459inter9), .O(gate459inter11));
  nor2  gate1259(.a(gate459inter11), .b(gate459inter6), .O(gate459inter12));
  nand2 gate1260(.a(gate459inter12), .b(gate459inter1), .O(G1268));
nand2 gate460( .a(G1096), .b(G1192), .O(G1269) );
nand2 gate461( .a(G22), .b(G1195), .O(G1270) );
nand2 gate462( .a(G1099), .b(G1195), .O(G1271) );
nand2 gate463( .a(G23), .b(G1198), .O(G1272) );
nand2 gate464( .a(G1102), .b(G1198), .O(G1273) );
nand2 gate465( .a(G24), .b(G1201), .O(G1274) );
nand2 gate466( .a(G1105), .b(G1201), .O(G1275) );
nand2 gate467( .a(G25), .b(G1204), .O(G1276) );

  xor2  gate1401(.a(G1204), .b(G1108), .O(gate468inter0));
  nand2 gate1402(.a(gate468inter0), .b(s_122), .O(gate468inter1));
  and2  gate1403(.a(G1204), .b(G1108), .O(gate468inter2));
  inv1  gate1404(.a(s_122), .O(gate468inter3));
  inv1  gate1405(.a(s_123), .O(gate468inter4));
  nand2 gate1406(.a(gate468inter4), .b(gate468inter3), .O(gate468inter5));
  nor2  gate1407(.a(gate468inter5), .b(gate468inter2), .O(gate468inter6));
  inv1  gate1408(.a(G1108), .O(gate468inter7));
  inv1  gate1409(.a(G1204), .O(gate468inter8));
  nand2 gate1410(.a(gate468inter8), .b(gate468inter7), .O(gate468inter9));
  nand2 gate1411(.a(s_123), .b(gate468inter3), .O(gate468inter10));
  nor2  gate1412(.a(gate468inter10), .b(gate468inter9), .O(gate468inter11));
  nor2  gate1413(.a(gate468inter11), .b(gate468inter6), .O(gate468inter12));
  nand2 gate1414(.a(gate468inter12), .b(gate468inter1), .O(G1277));
nand2 gate469( .a(G26), .b(G1207), .O(G1278) );
nand2 gate470( .a(G1111), .b(G1207), .O(G1279) );
nand2 gate471( .a(G27), .b(G1210), .O(G1280) );

  xor2  gate1387(.a(G1210), .b(G1114), .O(gate472inter0));
  nand2 gate1388(.a(gate472inter0), .b(s_120), .O(gate472inter1));
  and2  gate1389(.a(G1210), .b(G1114), .O(gate472inter2));
  inv1  gate1390(.a(s_120), .O(gate472inter3));
  inv1  gate1391(.a(s_121), .O(gate472inter4));
  nand2 gate1392(.a(gate472inter4), .b(gate472inter3), .O(gate472inter5));
  nor2  gate1393(.a(gate472inter5), .b(gate472inter2), .O(gate472inter6));
  inv1  gate1394(.a(G1114), .O(gate472inter7));
  inv1  gate1395(.a(G1210), .O(gate472inter8));
  nand2 gate1396(.a(gate472inter8), .b(gate472inter7), .O(gate472inter9));
  nand2 gate1397(.a(s_121), .b(gate472inter3), .O(gate472inter10));
  nor2  gate1398(.a(gate472inter10), .b(gate472inter9), .O(gate472inter11));
  nor2  gate1399(.a(gate472inter11), .b(gate472inter6), .O(gate472inter12));
  nand2 gate1400(.a(gate472inter12), .b(gate472inter1), .O(G1281));
nand2 gate473( .a(G28), .b(G1213), .O(G1282) );
nand2 gate474( .a(G1117), .b(G1213), .O(G1283) );

  xor2  gate631(.a(G1216), .b(G29), .O(gate475inter0));
  nand2 gate632(.a(gate475inter0), .b(s_12), .O(gate475inter1));
  and2  gate633(.a(G1216), .b(G29), .O(gate475inter2));
  inv1  gate634(.a(s_12), .O(gate475inter3));
  inv1  gate635(.a(s_13), .O(gate475inter4));
  nand2 gate636(.a(gate475inter4), .b(gate475inter3), .O(gate475inter5));
  nor2  gate637(.a(gate475inter5), .b(gate475inter2), .O(gate475inter6));
  inv1  gate638(.a(G29), .O(gate475inter7));
  inv1  gate639(.a(G1216), .O(gate475inter8));
  nand2 gate640(.a(gate475inter8), .b(gate475inter7), .O(gate475inter9));
  nand2 gate641(.a(s_13), .b(gate475inter3), .O(gate475inter10));
  nor2  gate642(.a(gate475inter10), .b(gate475inter9), .O(gate475inter11));
  nor2  gate643(.a(gate475inter11), .b(gate475inter6), .O(gate475inter12));
  nand2 gate644(.a(gate475inter12), .b(gate475inter1), .O(G1284));
nand2 gate476( .a(G1120), .b(G1216), .O(G1285) );
nand2 gate477( .a(G30), .b(G1219), .O(G1286) );

  xor2  gate743(.a(G1219), .b(G1123), .O(gate478inter0));
  nand2 gate744(.a(gate478inter0), .b(s_28), .O(gate478inter1));
  and2  gate745(.a(G1219), .b(G1123), .O(gate478inter2));
  inv1  gate746(.a(s_28), .O(gate478inter3));
  inv1  gate747(.a(s_29), .O(gate478inter4));
  nand2 gate748(.a(gate478inter4), .b(gate478inter3), .O(gate478inter5));
  nor2  gate749(.a(gate478inter5), .b(gate478inter2), .O(gate478inter6));
  inv1  gate750(.a(G1123), .O(gate478inter7));
  inv1  gate751(.a(G1219), .O(gate478inter8));
  nand2 gate752(.a(gate478inter8), .b(gate478inter7), .O(gate478inter9));
  nand2 gate753(.a(s_29), .b(gate478inter3), .O(gate478inter10));
  nor2  gate754(.a(gate478inter10), .b(gate478inter9), .O(gate478inter11));
  nor2  gate755(.a(gate478inter11), .b(gate478inter6), .O(gate478inter12));
  nand2 gate756(.a(gate478inter12), .b(gate478inter1), .O(G1287));
nand2 gate479( .a(G31), .b(G1222), .O(G1288) );
nand2 gate480( .a(G1126), .b(G1222), .O(G1289) );

  xor2  gate1499(.a(G1225), .b(G32), .O(gate481inter0));
  nand2 gate1500(.a(gate481inter0), .b(s_136), .O(gate481inter1));
  and2  gate1501(.a(G1225), .b(G32), .O(gate481inter2));
  inv1  gate1502(.a(s_136), .O(gate481inter3));
  inv1  gate1503(.a(s_137), .O(gate481inter4));
  nand2 gate1504(.a(gate481inter4), .b(gate481inter3), .O(gate481inter5));
  nor2  gate1505(.a(gate481inter5), .b(gate481inter2), .O(gate481inter6));
  inv1  gate1506(.a(G32), .O(gate481inter7));
  inv1  gate1507(.a(G1225), .O(gate481inter8));
  nand2 gate1508(.a(gate481inter8), .b(gate481inter7), .O(gate481inter9));
  nand2 gate1509(.a(s_137), .b(gate481inter3), .O(gate481inter10));
  nor2  gate1510(.a(gate481inter10), .b(gate481inter9), .O(gate481inter11));
  nor2  gate1511(.a(gate481inter11), .b(gate481inter6), .O(gate481inter12));
  nand2 gate1512(.a(gate481inter12), .b(gate481inter1), .O(G1290));
nand2 gate482( .a(G1129), .b(G1225), .O(G1291) );
nand2 gate483( .a(G1228), .b(G1229), .O(G1292) );
nand2 gate484( .a(G1230), .b(G1231), .O(G1293) );
nand2 gate485( .a(G1232), .b(G1233), .O(G1294) );

  xor2  gate911(.a(G1235), .b(G1234), .O(gate486inter0));
  nand2 gate912(.a(gate486inter0), .b(s_52), .O(gate486inter1));
  and2  gate913(.a(G1235), .b(G1234), .O(gate486inter2));
  inv1  gate914(.a(s_52), .O(gate486inter3));
  inv1  gate915(.a(s_53), .O(gate486inter4));
  nand2 gate916(.a(gate486inter4), .b(gate486inter3), .O(gate486inter5));
  nor2  gate917(.a(gate486inter5), .b(gate486inter2), .O(gate486inter6));
  inv1  gate918(.a(G1234), .O(gate486inter7));
  inv1  gate919(.a(G1235), .O(gate486inter8));
  nand2 gate920(.a(gate486inter8), .b(gate486inter7), .O(gate486inter9));
  nand2 gate921(.a(s_53), .b(gate486inter3), .O(gate486inter10));
  nor2  gate922(.a(gate486inter10), .b(gate486inter9), .O(gate486inter11));
  nor2  gate923(.a(gate486inter11), .b(gate486inter6), .O(gate486inter12));
  nand2 gate924(.a(gate486inter12), .b(gate486inter1), .O(G1295));
nand2 gate487( .a(G1236), .b(G1237), .O(G1296) );

  xor2  gate1513(.a(G1239), .b(G1238), .O(gate488inter0));
  nand2 gate1514(.a(gate488inter0), .b(s_138), .O(gate488inter1));
  and2  gate1515(.a(G1239), .b(G1238), .O(gate488inter2));
  inv1  gate1516(.a(s_138), .O(gate488inter3));
  inv1  gate1517(.a(s_139), .O(gate488inter4));
  nand2 gate1518(.a(gate488inter4), .b(gate488inter3), .O(gate488inter5));
  nor2  gate1519(.a(gate488inter5), .b(gate488inter2), .O(gate488inter6));
  inv1  gate1520(.a(G1238), .O(gate488inter7));
  inv1  gate1521(.a(G1239), .O(gate488inter8));
  nand2 gate1522(.a(gate488inter8), .b(gate488inter7), .O(gate488inter9));
  nand2 gate1523(.a(s_139), .b(gate488inter3), .O(gate488inter10));
  nor2  gate1524(.a(gate488inter10), .b(gate488inter9), .O(gate488inter11));
  nor2  gate1525(.a(gate488inter11), .b(gate488inter6), .O(gate488inter12));
  nand2 gate1526(.a(gate488inter12), .b(gate488inter1), .O(G1297));
nand2 gate489( .a(G1240), .b(G1241), .O(G1298) );
nand2 gate490( .a(G1242), .b(G1243), .O(G1299) );
nand2 gate491( .a(G1244), .b(G1245), .O(G1300) );
nand2 gate492( .a(G1246), .b(G1247), .O(G1301) );
nand2 gate493( .a(G1248), .b(G1249), .O(G1302) );
nand2 gate494( .a(G1250), .b(G1251), .O(G1303) );
nand2 gate495( .a(G1252), .b(G1253), .O(G1304) );
nand2 gate496( .a(G1254), .b(G1255), .O(G1305) );
nand2 gate497( .a(G1256), .b(G1257), .O(G1306) );
nand2 gate498( .a(G1258), .b(G1259), .O(G1307) );
nand2 gate499( .a(G1260), .b(G1261), .O(G1308) );
nand2 gate500( .a(G1262), .b(G1263), .O(G1309) );

  xor2  gate1667(.a(G1265), .b(G1264), .O(gate501inter0));
  nand2 gate1668(.a(gate501inter0), .b(s_160), .O(gate501inter1));
  and2  gate1669(.a(G1265), .b(G1264), .O(gate501inter2));
  inv1  gate1670(.a(s_160), .O(gate501inter3));
  inv1  gate1671(.a(s_161), .O(gate501inter4));
  nand2 gate1672(.a(gate501inter4), .b(gate501inter3), .O(gate501inter5));
  nor2  gate1673(.a(gate501inter5), .b(gate501inter2), .O(gate501inter6));
  inv1  gate1674(.a(G1264), .O(gate501inter7));
  inv1  gate1675(.a(G1265), .O(gate501inter8));
  nand2 gate1676(.a(gate501inter8), .b(gate501inter7), .O(gate501inter9));
  nand2 gate1677(.a(s_161), .b(gate501inter3), .O(gate501inter10));
  nor2  gate1678(.a(gate501inter10), .b(gate501inter9), .O(gate501inter11));
  nor2  gate1679(.a(gate501inter11), .b(gate501inter6), .O(gate501inter12));
  nand2 gate1680(.a(gate501inter12), .b(gate501inter1), .O(G1310));
nand2 gate502( .a(G1266), .b(G1267), .O(G1311) );
nand2 gate503( .a(G1268), .b(G1269), .O(G1312) );
nand2 gate504( .a(G1270), .b(G1271), .O(G1313) );
nand2 gate505( .a(G1272), .b(G1273), .O(G1314) );
nand2 gate506( .a(G1274), .b(G1275), .O(G1315) );

  xor2  gate1653(.a(G1277), .b(G1276), .O(gate507inter0));
  nand2 gate1654(.a(gate507inter0), .b(s_158), .O(gate507inter1));
  and2  gate1655(.a(G1277), .b(G1276), .O(gate507inter2));
  inv1  gate1656(.a(s_158), .O(gate507inter3));
  inv1  gate1657(.a(s_159), .O(gate507inter4));
  nand2 gate1658(.a(gate507inter4), .b(gate507inter3), .O(gate507inter5));
  nor2  gate1659(.a(gate507inter5), .b(gate507inter2), .O(gate507inter6));
  inv1  gate1660(.a(G1276), .O(gate507inter7));
  inv1  gate1661(.a(G1277), .O(gate507inter8));
  nand2 gate1662(.a(gate507inter8), .b(gate507inter7), .O(gate507inter9));
  nand2 gate1663(.a(s_159), .b(gate507inter3), .O(gate507inter10));
  nor2  gate1664(.a(gate507inter10), .b(gate507inter9), .O(gate507inter11));
  nor2  gate1665(.a(gate507inter11), .b(gate507inter6), .O(gate507inter12));
  nand2 gate1666(.a(gate507inter12), .b(gate507inter1), .O(G1316));
nand2 gate508( .a(G1278), .b(G1279), .O(G1317) );
nand2 gate509( .a(G1280), .b(G1281), .O(G1318) );
nand2 gate510( .a(G1282), .b(G1283), .O(G1319) );
nand2 gate511( .a(G1284), .b(G1285), .O(G1320) );
nand2 gate512( .a(G1286), .b(G1287), .O(G1321) );
nand2 gate513( .a(G1288), .b(G1289), .O(G1322) );
nand2 gate514( .a(G1290), .b(G1291), .O(G1323) );
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule