module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);

input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;//RE__PI;

input s_0,s_1;//RE__ALLOW(00,01,10,11);
input s_2,s_3;//RE__ALLOW(00,01,10,11);
input s_4,s_5;//RE__ALLOW(00,01,10,11);
input s_6,s_7;//RE__ALLOW(00,01,10,11);
input s_8,s_9;//RE__ALLOW(00,01,10,11);
input s_10,s_11;//RE__ALLOW(00,01,10,11);
input s_12,s_13;//RE__ALLOW(00,01,10,11);
input s_14,s_15;//RE__ALLOW(00,01,10,11);
input s_16,s_17;//RE__ALLOW(00,01,10,11);
input s_18,s_19;//RE__ALLOW(00,01,10,11);
input s_20,s_21;//RE__ALLOW(00,01,10,11);
input s_22,s_23;//RE__ALLOW(00,01,10,11);
input s_24,s_25;//RE__ALLOW(00,01,10,11);
input s_26,s_27;//RE__ALLOW(00,01,10,11);
input s_28,s_29;//RE__ALLOW(00,01,10,11);
input s_30,s_31;//RE__ALLOW(00,01,10,11);
input s_32,s_33;//RE__ALLOW(00,01,10,11);
input s_34,s_35;//RE__ALLOW(00,01,10,11);
input s_36,s_37;//RE__ALLOW(00,01,10,11);
input s_38,s_39;//RE__ALLOW(00,01,10,11);
input s_40,s_41;//RE__ALLOW(00,01,10,11);
input s_42,s_43;//RE__ALLOW(00,01,10,11);
input s_44,s_45;//RE__ALLOW(00,01,10,11);
input s_46,s_47;//RE__ALLOW(00,01,10,11);
input s_48,s_49;//RE__ALLOW(00,01,10,11);
input s_50,s_51;//RE__ALLOW(00,01,10,11);
input s_52,s_53;//RE__ALLOW(00,01,10,11);
input s_54,s_55;//RE__ALLOW(00,01,10,11);
input s_56,s_57;//RE__ALLOW(00,01,10,11);
input s_58,s_59;//RE__ALLOW(00,01,10,11);
input s_60,s_61;//RE__ALLOW(00,01,10,11);
input s_62,s_63;//RE__ALLOW(00,01,10,11);
input s_64,s_65;//RE__ALLOW(00,01,10,11);
input s_66,s_67;//RE__ALLOW(00,01,10,11);
input s_68,s_69;//RE__ALLOW(00,01,10,11);
input s_70,s_71;//RE__ALLOW(00,01,10,11);
input s_72,s_73;//RE__ALLOW(00,01,10,11);
input s_74,s_75;//RE__ALLOW(00,01,10,11);
input s_76,s_77;//RE__ALLOW(00,01,10,11);
input s_78,s_79;//RE__ALLOW(00,01,10,11);
input s_80,s_81;//RE__ALLOW(00,01,10,11);
input s_82,s_83;//RE__ALLOW(00,01,10,11);
input s_84,s_85;//RE__ALLOW(00,01,10,11);
input s_86,s_87;//RE__ALLOW(00,01,10,11);
input s_88,s_89;//RE__ALLOW(00,01,10,11);
input s_90,s_91;//RE__ALLOW(00,01,10,11);
input s_92,s_93;//RE__ALLOW(00,01,10,11);
input s_94,s_95;//RE__ALLOW(00,01,10,11);
input s_96,s_97;//RE__ALLOW(00,01,10,11);
input s_98,s_99;//RE__ALLOW(00,01,10,11);
input s_100,s_101;//RE__ALLOW(00,01,10,11);
input s_102,s_103;//RE__ALLOW(00,01,10,11);
input s_104,s_105;//RE__ALLOW(00,01,10,11);
input s_106,s_107;//RE__ALLOW(00,01,10,11);
input s_108,s_109;//RE__ALLOW(00,01,10,11);
input s_110,s_111;//RE__ALLOW(00,01,10,11);
input s_112,s_113;//RE__ALLOW(00,01,10,11);
input s_114,s_115;//RE__ALLOW(00,01,10,11);
input s_116,s_117;//RE__ALLOW(00,01,10,11);
input s_118,s_119;//RE__ALLOW(00,01,10,11);
input s_120,s_121;//RE__ALLOW(00,01,10,11);
input s_122,s_123;//RE__ALLOW(00,01,10,11);
input s_124,s_125;//RE__ALLOW(00,01,10,11);
input s_126,s_127;//RE__ALLOW(00,01,10,11);
input s_128,s_129;//RE__ALLOW(00,01,10,11);
input s_130,s_131;//RE__ALLOW(00,01,10,11);
input s_132,s_133;//RE__ALLOW(00,01,10,11);
input s_134,s_135;//RE__ALLOW(00,01,10,11);
input s_136,s_137;//RE__ALLOW(00,01,10,11);
input s_138,s_139;//RE__ALLOW(00,01,10,11);
input s_140,s_141;//RE__ALLOW(00,01,10,11);
input s_142,s_143;//RE__ALLOW(00,01,10,11);
input s_144,s_145;//RE__ALLOW(00,01,10,11);
input s_146,s_147;//RE__ALLOW(00,01,10,11);
input s_148,s_149;//RE__ALLOW(00,01,10,11);
input s_150,s_151;//RE__ALLOW(00,01,10,11);
input s_152,s_153;//RE__ALLOW(00,01,10,11);
input s_154,s_155;//RE__ALLOW(00,01,10,11);
input s_156,s_157;//RE__ALLOW(00,01,10,11);
input s_158,s_159;//RE__ALLOW(00,01,10,11);
input s_160,s_161;//RE__ALLOW(00,01,10,11);
input s_162,s_163;//RE__ALLOW(00,01,10,11);
input s_164,s_165;//RE__ALLOW(00,01,10,11);
input s_166,s_167;//RE__ALLOW(00,01,10,11);
input s_168,s_169;//RE__ALLOW(00,01,10,11);
input s_170,s_171;//RE__ALLOW(00,01,10,11);
input s_172,s_173;//RE__ALLOW(00,01,10,11);
input s_174,s_175;//RE__ALLOW(00,01,10,11);
input s_176,s_177;//RE__ALLOW(00,01,10,11);
input s_178,s_179;//RE__ALLOW(00,01,10,11);
input s_180,s_181;//RE__ALLOW(00,01,10,11);
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;

  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate401inter0, gate401inter1, gate401inter2, gate401inter3, gate401inter4, gate401inter5, gate401inter6, gate401inter7, gate401inter8, gate401inter9, gate401inter10, gate401inter11, gate401inter12, gate489inter0, gate489inter1, gate489inter2, gate489inter3, gate489inter4, gate489inter5, gate489inter6, gate489inter7, gate489inter8, gate489inter9, gate489inter10, gate489inter11, gate489inter12, gate186inter0, gate186inter1, gate186inter2, gate186inter3, gate186inter4, gate186inter5, gate186inter6, gate186inter7, gate186inter8, gate186inter9, gate186inter10, gate186inter11, gate186inter12, gate123inter0, gate123inter1, gate123inter2, gate123inter3, gate123inter4, gate123inter5, gate123inter6, gate123inter7, gate123inter8, gate123inter9, gate123inter10, gate123inter11, gate123inter12, gate206inter0, gate206inter1, gate206inter2, gate206inter3, gate206inter4, gate206inter5, gate206inter6, gate206inter7, gate206inter8, gate206inter9, gate206inter10, gate206inter11, gate206inter12, gate83inter0, gate83inter1, gate83inter2, gate83inter3, gate83inter4, gate83inter5, gate83inter6, gate83inter7, gate83inter8, gate83inter9, gate83inter10, gate83inter11, gate83inter12, gate196inter0, gate196inter1, gate196inter2, gate196inter3, gate196inter4, gate196inter5, gate196inter6, gate196inter7, gate196inter8, gate196inter9, gate196inter10, gate196inter11, gate196inter12, gate395inter0, gate395inter1, gate395inter2, gate395inter3, gate395inter4, gate395inter5, gate395inter6, gate395inter7, gate395inter8, gate395inter9, gate395inter10, gate395inter11, gate395inter12, gate465inter0, gate465inter1, gate465inter2, gate465inter3, gate465inter4, gate465inter5, gate465inter6, gate465inter7, gate465inter8, gate465inter9, gate465inter10, gate465inter11, gate465inter12, gate413inter0, gate413inter1, gate413inter2, gate413inter3, gate413inter4, gate413inter5, gate413inter6, gate413inter7, gate413inter8, gate413inter9, gate413inter10, gate413inter11, gate413inter12, gate512inter0, gate512inter1, gate512inter2, gate512inter3, gate512inter4, gate512inter5, gate512inter6, gate512inter7, gate512inter8, gate512inter9, gate512inter10, gate512inter11, gate512inter12, gate258inter0, gate258inter1, gate258inter2, gate258inter3, gate258inter4, gate258inter5, gate258inter6, gate258inter7, gate258inter8, gate258inter9, gate258inter10, gate258inter11, gate258inter12, gate226inter0, gate226inter1, gate226inter2, gate226inter3, gate226inter4, gate226inter5, gate226inter6, gate226inter7, gate226inter8, gate226inter9, gate226inter10, gate226inter11, gate226inter12, gate421inter0, gate421inter1, gate421inter2, gate421inter3, gate421inter4, gate421inter5, gate421inter6, gate421inter7, gate421inter8, gate421inter9, gate421inter10, gate421inter11, gate421inter12, gate56inter0, gate56inter1, gate56inter2, gate56inter3, gate56inter4, gate56inter5, gate56inter6, gate56inter7, gate56inter8, gate56inter9, gate56inter10, gate56inter11, gate56inter12, gate481inter0, gate481inter1, gate481inter2, gate481inter3, gate481inter4, gate481inter5, gate481inter6, gate481inter7, gate481inter8, gate481inter9, gate481inter10, gate481inter11, gate481inter12, gate40inter0, gate40inter1, gate40inter2, gate40inter3, gate40inter4, gate40inter5, gate40inter6, gate40inter7, gate40inter8, gate40inter9, gate40inter10, gate40inter11, gate40inter12, gate103inter0, gate103inter1, gate103inter2, gate103inter3, gate103inter4, gate103inter5, gate103inter6, gate103inter7, gate103inter8, gate103inter9, gate103inter10, gate103inter11, gate103inter12, gate16inter0, gate16inter1, gate16inter2, gate16inter3, gate16inter4, gate16inter5, gate16inter6, gate16inter7, gate16inter8, gate16inter9, gate16inter10, gate16inter11, gate16inter12, gate100inter0, gate100inter1, gate100inter2, gate100inter3, gate100inter4, gate100inter5, gate100inter6, gate100inter7, gate100inter8, gate100inter9, gate100inter10, gate100inter11, gate100inter12, gate441inter0, gate441inter1, gate441inter2, gate441inter3, gate441inter4, gate441inter5, gate441inter6, gate441inter7, gate441inter8, gate441inter9, gate441inter10, gate441inter11, gate441inter12, gate236inter0, gate236inter1, gate236inter2, gate236inter3, gate236inter4, gate236inter5, gate236inter6, gate236inter7, gate236inter8, gate236inter9, gate236inter10, gate236inter11, gate236inter12, gate387inter0, gate387inter1, gate387inter2, gate387inter3, gate387inter4, gate387inter5, gate387inter6, gate387inter7, gate387inter8, gate387inter9, gate387inter10, gate387inter11, gate387inter12, gate128inter0, gate128inter1, gate128inter2, gate128inter3, gate128inter4, gate128inter5, gate128inter6, gate128inter7, gate128inter8, gate128inter9, gate128inter10, gate128inter11, gate128inter12, gate392inter0, gate392inter1, gate392inter2, gate392inter3, gate392inter4, gate392inter5, gate392inter6, gate392inter7, gate392inter8, gate392inter9, gate392inter10, gate392inter11, gate392inter12, gate116inter0, gate116inter1, gate116inter2, gate116inter3, gate116inter4, gate116inter5, gate116inter6, gate116inter7, gate116inter8, gate116inter9, gate116inter10, gate116inter11, gate116inter12, gate51inter0, gate51inter1, gate51inter2, gate51inter3, gate51inter4, gate51inter5, gate51inter6, gate51inter7, gate51inter8, gate51inter9, gate51inter10, gate51inter11, gate51inter12, gate483inter0, gate483inter1, gate483inter2, gate483inter3, gate483inter4, gate483inter5, gate483inter6, gate483inter7, gate483inter8, gate483inter9, gate483inter10, gate483inter11, gate483inter12, gate29inter0, gate29inter1, gate29inter2, gate29inter3, gate29inter4, gate29inter5, gate29inter6, gate29inter7, gate29inter8, gate29inter9, gate29inter10, gate29inter11, gate29inter12, gate462inter0, gate462inter1, gate462inter2, gate462inter3, gate462inter4, gate462inter5, gate462inter6, gate462inter7, gate462inter8, gate462inter9, gate462inter10, gate462inter11, gate462inter12, gate470inter0, gate470inter1, gate470inter2, gate470inter3, gate470inter4, gate470inter5, gate470inter6, gate470inter7, gate470inter8, gate470inter9, gate470inter10, gate470inter11, gate470inter12, gate188inter0, gate188inter1, gate188inter2, gate188inter3, gate188inter4, gate188inter5, gate188inter6, gate188inter7, gate188inter8, gate188inter9, gate188inter10, gate188inter11, gate188inter12, gate132inter0, gate132inter1, gate132inter2, gate132inter3, gate132inter4, gate132inter5, gate132inter6, gate132inter7, gate132inter8, gate132inter9, gate132inter10, gate132inter11, gate132inter12, gate198inter0, gate198inter1, gate198inter2, gate198inter3, gate198inter4, gate198inter5, gate198inter6, gate198inter7, gate198inter8, gate198inter9, gate198inter10, gate198inter11, gate198inter12, gate244inter0, gate244inter1, gate244inter2, gate244inter3, gate244inter4, gate244inter5, gate244inter6, gate244inter7, gate244inter8, gate244inter9, gate244inter10, gate244inter11, gate244inter12, gate35inter0, gate35inter1, gate35inter2, gate35inter3, gate35inter4, gate35inter5, gate35inter6, gate35inter7, gate35inter8, gate35inter9, gate35inter10, gate35inter11, gate35inter12, gate487inter0, gate487inter1, gate487inter2, gate487inter3, gate487inter4, gate487inter5, gate487inter6, gate487inter7, gate487inter8, gate487inter9, gate487inter10, gate487inter11, gate487inter12, gate133inter0, gate133inter1, gate133inter2, gate133inter3, gate133inter4, gate133inter5, gate133inter6, gate133inter7, gate133inter8, gate133inter9, gate133inter10, gate133inter11, gate133inter12, gate216inter0, gate216inter1, gate216inter2, gate216inter3, gate216inter4, gate216inter5, gate216inter6, gate216inter7, gate216inter8, gate216inter9, gate216inter10, gate216inter11, gate216inter12, gate280inter0, gate280inter1, gate280inter2, gate280inter3, gate280inter4, gate280inter5, gate280inter6, gate280inter7, gate280inter8, gate280inter9, gate280inter10, gate280inter11, gate280inter12, gate131inter0, gate131inter1, gate131inter2, gate131inter3, gate131inter4, gate131inter5, gate131inter6, gate131inter7, gate131inter8, gate131inter9, gate131inter10, gate131inter11, gate131inter12, gate488inter0, gate488inter1, gate488inter2, gate488inter3, gate488inter4, gate488inter5, gate488inter6, gate488inter7, gate488inter8, gate488inter9, gate488inter10, gate488inter11, gate488inter12, gate493inter0, gate493inter1, gate493inter2, gate493inter3, gate493inter4, gate493inter5, gate493inter6, gate493inter7, gate493inter8, gate493inter9, gate493inter10, gate493inter11, gate493inter12, gate252inter0, gate252inter1, gate252inter2, gate252inter3, gate252inter4, gate252inter5, gate252inter6, gate252inter7, gate252inter8, gate252inter9, gate252inter10, gate252inter11, gate252inter12, gate24inter0, gate24inter1, gate24inter2, gate24inter3, gate24inter4, gate24inter5, gate24inter6, gate24inter7, gate24inter8, gate24inter9, gate24inter10, gate24inter11, gate24inter12, gate394inter0, gate394inter1, gate394inter2, gate394inter3, gate394inter4, gate394inter5, gate394inter6, gate394inter7, gate394inter8, gate394inter9, gate394inter10, gate394inter11, gate394inter12, gate156inter0, gate156inter1, gate156inter2, gate156inter3, gate156inter4, gate156inter5, gate156inter6, gate156inter7, gate156inter8, gate156inter9, gate156inter10, gate156inter11, gate156inter12, gate66inter0, gate66inter1, gate66inter2, gate66inter3, gate66inter4, gate66inter5, gate66inter6, gate66inter7, gate66inter8, gate66inter9, gate66inter10, gate66inter11, gate66inter12, gate64inter0, gate64inter1, gate64inter2, gate64inter3, gate64inter4, gate64inter5, gate64inter6, gate64inter7, gate64inter8, gate64inter9, gate64inter10, gate64inter11, gate64inter12, gate45inter0, gate45inter1, gate45inter2, gate45inter3, gate45inter4, gate45inter5, gate45inter6, gate45inter7, gate45inter8, gate45inter9, gate45inter10, gate45inter11, gate45inter12, gate65inter0, gate65inter1, gate65inter2, gate65inter3, gate65inter4, gate65inter5, gate65inter6, gate65inter7, gate65inter8, gate65inter9, gate65inter10, gate65inter11, gate65inter12, gate114inter0, gate114inter1, gate114inter2, gate114inter3, gate114inter4, gate114inter5, gate114inter6, gate114inter7, gate114inter8, gate114inter9, gate114inter10, gate114inter11, gate114inter12, gate283inter0, gate283inter1, gate283inter2, gate283inter3, gate283inter4, gate283inter5, gate283inter6, gate283inter7, gate283inter8, gate283inter9, gate283inter10, gate283inter11, gate283inter12, gate205inter0, gate205inter1, gate205inter2, gate205inter3, gate205inter4, gate205inter5, gate205inter6, gate205inter7, gate205inter8, gate205inter9, gate205inter10, gate205inter11, gate205inter12, gate504inter0, gate504inter1, gate504inter2, gate504inter3, gate504inter4, gate504inter5, gate504inter6, gate504inter7, gate504inter8, gate504inter9, gate504inter10, gate504inter11, gate504inter12, gate485inter0, gate485inter1, gate485inter2, gate485inter3, gate485inter4, gate485inter5, gate485inter6, gate485inter7, gate485inter8, gate485inter9, gate485inter10, gate485inter11, gate485inter12, gate259inter0, gate259inter1, gate259inter2, gate259inter3, gate259inter4, gate259inter5, gate259inter6, gate259inter7, gate259inter8, gate259inter9, gate259inter10, gate259inter11, gate259inter12, gate112inter0, gate112inter1, gate112inter2, gate112inter3, gate112inter4, gate112inter5, gate112inter6, gate112inter7, gate112inter8, gate112inter9, gate112inter10, gate112inter11, gate112inter12, gate91inter0, gate91inter1, gate91inter2, gate91inter3, gate91inter4, gate91inter5, gate91inter6, gate91inter7, gate91inter8, gate91inter9, gate91inter10, gate91inter11, gate91inter12, gate506inter0, gate506inter1, gate506inter2, gate506inter3, gate506inter4, gate506inter5, gate506inter6, gate506inter7, gate506inter8, gate506inter9, gate506inter10, gate506inter11, gate506inter12, gate251inter0, gate251inter1, gate251inter2, gate251inter3, gate251inter4, gate251inter5, gate251inter6, gate251inter7, gate251inter8, gate251inter9, gate251inter10, gate251inter11, gate251inter12, gate232inter0, gate232inter1, gate232inter2, gate232inter3, gate232inter4, gate232inter5, gate232inter6, gate232inter7, gate232inter8, gate232inter9, gate232inter10, gate232inter11, gate232inter12, gate90inter0, gate90inter1, gate90inter2, gate90inter3, gate90inter4, gate90inter5, gate90inter6, gate90inter7, gate90inter8, gate90inter9, gate90inter10, gate90inter11, gate90inter12, gate287inter0, gate287inter1, gate287inter2, gate287inter3, gate287inter4, gate287inter5, gate287inter6, gate287inter7, gate287inter8, gate287inter9, gate287inter10, gate287inter11, gate287inter12, gate169inter0, gate169inter1, gate169inter2, gate169inter3, gate169inter4, gate169inter5, gate169inter6, gate169inter7, gate169inter8, gate169inter9, gate169inter10, gate169inter11, gate169inter12, gate437inter0, gate437inter1, gate437inter2, gate437inter3, gate437inter4, gate437inter5, gate437inter6, gate437inter7, gate437inter8, gate437inter9, gate437inter10, gate437inter11, gate437inter12, gate39inter0, gate39inter1, gate39inter2, gate39inter3, gate39inter4, gate39inter5, gate39inter6, gate39inter7, gate39inter8, gate39inter9, gate39inter10, gate39inter11, gate39inter12, gate268inter0, gate268inter1, gate268inter2, gate268inter3, gate268inter4, gate268inter5, gate268inter6, gate268inter7, gate268inter8, gate268inter9, gate268inter10, gate268inter11, gate268inter12, gate111inter0, gate111inter1, gate111inter2, gate111inter3, gate111inter4, gate111inter5, gate111inter6, gate111inter7, gate111inter8, gate111inter9, gate111inter10, gate111inter11, gate111inter12, gate435inter0, gate435inter1, gate435inter2, gate435inter3, gate435inter4, gate435inter5, gate435inter6, gate435inter7, gate435inter8, gate435inter9, gate435inter10, gate435inter11, gate435inter12, gate195inter0, gate195inter1, gate195inter2, gate195inter3, gate195inter4, gate195inter5, gate195inter6, gate195inter7, gate195inter8, gate195inter9, gate195inter10, gate195inter11, gate195inter12, gate411inter0, gate411inter1, gate411inter2, gate411inter3, gate411inter4, gate411inter5, gate411inter6, gate411inter7, gate411inter8, gate411inter9, gate411inter10, gate411inter11, gate411inter12, gate514inter0, gate514inter1, gate514inter2, gate514inter3, gate514inter4, gate514inter5, gate514inter6, gate514inter7, gate514inter8, gate514inter9, gate514inter10, gate514inter11, gate514inter12, gate189inter0, gate189inter1, gate189inter2, gate189inter3, gate189inter4, gate189inter5, gate189inter6, gate189inter7, gate189inter8, gate189inter9, gate189inter10, gate189inter11, gate189inter12, gate135inter0, gate135inter1, gate135inter2, gate135inter3, gate135inter4, gate135inter5, gate135inter6, gate135inter7, gate135inter8, gate135inter9, gate135inter10, gate135inter11, gate135inter12, gate237inter0, gate237inter1, gate237inter2, gate237inter3, gate237inter4, gate237inter5, gate237inter6, gate237inter7, gate237inter8, gate237inter9, gate237inter10, gate237inter11, gate237inter12, gate104inter0, gate104inter1, gate104inter2, gate104inter3, gate104inter4, gate104inter5, gate104inter6, gate104inter7, gate104inter8, gate104inter9, gate104inter10, gate104inter11, gate104inter12, gate388inter0, gate388inter1, gate388inter2, gate388inter3, gate388inter4, gate388inter5, gate388inter6, gate388inter7, gate388inter8, gate388inter9, gate388inter10, gate388inter11, gate388inter12, gate36inter0, gate36inter1, gate36inter2, gate36inter3, gate36inter4, gate36inter5, gate36inter6, gate36inter7, gate36inter8, gate36inter9, gate36inter10, gate36inter11, gate36inter12, gate143inter0, gate143inter1, gate143inter2, gate143inter3, gate143inter4, gate143inter5, gate143inter6, gate143inter7, gate143inter8, gate143inter9, gate143inter10, gate143inter11, gate143inter12, gate107inter0, gate107inter1, gate107inter2, gate107inter3, gate107inter4, gate107inter5, gate107inter6, gate107inter7, gate107inter8, gate107inter9, gate107inter10, gate107inter11, gate107inter12, gate480inter0, gate480inter1, gate480inter2, gate480inter3, gate480inter4, gate480inter5, gate480inter6, gate480inter7, gate480inter8, gate480inter9, gate480inter10, gate480inter11, gate480inter12, gate443inter0, gate443inter1, gate443inter2, gate443inter3, gate443inter4, gate443inter5, gate443inter6, gate443inter7, gate443inter8, gate443inter9, gate443inter10, gate443inter11, gate443inter12, gate240inter0, gate240inter1, gate240inter2, gate240inter3, gate240inter4, gate240inter5, gate240inter6, gate240inter7, gate240inter8, gate240inter9, gate240inter10, gate240inter11, gate240inter12, gate257inter0, gate257inter1, gate257inter2, gate257inter3, gate257inter4, gate257inter5, gate257inter6, gate257inter7, gate257inter8, gate257inter9, gate257inter10, gate257inter11, gate257inter12, gate475inter0, gate475inter1, gate475inter2, gate475inter3, gate475inter4, gate475inter5, gate475inter6, gate475inter7, gate475inter8, gate475inter9, gate475inter10, gate475inter11, gate475inter12, gate101inter0, gate101inter1, gate101inter2, gate101inter3, gate101inter4, gate101inter5, gate101inter6, gate101inter7, gate101inter8, gate101inter9, gate101inter10, gate101inter11, gate101inter12, gate30inter0, gate30inter1, gate30inter2, gate30inter3, gate30inter4, gate30inter5, gate30inter6, gate30inter7, gate30inter8, gate30inter9, gate30inter10, gate30inter11, gate30inter12, gate474inter0, gate474inter1, gate474inter2, gate474inter3, gate474inter4, gate474inter5, gate474inter6, gate474inter7, gate474inter8, gate474inter9, gate474inter10, gate474inter11, gate474inter12, gate212inter0, gate212inter1, gate212inter2, gate212inter3, gate212inter4, gate212inter5, gate212inter6, gate212inter7, gate212inter8, gate212inter9, gate212inter10, gate212inter11, gate212inter12, gate223inter0, gate223inter1, gate223inter2, gate223inter3, gate223inter4, gate223inter5, gate223inter6, gate223inter7, gate223inter8, gate223inter9, gate223inter10, gate223inter11, gate223inter12;



and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );
nand2 gate9( .a(G1), .b(G2), .O(G266) );
nand2 gate10( .a(G3), .b(G4), .O(G269) );
nand2 gate11( .a(G5), .b(G6), .O(G272) );
nand2 gate12( .a(G7), .b(G8), .O(G275) );
nand2 gate13( .a(G9), .b(G10), .O(G278) );
nand2 gate14( .a(G11), .b(G12), .O(G281) );
nand2 gate15( .a(G13), .b(G14), .O(G284) );

  xor2  gate799(.a(G16), .b(G15), .O(gate16inter0));
  nand2 gate800(.a(gate16inter0), .b(s_36), .O(gate16inter1));
  and2  gate801(.a(G16), .b(G15), .O(gate16inter2));
  inv1  gate802(.a(s_36), .O(gate16inter3));
  inv1  gate803(.a(s_37), .O(gate16inter4));
  nand2 gate804(.a(gate16inter4), .b(gate16inter3), .O(gate16inter5));
  nor2  gate805(.a(gate16inter5), .b(gate16inter2), .O(gate16inter6));
  inv1  gate806(.a(G15), .O(gate16inter7));
  inv1  gate807(.a(G16), .O(gate16inter8));
  nand2 gate808(.a(gate16inter8), .b(gate16inter7), .O(gate16inter9));
  nand2 gate809(.a(s_37), .b(gate16inter3), .O(gate16inter10));
  nor2  gate810(.a(gate16inter10), .b(gate16inter9), .O(gate16inter11));
  nor2  gate811(.a(gate16inter11), .b(gate16inter6), .O(gate16inter12));
  nand2 gate812(.a(gate16inter12), .b(gate16inter1), .O(G287));
nand2 gate17( .a(G17), .b(G18), .O(G290) );
nand2 gate18( .a(G19), .b(G20), .O(G293) );
nand2 gate19( .a(G21), .b(G22), .O(G296) );
nand2 gate20( .a(G23), .b(G24), .O(G299) );
nand2 gate21( .a(G25), .b(G26), .O(G302) );
nand2 gate22( .a(G27), .b(G28), .O(G305) );
nand2 gate23( .a(G29), .b(G30), .O(G308) );

  xor2  gate1163(.a(G32), .b(G31), .O(gate24inter0));
  nand2 gate1164(.a(gate24inter0), .b(s_88), .O(gate24inter1));
  and2  gate1165(.a(G32), .b(G31), .O(gate24inter2));
  inv1  gate1166(.a(s_88), .O(gate24inter3));
  inv1  gate1167(.a(s_89), .O(gate24inter4));
  nand2 gate1168(.a(gate24inter4), .b(gate24inter3), .O(gate24inter5));
  nor2  gate1169(.a(gate24inter5), .b(gate24inter2), .O(gate24inter6));
  inv1  gate1170(.a(G31), .O(gate24inter7));
  inv1  gate1171(.a(G32), .O(gate24inter8));
  nand2 gate1172(.a(gate24inter8), .b(gate24inter7), .O(gate24inter9));
  nand2 gate1173(.a(s_89), .b(gate24inter3), .O(gate24inter10));
  nor2  gate1174(.a(gate24inter10), .b(gate24inter9), .O(gate24inter11));
  nor2  gate1175(.a(gate24inter11), .b(gate24inter6), .O(gate24inter12));
  nand2 gate1176(.a(gate24inter12), .b(gate24inter1), .O(G311));
nand2 gate25( .a(G1), .b(G5), .O(G314) );
nand2 gate26( .a(G9), .b(G13), .O(G317) );
nand2 gate27( .a(G2), .b(G6), .O(G320) );
nand2 gate28( .a(G10), .b(G14), .O(G323) );

  xor2  gate939(.a(G7), .b(G3), .O(gate29inter0));
  nand2 gate940(.a(gate29inter0), .b(s_56), .O(gate29inter1));
  and2  gate941(.a(G7), .b(G3), .O(gate29inter2));
  inv1  gate942(.a(s_56), .O(gate29inter3));
  inv1  gate943(.a(s_57), .O(gate29inter4));
  nand2 gate944(.a(gate29inter4), .b(gate29inter3), .O(gate29inter5));
  nor2  gate945(.a(gate29inter5), .b(gate29inter2), .O(gate29inter6));
  inv1  gate946(.a(G3), .O(gate29inter7));
  inv1  gate947(.a(G7), .O(gate29inter8));
  nand2 gate948(.a(gate29inter8), .b(gate29inter7), .O(gate29inter9));
  nand2 gate949(.a(s_57), .b(gate29inter3), .O(gate29inter10));
  nor2  gate950(.a(gate29inter10), .b(gate29inter9), .O(gate29inter11));
  nor2  gate951(.a(gate29inter11), .b(gate29inter6), .O(gate29inter12));
  nand2 gate952(.a(gate29inter12), .b(gate29inter1), .O(G326));

  xor2  gate1765(.a(G15), .b(G11), .O(gate30inter0));
  nand2 gate1766(.a(gate30inter0), .b(s_174), .O(gate30inter1));
  and2  gate1767(.a(G15), .b(G11), .O(gate30inter2));
  inv1  gate1768(.a(s_174), .O(gate30inter3));
  inv1  gate1769(.a(s_175), .O(gate30inter4));
  nand2 gate1770(.a(gate30inter4), .b(gate30inter3), .O(gate30inter5));
  nor2  gate1771(.a(gate30inter5), .b(gate30inter2), .O(gate30inter6));
  inv1  gate1772(.a(G11), .O(gate30inter7));
  inv1  gate1773(.a(G15), .O(gate30inter8));
  nand2 gate1774(.a(gate30inter8), .b(gate30inter7), .O(gate30inter9));
  nand2 gate1775(.a(s_175), .b(gate30inter3), .O(gate30inter10));
  nor2  gate1776(.a(gate30inter10), .b(gate30inter9), .O(gate30inter11));
  nor2  gate1777(.a(gate30inter11), .b(gate30inter6), .O(gate30inter12));
  nand2 gate1778(.a(gate30inter12), .b(gate30inter1), .O(G329));
nand2 gate31( .a(G4), .b(G8), .O(G332) );
nand2 gate32( .a(G12), .b(G16), .O(G335) );
nand2 gate33( .a(G17), .b(G21), .O(G338) );
nand2 gate34( .a(G25), .b(G29), .O(G341) );

  xor2  gate1037(.a(G22), .b(G18), .O(gate35inter0));
  nand2 gate1038(.a(gate35inter0), .b(s_70), .O(gate35inter1));
  and2  gate1039(.a(G22), .b(G18), .O(gate35inter2));
  inv1  gate1040(.a(s_70), .O(gate35inter3));
  inv1  gate1041(.a(s_71), .O(gate35inter4));
  nand2 gate1042(.a(gate35inter4), .b(gate35inter3), .O(gate35inter5));
  nor2  gate1043(.a(gate35inter5), .b(gate35inter2), .O(gate35inter6));
  inv1  gate1044(.a(G18), .O(gate35inter7));
  inv1  gate1045(.a(G22), .O(gate35inter8));
  nand2 gate1046(.a(gate35inter8), .b(gate35inter7), .O(gate35inter9));
  nand2 gate1047(.a(s_71), .b(gate35inter3), .O(gate35inter10));
  nor2  gate1048(.a(gate35inter10), .b(gate35inter9), .O(gate35inter11));
  nor2  gate1049(.a(gate35inter11), .b(gate35inter6), .O(gate35inter12));
  nand2 gate1050(.a(gate35inter12), .b(gate35inter1), .O(G344));

  xor2  gate1639(.a(G30), .b(G26), .O(gate36inter0));
  nand2 gate1640(.a(gate36inter0), .b(s_156), .O(gate36inter1));
  and2  gate1641(.a(G30), .b(G26), .O(gate36inter2));
  inv1  gate1642(.a(s_156), .O(gate36inter3));
  inv1  gate1643(.a(s_157), .O(gate36inter4));
  nand2 gate1644(.a(gate36inter4), .b(gate36inter3), .O(gate36inter5));
  nor2  gate1645(.a(gate36inter5), .b(gate36inter2), .O(gate36inter6));
  inv1  gate1646(.a(G26), .O(gate36inter7));
  inv1  gate1647(.a(G30), .O(gate36inter8));
  nand2 gate1648(.a(gate36inter8), .b(gate36inter7), .O(gate36inter9));
  nand2 gate1649(.a(s_157), .b(gate36inter3), .O(gate36inter10));
  nor2  gate1650(.a(gate36inter10), .b(gate36inter9), .O(gate36inter11));
  nor2  gate1651(.a(gate36inter11), .b(gate36inter6), .O(gate36inter12));
  nand2 gate1652(.a(gate36inter12), .b(gate36inter1), .O(G347));
nand2 gate37( .a(G19), .b(G23), .O(G350) );
nand2 gate38( .a(G27), .b(G31), .O(G353) );

  xor2  gate1471(.a(G24), .b(G20), .O(gate39inter0));
  nand2 gate1472(.a(gate39inter0), .b(s_132), .O(gate39inter1));
  and2  gate1473(.a(G24), .b(G20), .O(gate39inter2));
  inv1  gate1474(.a(s_132), .O(gate39inter3));
  inv1  gate1475(.a(s_133), .O(gate39inter4));
  nand2 gate1476(.a(gate39inter4), .b(gate39inter3), .O(gate39inter5));
  nor2  gate1477(.a(gate39inter5), .b(gate39inter2), .O(gate39inter6));
  inv1  gate1478(.a(G20), .O(gate39inter7));
  inv1  gate1479(.a(G24), .O(gate39inter8));
  nand2 gate1480(.a(gate39inter8), .b(gate39inter7), .O(gate39inter9));
  nand2 gate1481(.a(s_133), .b(gate39inter3), .O(gate39inter10));
  nor2  gate1482(.a(gate39inter10), .b(gate39inter9), .O(gate39inter11));
  nor2  gate1483(.a(gate39inter11), .b(gate39inter6), .O(gate39inter12));
  nand2 gate1484(.a(gate39inter12), .b(gate39inter1), .O(G356));

  xor2  gate771(.a(G32), .b(G28), .O(gate40inter0));
  nand2 gate772(.a(gate40inter0), .b(s_32), .O(gate40inter1));
  and2  gate773(.a(G32), .b(G28), .O(gate40inter2));
  inv1  gate774(.a(s_32), .O(gate40inter3));
  inv1  gate775(.a(s_33), .O(gate40inter4));
  nand2 gate776(.a(gate40inter4), .b(gate40inter3), .O(gate40inter5));
  nor2  gate777(.a(gate40inter5), .b(gate40inter2), .O(gate40inter6));
  inv1  gate778(.a(G28), .O(gate40inter7));
  inv1  gate779(.a(G32), .O(gate40inter8));
  nand2 gate780(.a(gate40inter8), .b(gate40inter7), .O(gate40inter9));
  nand2 gate781(.a(s_33), .b(gate40inter3), .O(gate40inter10));
  nor2  gate782(.a(gate40inter10), .b(gate40inter9), .O(gate40inter11));
  nor2  gate783(.a(gate40inter11), .b(gate40inter6), .O(gate40inter12));
  nand2 gate784(.a(gate40inter12), .b(gate40inter1), .O(G359));
nand2 gate41( .a(G1), .b(G266), .O(G362) );
nand2 gate42( .a(G2), .b(G266), .O(G363) );
nand2 gate43( .a(G3), .b(G269), .O(G364) );
nand2 gate44( .a(G4), .b(G269), .O(G365) );

  xor2  gate1233(.a(G272), .b(G5), .O(gate45inter0));
  nand2 gate1234(.a(gate45inter0), .b(s_98), .O(gate45inter1));
  and2  gate1235(.a(G272), .b(G5), .O(gate45inter2));
  inv1  gate1236(.a(s_98), .O(gate45inter3));
  inv1  gate1237(.a(s_99), .O(gate45inter4));
  nand2 gate1238(.a(gate45inter4), .b(gate45inter3), .O(gate45inter5));
  nor2  gate1239(.a(gate45inter5), .b(gate45inter2), .O(gate45inter6));
  inv1  gate1240(.a(G5), .O(gate45inter7));
  inv1  gate1241(.a(G272), .O(gate45inter8));
  nand2 gate1242(.a(gate45inter8), .b(gate45inter7), .O(gate45inter9));
  nand2 gate1243(.a(s_99), .b(gate45inter3), .O(gate45inter10));
  nor2  gate1244(.a(gate45inter10), .b(gate45inter9), .O(gate45inter11));
  nor2  gate1245(.a(gate45inter11), .b(gate45inter6), .O(gate45inter12));
  nand2 gate1246(.a(gate45inter12), .b(gate45inter1), .O(G366));
nand2 gate46( .a(G6), .b(G272), .O(G367) );
nand2 gate47( .a(G7), .b(G275), .O(G368) );
nand2 gate48( .a(G8), .b(G275), .O(G369) );
nand2 gate49( .a(G9), .b(G278), .O(G370) );
nand2 gate50( .a(G10), .b(G278), .O(G371) );

  xor2  gate911(.a(G281), .b(G11), .O(gate51inter0));
  nand2 gate912(.a(gate51inter0), .b(s_52), .O(gate51inter1));
  and2  gate913(.a(G281), .b(G11), .O(gate51inter2));
  inv1  gate914(.a(s_52), .O(gate51inter3));
  inv1  gate915(.a(s_53), .O(gate51inter4));
  nand2 gate916(.a(gate51inter4), .b(gate51inter3), .O(gate51inter5));
  nor2  gate917(.a(gate51inter5), .b(gate51inter2), .O(gate51inter6));
  inv1  gate918(.a(G11), .O(gate51inter7));
  inv1  gate919(.a(G281), .O(gate51inter8));
  nand2 gate920(.a(gate51inter8), .b(gate51inter7), .O(gate51inter9));
  nand2 gate921(.a(s_53), .b(gate51inter3), .O(gate51inter10));
  nor2  gate922(.a(gate51inter10), .b(gate51inter9), .O(gate51inter11));
  nor2  gate923(.a(gate51inter11), .b(gate51inter6), .O(gate51inter12));
  nand2 gate924(.a(gate51inter12), .b(gate51inter1), .O(G372));
nand2 gate52( .a(G12), .b(G281), .O(G373) );
nand2 gate53( .a(G13), .b(G284), .O(G374) );
nand2 gate54( .a(G14), .b(G284), .O(G375) );
nand2 gate55( .a(G15), .b(G287), .O(G376) );

  xor2  gate743(.a(G287), .b(G16), .O(gate56inter0));
  nand2 gate744(.a(gate56inter0), .b(s_28), .O(gate56inter1));
  and2  gate745(.a(G287), .b(G16), .O(gate56inter2));
  inv1  gate746(.a(s_28), .O(gate56inter3));
  inv1  gate747(.a(s_29), .O(gate56inter4));
  nand2 gate748(.a(gate56inter4), .b(gate56inter3), .O(gate56inter5));
  nor2  gate749(.a(gate56inter5), .b(gate56inter2), .O(gate56inter6));
  inv1  gate750(.a(G16), .O(gate56inter7));
  inv1  gate751(.a(G287), .O(gate56inter8));
  nand2 gate752(.a(gate56inter8), .b(gate56inter7), .O(gate56inter9));
  nand2 gate753(.a(s_29), .b(gate56inter3), .O(gate56inter10));
  nor2  gate754(.a(gate56inter10), .b(gate56inter9), .O(gate56inter11));
  nor2  gate755(.a(gate56inter11), .b(gate56inter6), .O(gate56inter12));
  nand2 gate756(.a(gate56inter12), .b(gate56inter1), .O(G377));
nand2 gate57( .a(G17), .b(G290), .O(G378) );
nand2 gate58( .a(G18), .b(G290), .O(G379) );
nand2 gate59( .a(G19), .b(G293), .O(G380) );
nand2 gate60( .a(G20), .b(G293), .O(G381) );
nand2 gate61( .a(G21), .b(G296), .O(G382) );
nand2 gate62( .a(G22), .b(G296), .O(G383) );
nand2 gate63( .a(G23), .b(G299), .O(G384) );

  xor2  gate1219(.a(G299), .b(G24), .O(gate64inter0));
  nand2 gate1220(.a(gate64inter0), .b(s_96), .O(gate64inter1));
  and2  gate1221(.a(G299), .b(G24), .O(gate64inter2));
  inv1  gate1222(.a(s_96), .O(gate64inter3));
  inv1  gate1223(.a(s_97), .O(gate64inter4));
  nand2 gate1224(.a(gate64inter4), .b(gate64inter3), .O(gate64inter5));
  nor2  gate1225(.a(gate64inter5), .b(gate64inter2), .O(gate64inter6));
  inv1  gate1226(.a(G24), .O(gate64inter7));
  inv1  gate1227(.a(G299), .O(gate64inter8));
  nand2 gate1228(.a(gate64inter8), .b(gate64inter7), .O(gate64inter9));
  nand2 gate1229(.a(s_97), .b(gate64inter3), .O(gate64inter10));
  nor2  gate1230(.a(gate64inter10), .b(gate64inter9), .O(gate64inter11));
  nor2  gate1231(.a(gate64inter11), .b(gate64inter6), .O(gate64inter12));
  nand2 gate1232(.a(gate64inter12), .b(gate64inter1), .O(G385));

  xor2  gate1247(.a(G302), .b(G25), .O(gate65inter0));
  nand2 gate1248(.a(gate65inter0), .b(s_100), .O(gate65inter1));
  and2  gate1249(.a(G302), .b(G25), .O(gate65inter2));
  inv1  gate1250(.a(s_100), .O(gate65inter3));
  inv1  gate1251(.a(s_101), .O(gate65inter4));
  nand2 gate1252(.a(gate65inter4), .b(gate65inter3), .O(gate65inter5));
  nor2  gate1253(.a(gate65inter5), .b(gate65inter2), .O(gate65inter6));
  inv1  gate1254(.a(G25), .O(gate65inter7));
  inv1  gate1255(.a(G302), .O(gate65inter8));
  nand2 gate1256(.a(gate65inter8), .b(gate65inter7), .O(gate65inter9));
  nand2 gate1257(.a(s_101), .b(gate65inter3), .O(gate65inter10));
  nor2  gate1258(.a(gate65inter10), .b(gate65inter9), .O(gate65inter11));
  nor2  gate1259(.a(gate65inter11), .b(gate65inter6), .O(gate65inter12));
  nand2 gate1260(.a(gate65inter12), .b(gate65inter1), .O(G386));

  xor2  gate1205(.a(G302), .b(G26), .O(gate66inter0));
  nand2 gate1206(.a(gate66inter0), .b(s_94), .O(gate66inter1));
  and2  gate1207(.a(G302), .b(G26), .O(gate66inter2));
  inv1  gate1208(.a(s_94), .O(gate66inter3));
  inv1  gate1209(.a(s_95), .O(gate66inter4));
  nand2 gate1210(.a(gate66inter4), .b(gate66inter3), .O(gate66inter5));
  nor2  gate1211(.a(gate66inter5), .b(gate66inter2), .O(gate66inter6));
  inv1  gate1212(.a(G26), .O(gate66inter7));
  inv1  gate1213(.a(G302), .O(gate66inter8));
  nand2 gate1214(.a(gate66inter8), .b(gate66inter7), .O(gate66inter9));
  nand2 gate1215(.a(s_95), .b(gate66inter3), .O(gate66inter10));
  nor2  gate1216(.a(gate66inter10), .b(gate66inter9), .O(gate66inter11));
  nor2  gate1217(.a(gate66inter11), .b(gate66inter6), .O(gate66inter12));
  nand2 gate1218(.a(gate66inter12), .b(gate66inter1), .O(G387));
nand2 gate67( .a(G27), .b(G305), .O(G388) );
nand2 gate68( .a(G28), .b(G305), .O(G389) );
nand2 gate69( .a(G29), .b(G308), .O(G390) );
nand2 gate70( .a(G30), .b(G308), .O(G391) );
nand2 gate71( .a(G31), .b(G311), .O(G392) );
nand2 gate72( .a(G32), .b(G311), .O(G393) );
nand2 gate73( .a(G1), .b(G314), .O(G394) );
nand2 gate74( .a(G5), .b(G314), .O(G395) );
nand2 gate75( .a(G9), .b(G317), .O(G396) );
nand2 gate76( .a(G13), .b(G317), .O(G397) );
nand2 gate77( .a(G2), .b(G320), .O(G398) );
nand2 gate78( .a(G6), .b(G320), .O(G399) );
nand2 gate79( .a(G10), .b(G323), .O(G400) );
nand2 gate80( .a(G14), .b(G323), .O(G401) );
nand2 gate81( .a(G3), .b(G326), .O(G402) );
nand2 gate82( .a(G7), .b(G326), .O(G403) );

  xor2  gate617(.a(G329), .b(G11), .O(gate83inter0));
  nand2 gate618(.a(gate83inter0), .b(s_10), .O(gate83inter1));
  and2  gate619(.a(G329), .b(G11), .O(gate83inter2));
  inv1  gate620(.a(s_10), .O(gate83inter3));
  inv1  gate621(.a(s_11), .O(gate83inter4));
  nand2 gate622(.a(gate83inter4), .b(gate83inter3), .O(gate83inter5));
  nor2  gate623(.a(gate83inter5), .b(gate83inter2), .O(gate83inter6));
  inv1  gate624(.a(G11), .O(gate83inter7));
  inv1  gate625(.a(G329), .O(gate83inter8));
  nand2 gate626(.a(gate83inter8), .b(gate83inter7), .O(gate83inter9));
  nand2 gate627(.a(s_11), .b(gate83inter3), .O(gate83inter10));
  nor2  gate628(.a(gate83inter10), .b(gate83inter9), .O(gate83inter11));
  nor2  gate629(.a(gate83inter11), .b(gate83inter6), .O(gate83inter12));
  nand2 gate630(.a(gate83inter12), .b(gate83inter1), .O(G404));
nand2 gate84( .a(G15), .b(G329), .O(G405) );
nand2 gate85( .a(G4), .b(G332), .O(G406) );
nand2 gate86( .a(G8), .b(G332), .O(G407) );
nand2 gate87( .a(G12), .b(G335), .O(G408) );
nand2 gate88( .a(G16), .b(G335), .O(G409) );
nand2 gate89( .a(G17), .b(G338), .O(G410) );

  xor2  gate1415(.a(G338), .b(G21), .O(gate90inter0));
  nand2 gate1416(.a(gate90inter0), .b(s_124), .O(gate90inter1));
  and2  gate1417(.a(G338), .b(G21), .O(gate90inter2));
  inv1  gate1418(.a(s_124), .O(gate90inter3));
  inv1  gate1419(.a(s_125), .O(gate90inter4));
  nand2 gate1420(.a(gate90inter4), .b(gate90inter3), .O(gate90inter5));
  nor2  gate1421(.a(gate90inter5), .b(gate90inter2), .O(gate90inter6));
  inv1  gate1422(.a(G21), .O(gate90inter7));
  inv1  gate1423(.a(G338), .O(gate90inter8));
  nand2 gate1424(.a(gate90inter8), .b(gate90inter7), .O(gate90inter9));
  nand2 gate1425(.a(s_125), .b(gate90inter3), .O(gate90inter10));
  nor2  gate1426(.a(gate90inter10), .b(gate90inter9), .O(gate90inter11));
  nor2  gate1427(.a(gate90inter11), .b(gate90inter6), .O(gate90inter12));
  nand2 gate1428(.a(gate90inter12), .b(gate90inter1), .O(G411));

  xor2  gate1359(.a(G341), .b(G25), .O(gate91inter0));
  nand2 gate1360(.a(gate91inter0), .b(s_116), .O(gate91inter1));
  and2  gate1361(.a(G341), .b(G25), .O(gate91inter2));
  inv1  gate1362(.a(s_116), .O(gate91inter3));
  inv1  gate1363(.a(s_117), .O(gate91inter4));
  nand2 gate1364(.a(gate91inter4), .b(gate91inter3), .O(gate91inter5));
  nor2  gate1365(.a(gate91inter5), .b(gate91inter2), .O(gate91inter6));
  inv1  gate1366(.a(G25), .O(gate91inter7));
  inv1  gate1367(.a(G341), .O(gate91inter8));
  nand2 gate1368(.a(gate91inter8), .b(gate91inter7), .O(gate91inter9));
  nand2 gate1369(.a(s_117), .b(gate91inter3), .O(gate91inter10));
  nor2  gate1370(.a(gate91inter10), .b(gate91inter9), .O(gate91inter11));
  nor2  gate1371(.a(gate91inter11), .b(gate91inter6), .O(gate91inter12));
  nand2 gate1372(.a(gate91inter12), .b(gate91inter1), .O(G412));
nand2 gate92( .a(G29), .b(G341), .O(G413) );
nand2 gate93( .a(G18), .b(G344), .O(G414) );
nand2 gate94( .a(G22), .b(G344), .O(G415) );
nand2 gate95( .a(G26), .b(G347), .O(G416) );
nand2 gate96( .a(G30), .b(G347), .O(G417) );
nand2 gate97( .a(G19), .b(G350), .O(G418) );
nand2 gate98( .a(G23), .b(G350), .O(G419) );
nand2 gate99( .a(G27), .b(G353), .O(G420) );

  xor2  gate813(.a(G353), .b(G31), .O(gate100inter0));
  nand2 gate814(.a(gate100inter0), .b(s_38), .O(gate100inter1));
  and2  gate815(.a(G353), .b(G31), .O(gate100inter2));
  inv1  gate816(.a(s_38), .O(gate100inter3));
  inv1  gate817(.a(s_39), .O(gate100inter4));
  nand2 gate818(.a(gate100inter4), .b(gate100inter3), .O(gate100inter5));
  nor2  gate819(.a(gate100inter5), .b(gate100inter2), .O(gate100inter6));
  inv1  gate820(.a(G31), .O(gate100inter7));
  inv1  gate821(.a(G353), .O(gate100inter8));
  nand2 gate822(.a(gate100inter8), .b(gate100inter7), .O(gate100inter9));
  nand2 gate823(.a(s_39), .b(gate100inter3), .O(gate100inter10));
  nor2  gate824(.a(gate100inter10), .b(gate100inter9), .O(gate100inter11));
  nor2  gate825(.a(gate100inter11), .b(gate100inter6), .O(gate100inter12));
  nand2 gate826(.a(gate100inter12), .b(gate100inter1), .O(G421));

  xor2  gate1751(.a(G356), .b(G20), .O(gate101inter0));
  nand2 gate1752(.a(gate101inter0), .b(s_172), .O(gate101inter1));
  and2  gate1753(.a(G356), .b(G20), .O(gate101inter2));
  inv1  gate1754(.a(s_172), .O(gate101inter3));
  inv1  gate1755(.a(s_173), .O(gate101inter4));
  nand2 gate1756(.a(gate101inter4), .b(gate101inter3), .O(gate101inter5));
  nor2  gate1757(.a(gate101inter5), .b(gate101inter2), .O(gate101inter6));
  inv1  gate1758(.a(G20), .O(gate101inter7));
  inv1  gate1759(.a(G356), .O(gate101inter8));
  nand2 gate1760(.a(gate101inter8), .b(gate101inter7), .O(gate101inter9));
  nand2 gate1761(.a(s_173), .b(gate101inter3), .O(gate101inter10));
  nor2  gate1762(.a(gate101inter10), .b(gate101inter9), .O(gate101inter11));
  nor2  gate1763(.a(gate101inter11), .b(gate101inter6), .O(gate101inter12));
  nand2 gate1764(.a(gate101inter12), .b(gate101inter1), .O(G422));
nand2 gate102( .a(G24), .b(G356), .O(G423) );

  xor2  gate785(.a(G359), .b(G28), .O(gate103inter0));
  nand2 gate786(.a(gate103inter0), .b(s_34), .O(gate103inter1));
  and2  gate787(.a(G359), .b(G28), .O(gate103inter2));
  inv1  gate788(.a(s_34), .O(gate103inter3));
  inv1  gate789(.a(s_35), .O(gate103inter4));
  nand2 gate790(.a(gate103inter4), .b(gate103inter3), .O(gate103inter5));
  nor2  gate791(.a(gate103inter5), .b(gate103inter2), .O(gate103inter6));
  inv1  gate792(.a(G28), .O(gate103inter7));
  inv1  gate793(.a(G359), .O(gate103inter8));
  nand2 gate794(.a(gate103inter8), .b(gate103inter7), .O(gate103inter9));
  nand2 gate795(.a(s_35), .b(gate103inter3), .O(gate103inter10));
  nor2  gate796(.a(gate103inter10), .b(gate103inter9), .O(gate103inter11));
  nor2  gate797(.a(gate103inter11), .b(gate103inter6), .O(gate103inter12));
  nand2 gate798(.a(gate103inter12), .b(gate103inter1), .O(G424));

  xor2  gate1611(.a(G359), .b(G32), .O(gate104inter0));
  nand2 gate1612(.a(gate104inter0), .b(s_152), .O(gate104inter1));
  and2  gate1613(.a(G359), .b(G32), .O(gate104inter2));
  inv1  gate1614(.a(s_152), .O(gate104inter3));
  inv1  gate1615(.a(s_153), .O(gate104inter4));
  nand2 gate1616(.a(gate104inter4), .b(gate104inter3), .O(gate104inter5));
  nor2  gate1617(.a(gate104inter5), .b(gate104inter2), .O(gate104inter6));
  inv1  gate1618(.a(G32), .O(gate104inter7));
  inv1  gate1619(.a(G359), .O(gate104inter8));
  nand2 gate1620(.a(gate104inter8), .b(gate104inter7), .O(gate104inter9));
  nand2 gate1621(.a(s_153), .b(gate104inter3), .O(gate104inter10));
  nor2  gate1622(.a(gate104inter10), .b(gate104inter9), .O(gate104inter11));
  nor2  gate1623(.a(gate104inter11), .b(gate104inter6), .O(gate104inter12));
  nand2 gate1624(.a(gate104inter12), .b(gate104inter1), .O(G425));
nand2 gate105( .a(G362), .b(G363), .O(G426) );
nand2 gate106( .a(G364), .b(G365), .O(G429) );

  xor2  gate1667(.a(G367), .b(G366), .O(gate107inter0));
  nand2 gate1668(.a(gate107inter0), .b(s_160), .O(gate107inter1));
  and2  gate1669(.a(G367), .b(G366), .O(gate107inter2));
  inv1  gate1670(.a(s_160), .O(gate107inter3));
  inv1  gate1671(.a(s_161), .O(gate107inter4));
  nand2 gate1672(.a(gate107inter4), .b(gate107inter3), .O(gate107inter5));
  nor2  gate1673(.a(gate107inter5), .b(gate107inter2), .O(gate107inter6));
  inv1  gate1674(.a(G366), .O(gate107inter7));
  inv1  gate1675(.a(G367), .O(gate107inter8));
  nand2 gate1676(.a(gate107inter8), .b(gate107inter7), .O(gate107inter9));
  nand2 gate1677(.a(s_161), .b(gate107inter3), .O(gate107inter10));
  nor2  gate1678(.a(gate107inter10), .b(gate107inter9), .O(gate107inter11));
  nor2  gate1679(.a(gate107inter11), .b(gate107inter6), .O(gate107inter12));
  nand2 gate1680(.a(gate107inter12), .b(gate107inter1), .O(G432));
nand2 gate108( .a(G368), .b(G369), .O(G435) );
nand2 gate109( .a(G370), .b(G371), .O(G438) );
nand2 gate110( .a(G372), .b(G373), .O(G441) );

  xor2  gate1499(.a(G375), .b(G374), .O(gate111inter0));
  nand2 gate1500(.a(gate111inter0), .b(s_136), .O(gate111inter1));
  and2  gate1501(.a(G375), .b(G374), .O(gate111inter2));
  inv1  gate1502(.a(s_136), .O(gate111inter3));
  inv1  gate1503(.a(s_137), .O(gate111inter4));
  nand2 gate1504(.a(gate111inter4), .b(gate111inter3), .O(gate111inter5));
  nor2  gate1505(.a(gate111inter5), .b(gate111inter2), .O(gate111inter6));
  inv1  gate1506(.a(G374), .O(gate111inter7));
  inv1  gate1507(.a(G375), .O(gate111inter8));
  nand2 gate1508(.a(gate111inter8), .b(gate111inter7), .O(gate111inter9));
  nand2 gate1509(.a(s_137), .b(gate111inter3), .O(gate111inter10));
  nor2  gate1510(.a(gate111inter10), .b(gate111inter9), .O(gate111inter11));
  nor2  gate1511(.a(gate111inter11), .b(gate111inter6), .O(gate111inter12));
  nand2 gate1512(.a(gate111inter12), .b(gate111inter1), .O(G444));

  xor2  gate1345(.a(G377), .b(G376), .O(gate112inter0));
  nand2 gate1346(.a(gate112inter0), .b(s_114), .O(gate112inter1));
  and2  gate1347(.a(G377), .b(G376), .O(gate112inter2));
  inv1  gate1348(.a(s_114), .O(gate112inter3));
  inv1  gate1349(.a(s_115), .O(gate112inter4));
  nand2 gate1350(.a(gate112inter4), .b(gate112inter3), .O(gate112inter5));
  nor2  gate1351(.a(gate112inter5), .b(gate112inter2), .O(gate112inter6));
  inv1  gate1352(.a(G376), .O(gate112inter7));
  inv1  gate1353(.a(G377), .O(gate112inter8));
  nand2 gate1354(.a(gate112inter8), .b(gate112inter7), .O(gate112inter9));
  nand2 gate1355(.a(s_115), .b(gate112inter3), .O(gate112inter10));
  nor2  gate1356(.a(gate112inter10), .b(gate112inter9), .O(gate112inter11));
  nor2  gate1357(.a(gate112inter11), .b(gate112inter6), .O(gate112inter12));
  nand2 gate1358(.a(gate112inter12), .b(gate112inter1), .O(G447));
nand2 gate113( .a(G378), .b(G379), .O(G450) );

  xor2  gate1261(.a(G381), .b(G380), .O(gate114inter0));
  nand2 gate1262(.a(gate114inter0), .b(s_102), .O(gate114inter1));
  and2  gate1263(.a(G381), .b(G380), .O(gate114inter2));
  inv1  gate1264(.a(s_102), .O(gate114inter3));
  inv1  gate1265(.a(s_103), .O(gate114inter4));
  nand2 gate1266(.a(gate114inter4), .b(gate114inter3), .O(gate114inter5));
  nor2  gate1267(.a(gate114inter5), .b(gate114inter2), .O(gate114inter6));
  inv1  gate1268(.a(G380), .O(gate114inter7));
  inv1  gate1269(.a(G381), .O(gate114inter8));
  nand2 gate1270(.a(gate114inter8), .b(gate114inter7), .O(gate114inter9));
  nand2 gate1271(.a(s_103), .b(gate114inter3), .O(gate114inter10));
  nor2  gate1272(.a(gate114inter10), .b(gate114inter9), .O(gate114inter11));
  nor2  gate1273(.a(gate114inter11), .b(gate114inter6), .O(gate114inter12));
  nand2 gate1274(.a(gate114inter12), .b(gate114inter1), .O(G453));
nand2 gate115( .a(G382), .b(G383), .O(G456) );

  xor2  gate897(.a(G385), .b(G384), .O(gate116inter0));
  nand2 gate898(.a(gate116inter0), .b(s_50), .O(gate116inter1));
  and2  gate899(.a(G385), .b(G384), .O(gate116inter2));
  inv1  gate900(.a(s_50), .O(gate116inter3));
  inv1  gate901(.a(s_51), .O(gate116inter4));
  nand2 gate902(.a(gate116inter4), .b(gate116inter3), .O(gate116inter5));
  nor2  gate903(.a(gate116inter5), .b(gate116inter2), .O(gate116inter6));
  inv1  gate904(.a(G384), .O(gate116inter7));
  inv1  gate905(.a(G385), .O(gate116inter8));
  nand2 gate906(.a(gate116inter8), .b(gate116inter7), .O(gate116inter9));
  nand2 gate907(.a(s_51), .b(gate116inter3), .O(gate116inter10));
  nor2  gate908(.a(gate116inter10), .b(gate116inter9), .O(gate116inter11));
  nor2  gate909(.a(gate116inter11), .b(gate116inter6), .O(gate116inter12));
  nand2 gate910(.a(gate116inter12), .b(gate116inter1), .O(G459));
nand2 gate117( .a(G386), .b(G387), .O(G462) );
nand2 gate118( .a(G388), .b(G389), .O(G465) );
nand2 gate119( .a(G390), .b(G391), .O(G468) );
nand2 gate120( .a(G392), .b(G393), .O(G471) );
nand2 gate121( .a(G394), .b(G395), .O(G474) );
nand2 gate122( .a(G396), .b(G397), .O(G477) );

  xor2  gate589(.a(G399), .b(G398), .O(gate123inter0));
  nand2 gate590(.a(gate123inter0), .b(s_6), .O(gate123inter1));
  and2  gate591(.a(G399), .b(G398), .O(gate123inter2));
  inv1  gate592(.a(s_6), .O(gate123inter3));
  inv1  gate593(.a(s_7), .O(gate123inter4));
  nand2 gate594(.a(gate123inter4), .b(gate123inter3), .O(gate123inter5));
  nor2  gate595(.a(gate123inter5), .b(gate123inter2), .O(gate123inter6));
  inv1  gate596(.a(G398), .O(gate123inter7));
  inv1  gate597(.a(G399), .O(gate123inter8));
  nand2 gate598(.a(gate123inter8), .b(gate123inter7), .O(gate123inter9));
  nand2 gate599(.a(s_7), .b(gate123inter3), .O(gate123inter10));
  nor2  gate600(.a(gate123inter10), .b(gate123inter9), .O(gate123inter11));
  nor2  gate601(.a(gate123inter11), .b(gate123inter6), .O(gate123inter12));
  nand2 gate602(.a(gate123inter12), .b(gate123inter1), .O(G480));
nand2 gate124( .a(G400), .b(G401), .O(G483) );
nand2 gate125( .a(G402), .b(G403), .O(G486) );
nand2 gate126( .a(G404), .b(G405), .O(G489) );
nand2 gate127( .a(G406), .b(G407), .O(G492) );

  xor2  gate869(.a(G409), .b(G408), .O(gate128inter0));
  nand2 gate870(.a(gate128inter0), .b(s_46), .O(gate128inter1));
  and2  gate871(.a(G409), .b(G408), .O(gate128inter2));
  inv1  gate872(.a(s_46), .O(gate128inter3));
  inv1  gate873(.a(s_47), .O(gate128inter4));
  nand2 gate874(.a(gate128inter4), .b(gate128inter3), .O(gate128inter5));
  nor2  gate875(.a(gate128inter5), .b(gate128inter2), .O(gate128inter6));
  inv1  gate876(.a(G408), .O(gate128inter7));
  inv1  gate877(.a(G409), .O(gate128inter8));
  nand2 gate878(.a(gate128inter8), .b(gate128inter7), .O(gate128inter9));
  nand2 gate879(.a(s_47), .b(gate128inter3), .O(gate128inter10));
  nor2  gate880(.a(gate128inter10), .b(gate128inter9), .O(gate128inter11));
  nor2  gate881(.a(gate128inter11), .b(gate128inter6), .O(gate128inter12));
  nand2 gate882(.a(gate128inter12), .b(gate128inter1), .O(G495));
nand2 gate129( .a(G410), .b(G411), .O(G498) );
nand2 gate130( .a(G412), .b(G413), .O(G501) );

  xor2  gate1107(.a(G415), .b(G414), .O(gate131inter0));
  nand2 gate1108(.a(gate131inter0), .b(s_80), .O(gate131inter1));
  and2  gate1109(.a(G415), .b(G414), .O(gate131inter2));
  inv1  gate1110(.a(s_80), .O(gate131inter3));
  inv1  gate1111(.a(s_81), .O(gate131inter4));
  nand2 gate1112(.a(gate131inter4), .b(gate131inter3), .O(gate131inter5));
  nor2  gate1113(.a(gate131inter5), .b(gate131inter2), .O(gate131inter6));
  inv1  gate1114(.a(G414), .O(gate131inter7));
  inv1  gate1115(.a(G415), .O(gate131inter8));
  nand2 gate1116(.a(gate131inter8), .b(gate131inter7), .O(gate131inter9));
  nand2 gate1117(.a(s_81), .b(gate131inter3), .O(gate131inter10));
  nor2  gate1118(.a(gate131inter10), .b(gate131inter9), .O(gate131inter11));
  nor2  gate1119(.a(gate131inter11), .b(gate131inter6), .O(gate131inter12));
  nand2 gate1120(.a(gate131inter12), .b(gate131inter1), .O(G504));

  xor2  gate995(.a(G417), .b(G416), .O(gate132inter0));
  nand2 gate996(.a(gate132inter0), .b(s_64), .O(gate132inter1));
  and2  gate997(.a(G417), .b(G416), .O(gate132inter2));
  inv1  gate998(.a(s_64), .O(gate132inter3));
  inv1  gate999(.a(s_65), .O(gate132inter4));
  nand2 gate1000(.a(gate132inter4), .b(gate132inter3), .O(gate132inter5));
  nor2  gate1001(.a(gate132inter5), .b(gate132inter2), .O(gate132inter6));
  inv1  gate1002(.a(G416), .O(gate132inter7));
  inv1  gate1003(.a(G417), .O(gate132inter8));
  nand2 gate1004(.a(gate132inter8), .b(gate132inter7), .O(gate132inter9));
  nand2 gate1005(.a(s_65), .b(gate132inter3), .O(gate132inter10));
  nor2  gate1006(.a(gate132inter10), .b(gate132inter9), .O(gate132inter11));
  nor2  gate1007(.a(gate132inter11), .b(gate132inter6), .O(gate132inter12));
  nand2 gate1008(.a(gate132inter12), .b(gate132inter1), .O(G507));

  xor2  gate1065(.a(G419), .b(G418), .O(gate133inter0));
  nand2 gate1066(.a(gate133inter0), .b(s_74), .O(gate133inter1));
  and2  gate1067(.a(G419), .b(G418), .O(gate133inter2));
  inv1  gate1068(.a(s_74), .O(gate133inter3));
  inv1  gate1069(.a(s_75), .O(gate133inter4));
  nand2 gate1070(.a(gate133inter4), .b(gate133inter3), .O(gate133inter5));
  nor2  gate1071(.a(gate133inter5), .b(gate133inter2), .O(gate133inter6));
  inv1  gate1072(.a(G418), .O(gate133inter7));
  inv1  gate1073(.a(G419), .O(gate133inter8));
  nand2 gate1074(.a(gate133inter8), .b(gate133inter7), .O(gate133inter9));
  nand2 gate1075(.a(s_75), .b(gate133inter3), .O(gate133inter10));
  nor2  gate1076(.a(gate133inter10), .b(gate133inter9), .O(gate133inter11));
  nor2  gate1077(.a(gate133inter11), .b(gate133inter6), .O(gate133inter12));
  nand2 gate1078(.a(gate133inter12), .b(gate133inter1), .O(G510));
nand2 gate134( .a(G420), .b(G421), .O(G513) );

  xor2  gate1583(.a(G423), .b(G422), .O(gate135inter0));
  nand2 gate1584(.a(gate135inter0), .b(s_148), .O(gate135inter1));
  and2  gate1585(.a(G423), .b(G422), .O(gate135inter2));
  inv1  gate1586(.a(s_148), .O(gate135inter3));
  inv1  gate1587(.a(s_149), .O(gate135inter4));
  nand2 gate1588(.a(gate135inter4), .b(gate135inter3), .O(gate135inter5));
  nor2  gate1589(.a(gate135inter5), .b(gate135inter2), .O(gate135inter6));
  inv1  gate1590(.a(G422), .O(gate135inter7));
  inv1  gate1591(.a(G423), .O(gate135inter8));
  nand2 gate1592(.a(gate135inter8), .b(gate135inter7), .O(gate135inter9));
  nand2 gate1593(.a(s_149), .b(gate135inter3), .O(gate135inter10));
  nor2  gate1594(.a(gate135inter10), .b(gate135inter9), .O(gate135inter11));
  nor2  gate1595(.a(gate135inter11), .b(gate135inter6), .O(gate135inter12));
  nand2 gate1596(.a(gate135inter12), .b(gate135inter1), .O(G516));
nand2 gate136( .a(G424), .b(G425), .O(G519) );
nand2 gate137( .a(G426), .b(G429), .O(G522) );
nand2 gate138( .a(G432), .b(G435), .O(G525) );
nand2 gate139( .a(G438), .b(G441), .O(G528) );
nand2 gate140( .a(G444), .b(G447), .O(G531) );
nand2 gate141( .a(G450), .b(G453), .O(G534) );
nand2 gate142( .a(G456), .b(G459), .O(G537) );

  xor2  gate1653(.a(G465), .b(G462), .O(gate143inter0));
  nand2 gate1654(.a(gate143inter0), .b(s_158), .O(gate143inter1));
  and2  gate1655(.a(G465), .b(G462), .O(gate143inter2));
  inv1  gate1656(.a(s_158), .O(gate143inter3));
  inv1  gate1657(.a(s_159), .O(gate143inter4));
  nand2 gate1658(.a(gate143inter4), .b(gate143inter3), .O(gate143inter5));
  nor2  gate1659(.a(gate143inter5), .b(gate143inter2), .O(gate143inter6));
  inv1  gate1660(.a(G462), .O(gate143inter7));
  inv1  gate1661(.a(G465), .O(gate143inter8));
  nand2 gate1662(.a(gate143inter8), .b(gate143inter7), .O(gate143inter9));
  nand2 gate1663(.a(s_159), .b(gate143inter3), .O(gate143inter10));
  nor2  gate1664(.a(gate143inter10), .b(gate143inter9), .O(gate143inter11));
  nor2  gate1665(.a(gate143inter11), .b(gate143inter6), .O(gate143inter12));
  nand2 gate1666(.a(gate143inter12), .b(gate143inter1), .O(G540));
nand2 gate144( .a(G468), .b(G471), .O(G543) );
nand2 gate145( .a(G474), .b(G477), .O(G546) );
nand2 gate146( .a(G480), .b(G483), .O(G549) );
nand2 gate147( .a(G486), .b(G489), .O(G552) );
nand2 gate148( .a(G492), .b(G495), .O(G555) );
nand2 gate149( .a(G498), .b(G501), .O(G558) );
nand2 gate150( .a(G504), .b(G507), .O(G561) );
nand2 gate151( .a(G510), .b(G513), .O(G564) );
nand2 gate152( .a(G516), .b(G519), .O(G567) );
nand2 gate153( .a(G426), .b(G522), .O(G570) );
nand2 gate154( .a(G429), .b(G522), .O(G571) );
nand2 gate155( .a(G432), .b(G525), .O(G572) );

  xor2  gate1191(.a(G525), .b(G435), .O(gate156inter0));
  nand2 gate1192(.a(gate156inter0), .b(s_92), .O(gate156inter1));
  and2  gate1193(.a(G525), .b(G435), .O(gate156inter2));
  inv1  gate1194(.a(s_92), .O(gate156inter3));
  inv1  gate1195(.a(s_93), .O(gate156inter4));
  nand2 gate1196(.a(gate156inter4), .b(gate156inter3), .O(gate156inter5));
  nor2  gate1197(.a(gate156inter5), .b(gate156inter2), .O(gate156inter6));
  inv1  gate1198(.a(G435), .O(gate156inter7));
  inv1  gate1199(.a(G525), .O(gate156inter8));
  nand2 gate1200(.a(gate156inter8), .b(gate156inter7), .O(gate156inter9));
  nand2 gate1201(.a(s_93), .b(gate156inter3), .O(gate156inter10));
  nor2  gate1202(.a(gate156inter10), .b(gate156inter9), .O(gate156inter11));
  nor2  gate1203(.a(gate156inter11), .b(gate156inter6), .O(gate156inter12));
  nand2 gate1204(.a(gate156inter12), .b(gate156inter1), .O(G573));
nand2 gate157( .a(G438), .b(G528), .O(G574) );
nand2 gate158( .a(G441), .b(G528), .O(G575) );
nand2 gate159( .a(G444), .b(G531), .O(G576) );
nand2 gate160( .a(G447), .b(G531), .O(G577) );
nand2 gate161( .a(G450), .b(G534), .O(G578) );
nand2 gate162( .a(G453), .b(G534), .O(G579) );
nand2 gate163( .a(G456), .b(G537), .O(G580) );
nand2 gate164( .a(G459), .b(G537), .O(G581) );
nand2 gate165( .a(G462), .b(G540), .O(G582) );
nand2 gate166( .a(G465), .b(G540), .O(G583) );
nand2 gate167( .a(G468), .b(G543), .O(G584) );
nand2 gate168( .a(G471), .b(G543), .O(G585) );

  xor2  gate1443(.a(G546), .b(G474), .O(gate169inter0));
  nand2 gate1444(.a(gate169inter0), .b(s_128), .O(gate169inter1));
  and2  gate1445(.a(G546), .b(G474), .O(gate169inter2));
  inv1  gate1446(.a(s_128), .O(gate169inter3));
  inv1  gate1447(.a(s_129), .O(gate169inter4));
  nand2 gate1448(.a(gate169inter4), .b(gate169inter3), .O(gate169inter5));
  nor2  gate1449(.a(gate169inter5), .b(gate169inter2), .O(gate169inter6));
  inv1  gate1450(.a(G474), .O(gate169inter7));
  inv1  gate1451(.a(G546), .O(gate169inter8));
  nand2 gate1452(.a(gate169inter8), .b(gate169inter7), .O(gate169inter9));
  nand2 gate1453(.a(s_129), .b(gate169inter3), .O(gate169inter10));
  nor2  gate1454(.a(gate169inter10), .b(gate169inter9), .O(gate169inter11));
  nor2  gate1455(.a(gate169inter11), .b(gate169inter6), .O(gate169inter12));
  nand2 gate1456(.a(gate169inter12), .b(gate169inter1), .O(G586));
nand2 gate170( .a(G477), .b(G546), .O(G587) );
nand2 gate171( .a(G480), .b(G549), .O(G588) );
nand2 gate172( .a(G483), .b(G549), .O(G589) );
nand2 gate173( .a(G486), .b(G552), .O(G590) );
nand2 gate174( .a(G489), .b(G552), .O(G591) );
nand2 gate175( .a(G492), .b(G555), .O(G592) );
nand2 gate176( .a(G495), .b(G555), .O(G593) );
nand2 gate177( .a(G498), .b(G558), .O(G594) );
nand2 gate178( .a(G501), .b(G558), .O(G595) );
nand2 gate179( .a(G504), .b(G561), .O(G596) );
nand2 gate180( .a(G507), .b(G561), .O(G597) );
nand2 gate181( .a(G510), .b(G564), .O(G598) );
nand2 gate182( .a(G513), .b(G564), .O(G599) );
nand2 gate183( .a(G516), .b(G567), .O(G600) );
nand2 gate184( .a(G519), .b(G567), .O(G601) );
nand2 gate185( .a(G570), .b(G571), .O(G602) );

  xor2  gate575(.a(G573), .b(G572), .O(gate186inter0));
  nand2 gate576(.a(gate186inter0), .b(s_4), .O(gate186inter1));
  and2  gate577(.a(G573), .b(G572), .O(gate186inter2));
  inv1  gate578(.a(s_4), .O(gate186inter3));
  inv1  gate579(.a(s_5), .O(gate186inter4));
  nand2 gate580(.a(gate186inter4), .b(gate186inter3), .O(gate186inter5));
  nor2  gate581(.a(gate186inter5), .b(gate186inter2), .O(gate186inter6));
  inv1  gate582(.a(G572), .O(gate186inter7));
  inv1  gate583(.a(G573), .O(gate186inter8));
  nand2 gate584(.a(gate186inter8), .b(gate186inter7), .O(gate186inter9));
  nand2 gate585(.a(s_5), .b(gate186inter3), .O(gate186inter10));
  nor2  gate586(.a(gate186inter10), .b(gate186inter9), .O(gate186inter11));
  nor2  gate587(.a(gate186inter11), .b(gate186inter6), .O(gate186inter12));
  nand2 gate588(.a(gate186inter12), .b(gate186inter1), .O(G607));
nand2 gate187( .a(G574), .b(G575), .O(G612) );

  xor2  gate981(.a(G577), .b(G576), .O(gate188inter0));
  nand2 gate982(.a(gate188inter0), .b(s_62), .O(gate188inter1));
  and2  gate983(.a(G577), .b(G576), .O(gate188inter2));
  inv1  gate984(.a(s_62), .O(gate188inter3));
  inv1  gate985(.a(s_63), .O(gate188inter4));
  nand2 gate986(.a(gate188inter4), .b(gate188inter3), .O(gate188inter5));
  nor2  gate987(.a(gate188inter5), .b(gate188inter2), .O(gate188inter6));
  inv1  gate988(.a(G576), .O(gate188inter7));
  inv1  gate989(.a(G577), .O(gate188inter8));
  nand2 gate990(.a(gate188inter8), .b(gate188inter7), .O(gate188inter9));
  nand2 gate991(.a(s_63), .b(gate188inter3), .O(gate188inter10));
  nor2  gate992(.a(gate188inter10), .b(gate188inter9), .O(gate188inter11));
  nor2  gate993(.a(gate188inter11), .b(gate188inter6), .O(gate188inter12));
  nand2 gate994(.a(gate188inter12), .b(gate188inter1), .O(G617));

  xor2  gate1569(.a(G579), .b(G578), .O(gate189inter0));
  nand2 gate1570(.a(gate189inter0), .b(s_146), .O(gate189inter1));
  and2  gate1571(.a(G579), .b(G578), .O(gate189inter2));
  inv1  gate1572(.a(s_146), .O(gate189inter3));
  inv1  gate1573(.a(s_147), .O(gate189inter4));
  nand2 gate1574(.a(gate189inter4), .b(gate189inter3), .O(gate189inter5));
  nor2  gate1575(.a(gate189inter5), .b(gate189inter2), .O(gate189inter6));
  inv1  gate1576(.a(G578), .O(gate189inter7));
  inv1  gate1577(.a(G579), .O(gate189inter8));
  nand2 gate1578(.a(gate189inter8), .b(gate189inter7), .O(gate189inter9));
  nand2 gate1579(.a(s_147), .b(gate189inter3), .O(gate189inter10));
  nor2  gate1580(.a(gate189inter10), .b(gate189inter9), .O(gate189inter11));
  nor2  gate1581(.a(gate189inter11), .b(gate189inter6), .O(gate189inter12));
  nand2 gate1582(.a(gate189inter12), .b(gate189inter1), .O(G622));
nand2 gate190( .a(G580), .b(G581), .O(G627) );
nand2 gate191( .a(G582), .b(G583), .O(G632) );
nand2 gate192( .a(G584), .b(G585), .O(G637) );
nand2 gate193( .a(G586), .b(G587), .O(G642) );
nand2 gate194( .a(G588), .b(G589), .O(G645) );

  xor2  gate1527(.a(G591), .b(G590), .O(gate195inter0));
  nand2 gate1528(.a(gate195inter0), .b(s_140), .O(gate195inter1));
  and2  gate1529(.a(G591), .b(G590), .O(gate195inter2));
  inv1  gate1530(.a(s_140), .O(gate195inter3));
  inv1  gate1531(.a(s_141), .O(gate195inter4));
  nand2 gate1532(.a(gate195inter4), .b(gate195inter3), .O(gate195inter5));
  nor2  gate1533(.a(gate195inter5), .b(gate195inter2), .O(gate195inter6));
  inv1  gate1534(.a(G590), .O(gate195inter7));
  inv1  gate1535(.a(G591), .O(gate195inter8));
  nand2 gate1536(.a(gate195inter8), .b(gate195inter7), .O(gate195inter9));
  nand2 gate1537(.a(s_141), .b(gate195inter3), .O(gate195inter10));
  nor2  gate1538(.a(gate195inter10), .b(gate195inter9), .O(gate195inter11));
  nor2  gate1539(.a(gate195inter11), .b(gate195inter6), .O(gate195inter12));
  nand2 gate1540(.a(gate195inter12), .b(gate195inter1), .O(G648));

  xor2  gate631(.a(G593), .b(G592), .O(gate196inter0));
  nand2 gate632(.a(gate196inter0), .b(s_12), .O(gate196inter1));
  and2  gate633(.a(G593), .b(G592), .O(gate196inter2));
  inv1  gate634(.a(s_12), .O(gate196inter3));
  inv1  gate635(.a(s_13), .O(gate196inter4));
  nand2 gate636(.a(gate196inter4), .b(gate196inter3), .O(gate196inter5));
  nor2  gate637(.a(gate196inter5), .b(gate196inter2), .O(gate196inter6));
  inv1  gate638(.a(G592), .O(gate196inter7));
  inv1  gate639(.a(G593), .O(gate196inter8));
  nand2 gate640(.a(gate196inter8), .b(gate196inter7), .O(gate196inter9));
  nand2 gate641(.a(s_13), .b(gate196inter3), .O(gate196inter10));
  nor2  gate642(.a(gate196inter10), .b(gate196inter9), .O(gate196inter11));
  nor2  gate643(.a(gate196inter11), .b(gate196inter6), .O(gate196inter12));
  nand2 gate644(.a(gate196inter12), .b(gate196inter1), .O(G651));
nand2 gate197( .a(G594), .b(G595), .O(G654) );

  xor2  gate1009(.a(G597), .b(G596), .O(gate198inter0));
  nand2 gate1010(.a(gate198inter0), .b(s_66), .O(gate198inter1));
  and2  gate1011(.a(G597), .b(G596), .O(gate198inter2));
  inv1  gate1012(.a(s_66), .O(gate198inter3));
  inv1  gate1013(.a(s_67), .O(gate198inter4));
  nand2 gate1014(.a(gate198inter4), .b(gate198inter3), .O(gate198inter5));
  nor2  gate1015(.a(gate198inter5), .b(gate198inter2), .O(gate198inter6));
  inv1  gate1016(.a(G596), .O(gate198inter7));
  inv1  gate1017(.a(G597), .O(gate198inter8));
  nand2 gate1018(.a(gate198inter8), .b(gate198inter7), .O(gate198inter9));
  nand2 gate1019(.a(s_67), .b(gate198inter3), .O(gate198inter10));
  nor2  gate1020(.a(gate198inter10), .b(gate198inter9), .O(gate198inter11));
  nor2  gate1021(.a(gate198inter11), .b(gate198inter6), .O(gate198inter12));
  nand2 gate1022(.a(gate198inter12), .b(gate198inter1), .O(G657));
nand2 gate199( .a(G598), .b(G599), .O(G660) );
nand2 gate200( .a(G600), .b(G601), .O(G663) );
nand2 gate201( .a(G602), .b(G607), .O(G666) );
nand2 gate202( .a(G612), .b(G617), .O(G669) );
nand2 gate203( .a(G602), .b(G612), .O(G672) );
nand2 gate204( .a(G607), .b(G617), .O(G675) );

  xor2  gate1289(.a(G627), .b(G622), .O(gate205inter0));
  nand2 gate1290(.a(gate205inter0), .b(s_106), .O(gate205inter1));
  and2  gate1291(.a(G627), .b(G622), .O(gate205inter2));
  inv1  gate1292(.a(s_106), .O(gate205inter3));
  inv1  gate1293(.a(s_107), .O(gate205inter4));
  nand2 gate1294(.a(gate205inter4), .b(gate205inter3), .O(gate205inter5));
  nor2  gate1295(.a(gate205inter5), .b(gate205inter2), .O(gate205inter6));
  inv1  gate1296(.a(G622), .O(gate205inter7));
  inv1  gate1297(.a(G627), .O(gate205inter8));
  nand2 gate1298(.a(gate205inter8), .b(gate205inter7), .O(gate205inter9));
  nand2 gate1299(.a(s_107), .b(gate205inter3), .O(gate205inter10));
  nor2  gate1300(.a(gate205inter10), .b(gate205inter9), .O(gate205inter11));
  nor2  gate1301(.a(gate205inter11), .b(gate205inter6), .O(gate205inter12));
  nand2 gate1302(.a(gate205inter12), .b(gate205inter1), .O(G678));

  xor2  gate603(.a(G637), .b(G632), .O(gate206inter0));
  nand2 gate604(.a(gate206inter0), .b(s_8), .O(gate206inter1));
  and2  gate605(.a(G637), .b(G632), .O(gate206inter2));
  inv1  gate606(.a(s_8), .O(gate206inter3));
  inv1  gate607(.a(s_9), .O(gate206inter4));
  nand2 gate608(.a(gate206inter4), .b(gate206inter3), .O(gate206inter5));
  nor2  gate609(.a(gate206inter5), .b(gate206inter2), .O(gate206inter6));
  inv1  gate610(.a(G632), .O(gate206inter7));
  inv1  gate611(.a(G637), .O(gate206inter8));
  nand2 gate612(.a(gate206inter8), .b(gate206inter7), .O(gate206inter9));
  nand2 gate613(.a(s_9), .b(gate206inter3), .O(gate206inter10));
  nor2  gate614(.a(gate206inter10), .b(gate206inter9), .O(gate206inter11));
  nor2  gate615(.a(gate206inter11), .b(gate206inter6), .O(gate206inter12));
  nand2 gate616(.a(gate206inter12), .b(gate206inter1), .O(G681));
nand2 gate207( .a(G622), .b(G632), .O(G684) );
nand2 gate208( .a(G627), .b(G637), .O(G687) );
nand2 gate209( .a(G602), .b(G666), .O(G690) );
nand2 gate210( .a(G607), .b(G666), .O(G691) );
nand2 gate211( .a(G612), .b(G669), .O(G692) );

  xor2  gate1793(.a(G669), .b(G617), .O(gate212inter0));
  nand2 gate1794(.a(gate212inter0), .b(s_178), .O(gate212inter1));
  and2  gate1795(.a(G669), .b(G617), .O(gate212inter2));
  inv1  gate1796(.a(s_178), .O(gate212inter3));
  inv1  gate1797(.a(s_179), .O(gate212inter4));
  nand2 gate1798(.a(gate212inter4), .b(gate212inter3), .O(gate212inter5));
  nor2  gate1799(.a(gate212inter5), .b(gate212inter2), .O(gate212inter6));
  inv1  gate1800(.a(G617), .O(gate212inter7));
  inv1  gate1801(.a(G669), .O(gate212inter8));
  nand2 gate1802(.a(gate212inter8), .b(gate212inter7), .O(gate212inter9));
  nand2 gate1803(.a(s_179), .b(gate212inter3), .O(gate212inter10));
  nor2  gate1804(.a(gate212inter10), .b(gate212inter9), .O(gate212inter11));
  nor2  gate1805(.a(gate212inter11), .b(gate212inter6), .O(gate212inter12));
  nand2 gate1806(.a(gate212inter12), .b(gate212inter1), .O(G693));
nand2 gate213( .a(G602), .b(G672), .O(G694) );
nand2 gate214( .a(G612), .b(G672), .O(G695) );
nand2 gate215( .a(G607), .b(G675), .O(G696) );

  xor2  gate1079(.a(G675), .b(G617), .O(gate216inter0));
  nand2 gate1080(.a(gate216inter0), .b(s_76), .O(gate216inter1));
  and2  gate1081(.a(G675), .b(G617), .O(gate216inter2));
  inv1  gate1082(.a(s_76), .O(gate216inter3));
  inv1  gate1083(.a(s_77), .O(gate216inter4));
  nand2 gate1084(.a(gate216inter4), .b(gate216inter3), .O(gate216inter5));
  nor2  gate1085(.a(gate216inter5), .b(gate216inter2), .O(gate216inter6));
  inv1  gate1086(.a(G617), .O(gate216inter7));
  inv1  gate1087(.a(G675), .O(gate216inter8));
  nand2 gate1088(.a(gate216inter8), .b(gate216inter7), .O(gate216inter9));
  nand2 gate1089(.a(s_77), .b(gate216inter3), .O(gate216inter10));
  nor2  gate1090(.a(gate216inter10), .b(gate216inter9), .O(gate216inter11));
  nor2  gate1091(.a(gate216inter11), .b(gate216inter6), .O(gate216inter12));
  nand2 gate1092(.a(gate216inter12), .b(gate216inter1), .O(G697));
nand2 gate217( .a(G622), .b(G678), .O(G698) );
nand2 gate218( .a(G627), .b(G678), .O(G699) );
nand2 gate219( .a(G632), .b(G681), .O(G700) );
nand2 gate220( .a(G637), .b(G681), .O(G701) );
nand2 gate221( .a(G622), .b(G684), .O(G702) );
nand2 gate222( .a(G632), .b(G684), .O(G703) );

  xor2  gate1807(.a(G687), .b(G627), .O(gate223inter0));
  nand2 gate1808(.a(gate223inter0), .b(s_180), .O(gate223inter1));
  and2  gate1809(.a(G687), .b(G627), .O(gate223inter2));
  inv1  gate1810(.a(s_180), .O(gate223inter3));
  inv1  gate1811(.a(s_181), .O(gate223inter4));
  nand2 gate1812(.a(gate223inter4), .b(gate223inter3), .O(gate223inter5));
  nor2  gate1813(.a(gate223inter5), .b(gate223inter2), .O(gate223inter6));
  inv1  gate1814(.a(G627), .O(gate223inter7));
  inv1  gate1815(.a(G687), .O(gate223inter8));
  nand2 gate1816(.a(gate223inter8), .b(gate223inter7), .O(gate223inter9));
  nand2 gate1817(.a(s_181), .b(gate223inter3), .O(gate223inter10));
  nor2  gate1818(.a(gate223inter10), .b(gate223inter9), .O(gate223inter11));
  nor2  gate1819(.a(gate223inter11), .b(gate223inter6), .O(gate223inter12));
  nand2 gate1820(.a(gate223inter12), .b(gate223inter1), .O(G704));
nand2 gate224( .a(G637), .b(G687), .O(G705) );
nand2 gate225( .a(G690), .b(G691), .O(G706) );

  xor2  gate715(.a(G693), .b(G692), .O(gate226inter0));
  nand2 gate716(.a(gate226inter0), .b(s_24), .O(gate226inter1));
  and2  gate717(.a(G693), .b(G692), .O(gate226inter2));
  inv1  gate718(.a(s_24), .O(gate226inter3));
  inv1  gate719(.a(s_25), .O(gate226inter4));
  nand2 gate720(.a(gate226inter4), .b(gate226inter3), .O(gate226inter5));
  nor2  gate721(.a(gate226inter5), .b(gate226inter2), .O(gate226inter6));
  inv1  gate722(.a(G692), .O(gate226inter7));
  inv1  gate723(.a(G693), .O(gate226inter8));
  nand2 gate724(.a(gate226inter8), .b(gate226inter7), .O(gate226inter9));
  nand2 gate725(.a(s_25), .b(gate226inter3), .O(gate226inter10));
  nor2  gate726(.a(gate226inter10), .b(gate226inter9), .O(gate226inter11));
  nor2  gate727(.a(gate226inter11), .b(gate226inter6), .O(gate226inter12));
  nand2 gate728(.a(gate226inter12), .b(gate226inter1), .O(G709));
nand2 gate227( .a(G694), .b(G695), .O(G712) );
nand2 gate228( .a(G696), .b(G697), .O(G715) );
nand2 gate229( .a(G698), .b(G699), .O(G718) );
nand2 gate230( .a(G700), .b(G701), .O(G721) );
nand2 gate231( .a(G702), .b(G703), .O(G724) );

  xor2  gate1401(.a(G705), .b(G704), .O(gate232inter0));
  nand2 gate1402(.a(gate232inter0), .b(s_122), .O(gate232inter1));
  and2  gate1403(.a(G705), .b(G704), .O(gate232inter2));
  inv1  gate1404(.a(s_122), .O(gate232inter3));
  inv1  gate1405(.a(s_123), .O(gate232inter4));
  nand2 gate1406(.a(gate232inter4), .b(gate232inter3), .O(gate232inter5));
  nor2  gate1407(.a(gate232inter5), .b(gate232inter2), .O(gate232inter6));
  inv1  gate1408(.a(G704), .O(gate232inter7));
  inv1  gate1409(.a(G705), .O(gate232inter8));
  nand2 gate1410(.a(gate232inter8), .b(gate232inter7), .O(gate232inter9));
  nand2 gate1411(.a(s_123), .b(gate232inter3), .O(gate232inter10));
  nor2  gate1412(.a(gate232inter10), .b(gate232inter9), .O(gate232inter11));
  nor2  gate1413(.a(gate232inter11), .b(gate232inter6), .O(gate232inter12));
  nand2 gate1414(.a(gate232inter12), .b(gate232inter1), .O(G727));
nand2 gate233( .a(G242), .b(G718), .O(G730) );
nand2 gate234( .a(G245), .b(G721), .O(G733) );
nand2 gate235( .a(G248), .b(G724), .O(G736) );

  xor2  gate841(.a(G727), .b(G251), .O(gate236inter0));
  nand2 gate842(.a(gate236inter0), .b(s_42), .O(gate236inter1));
  and2  gate843(.a(G727), .b(G251), .O(gate236inter2));
  inv1  gate844(.a(s_42), .O(gate236inter3));
  inv1  gate845(.a(s_43), .O(gate236inter4));
  nand2 gate846(.a(gate236inter4), .b(gate236inter3), .O(gate236inter5));
  nor2  gate847(.a(gate236inter5), .b(gate236inter2), .O(gate236inter6));
  inv1  gate848(.a(G251), .O(gate236inter7));
  inv1  gate849(.a(G727), .O(gate236inter8));
  nand2 gate850(.a(gate236inter8), .b(gate236inter7), .O(gate236inter9));
  nand2 gate851(.a(s_43), .b(gate236inter3), .O(gate236inter10));
  nor2  gate852(.a(gate236inter10), .b(gate236inter9), .O(gate236inter11));
  nor2  gate853(.a(gate236inter11), .b(gate236inter6), .O(gate236inter12));
  nand2 gate854(.a(gate236inter12), .b(gate236inter1), .O(G739));

  xor2  gate1597(.a(G706), .b(G254), .O(gate237inter0));
  nand2 gate1598(.a(gate237inter0), .b(s_150), .O(gate237inter1));
  and2  gate1599(.a(G706), .b(G254), .O(gate237inter2));
  inv1  gate1600(.a(s_150), .O(gate237inter3));
  inv1  gate1601(.a(s_151), .O(gate237inter4));
  nand2 gate1602(.a(gate237inter4), .b(gate237inter3), .O(gate237inter5));
  nor2  gate1603(.a(gate237inter5), .b(gate237inter2), .O(gate237inter6));
  inv1  gate1604(.a(G254), .O(gate237inter7));
  inv1  gate1605(.a(G706), .O(gate237inter8));
  nand2 gate1606(.a(gate237inter8), .b(gate237inter7), .O(gate237inter9));
  nand2 gate1607(.a(s_151), .b(gate237inter3), .O(gate237inter10));
  nor2  gate1608(.a(gate237inter10), .b(gate237inter9), .O(gate237inter11));
  nor2  gate1609(.a(gate237inter11), .b(gate237inter6), .O(gate237inter12));
  nand2 gate1610(.a(gate237inter12), .b(gate237inter1), .O(G742));
nand2 gate238( .a(G257), .b(G709), .O(G745) );
nand2 gate239( .a(G260), .b(G712), .O(G748) );

  xor2  gate1709(.a(G715), .b(G263), .O(gate240inter0));
  nand2 gate1710(.a(gate240inter0), .b(s_166), .O(gate240inter1));
  and2  gate1711(.a(G715), .b(G263), .O(gate240inter2));
  inv1  gate1712(.a(s_166), .O(gate240inter3));
  inv1  gate1713(.a(s_167), .O(gate240inter4));
  nand2 gate1714(.a(gate240inter4), .b(gate240inter3), .O(gate240inter5));
  nor2  gate1715(.a(gate240inter5), .b(gate240inter2), .O(gate240inter6));
  inv1  gate1716(.a(G263), .O(gate240inter7));
  inv1  gate1717(.a(G715), .O(gate240inter8));
  nand2 gate1718(.a(gate240inter8), .b(gate240inter7), .O(gate240inter9));
  nand2 gate1719(.a(s_167), .b(gate240inter3), .O(gate240inter10));
  nor2  gate1720(.a(gate240inter10), .b(gate240inter9), .O(gate240inter11));
  nor2  gate1721(.a(gate240inter11), .b(gate240inter6), .O(gate240inter12));
  nand2 gate1722(.a(gate240inter12), .b(gate240inter1), .O(G751));
nand2 gate241( .a(G242), .b(G730), .O(G754) );
nand2 gate242( .a(G718), .b(G730), .O(G755) );
nand2 gate243( .a(G245), .b(G733), .O(G756) );

  xor2  gate1023(.a(G733), .b(G721), .O(gate244inter0));
  nand2 gate1024(.a(gate244inter0), .b(s_68), .O(gate244inter1));
  and2  gate1025(.a(G733), .b(G721), .O(gate244inter2));
  inv1  gate1026(.a(s_68), .O(gate244inter3));
  inv1  gate1027(.a(s_69), .O(gate244inter4));
  nand2 gate1028(.a(gate244inter4), .b(gate244inter3), .O(gate244inter5));
  nor2  gate1029(.a(gate244inter5), .b(gate244inter2), .O(gate244inter6));
  inv1  gate1030(.a(G721), .O(gate244inter7));
  inv1  gate1031(.a(G733), .O(gate244inter8));
  nand2 gate1032(.a(gate244inter8), .b(gate244inter7), .O(gate244inter9));
  nand2 gate1033(.a(s_69), .b(gate244inter3), .O(gate244inter10));
  nor2  gate1034(.a(gate244inter10), .b(gate244inter9), .O(gate244inter11));
  nor2  gate1035(.a(gate244inter11), .b(gate244inter6), .O(gate244inter12));
  nand2 gate1036(.a(gate244inter12), .b(gate244inter1), .O(G757));
nand2 gate245( .a(G248), .b(G736), .O(G758) );
nand2 gate246( .a(G724), .b(G736), .O(G759) );
nand2 gate247( .a(G251), .b(G739), .O(G760) );
nand2 gate248( .a(G727), .b(G739), .O(G761) );
nand2 gate249( .a(G254), .b(G742), .O(G762) );
nand2 gate250( .a(G706), .b(G742), .O(G763) );

  xor2  gate1387(.a(G745), .b(G257), .O(gate251inter0));
  nand2 gate1388(.a(gate251inter0), .b(s_120), .O(gate251inter1));
  and2  gate1389(.a(G745), .b(G257), .O(gate251inter2));
  inv1  gate1390(.a(s_120), .O(gate251inter3));
  inv1  gate1391(.a(s_121), .O(gate251inter4));
  nand2 gate1392(.a(gate251inter4), .b(gate251inter3), .O(gate251inter5));
  nor2  gate1393(.a(gate251inter5), .b(gate251inter2), .O(gate251inter6));
  inv1  gate1394(.a(G257), .O(gate251inter7));
  inv1  gate1395(.a(G745), .O(gate251inter8));
  nand2 gate1396(.a(gate251inter8), .b(gate251inter7), .O(gate251inter9));
  nand2 gate1397(.a(s_121), .b(gate251inter3), .O(gate251inter10));
  nor2  gate1398(.a(gate251inter10), .b(gate251inter9), .O(gate251inter11));
  nor2  gate1399(.a(gate251inter11), .b(gate251inter6), .O(gate251inter12));
  nand2 gate1400(.a(gate251inter12), .b(gate251inter1), .O(G764));

  xor2  gate1149(.a(G745), .b(G709), .O(gate252inter0));
  nand2 gate1150(.a(gate252inter0), .b(s_86), .O(gate252inter1));
  and2  gate1151(.a(G745), .b(G709), .O(gate252inter2));
  inv1  gate1152(.a(s_86), .O(gate252inter3));
  inv1  gate1153(.a(s_87), .O(gate252inter4));
  nand2 gate1154(.a(gate252inter4), .b(gate252inter3), .O(gate252inter5));
  nor2  gate1155(.a(gate252inter5), .b(gate252inter2), .O(gate252inter6));
  inv1  gate1156(.a(G709), .O(gate252inter7));
  inv1  gate1157(.a(G745), .O(gate252inter8));
  nand2 gate1158(.a(gate252inter8), .b(gate252inter7), .O(gate252inter9));
  nand2 gate1159(.a(s_87), .b(gate252inter3), .O(gate252inter10));
  nor2  gate1160(.a(gate252inter10), .b(gate252inter9), .O(gate252inter11));
  nor2  gate1161(.a(gate252inter11), .b(gate252inter6), .O(gate252inter12));
  nand2 gate1162(.a(gate252inter12), .b(gate252inter1), .O(G765));
nand2 gate253( .a(G260), .b(G748), .O(G766) );
nand2 gate254( .a(G712), .b(G748), .O(G767) );
nand2 gate255( .a(G263), .b(G751), .O(G768) );
nand2 gate256( .a(G715), .b(G751), .O(G769) );

  xor2  gate1723(.a(G755), .b(G754), .O(gate257inter0));
  nand2 gate1724(.a(gate257inter0), .b(s_168), .O(gate257inter1));
  and2  gate1725(.a(G755), .b(G754), .O(gate257inter2));
  inv1  gate1726(.a(s_168), .O(gate257inter3));
  inv1  gate1727(.a(s_169), .O(gate257inter4));
  nand2 gate1728(.a(gate257inter4), .b(gate257inter3), .O(gate257inter5));
  nor2  gate1729(.a(gate257inter5), .b(gate257inter2), .O(gate257inter6));
  inv1  gate1730(.a(G754), .O(gate257inter7));
  inv1  gate1731(.a(G755), .O(gate257inter8));
  nand2 gate1732(.a(gate257inter8), .b(gate257inter7), .O(gate257inter9));
  nand2 gate1733(.a(s_169), .b(gate257inter3), .O(gate257inter10));
  nor2  gate1734(.a(gate257inter10), .b(gate257inter9), .O(gate257inter11));
  nor2  gate1735(.a(gate257inter11), .b(gate257inter6), .O(gate257inter12));
  nand2 gate1736(.a(gate257inter12), .b(gate257inter1), .O(G770));

  xor2  gate701(.a(G757), .b(G756), .O(gate258inter0));
  nand2 gate702(.a(gate258inter0), .b(s_22), .O(gate258inter1));
  and2  gate703(.a(G757), .b(G756), .O(gate258inter2));
  inv1  gate704(.a(s_22), .O(gate258inter3));
  inv1  gate705(.a(s_23), .O(gate258inter4));
  nand2 gate706(.a(gate258inter4), .b(gate258inter3), .O(gate258inter5));
  nor2  gate707(.a(gate258inter5), .b(gate258inter2), .O(gate258inter6));
  inv1  gate708(.a(G756), .O(gate258inter7));
  inv1  gate709(.a(G757), .O(gate258inter8));
  nand2 gate710(.a(gate258inter8), .b(gate258inter7), .O(gate258inter9));
  nand2 gate711(.a(s_23), .b(gate258inter3), .O(gate258inter10));
  nor2  gate712(.a(gate258inter10), .b(gate258inter9), .O(gate258inter11));
  nor2  gate713(.a(gate258inter11), .b(gate258inter6), .O(gate258inter12));
  nand2 gate714(.a(gate258inter12), .b(gate258inter1), .O(G773));

  xor2  gate1331(.a(G759), .b(G758), .O(gate259inter0));
  nand2 gate1332(.a(gate259inter0), .b(s_112), .O(gate259inter1));
  and2  gate1333(.a(G759), .b(G758), .O(gate259inter2));
  inv1  gate1334(.a(s_112), .O(gate259inter3));
  inv1  gate1335(.a(s_113), .O(gate259inter4));
  nand2 gate1336(.a(gate259inter4), .b(gate259inter3), .O(gate259inter5));
  nor2  gate1337(.a(gate259inter5), .b(gate259inter2), .O(gate259inter6));
  inv1  gate1338(.a(G758), .O(gate259inter7));
  inv1  gate1339(.a(G759), .O(gate259inter8));
  nand2 gate1340(.a(gate259inter8), .b(gate259inter7), .O(gate259inter9));
  nand2 gate1341(.a(s_113), .b(gate259inter3), .O(gate259inter10));
  nor2  gate1342(.a(gate259inter10), .b(gate259inter9), .O(gate259inter11));
  nor2  gate1343(.a(gate259inter11), .b(gate259inter6), .O(gate259inter12));
  nand2 gate1344(.a(gate259inter12), .b(gate259inter1), .O(G776));
nand2 gate260( .a(G760), .b(G761), .O(G779) );
nand2 gate261( .a(G762), .b(G763), .O(G782) );
nand2 gate262( .a(G764), .b(G765), .O(G785) );
nand2 gate263( .a(G766), .b(G767), .O(G788) );
nand2 gate264( .a(G768), .b(G769), .O(G791) );
nand2 gate265( .a(G642), .b(G770), .O(G794) );
nand2 gate266( .a(G645), .b(G773), .O(G797) );
nand2 gate267( .a(G648), .b(G776), .O(G800) );

  xor2  gate1485(.a(G779), .b(G651), .O(gate268inter0));
  nand2 gate1486(.a(gate268inter0), .b(s_134), .O(gate268inter1));
  and2  gate1487(.a(G779), .b(G651), .O(gate268inter2));
  inv1  gate1488(.a(s_134), .O(gate268inter3));
  inv1  gate1489(.a(s_135), .O(gate268inter4));
  nand2 gate1490(.a(gate268inter4), .b(gate268inter3), .O(gate268inter5));
  nor2  gate1491(.a(gate268inter5), .b(gate268inter2), .O(gate268inter6));
  inv1  gate1492(.a(G651), .O(gate268inter7));
  inv1  gate1493(.a(G779), .O(gate268inter8));
  nand2 gate1494(.a(gate268inter8), .b(gate268inter7), .O(gate268inter9));
  nand2 gate1495(.a(s_135), .b(gate268inter3), .O(gate268inter10));
  nor2  gate1496(.a(gate268inter10), .b(gate268inter9), .O(gate268inter11));
  nor2  gate1497(.a(gate268inter11), .b(gate268inter6), .O(gate268inter12));
  nand2 gate1498(.a(gate268inter12), .b(gate268inter1), .O(G803));
nand2 gate269( .a(G654), .b(G782), .O(G806) );
nand2 gate270( .a(G657), .b(G785), .O(G809) );
nand2 gate271( .a(G660), .b(G788), .O(G812) );
nand2 gate272( .a(G663), .b(G791), .O(G815) );
nand2 gate273( .a(G642), .b(G794), .O(G818) );
nand2 gate274( .a(G770), .b(G794), .O(G819) );
nand2 gate275( .a(G645), .b(G797), .O(G820) );
nand2 gate276( .a(G773), .b(G797), .O(G821) );
nand2 gate277( .a(G648), .b(G800), .O(G822) );
nand2 gate278( .a(G776), .b(G800), .O(G823) );
nand2 gate279( .a(G651), .b(G803), .O(G824) );

  xor2  gate1093(.a(G803), .b(G779), .O(gate280inter0));
  nand2 gate1094(.a(gate280inter0), .b(s_78), .O(gate280inter1));
  and2  gate1095(.a(G803), .b(G779), .O(gate280inter2));
  inv1  gate1096(.a(s_78), .O(gate280inter3));
  inv1  gate1097(.a(s_79), .O(gate280inter4));
  nand2 gate1098(.a(gate280inter4), .b(gate280inter3), .O(gate280inter5));
  nor2  gate1099(.a(gate280inter5), .b(gate280inter2), .O(gate280inter6));
  inv1  gate1100(.a(G779), .O(gate280inter7));
  inv1  gate1101(.a(G803), .O(gate280inter8));
  nand2 gate1102(.a(gate280inter8), .b(gate280inter7), .O(gate280inter9));
  nand2 gate1103(.a(s_79), .b(gate280inter3), .O(gate280inter10));
  nor2  gate1104(.a(gate280inter10), .b(gate280inter9), .O(gate280inter11));
  nor2  gate1105(.a(gate280inter11), .b(gate280inter6), .O(gate280inter12));
  nand2 gate1106(.a(gate280inter12), .b(gate280inter1), .O(G825));
nand2 gate281( .a(G654), .b(G806), .O(G826) );
nand2 gate282( .a(G782), .b(G806), .O(G827) );

  xor2  gate1275(.a(G809), .b(G657), .O(gate283inter0));
  nand2 gate1276(.a(gate283inter0), .b(s_104), .O(gate283inter1));
  and2  gate1277(.a(G809), .b(G657), .O(gate283inter2));
  inv1  gate1278(.a(s_104), .O(gate283inter3));
  inv1  gate1279(.a(s_105), .O(gate283inter4));
  nand2 gate1280(.a(gate283inter4), .b(gate283inter3), .O(gate283inter5));
  nor2  gate1281(.a(gate283inter5), .b(gate283inter2), .O(gate283inter6));
  inv1  gate1282(.a(G657), .O(gate283inter7));
  inv1  gate1283(.a(G809), .O(gate283inter8));
  nand2 gate1284(.a(gate283inter8), .b(gate283inter7), .O(gate283inter9));
  nand2 gate1285(.a(s_105), .b(gate283inter3), .O(gate283inter10));
  nor2  gate1286(.a(gate283inter10), .b(gate283inter9), .O(gate283inter11));
  nor2  gate1287(.a(gate283inter11), .b(gate283inter6), .O(gate283inter12));
  nand2 gate1288(.a(gate283inter12), .b(gate283inter1), .O(G828));
nand2 gate284( .a(G785), .b(G809), .O(G829) );
nand2 gate285( .a(G660), .b(G812), .O(G830) );
nand2 gate286( .a(G788), .b(G812), .O(G831) );

  xor2  gate1429(.a(G815), .b(G663), .O(gate287inter0));
  nand2 gate1430(.a(gate287inter0), .b(s_126), .O(gate287inter1));
  and2  gate1431(.a(G815), .b(G663), .O(gate287inter2));
  inv1  gate1432(.a(s_126), .O(gate287inter3));
  inv1  gate1433(.a(s_127), .O(gate287inter4));
  nand2 gate1434(.a(gate287inter4), .b(gate287inter3), .O(gate287inter5));
  nor2  gate1435(.a(gate287inter5), .b(gate287inter2), .O(gate287inter6));
  inv1  gate1436(.a(G663), .O(gate287inter7));
  inv1  gate1437(.a(G815), .O(gate287inter8));
  nand2 gate1438(.a(gate287inter8), .b(gate287inter7), .O(gate287inter9));
  nand2 gate1439(.a(s_127), .b(gate287inter3), .O(gate287inter10));
  nor2  gate1440(.a(gate287inter10), .b(gate287inter9), .O(gate287inter11));
  nor2  gate1441(.a(gate287inter11), .b(gate287inter6), .O(gate287inter12));
  nand2 gate1442(.a(gate287inter12), .b(gate287inter1), .O(G832));
nand2 gate288( .a(G791), .b(G815), .O(G833) );
nand2 gate289( .a(G818), .b(G819), .O(G834) );
nand2 gate290( .a(G820), .b(G821), .O(G847) );
nand2 gate291( .a(G822), .b(G823), .O(G860) );
nand2 gate292( .a(G824), .b(G825), .O(G873) );
nand2 gate293( .a(G828), .b(G829), .O(G886) );
nand2 gate294( .a(G832), .b(G833), .O(G899) );
nand2 gate295( .a(G830), .b(G831), .O(G912) );
nand2 gate296( .a(G826), .b(G827), .O(G925) );
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );

  xor2  gate855(.a(G1036), .b(G1), .O(gate387inter0));
  nand2 gate856(.a(gate387inter0), .b(s_44), .O(gate387inter1));
  and2  gate857(.a(G1036), .b(G1), .O(gate387inter2));
  inv1  gate858(.a(s_44), .O(gate387inter3));
  inv1  gate859(.a(s_45), .O(gate387inter4));
  nand2 gate860(.a(gate387inter4), .b(gate387inter3), .O(gate387inter5));
  nor2  gate861(.a(gate387inter5), .b(gate387inter2), .O(gate387inter6));
  inv1  gate862(.a(G1), .O(gate387inter7));
  inv1  gate863(.a(G1036), .O(gate387inter8));
  nand2 gate864(.a(gate387inter8), .b(gate387inter7), .O(gate387inter9));
  nand2 gate865(.a(s_45), .b(gate387inter3), .O(gate387inter10));
  nor2  gate866(.a(gate387inter10), .b(gate387inter9), .O(gate387inter11));
  nor2  gate867(.a(gate387inter11), .b(gate387inter6), .O(gate387inter12));
  nand2 gate868(.a(gate387inter12), .b(gate387inter1), .O(G1132));

  xor2  gate1625(.a(G1039), .b(G2), .O(gate388inter0));
  nand2 gate1626(.a(gate388inter0), .b(s_154), .O(gate388inter1));
  and2  gate1627(.a(G1039), .b(G2), .O(gate388inter2));
  inv1  gate1628(.a(s_154), .O(gate388inter3));
  inv1  gate1629(.a(s_155), .O(gate388inter4));
  nand2 gate1630(.a(gate388inter4), .b(gate388inter3), .O(gate388inter5));
  nor2  gate1631(.a(gate388inter5), .b(gate388inter2), .O(gate388inter6));
  inv1  gate1632(.a(G2), .O(gate388inter7));
  inv1  gate1633(.a(G1039), .O(gate388inter8));
  nand2 gate1634(.a(gate388inter8), .b(gate388inter7), .O(gate388inter9));
  nand2 gate1635(.a(s_155), .b(gate388inter3), .O(gate388inter10));
  nor2  gate1636(.a(gate388inter10), .b(gate388inter9), .O(gate388inter11));
  nor2  gate1637(.a(gate388inter11), .b(gate388inter6), .O(gate388inter12));
  nand2 gate1638(.a(gate388inter12), .b(gate388inter1), .O(G1135));
nand2 gate389( .a(G3), .b(G1042), .O(G1138) );
nand2 gate390( .a(G4), .b(G1045), .O(G1141) );
nand2 gate391( .a(G5), .b(G1048), .O(G1144) );

  xor2  gate883(.a(G1051), .b(G6), .O(gate392inter0));
  nand2 gate884(.a(gate392inter0), .b(s_48), .O(gate392inter1));
  and2  gate885(.a(G1051), .b(G6), .O(gate392inter2));
  inv1  gate886(.a(s_48), .O(gate392inter3));
  inv1  gate887(.a(s_49), .O(gate392inter4));
  nand2 gate888(.a(gate392inter4), .b(gate392inter3), .O(gate392inter5));
  nor2  gate889(.a(gate392inter5), .b(gate392inter2), .O(gate392inter6));
  inv1  gate890(.a(G6), .O(gate392inter7));
  inv1  gate891(.a(G1051), .O(gate392inter8));
  nand2 gate892(.a(gate392inter8), .b(gate392inter7), .O(gate392inter9));
  nand2 gate893(.a(s_49), .b(gate392inter3), .O(gate392inter10));
  nor2  gate894(.a(gate392inter10), .b(gate392inter9), .O(gate392inter11));
  nor2  gate895(.a(gate392inter11), .b(gate392inter6), .O(gate392inter12));
  nand2 gate896(.a(gate392inter12), .b(gate392inter1), .O(G1147));
nand2 gate393( .a(G7), .b(G1054), .O(G1150) );

  xor2  gate1177(.a(G1057), .b(G8), .O(gate394inter0));
  nand2 gate1178(.a(gate394inter0), .b(s_90), .O(gate394inter1));
  and2  gate1179(.a(G1057), .b(G8), .O(gate394inter2));
  inv1  gate1180(.a(s_90), .O(gate394inter3));
  inv1  gate1181(.a(s_91), .O(gate394inter4));
  nand2 gate1182(.a(gate394inter4), .b(gate394inter3), .O(gate394inter5));
  nor2  gate1183(.a(gate394inter5), .b(gate394inter2), .O(gate394inter6));
  inv1  gate1184(.a(G8), .O(gate394inter7));
  inv1  gate1185(.a(G1057), .O(gate394inter8));
  nand2 gate1186(.a(gate394inter8), .b(gate394inter7), .O(gate394inter9));
  nand2 gate1187(.a(s_91), .b(gate394inter3), .O(gate394inter10));
  nor2  gate1188(.a(gate394inter10), .b(gate394inter9), .O(gate394inter11));
  nor2  gate1189(.a(gate394inter11), .b(gate394inter6), .O(gate394inter12));
  nand2 gate1190(.a(gate394inter12), .b(gate394inter1), .O(G1153));

  xor2  gate645(.a(G1060), .b(G9), .O(gate395inter0));
  nand2 gate646(.a(gate395inter0), .b(s_14), .O(gate395inter1));
  and2  gate647(.a(G1060), .b(G9), .O(gate395inter2));
  inv1  gate648(.a(s_14), .O(gate395inter3));
  inv1  gate649(.a(s_15), .O(gate395inter4));
  nand2 gate650(.a(gate395inter4), .b(gate395inter3), .O(gate395inter5));
  nor2  gate651(.a(gate395inter5), .b(gate395inter2), .O(gate395inter6));
  inv1  gate652(.a(G9), .O(gate395inter7));
  inv1  gate653(.a(G1060), .O(gate395inter8));
  nand2 gate654(.a(gate395inter8), .b(gate395inter7), .O(gate395inter9));
  nand2 gate655(.a(s_15), .b(gate395inter3), .O(gate395inter10));
  nor2  gate656(.a(gate395inter10), .b(gate395inter9), .O(gate395inter11));
  nor2  gate657(.a(gate395inter11), .b(gate395inter6), .O(gate395inter12));
  nand2 gate658(.a(gate395inter12), .b(gate395inter1), .O(G1156));
nand2 gate396( .a(G10), .b(G1063), .O(G1159) );
nand2 gate397( .a(G11), .b(G1066), .O(G1162) );
nand2 gate398( .a(G12), .b(G1069), .O(G1165) );
nand2 gate399( .a(G13), .b(G1072), .O(G1168) );
nand2 gate400( .a(G14), .b(G1075), .O(G1171) );

  xor2  gate547(.a(G1078), .b(G15), .O(gate401inter0));
  nand2 gate548(.a(gate401inter0), .b(s_0), .O(gate401inter1));
  and2  gate549(.a(G1078), .b(G15), .O(gate401inter2));
  inv1  gate550(.a(s_0), .O(gate401inter3));
  inv1  gate551(.a(s_1), .O(gate401inter4));
  nand2 gate552(.a(gate401inter4), .b(gate401inter3), .O(gate401inter5));
  nor2  gate553(.a(gate401inter5), .b(gate401inter2), .O(gate401inter6));
  inv1  gate554(.a(G15), .O(gate401inter7));
  inv1  gate555(.a(G1078), .O(gate401inter8));
  nand2 gate556(.a(gate401inter8), .b(gate401inter7), .O(gate401inter9));
  nand2 gate557(.a(s_1), .b(gate401inter3), .O(gate401inter10));
  nor2  gate558(.a(gate401inter10), .b(gate401inter9), .O(gate401inter11));
  nor2  gate559(.a(gate401inter11), .b(gate401inter6), .O(gate401inter12));
  nand2 gate560(.a(gate401inter12), .b(gate401inter1), .O(G1174));
nand2 gate402( .a(G16), .b(G1081), .O(G1177) );
nand2 gate403( .a(G17), .b(G1084), .O(G1180) );
nand2 gate404( .a(G18), .b(G1087), .O(G1183) );
nand2 gate405( .a(G19), .b(G1090), .O(G1186) );
nand2 gate406( .a(G20), .b(G1093), .O(G1189) );
nand2 gate407( .a(G21), .b(G1096), .O(G1192) );
nand2 gate408( .a(G22), .b(G1099), .O(G1195) );
nand2 gate409( .a(G23), .b(G1102), .O(G1198) );
nand2 gate410( .a(G24), .b(G1105), .O(G1201) );

  xor2  gate1541(.a(G1108), .b(G25), .O(gate411inter0));
  nand2 gate1542(.a(gate411inter0), .b(s_142), .O(gate411inter1));
  and2  gate1543(.a(G1108), .b(G25), .O(gate411inter2));
  inv1  gate1544(.a(s_142), .O(gate411inter3));
  inv1  gate1545(.a(s_143), .O(gate411inter4));
  nand2 gate1546(.a(gate411inter4), .b(gate411inter3), .O(gate411inter5));
  nor2  gate1547(.a(gate411inter5), .b(gate411inter2), .O(gate411inter6));
  inv1  gate1548(.a(G25), .O(gate411inter7));
  inv1  gate1549(.a(G1108), .O(gate411inter8));
  nand2 gate1550(.a(gate411inter8), .b(gate411inter7), .O(gate411inter9));
  nand2 gate1551(.a(s_143), .b(gate411inter3), .O(gate411inter10));
  nor2  gate1552(.a(gate411inter10), .b(gate411inter9), .O(gate411inter11));
  nor2  gate1553(.a(gate411inter11), .b(gate411inter6), .O(gate411inter12));
  nand2 gate1554(.a(gate411inter12), .b(gate411inter1), .O(G1204));
nand2 gate412( .a(G26), .b(G1111), .O(G1207) );

  xor2  gate673(.a(G1114), .b(G27), .O(gate413inter0));
  nand2 gate674(.a(gate413inter0), .b(s_18), .O(gate413inter1));
  and2  gate675(.a(G1114), .b(G27), .O(gate413inter2));
  inv1  gate676(.a(s_18), .O(gate413inter3));
  inv1  gate677(.a(s_19), .O(gate413inter4));
  nand2 gate678(.a(gate413inter4), .b(gate413inter3), .O(gate413inter5));
  nor2  gate679(.a(gate413inter5), .b(gate413inter2), .O(gate413inter6));
  inv1  gate680(.a(G27), .O(gate413inter7));
  inv1  gate681(.a(G1114), .O(gate413inter8));
  nand2 gate682(.a(gate413inter8), .b(gate413inter7), .O(gate413inter9));
  nand2 gate683(.a(s_19), .b(gate413inter3), .O(gate413inter10));
  nor2  gate684(.a(gate413inter10), .b(gate413inter9), .O(gate413inter11));
  nor2  gate685(.a(gate413inter11), .b(gate413inter6), .O(gate413inter12));
  nand2 gate686(.a(gate413inter12), .b(gate413inter1), .O(G1210));
nand2 gate414( .a(G28), .b(G1117), .O(G1213) );
nand2 gate415( .a(G29), .b(G1120), .O(G1216) );
nand2 gate416( .a(G30), .b(G1123), .O(G1219) );
nand2 gate417( .a(G31), .b(G1126), .O(G1222) );
nand2 gate418( .a(G32), .b(G1129), .O(G1225) );
nand2 gate419( .a(G1), .b(G1132), .O(G1228) );
nand2 gate420( .a(G1036), .b(G1132), .O(G1229) );

  xor2  gate729(.a(G1135), .b(G2), .O(gate421inter0));
  nand2 gate730(.a(gate421inter0), .b(s_26), .O(gate421inter1));
  and2  gate731(.a(G1135), .b(G2), .O(gate421inter2));
  inv1  gate732(.a(s_26), .O(gate421inter3));
  inv1  gate733(.a(s_27), .O(gate421inter4));
  nand2 gate734(.a(gate421inter4), .b(gate421inter3), .O(gate421inter5));
  nor2  gate735(.a(gate421inter5), .b(gate421inter2), .O(gate421inter6));
  inv1  gate736(.a(G2), .O(gate421inter7));
  inv1  gate737(.a(G1135), .O(gate421inter8));
  nand2 gate738(.a(gate421inter8), .b(gate421inter7), .O(gate421inter9));
  nand2 gate739(.a(s_27), .b(gate421inter3), .O(gate421inter10));
  nor2  gate740(.a(gate421inter10), .b(gate421inter9), .O(gate421inter11));
  nor2  gate741(.a(gate421inter11), .b(gate421inter6), .O(gate421inter12));
  nand2 gate742(.a(gate421inter12), .b(gate421inter1), .O(G1230));
nand2 gate422( .a(G1039), .b(G1135), .O(G1231) );
nand2 gate423( .a(G3), .b(G1138), .O(G1232) );
nand2 gate424( .a(G1042), .b(G1138), .O(G1233) );
nand2 gate425( .a(G4), .b(G1141), .O(G1234) );
nand2 gate426( .a(G1045), .b(G1141), .O(G1235) );
nand2 gate427( .a(G5), .b(G1144), .O(G1236) );
nand2 gate428( .a(G1048), .b(G1144), .O(G1237) );
nand2 gate429( .a(G6), .b(G1147), .O(G1238) );
nand2 gate430( .a(G1051), .b(G1147), .O(G1239) );
nand2 gate431( .a(G7), .b(G1150), .O(G1240) );
nand2 gate432( .a(G1054), .b(G1150), .O(G1241) );
nand2 gate433( .a(G8), .b(G1153), .O(G1242) );
nand2 gate434( .a(G1057), .b(G1153), .O(G1243) );

  xor2  gate1513(.a(G1156), .b(G9), .O(gate435inter0));
  nand2 gate1514(.a(gate435inter0), .b(s_138), .O(gate435inter1));
  and2  gate1515(.a(G1156), .b(G9), .O(gate435inter2));
  inv1  gate1516(.a(s_138), .O(gate435inter3));
  inv1  gate1517(.a(s_139), .O(gate435inter4));
  nand2 gate1518(.a(gate435inter4), .b(gate435inter3), .O(gate435inter5));
  nor2  gate1519(.a(gate435inter5), .b(gate435inter2), .O(gate435inter6));
  inv1  gate1520(.a(G9), .O(gate435inter7));
  inv1  gate1521(.a(G1156), .O(gate435inter8));
  nand2 gate1522(.a(gate435inter8), .b(gate435inter7), .O(gate435inter9));
  nand2 gate1523(.a(s_139), .b(gate435inter3), .O(gate435inter10));
  nor2  gate1524(.a(gate435inter10), .b(gate435inter9), .O(gate435inter11));
  nor2  gate1525(.a(gate435inter11), .b(gate435inter6), .O(gate435inter12));
  nand2 gate1526(.a(gate435inter12), .b(gate435inter1), .O(G1244));
nand2 gate436( .a(G1060), .b(G1156), .O(G1245) );

  xor2  gate1457(.a(G1159), .b(G10), .O(gate437inter0));
  nand2 gate1458(.a(gate437inter0), .b(s_130), .O(gate437inter1));
  and2  gate1459(.a(G1159), .b(G10), .O(gate437inter2));
  inv1  gate1460(.a(s_130), .O(gate437inter3));
  inv1  gate1461(.a(s_131), .O(gate437inter4));
  nand2 gate1462(.a(gate437inter4), .b(gate437inter3), .O(gate437inter5));
  nor2  gate1463(.a(gate437inter5), .b(gate437inter2), .O(gate437inter6));
  inv1  gate1464(.a(G10), .O(gate437inter7));
  inv1  gate1465(.a(G1159), .O(gate437inter8));
  nand2 gate1466(.a(gate437inter8), .b(gate437inter7), .O(gate437inter9));
  nand2 gate1467(.a(s_131), .b(gate437inter3), .O(gate437inter10));
  nor2  gate1468(.a(gate437inter10), .b(gate437inter9), .O(gate437inter11));
  nor2  gate1469(.a(gate437inter11), .b(gate437inter6), .O(gate437inter12));
  nand2 gate1470(.a(gate437inter12), .b(gate437inter1), .O(G1246));
nand2 gate438( .a(G1063), .b(G1159), .O(G1247) );
nand2 gate439( .a(G11), .b(G1162), .O(G1248) );
nand2 gate440( .a(G1066), .b(G1162), .O(G1249) );

  xor2  gate827(.a(G1165), .b(G12), .O(gate441inter0));
  nand2 gate828(.a(gate441inter0), .b(s_40), .O(gate441inter1));
  and2  gate829(.a(G1165), .b(G12), .O(gate441inter2));
  inv1  gate830(.a(s_40), .O(gate441inter3));
  inv1  gate831(.a(s_41), .O(gate441inter4));
  nand2 gate832(.a(gate441inter4), .b(gate441inter3), .O(gate441inter5));
  nor2  gate833(.a(gate441inter5), .b(gate441inter2), .O(gate441inter6));
  inv1  gate834(.a(G12), .O(gate441inter7));
  inv1  gate835(.a(G1165), .O(gate441inter8));
  nand2 gate836(.a(gate441inter8), .b(gate441inter7), .O(gate441inter9));
  nand2 gate837(.a(s_41), .b(gate441inter3), .O(gate441inter10));
  nor2  gate838(.a(gate441inter10), .b(gate441inter9), .O(gate441inter11));
  nor2  gate839(.a(gate441inter11), .b(gate441inter6), .O(gate441inter12));
  nand2 gate840(.a(gate441inter12), .b(gate441inter1), .O(G1250));
nand2 gate442( .a(G1069), .b(G1165), .O(G1251) );

  xor2  gate1695(.a(G1168), .b(G13), .O(gate443inter0));
  nand2 gate1696(.a(gate443inter0), .b(s_164), .O(gate443inter1));
  and2  gate1697(.a(G1168), .b(G13), .O(gate443inter2));
  inv1  gate1698(.a(s_164), .O(gate443inter3));
  inv1  gate1699(.a(s_165), .O(gate443inter4));
  nand2 gate1700(.a(gate443inter4), .b(gate443inter3), .O(gate443inter5));
  nor2  gate1701(.a(gate443inter5), .b(gate443inter2), .O(gate443inter6));
  inv1  gate1702(.a(G13), .O(gate443inter7));
  inv1  gate1703(.a(G1168), .O(gate443inter8));
  nand2 gate1704(.a(gate443inter8), .b(gate443inter7), .O(gate443inter9));
  nand2 gate1705(.a(s_165), .b(gate443inter3), .O(gate443inter10));
  nor2  gate1706(.a(gate443inter10), .b(gate443inter9), .O(gate443inter11));
  nor2  gate1707(.a(gate443inter11), .b(gate443inter6), .O(gate443inter12));
  nand2 gate1708(.a(gate443inter12), .b(gate443inter1), .O(G1252));
nand2 gate444( .a(G1072), .b(G1168), .O(G1253) );
nand2 gate445( .a(G14), .b(G1171), .O(G1254) );
nand2 gate446( .a(G1075), .b(G1171), .O(G1255) );
nand2 gate447( .a(G15), .b(G1174), .O(G1256) );
nand2 gate448( .a(G1078), .b(G1174), .O(G1257) );
nand2 gate449( .a(G16), .b(G1177), .O(G1258) );
nand2 gate450( .a(G1081), .b(G1177), .O(G1259) );
nand2 gate451( .a(G17), .b(G1180), .O(G1260) );
nand2 gate452( .a(G1084), .b(G1180), .O(G1261) );
nand2 gate453( .a(G18), .b(G1183), .O(G1262) );
nand2 gate454( .a(G1087), .b(G1183), .O(G1263) );
nand2 gate455( .a(G19), .b(G1186), .O(G1264) );
nand2 gate456( .a(G1090), .b(G1186), .O(G1265) );
nand2 gate457( .a(G20), .b(G1189), .O(G1266) );
nand2 gate458( .a(G1093), .b(G1189), .O(G1267) );
nand2 gate459( .a(G21), .b(G1192), .O(G1268) );
nand2 gate460( .a(G1096), .b(G1192), .O(G1269) );
nand2 gate461( .a(G22), .b(G1195), .O(G1270) );

  xor2  gate953(.a(G1195), .b(G1099), .O(gate462inter0));
  nand2 gate954(.a(gate462inter0), .b(s_58), .O(gate462inter1));
  and2  gate955(.a(G1195), .b(G1099), .O(gate462inter2));
  inv1  gate956(.a(s_58), .O(gate462inter3));
  inv1  gate957(.a(s_59), .O(gate462inter4));
  nand2 gate958(.a(gate462inter4), .b(gate462inter3), .O(gate462inter5));
  nor2  gate959(.a(gate462inter5), .b(gate462inter2), .O(gate462inter6));
  inv1  gate960(.a(G1099), .O(gate462inter7));
  inv1  gate961(.a(G1195), .O(gate462inter8));
  nand2 gate962(.a(gate462inter8), .b(gate462inter7), .O(gate462inter9));
  nand2 gate963(.a(s_59), .b(gate462inter3), .O(gate462inter10));
  nor2  gate964(.a(gate462inter10), .b(gate462inter9), .O(gate462inter11));
  nor2  gate965(.a(gate462inter11), .b(gate462inter6), .O(gate462inter12));
  nand2 gate966(.a(gate462inter12), .b(gate462inter1), .O(G1271));
nand2 gate463( .a(G23), .b(G1198), .O(G1272) );
nand2 gate464( .a(G1102), .b(G1198), .O(G1273) );

  xor2  gate659(.a(G1201), .b(G24), .O(gate465inter0));
  nand2 gate660(.a(gate465inter0), .b(s_16), .O(gate465inter1));
  and2  gate661(.a(G1201), .b(G24), .O(gate465inter2));
  inv1  gate662(.a(s_16), .O(gate465inter3));
  inv1  gate663(.a(s_17), .O(gate465inter4));
  nand2 gate664(.a(gate465inter4), .b(gate465inter3), .O(gate465inter5));
  nor2  gate665(.a(gate465inter5), .b(gate465inter2), .O(gate465inter6));
  inv1  gate666(.a(G24), .O(gate465inter7));
  inv1  gate667(.a(G1201), .O(gate465inter8));
  nand2 gate668(.a(gate465inter8), .b(gate465inter7), .O(gate465inter9));
  nand2 gate669(.a(s_17), .b(gate465inter3), .O(gate465inter10));
  nor2  gate670(.a(gate465inter10), .b(gate465inter9), .O(gate465inter11));
  nor2  gate671(.a(gate465inter11), .b(gate465inter6), .O(gate465inter12));
  nand2 gate672(.a(gate465inter12), .b(gate465inter1), .O(G1274));
nand2 gate466( .a(G1105), .b(G1201), .O(G1275) );
nand2 gate467( .a(G25), .b(G1204), .O(G1276) );
nand2 gate468( .a(G1108), .b(G1204), .O(G1277) );
nand2 gate469( .a(G26), .b(G1207), .O(G1278) );

  xor2  gate967(.a(G1207), .b(G1111), .O(gate470inter0));
  nand2 gate968(.a(gate470inter0), .b(s_60), .O(gate470inter1));
  and2  gate969(.a(G1207), .b(G1111), .O(gate470inter2));
  inv1  gate970(.a(s_60), .O(gate470inter3));
  inv1  gate971(.a(s_61), .O(gate470inter4));
  nand2 gate972(.a(gate470inter4), .b(gate470inter3), .O(gate470inter5));
  nor2  gate973(.a(gate470inter5), .b(gate470inter2), .O(gate470inter6));
  inv1  gate974(.a(G1111), .O(gate470inter7));
  inv1  gate975(.a(G1207), .O(gate470inter8));
  nand2 gate976(.a(gate470inter8), .b(gate470inter7), .O(gate470inter9));
  nand2 gate977(.a(s_61), .b(gate470inter3), .O(gate470inter10));
  nor2  gate978(.a(gate470inter10), .b(gate470inter9), .O(gate470inter11));
  nor2  gate979(.a(gate470inter11), .b(gate470inter6), .O(gate470inter12));
  nand2 gate980(.a(gate470inter12), .b(gate470inter1), .O(G1279));
nand2 gate471( .a(G27), .b(G1210), .O(G1280) );
nand2 gate472( .a(G1114), .b(G1210), .O(G1281) );
nand2 gate473( .a(G28), .b(G1213), .O(G1282) );

  xor2  gate1779(.a(G1213), .b(G1117), .O(gate474inter0));
  nand2 gate1780(.a(gate474inter0), .b(s_176), .O(gate474inter1));
  and2  gate1781(.a(G1213), .b(G1117), .O(gate474inter2));
  inv1  gate1782(.a(s_176), .O(gate474inter3));
  inv1  gate1783(.a(s_177), .O(gate474inter4));
  nand2 gate1784(.a(gate474inter4), .b(gate474inter3), .O(gate474inter5));
  nor2  gate1785(.a(gate474inter5), .b(gate474inter2), .O(gate474inter6));
  inv1  gate1786(.a(G1117), .O(gate474inter7));
  inv1  gate1787(.a(G1213), .O(gate474inter8));
  nand2 gate1788(.a(gate474inter8), .b(gate474inter7), .O(gate474inter9));
  nand2 gate1789(.a(s_177), .b(gate474inter3), .O(gate474inter10));
  nor2  gate1790(.a(gate474inter10), .b(gate474inter9), .O(gate474inter11));
  nor2  gate1791(.a(gate474inter11), .b(gate474inter6), .O(gate474inter12));
  nand2 gate1792(.a(gate474inter12), .b(gate474inter1), .O(G1283));

  xor2  gate1737(.a(G1216), .b(G29), .O(gate475inter0));
  nand2 gate1738(.a(gate475inter0), .b(s_170), .O(gate475inter1));
  and2  gate1739(.a(G1216), .b(G29), .O(gate475inter2));
  inv1  gate1740(.a(s_170), .O(gate475inter3));
  inv1  gate1741(.a(s_171), .O(gate475inter4));
  nand2 gate1742(.a(gate475inter4), .b(gate475inter3), .O(gate475inter5));
  nor2  gate1743(.a(gate475inter5), .b(gate475inter2), .O(gate475inter6));
  inv1  gate1744(.a(G29), .O(gate475inter7));
  inv1  gate1745(.a(G1216), .O(gate475inter8));
  nand2 gate1746(.a(gate475inter8), .b(gate475inter7), .O(gate475inter9));
  nand2 gate1747(.a(s_171), .b(gate475inter3), .O(gate475inter10));
  nor2  gate1748(.a(gate475inter10), .b(gate475inter9), .O(gate475inter11));
  nor2  gate1749(.a(gate475inter11), .b(gate475inter6), .O(gate475inter12));
  nand2 gate1750(.a(gate475inter12), .b(gate475inter1), .O(G1284));
nand2 gate476( .a(G1120), .b(G1216), .O(G1285) );
nand2 gate477( .a(G30), .b(G1219), .O(G1286) );
nand2 gate478( .a(G1123), .b(G1219), .O(G1287) );
nand2 gate479( .a(G31), .b(G1222), .O(G1288) );

  xor2  gate1681(.a(G1222), .b(G1126), .O(gate480inter0));
  nand2 gate1682(.a(gate480inter0), .b(s_162), .O(gate480inter1));
  and2  gate1683(.a(G1222), .b(G1126), .O(gate480inter2));
  inv1  gate1684(.a(s_162), .O(gate480inter3));
  inv1  gate1685(.a(s_163), .O(gate480inter4));
  nand2 gate1686(.a(gate480inter4), .b(gate480inter3), .O(gate480inter5));
  nor2  gate1687(.a(gate480inter5), .b(gate480inter2), .O(gate480inter6));
  inv1  gate1688(.a(G1126), .O(gate480inter7));
  inv1  gate1689(.a(G1222), .O(gate480inter8));
  nand2 gate1690(.a(gate480inter8), .b(gate480inter7), .O(gate480inter9));
  nand2 gate1691(.a(s_163), .b(gate480inter3), .O(gate480inter10));
  nor2  gate1692(.a(gate480inter10), .b(gate480inter9), .O(gate480inter11));
  nor2  gate1693(.a(gate480inter11), .b(gate480inter6), .O(gate480inter12));
  nand2 gate1694(.a(gate480inter12), .b(gate480inter1), .O(G1289));

  xor2  gate757(.a(G1225), .b(G32), .O(gate481inter0));
  nand2 gate758(.a(gate481inter0), .b(s_30), .O(gate481inter1));
  and2  gate759(.a(G1225), .b(G32), .O(gate481inter2));
  inv1  gate760(.a(s_30), .O(gate481inter3));
  inv1  gate761(.a(s_31), .O(gate481inter4));
  nand2 gate762(.a(gate481inter4), .b(gate481inter3), .O(gate481inter5));
  nor2  gate763(.a(gate481inter5), .b(gate481inter2), .O(gate481inter6));
  inv1  gate764(.a(G32), .O(gate481inter7));
  inv1  gate765(.a(G1225), .O(gate481inter8));
  nand2 gate766(.a(gate481inter8), .b(gate481inter7), .O(gate481inter9));
  nand2 gate767(.a(s_31), .b(gate481inter3), .O(gate481inter10));
  nor2  gate768(.a(gate481inter10), .b(gate481inter9), .O(gate481inter11));
  nor2  gate769(.a(gate481inter11), .b(gate481inter6), .O(gate481inter12));
  nand2 gate770(.a(gate481inter12), .b(gate481inter1), .O(G1290));
nand2 gate482( .a(G1129), .b(G1225), .O(G1291) );

  xor2  gate925(.a(G1229), .b(G1228), .O(gate483inter0));
  nand2 gate926(.a(gate483inter0), .b(s_54), .O(gate483inter1));
  and2  gate927(.a(G1229), .b(G1228), .O(gate483inter2));
  inv1  gate928(.a(s_54), .O(gate483inter3));
  inv1  gate929(.a(s_55), .O(gate483inter4));
  nand2 gate930(.a(gate483inter4), .b(gate483inter3), .O(gate483inter5));
  nor2  gate931(.a(gate483inter5), .b(gate483inter2), .O(gate483inter6));
  inv1  gate932(.a(G1228), .O(gate483inter7));
  inv1  gate933(.a(G1229), .O(gate483inter8));
  nand2 gate934(.a(gate483inter8), .b(gate483inter7), .O(gate483inter9));
  nand2 gate935(.a(s_55), .b(gate483inter3), .O(gate483inter10));
  nor2  gate936(.a(gate483inter10), .b(gate483inter9), .O(gate483inter11));
  nor2  gate937(.a(gate483inter11), .b(gate483inter6), .O(gate483inter12));
  nand2 gate938(.a(gate483inter12), .b(gate483inter1), .O(G1292));
nand2 gate484( .a(G1230), .b(G1231), .O(G1293) );

  xor2  gate1317(.a(G1233), .b(G1232), .O(gate485inter0));
  nand2 gate1318(.a(gate485inter0), .b(s_110), .O(gate485inter1));
  and2  gate1319(.a(G1233), .b(G1232), .O(gate485inter2));
  inv1  gate1320(.a(s_110), .O(gate485inter3));
  inv1  gate1321(.a(s_111), .O(gate485inter4));
  nand2 gate1322(.a(gate485inter4), .b(gate485inter3), .O(gate485inter5));
  nor2  gate1323(.a(gate485inter5), .b(gate485inter2), .O(gate485inter6));
  inv1  gate1324(.a(G1232), .O(gate485inter7));
  inv1  gate1325(.a(G1233), .O(gate485inter8));
  nand2 gate1326(.a(gate485inter8), .b(gate485inter7), .O(gate485inter9));
  nand2 gate1327(.a(s_111), .b(gate485inter3), .O(gate485inter10));
  nor2  gate1328(.a(gate485inter10), .b(gate485inter9), .O(gate485inter11));
  nor2  gate1329(.a(gate485inter11), .b(gate485inter6), .O(gate485inter12));
  nand2 gate1330(.a(gate485inter12), .b(gate485inter1), .O(G1294));
nand2 gate486( .a(G1234), .b(G1235), .O(G1295) );

  xor2  gate1051(.a(G1237), .b(G1236), .O(gate487inter0));
  nand2 gate1052(.a(gate487inter0), .b(s_72), .O(gate487inter1));
  and2  gate1053(.a(G1237), .b(G1236), .O(gate487inter2));
  inv1  gate1054(.a(s_72), .O(gate487inter3));
  inv1  gate1055(.a(s_73), .O(gate487inter4));
  nand2 gate1056(.a(gate487inter4), .b(gate487inter3), .O(gate487inter5));
  nor2  gate1057(.a(gate487inter5), .b(gate487inter2), .O(gate487inter6));
  inv1  gate1058(.a(G1236), .O(gate487inter7));
  inv1  gate1059(.a(G1237), .O(gate487inter8));
  nand2 gate1060(.a(gate487inter8), .b(gate487inter7), .O(gate487inter9));
  nand2 gate1061(.a(s_73), .b(gate487inter3), .O(gate487inter10));
  nor2  gate1062(.a(gate487inter10), .b(gate487inter9), .O(gate487inter11));
  nor2  gate1063(.a(gate487inter11), .b(gate487inter6), .O(gate487inter12));
  nand2 gate1064(.a(gate487inter12), .b(gate487inter1), .O(G1296));

  xor2  gate1121(.a(G1239), .b(G1238), .O(gate488inter0));
  nand2 gate1122(.a(gate488inter0), .b(s_82), .O(gate488inter1));
  and2  gate1123(.a(G1239), .b(G1238), .O(gate488inter2));
  inv1  gate1124(.a(s_82), .O(gate488inter3));
  inv1  gate1125(.a(s_83), .O(gate488inter4));
  nand2 gate1126(.a(gate488inter4), .b(gate488inter3), .O(gate488inter5));
  nor2  gate1127(.a(gate488inter5), .b(gate488inter2), .O(gate488inter6));
  inv1  gate1128(.a(G1238), .O(gate488inter7));
  inv1  gate1129(.a(G1239), .O(gate488inter8));
  nand2 gate1130(.a(gate488inter8), .b(gate488inter7), .O(gate488inter9));
  nand2 gate1131(.a(s_83), .b(gate488inter3), .O(gate488inter10));
  nor2  gate1132(.a(gate488inter10), .b(gate488inter9), .O(gate488inter11));
  nor2  gate1133(.a(gate488inter11), .b(gate488inter6), .O(gate488inter12));
  nand2 gate1134(.a(gate488inter12), .b(gate488inter1), .O(G1297));

  xor2  gate561(.a(G1241), .b(G1240), .O(gate489inter0));
  nand2 gate562(.a(gate489inter0), .b(s_2), .O(gate489inter1));
  and2  gate563(.a(G1241), .b(G1240), .O(gate489inter2));
  inv1  gate564(.a(s_2), .O(gate489inter3));
  inv1  gate565(.a(s_3), .O(gate489inter4));
  nand2 gate566(.a(gate489inter4), .b(gate489inter3), .O(gate489inter5));
  nor2  gate567(.a(gate489inter5), .b(gate489inter2), .O(gate489inter6));
  inv1  gate568(.a(G1240), .O(gate489inter7));
  inv1  gate569(.a(G1241), .O(gate489inter8));
  nand2 gate570(.a(gate489inter8), .b(gate489inter7), .O(gate489inter9));
  nand2 gate571(.a(s_3), .b(gate489inter3), .O(gate489inter10));
  nor2  gate572(.a(gate489inter10), .b(gate489inter9), .O(gate489inter11));
  nor2  gate573(.a(gate489inter11), .b(gate489inter6), .O(gate489inter12));
  nand2 gate574(.a(gate489inter12), .b(gate489inter1), .O(G1298));
nand2 gate490( .a(G1242), .b(G1243), .O(G1299) );
nand2 gate491( .a(G1244), .b(G1245), .O(G1300) );
nand2 gate492( .a(G1246), .b(G1247), .O(G1301) );

  xor2  gate1135(.a(G1249), .b(G1248), .O(gate493inter0));
  nand2 gate1136(.a(gate493inter0), .b(s_84), .O(gate493inter1));
  and2  gate1137(.a(G1249), .b(G1248), .O(gate493inter2));
  inv1  gate1138(.a(s_84), .O(gate493inter3));
  inv1  gate1139(.a(s_85), .O(gate493inter4));
  nand2 gate1140(.a(gate493inter4), .b(gate493inter3), .O(gate493inter5));
  nor2  gate1141(.a(gate493inter5), .b(gate493inter2), .O(gate493inter6));
  inv1  gate1142(.a(G1248), .O(gate493inter7));
  inv1  gate1143(.a(G1249), .O(gate493inter8));
  nand2 gate1144(.a(gate493inter8), .b(gate493inter7), .O(gate493inter9));
  nand2 gate1145(.a(s_85), .b(gate493inter3), .O(gate493inter10));
  nor2  gate1146(.a(gate493inter10), .b(gate493inter9), .O(gate493inter11));
  nor2  gate1147(.a(gate493inter11), .b(gate493inter6), .O(gate493inter12));
  nand2 gate1148(.a(gate493inter12), .b(gate493inter1), .O(G1302));
nand2 gate494( .a(G1250), .b(G1251), .O(G1303) );
nand2 gate495( .a(G1252), .b(G1253), .O(G1304) );
nand2 gate496( .a(G1254), .b(G1255), .O(G1305) );
nand2 gate497( .a(G1256), .b(G1257), .O(G1306) );
nand2 gate498( .a(G1258), .b(G1259), .O(G1307) );
nand2 gate499( .a(G1260), .b(G1261), .O(G1308) );
nand2 gate500( .a(G1262), .b(G1263), .O(G1309) );
nand2 gate501( .a(G1264), .b(G1265), .O(G1310) );
nand2 gate502( .a(G1266), .b(G1267), .O(G1311) );
nand2 gate503( .a(G1268), .b(G1269), .O(G1312) );

  xor2  gate1303(.a(G1271), .b(G1270), .O(gate504inter0));
  nand2 gate1304(.a(gate504inter0), .b(s_108), .O(gate504inter1));
  and2  gate1305(.a(G1271), .b(G1270), .O(gate504inter2));
  inv1  gate1306(.a(s_108), .O(gate504inter3));
  inv1  gate1307(.a(s_109), .O(gate504inter4));
  nand2 gate1308(.a(gate504inter4), .b(gate504inter3), .O(gate504inter5));
  nor2  gate1309(.a(gate504inter5), .b(gate504inter2), .O(gate504inter6));
  inv1  gate1310(.a(G1270), .O(gate504inter7));
  inv1  gate1311(.a(G1271), .O(gate504inter8));
  nand2 gate1312(.a(gate504inter8), .b(gate504inter7), .O(gate504inter9));
  nand2 gate1313(.a(s_109), .b(gate504inter3), .O(gate504inter10));
  nor2  gate1314(.a(gate504inter10), .b(gate504inter9), .O(gate504inter11));
  nor2  gate1315(.a(gate504inter11), .b(gate504inter6), .O(gate504inter12));
  nand2 gate1316(.a(gate504inter12), .b(gate504inter1), .O(G1313));
nand2 gate505( .a(G1272), .b(G1273), .O(G1314) );

  xor2  gate1373(.a(G1275), .b(G1274), .O(gate506inter0));
  nand2 gate1374(.a(gate506inter0), .b(s_118), .O(gate506inter1));
  and2  gate1375(.a(G1275), .b(G1274), .O(gate506inter2));
  inv1  gate1376(.a(s_118), .O(gate506inter3));
  inv1  gate1377(.a(s_119), .O(gate506inter4));
  nand2 gate1378(.a(gate506inter4), .b(gate506inter3), .O(gate506inter5));
  nor2  gate1379(.a(gate506inter5), .b(gate506inter2), .O(gate506inter6));
  inv1  gate1380(.a(G1274), .O(gate506inter7));
  inv1  gate1381(.a(G1275), .O(gate506inter8));
  nand2 gate1382(.a(gate506inter8), .b(gate506inter7), .O(gate506inter9));
  nand2 gate1383(.a(s_119), .b(gate506inter3), .O(gate506inter10));
  nor2  gate1384(.a(gate506inter10), .b(gate506inter9), .O(gate506inter11));
  nor2  gate1385(.a(gate506inter11), .b(gate506inter6), .O(gate506inter12));
  nand2 gate1386(.a(gate506inter12), .b(gate506inter1), .O(G1315));
nand2 gate507( .a(G1276), .b(G1277), .O(G1316) );
nand2 gate508( .a(G1278), .b(G1279), .O(G1317) );
nand2 gate509( .a(G1280), .b(G1281), .O(G1318) );
nand2 gate510( .a(G1282), .b(G1283), .O(G1319) );
nand2 gate511( .a(G1284), .b(G1285), .O(G1320) );

  xor2  gate687(.a(G1287), .b(G1286), .O(gate512inter0));
  nand2 gate688(.a(gate512inter0), .b(s_20), .O(gate512inter1));
  and2  gate689(.a(G1287), .b(G1286), .O(gate512inter2));
  inv1  gate690(.a(s_20), .O(gate512inter3));
  inv1  gate691(.a(s_21), .O(gate512inter4));
  nand2 gate692(.a(gate512inter4), .b(gate512inter3), .O(gate512inter5));
  nor2  gate693(.a(gate512inter5), .b(gate512inter2), .O(gate512inter6));
  inv1  gate694(.a(G1286), .O(gate512inter7));
  inv1  gate695(.a(G1287), .O(gate512inter8));
  nand2 gate696(.a(gate512inter8), .b(gate512inter7), .O(gate512inter9));
  nand2 gate697(.a(s_21), .b(gate512inter3), .O(gate512inter10));
  nor2  gate698(.a(gate512inter10), .b(gate512inter9), .O(gate512inter11));
  nor2  gate699(.a(gate512inter11), .b(gate512inter6), .O(gate512inter12));
  nand2 gate700(.a(gate512inter12), .b(gate512inter1), .O(G1321));
nand2 gate513( .a(G1288), .b(G1289), .O(G1322) );

  xor2  gate1555(.a(G1291), .b(G1290), .O(gate514inter0));
  nand2 gate1556(.a(gate514inter0), .b(s_144), .O(gate514inter1));
  and2  gate1557(.a(G1291), .b(G1290), .O(gate514inter2));
  inv1  gate1558(.a(s_144), .O(gate514inter3));
  inv1  gate1559(.a(s_145), .O(gate514inter4));
  nand2 gate1560(.a(gate514inter4), .b(gate514inter3), .O(gate514inter5));
  nor2  gate1561(.a(gate514inter5), .b(gate514inter2), .O(gate514inter6));
  inv1  gate1562(.a(G1290), .O(gate514inter7));
  inv1  gate1563(.a(G1291), .O(gate514inter8));
  nand2 gate1564(.a(gate514inter8), .b(gate514inter7), .O(gate514inter9));
  nand2 gate1565(.a(s_145), .b(gate514inter3), .O(gate514inter10));
  nor2  gate1566(.a(gate514inter10), .b(gate514inter9), .O(gate514inter11));
  nor2  gate1567(.a(gate514inter11), .b(gate514inter6), .O(gate514inter12));
  nand2 gate1568(.a(gate514inter12), .b(gate514inter1), .O(G1323));
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule