module c7552 (N1,N5,N9,N12,N15,N18,N23,N26,N29,N32,
              N35,N38,N41,N44,N47,N50,N53,N54,N55,N56,
              N57,N58,N59,N60,N61,N62,N63,N64,N65,N66,
              N69,N70,N73,N74,N75,N76,N77,N78,N79,N80,
              N81,N82,N83,N84,N85,N86,N87,N88,N89,N94,
              N97,N100,N103,N106,N109,N110,N111,N112,N113,N114,
              N115,N118,N121,N124,N127,N130,N133,N134,N135,N138,
              N141,N144,N147,N150,N151,N152,N153,N154,N155,N156,
              N157,N158,N159,N160,N161,N162,N163,N164,N165,N166,
              N167,N168,N169,N170,N171,N172,N173,N174,N175,N176,
              N177,N178,N179,N180,N181,N182,N183,N184,N185,N186,
              N187,N188,N189,N190,N191,N192,N193,N194,N195,N196,
              N197,N198,N199,N200,N201,N202,N203,N204,N205,N206,
              N207,N208,N209,N210,N211,N212,N213,N214,N215,N216,
              N217,N218,N219,N220,N221,N222,N223,N224,N225,N226,
              N227,N228,N229,N230,N231,N232,N233,N234,N235,N236,
              N237,N238,N239,N240,N242,N245,N248,N251,N254,N257,
              N260,N263,N267,N271,N274,N277,N280,N283,N286,N289,
              N293,N296,N299,N303,N307,N310,N313,N316,N319,N322,
              N325,N328,N331,N334,N337,N340,N343,N346,N349,N352,
              N355,N358,N361,N364,N367,N382,N241_I,N387,N388,N478,
              N482,N484,N486,N489,N492,N501,N505,N507,N509,N511,
              N513,N515,N517,N519,N535,N537,N539,N541,N543,N545,
              N547,N549,N551,N553,N556,N559,N561,N563,N565,N567,
              N569,N571,N573,N582,N643,N707,N813,N881,N882,N883,
              N884,N885,N889,N945,N1110,N1111,N1112,N1113,N1114,N1489,
              N1490,N1781,N10025,N10101,N10102,N10103,N10104,N10109,N10110,N10111,
              N10112,N10350,N10351,N10352,N10353,N10574,N10575,N10576,N10628,N10632,
              N10641,N10704,N10706,N10711,N10712,N10713,N10714,N10715,N10716,N10717,
              N10718,N10729,N10759,N10760,N10761,N10762,N10763,N10827,N10837,N10838,
              N10839,N10840,N10868,N10869,N10870,N10871,N10905,N10906,N10907,N10908,
              N11333,N11334,N11340,N11342,N241_O);

input N1,N5,N9,N12,N15,N18,N23,N26,N29,N32,
      N35,N38,N41,N44,N47,N50,N53,N54,N55,N56,
      N57,N58,N59,N60,N61,N62,N63,N64,N65,N66,
      N69,N70,N73,N74,N75,N76,N77,N78,N79,N80,
      N81,N82,N83,N84,N85,N86,N87,N88,N89,N94,
      N97,N100,N103,N106,N109,N110,N111,N112,N113,N114,
      N115,N118,N121,N124,N127,N130,N133,N134,N135,N138,
      N141,N144,N147,N150,N151,N152,N153,N154,N155,N156,
      N157,N158,N159,N160,N161,N162,N163,N164,N165,N166,
      N167,N168,N169,N170,N171,N172,N173,N174,N175,N176,
      N177,N178,N179,N180,N181,N182,N183,N184,N185,N186,
      N187,N188,N189,N190,N191,N192,N193,N194,N195,N196,
      N197,N198,N199,N200,N201,N202,N203,N204,N205,N206,
      N207,N208,N209,N210,N211,N212,N213,N214,N215,N216,
      N217,N218,N219,N220,N221,N222,N223,N224,N225,N226,
      N227,N228,N229,N230,N231,N232,N233,N234,N235,N236,
      N237,N238,N239,N240,N242,N245,N248,N251,N254,N257,
      N260,N263,N267,N271,N274,N277,N280,N283,N286,N289,
      N293,N296,N299,N303,N307,N310,N313,N316,N319,N322,
      N325,N328,N331,N334,N337,N340,N343,N346,N349,N352,
      N355,N358,N361,N364,N367,N382,N241_I;//RE__PI;

input s_0,s_1;//RE__ALLOW(00,01,10,11);
input s_2,s_3;//RE__ALLOW(00,01,10,11);
input s_4,s_5;//RE__ALLOW(00,01,10,11);
input s_6,s_7;//RE__ALLOW(00,01,10,11);
input s_8,s_9;//RE__ALLOW(00,01,10,11);
input s_10,s_11;//RE__ALLOW(00,01,10,11);
input s_12,s_13;//RE__ALLOW(00,01,10,11);
input s_14,s_15;//RE__ALLOW(00,01,10,11);
input s_16,s_17;//RE__ALLOW(00,01,10,11);
input s_18,s_19;//RE__ALLOW(00,01,10,11);
input s_20,s_21;//RE__ALLOW(00,01,10,11);
input s_22,s_23;//RE__ALLOW(00,01,10,11);
input s_24,s_25;//RE__ALLOW(00,01,10,11);
input s_26,s_27;//RE__ALLOW(00,01,10,11);
input s_28,s_29;//RE__ALLOW(00,01,10,11);
input s_30,s_31;//RE__ALLOW(00,01,10,11);
input s_32,s_33;//RE__ALLOW(00,01,10,11);
input s_34,s_35;//RE__ALLOW(00,01,10,11);
input s_36,s_37;//RE__ALLOW(00,01,10,11);
input s_38,s_39;//RE__ALLOW(00,01,10,11);
input s_40,s_41;//RE__ALLOW(00,01,10,11);
input s_42,s_43;//RE__ALLOW(00,01,10,11);
input s_44,s_45;//RE__ALLOW(00,01,10,11);
input s_46,s_47;//RE__ALLOW(00,01,10,11);
input s_48,s_49;//RE__ALLOW(00,01,10,11);
input s_50,s_51;//RE__ALLOW(00,01,10,11);
input s_52,s_53;//RE__ALLOW(00,01,10,11);
input s_54,s_55;//RE__ALLOW(00,01,10,11);
input s_56,s_57;//RE__ALLOW(00,01,10,11);
input s_58,s_59;//RE__ALLOW(00,01,10,11);
input s_60,s_61;//RE__ALLOW(00,01,10,11);
input s_62,s_63;//RE__ALLOW(00,01,10,11);
input s_64,s_65;//RE__ALLOW(00,01,10,11);
input s_66,s_67;//RE__ALLOW(00,01,10,11);
input s_68,s_69;//RE__ALLOW(00,01,10,11);
input s_70,s_71;//RE__ALLOW(00,01,10,11);
input s_72,s_73;//RE__ALLOW(00,01,10,11);
input s_74,s_75;//RE__ALLOW(00,01,10,11);
input s_76,s_77;//RE__ALLOW(00,01,10,11);
input s_78,s_79;//RE__ALLOW(00,01,10,11);
input s_80,s_81;//RE__ALLOW(00,01,10,11);
input s_82,s_83;//RE__ALLOW(00,01,10,11);
input s_84,s_85;//RE__ALLOW(00,01,10,11);
input s_86,s_87;//RE__ALLOW(00,01,10,11);
input s_88,s_89;//RE__ALLOW(00,01,10,11);
input s_90,s_91;//RE__ALLOW(00,01,10,11);
input s_92,s_93;//RE__ALLOW(00,01,10,11);
input s_94,s_95;//RE__ALLOW(00,01,10,11);
input s_96,s_97;//RE__ALLOW(00,01,10,11);
input s_98,s_99;//RE__ALLOW(00,01,10,11);
input s_100,s_101;//RE__ALLOW(00,01,10,11);
input s_102,s_103;//RE__ALLOW(00,01,10,11);
input s_104,s_105;//RE__ALLOW(00,01,10,11);
input s_106,s_107;//RE__ALLOW(00,01,10,11);
input s_108,s_109;//RE__ALLOW(00,01,10,11);
input s_110,s_111;//RE__ALLOW(00,01,10,11);
input s_112,s_113;//RE__ALLOW(00,01,10,11);
input s_114,s_115;//RE__ALLOW(00,01,10,11);
input s_116,s_117;//RE__ALLOW(00,01,10,11);
input s_118,s_119;//RE__ALLOW(00,01,10,11);
input s_120,s_121;//RE__ALLOW(00,01,10,11);
input s_122,s_123;//RE__ALLOW(00,01,10,11);
input s_124,s_125;//RE__ALLOW(00,01,10,11);
input s_126,s_127;//RE__ALLOW(00,01,10,11);
input s_128,s_129;//RE__ALLOW(00,01,10,11);
input s_130,s_131;//RE__ALLOW(00,01,10,11);
input s_132,s_133;//RE__ALLOW(00,01,10,11);
input s_134,s_135;//RE__ALLOW(00,01,10,11);
input s_136,s_137;//RE__ALLOW(00,01,10,11);
input s_138,s_139;//RE__ALLOW(00,01,10,11);
input s_140,s_141;//RE__ALLOW(00,01,10,11);
input s_142,s_143;//RE__ALLOW(00,01,10,11);
input s_144,s_145;//RE__ALLOW(00,01,10,11);
input s_146,s_147;//RE__ALLOW(00,01,10,11);
input s_148,s_149;//RE__ALLOW(00,01,10,11);
input s_150,s_151;//RE__ALLOW(00,01,10,11);
input s_152,s_153;//RE__ALLOW(00,01,10,11);
input s_154,s_155;//RE__ALLOW(00,01,10,11);
input s_156,s_157;//RE__ALLOW(00,01,10,11);
input s_158,s_159;//RE__ALLOW(00,01,10,11);
input s_160,s_161;//RE__ALLOW(00,01,10,11);
input s_162,s_163;//RE__ALLOW(00,01,10,11);
input s_164,s_165;//RE__ALLOW(00,01,10,11);
input s_166,s_167;//RE__ALLOW(00,01,10,11);
input s_168,s_169;//RE__ALLOW(00,01,10,11);
input s_170,s_171;//RE__ALLOW(00,01,10,11);
input s_172,s_173;//RE__ALLOW(00,01,10,11);
input s_174,s_175;//RE__ALLOW(00,01,10,11);
input s_176,s_177;//RE__ALLOW(00,01,10,11);
input s_178,s_179;//RE__ALLOW(00,01,10,11);
input s_180,s_181;//RE__ALLOW(00,01,10,11);
input s_182,s_183;//RE__ALLOW(00,01,10,11);
input s_184,s_185;//RE__ALLOW(00,01,10,11);
input s_186,s_187;//RE__ALLOW(00,01,10,11);
input s_188,s_189;//RE__ALLOW(00,01,10,11);
input s_190,s_191;//RE__ALLOW(00,01,10,11);
input s_192,s_193;//RE__ALLOW(00,01,10,11);
input s_194,s_195;//RE__ALLOW(00,01,10,11);
input s_196,s_197;//RE__ALLOW(00,01,10,11);
input s_198,s_199;//RE__ALLOW(00,01,10,11);
input s_200,s_201;//RE__ALLOW(00,01,10,11);
input s_202,s_203;//RE__ALLOW(00,01,10,11);
input s_204,s_205;//RE__ALLOW(00,01,10,11);
input s_206,s_207;//RE__ALLOW(00,01,10,11);
input s_208,s_209;//RE__ALLOW(00,01,10,11);
input s_210,s_211;//RE__ALLOW(00,01,10,11);
input s_212,s_213;//RE__ALLOW(00,01,10,11);
input s_214,s_215;//RE__ALLOW(00,01,10,11);
input s_216,s_217;//RE__ALLOW(00,01,10,11);
input s_218,s_219;//RE__ALLOW(00,01,10,11);
input s_220,s_221;//RE__ALLOW(00,01,10,11);
input s_222,s_223;//RE__ALLOW(00,01,10,11);
input s_224,s_225;//RE__ALLOW(00,01,10,11);
input s_226,s_227;//RE__ALLOW(00,01,10,11);
input s_228,s_229;//RE__ALLOW(00,01,10,11);
input s_230,s_231;//RE__ALLOW(00,01,10,11);
input s_232,s_233;//RE__ALLOW(00,01,10,11);
input s_234,s_235;//RE__ALLOW(00,01,10,11);
input s_236,s_237;//RE__ALLOW(00,01,10,11);
input s_238,s_239;//RE__ALLOW(00,01,10,11);
input s_240,s_241;//RE__ALLOW(00,01,10,11);
input s_242,s_243;//RE__ALLOW(00,01,10,11);
input s_244,s_245;//RE__ALLOW(00,01,10,11);
input s_246,s_247;//RE__ALLOW(00,01,10,11);
input s_248,s_249;//RE__ALLOW(00,01,10,11);
input s_250,s_251;//RE__ALLOW(00,01,10,11);
input s_252,s_253;//RE__ALLOW(00,01,10,11);
input s_254,s_255;//RE__ALLOW(00,01,10,11);
input s_256,s_257;//RE__ALLOW(00,01,10,11);
input s_258,s_259;//RE__ALLOW(00,01,10,11);
input s_260,s_261;//RE__ALLOW(00,01,10,11);
output N387,N388,N478,N482,N484,N486,N489,N492,N501,N505,
       N507,N509,N511,N513,N515,N517,N519,N535,N537,N539,
       N541,N543,N545,N547,N549,N551,N553,N556,N559,N561,
       N563,N565,N567,N569,N571,N573,N582,N643,N707,N813,
       N881,N882,N883,N884,N885,N889,N945,N1110,N1111,N1112,
       N1113,N1114,N1489,N1490,N1781,N10025,N10101,N10102,N10103,N10104,
       N10109,N10110,N10111,N10112,N10350,N10351,N10352,N10353,N10574,N10575,
       N10576,N10628,N10632,N10641,N10704,N10706,N10711,N10712,N10713,N10714,
       N10715,N10716,N10717,N10718,N10729,N10759,N10760,N10761,N10762,N10763,
       N10827,N10837,N10838,N10839,N10840,N10868,N10869,N10870,N10871,N10905,
       N10906,N10907,N10908,N11333,N11334,N11340,N11342,N241_O;

wire N467,N469,N494,N528,N575,N578,N585,N590,N593,N596,
     N599,N604,N609,N614,N625,N628,N632,N636,N641,N642,
     N644,N651,N657,N660,N666,N672,N673,N674,N676,N682,
     N688,N689,N695,N700,N705,N706,N708,N715,N721,N727,
     N733,N734,N742,N748,N749,N750,N758,N759,N762,N768,
     N774,N780,N786,N794,N800,N806,N812,N814,N821,N827,
     N833,N839,N845,N853,N859,N865,N871,N886,N887,N957,
     N1028,N1029,N1109,N1115,N1116,N1119,N1125,N1132,N1136,N1141,
     N1147,N1154,N1160,N1167,N1174,N1175,N1182,N1189,N1194,N1199,
     N1206,N1211,N1218,N1222,N1227,N1233,N1240,N1244,N1249,N1256,
     N1263,N1270,N1277,N1284,N1287,N1290,N1293,N1296,N1299,N1302,
     N1305,N1308,N1311,N1314,N1317,N1320,N1323,N1326,N1329,N1332,
     N1335,N1338,N1341,N1344,N1347,N1350,N1353,N1356,N1359,N1362,
     N1365,N1368,N1371,N1374,N1377,N1380,N1383,N1386,N1389,N1392,
     N1395,N1398,N1401,N1404,N1407,N1410,N1413,N1416,N1419,N1422,
     N1425,N1428,N1431,N1434,N1437,N1440,N1443,N1446,N1449,N1452,
     N1455,N1458,N1461,N1464,N1467,N1470,N1473,N1476,N1479,N1482,
     N1485,N1537,N1551,N1649,N1703,N1708,N1713,N1721,N1758,N1782,
     N1783,N1789,N1793,N1794,N1795,N1796,N1797,N1798,N1799,N1805,
     N1811,N1812,N1813,N1814,N1815,N1816,N1817,N1818,N1819,N1820,
     N1821,N1822,N1828,N1829,N1830,N1832,N1833,N1834,N1835,N1839,
     N1840,N1841,N1842,N1843,N1845,N1851,N1857,N1858,N1859,N1860,
     N1861,N1862,N1863,N1864,N1865,N1866,N1867,N1868,N1869,N1870,
     N1871,N1872,N1873,N1874,N1875,N1876,N1877,N1878,N1879,N1880,
     N1881,N1882,N1883,N1884,N1885,N1892,N1899,N1906,N1913,N1919,
     N1926,N1927,N1928,N1929,N1930,N1931,N1932,N1933,N1934,N1935,
     N1936,N1937,N1938,N1939,N1940,N1941,N1942,N1943,N1944,N1945,
     N1946,N1947,N1953,N1957,N1958,N1959,N1960,N1961,N1962,N1963,
     N1965,N1966,N1967,N1968,N1969,N1970,N1971,N1972,N1973,N1974,
     N1975,N1976,N1977,N1983,N1989,N1990,N1991,N1992,N1993,N1994,
     N1995,N1996,N1997,N2003,N2010,N2011,N2012,N2013,N2014,N2015,
     N2016,N2017,N2018,N2019,N2020,N2021,N2022,N2023,N2024,N2031,
     N2038,N2045,N2052,N2058,N2064,N2065,N2066,N2067,N2068,N2069,
     N2070,N2071,N2072,N2073,N2074,N2081,N2086,N2107,N2108,N2110,
     N2111,N2112,N2113,N2114,N2115,N2117,N2171,N2172,N2230,N2231,
     N2235,N2239,N2240,N2241,N2242,N2243,N2244,N2245,N2246,N2247,
     N2248,N2249,N2250,N2251,N2252,N2253,N2254,N2255,N2256,N2257,
     N2267,N2268,N2269,N2274,N2275,N2277,N2278,N2279,N2280,N2281,
     N2282,N2283,N2284,N2285,N2286,N2287,N2293,N2299,N2300,N2301,
     N2302,N2303,N2304,N2305,N2306,N2307,N2308,N2309,N2315,N2321,
     N2322,N2323,N2324,N2325,N2326,N2327,N2328,N2329,N2330,N2331,
     N2337,N2338,N2339,N2340,N2341,N2342,N2343,N2344,N2345,N2346,
     N2347,N2348,N2349,N2350,N2351,N2352,N2353,N2354,N2355,N2356,
     N2357,N2358,N2359,N2360,N2361,N2362,N2363,N2364,N2365,N2366,
     N2367,N2368,N2374,N2375,N2376,N2377,N2378,N2379,N2380,N2381,
     N2382,N2383,N2384,N2390,N2396,N2397,N2398,N2399,N2400,N2401,
     N2402,N2403,N2404,N2405,N2406,N2412,N2418,N2419,N2420,N2421,
     N2422,N2423,N2424,N2425,N2426,N2427,N2428,N2429,N2430,N2431,
     N2432,N2433,N2434,N2435,N2436,N2437,N2441,N2442,N2446,N2450,
     N2454,N2458,N2462,N2466,N2470,N2474,N2478,N2482,N2488,N2496,
     N2502,N2508,N2523,N2533,N2537,N2538,N2542,N2546,N2550,N2554,
     N2561,N2567,N2573,N2604,N2607,N2611,N2615,N2619,N2626,N2632,
     N2638,N2644,N2650,N2653,N2654,N2658,N2662,N2666,N2670,N2674,
     N2680,N2688,N2692,N2696,N2700,N2704,N2728,N2729,N2733,N2737,
     N2741,N2745,N2749,N2753,N2757,N2761,N2765,N2766,N2769,N2772,
     N2775,N2778,N2781,N2784,N2787,N2790,N2793,N2796,N2866,N2867,
     N2868,N2869,N2878,N2913,N2914,N2915,N2916,N2917,N2918,N2919,
     N2920,N2921,N2922,N2923,N2924,N2925,N2926,N2927,N2928,N2929,
     N2930,N2931,N2932,N2933,N2934,N2935,N2936,N2937,N2988,N3005,
     N3006,N3007,N3008,N3009,N3020,N3021,N3022,N3023,N3024,N3025,
     N3026,N3027,N3028,N3029,N3032,N3033,N3034,N3035,N3036,N3037,
     N3038,N3039,N3040,N3041,N3061,N3064,N3067,N3070,N3073,N3080,
     N3096,N3097,N3101,N3107,N3114,N3122,N3126,N3130,N3131,N3134,
     N3135,N3136,N3137,N3140,N3144,N3149,N3155,N3159,N3167,N3168,
     N3169,N3173,N3178,N3184,N3185,N3189,N3195,N3202,N3210,N3211,
     N3215,N3221,N3228,N3229,N3232,N3236,N3241,N3247,N3251,N3255,
     N3259,N3263,N3267,N3273,N3281,N3287,N3293,N3299,N3303,N3307,
     N3311,N3315,N3322,N3328,N3334,N3340,N3343,N3349,N3355,N3361,
     N3362,N3363,N3364,N3365,N3366,N3367,N3368,N3369,N3370,N3371,
     N3372,N3373,N3374,N3375,N3379,N3380,N3381,N3384,N3390,N3398,
     N3404,N3410,N3416,N3420,N3424,N3428,N3432,N3436,N3440,N3444,
     N3448,N3452,N3453,N3454,N3458,N3462,N3466,N3470,N3474,N3478,
     N3482,N3486,N3487,N3490,N3493,N3496,N3499,N3502,N3507,N3510,
     N3515,N3518,N3521,N3524,N3527,N3530,N3535,N3539,N3542,N3545,
     N3548,N3551,N3552,N3553,N3557,N3560,N3563,N3566,N3569,N3570,
     N3571,N3574,N3577,N3580,N3583,N3586,N3589,N3592,N3595,N3598,
     N3601,N3604,N3607,N3610,N3613,N3616,N3619,N3622,N3625,N3628,
     N3631,N3634,N3637,N3640,N3643,N3646,N3649,N3652,N3655,N3658,
     N3661,N3664,N3667,N3670,N3673,N3676,N3679,N3682,N3685,N3688,
     N3691,N3694,N3697,N3700,N3703,N3706,N3709,N3712,N3715,N3718,
     N3721,N3724,N3727,N3730,N3733,N3736,N3739,N3742,N3745,N3748,
     N3751,N3754,N3757,N3760,N3763,N3766,N3769,N3772,N3775,N3778,
     N3781,N3782,N3783,N3786,N3789,N3792,N3795,N3798,N3801,N3804,
     N3807,N3810,N3813,N3816,N3819,N3822,N3825,N3828,N3831,N3834,
     N3837,N3840,N3843,N3846,N3849,N3852,N3855,N3858,N3861,N3864,
     N3867,N3870,N3873,N3876,N3879,N3882,N3885,N3888,N3891,N3953,
     N3954,N3955,N3956,N3958,N3964,N4193,N4303,N4308,N4313,N4326,
     N4327,N4333,N4334,N4411,N4412,N4463,N4464,N4465,N4466,N4467,
     N4468,N4469,N4470,N4471,N4472,N4473,N4474,N4475,N4476,N4477,
     N4478,N4479,N4480,N4481,N4482,N4483,N4484,N4485,N4486,N4487,
     N4488,N4489,N4490,N4491,N4492,N4493,N4494,N4495,N4496,N4497,
     N4498,N4499,N4500,N4501,N4502,N4503,N4504,N4505,N4506,N4507,
     N4508,N4509,N4510,N4511,N4512,N4513,N4514,N4515,N4516,N4517,
     N4518,N4519,N4520,N4521,N4522,N4523,N4524,N4525,N4526,N4527,
     N4528,N4529,N4530,N4531,N4532,N4533,N4534,N4535,N4536,N4537,
     N4538,N4539,N4540,N4541,N4542,N4543,N4544,N4545,N4549,N4555,
     N4562,N4563,N4566,N4570,N4575,N4576,N4577,N4581,N4586,N4592,
     N4593,N4597,N4603,N4610,N4611,N4612,N4613,N4614,N4615,N4616,
     N4617,N4618,N4619,N4620,N4621,N4622,N4623,N4624,N4625,N4626,
     N4627,N4628,N4629,N4630,N4631,N4632,N4633,N4634,N4635,N4636,
     N4637,N4638,N4639,N4640,N4641,N4642,N4643,N4644,N4645,N4646,
     N4647,N4648,N4649,N4650,N4651,N4652,N4653,N4656,N4657,N4661,
     N4667,N4674,N4675,N4678,N4682,N4687,N4693,N4694,N4695,N4696,
     N4697,N4698,N4699,N4700,N4701,N4702,N4706,N4711,N4717,N4718,
     N4722,N4728,N4735,N4743,N4744,N4745,N4746,N4747,N4748,N4749,
     N4750,N4751,N4752,N4753,N4754,N4755,N4756,N4757,N4758,N4759,
     N4760,N4761,N4762,N4763,N4764,N4765,N4766,N4767,N4768,N4769,
     N4775,N4776,N4777,N4778,N4779,N4780,N4781,N4782,N4783,N4784,
     N4789,N4790,N4793,N4794,N4795,N4796,N4799,N4800,N4801,N4802,
     N4803,N4806,N4809,N4810,N4813,N4814,N4817,N4820,N4823,N4826,
     N4829,N4832,N4835,N4838,N4841,N4844,N4847,N4850,N4853,N4856,
     N4859,N4862,N4865,N4868,N4871,N4874,N4877,N4880,N4883,N4886,
     N4889,N4892,N4895,N4898,N4901,N4904,N4907,N4910,N4913,N4916,
     N4919,N4922,N4925,N4928,N4931,N4934,N4937,N4940,N4943,N4946,
     N4949,N4952,N4955,N4958,N4961,N4964,N4967,N4970,N4973,N4976,
     N4979,N4982,N4985,N4988,N4991,N4994,N4997,N5000,N5003,N5006,
     N5009,N5012,N5015,N5018,N5021,N5024,N5027,N5030,N5033,N5036,
     N5039,N5042,N5045,N5046,N5047,N5048,N5049,N5052,N5055,N5058,
     N5061,N5064,N5065,N5066,N5067,N5068,N5071,N5074,N5077,N5080,
     N5083,N5086,N5089,N5092,N5095,N5098,N5101,N5104,N5107,N5110,
     N5111,N5112,N5113,N5114,N5117,N5120,N5123,N5126,N5129,N5132,
     N5135,N5138,N5141,N5144,N5147,N5150,N5153,N5156,N5159,N5162,
     N5165,N5166,N5167,N5168,N5169,N5170,N5171,N5172,N5173,N5174,
     N5175,N5176,N5177,N5178,N5179,N5180,N5181,N5182,N5183,N5184,
     N5185,N5186,N5187,N5188,N5189,N5190,N5191,N5192,N5193,N5196,
     N5197,N5198,N5199,N5200,N5201,N5202,N5203,N5204,N5205,N5206,
     N5207,N5208,N5209,N5210,N5211,N5212,N5213,N5283,N5284,N5285,
     N5286,N5287,N5288,N5289,N5290,N5291,N5292,N5293,N5294,N5295,
     N5296,N5297,N5298,N5299,N5300,N5314,N5315,N5316,N5317,N5318,
     N5319,N5320,N5321,N5322,N5323,N5324,N5363,N5364,N5365,N5366,
     N5367,N5425,N5426,N5427,N5429,N5430,N5431,N5432,N5433,N5451,
     N5452,N5453,N5454,N5455,N5456,N5457,N5469,N5474,N5475,N5476,
     N5477,N5571,N5572,N5573,N5574,N5584,N5585,N5586,N5587,N5602,
     N5603,N5604,N5605,N5631,N5632,N5640,N5654,N5670,N5683,N5690,
     N5697,N5707,N5718,N5728,N5735,N5736,N5740,N5744,N5747,N5751,
     N5755,N5758,N5762,N5766,N5769,N5770,N5771,N5778,N5789,N5799,
     N5807,N5821,N5837,N5850,N5856,N5863,N5870,N5881,N5892,N5898,
     N5905,N5915,N5926,N5936,N5943,N5944,N5945,N5946,N5947,N5948,
     N5949,N5950,N5951,N5952,N5953,N5954,N5955,N5956,N5957,N5958,
     N5959,N5960,N5966,N5967,N5968,N5969,N5970,N5971,N5972,N5973,
     N5974,N5975,N5976,N5977,N5978,N5979,N5980,N5981,N5989,N5990,
     N5991,N5996,N6000,N6003,N6009,N6014,N6018,N6021,N6022,N6023,
     N6024,N6025,N6026,N6027,N6028,N6029,N6030,N6031,N6032,N6033,
     N6034,N6035,N6036,N6037,N6038,N6039,N6040,N6041,N6047,N6052,
     N6056,N6059,N6060,N6061,N6062,N6063,N6064,N6065,N6066,N6067,
     N6068,N6069,N6070,N6071,N6072,N6073,N6074,N6075,N6076,N6077,
     N6078,N6079,N6083,N6087,N6090,N6091,N6092,N6093,N6094,N6095,
     N6096,N6097,N6098,N6099,N6100,N6101,N6102,N6103,N6104,N6105,
     N6106,N6107,N6108,N6109,N6110,N6111,N6112,N6113,N6114,N6115,
     N6116,N6117,N6118,N6119,N6120,N6121,N6122,N6123,N6124,N6125,
     N6126,N6127,N6131,N6135,N6136,N6137,N6141,N6145,N6148,N6149,
     N6150,N6151,N6152,N6153,N6154,N6155,N6156,N6157,N6158,N6159,
     N6160,N6161,N6162,N6163,N6164,N6165,N6166,N6170,N6174,N6177,
     N6181,N6182,N6183,N6184,N6185,N6186,N6187,N6188,N6189,N6190,
     N6191,N6192,N6193,N6194,N6195,N6196,N6199,N6202,N6203,N6204,
     N6207,N6210,N6213,N6214,N6217,N6220,N6223,N6224,N6225,N6226,
     N6227,N6228,N6229,N6230,N6231,N6232,N6235,N6236,N6239,N6240,
     N6241,N6242,N6243,N6246,N6249,N6252,N6255,N6256,N6257,N6258,
     N6259,N6260,N6261,N6262,N6263,N6266,N6540,N6541,N6542,N6543,
     N6544,N6545,N6546,N6547,N6555,N6556,N6557,N6558,N6559,N6560,
     N6561,N6569,N6594,N6595,N6596,N6597,N6598,N6599,N6600,N6601,
     N6602,N6603,N6604,N6605,N6606,N6621,N6622,N6623,N6624,N6625,
     N6626,N6627,N6628,N6629,N6639,N6640,N6641,N6642,N6643,N6644,
     N6645,N6646,N6647,N6648,N6649,N6650,N6651,N6652,N6653,N6654,
     N6655,N6656,N6657,N6658,N6659,N6660,N6661,N6668,N6677,N6678,
     N6679,N6680,N6681,N6682,N6683,N6684,N6685,N6686,N6687,N6688,
     N6689,N6690,N6702,N6703,N6704,N6705,N6706,N6707,N6708,N6709,
     N6710,N6711,N6712,N6729,N6730,N6731,N6732,N6733,N6734,N6735,
     N6736,N6741,N6742,N6743,N6744,N6751,N6752,N6753,N6754,N6755,
     N6756,N6757,N6758,N6761,N6762,N6766,N6767,N6768,N6769,N6770,
     N6771,N6772,N6773,N6774,N6775,N6776,N6777,N6778,N6779,N6780,
     N6781,N6782,N6783,N6784,N6787,N6788,N6789,N6790,N6791,N6792,
     N6793,N6794,N6795,N6796,N6797,N6800,N6803,N6806,N6809,N6812,
     N6815,N6818,N6821,N6824,N6827,N6830,N6833,N6836,N6837,N6838,
     N6839,N6840,N6841,N6842,N6843,N6844,N6845,N6848,N6849,N6850,
     N6851,N6852,N6853,N6854,N6855,N6856,N6857,N6858,N6859,N6860,
     N6861,N6862,N6863,N6864,N6865,N6866,N6867,N6870,N6871,N6872,
     N6873,N6874,N6875,N6876,N6877,N6878,N6879,N6880,N6881,N6884,
     N6885,N6886,N6887,N6888,N6889,N6890,N6891,N6892,N6893,N6894,
     N6901,N6912,N6923,N6929,N6936,N6946,N6957,N6967,N6968,N6969,
     N6970,N6977,N6988,N6998,N7006,N7020,N7036,N7049,N7055,N7056,
     N7057,N7060,N7061,N7062,N7063,N7064,N7065,N7066,N7067,N7068,
     N7073,N7077,N7080,N7086,N7091,N7095,N7098,N7099,N7100,N7103,
     N7104,N7105,N7106,N7107,N7114,N7125,N7136,N7142,N7149,N7159,
     N7170,N7180,N7187,N7188,N7191,N7194,N7198,N7202,N7205,N7209,
     N7213,N7216,N7219,N7222,N7229,N7240,N7250,N7258,N7272,N7288,
     N7301,N7307,N7314,N7318,N7322,N7325,N7328,N7331,N7334,N7337,
     N7340,N7343,N7346,N7351,N7355,N7358,N7364,N7369,N7373,N7376,
     N7377,N7378,N7381,N7384,N7387,N7391,N7394,N7398,N7402,N7405,
     N7408,N7411,N7414,N7417,N7420,N7423,N7426,N7429,N7432,N7435,
     N7438,N7441,N7444,N7447,N7450,N7453,N7456,N7459,N7462,N7465,
     N7468,N7471,N7474,N7477,N7478,N7479,N7482,N7485,N7488,N7491,
     N7494,N7497,N7500,N7503,N7506,N7509,N7512,N7515,N7518,N7521,
     N7524,N7527,N7530,N7533,N7536,N7539,N7542,N7545,N7548,N7551,
     N7552,N7553,N7556,N7557,N7558,N7559,N7560,N7563,N7566,N7569,
     N7572,N7573,N7574,N7577,N7580,N7581,N7582,N7585,N7588,N7591,
     N7609,N7613,N7620,N7649,N7650,N7655,N7659,N7668,N7671,N7744,
     N7822,N7825,N7826,N7852,N8114,N8117,N8131,N8134,N8144,N8145,
     N8146,N8156,N8166,N8169,N8183,N8186,N8196,N8200,N8204,N8208,
     N8216,N8217,N8218,N8219,N8232,N8233,N8242,N8243,N8244,N8245,
     N8246,N8247,N8248,N8249,N8250,N8251,N8252,N8253,N8254,N8260,
     N8261,N8262,N8269,N8274,N8275,N8276,N8277,N8278,N8279,N8280,
     N8281,N8282,N8283,N8284,N8285,N8288,N8294,N8295,N8296,N8297,
     N8298,N8307,N8315,N8317,N8319,N8321,N8322,N8323,N8324,N8325,
     N8326,N8333,N8337,N8338,N8339,N8340,N8341,N8342,N8343,N8344,
     N8345,N8346,N8347,N8348,N8349,N8350,N8351,N8352,N8353,N8354,
     N8355,N8356,N8357,N8358,N8365,N8369,N8370,N8371,N8372,N8373,
     N8374,N8375,N8376,N8377,N8378,N8379,N8380,N8381,N8382,N8383,
     N8384,N8385,N8386,N8387,N8388,N8389,N8390,N8391,N8392,N8393,
     N8394,N8404,N8405,N8409,N8410,N8411,N8412,N8415,N8416,N8417,
     N8418,N8421,N8430,N8433,N8434,N8435,N8436,N8437,N8438,N8439,
     N8440,N8441,N8442,N8443,N8444,N8447,N8448,N8449,N8450,N8451,
     N8452,N8453,N8454,N8455,N8456,N8457,N8460,N8463,N8466,N8469,
     N8470,N8471,N8474,N8477,N8480,N8483,N8484,N8485,N8488,N8489,
     N8490,N8491,N8492,N8493,N8494,N8495,N8496,N8497,N8500,N8501,
     N8502,N8503,N8504,N8505,N8506,N8507,N8508,N8509,N8510,N8511,
     N8512,N8513,N8514,N8515,N8516,N8517,N8518,N8519,N8522,N8525,
     N8528,N8531,N8534,N8537,N8538,N8539,N8540,N8541,N8545,N8546,
     N8547,N8548,N8551,N8552,N8553,N8554,N8555,N8558,N8561,N8564,
     N8565,N8566,N8569,N8572,N8575,N8578,N8579,N8580,N8583,N8586,
     N8589,N8592,N8595,N8598,N8601,N8604,N8607,N8608,N8609,N8610,
     N8615,N8616,N8617,N8618,N8619,N8624,N8625,N8626,N8627,N8632,
     N8633,N8634,N8637,N8638,N8639,N8644,N8645,N8646,N8647,N8648,
     N8653,N8654,N8655,N8660,N8663,N8666,N8669,N8672,N8675,N8678,
     N8681,N8684,N8687,N8690,N8693,N8696,N8699,N8702,N8705,N8708,
     N8711,N8714,N8717,N8718,N8721,N8724,N8727,N8730,N8733,N8734,
     N8735,N8738,N8741,N8744,N8747,N8750,N8753,N8754,N8755,N8756,
     N8757,N8760,N8763,N8766,N8769,N8772,N8775,N8778,N8781,N8784,
     N8787,N8790,N8793,N8796,N8799,N8802,N8805,N8808,N8811,N8814,
     N8815,N8816,N8817,N8818,N8840,N8857,N8861,N8862,N8863,N8864,
     N8865,N8866,N8871,N8874,N8878,N8879,N8880,N8881,N8882,N8883,
     N8884,N8885,N8886,N8887,N8888,N8898,N8902,N8920,N8924,N8927,
     N8931,N8943,N8950,N8956,N8959,N8960,N8963,N8966,N8991,N8992,
     N8995,N8996,N9001,N9005,N9024,N9025,N9029,N9035,N9053,N9054,
     N9064,N9065,N9066,N9067,N9068,N9071,N9072,N9073,N9074,N9077,
     N9079,N9082,N9083,N9086,N9087,N9088,N9089,N9092,N9093,N9094,
     N9095,N9098,N9099,N9103,N9107,N9111,N9117,N9127,N9146,N9149,
     N9159,N9160,N9161,N9165,N9169,N9173,N9179,N9180,N9181,N9182,
     N9183,N9193,N9203,N9206,N9220,N9223,N9234,N9235,N9236,N9237,
     N9238,N9242,N9243,N9244,N9245,N9246,N9247,N9248,N9249,N9250,
     N9251,N9252,N9256,N9257,N9258,N9259,N9260,N9261,N9262,N9265,
     N9268,N9271,N9272,N9273,N9274,N9275,N9276,N9280,N9285,N9286,
     N9287,N9288,N9290,N9292,N9294,N9296,N9297,N9298,N9299,N9300,
     N9301,N9307,N9314,N9315,N9318,N9319,N9320,N9321,N9322,N9323,
     N9324,N9326,N9332,N9339,N9344,N9352,N9354,N9356,N9358,N9359,
     N9360,N9361,N9362,N9363,N9364,N9365,N9366,N9367,N9368,N9369,
     N9370,N9371,N9372,N9375,N9381,N9382,N9383,N9384,N9385,N9392,
     N9393,N9394,N9395,N9396,N9397,N9398,N9399,N9400,N9401,N9402,
     N9407,N9408,N9412,N9413,N9414,N9415,N9416,N9417,N9418,N9419,
     N9420,N9421,N9422,N9423,N9426,N9429,N9432,N9435,N9442,N9445,
     N9454,N9455,N9456,N9459,N9460,N9461,N9462,N9465,N9466,N9467,
     N9468,N9473,N9476,N9477,N9478,N9485,N9488,N9493,N9494,N9495,
     N9498,N9499,N9500,N9505,N9506,N9507,N9508,N9509,N9514,N9515,
     N9516,N9517,N9520,N9526,N9531,N9539,N9540,N9541,N9543,N9551,
     N9555,N9556,N9557,N9560,N9561,N9562,N9563,N9564,N9565,N9566,
     N9567,N9568,N9569,N9570,N9571,N9575,N9579,N9581,N9582,N9585,
     N9591,N9592,N9593,N9594,N9595,N9596,N9597,N9598,N9599,N9600,
     N9601,N9602,N9603,N9604,N9605,N9608,N9611,N9612,N9613,N9614,
     N9615,N9616,N9617,N9618,N9621,N9622,N9623,N9624,N9626,N9629,
     N9632,N9635,N9642,N9645,N9646,N9649,N9650,N9653,N9656,N9659,
     N9660,N9661,N9662,N9663,N9666,N9667,N9670,N9671,N9674,N9675,
     N9678,N9679,N9682,N9685,N9690,N9691,N9692,N9695,N9698,N9702,
     N9707,N9710,N9711,N9714,N9715,N9716,N9717,N9720,N9721,N9722,
     N9723,N9726,N9727,N9732,N9733,N9734,N9735,N9736,N9737,N9738,
     N9739,N9740,N9741,N9742,N9754,N9758,N9762,N9763,N9764,N9765,
     N9766,N9767,N9768,N9769,N9773,N9774,N9775,N9779,N9784,N9785,
     N9786,N9790,N9791,N9795,N9796,N9797,N9798,N9799,N9800,N9801,
     N9802,N9803,N9805,N9806,N9809,N9813,N9814,N9815,N9816,N9817,
     N9820,N9825,N9826,N9827,N9828,N9829,N9830,N9835,N9836,N9837,
     N9838,N9846,N9847,N9862,N9863,N9866,N9873,N9876,N9890,N9891,
     N9892,N9893,N9894,N9895,N9896,N9897,N9898,N9899,N9900,N9901,
     N9902,N9903,N9904,N9905,N9906,N9907,N9908,N9909,N9910,N9911,
     N9917,N9923,N9924,N9925,N9932,N9935,N9938,N9939,N9945,N9946,
     N9947,N9948,N9949,N9953,N9954,N9955,N9956,N9957,N9958,N9959,
     N9960,N9961,N9964,N9967,N9968,N9969,N9970,N9971,N9972,N9973,
     N9974,N9975,N9976,N9977,N9978,N9979,N9982,N9983,N9986,N9989,
     N9992,N9995,N9996,N9997,N9998,N9999,N10002,N10003,N10006,N10007,
     N10010,N10013,N10014,N10015,N10016,N10017,N10018,N10019,N10020,N10021,
     N10022,N10023,N10024,N10026,N10028,N10032,N10033,N10034,N10035,N10036,
     N10037,N10038,N10039,N10040,N10041,N10042,N10043,N10050,N10053,N10054,
     N10055,N10056,N10057,N10058,N10059,N10060,N10061,N10062,N10067,N10070,
     N10073,N10076,N10077,N10082,N10083,N10084,N10085,N10086,N10093,N10094,
     N10105,N10106,N10107,N10108,N10113,N10114,N10115,N10116,N10119,N10124,
     N10130,N10131,N10132,N10133,N10134,N10135,N10136,N10137,N10138,N10139,
     N10140,N10141,N10148,N10155,N10156,N10157,N10158,N10159,N10160,N10161,
     N10162,N10163,N10164,N10165,N10170,N10173,N10176,N10177,N10178,N10179,
     N10180,N10183,N10186,N10189,N10192,N10195,N10196,N10197,N10200,N10203,
     N10204,N10205,N10206,N10212,N10213,N10230,N10231,N10232,N10233,N10234,
     N10237,N10238,N10239,N10240,N10241,N10242,N10247,N10248,N10259,N10264,
     N10265,N10266,N10267,N10268,N10269,N10270,N10271,N10272,N10273,N10278,
     N10279,N10280,N10281,N10282,N10283,N10287,N10288,N10289,N10290,N10291,
     N10292,N10293,N10294,N10295,N10296,N10299,N10300,N10301,N10306,N10307,
     N10308,N10311,N10314,N10315,N10316,N10317,N10318,N10321,N10324,N10325,
     N10326,N10327,N10328,N10329,N10330,N10331,N10332,N10333,N10334,N10337,
     N10338,N10339,N10340,N10341,N10344,N10354,N10357,N10360,N10367,N10375,
     N10381,N10388,N10391,N10399,N10402,N10406,N10409,N10412,N10415,N10419,
     N10422,N10425,N10428,N10431,N10432,N10437,N10438,N10439,N10440,N10441,
     N10444,N10445,N10450,N10451,N10455,N10456,N10465,N10466,N10479,N10497,
     N10509,N10512,N10515,N10516,N10517,N10518,N10519,N10522,N10525,N10528,
     N10531,N10534,N10535,N10536,N10539,N10542,N10543,N10544,N10545,N10546,
     N10547,N10548,N10549,N10550,N10551,N10552,N10553,N10554,N10555,N10556,
     N10557,N10558,N10559,N10560,N10561,N10562,N10563,N10564,N10565,N10566,
     N10567,N10568,N10569,N10570,N10571,N10572,N10573,N10577,N10581,N10582,
     N10583,N10587,N10588,N10589,N10594,N10595,N10596,N10597,N10598,N10602,
     N10609,N10610,N10621,N10626,N10627,N10629,N10631,N10637,N10638,N10639,
     N10640,N10642,N10643,N10644,N10645,N10647,N10648,N10649,N10652,N10659,
     N10662,N10665,N10668,N10671,N10672,N10673,N10674,N10675,N10678,N10681,
     N10682,N10683,N10684,N10685,N10686,N10687,N10688,N10689,N10690,N10691,
     N10694,N10695,N10696,N10697,N10698,N10701,N10705,N10707,N10708,N10709,
     N10710,N10719,N10720,N10730,N10731,N10737,N10738,N10739,N10746,N10747,
     N10748,N10749,N10750,N10753,N10754,N10764,N10765,N10766,N10767,N10768,
     N10769,N10770,N10771,N10772,N10773,N10774,N10775,N10776,N10778,N10781,
     N10784,N10789,N10792,N10796,N10797,N10798,N10799,N10800,N10803,N10806,
     N10809,N10812,N10815,N10816,N10817,N10820,N10823,N10824,N10825,N10826,
     N10832,N10833,N10834,N10835,N10836,N10845,N10846,N10857,N10862,N10863,
     N10864,N10865,N10866,N10867,N10872,N10873,N10874,N10875,N10876,N10879,
     N10882,N10883,N10884,N10885,N10886,N10887,N10888,N10889,N10890,N10891,
     N10892,N10895,N10896,N10897,N10898,N10899,N10902,N10909,N10910,N10915,
     N10916,N10917,N10918,N10919,N10922,N10923,N10928,N10931,N10934,N10935,
     N10936,N10937,N10938,N10941,N10944,N10947,N10950,N10953,N10954,N10955,
     N10958,N10961,N10962,N10963,N10964,N10969,N10970,N10981,N10986,N10987,
     N10988,N10989,N10990,N10991,N10992,N10995,N10998,N10999,N11000,N11001,
     N11002,N11003,N11004,N11005,N11006,N11007,N11008,N11011,N11012,N11013,
     N11014,N11015,N11018,N11023,N11024,N11027,N11028,N11029,N11030,N11031,
     N11034,N11035,N11040,N11041,N11042,N11043,N11044,N11047,N11050,N11053,
     N11056,N11059,N11062,N11065,N11066,N11067,N11070,N11073,N11074,N11075,
     N11076,N11077,N11078,N11095,N11098,N11099,N11100,N11103,N11106,N11107,
     N11108,N11109,N11110,N11111,N11112,N11113,N11114,N11115,N11116,N11117,
     N11118,N11119,N11120,N11121,N11122,N11123,N11124,N11127,N11130,N11137,
     N11138,N11139,N11140,N11141,N11142,N11143,N11144,N11145,N11152,N11153,
     N11154,N11155,N11156,N11159,N11162,N11165,N11168,N11171,N11174,N11177,
     N11180,N11183,N11184,N11185,N11186,N11187,N11188,N11205,N11210,N11211,
     N11212,N11213,N11214,N11215,N11216,N11217,N11218,N11219,N11220,N11222,
     N11223,N11224,N11225,N11226,N11227,N11228,N11229,N11231,N11232,N11233,
     N11236,N11239,N11242,N11243,N11244,N11245,N11246,N11250,N11252,N11257,
     N11260,N11261,N11262,N11263,N11264,N11265,N11267,N11268,N11269,N11270,
     N11272,N11277,N11278,N11279,N11280,N11282,N11283,N11284,N11285,N11286,
     N11288,N11289,N11290,N11291,N11292,N11293,N11294,N11295,N11296,N11297,
     N11298,N11299,N11302,N11307,N11308,N11309,N11312,N11313,N11314,N11315,
     N11316,N11317,N11320,N11321,N11323,N11327,N11328,N11329,N11331,N11335,
     N11336,N11337,N11338,N11339,N11341, gate3184inter0, gate3184inter1, gate3184inter2, gate3184inter3, gate3184inter4, gate3184inter5, gate3184inter6, gate3184inter7, gate3184inter8, gate3184inter9, gate3184inter10, gate3184inter11, gate3184inter12, gate3154inter0, gate3154inter1, gate3154inter2, gate3154inter3, gate3154inter4, gate3154inter5, gate3154inter6, gate3154inter7, gate3154inter8, gate3154inter9, gate3154inter10, gate3154inter11, gate3154inter12, gate2263inter0, gate2263inter1, gate2263inter2, gate2263inter3, gate2263inter4, gate2263inter5, gate2263inter6, gate2263inter7, gate2263inter8, gate2263inter9, gate2263inter10, gate2263inter11, gate2263inter12, gate484inter0, gate484inter1, gate484inter2, gate484inter3, gate484inter4, gate484inter5, gate484inter6, gate484inter7, gate484inter8, gate484inter9, gate484inter10, gate484inter11, gate484inter12, gate1495inter0, gate1495inter1, gate1495inter2, gate1495inter3, gate1495inter4, gate1495inter5, gate1495inter6, gate1495inter7, gate1495inter8, gate1495inter9, gate1495inter10, gate1495inter11, gate1495inter12, gate1669inter0, gate1669inter1, gate1669inter2, gate1669inter3, gate1669inter4, gate1669inter5, gate1669inter6, gate1669inter7, gate1669inter8, gate1669inter9, gate1669inter10, gate1669inter11, gate1669inter12, gate1421inter0, gate1421inter1, gate1421inter2, gate1421inter3, gate1421inter4, gate1421inter5, gate1421inter6, gate1421inter7, gate1421inter8, gate1421inter9, gate1421inter10, gate1421inter11, gate1421inter12, gate3413inter0, gate3413inter1, gate3413inter2, gate3413inter3, gate3413inter4, gate3413inter5, gate3413inter6, gate3413inter7, gate3413inter8, gate3413inter9, gate3413inter10, gate3413inter11, gate3413inter12, gate3082inter0, gate3082inter1, gate3082inter2, gate3082inter3, gate3082inter4, gate3082inter5, gate3082inter6, gate3082inter7, gate3082inter8, gate3082inter9, gate3082inter10, gate3082inter11, gate3082inter12, gate1405inter0, gate1405inter1, gate1405inter2, gate1405inter3, gate1405inter4, gate1405inter5, gate1405inter6, gate1405inter7, gate1405inter8, gate1405inter9, gate1405inter10, gate1405inter11, gate1405inter12, gate2459inter0, gate2459inter1, gate2459inter2, gate2459inter3, gate2459inter4, gate2459inter5, gate2459inter6, gate2459inter7, gate2459inter8, gate2459inter9, gate2459inter10, gate2459inter11, gate2459inter12, gate2885inter0, gate2885inter1, gate2885inter2, gate2885inter3, gate2885inter4, gate2885inter5, gate2885inter6, gate2885inter7, gate2885inter8, gate2885inter9, gate2885inter10, gate2885inter11, gate2885inter12, gate958inter0, gate958inter1, gate958inter2, gate958inter3, gate958inter4, gate958inter5, gate958inter6, gate958inter7, gate958inter8, gate958inter9, gate958inter10, gate958inter11, gate958inter12, gate1687inter0, gate1687inter1, gate1687inter2, gate1687inter3, gate1687inter4, gate1687inter5, gate1687inter6, gate1687inter7, gate1687inter8, gate1687inter9, gate1687inter10, gate1687inter11, gate1687inter12, gate3175inter0, gate3175inter1, gate3175inter2, gate3175inter3, gate3175inter4, gate3175inter5, gate3175inter6, gate3175inter7, gate3175inter8, gate3175inter9, gate3175inter10, gate3175inter11, gate3175inter12, gate2920inter0, gate2920inter1, gate2920inter2, gate2920inter3, gate2920inter4, gate2920inter5, gate2920inter6, gate2920inter7, gate2920inter8, gate2920inter9, gate2920inter10, gate2920inter11, gate2920inter12, gate835inter0, gate835inter1, gate835inter2, gate835inter3, gate835inter4, gate835inter5, gate835inter6, gate835inter7, gate835inter8, gate835inter9, gate835inter10, gate835inter11, gate835inter12, gate2571inter0, gate2571inter1, gate2571inter2, gate2571inter3, gate2571inter4, gate2571inter5, gate2571inter6, gate2571inter7, gate2571inter8, gate2571inter9, gate2571inter10, gate2571inter11, gate2571inter12, gate784inter0, gate784inter1, gate784inter2, gate784inter3, gate784inter4, gate784inter5, gate784inter6, gate784inter7, gate784inter8, gate784inter9, gate784inter10, gate784inter11, gate784inter12, gate3003inter0, gate3003inter1, gate3003inter2, gate3003inter3, gate3003inter4, gate3003inter5, gate3003inter6, gate3003inter7, gate3003inter8, gate3003inter9, gate3003inter10, gate3003inter11, gate3003inter12, gate2976inter0, gate2976inter1, gate2976inter2, gate2976inter3, gate2976inter4, gate2976inter5, gate2976inter6, gate2976inter7, gate2976inter8, gate2976inter9, gate2976inter10, gate2976inter11, gate2976inter12, gate3377inter0, gate3377inter1, gate3377inter2, gate3377inter3, gate3377inter4, gate3377inter5, gate3377inter6, gate3377inter7, gate3377inter8, gate3377inter9, gate3377inter10, gate3377inter11, gate3377inter12, gate2870inter0, gate2870inter1, gate2870inter2, gate2870inter3, gate2870inter4, gate2870inter5, gate2870inter6, gate2870inter7, gate2870inter8, gate2870inter9, gate2870inter10, gate2870inter11, gate2870inter12, gate1003inter0, gate1003inter1, gate1003inter2, gate1003inter3, gate1003inter4, gate1003inter5, gate1003inter6, gate1003inter7, gate1003inter8, gate1003inter9, gate1003inter10, gate1003inter11, gate1003inter12, gate1379inter0, gate1379inter1, gate1379inter2, gate1379inter3, gate1379inter4, gate1379inter5, gate1379inter6, gate1379inter7, gate1379inter8, gate1379inter9, gate1379inter10, gate1379inter11, gate1379inter12, gate2653inter0, gate2653inter1, gate2653inter2, gate2653inter3, gate2653inter4, gate2653inter5, gate2653inter6, gate2653inter7, gate2653inter8, gate2653inter9, gate2653inter10, gate2653inter11, gate2653inter12, gate1329inter0, gate1329inter1, gate1329inter2, gate1329inter3, gate1329inter4, gate1329inter5, gate1329inter6, gate1329inter7, gate1329inter8, gate1329inter9, gate1329inter10, gate1329inter11, gate1329inter12, gate3497inter0, gate3497inter1, gate3497inter2, gate3497inter3, gate3497inter4, gate3497inter5, gate3497inter6, gate3497inter7, gate3497inter8, gate3497inter9, gate3497inter10, gate3497inter11, gate3497inter12, gate3464inter0, gate3464inter1, gate3464inter2, gate3464inter3, gate3464inter4, gate3464inter5, gate3464inter6, gate3464inter7, gate3464inter8, gate3464inter9, gate3464inter10, gate3464inter11, gate3464inter12, gate2747inter0, gate2747inter1, gate2747inter2, gate2747inter3, gate2747inter4, gate2747inter5, gate2747inter6, gate2747inter7, gate2747inter8, gate2747inter9, gate2747inter10, gate2747inter11, gate2747inter12, gate3243inter0, gate3243inter1, gate3243inter2, gate3243inter3, gate3243inter4, gate3243inter5, gate3243inter6, gate3243inter7, gate3243inter8, gate3243inter9, gate3243inter10, gate3243inter11, gate3243inter12, gate1610inter0, gate1610inter1, gate1610inter2, gate1610inter3, gate1610inter4, gate1610inter5, gate1610inter6, gate1610inter7, gate1610inter8, gate1610inter9, gate1610inter10, gate1610inter11, gate1610inter12, gate1412inter0, gate1412inter1, gate1412inter2, gate1412inter3, gate1412inter4, gate1412inter5, gate1412inter6, gate1412inter7, gate1412inter8, gate1412inter9, gate1412inter10, gate1412inter11, gate1412inter12, gate3147inter0, gate3147inter1, gate3147inter2, gate3147inter3, gate3147inter4, gate3147inter5, gate3147inter6, gate3147inter7, gate3147inter8, gate3147inter9, gate3147inter10, gate3147inter11, gate3147inter12, gate3336inter0, gate3336inter1, gate3336inter2, gate3336inter3, gate3336inter4, gate3336inter5, gate3336inter6, gate3336inter7, gate3336inter8, gate3336inter9, gate3336inter10, gate3336inter11, gate3336inter12, gate1861inter0, gate1861inter1, gate1861inter2, gate1861inter3, gate1861inter4, gate1861inter5, gate1861inter6, gate1861inter7, gate1861inter8, gate1861inter9, gate1861inter10, gate1861inter11, gate1861inter12, gate1744inter0, gate1744inter1, gate1744inter2, gate1744inter3, gate1744inter4, gate1744inter5, gate1744inter6, gate1744inter7, gate1744inter8, gate1744inter9, gate1744inter10, gate1744inter11, gate1744inter12, gate3145inter0, gate3145inter1, gate3145inter2, gate3145inter3, gate3145inter4, gate3145inter5, gate3145inter6, gate3145inter7, gate3145inter8, gate3145inter9, gate3145inter10, gate3145inter11, gate3145inter12, gate2572inter0, gate2572inter1, gate2572inter2, gate2572inter3, gate2572inter4, gate2572inter5, gate2572inter6, gate2572inter7, gate2572inter8, gate2572inter9, gate2572inter10, gate2572inter11, gate2572inter12, gate1557inter0, gate1557inter1, gate1557inter2, gate1557inter3, gate1557inter4, gate1557inter5, gate1557inter6, gate1557inter7, gate1557inter8, gate1557inter9, gate1557inter10, gate1557inter11, gate1557inter12, gate1846inter0, gate1846inter1, gate1846inter2, gate1846inter3, gate1846inter4, gate1846inter5, gate1846inter6, gate1846inter7, gate1846inter8, gate1846inter9, gate1846inter10, gate1846inter11, gate1846inter12, gate2757inter0, gate2757inter1, gate2757inter2, gate2757inter3, gate2757inter4, gate2757inter5, gate2757inter6, gate2757inter7, gate2757inter8, gate2757inter9, gate2757inter10, gate2757inter11, gate2757inter12, gate917inter0, gate917inter1, gate917inter2, gate917inter3, gate917inter4, gate917inter5, gate917inter6, gate917inter7, gate917inter8, gate917inter9, gate917inter10, gate917inter11, gate917inter12, gate1312inter0, gate1312inter1, gate1312inter2, gate1312inter3, gate1312inter4, gate1312inter5, gate1312inter6, gate1312inter7, gate1312inter8, gate1312inter9, gate1312inter10, gate1312inter11, gate1312inter12, gate1510inter0, gate1510inter1, gate1510inter2, gate1510inter3, gate1510inter4, gate1510inter5, gate1510inter6, gate1510inter7, gate1510inter8, gate1510inter9, gate1510inter10, gate1510inter11, gate1510inter12, gate1672inter0, gate1672inter1, gate1672inter2, gate1672inter3, gate1672inter4, gate1672inter5, gate1672inter6, gate1672inter7, gate1672inter8, gate1672inter9, gate1672inter10, gate1672inter11, gate1672inter12, gate3244inter0, gate3244inter1, gate3244inter2, gate3244inter3, gate3244inter4, gate3244inter5, gate3244inter6, gate3244inter7, gate3244inter8, gate3244inter9, gate3244inter10, gate3244inter11, gate3244inter12, gate1730inter0, gate1730inter1, gate1730inter2, gate1730inter3, gate1730inter4, gate1730inter5, gate1730inter6, gate1730inter7, gate1730inter8, gate1730inter9, gate1730inter10, gate1730inter11, gate1730inter12, gate1367inter0, gate1367inter1, gate1367inter2, gate1367inter3, gate1367inter4, gate1367inter5, gate1367inter6, gate1367inter7, gate1367inter8, gate1367inter9, gate1367inter10, gate1367inter11, gate1367inter12, gate3455inter0, gate3455inter1, gate3455inter2, gate3455inter3, gate3455inter4, gate3455inter5, gate3455inter6, gate3455inter7, gate3455inter8, gate3455inter9, gate3455inter10, gate3455inter11, gate3455inter12, gate2696inter0, gate2696inter1, gate2696inter2, gate2696inter3, gate2696inter4, gate2696inter5, gate2696inter6, gate2696inter7, gate2696inter8, gate2696inter9, gate2696inter10, gate2696inter11, gate2696inter12, gate1913inter0, gate1913inter1, gate1913inter2, gate1913inter3, gate1913inter4, gate1913inter5, gate1913inter6, gate1913inter7, gate1913inter8, gate1913inter9, gate1913inter10, gate1913inter11, gate1913inter12, gate1362inter0, gate1362inter1, gate1362inter2, gate1362inter3, gate1362inter4, gate1362inter5, gate1362inter6, gate1362inter7, gate1362inter8, gate1362inter9, gate1362inter10, gate1362inter11, gate1362inter12, gate2946inter0, gate2946inter1, gate2946inter2, gate2946inter3, gate2946inter4, gate2946inter5, gate2946inter6, gate2946inter7, gate2946inter8, gate2946inter9, gate2946inter10, gate2946inter11, gate2946inter12, gate2047inter0, gate2047inter1, gate2047inter2, gate2047inter3, gate2047inter4, gate2047inter5, gate2047inter6, gate2047inter7, gate2047inter8, gate2047inter9, gate2047inter10, gate2047inter11, gate2047inter12, gate1643inter0, gate1643inter1, gate1643inter2, gate1643inter3, gate1643inter4, gate1643inter5, gate1643inter6, gate1643inter7, gate1643inter8, gate1643inter9, gate1643inter10, gate1643inter11, gate1643inter12, gate2715inter0, gate2715inter1, gate2715inter2, gate2715inter3, gate2715inter4, gate2715inter5, gate2715inter6, gate2715inter7, gate2715inter8, gate2715inter9, gate2715inter10, gate2715inter11, gate2715inter12, gate2661inter0, gate2661inter1, gate2661inter2, gate2661inter3, gate2661inter4, gate2661inter5, gate2661inter6, gate2661inter7, gate2661inter8, gate2661inter9, gate2661inter10, gate2661inter11, gate2661inter12, gate1147inter0, gate1147inter1, gate1147inter2, gate1147inter3, gate1147inter4, gate1147inter5, gate1147inter6, gate1147inter7, gate1147inter8, gate1147inter9, gate1147inter10, gate1147inter11, gate1147inter12, gate3054inter0, gate3054inter1, gate3054inter2, gate3054inter3, gate3054inter4, gate3054inter5, gate3054inter6, gate3054inter7, gate3054inter8, gate3054inter9, gate3054inter10, gate3054inter11, gate3054inter12, gate2620inter0, gate2620inter1, gate2620inter2, gate2620inter3, gate2620inter4, gate2620inter5, gate2620inter6, gate2620inter7, gate2620inter8, gate2620inter9, gate2620inter10, gate2620inter11, gate2620inter12, gate1652inter0, gate1652inter1, gate1652inter2, gate1652inter3, gate1652inter4, gate1652inter5, gate1652inter6, gate1652inter7, gate1652inter8, gate1652inter9, gate1652inter10, gate1652inter11, gate1652inter12, gate1890inter0, gate1890inter1, gate1890inter2, gate1890inter3, gate1890inter4, gate1890inter5, gate1890inter6, gate1890inter7, gate1890inter8, gate1890inter9, gate1890inter10, gate1890inter11, gate1890inter12, gate3367inter0, gate3367inter1, gate3367inter2, gate3367inter3, gate3367inter4, gate3367inter5, gate3367inter6, gate3367inter7, gate3367inter8, gate3367inter9, gate3367inter10, gate3367inter11, gate3367inter12, gate1740inter0, gate1740inter1, gate1740inter2, gate1740inter3, gate1740inter4, gate1740inter5, gate1740inter6, gate1740inter7, gate1740inter8, gate1740inter9, gate1740inter10, gate1740inter11, gate1740inter12, gate1674inter0, gate1674inter1, gate1674inter2, gate1674inter3, gate1674inter4, gate1674inter5, gate1674inter6, gate1674inter7, gate1674inter8, gate1674inter9, gate1674inter10, gate1674inter11, gate1674inter12, gate3461inter0, gate3461inter1, gate3461inter2, gate3461inter3, gate3461inter4, gate3461inter5, gate3461inter6, gate3461inter7, gate3461inter8, gate3461inter9, gate3461inter10, gate3461inter11, gate3461inter12, gate3186inter0, gate3186inter1, gate3186inter2, gate3186inter3, gate3186inter4, gate3186inter5, gate3186inter6, gate3186inter7, gate3186inter8, gate3186inter9, gate3186inter10, gate3186inter11, gate3186inter12, gate2947inter0, gate2947inter1, gate2947inter2, gate2947inter3, gate2947inter4, gate2947inter5, gate2947inter6, gate2947inter7, gate2947inter8, gate2947inter9, gate2947inter10, gate2947inter11, gate2947inter12, gate1690inter0, gate1690inter1, gate1690inter2, gate1690inter3, gate1690inter4, gate1690inter5, gate1690inter6, gate1690inter7, gate1690inter8, gate1690inter9, gate1690inter10, gate1690inter11, gate1690inter12, gate3381inter0, gate3381inter1, gate3381inter2, gate3381inter3, gate3381inter4, gate3381inter5, gate3381inter6, gate3381inter7, gate3381inter8, gate3381inter9, gate3381inter10, gate3381inter11, gate3381inter12, gate1930inter0, gate1930inter1, gate1930inter2, gate1930inter3, gate1930inter4, gate1930inter5, gate1930inter6, gate1930inter7, gate1930inter8, gate1930inter9, gate1930inter10, gate1930inter11, gate1930inter12, gate2891inter0, gate2891inter1, gate2891inter2, gate2891inter3, gate2891inter4, gate2891inter5, gate2891inter6, gate2891inter7, gate2891inter8, gate2891inter9, gate2891inter10, gate2891inter11, gate2891inter12, gate1537inter0, gate1537inter1, gate1537inter2, gate1537inter3, gate1537inter4, gate1537inter5, gate1537inter6, gate1537inter7, gate1537inter8, gate1537inter9, gate1537inter10, gate1537inter11, gate1537inter12, gate2802inter0, gate2802inter1, gate2802inter2, gate2802inter3, gate2802inter4, gate2802inter5, gate2802inter6, gate2802inter7, gate2802inter8, gate2802inter9, gate2802inter10, gate2802inter11, gate2802inter12, gate1359inter0, gate1359inter1, gate1359inter2, gate1359inter3, gate1359inter4, gate1359inter5, gate1359inter6, gate1359inter7, gate1359inter8, gate1359inter9, gate1359inter10, gate1359inter11, gate1359inter12, gate1535inter0, gate1535inter1, gate1535inter2, gate1535inter3, gate1535inter4, gate1535inter5, gate1535inter6, gate1535inter7, gate1535inter8, gate1535inter9, gate1535inter10, gate1535inter11, gate1535inter12, gate3050inter0, gate3050inter1, gate3050inter2, gate3050inter3, gate3050inter4, gate3050inter5, gate3050inter6, gate3050inter7, gate3050inter8, gate3050inter9, gate3050inter10, gate3050inter11, gate3050inter12, gate1356inter0, gate1356inter1, gate1356inter2, gate1356inter3, gate1356inter4, gate1356inter5, gate1356inter6, gate1356inter7, gate1356inter8, gate1356inter9, gate1356inter10, gate1356inter11, gate1356inter12, gate1555inter0, gate1555inter1, gate1555inter2, gate1555inter3, gate1555inter4, gate1555inter5, gate1555inter6, gate1555inter7, gate1555inter8, gate1555inter9, gate1555inter10, gate1555inter11, gate1555inter12, gate2312inter0, gate2312inter1, gate2312inter2, gate2312inter3, gate2312inter4, gate2312inter5, gate2312inter6, gate2312inter7, gate2312inter8, gate2312inter9, gate2312inter10, gate2312inter11, gate2312inter12, gate2796inter0, gate2796inter1, gate2796inter2, gate2796inter3, gate2796inter4, gate2796inter5, gate2796inter6, gate2796inter7, gate2796inter8, gate2796inter9, gate2796inter10, gate2796inter11, gate2796inter12, gate1649inter0, gate1649inter1, gate1649inter2, gate1649inter3, gate1649inter4, gate1649inter5, gate1649inter6, gate1649inter7, gate1649inter8, gate1649inter9, gate1649inter10, gate1649inter11, gate1649inter12, gate1397inter0, gate1397inter1, gate1397inter2, gate1397inter3, gate1397inter4, gate1397inter5, gate1397inter6, gate1397inter7, gate1397inter8, gate1397inter9, gate1397inter10, gate1397inter11, gate1397inter12, gate1347inter0, gate1347inter1, gate1347inter2, gate1347inter3, gate1347inter4, gate1347inter5, gate1347inter6, gate1347inter7, gate1347inter8, gate1347inter9, gate1347inter10, gate1347inter11, gate1347inter12, gate1478inter0, gate1478inter1, gate1478inter2, gate1478inter3, gate1478inter4, gate1478inter5, gate1478inter6, gate1478inter7, gate1478inter8, gate1478inter9, gate1478inter10, gate1478inter11, gate1478inter12, gate1920inter0, gate1920inter1, gate1920inter2, gate1920inter3, gate1920inter4, gate1920inter5, gate1920inter6, gate1920inter7, gate1920inter8, gate1920inter9, gate1920inter10, gate1920inter11, gate1920inter12, gate3329inter0, gate3329inter1, gate3329inter2, gate3329inter3, gate3329inter4, gate3329inter5, gate3329inter6, gate3329inter7, gate3329inter8, gate3329inter9, gate3329inter10, gate3329inter11, gate3329inter12, gate1102inter0, gate1102inter1, gate1102inter2, gate1102inter3, gate1102inter4, gate1102inter5, gate1102inter6, gate1102inter7, gate1102inter8, gate1102inter9, gate1102inter10, gate1102inter11, gate1102inter12, gate2050inter0, gate2050inter1, gate2050inter2, gate2050inter3, gate2050inter4, gate2050inter5, gate2050inter6, gate2050inter7, gate2050inter8, gate2050inter9, gate2050inter10, gate2050inter11, gate2050inter12, gate3204inter0, gate3204inter1, gate3204inter2, gate3204inter3, gate3204inter4, gate3204inter5, gate3204inter6, gate3204inter7, gate3204inter8, gate3204inter9, gate3204inter10, gate3204inter11, gate3204inter12, gate1655inter0, gate1655inter1, gate1655inter2, gate1655inter3, gate1655inter4, gate1655inter5, gate1655inter6, gate1655inter7, gate1655inter8, gate1655inter9, gate1655inter10, gate1655inter11, gate1655inter12, gate3217inter0, gate3217inter1, gate3217inter2, gate3217inter3, gate3217inter4, gate3217inter5, gate3217inter6, gate3217inter7, gate3217inter8, gate3217inter9, gate3217inter10, gate3217inter11, gate3217inter12, gate579inter0, gate579inter1, gate579inter2, gate579inter3, gate579inter4, gate579inter5, gate579inter6, gate579inter7, gate579inter8, gate579inter9, gate579inter10, gate579inter11, gate579inter12, gate1630inter0, gate1630inter1, gate1630inter2, gate1630inter3, gate1630inter4, gate1630inter5, gate1630inter6, gate1630inter7, gate1630inter8, gate1630inter9, gate1630inter10, gate1630inter11, gate1630inter12, gate2426inter0, gate2426inter1, gate2426inter2, gate2426inter3, gate2426inter4, gate2426inter5, gate2426inter6, gate2426inter7, gate2426inter8, gate2426inter9, gate2426inter10, gate2426inter11, gate2426inter12, gate3038inter0, gate3038inter1, gate3038inter2, gate3038inter3, gate3038inter4, gate3038inter5, gate3038inter6, gate3038inter7, gate3038inter8, gate3038inter9, gate3038inter10, gate3038inter11, gate3038inter12, gate1364inter0, gate1364inter1, gate1364inter2, gate1364inter3, gate1364inter4, gate1364inter5, gate1364inter6, gate1364inter7, gate1364inter8, gate1364inter9, gate1364inter10, gate1364inter11, gate1364inter12, gate2932inter0, gate2932inter1, gate2932inter2, gate2932inter3, gate2932inter4, gate2932inter5, gate2932inter6, gate2932inter7, gate2932inter8, gate2932inter9, gate2932inter10, gate2932inter11, gate2932inter12, gate2656inter0, gate2656inter1, gate2656inter2, gate2656inter3, gate2656inter4, gate2656inter5, gate2656inter6, gate2656inter7, gate2656inter8, gate2656inter9, gate2656inter10, gate2656inter11, gate2656inter12, gate1879inter0, gate1879inter1, gate1879inter2, gate1879inter3, gate1879inter4, gate1879inter5, gate1879inter6, gate1879inter7, gate1879inter8, gate1879inter9, gate1879inter10, gate1879inter11, gate1879inter12, gate1391inter0, gate1391inter1, gate1391inter2, gate1391inter3, gate1391inter4, gate1391inter5, gate1391inter6, gate1391inter7, gate1391inter8, gate1391inter9, gate1391inter10, gate1391inter11, gate1391inter12, gate3046inter0, gate3046inter1, gate3046inter2, gate3046inter3, gate3046inter4, gate3046inter5, gate3046inter6, gate3046inter7, gate3046inter8, gate3046inter9, gate3046inter10, gate3046inter11, gate3046inter12, gate1466inter0, gate1466inter1, gate1466inter2, gate1466inter3, gate1466inter4, gate1466inter5, gate1466inter6, gate1466inter7, gate1466inter8, gate1466inter9, gate1466inter10, gate1466inter11, gate1466inter12, gate3122inter0, gate3122inter1, gate3122inter2, gate3122inter3, gate3122inter4, gate3122inter5, gate3122inter6, gate3122inter7, gate3122inter8, gate3122inter9, gate3122inter10, gate3122inter11, gate3122inter12, gate3304inter0, gate3304inter1, gate3304inter2, gate3304inter3, gate3304inter4, gate3304inter5, gate3304inter6, gate3304inter7, gate3304inter8, gate3304inter9, gate3304inter10, gate3304inter11, gate3304inter12, gate2411inter0, gate2411inter1, gate2411inter2, gate2411inter3, gate2411inter4, gate2411inter5, gate2411inter6, gate2411inter7, gate2411inter8, gate2411inter9, gate2411inter10, gate2411inter11, gate2411inter12, gate1371inter0, gate1371inter1, gate1371inter2, gate1371inter3, gate1371inter4, gate1371inter5, gate1371inter6, gate1371inter7, gate1371inter8, gate1371inter9, gate1371inter10, gate1371inter11, gate1371inter12, gate1289inter0, gate1289inter1, gate1289inter2, gate1289inter3, gate1289inter4, gate1289inter5, gate1289inter6, gate1289inter7, gate1289inter8, gate1289inter9, gate1289inter10, gate1289inter11, gate1289inter12, gate3296inter0, gate3296inter1, gate3296inter2, gate3296inter3, gate3296inter4, gate3296inter5, gate3296inter6, gate3296inter7, gate3296inter8, gate3296inter9, gate3296inter10, gate3296inter11, gate3296inter12, gate1330inter0, gate1330inter1, gate1330inter2, gate1330inter3, gate1330inter4, gate1330inter5, gate1330inter6, gate1330inter7, gate1330inter8, gate1330inter9, gate1330inter10, gate1330inter11, gate1330inter12, gate1859inter0, gate1859inter1, gate1859inter2, gate1859inter3, gate1859inter4, gate1859inter5, gate1859inter6, gate1859inter7, gate1859inter8, gate1859inter9, gate1859inter10, gate1859inter11, gate1859inter12, gate1328inter0, gate1328inter1, gate1328inter2, gate1328inter3, gate1328inter4, gate1328inter5, gate1328inter6, gate1328inter7, gate1328inter8, gate1328inter9, gate1328inter10, gate1328inter11, gate1328inter12, gate1727inter0, gate1727inter1, gate1727inter2, gate1727inter3, gate1727inter4, gate1727inter5, gate1727inter6, gate1727inter7, gate1727inter8, gate1727inter9, gate1727inter10, gate1727inter11, gate1727inter12, gate3084inter0, gate3084inter1, gate3084inter2, gate3084inter3, gate3084inter4, gate3084inter5, gate3084inter6, gate3084inter7, gate3084inter8, gate3084inter9, gate3084inter10, gate3084inter11, gate3084inter12, gate3215inter0, gate3215inter1, gate3215inter2, gate3215inter3, gate3215inter4, gate3215inter5, gate3215inter6, gate3215inter7, gate3215inter8, gate3215inter9, gate3215inter10, gate3215inter11, gate3215inter12, gate935inter0, gate935inter1, gate935inter2, gate935inter3, gate935inter4, gate935inter5, gate935inter6, gate935inter7, gate935inter8, gate935inter9, gate935inter10, gate935inter11, gate935inter12, gate1286inter0, gate1286inter1, gate1286inter2, gate1286inter3, gate1286inter4, gate1286inter5, gate1286inter6, gate1286inter7, gate1286inter8, gate1286inter9, gate1286inter10, gate1286inter11, gate1286inter12, gate3212inter0, gate3212inter1, gate3212inter2, gate3212inter3, gate3212inter4, gate3212inter5, gate3212inter6, gate3212inter7, gate3212inter8, gate3212inter9, gate3212inter10, gate3212inter11, gate3212inter12, gate3500inter0, gate3500inter1, gate3500inter2, gate3500inter3, gate3500inter4, gate3500inter5, gate3500inter6, gate3500inter7, gate3500inter8, gate3500inter9, gate3500inter10, gate3500inter11, gate3500inter12, gate3120inter0, gate3120inter1, gate3120inter2, gate3120inter3, gate3120inter4, gate3120inter5, gate3120inter6, gate3120inter7, gate3120inter8, gate3120inter9, gate3120inter10, gate3120inter11, gate3120inter12, gate1558inter0, gate1558inter1, gate1558inter2, gate1558inter3, gate1558inter4, gate1558inter5, gate1558inter6, gate1558inter7, gate1558inter8, gate1558inter9, gate1558inter10, gate1558inter11, gate1558inter12, gate3298inter0, gate3298inter1, gate3298inter2, gate3298inter3, gate3298inter4, gate3298inter5, gate3298inter6, gate3298inter7, gate3298inter8, gate3298inter9, gate3298inter10, gate3298inter11, gate3298inter12, gate2823inter0, gate2823inter1, gate2823inter2, gate2823inter3, gate2823inter4, gate2823inter5, gate2823inter6, gate2823inter7, gate2823inter8, gate2823inter9, gate2823inter10, gate2823inter11, gate2823inter12, gate3396inter0, gate3396inter1, gate3396inter2, gate3396inter3, gate3396inter4, gate3396inter5, gate3396inter6, gate3396inter7, gate3396inter8, gate3396inter9, gate3396inter10, gate3396inter11, gate3396inter12, gate1726inter0, gate1726inter1, gate1726inter2, gate1726inter3, gate1726inter4, gate1726inter5, gate1726inter6, gate1726inter7, gate1726inter8, gate1726inter9, gate1726inter10, gate1726inter11, gate1726inter12, gate121inter0, gate121inter1, gate121inter2, gate121inter3, gate121inter4, gate121inter5, gate121inter6, gate121inter7, gate121inter8, gate121inter9, gate121inter10, gate121inter11, gate121inter12, gate1314inter0, gate1314inter1, gate1314inter2, gate1314inter3, gate1314inter4, gate1314inter5, gate1314inter6, gate1314inter7, gate1314inter8, gate1314inter9, gate1314inter10, gate1314inter11, gate1314inter12, gate2443inter0, gate2443inter1, gate2443inter2, gate2443inter3, gate2443inter4, gate2443inter5, gate2443inter6, gate2443inter7, gate2443inter8, gate2443inter9, gate2443inter10, gate2443inter11, gate2443inter12, gate1474inter0, gate1474inter1, gate1474inter2, gate1474inter3, gate1474inter4, gate1474inter5, gate1474inter6, gate1474inter7, gate1474inter8, gate1474inter9, gate1474inter10, gate1474inter11, gate1474inter12, gate2797inter0, gate2797inter1, gate2797inter2, gate2797inter3, gate2797inter4, gate2797inter5, gate2797inter6, gate2797inter7, gate2797inter8, gate2797inter9, gate2797inter10, gate2797inter11, gate2797inter12;



buf1 gate1( .a(N1), .O(N387) );
buf1 gate2( .a(N1), .O(N388) );
inv1 gate3( .a(N57), .O(N467) );
and2 gate4( .a(N134), .b(N133), .O(N469) );
buf1 gate5( .a(N248), .O(N478) );
buf1 gate6( .a(N254), .O(N482) );
buf1 gate7( .a(N257), .O(N484) );
buf1 gate8( .a(N260), .O(N486) );
buf1 gate9( .a(N263), .O(N489) );
buf1 gate10( .a(N267), .O(N492) );
and4 gate11( .a(N162), .b(N172), .c(N188), .d(N199), .O(N494) );
buf1 gate12( .a(N274), .O(N501) );
buf1 gate13( .a(N280), .O(N505) );
buf1 gate14( .a(N283), .O(N507) );
buf1 gate15( .a(N286), .O(N509) );
buf1 gate16( .a(N289), .O(N511) );
buf1 gate17( .a(N293), .O(N513) );
buf1 gate18( .a(N296), .O(N515) );
buf1 gate19( .a(N299), .O(N517) );
buf1 gate20( .a(N303), .O(N519) );
and4 gate21( .a(N150), .b(N184), .c(N228), .d(N240), .O(N528) );
buf1 gate22( .a(N307), .O(N535) );
buf1 gate23( .a(N310), .O(N537) );
buf1 gate24( .a(N313), .O(N539) );
buf1 gate25( .a(N316), .O(N541) );
buf1 gate26( .a(N319), .O(N543) );
buf1 gate27( .a(N322), .O(N545) );
buf1 gate28( .a(N325), .O(N547) );
buf1 gate29( .a(N328), .O(N549) );
buf1 gate30( .a(N331), .O(N551) );
buf1 gate31( .a(N334), .O(N553) );
buf1 gate32( .a(N337), .O(N556) );
buf1 gate33( .a(N343), .O(N559) );
buf1 gate34( .a(N346), .O(N561) );
buf1 gate35( .a(N349), .O(N563) );
buf1 gate36( .a(N352), .O(N565) );
buf1 gate37( .a(N355), .O(N567) );
buf1 gate38( .a(N358), .O(N569) );
buf1 gate39( .a(N361), .O(N571) );
buf1 gate40( .a(N364), .O(N573) );
and4 gate41( .a(N183), .b(N182), .c(N185), .d(N186), .O(N575) );
and4 gate42( .a(N210), .b(N152), .c(N218), .d(N230), .O(N578) );
inv1 gate43( .a(N15), .O(N582) );
inv1 gate44( .a(N5), .O(N585) );
buf1 gate45( .a(N1), .O(N590) );
inv1 gate46( .a(N5), .O(N593) );
inv1 gate47( .a(N5), .O(N596) );
inv1 gate48( .a(N289), .O(N599) );
inv1 gate49( .a(N299), .O(N604) );
inv1 gate50( .a(N303), .O(N609) );
buf1 gate51( .a(N38), .O(N614) );
buf1 gate52( .a(N15), .O(N625) );
nand2 gate53( .a(N12), .b(N9), .O(N628) );
nand2 gate54( .a(N12), .b(N9), .O(N632) );
buf1 gate55( .a(N38), .O(N636) );
inv1 gate56( .a(N245), .O(N641) );
inv1 gate57( .a(N248), .O(N642) );
buf1 gate58( .a(N251), .O(N643) );
inv1 gate59( .a(N251), .O(N644) );
inv1 gate60( .a(N254), .O(N651) );
buf1 gate61( .a(N106), .O(N657) );
inv1 gate62( .a(N257), .O(N660) );
inv1 gate63( .a(N260), .O(N666) );
inv1 gate64( .a(N263), .O(N672) );
inv1 gate65( .a(N267), .O(N673) );
inv1 gate66( .a(N106), .O(N674) );
buf1 gate67( .a(N18), .O(N676) );
buf1 gate68( .a(N18), .O(N682) );
and2 gate69( .a(N382), .b(N263), .O(N688) );
buf1 gate70( .a(N18), .O(N689) );
inv1 gate71( .a(N18), .O(N695) );
nand2 gate72( .a(N382), .b(N267), .O(N700) );
inv1 gate73( .a(N271), .O(N705) );
inv1 gate74( .a(N274), .O(N706) );
buf1 gate75( .a(N277), .O(N707) );
inv1 gate76( .a(N277), .O(N708) );
inv1 gate77( .a(N280), .O(N715) );
inv1 gate78( .a(N283), .O(N721) );
inv1 gate79( .a(N286), .O(N727) );
inv1 gate80( .a(N289), .O(N733) );
inv1 gate81( .a(N293), .O(N734) );
inv1 gate82( .a(N296), .O(N742) );
inv1 gate83( .a(N299), .O(N748) );
inv1 gate84( .a(N303), .O(N749) );
buf1 gate85( .a(N367), .O(N750) );
inv1 gate86( .a(N307), .O(N758) );
inv1 gate87( .a(N310), .O(N759) );
inv1 gate88( .a(N313), .O(N762) );
inv1 gate89( .a(N316), .O(N768) );
inv1 gate90( .a(N319), .O(N774) );
inv1 gate91( .a(N322), .O(N780) );
inv1 gate92( .a(N325), .O(N786) );
inv1 gate93( .a(N328), .O(N794) );
inv1 gate94( .a(N331), .O(N800) );
inv1 gate95( .a(N334), .O(N806) );
inv1 gate96( .a(N337), .O(N812) );
buf1 gate97( .a(N340), .O(N813) );
inv1 gate98( .a(N340), .O(N814) );
inv1 gate99( .a(N343), .O(N821) );
inv1 gate100( .a(N346), .O(N827) );
inv1 gate101( .a(N349), .O(N833) );
inv1 gate102( .a(N352), .O(N839) );
inv1 gate103( .a(N355), .O(N845) );
inv1 gate104( .a(N358), .O(N853) );
inv1 gate105( .a(N361), .O(N859) );
inv1 gate106( .a(N364), .O(N865) );
buf1 gate107( .a(N367), .O(N871) );
nand2 gate108( .a(N467), .b(N585), .O(N881) );
inv1 gate109( .a(N528), .O(N882) );
inv1 gate110( .a(N578), .O(N883) );
inv1 gate111( .a(N575), .O(N884) );
inv1 gate112( .a(N494), .O(N885) );
and2 gate113( .a(N528), .b(N578), .O(N886) );
and2 gate114( .a(N575), .b(N494), .O(N887) );
buf1 gate115( .a(N590), .O(N889) );
buf1 gate116( .a(N657), .O(N945) );
inv1 gate117( .a(N688), .O(N957) );
and2 gate118( .a(N382), .b(N641), .O(N1028) );
nand2 gate119( .a(N382), .b(N705), .O(N1029) );
and2 gate120( .a(N469), .b(N596), .O(N1109) );

  xor2  gate5278(.a(N593), .b(N242), .O(gate121inter0));
  nand2 gate5279(.a(gate121inter0), .b(s_252), .O(gate121inter1));
  and2  gate5280(.a(N593), .b(N242), .O(gate121inter2));
  inv1  gate5281(.a(s_252), .O(gate121inter3));
  inv1  gate5282(.a(s_253), .O(gate121inter4));
  nand2 gate5283(.a(gate121inter4), .b(gate121inter3), .O(gate121inter5));
  nor2  gate5284(.a(gate121inter5), .b(gate121inter2), .O(gate121inter6));
  inv1  gate5285(.a(N242), .O(gate121inter7));
  inv1  gate5286(.a(N593), .O(gate121inter8));
  nand2 gate5287(.a(gate121inter8), .b(gate121inter7), .O(gate121inter9));
  nand2 gate5288(.a(s_253), .b(gate121inter3), .O(gate121inter10));
  nor2  gate5289(.a(gate121inter10), .b(gate121inter9), .O(gate121inter11));
  nor2  gate5290(.a(gate121inter11), .b(gate121inter6), .O(gate121inter12));
  nand2 gate5291(.a(gate121inter12), .b(gate121inter1), .O(N1110));
inv1 gate122( .a(N625), .O(N1111) );
nand2 gate123( .a(N242), .b(N593), .O(N1112) );
nand2 gate124( .a(N469), .b(N596), .O(N1113) );
inv1 gate125( .a(N625), .O(N1114) );
inv1 gate126( .a(N871), .O(N1115) );
buf1 gate127( .a(N590), .O(N1116) );
buf1 gate128( .a(N628), .O(N1119) );
buf1 gate129( .a(N682), .O(N1125) );
buf1 gate130( .a(N628), .O(N1132) );
buf1 gate131( .a(N682), .O(N1136) );
buf1 gate132( .a(N628), .O(N1141) );
buf1 gate133( .a(N682), .O(N1147) );
buf1 gate134( .a(N632), .O(N1154) );
buf1 gate135( .a(N676), .O(N1160) );
and2 gate136( .a(N700), .b(N614), .O(N1167) );
and2 gate137( .a(N700), .b(N614), .O(N1174) );
buf1 gate138( .a(N682), .O(N1175) );
buf1 gate139( .a(N676), .O(N1182) );
inv1 gate140( .a(N657), .O(N1189) );
inv1 gate141( .a(N676), .O(N1194) );
inv1 gate142( .a(N682), .O(N1199) );
inv1 gate143( .a(N689), .O(N1206) );
buf1 gate144( .a(N695), .O(N1211) );
inv1 gate145( .a(N750), .O(N1218) );
inv1 gate146( .a(N1028), .O(N1222) );
buf1 gate147( .a(N632), .O(N1227) );
buf1 gate148( .a(N676), .O(N1233) );
buf1 gate149( .a(N632), .O(N1240) );
buf1 gate150( .a(N676), .O(N1244) );
buf1 gate151( .a(N689), .O(N1249) );
buf1 gate152( .a(N689), .O(N1256) );
buf1 gate153( .a(N695), .O(N1263) );
buf1 gate154( .a(N689), .O(N1270) );
buf1 gate155( .a(N689), .O(N1277) );
buf1 gate156( .a(N700), .O(N1284) );
buf1 gate157( .a(N614), .O(N1287) );
buf1 gate158( .a(N666), .O(N1290) );
buf1 gate159( .a(N660), .O(N1293) );
buf1 gate160( .a(N651), .O(N1296) );
buf1 gate161( .a(N614), .O(N1299) );
buf1 gate162( .a(N644), .O(N1302) );
buf1 gate163( .a(N700), .O(N1305) );
buf1 gate164( .a(N614), .O(N1308) );
buf1 gate165( .a(N614), .O(N1311) );
buf1 gate166( .a(N666), .O(N1314) );
buf1 gate167( .a(N660), .O(N1317) );
buf1 gate168( .a(N651), .O(N1320) );
buf1 gate169( .a(N644), .O(N1323) );
buf1 gate170( .a(N609), .O(N1326) );
buf1 gate171( .a(N604), .O(N1329) );
buf1 gate172( .a(N742), .O(N1332) );
buf1 gate173( .a(N599), .O(N1335) );
buf1 gate174( .a(N727), .O(N1338) );
buf1 gate175( .a(N721), .O(N1341) );
buf1 gate176( .a(N715), .O(N1344) );
buf1 gate177( .a(N734), .O(N1347) );
buf1 gate178( .a(N708), .O(N1350) );
buf1 gate179( .a(N609), .O(N1353) );
buf1 gate180( .a(N604), .O(N1356) );
buf1 gate181( .a(N742), .O(N1359) );
buf1 gate182( .a(N734), .O(N1362) );
buf1 gate183( .a(N599), .O(N1365) );
buf1 gate184( .a(N727), .O(N1368) );
buf1 gate185( .a(N721), .O(N1371) );
buf1 gate186( .a(N715), .O(N1374) );
buf1 gate187( .a(N708), .O(N1377) );
buf1 gate188( .a(N806), .O(N1380) );
buf1 gate189( .a(N800), .O(N1383) );
buf1 gate190( .a(N794), .O(N1386) );
buf1 gate191( .a(N786), .O(N1389) );
buf1 gate192( .a(N780), .O(N1392) );
buf1 gate193( .a(N774), .O(N1395) );
buf1 gate194( .a(N768), .O(N1398) );
buf1 gate195( .a(N762), .O(N1401) );
buf1 gate196( .a(N806), .O(N1404) );
buf1 gate197( .a(N800), .O(N1407) );
buf1 gate198( .a(N794), .O(N1410) );
buf1 gate199( .a(N780), .O(N1413) );
buf1 gate200( .a(N774), .O(N1416) );
buf1 gate201( .a(N768), .O(N1419) );
buf1 gate202( .a(N762), .O(N1422) );
buf1 gate203( .a(N786), .O(N1425) );
buf1 gate204( .a(N636), .O(N1428) );
buf1 gate205( .a(N636), .O(N1431) );
buf1 gate206( .a(N865), .O(N1434) );
buf1 gate207( .a(N859), .O(N1437) );
buf1 gate208( .a(N853), .O(N1440) );
buf1 gate209( .a(N845), .O(N1443) );
buf1 gate210( .a(N839), .O(N1446) );
buf1 gate211( .a(N833), .O(N1449) );
buf1 gate212( .a(N827), .O(N1452) );
buf1 gate213( .a(N821), .O(N1455) );
buf1 gate214( .a(N814), .O(N1458) );
buf1 gate215( .a(N865), .O(N1461) );
buf1 gate216( .a(N859), .O(N1464) );
buf1 gate217( .a(N853), .O(N1467) );
buf1 gate218( .a(N839), .O(N1470) );
buf1 gate219( .a(N833), .O(N1473) );
buf1 gate220( .a(N827), .O(N1476) );
buf1 gate221( .a(N821), .O(N1479) );
buf1 gate222( .a(N845), .O(N1482) );
buf1 gate223( .a(N814), .O(N1485) );
inv1 gate224( .a(N1109), .O(N1489) );
buf1 gate225( .a(N1116), .O(N1490) );
and2 gate226( .a(N957), .b(N614), .O(N1537) );
and2 gate227( .a(N614), .b(N957), .O(N1551) );
and2 gate228( .a(N1029), .b(N636), .O(N1649) );
buf1 gate229( .a(N957), .O(N1703) );
nor2 gate230( .a(N957), .b(N614), .O(N1708) );
buf1 gate231( .a(N957), .O(N1713) );
nor2 gate232( .a(N614), .b(N957), .O(N1721) );
buf1 gate233( .a(N1029), .O(N1758) );
and2 gate234( .a(N163), .b(N1116), .O(N1781) );
and2 gate235( .a(N170), .b(N1125), .O(N1782) );
inv1 gate236( .a(N1125), .O(N1783) );
inv1 gate237( .a(N1136), .O(N1789) );
and2 gate238( .a(N169), .b(N1125), .O(N1793) );
and2 gate239( .a(N168), .b(N1125), .O(N1794) );
and2 gate240( .a(N167), .b(N1125), .O(N1795) );
and2 gate241( .a(N166), .b(N1136), .O(N1796) );
and2 gate242( .a(N165), .b(N1136), .O(N1797) );
and2 gate243( .a(N164), .b(N1136), .O(N1798) );
inv1 gate244( .a(N1147), .O(N1799) );
inv1 gate245( .a(N1160), .O(N1805) );
and2 gate246( .a(N177), .b(N1147), .O(N1811) );
and2 gate247( .a(N176), .b(N1147), .O(N1812) );
and2 gate248( .a(N175), .b(N1147), .O(N1813) );
and2 gate249( .a(N174), .b(N1147), .O(N1814) );
and2 gate250( .a(N173), .b(N1147), .O(N1815) );
and2 gate251( .a(N157), .b(N1160), .O(N1816) );
and2 gate252( .a(N156), .b(N1160), .O(N1817) );
and2 gate253( .a(N155), .b(N1160), .O(N1818) );
and2 gate254( .a(N154), .b(N1160), .O(N1819) );
and2 gate255( .a(N153), .b(N1160), .O(N1820) );
inv1 gate256( .a(N1284), .O(N1821) );
inv1 gate257( .a(N1287), .O(N1822) );
inv1 gate258( .a(N1290), .O(N1828) );
inv1 gate259( .a(N1293), .O(N1829) );
inv1 gate260( .a(N1296), .O(N1830) );
inv1 gate261( .a(N1299), .O(N1832) );
inv1 gate262( .a(N1302), .O(N1833) );
inv1 gate263( .a(N1305), .O(N1834) );
inv1 gate264( .a(N1308), .O(N1835) );
inv1 gate265( .a(N1311), .O(N1839) );
inv1 gate266( .a(N1314), .O(N1840) );
inv1 gate267( .a(N1317), .O(N1841) );
inv1 gate268( .a(N1320), .O(N1842) );
inv1 gate269( .a(N1323), .O(N1843) );
inv1 gate270( .a(N1175), .O(N1845) );
inv1 gate271( .a(N1182), .O(N1851) );
and2 gate272( .a(N181), .b(N1175), .O(N1857) );
and2 gate273( .a(N171), .b(N1175), .O(N1858) );
and2 gate274( .a(N180), .b(N1175), .O(N1859) );
and2 gate275( .a(N179), .b(N1175), .O(N1860) );
and2 gate276( .a(N178), .b(N1175), .O(N1861) );
and2 gate277( .a(N161), .b(N1182), .O(N1862) );
and2 gate278( .a(N151), .b(N1182), .O(N1863) );
and2 gate279( .a(N160), .b(N1182), .O(N1864) );
and2 gate280( .a(N159), .b(N1182), .O(N1865) );
and2 gate281( .a(N158), .b(N1182), .O(N1866) );
inv1 gate282( .a(N1326), .O(N1867) );
inv1 gate283( .a(N1329), .O(N1868) );
inv1 gate284( .a(N1332), .O(N1869) );
inv1 gate285( .a(N1335), .O(N1870) );
inv1 gate286( .a(N1338), .O(N1871) );
inv1 gate287( .a(N1341), .O(N1872) );
inv1 gate288( .a(N1344), .O(N1873) );
inv1 gate289( .a(N1347), .O(N1874) );
inv1 gate290( .a(N1350), .O(N1875) );
inv1 gate291( .a(N1353), .O(N1876) );
inv1 gate292( .a(N1356), .O(N1877) );
inv1 gate293( .a(N1359), .O(N1878) );
inv1 gate294( .a(N1362), .O(N1879) );
inv1 gate295( .a(N1365), .O(N1880) );
inv1 gate296( .a(N1368), .O(N1881) );
inv1 gate297( .a(N1371), .O(N1882) );
inv1 gate298( .a(N1374), .O(N1883) );
inv1 gate299( .a(N1377), .O(N1884) );
buf1 gate300( .a(N1199), .O(N1885) );
buf1 gate301( .a(N1194), .O(N1892) );
buf1 gate302( .a(N1199), .O(N1899) );
buf1 gate303( .a(N1194), .O(N1906) );
inv1 gate304( .a(N1211), .O(N1913) );
buf1 gate305( .a(N1194), .O(N1919) );
and2 gate306( .a(N44), .b(N1211), .O(N1926) );
and2 gate307( .a(N41), .b(N1211), .O(N1927) );
and2 gate308( .a(N29), .b(N1211), .O(N1928) );
and2 gate309( .a(N26), .b(N1211), .O(N1929) );
and2 gate310( .a(N23), .b(N1211), .O(N1930) );
inv1 gate311( .a(N1380), .O(N1931) );
inv1 gate312( .a(N1383), .O(N1932) );
inv1 gate313( .a(N1386), .O(N1933) );
inv1 gate314( .a(N1389), .O(N1934) );
inv1 gate315( .a(N1392), .O(N1935) );
inv1 gate316( .a(N1395), .O(N1936) );
inv1 gate317( .a(N1398), .O(N1937) );
inv1 gate318( .a(N1401), .O(N1938) );
inv1 gate319( .a(N1404), .O(N1939) );
inv1 gate320( .a(N1407), .O(N1940) );
inv1 gate321( .a(N1410), .O(N1941) );
inv1 gate322( .a(N1413), .O(N1942) );
inv1 gate323( .a(N1416), .O(N1943) );
inv1 gate324( .a(N1419), .O(N1944) );
inv1 gate325( .a(N1422), .O(N1945) );
inv1 gate326( .a(N1425), .O(N1946) );
inv1 gate327( .a(N1233), .O(N1947) );
inv1 gate328( .a(N1244), .O(N1953) );
and2 gate329( .a(N209), .b(N1233), .O(N1957) );
and2 gate330( .a(N216), .b(N1233), .O(N1958) );
and2 gate331( .a(N215), .b(N1233), .O(N1959) );
and2 gate332( .a(N214), .b(N1233), .O(N1960) );
and2 gate333( .a(N213), .b(N1244), .O(N1961) );
and2 gate334( .a(N212), .b(N1244), .O(N1962) );
and2 gate335( .a(N211), .b(N1244), .O(N1963) );
inv1 gate336( .a(N1428), .O(N1965) );
and2 gate337( .a(N1222), .b(N636), .O(N1966) );
inv1 gate338( .a(N1431), .O(N1967) );
inv1 gate339( .a(N1434), .O(N1968) );
inv1 gate340( .a(N1437), .O(N1969) );
inv1 gate341( .a(N1440), .O(N1970) );
inv1 gate342( .a(N1443), .O(N1971) );
inv1 gate343( .a(N1446), .O(N1972) );
inv1 gate344( .a(N1449), .O(N1973) );
inv1 gate345( .a(N1452), .O(N1974) );
inv1 gate346( .a(N1455), .O(N1975) );
inv1 gate347( .a(N1458), .O(N1976) );
inv1 gate348( .a(N1249), .O(N1977) );
inv1 gate349( .a(N1256), .O(N1983) );
and2 gate350( .a(N642), .b(N1249), .O(N1989) );
and2 gate351( .a(N644), .b(N1249), .O(N1990) );
and2 gate352( .a(N651), .b(N1249), .O(N1991) );
and2 gate353( .a(N674), .b(N1249), .O(N1992) );
and2 gate354( .a(N660), .b(N1249), .O(N1993) );
and2 gate355( .a(N666), .b(N1256), .O(N1994) );
and2 gate356( .a(N672), .b(N1256), .O(N1995) );
and2 gate357( .a(N673), .b(N1256), .O(N1996) );
inv1 gate358( .a(N1263), .O(N1997) );
buf1 gate359( .a(N1194), .O(N2003) );
and2 gate360( .a(N47), .b(N1263), .O(N2010) );
and2 gate361( .a(N35), .b(N1263), .O(N2011) );
and2 gate362( .a(N32), .b(N1263), .O(N2012) );
and2 gate363( .a(N50), .b(N1263), .O(N2013) );
and2 gate364( .a(N66), .b(N1263), .O(N2014) );
inv1 gate365( .a(N1461), .O(N2015) );
inv1 gate366( .a(N1464), .O(N2016) );
inv1 gate367( .a(N1467), .O(N2017) );
inv1 gate368( .a(N1470), .O(N2018) );
inv1 gate369( .a(N1473), .O(N2019) );
inv1 gate370( .a(N1476), .O(N2020) );
inv1 gate371( .a(N1479), .O(N2021) );
inv1 gate372( .a(N1482), .O(N2022) );
inv1 gate373( .a(N1485), .O(N2023) );
buf1 gate374( .a(N1206), .O(N2024) );
buf1 gate375( .a(N1206), .O(N2031) );
buf1 gate376( .a(N1206), .O(N2038) );
buf1 gate377( .a(N1206), .O(N2045) );
inv1 gate378( .a(N1270), .O(N2052) );
inv1 gate379( .a(N1277), .O(N2058) );
and2 gate380( .a(N706), .b(N1270), .O(N2064) );
and2 gate381( .a(N708), .b(N1270), .O(N2065) );
and2 gate382( .a(N715), .b(N1270), .O(N2066) );
and2 gate383( .a(N721), .b(N1270), .O(N2067) );
and2 gate384( .a(N727), .b(N1270), .O(N2068) );
and2 gate385( .a(N733), .b(N1277), .O(N2069) );
and2 gate386( .a(N734), .b(N1277), .O(N2070) );
and2 gate387( .a(N742), .b(N1277), .O(N2071) );
and2 gate388( .a(N748), .b(N1277), .O(N2072) );
and2 gate389( .a(N749), .b(N1277), .O(N2073) );
buf1 gate390( .a(N1189), .O(N2074) );
buf1 gate391( .a(N1189), .O(N2081) );
buf1 gate392( .a(N1222), .O(N2086) );
nand2 gate393( .a(N1287), .b(N1821), .O(N2107) );
nand2 gate394( .a(N1284), .b(N1822), .O(N2108) );
inv1 gate395( .a(N1703), .O(N2110) );
nand2 gate396( .a(N1703), .b(N1832), .O(N2111) );
nand2 gate397( .a(N1308), .b(N1834), .O(N2112) );
nand2 gate398( .a(N1305), .b(N1835), .O(N2113) );
inv1 gate399( .a(N1713), .O(N2114) );
nand2 gate400( .a(N1713), .b(N1839), .O(N2115) );
inv1 gate401( .a(N1721), .O(N2117) );
inv1 gate402( .a(N1758), .O(N2171) );
nand2 gate403( .a(N1758), .b(N1965), .O(N2172) );
inv1 gate404( .a(N1708), .O(N2230) );
buf1 gate405( .a(N1537), .O(N2231) );
buf1 gate406( .a(N1551), .O(N2235) );
or2 gate407( .a(N1783), .b(N1782), .O(N2239) );
or2 gate408( .a(N1783), .b(N1125), .O(N2240) );
or2 gate409( .a(N1783), .b(N1793), .O(N2241) );
or2 gate410( .a(N1783), .b(N1794), .O(N2242) );
or2 gate411( .a(N1783), .b(N1795), .O(N2243) );
or2 gate412( .a(N1789), .b(N1796), .O(N2244) );
or2 gate413( .a(N1789), .b(N1797), .O(N2245) );
or2 gate414( .a(N1789), .b(N1798), .O(N2246) );
or2 gate415( .a(N1799), .b(N1811), .O(N2247) );
or2 gate416( .a(N1799), .b(N1812), .O(N2248) );
or2 gate417( .a(N1799), .b(N1813), .O(N2249) );
or2 gate418( .a(N1799), .b(N1814), .O(N2250) );
or2 gate419( .a(N1799), .b(N1815), .O(N2251) );
or2 gate420( .a(N1805), .b(N1816), .O(N2252) );
or2 gate421( .a(N1805), .b(N1817), .O(N2253) );
or2 gate422( .a(N1805), .b(N1818), .O(N2254) );
or2 gate423( .a(N1805), .b(N1819), .O(N2255) );
or2 gate424( .a(N1805), .b(N1820), .O(N2256) );
nand2 gate425( .a(N2107), .b(N2108), .O(N2257) );
inv1 gate426( .a(N2074), .O(N2267) );
nand2 gate427( .a(N1299), .b(N2110), .O(N2268) );
nand2 gate428( .a(N2112), .b(N2113), .O(N2269) );
nand2 gate429( .a(N1311), .b(N2114), .O(N2274) );
inv1 gate430( .a(N2081), .O(N2275) );
and2 gate431( .a(N141), .b(N1845), .O(N2277) );
and2 gate432( .a(N147), .b(N1845), .O(N2278) );
and2 gate433( .a(N138), .b(N1845), .O(N2279) );
and2 gate434( .a(N144), .b(N1845), .O(N2280) );
and2 gate435( .a(N135), .b(N1845), .O(N2281) );
and2 gate436( .a(N141), .b(N1851), .O(N2282) );
and2 gate437( .a(N147), .b(N1851), .O(N2283) );
and2 gate438( .a(N138), .b(N1851), .O(N2284) );
and2 gate439( .a(N144), .b(N1851), .O(N2285) );
and2 gate440( .a(N135), .b(N1851), .O(N2286) );
inv1 gate441( .a(N1885), .O(N2287) );
inv1 gate442( .a(N1892), .O(N2293) );
and2 gate443( .a(N103), .b(N1885), .O(N2299) );
and2 gate444( .a(N130), .b(N1885), .O(N2300) );
and2 gate445( .a(N127), .b(N1885), .O(N2301) );
and2 gate446( .a(N124), .b(N1885), .O(N2302) );
and2 gate447( .a(N100), .b(N1885), .O(N2303) );
and2 gate448( .a(N103), .b(N1892), .O(N2304) );
and2 gate449( .a(N130), .b(N1892), .O(N2305) );
and2 gate450( .a(N127), .b(N1892), .O(N2306) );
and2 gate451( .a(N124), .b(N1892), .O(N2307) );
and2 gate452( .a(N100), .b(N1892), .O(N2308) );
inv1 gate453( .a(N1899), .O(N2309) );
inv1 gate454( .a(N1906), .O(N2315) );
and2 gate455( .a(N115), .b(N1899), .O(N2321) );
and2 gate456( .a(N118), .b(N1899), .O(N2322) );
and2 gate457( .a(N97), .b(N1899), .O(N2323) );
and2 gate458( .a(N94), .b(N1899), .O(N2324) );
and2 gate459( .a(N121), .b(N1899), .O(N2325) );
and2 gate460( .a(N115), .b(N1906), .O(N2326) );
and2 gate461( .a(N118), .b(N1906), .O(N2327) );
and2 gate462( .a(N97), .b(N1906), .O(N2328) );
and2 gate463( .a(N94), .b(N1906), .O(N2329) );
and2 gate464( .a(N121), .b(N1906), .O(N2330) );
inv1 gate465( .a(N1919), .O(N2331) );
and2 gate466( .a(N208), .b(N1913), .O(N2337) );
and2 gate467( .a(N198), .b(N1913), .O(N2338) );
and2 gate468( .a(N207), .b(N1913), .O(N2339) );
and2 gate469( .a(N206), .b(N1913), .O(N2340) );
and2 gate470( .a(N205), .b(N1913), .O(N2341) );
and2 gate471( .a(N44), .b(N1919), .O(N2342) );
and2 gate472( .a(N41), .b(N1919), .O(N2343) );
and2 gate473( .a(N29), .b(N1919), .O(N2344) );
and2 gate474( .a(N26), .b(N1919), .O(N2345) );
and2 gate475( .a(N23), .b(N1919), .O(N2346) );
or2 gate476( .a(N1947), .b(N1233), .O(N2347) );
or2 gate477( .a(N1947), .b(N1957), .O(N2348) );
or2 gate478( .a(N1947), .b(N1958), .O(N2349) );
or2 gate479( .a(N1947), .b(N1959), .O(N2350) );
or2 gate480( .a(N1947), .b(N1960), .O(N2351) );
or2 gate481( .a(N1953), .b(N1961), .O(N2352) );
or2 gate482( .a(N1953), .b(N1962), .O(N2353) );
or2 gate483( .a(N1953), .b(N1963), .O(N2354) );

  xor2  gate3556(.a(N2171), .b(N1428), .O(gate484inter0));
  nand2 gate3557(.a(gate484inter0), .b(s_6), .O(gate484inter1));
  and2  gate3558(.a(N2171), .b(N1428), .O(gate484inter2));
  inv1  gate3559(.a(s_6), .O(gate484inter3));
  inv1  gate3560(.a(s_7), .O(gate484inter4));
  nand2 gate3561(.a(gate484inter4), .b(gate484inter3), .O(gate484inter5));
  nor2  gate3562(.a(gate484inter5), .b(gate484inter2), .O(gate484inter6));
  inv1  gate3563(.a(N1428), .O(gate484inter7));
  inv1  gate3564(.a(N2171), .O(gate484inter8));
  nand2 gate3565(.a(gate484inter8), .b(gate484inter7), .O(gate484inter9));
  nand2 gate3566(.a(s_7), .b(gate484inter3), .O(gate484inter10));
  nor2  gate3567(.a(gate484inter10), .b(gate484inter9), .O(gate484inter11));
  nor2  gate3568(.a(gate484inter11), .b(gate484inter6), .O(gate484inter12));
  nand2 gate3569(.a(gate484inter12), .b(gate484inter1), .O(N2355));
inv1 gate485( .a(N2086), .O(N2356) );
nand2 gate486( .a(N2086), .b(N1967), .O(N2357) );
and2 gate487( .a(N114), .b(N1977), .O(N2358) );
and2 gate488( .a(N113), .b(N1977), .O(N2359) );
and2 gate489( .a(N111), .b(N1977), .O(N2360) );
and2 gate490( .a(N87), .b(N1977), .O(N2361) );
and2 gate491( .a(N112), .b(N1977), .O(N2362) );
and2 gate492( .a(N88), .b(N1983), .O(N2363) );
and2 gate493( .a(N245), .b(N1983), .O(N2364) );
and2 gate494( .a(N271), .b(N1983), .O(N2365) );
and2 gate495( .a(N759), .b(N1983), .O(N2366) );
and2 gate496( .a(N70), .b(N1983), .O(N2367) );
inv1 gate497( .a(N2003), .O(N2368) );
and2 gate498( .a(N193), .b(N1997), .O(N2374) );
and2 gate499( .a(N192), .b(N1997), .O(N2375) );
and2 gate500( .a(N191), .b(N1997), .O(N2376) );
and2 gate501( .a(N190), .b(N1997), .O(N2377) );
and2 gate502( .a(N189), .b(N1997), .O(N2378) );
and2 gate503( .a(N47), .b(N2003), .O(N2379) );
and2 gate504( .a(N35), .b(N2003), .O(N2380) );
and2 gate505( .a(N32), .b(N2003), .O(N2381) );
and2 gate506( .a(N50), .b(N2003), .O(N2382) );
and2 gate507( .a(N66), .b(N2003), .O(N2383) );
inv1 gate508( .a(N2024), .O(N2384) );
inv1 gate509( .a(N2031), .O(N2390) );
and2 gate510( .a(N58), .b(N2024), .O(N2396) );
and2 gate511( .a(N77), .b(N2024), .O(N2397) );
and2 gate512( .a(N78), .b(N2024), .O(N2398) );
and2 gate513( .a(N59), .b(N2024), .O(N2399) );
and2 gate514( .a(N81), .b(N2024), .O(N2400) );
and2 gate515( .a(N80), .b(N2031), .O(N2401) );
and2 gate516( .a(N79), .b(N2031), .O(N2402) );
and2 gate517( .a(N60), .b(N2031), .O(N2403) );
and2 gate518( .a(N61), .b(N2031), .O(N2404) );
and2 gate519( .a(N62), .b(N2031), .O(N2405) );
inv1 gate520( .a(N2038), .O(N2406) );
inv1 gate521( .a(N2045), .O(N2412) );
and2 gate522( .a(N69), .b(N2038), .O(N2418) );
and2 gate523( .a(N70), .b(N2038), .O(N2419) );
and2 gate524( .a(N74), .b(N2038), .O(N2420) );
and2 gate525( .a(N76), .b(N2038), .O(N2421) );
and2 gate526( .a(N75), .b(N2038), .O(N2422) );
and2 gate527( .a(N73), .b(N2045), .O(N2423) );
and2 gate528( .a(N53), .b(N2045), .O(N2424) );
and2 gate529( .a(N54), .b(N2045), .O(N2425) );
and2 gate530( .a(N55), .b(N2045), .O(N2426) );
and2 gate531( .a(N56), .b(N2045), .O(N2427) );
and2 gate532( .a(N82), .b(N2052), .O(N2428) );
and2 gate533( .a(N65), .b(N2052), .O(N2429) );
and2 gate534( .a(N83), .b(N2052), .O(N2430) );
and2 gate535( .a(N84), .b(N2052), .O(N2431) );
and2 gate536( .a(N85), .b(N2052), .O(N2432) );
and2 gate537( .a(N64), .b(N2058), .O(N2433) );
and2 gate538( .a(N63), .b(N2058), .O(N2434) );
and2 gate539( .a(N86), .b(N2058), .O(N2435) );
and2 gate540( .a(N109), .b(N2058), .O(N2436) );
and2 gate541( .a(N110), .b(N2058), .O(N2437) );
and2 gate542( .a(N2239), .b(N1119), .O(N2441) );
and2 gate543( .a(N2240), .b(N1119), .O(N2442) );
and2 gate544( .a(N2241), .b(N1119), .O(N2446) );
and2 gate545( .a(N2242), .b(N1119), .O(N2450) );
and2 gate546( .a(N2243), .b(N1119), .O(N2454) );
and2 gate547( .a(N2244), .b(N1132), .O(N2458) );
and2 gate548( .a(N2247), .b(N1141), .O(N2462) );
and2 gate549( .a(N2248), .b(N1141), .O(N2466) );
and2 gate550( .a(N2249), .b(N1141), .O(N2470) );
and2 gate551( .a(N2250), .b(N1141), .O(N2474) );
and2 gate552( .a(N2251), .b(N1141), .O(N2478) );
and2 gate553( .a(N2252), .b(N1154), .O(N2482) );
and2 gate554( .a(N2253), .b(N1154), .O(N2488) );
and2 gate555( .a(N2254), .b(N1154), .O(N2496) );
and2 gate556( .a(N2255), .b(N1154), .O(N2502) );
and2 gate557( .a(N2256), .b(N1154), .O(N2508) );
nand2 gate558( .a(N2268), .b(N2111), .O(N2523) );
nand2 gate559( .a(N2274), .b(N2115), .O(N2533) );
inv1 gate560( .a(N2235), .O(N2537) );
or2 gate561( .a(N2278), .b(N1858), .O(N2538) );
or2 gate562( .a(N2279), .b(N1859), .O(N2542) );
or2 gate563( .a(N2280), .b(N1860), .O(N2546) );
or2 gate564( .a(N2281), .b(N1861), .O(N2550) );
or2 gate565( .a(N2283), .b(N1863), .O(N2554) );
or2 gate566( .a(N2284), .b(N1864), .O(N2561) );
or2 gate567( .a(N2285), .b(N1865), .O(N2567) );
or2 gate568( .a(N2286), .b(N1866), .O(N2573) );
or2 gate569( .a(N2338), .b(N1927), .O(N2604) );
or2 gate570( .a(N2339), .b(N1928), .O(N2607) );
or2 gate571( .a(N2340), .b(N1929), .O(N2611) );
or2 gate572( .a(N2341), .b(N1930), .O(N2615) );
and2 gate573( .a(N2348), .b(N1227), .O(N2619) );
and2 gate574( .a(N2349), .b(N1227), .O(N2626) );
and2 gate575( .a(N2350), .b(N1227), .O(N2632) );
and2 gate576( .a(N2351), .b(N1227), .O(N2638) );
and2 gate577( .a(N2352), .b(N1240), .O(N2644) );
nand2 gate578( .a(N2355), .b(N2172), .O(N2650) );

  xor2  gate4816(.a(N2356), .b(N1431), .O(gate579inter0));
  nand2 gate4817(.a(gate579inter0), .b(s_186), .O(gate579inter1));
  and2  gate4818(.a(N2356), .b(N1431), .O(gate579inter2));
  inv1  gate4819(.a(s_186), .O(gate579inter3));
  inv1  gate4820(.a(s_187), .O(gate579inter4));
  nand2 gate4821(.a(gate579inter4), .b(gate579inter3), .O(gate579inter5));
  nor2  gate4822(.a(gate579inter5), .b(gate579inter2), .O(gate579inter6));
  inv1  gate4823(.a(N1431), .O(gate579inter7));
  inv1  gate4824(.a(N2356), .O(gate579inter8));
  nand2 gate4825(.a(gate579inter8), .b(gate579inter7), .O(gate579inter9));
  nand2 gate4826(.a(s_187), .b(gate579inter3), .O(gate579inter10));
  nor2  gate4827(.a(gate579inter10), .b(gate579inter9), .O(gate579inter11));
  nor2  gate4828(.a(gate579inter11), .b(gate579inter6), .O(gate579inter12));
  nand2 gate4829(.a(gate579inter12), .b(gate579inter1), .O(N2653));
or2 gate580( .a(N2359), .b(N1990), .O(N2654) );
or2 gate581( .a(N2360), .b(N1991), .O(N2658) );
or2 gate582( .a(N2361), .b(N1992), .O(N2662) );
or2 gate583( .a(N2362), .b(N1993), .O(N2666) );
or2 gate584( .a(N2363), .b(N1994), .O(N2670) );
or2 gate585( .a(N2366), .b(N1256), .O(N2674) );
or2 gate586( .a(N2367), .b(N1256), .O(N2680) );
or2 gate587( .a(N2374), .b(N2010), .O(N2688) );
or2 gate588( .a(N2375), .b(N2011), .O(N2692) );
or2 gate589( .a(N2376), .b(N2012), .O(N2696) );
or2 gate590( .a(N2377), .b(N2013), .O(N2700) );
or2 gate591( .a(N2378), .b(N2014), .O(N2704) );
and2 gate592( .a(N2347), .b(N1227), .O(N2728) );
or2 gate593( .a(N2429), .b(N2065), .O(N2729) );
or2 gate594( .a(N2430), .b(N2066), .O(N2733) );
or2 gate595( .a(N2431), .b(N2067), .O(N2737) );
or2 gate596( .a(N2432), .b(N2068), .O(N2741) );
or2 gate597( .a(N2433), .b(N2069), .O(N2745) );
or2 gate598( .a(N2434), .b(N2070), .O(N2749) );
or2 gate599( .a(N2435), .b(N2071), .O(N2753) );
or2 gate600( .a(N2436), .b(N2072), .O(N2757) );
or2 gate601( .a(N2437), .b(N2073), .O(N2761) );
inv1 gate602( .a(N2231), .O(N2765) );
and2 gate603( .a(N2354), .b(N1240), .O(N2766) );
and2 gate604( .a(N2353), .b(N1240), .O(N2769) );
and2 gate605( .a(N2246), .b(N1132), .O(N2772) );
and2 gate606( .a(N2245), .b(N1132), .O(N2775) );
or2 gate607( .a(N2282), .b(N1862), .O(N2778) );
or2 gate608( .a(N2358), .b(N1989), .O(N2781) );
or2 gate609( .a(N2365), .b(N1996), .O(N2784) );
or2 gate610( .a(N2364), .b(N1995), .O(N2787) );
or2 gate611( .a(N2337), .b(N1926), .O(N2790) );
or2 gate612( .a(N2277), .b(N1857), .O(N2793) );
or2 gate613( .a(N2428), .b(N2064), .O(N2796) );
and2 gate614( .a(N2257), .b(N1537), .O(N2866) );
and2 gate615( .a(N2257), .b(N1537), .O(N2867) );
and2 gate616( .a(N2257), .b(N1537), .O(N2868) );
and2 gate617( .a(N2257), .b(N1537), .O(N2869) );
and2 gate618( .a(N2269), .b(N1551), .O(N2878) );
and2 gate619( .a(N204), .b(N2287), .O(N2913) );
and2 gate620( .a(N203), .b(N2287), .O(N2914) );
and2 gate621( .a(N202), .b(N2287), .O(N2915) );
and2 gate622( .a(N201), .b(N2287), .O(N2916) );
and2 gate623( .a(N200), .b(N2287), .O(N2917) );
and2 gate624( .a(N235), .b(N2293), .O(N2918) );
and2 gate625( .a(N234), .b(N2293), .O(N2919) );
and2 gate626( .a(N233), .b(N2293), .O(N2920) );
and2 gate627( .a(N232), .b(N2293), .O(N2921) );
and2 gate628( .a(N231), .b(N2293), .O(N2922) );
and2 gate629( .a(N197), .b(N2309), .O(N2923) );
and2 gate630( .a(N187), .b(N2309), .O(N2924) );
and2 gate631( .a(N196), .b(N2309), .O(N2925) );
and2 gate632( .a(N195), .b(N2309), .O(N2926) );
and2 gate633( .a(N194), .b(N2309), .O(N2927) );
and2 gate634( .a(N227), .b(N2315), .O(N2928) );
and2 gate635( .a(N217), .b(N2315), .O(N2929) );
and2 gate636( .a(N226), .b(N2315), .O(N2930) );
and2 gate637( .a(N225), .b(N2315), .O(N2931) );
and2 gate638( .a(N224), .b(N2315), .O(N2932) );
and2 gate639( .a(N239), .b(N2331), .O(N2933) );
and2 gate640( .a(N229), .b(N2331), .O(N2934) );
and2 gate641( .a(N238), .b(N2331), .O(N2935) );
and2 gate642( .a(N237), .b(N2331), .O(N2936) );
and2 gate643( .a(N236), .b(N2331), .O(N2937) );
nand2 gate644( .a(N2653), .b(N2357), .O(N2988) );
and2 gate645( .a(N223), .b(N2368), .O(N3005) );
and2 gate646( .a(N222), .b(N2368), .O(N3006) );
and2 gate647( .a(N221), .b(N2368), .O(N3007) );
and2 gate648( .a(N220), .b(N2368), .O(N3008) );
and2 gate649( .a(N219), .b(N2368), .O(N3009) );
and2 gate650( .a(N812), .b(N2384), .O(N3020) );
and2 gate651( .a(N814), .b(N2384), .O(N3021) );
and2 gate652( .a(N821), .b(N2384), .O(N3022) );
and2 gate653( .a(N827), .b(N2384), .O(N3023) );
and2 gate654( .a(N833), .b(N2384), .O(N3024) );
and2 gate655( .a(N839), .b(N2390), .O(N3025) );
and2 gate656( .a(N845), .b(N2390), .O(N3026) );
and2 gate657( .a(N853), .b(N2390), .O(N3027) );
and2 gate658( .a(N859), .b(N2390), .O(N3028) );
and2 gate659( .a(N865), .b(N2390), .O(N3029) );
and2 gate660( .a(N758), .b(N2406), .O(N3032) );
and2 gate661( .a(N759), .b(N2406), .O(N3033) );
and2 gate662( .a(N762), .b(N2406), .O(N3034) );
and2 gate663( .a(N768), .b(N2406), .O(N3035) );
and2 gate664( .a(N774), .b(N2406), .O(N3036) );
and2 gate665( .a(N780), .b(N2412), .O(N3037) );
and2 gate666( .a(N786), .b(N2412), .O(N3038) );
and2 gate667( .a(N794), .b(N2412), .O(N3039) );
and2 gate668( .a(N800), .b(N2412), .O(N3040) );
and2 gate669( .a(N806), .b(N2412), .O(N3041) );
buf1 gate670( .a(N2257), .O(N3061) );
buf1 gate671( .a(N2257), .O(N3064) );
buf1 gate672( .a(N2269), .O(N3067) );
buf1 gate673( .a(N2269), .O(N3070) );
inv1 gate674( .a(N2728), .O(N3073) );
inv1 gate675( .a(N2441), .O(N3080) );
and2 gate676( .a(N666), .b(N2644), .O(N3096) );
and2 gate677( .a(N660), .b(N2638), .O(N3097) );
and2 gate678( .a(N1189), .b(N2632), .O(N3101) );
and2 gate679( .a(N651), .b(N2626), .O(N3107) );
and2 gate680( .a(N644), .b(N2619), .O(N3114) );
and2 gate681( .a(N2523), .b(N2257), .O(N3122) );
or2 gate682( .a(N1167), .b(N2866), .O(N3126) );
and2 gate683( .a(N2523), .b(N2257), .O(N3130) );
or2 gate684( .a(N1167), .b(N2869), .O(N3131) );
and2 gate685( .a(N2523), .b(N2257), .O(N3134) );
inv1 gate686( .a(N2533), .O(N3135) );
and2 gate687( .a(N666), .b(N2644), .O(N3136) );
and2 gate688( .a(N660), .b(N2638), .O(N3137) );
and2 gate689( .a(N1189), .b(N2632), .O(N3140) );
and2 gate690( .a(N651), .b(N2626), .O(N3144) );
and2 gate691( .a(N644), .b(N2619), .O(N3149) );
and2 gate692( .a(N2533), .b(N2269), .O(N3155) );
or2 gate693( .a(N1174), .b(N2878), .O(N3159) );
inv1 gate694( .a(N2778), .O(N3167) );
and2 gate695( .a(N609), .b(N2508), .O(N3168) );
and2 gate696( .a(N604), .b(N2502), .O(N3169) );
and2 gate697( .a(N742), .b(N2496), .O(N3173) );
and2 gate698( .a(N734), .b(N2488), .O(N3178) );
and2 gate699( .a(N599), .b(N2482), .O(N3184) );
and2 gate700( .a(N727), .b(N2573), .O(N3185) );
and2 gate701( .a(N721), .b(N2567), .O(N3189) );
and2 gate702( .a(N715), .b(N2561), .O(N3195) );
and2 gate703( .a(N708), .b(N2554), .O(N3202) );
and2 gate704( .a(N609), .b(N2508), .O(N3210) );
and2 gate705( .a(N604), .b(N2502), .O(N3211) );
and2 gate706( .a(N742), .b(N2496), .O(N3215) );
and2 gate707( .a(N2488), .b(N734), .O(N3221) );
and2 gate708( .a(N599), .b(N2482), .O(N3228) );
and2 gate709( .a(N727), .b(N2573), .O(N3229) );
and2 gate710( .a(N721), .b(N2567), .O(N3232) );
and2 gate711( .a(N715), .b(N2561), .O(N3236) );
and2 gate712( .a(N708), .b(N2554), .O(N3241) );
or2 gate713( .a(N2913), .b(N2299), .O(N3247) );
or2 gate714( .a(N2914), .b(N2300), .O(N3251) );
or2 gate715( .a(N2915), .b(N2301), .O(N3255) );
or2 gate716( .a(N2916), .b(N2302), .O(N3259) );
or2 gate717( .a(N2917), .b(N2303), .O(N3263) );
or2 gate718( .a(N2918), .b(N2304), .O(N3267) );
or2 gate719( .a(N2919), .b(N2305), .O(N3273) );
or2 gate720( .a(N2920), .b(N2306), .O(N3281) );
or2 gate721( .a(N2921), .b(N2307), .O(N3287) );
or2 gate722( .a(N2922), .b(N2308), .O(N3293) );
or2 gate723( .a(N2924), .b(N2322), .O(N3299) );
or2 gate724( .a(N2925), .b(N2323), .O(N3303) );
or2 gate725( .a(N2926), .b(N2324), .O(N3307) );
or2 gate726( .a(N2927), .b(N2325), .O(N3311) );
or2 gate727( .a(N2929), .b(N2327), .O(N3315) );
or2 gate728( .a(N2930), .b(N2328), .O(N3322) );
or2 gate729( .a(N2931), .b(N2329), .O(N3328) );
or2 gate730( .a(N2932), .b(N2330), .O(N3334) );
or2 gate731( .a(N2934), .b(N2343), .O(N3340) );
or2 gate732( .a(N2935), .b(N2344), .O(N3343) );
or2 gate733( .a(N2936), .b(N2345), .O(N3349) );
or2 gate734( .a(N2937), .b(N2346), .O(N3355) );
and2 gate735( .a(N2761), .b(N2478), .O(N3361) );
and2 gate736( .a(N2757), .b(N2474), .O(N3362) );
and2 gate737( .a(N2753), .b(N2470), .O(N3363) );
and2 gate738( .a(N2749), .b(N2466), .O(N3364) );
and2 gate739( .a(N2745), .b(N2462), .O(N3365) );
and2 gate740( .a(N2741), .b(N2550), .O(N3366) );
and2 gate741( .a(N2737), .b(N2546), .O(N3367) );
and2 gate742( .a(N2733), .b(N2542), .O(N3368) );
and2 gate743( .a(N2729), .b(N2538), .O(N3369) );
and2 gate744( .a(N2670), .b(N2458), .O(N3370) );
and2 gate745( .a(N2666), .b(N2454), .O(N3371) );
and2 gate746( .a(N2662), .b(N2450), .O(N3372) );
and2 gate747( .a(N2658), .b(N2446), .O(N3373) );
and2 gate748( .a(N2654), .b(N2442), .O(N3374) );
and2 gate749( .a(N2988), .b(N2650), .O(N3375) );
and2 gate750( .a(N2650), .b(N1966), .O(N3379) );
inv1 gate751( .a(N2781), .O(N3380) );
and2 gate752( .a(N695), .b(N2604), .O(N3381) );
or2 gate753( .a(N3005), .b(N2379), .O(N3384) );
or2 gate754( .a(N3006), .b(N2380), .O(N3390) );
or2 gate755( .a(N3007), .b(N2381), .O(N3398) );
or2 gate756( .a(N3008), .b(N2382), .O(N3404) );
or2 gate757( .a(N3009), .b(N2383), .O(N3410) );
or2 gate758( .a(N3021), .b(N2397), .O(N3416) );
or2 gate759( .a(N3022), .b(N2398), .O(N3420) );
or2 gate760( .a(N3023), .b(N2399), .O(N3424) );
or2 gate761( .a(N3024), .b(N2400), .O(N3428) );
or2 gate762( .a(N3025), .b(N2401), .O(N3432) );
or2 gate763( .a(N3026), .b(N2402), .O(N3436) );
or2 gate764( .a(N3027), .b(N2403), .O(N3440) );
or2 gate765( .a(N3028), .b(N2404), .O(N3444) );
or2 gate766( .a(N3029), .b(N2405), .O(N3448) );
inv1 gate767( .a(N2790), .O(N3452) );
inv1 gate768( .a(N2793), .O(N3453) );
or2 gate769( .a(N3034), .b(N2420), .O(N3454) );
or2 gate770( .a(N3035), .b(N2421), .O(N3458) );
or2 gate771( .a(N3036), .b(N2422), .O(N3462) );
or2 gate772( .a(N3037), .b(N2423), .O(N3466) );
or2 gate773( .a(N3038), .b(N2424), .O(N3470) );
or2 gate774( .a(N3039), .b(N2425), .O(N3474) );
or2 gate775( .a(N3040), .b(N2426), .O(N3478) );
or2 gate776( .a(N3041), .b(N2427), .O(N3482) );
inv1 gate777( .a(N2796), .O(N3486) );
buf1 gate778( .a(N2644), .O(N3487) );
buf1 gate779( .a(N2638), .O(N3490) );
buf1 gate780( .a(N2632), .O(N3493) );
buf1 gate781( .a(N2626), .O(N3496) );
buf1 gate782( .a(N2619), .O(N3499) );
buf1 gate783( .a(N2523), .O(N3502) );

  xor2  gate3766(.a(N2868), .b(N1167), .O(gate784inter0));
  nand2 gate3767(.a(gate784inter0), .b(s_36), .O(gate784inter1));
  and2  gate3768(.a(N2868), .b(N1167), .O(gate784inter2));
  inv1  gate3769(.a(s_36), .O(gate784inter3));
  inv1  gate3770(.a(s_37), .O(gate784inter4));
  nand2 gate3771(.a(gate784inter4), .b(gate784inter3), .O(gate784inter5));
  nor2  gate3772(.a(gate784inter5), .b(gate784inter2), .O(gate784inter6));
  inv1  gate3773(.a(N1167), .O(gate784inter7));
  inv1  gate3774(.a(N2868), .O(gate784inter8));
  nand2 gate3775(.a(gate784inter8), .b(gate784inter7), .O(gate784inter9));
  nand2 gate3776(.a(s_37), .b(gate784inter3), .O(gate784inter10));
  nor2  gate3777(.a(gate784inter10), .b(gate784inter9), .O(gate784inter11));
  nor2  gate3778(.a(gate784inter11), .b(gate784inter6), .O(gate784inter12));
  nand2 gate3779(.a(gate784inter12), .b(gate784inter1), .O(N3507));
buf1 gate785( .a(N2523), .O(N3510) );
nor2 gate786( .a(N644), .b(N2619), .O(N3515) );
buf1 gate787( .a(N2644), .O(N3518) );
buf1 gate788( .a(N2638), .O(N3521) );
buf1 gate789( .a(N2632), .O(N3524) );
buf1 gate790( .a(N2626), .O(N3527) );
buf1 gate791( .a(N2619), .O(N3530) );
buf1 gate792( .a(N2619), .O(N3535) );
buf1 gate793( .a(N2632), .O(N3539) );
buf1 gate794( .a(N2626), .O(N3542) );
buf1 gate795( .a(N2644), .O(N3545) );
buf1 gate796( .a(N2638), .O(N3548) );
inv1 gate797( .a(N2766), .O(N3551) );
inv1 gate798( .a(N2769), .O(N3552) );
buf1 gate799( .a(N2442), .O(N3553) );
buf1 gate800( .a(N2450), .O(N3557) );
buf1 gate801( .a(N2446), .O(N3560) );
buf1 gate802( .a(N2458), .O(N3563) );
buf1 gate803( .a(N2454), .O(N3566) );
inv1 gate804( .a(N2772), .O(N3569) );
inv1 gate805( .a(N2775), .O(N3570) );
buf1 gate806( .a(N2554), .O(N3571) );
buf1 gate807( .a(N2567), .O(N3574) );
buf1 gate808( .a(N2561), .O(N3577) );
buf1 gate809( .a(N2482), .O(N3580) );
buf1 gate810( .a(N2573), .O(N3583) );
buf1 gate811( .a(N2496), .O(N3586) );
buf1 gate812( .a(N2488), .O(N3589) );
buf1 gate813( .a(N2508), .O(N3592) );
buf1 gate814( .a(N2502), .O(N3595) );
buf1 gate815( .a(N2508), .O(N3598) );
buf1 gate816( .a(N2502), .O(N3601) );
buf1 gate817( .a(N2496), .O(N3604) );
buf1 gate818( .a(N2482), .O(N3607) );
buf1 gate819( .a(N2573), .O(N3610) );
buf1 gate820( .a(N2567), .O(N3613) );
buf1 gate821( .a(N2561), .O(N3616) );
buf1 gate822( .a(N2488), .O(N3619) );
buf1 gate823( .a(N2554), .O(N3622) );
nor2 gate824( .a(N734), .b(N2488), .O(N3625) );
nor2 gate825( .a(N708), .b(N2554), .O(N3628) );
buf1 gate826( .a(N2508), .O(N3631) );
buf1 gate827( .a(N2502), .O(N3634) );
buf1 gate828( .a(N2496), .O(N3637) );
buf1 gate829( .a(N2488), .O(N3640) );
buf1 gate830( .a(N2482), .O(N3643) );
buf1 gate831( .a(N2573), .O(N3646) );
buf1 gate832( .a(N2567), .O(N3649) );
buf1 gate833( .a(N2561), .O(N3652) );
buf1 gate834( .a(N2554), .O(N3655) );

  xor2  gate3738(.a(N734), .b(N2488), .O(gate835inter0));
  nand2 gate3739(.a(gate835inter0), .b(s_32), .O(gate835inter1));
  and2  gate3740(.a(N734), .b(N2488), .O(gate835inter2));
  inv1  gate3741(.a(s_32), .O(gate835inter3));
  inv1  gate3742(.a(s_33), .O(gate835inter4));
  nand2 gate3743(.a(gate835inter4), .b(gate835inter3), .O(gate835inter5));
  nor2  gate3744(.a(gate835inter5), .b(gate835inter2), .O(gate835inter6));
  inv1  gate3745(.a(N2488), .O(gate835inter7));
  inv1  gate3746(.a(N734), .O(gate835inter8));
  nand2 gate3747(.a(gate835inter8), .b(gate835inter7), .O(gate835inter9));
  nand2 gate3748(.a(s_33), .b(gate835inter3), .O(gate835inter10));
  nor2  gate3749(.a(gate835inter10), .b(gate835inter9), .O(gate835inter11));
  nor2  gate3750(.a(gate835inter11), .b(gate835inter6), .O(gate835inter12));
  nand2 gate3751(.a(gate835inter12), .b(gate835inter1), .O(N3658));
buf1 gate836( .a(N2674), .O(N3661) );
buf1 gate837( .a(N2674), .O(N3664) );
buf1 gate838( .a(N2761), .O(N3667) );
buf1 gate839( .a(N2478), .O(N3670) );
buf1 gate840( .a(N2757), .O(N3673) );
buf1 gate841( .a(N2474), .O(N3676) );
buf1 gate842( .a(N2753), .O(N3679) );
buf1 gate843( .a(N2470), .O(N3682) );
buf1 gate844( .a(N2745), .O(N3685) );
buf1 gate845( .a(N2462), .O(N3688) );
buf1 gate846( .a(N2741), .O(N3691) );
buf1 gate847( .a(N2550), .O(N3694) );
buf1 gate848( .a(N2737), .O(N3697) );
buf1 gate849( .a(N2546), .O(N3700) );
buf1 gate850( .a(N2733), .O(N3703) );
buf1 gate851( .a(N2542), .O(N3706) );
buf1 gate852( .a(N2749), .O(N3709) );
buf1 gate853( .a(N2466), .O(N3712) );
buf1 gate854( .a(N2729), .O(N3715) );
buf1 gate855( .a(N2538), .O(N3718) );
buf1 gate856( .a(N2704), .O(N3721) );
buf1 gate857( .a(N2700), .O(N3724) );
buf1 gate858( .a(N2696), .O(N3727) );
buf1 gate859( .a(N2688), .O(N3730) );
buf1 gate860( .a(N2692), .O(N3733) );
buf1 gate861( .a(N2670), .O(N3736) );
buf1 gate862( .a(N2458), .O(N3739) );
buf1 gate863( .a(N2666), .O(N3742) );
buf1 gate864( .a(N2454), .O(N3745) );
buf1 gate865( .a(N2662), .O(N3748) );
buf1 gate866( .a(N2450), .O(N3751) );
buf1 gate867( .a(N2658), .O(N3754) );
buf1 gate868( .a(N2446), .O(N3757) );
buf1 gate869( .a(N2654), .O(N3760) );
buf1 gate870( .a(N2442), .O(N3763) );
buf1 gate871( .a(N2654), .O(N3766) );
buf1 gate872( .a(N2662), .O(N3769) );
buf1 gate873( .a(N2658), .O(N3772) );
buf1 gate874( .a(N2670), .O(N3775) );
buf1 gate875( .a(N2666), .O(N3778) );
inv1 gate876( .a(N2784), .O(N3781) );
inv1 gate877( .a(N2787), .O(N3782) );
or2 gate878( .a(N2928), .b(N2326), .O(N3783) );
or2 gate879( .a(N2933), .b(N2342), .O(N3786) );
or2 gate880( .a(N2923), .b(N2321), .O(N3789) );
buf1 gate881( .a(N2688), .O(N3792) );
buf1 gate882( .a(N2696), .O(N3795) );
buf1 gate883( .a(N2692), .O(N3798) );
buf1 gate884( .a(N2704), .O(N3801) );
buf1 gate885( .a(N2700), .O(N3804) );
buf1 gate886( .a(N2604), .O(N3807) );
buf1 gate887( .a(N2611), .O(N3810) );
buf1 gate888( .a(N2607), .O(N3813) );
buf1 gate889( .a(N2615), .O(N3816) );
buf1 gate890( .a(N2538), .O(N3819) );
buf1 gate891( .a(N2546), .O(N3822) );
buf1 gate892( .a(N2542), .O(N3825) );
buf1 gate893( .a(N2462), .O(N3828) );
buf1 gate894( .a(N2550), .O(N3831) );
buf1 gate895( .a(N2470), .O(N3834) );
buf1 gate896( .a(N2466), .O(N3837) );
buf1 gate897( .a(N2478), .O(N3840) );
buf1 gate898( .a(N2474), .O(N3843) );
buf1 gate899( .a(N2615), .O(N3846) );
buf1 gate900( .a(N2611), .O(N3849) );
buf1 gate901( .a(N2607), .O(N3852) );
buf1 gate902( .a(N2680), .O(N3855) );
buf1 gate903( .a(N2729), .O(N3858) );
buf1 gate904( .a(N2737), .O(N3861) );
buf1 gate905( .a(N2733), .O(N3864) );
buf1 gate906( .a(N2745), .O(N3867) );
buf1 gate907( .a(N2741), .O(N3870) );
buf1 gate908( .a(N2753), .O(N3873) );
buf1 gate909( .a(N2749), .O(N3876) );
buf1 gate910( .a(N2761), .O(N3879) );
buf1 gate911( .a(N2757), .O(N3882) );
or2 gate912( .a(N3033), .b(N2419), .O(N3885) );
or2 gate913( .a(N3032), .b(N2418), .O(N3888) );
or2 gate914( .a(N3020), .b(N2396), .O(N3891) );
nand2 gate915( .a(N3067), .b(N2117), .O(N3953) );
inv1 gate916( .a(N3067), .O(N3954) );

  xor2  gate4102(.a(N2537), .b(N3070), .O(gate917inter0));
  nand2 gate4103(.a(gate917inter0), .b(s_84), .O(gate917inter1));
  and2  gate4104(.a(N2537), .b(N3070), .O(gate917inter2));
  inv1  gate4105(.a(s_84), .O(gate917inter3));
  inv1  gate4106(.a(s_85), .O(gate917inter4));
  nand2 gate4107(.a(gate917inter4), .b(gate917inter3), .O(gate917inter5));
  nor2  gate4108(.a(gate917inter5), .b(gate917inter2), .O(gate917inter6));
  inv1  gate4109(.a(N3070), .O(gate917inter7));
  inv1  gate4110(.a(N2537), .O(gate917inter8));
  nand2 gate4111(.a(gate917inter8), .b(gate917inter7), .O(gate917inter9));
  nand2 gate4112(.a(s_85), .b(gate917inter3), .O(gate917inter10));
  nor2  gate4113(.a(gate917inter10), .b(gate917inter9), .O(gate917inter11));
  nor2  gate4114(.a(gate917inter11), .b(gate917inter6), .O(gate917inter12));
  nand2 gate4115(.a(gate917inter12), .b(gate917inter1), .O(N3955));
inv1 gate918( .a(N3070), .O(N3956) );
inv1 gate919( .a(N3073), .O(N3958) );
inv1 gate920( .a(N3080), .O(N3964) );
or2 gate921( .a(N1649), .b(N3379), .O(N4193) );
or3 gate922( .a(N1167), .b(N2867), .c(N3130), .O(N4303) );
inv1 gate923( .a(N3061), .O(N4308) );
inv1 gate924( .a(N3064), .O(N4313) );
nand2 gate925( .a(N2769), .b(N3551), .O(N4326) );
nand2 gate926( .a(N2766), .b(N3552), .O(N4327) );
nand2 gate927( .a(N2775), .b(N3569), .O(N4333) );
nand2 gate928( .a(N2772), .b(N3570), .O(N4334) );
nand2 gate929( .a(N2787), .b(N3781), .O(N4411) );
nand2 gate930( .a(N2784), .b(N3782), .O(N4412) );
nand2 gate931( .a(N3487), .b(N1828), .O(N4463) );
inv1 gate932( .a(N3487), .O(N4464) );
nand2 gate933( .a(N3490), .b(N1829), .O(N4465) );
inv1 gate934( .a(N3490), .O(N4466) );

  xor2  gate5138(.a(N2267), .b(N3493), .O(gate935inter0));
  nand2 gate5139(.a(gate935inter0), .b(s_232), .O(gate935inter1));
  and2  gate5140(.a(N2267), .b(N3493), .O(gate935inter2));
  inv1  gate5141(.a(s_232), .O(gate935inter3));
  inv1  gate5142(.a(s_233), .O(gate935inter4));
  nand2 gate5143(.a(gate935inter4), .b(gate935inter3), .O(gate935inter5));
  nor2  gate5144(.a(gate935inter5), .b(gate935inter2), .O(gate935inter6));
  inv1  gate5145(.a(N3493), .O(gate935inter7));
  inv1  gate5146(.a(N2267), .O(gate935inter8));
  nand2 gate5147(.a(gate935inter8), .b(gate935inter7), .O(gate935inter9));
  nand2 gate5148(.a(s_233), .b(gate935inter3), .O(gate935inter10));
  nor2  gate5149(.a(gate935inter10), .b(gate935inter9), .O(gate935inter11));
  nor2  gate5150(.a(gate935inter11), .b(gate935inter6), .O(gate935inter12));
  nand2 gate5151(.a(gate935inter12), .b(gate935inter1), .O(N4467));
inv1 gate936( .a(N3493), .O(N4468) );
nand2 gate937( .a(N3496), .b(N1830), .O(N4469) );
inv1 gate938( .a(N3496), .O(N4470) );
nand2 gate939( .a(N3499), .b(N1833), .O(N4471) );
inv1 gate940( .a(N3499), .O(N4472) );
inv1 gate941( .a(N3122), .O(N4473) );
inv1 gate942( .a(N3126), .O(N4474) );
nand2 gate943( .a(N3518), .b(N1840), .O(N4475) );
inv1 gate944( .a(N3518), .O(N4476) );
nand2 gate945( .a(N3521), .b(N1841), .O(N4477) );
inv1 gate946( .a(N3521), .O(N4478) );
nand2 gate947( .a(N3524), .b(N2275), .O(N4479) );
inv1 gate948( .a(N3524), .O(N4480) );
nand2 gate949( .a(N3527), .b(N1842), .O(N4481) );
inv1 gate950( .a(N3527), .O(N4482) );
nand2 gate951( .a(N3530), .b(N1843), .O(N4483) );
inv1 gate952( .a(N3530), .O(N4484) );
inv1 gate953( .a(N3155), .O(N4485) );
inv1 gate954( .a(N3159), .O(N4486) );
nand2 gate955( .a(N1721), .b(N3954), .O(N4487) );
nand2 gate956( .a(N2235), .b(N3956), .O(N4488) );
inv1 gate957( .a(N3535), .O(N4489) );

  xor2  gate3682(.a(N3958), .b(N3535), .O(gate958inter0));
  nand2 gate3683(.a(gate958inter0), .b(s_24), .O(gate958inter1));
  and2  gate3684(.a(N3958), .b(N3535), .O(gate958inter2));
  inv1  gate3685(.a(s_24), .O(gate958inter3));
  inv1  gate3686(.a(s_25), .O(gate958inter4));
  nand2 gate3687(.a(gate958inter4), .b(gate958inter3), .O(gate958inter5));
  nor2  gate3688(.a(gate958inter5), .b(gate958inter2), .O(gate958inter6));
  inv1  gate3689(.a(N3535), .O(gate958inter7));
  inv1  gate3690(.a(N3958), .O(gate958inter8));
  nand2 gate3691(.a(gate958inter8), .b(gate958inter7), .O(gate958inter9));
  nand2 gate3692(.a(s_25), .b(gate958inter3), .O(gate958inter10));
  nor2  gate3693(.a(gate958inter10), .b(gate958inter9), .O(gate958inter11));
  nor2  gate3694(.a(gate958inter11), .b(gate958inter6), .O(gate958inter12));
  nand2 gate3695(.a(gate958inter12), .b(gate958inter1), .O(N4490));
inv1 gate959( .a(N3539), .O(N4491) );
inv1 gate960( .a(N3542), .O(N4492) );
inv1 gate961( .a(N3545), .O(N4493) );
inv1 gate962( .a(N3548), .O(N4494) );
inv1 gate963( .a(N3553), .O(N4495) );
nand2 gate964( .a(N3553), .b(N3964), .O(N4496) );
inv1 gate965( .a(N3557), .O(N4497) );
inv1 gate966( .a(N3560), .O(N4498) );
inv1 gate967( .a(N3563), .O(N4499) );
inv1 gate968( .a(N3566), .O(N4500) );
inv1 gate969( .a(N3571), .O(N4501) );
nand2 gate970( .a(N3571), .b(N3167), .O(N4502) );
inv1 gate971( .a(N3574), .O(N4503) );
inv1 gate972( .a(N3577), .O(N4504) );
inv1 gate973( .a(N3580), .O(N4505) );
inv1 gate974( .a(N3583), .O(N4506) );
nand2 gate975( .a(N3598), .b(N1867), .O(N4507) );
inv1 gate976( .a(N3598), .O(N4508) );
nand2 gate977( .a(N3601), .b(N1868), .O(N4509) );
inv1 gate978( .a(N3601), .O(N4510) );
nand2 gate979( .a(N3604), .b(N1869), .O(N4511) );
inv1 gate980( .a(N3604), .O(N4512) );
nand2 gate981( .a(N3607), .b(N1870), .O(N4513) );
inv1 gate982( .a(N3607), .O(N4514) );
nand2 gate983( .a(N3610), .b(N1871), .O(N4515) );
inv1 gate984( .a(N3610), .O(N4516) );
nand2 gate985( .a(N3613), .b(N1872), .O(N4517) );
inv1 gate986( .a(N3613), .O(N4518) );
nand2 gate987( .a(N3616), .b(N1873), .O(N4519) );
inv1 gate988( .a(N3616), .O(N4520) );
nand2 gate989( .a(N3619), .b(N1874), .O(N4521) );
inv1 gate990( .a(N3619), .O(N4522) );
nand2 gate991( .a(N3622), .b(N1875), .O(N4523) );
inv1 gate992( .a(N3622), .O(N4524) );
nand2 gate993( .a(N3631), .b(N1876), .O(N4525) );
inv1 gate994( .a(N3631), .O(N4526) );
nand2 gate995( .a(N3634), .b(N1877), .O(N4527) );
inv1 gate996( .a(N3634), .O(N4528) );
nand2 gate997( .a(N3637), .b(N1878), .O(N4529) );
inv1 gate998( .a(N3637), .O(N4530) );
nand2 gate999( .a(N3640), .b(N1879), .O(N4531) );
inv1 gate1000( .a(N3640), .O(N4532) );
nand2 gate1001( .a(N3643), .b(N1880), .O(N4533) );
inv1 gate1002( .a(N3643), .O(N4534) );

  xor2  gate3836(.a(N1881), .b(N3646), .O(gate1003inter0));
  nand2 gate3837(.a(gate1003inter0), .b(s_46), .O(gate1003inter1));
  and2  gate3838(.a(N1881), .b(N3646), .O(gate1003inter2));
  inv1  gate3839(.a(s_46), .O(gate1003inter3));
  inv1  gate3840(.a(s_47), .O(gate1003inter4));
  nand2 gate3841(.a(gate1003inter4), .b(gate1003inter3), .O(gate1003inter5));
  nor2  gate3842(.a(gate1003inter5), .b(gate1003inter2), .O(gate1003inter6));
  inv1  gate3843(.a(N3646), .O(gate1003inter7));
  inv1  gate3844(.a(N1881), .O(gate1003inter8));
  nand2 gate3845(.a(gate1003inter8), .b(gate1003inter7), .O(gate1003inter9));
  nand2 gate3846(.a(s_47), .b(gate1003inter3), .O(gate1003inter10));
  nor2  gate3847(.a(gate1003inter10), .b(gate1003inter9), .O(gate1003inter11));
  nor2  gate3848(.a(gate1003inter11), .b(gate1003inter6), .O(gate1003inter12));
  nand2 gate3849(.a(gate1003inter12), .b(gate1003inter1), .O(N4535));
inv1 gate1004( .a(N3646), .O(N4536) );
nand2 gate1005( .a(N3649), .b(N1882), .O(N4537) );
inv1 gate1006( .a(N3649), .O(N4538) );
nand2 gate1007( .a(N3652), .b(N1883), .O(N4539) );
inv1 gate1008( .a(N3652), .O(N4540) );
nand2 gate1009( .a(N3655), .b(N1884), .O(N4541) );
inv1 gate1010( .a(N3655), .O(N4542) );
inv1 gate1011( .a(N3658), .O(N4543) );
and2 gate1012( .a(N806), .b(N3293), .O(N4544) );
and2 gate1013( .a(N800), .b(N3287), .O(N4545) );
and2 gate1014( .a(N794), .b(N3281), .O(N4549) );
and2 gate1015( .a(N3273), .b(N786), .O(N4555) );
and2 gate1016( .a(N780), .b(N3267), .O(N4562) );
and2 gate1017( .a(N774), .b(N3355), .O(N4563) );
and2 gate1018( .a(N768), .b(N3349), .O(N4566) );
and2 gate1019( .a(N762), .b(N3343), .O(N4570) );
inv1 gate1020( .a(N3661), .O(N4575) );
and2 gate1021( .a(N806), .b(N3293), .O(N4576) );
and2 gate1022( .a(N800), .b(N3287), .O(N4577) );
and2 gate1023( .a(N794), .b(N3281), .O(N4581) );
and2 gate1024( .a(N786), .b(N3273), .O(N4586) );
and2 gate1025( .a(N780), .b(N3267), .O(N4592) );
and2 gate1026( .a(N774), .b(N3355), .O(N4593) );
and2 gate1027( .a(N768), .b(N3349), .O(N4597) );
and2 gate1028( .a(N762), .b(N3343), .O(N4603) );
inv1 gate1029( .a(N3664), .O(N4610) );
inv1 gate1030( .a(N3667), .O(N4611) );
inv1 gate1031( .a(N3670), .O(N4612) );
inv1 gate1032( .a(N3673), .O(N4613) );
inv1 gate1033( .a(N3676), .O(N4614) );
inv1 gate1034( .a(N3679), .O(N4615) );
inv1 gate1035( .a(N3682), .O(N4616) );
inv1 gate1036( .a(N3685), .O(N4617) );
inv1 gate1037( .a(N3688), .O(N4618) );
inv1 gate1038( .a(N3691), .O(N4619) );
inv1 gate1039( .a(N3694), .O(N4620) );
inv1 gate1040( .a(N3697), .O(N4621) );
inv1 gate1041( .a(N3700), .O(N4622) );
inv1 gate1042( .a(N3703), .O(N4623) );
inv1 gate1043( .a(N3706), .O(N4624) );
inv1 gate1044( .a(N3709), .O(N4625) );
inv1 gate1045( .a(N3712), .O(N4626) );
inv1 gate1046( .a(N3715), .O(N4627) );
inv1 gate1047( .a(N3718), .O(N4628) );
inv1 gate1048( .a(N3721), .O(N4629) );
and2 gate1049( .a(N3448), .b(N2704), .O(N4630) );
inv1 gate1050( .a(N3724), .O(N4631) );
and2 gate1051( .a(N3444), .b(N2700), .O(N4632) );
inv1 gate1052( .a(N3727), .O(N4633) );
and2 gate1053( .a(N3440), .b(N2696), .O(N4634) );
and2 gate1054( .a(N3436), .b(N2692), .O(N4635) );
inv1 gate1055( .a(N3730), .O(N4636) );
and2 gate1056( .a(N3432), .b(N2688), .O(N4637) );
and2 gate1057( .a(N3428), .b(N3311), .O(N4638) );
and2 gate1058( .a(N3424), .b(N3307), .O(N4639) );
and2 gate1059( .a(N3420), .b(N3303), .O(N4640) );
and2 gate1060( .a(N3416), .b(N3299), .O(N4641) );
inv1 gate1061( .a(N3733), .O(N4642) );
inv1 gate1062( .a(N3736), .O(N4643) );
inv1 gate1063( .a(N3739), .O(N4644) );
inv1 gate1064( .a(N3742), .O(N4645) );
inv1 gate1065( .a(N3745), .O(N4646) );
inv1 gate1066( .a(N3748), .O(N4647) );
inv1 gate1067( .a(N3751), .O(N4648) );
inv1 gate1068( .a(N3754), .O(N4649) );
inv1 gate1069( .a(N3757), .O(N4650) );
inv1 gate1070( .a(N3760), .O(N4651) );
inv1 gate1071( .a(N3763), .O(N4652) );
inv1 gate1072( .a(N3375), .O(N4653) );
and2 gate1073( .a(N865), .b(N3410), .O(N4656) );
and2 gate1074( .a(N859), .b(N3404), .O(N4657) );
and2 gate1075( .a(N853), .b(N3398), .O(N4661) );
and2 gate1076( .a(N3390), .b(N845), .O(N4667) );
and2 gate1077( .a(N839), .b(N3384), .O(N4674) );
and2 gate1078( .a(N833), .b(N3334), .O(N4675) );
and2 gate1079( .a(N827), .b(N3328), .O(N4678) );
and2 gate1080( .a(N821), .b(N3322), .O(N4682) );
and2 gate1081( .a(N814), .b(N3315), .O(N4687) );
inv1 gate1082( .a(N3766), .O(N4693) );
nand2 gate1083( .a(N3766), .b(N3380), .O(N4694) );
inv1 gate1084( .a(N3769), .O(N4695) );
inv1 gate1085( .a(N3772), .O(N4696) );
inv1 gate1086( .a(N3775), .O(N4697) );
inv1 gate1087( .a(N3778), .O(N4698) );
inv1 gate1088( .a(N3783), .O(N4699) );
inv1 gate1089( .a(N3786), .O(N4700) );
and2 gate1090( .a(N865), .b(N3410), .O(N4701) );
and2 gate1091( .a(N859), .b(N3404), .O(N4702) );
and2 gate1092( .a(N853), .b(N3398), .O(N4706) );
and2 gate1093( .a(N845), .b(N3390), .O(N4711) );
and2 gate1094( .a(N839), .b(N3384), .O(N4717) );
and2 gate1095( .a(N833), .b(N3334), .O(N4718) );
and2 gate1096( .a(N827), .b(N3328), .O(N4722) );
and2 gate1097( .a(N821), .b(N3322), .O(N4728) );
and2 gate1098( .a(N814), .b(N3315), .O(N4735) );
inv1 gate1099( .a(N3789), .O(N4743) );
inv1 gate1100( .a(N3792), .O(N4744) );
inv1 gate1101( .a(N3807), .O(N4745) );

  xor2  gate4746(.a(N3452), .b(N3807), .O(gate1102inter0));
  nand2 gate4747(.a(gate1102inter0), .b(s_176), .O(gate1102inter1));
  and2  gate4748(.a(N3452), .b(N3807), .O(gate1102inter2));
  inv1  gate4749(.a(s_176), .O(gate1102inter3));
  inv1  gate4750(.a(s_177), .O(gate1102inter4));
  nand2 gate4751(.a(gate1102inter4), .b(gate1102inter3), .O(gate1102inter5));
  nor2  gate4752(.a(gate1102inter5), .b(gate1102inter2), .O(gate1102inter6));
  inv1  gate4753(.a(N3807), .O(gate1102inter7));
  inv1  gate4754(.a(N3452), .O(gate1102inter8));
  nand2 gate4755(.a(gate1102inter8), .b(gate1102inter7), .O(gate1102inter9));
  nand2 gate4756(.a(s_177), .b(gate1102inter3), .O(gate1102inter10));
  nor2  gate4757(.a(gate1102inter10), .b(gate1102inter9), .O(gate1102inter11));
  nor2  gate4758(.a(gate1102inter11), .b(gate1102inter6), .O(gate1102inter12));
  nand2 gate4759(.a(gate1102inter12), .b(gate1102inter1), .O(N4746));
inv1 gate1103( .a(N3810), .O(N4747) );
inv1 gate1104( .a(N3813), .O(N4748) );
inv1 gate1105( .a(N3816), .O(N4749) );
inv1 gate1106( .a(N3819), .O(N4750) );
nand2 gate1107( .a(N3819), .b(N3453), .O(N4751) );
inv1 gate1108( .a(N3822), .O(N4752) );
inv1 gate1109( .a(N3825), .O(N4753) );
inv1 gate1110( .a(N3828), .O(N4754) );
inv1 gate1111( .a(N3831), .O(N4755) );
and2 gate1112( .a(N3482), .b(N3263), .O(N4756) );
and2 gate1113( .a(N3478), .b(N3259), .O(N4757) );
and2 gate1114( .a(N3474), .b(N3255), .O(N4758) );
and2 gate1115( .a(N3470), .b(N3251), .O(N4759) );
and2 gate1116( .a(N3466), .b(N3247), .O(N4760) );
inv1 gate1117( .a(N3846), .O(N4761) );
and2 gate1118( .a(N3462), .b(N2615), .O(N4762) );
inv1 gate1119( .a(N3849), .O(N4763) );
and2 gate1120( .a(N3458), .b(N2611), .O(N4764) );
inv1 gate1121( .a(N3852), .O(N4765) );
and2 gate1122( .a(N3454), .b(N2607), .O(N4766) );
and2 gate1123( .a(N2680), .b(N3381), .O(N4767) );
inv1 gate1124( .a(N3855), .O(N4768) );
and2 gate1125( .a(N3340), .b(N695), .O(N4769) );
inv1 gate1126( .a(N3858), .O(N4775) );
nand2 gate1127( .a(N3858), .b(N3486), .O(N4776) );
inv1 gate1128( .a(N3861), .O(N4777) );
inv1 gate1129( .a(N3864), .O(N4778) );
inv1 gate1130( .a(N3867), .O(N4779) );
inv1 gate1131( .a(N3870), .O(N4780) );
inv1 gate1132( .a(N3885), .O(N4781) );
inv1 gate1133( .a(N3888), .O(N4782) );
inv1 gate1134( .a(N3891), .O(N4783) );
or2 gate1135( .a(N3131), .b(N3134), .O(N4784) );
inv1 gate1136( .a(N3502), .O(N4789) );
inv1 gate1137( .a(N3131), .O(N4790) );
inv1 gate1138( .a(N3507), .O(N4793) );
inv1 gate1139( .a(N3510), .O(N4794) );
inv1 gate1140( .a(N3515), .O(N4795) );
buf1 gate1141( .a(N3114), .O(N4796) );
inv1 gate1142( .a(N3586), .O(N4799) );
inv1 gate1143( .a(N3589), .O(N4800) );
inv1 gate1144( .a(N3592), .O(N4801) );
inv1 gate1145( .a(N3595), .O(N4802) );
nand2 gate1146( .a(N4326), .b(N4327), .O(N4803) );

  xor2  gate4326(.a(N4334), .b(N4333), .O(gate1147inter0));
  nand2 gate4327(.a(gate1147inter0), .b(s_116), .O(gate1147inter1));
  and2  gate4328(.a(N4334), .b(N4333), .O(gate1147inter2));
  inv1  gate4329(.a(s_116), .O(gate1147inter3));
  inv1  gate4330(.a(s_117), .O(gate1147inter4));
  nand2 gate4331(.a(gate1147inter4), .b(gate1147inter3), .O(gate1147inter5));
  nor2  gate4332(.a(gate1147inter5), .b(gate1147inter2), .O(gate1147inter6));
  inv1  gate4333(.a(N4333), .O(gate1147inter7));
  inv1  gate4334(.a(N4334), .O(gate1147inter8));
  nand2 gate4335(.a(gate1147inter8), .b(gate1147inter7), .O(gate1147inter9));
  nand2 gate4336(.a(s_117), .b(gate1147inter3), .O(gate1147inter10));
  nor2  gate4337(.a(gate1147inter10), .b(gate1147inter9), .O(gate1147inter11));
  nor2  gate4338(.a(gate1147inter11), .b(gate1147inter6), .O(gate1147inter12));
  nand2 gate4339(.a(gate1147inter12), .b(gate1147inter1), .O(N4806));
inv1 gate1148( .a(N3625), .O(N4809) );
buf1 gate1149( .a(N3178), .O(N4810) );
inv1 gate1150( .a(N3628), .O(N4813) );
buf1 gate1151( .a(N3202), .O(N4814) );
buf1 gate1152( .a(N3221), .O(N4817) );
buf1 gate1153( .a(N3293), .O(N4820) );
buf1 gate1154( .a(N3287), .O(N4823) );
buf1 gate1155( .a(N3281), .O(N4826) );
buf1 gate1156( .a(N3273), .O(N4829) );
buf1 gate1157( .a(N3267), .O(N4832) );
buf1 gate1158( .a(N3355), .O(N4835) );
buf1 gate1159( .a(N3349), .O(N4838) );
buf1 gate1160( .a(N3343), .O(N4841) );
nor2 gate1161( .a(N3273), .b(N786), .O(N4844) );
buf1 gate1162( .a(N3293), .O(N4847) );
buf1 gate1163( .a(N3287), .O(N4850) );
buf1 gate1164( .a(N3281), .O(N4853) );
buf1 gate1165( .a(N3267), .O(N4856) );
buf1 gate1166( .a(N3355), .O(N4859) );
buf1 gate1167( .a(N3349), .O(N4862) );
buf1 gate1168( .a(N3343), .O(N4865) );
buf1 gate1169( .a(N3273), .O(N4868) );
nor2 gate1170( .a(N786), .b(N3273), .O(N4871) );
buf1 gate1171( .a(N3448), .O(N4874) );
buf1 gate1172( .a(N3444), .O(N4877) );
buf1 gate1173( .a(N3440), .O(N4880) );
buf1 gate1174( .a(N3432), .O(N4883) );
buf1 gate1175( .a(N3428), .O(N4886) );
buf1 gate1176( .a(N3311), .O(N4889) );
buf1 gate1177( .a(N3424), .O(N4892) );
buf1 gate1178( .a(N3307), .O(N4895) );
buf1 gate1179( .a(N3420), .O(N4898) );
buf1 gate1180( .a(N3303), .O(N4901) );
buf1 gate1181( .a(N3436), .O(N4904) );
buf1 gate1182( .a(N3416), .O(N4907) );
buf1 gate1183( .a(N3299), .O(N4910) );
buf1 gate1184( .a(N3410), .O(N4913) );
buf1 gate1185( .a(N3404), .O(N4916) );
buf1 gate1186( .a(N3398), .O(N4919) );
buf1 gate1187( .a(N3390), .O(N4922) );
buf1 gate1188( .a(N3384), .O(N4925) );
buf1 gate1189( .a(N3334), .O(N4928) );
buf1 gate1190( .a(N3328), .O(N4931) );
buf1 gate1191( .a(N3322), .O(N4934) );
buf1 gate1192( .a(N3315), .O(N4937) );
nor2 gate1193( .a(N3390), .b(N845), .O(N4940) );
buf1 gate1194( .a(N3315), .O(N4943) );
buf1 gate1195( .a(N3328), .O(N4946) );
buf1 gate1196( .a(N3322), .O(N4949) );
buf1 gate1197( .a(N3384), .O(N4952) );
buf1 gate1198( .a(N3334), .O(N4955) );
buf1 gate1199( .a(N3398), .O(N4958) );
buf1 gate1200( .a(N3390), .O(N4961) );
buf1 gate1201( .a(N3410), .O(N4964) );
buf1 gate1202( .a(N3404), .O(N4967) );
buf1 gate1203( .a(N3340), .O(N4970) );
buf1 gate1204( .a(N3349), .O(N4973) );
buf1 gate1205( .a(N3343), .O(N4976) );
buf1 gate1206( .a(N3267), .O(N4979) );
buf1 gate1207( .a(N3355), .O(N4982) );
buf1 gate1208( .a(N3281), .O(N4985) );
buf1 gate1209( .a(N3273), .O(N4988) );
buf1 gate1210( .a(N3293), .O(N4991) );
buf1 gate1211( .a(N3287), .O(N4994) );
nand2 gate1212( .a(N4411), .b(N4412), .O(N4997) );
buf1 gate1213( .a(N3410), .O(N5000) );
buf1 gate1214( .a(N3404), .O(N5003) );
buf1 gate1215( .a(N3398), .O(N5006) );
buf1 gate1216( .a(N3384), .O(N5009) );
buf1 gate1217( .a(N3334), .O(N5012) );
buf1 gate1218( .a(N3328), .O(N5015) );
buf1 gate1219( .a(N3322), .O(N5018) );
buf1 gate1220( .a(N3390), .O(N5021) );
buf1 gate1221( .a(N3315), .O(N5024) );
nor2 gate1222( .a(N845), .b(N3390), .O(N5027) );
nor2 gate1223( .a(N814), .b(N3315), .O(N5030) );
buf1 gate1224( .a(N3299), .O(N5033) );
buf1 gate1225( .a(N3307), .O(N5036) );
buf1 gate1226( .a(N3303), .O(N5039) );
buf1 gate1227( .a(N3311), .O(N5042) );
inv1 gate1228( .a(N3795), .O(N5045) );
inv1 gate1229( .a(N3798), .O(N5046) );
inv1 gate1230( .a(N3801), .O(N5047) );
inv1 gate1231( .a(N3804), .O(N5048) );
buf1 gate1232( .a(N3247), .O(N5049) );
buf1 gate1233( .a(N3255), .O(N5052) );
buf1 gate1234( .a(N3251), .O(N5055) );
buf1 gate1235( .a(N3263), .O(N5058) );
buf1 gate1236( .a(N3259), .O(N5061) );
inv1 gate1237( .a(N3834), .O(N5064) );
inv1 gate1238( .a(N3837), .O(N5065) );
inv1 gate1239( .a(N3840), .O(N5066) );
inv1 gate1240( .a(N3843), .O(N5067) );
buf1 gate1241( .a(N3482), .O(N5068) );
buf1 gate1242( .a(N3263), .O(N5071) );
buf1 gate1243( .a(N3478), .O(N5074) );
buf1 gate1244( .a(N3259), .O(N5077) );
buf1 gate1245( .a(N3474), .O(N5080) );
buf1 gate1246( .a(N3255), .O(N5083) );
buf1 gate1247( .a(N3466), .O(N5086) );
buf1 gate1248( .a(N3247), .O(N5089) );
buf1 gate1249( .a(N3462), .O(N5092) );
buf1 gate1250( .a(N3458), .O(N5095) );
buf1 gate1251( .a(N3454), .O(N5098) );
buf1 gate1252( .a(N3470), .O(N5101) );
buf1 gate1253( .a(N3251), .O(N5104) );
buf1 gate1254( .a(N3381), .O(N5107) );
inv1 gate1255( .a(N3873), .O(N5110) );
inv1 gate1256( .a(N3876), .O(N5111) );
inv1 gate1257( .a(N3879), .O(N5112) );
inv1 gate1258( .a(N3882), .O(N5113) );
buf1 gate1259( .a(N3458), .O(N5114) );
buf1 gate1260( .a(N3454), .O(N5117) );
buf1 gate1261( .a(N3466), .O(N5120) );
buf1 gate1262( .a(N3462), .O(N5123) );
buf1 gate1263( .a(N3474), .O(N5126) );
buf1 gate1264( .a(N3470), .O(N5129) );
buf1 gate1265( .a(N3482), .O(N5132) );
buf1 gate1266( .a(N3478), .O(N5135) );
buf1 gate1267( .a(N3416), .O(N5138) );
buf1 gate1268( .a(N3424), .O(N5141) );
buf1 gate1269( .a(N3420), .O(N5144) );
buf1 gate1270( .a(N3432), .O(N5147) );
buf1 gate1271( .a(N3428), .O(N5150) );
buf1 gate1272( .a(N3440), .O(N5153) );
buf1 gate1273( .a(N3436), .O(N5156) );
buf1 gate1274( .a(N3448), .O(N5159) );
buf1 gate1275( .a(N3444), .O(N5162) );
nand2 gate1276( .a(N4486), .b(N4485), .O(N5165) );
nand2 gate1277( .a(N4474), .b(N4473), .O(N5166) );
nand2 gate1278( .a(N1290), .b(N4464), .O(N5167) );
nand2 gate1279( .a(N1293), .b(N4466), .O(N5168) );
nand2 gate1280( .a(N2074), .b(N4468), .O(N5169) );
nand2 gate1281( .a(N1296), .b(N4470), .O(N5170) );
nand2 gate1282( .a(N1302), .b(N4472), .O(N5171) );
nand2 gate1283( .a(N1314), .b(N4476), .O(N5172) );
nand2 gate1284( .a(N1317), .b(N4478), .O(N5173) );
nand2 gate1285( .a(N2081), .b(N4480), .O(N5174) );

  xor2  gate5152(.a(N4482), .b(N1320), .O(gate1286inter0));
  nand2 gate5153(.a(gate1286inter0), .b(s_234), .O(gate1286inter1));
  and2  gate5154(.a(N4482), .b(N1320), .O(gate1286inter2));
  inv1  gate5155(.a(s_234), .O(gate1286inter3));
  inv1  gate5156(.a(s_235), .O(gate1286inter4));
  nand2 gate5157(.a(gate1286inter4), .b(gate1286inter3), .O(gate1286inter5));
  nor2  gate5158(.a(gate1286inter5), .b(gate1286inter2), .O(gate1286inter6));
  inv1  gate5159(.a(N1320), .O(gate1286inter7));
  inv1  gate5160(.a(N4482), .O(gate1286inter8));
  nand2 gate5161(.a(gate1286inter8), .b(gate1286inter7), .O(gate1286inter9));
  nand2 gate5162(.a(s_235), .b(gate1286inter3), .O(gate1286inter10));
  nor2  gate5163(.a(gate1286inter10), .b(gate1286inter9), .O(gate1286inter11));
  nor2  gate5164(.a(gate1286inter11), .b(gate1286inter6), .O(gate1286inter12));
  nand2 gate5165(.a(gate1286inter12), .b(gate1286inter1), .O(N5175));
nand2 gate1287( .a(N1323), .b(N4484), .O(N5176) );
nand2 gate1288( .a(N3953), .b(N4487), .O(N5177) );

  xor2  gate5026(.a(N4488), .b(N3955), .O(gate1289inter0));
  nand2 gate5027(.a(gate1289inter0), .b(s_216), .O(gate1289inter1));
  and2  gate5028(.a(N4488), .b(N3955), .O(gate1289inter2));
  inv1  gate5029(.a(s_216), .O(gate1289inter3));
  inv1  gate5030(.a(s_217), .O(gate1289inter4));
  nand2 gate5031(.a(gate1289inter4), .b(gate1289inter3), .O(gate1289inter5));
  nor2  gate5032(.a(gate1289inter5), .b(gate1289inter2), .O(gate1289inter6));
  inv1  gate5033(.a(N3955), .O(gate1289inter7));
  inv1  gate5034(.a(N4488), .O(gate1289inter8));
  nand2 gate5035(.a(gate1289inter8), .b(gate1289inter7), .O(gate1289inter9));
  nand2 gate5036(.a(s_217), .b(gate1289inter3), .O(gate1289inter10));
  nor2  gate5037(.a(gate1289inter10), .b(gate1289inter9), .O(gate1289inter11));
  nor2  gate5038(.a(gate1289inter11), .b(gate1289inter6), .O(gate1289inter12));
  nand2 gate5039(.a(gate1289inter12), .b(gate1289inter1), .O(N5178));
nand2 gate1290( .a(N3073), .b(N4489), .O(N5179) );
nand2 gate1291( .a(N3542), .b(N4491), .O(N5180) );
nand2 gate1292( .a(N3539), .b(N4492), .O(N5181) );
nand2 gate1293( .a(N3548), .b(N4493), .O(N5182) );
nand2 gate1294( .a(N3545), .b(N4494), .O(N5183) );
nand2 gate1295( .a(N3080), .b(N4495), .O(N5184) );
nand2 gate1296( .a(N3560), .b(N4497), .O(N5185) );
nand2 gate1297( .a(N3557), .b(N4498), .O(N5186) );
nand2 gate1298( .a(N3566), .b(N4499), .O(N5187) );
nand2 gate1299( .a(N3563), .b(N4500), .O(N5188) );
nand2 gate1300( .a(N2778), .b(N4501), .O(N5189) );
nand2 gate1301( .a(N3577), .b(N4503), .O(N5190) );
nand2 gate1302( .a(N3574), .b(N4504), .O(N5191) );
nand2 gate1303( .a(N3583), .b(N4505), .O(N5192) );
nand2 gate1304( .a(N3580), .b(N4506), .O(N5193) );
nand2 gate1305( .a(N1326), .b(N4508), .O(N5196) );
nand2 gate1306( .a(N1329), .b(N4510), .O(N5197) );
nand2 gate1307( .a(N1332), .b(N4512), .O(N5198) );
nand2 gate1308( .a(N1335), .b(N4514), .O(N5199) );
nand2 gate1309( .a(N1338), .b(N4516), .O(N5200) );
nand2 gate1310( .a(N1341), .b(N4518), .O(N5201) );
nand2 gate1311( .a(N1344), .b(N4520), .O(N5202) );

  xor2  gate4116(.a(N4522), .b(N1347), .O(gate1312inter0));
  nand2 gate4117(.a(gate1312inter0), .b(s_86), .O(gate1312inter1));
  and2  gate4118(.a(N4522), .b(N1347), .O(gate1312inter2));
  inv1  gate4119(.a(s_86), .O(gate1312inter3));
  inv1  gate4120(.a(s_87), .O(gate1312inter4));
  nand2 gate4121(.a(gate1312inter4), .b(gate1312inter3), .O(gate1312inter5));
  nor2  gate4122(.a(gate1312inter5), .b(gate1312inter2), .O(gate1312inter6));
  inv1  gate4123(.a(N1347), .O(gate1312inter7));
  inv1  gate4124(.a(N4522), .O(gate1312inter8));
  nand2 gate4125(.a(gate1312inter8), .b(gate1312inter7), .O(gate1312inter9));
  nand2 gate4126(.a(s_87), .b(gate1312inter3), .O(gate1312inter10));
  nor2  gate4127(.a(gate1312inter10), .b(gate1312inter9), .O(gate1312inter11));
  nor2  gate4128(.a(gate1312inter11), .b(gate1312inter6), .O(gate1312inter12));
  nand2 gate4129(.a(gate1312inter12), .b(gate1312inter1), .O(N5203));
nand2 gate1313( .a(N1350), .b(N4524), .O(N5204) );

  xor2  gate5292(.a(N4526), .b(N1353), .O(gate1314inter0));
  nand2 gate5293(.a(gate1314inter0), .b(s_254), .O(gate1314inter1));
  and2  gate5294(.a(N4526), .b(N1353), .O(gate1314inter2));
  inv1  gate5295(.a(s_254), .O(gate1314inter3));
  inv1  gate5296(.a(s_255), .O(gate1314inter4));
  nand2 gate5297(.a(gate1314inter4), .b(gate1314inter3), .O(gate1314inter5));
  nor2  gate5298(.a(gate1314inter5), .b(gate1314inter2), .O(gate1314inter6));
  inv1  gate5299(.a(N1353), .O(gate1314inter7));
  inv1  gate5300(.a(N4526), .O(gate1314inter8));
  nand2 gate5301(.a(gate1314inter8), .b(gate1314inter7), .O(gate1314inter9));
  nand2 gate5302(.a(s_255), .b(gate1314inter3), .O(gate1314inter10));
  nor2  gate5303(.a(gate1314inter10), .b(gate1314inter9), .O(gate1314inter11));
  nor2  gate5304(.a(gate1314inter11), .b(gate1314inter6), .O(gate1314inter12));
  nand2 gate5305(.a(gate1314inter12), .b(gate1314inter1), .O(N5205));
nand2 gate1315( .a(N1356), .b(N4528), .O(N5206) );
nand2 gate1316( .a(N1359), .b(N4530), .O(N5207) );
nand2 gate1317( .a(N1362), .b(N4532), .O(N5208) );
nand2 gate1318( .a(N1365), .b(N4534), .O(N5209) );
nand2 gate1319( .a(N1368), .b(N4536), .O(N5210) );
nand2 gate1320( .a(N1371), .b(N4538), .O(N5211) );
nand2 gate1321( .a(N1374), .b(N4540), .O(N5212) );
nand2 gate1322( .a(N1377), .b(N4542), .O(N5213) );
nand2 gate1323( .a(N3670), .b(N4611), .O(N5283) );
nand2 gate1324( .a(N3667), .b(N4612), .O(N5284) );
nand2 gate1325( .a(N3676), .b(N4613), .O(N5285) );
nand2 gate1326( .a(N3673), .b(N4614), .O(N5286) );
nand2 gate1327( .a(N3682), .b(N4615), .O(N5287) );

  xor2  gate5082(.a(N4616), .b(N3679), .O(gate1328inter0));
  nand2 gate5083(.a(gate1328inter0), .b(s_224), .O(gate1328inter1));
  and2  gate5084(.a(N4616), .b(N3679), .O(gate1328inter2));
  inv1  gate5085(.a(s_224), .O(gate1328inter3));
  inv1  gate5086(.a(s_225), .O(gate1328inter4));
  nand2 gate5087(.a(gate1328inter4), .b(gate1328inter3), .O(gate1328inter5));
  nor2  gate5088(.a(gate1328inter5), .b(gate1328inter2), .O(gate1328inter6));
  inv1  gate5089(.a(N3679), .O(gate1328inter7));
  inv1  gate5090(.a(N4616), .O(gate1328inter8));
  nand2 gate5091(.a(gate1328inter8), .b(gate1328inter7), .O(gate1328inter9));
  nand2 gate5092(.a(s_225), .b(gate1328inter3), .O(gate1328inter10));
  nor2  gate5093(.a(gate1328inter10), .b(gate1328inter9), .O(gate1328inter11));
  nor2  gate5094(.a(gate1328inter11), .b(gate1328inter6), .O(gate1328inter12));
  nand2 gate5095(.a(gate1328inter12), .b(gate1328inter1), .O(N5288));

  xor2  gate3878(.a(N4617), .b(N3688), .O(gate1329inter0));
  nand2 gate3879(.a(gate1329inter0), .b(s_52), .O(gate1329inter1));
  and2  gate3880(.a(N4617), .b(N3688), .O(gate1329inter2));
  inv1  gate3881(.a(s_52), .O(gate1329inter3));
  inv1  gate3882(.a(s_53), .O(gate1329inter4));
  nand2 gate3883(.a(gate1329inter4), .b(gate1329inter3), .O(gate1329inter5));
  nor2  gate3884(.a(gate1329inter5), .b(gate1329inter2), .O(gate1329inter6));
  inv1  gate3885(.a(N3688), .O(gate1329inter7));
  inv1  gate3886(.a(N4617), .O(gate1329inter8));
  nand2 gate3887(.a(gate1329inter8), .b(gate1329inter7), .O(gate1329inter9));
  nand2 gate3888(.a(s_53), .b(gate1329inter3), .O(gate1329inter10));
  nor2  gate3889(.a(gate1329inter10), .b(gate1329inter9), .O(gate1329inter11));
  nor2  gate3890(.a(gate1329inter11), .b(gate1329inter6), .O(gate1329inter12));
  nand2 gate3891(.a(gate1329inter12), .b(gate1329inter1), .O(N5289));

  xor2  gate5054(.a(N4618), .b(N3685), .O(gate1330inter0));
  nand2 gate5055(.a(gate1330inter0), .b(s_220), .O(gate1330inter1));
  and2  gate5056(.a(N4618), .b(N3685), .O(gate1330inter2));
  inv1  gate5057(.a(s_220), .O(gate1330inter3));
  inv1  gate5058(.a(s_221), .O(gate1330inter4));
  nand2 gate5059(.a(gate1330inter4), .b(gate1330inter3), .O(gate1330inter5));
  nor2  gate5060(.a(gate1330inter5), .b(gate1330inter2), .O(gate1330inter6));
  inv1  gate5061(.a(N3685), .O(gate1330inter7));
  inv1  gate5062(.a(N4618), .O(gate1330inter8));
  nand2 gate5063(.a(gate1330inter8), .b(gate1330inter7), .O(gate1330inter9));
  nand2 gate5064(.a(s_221), .b(gate1330inter3), .O(gate1330inter10));
  nor2  gate5065(.a(gate1330inter10), .b(gate1330inter9), .O(gate1330inter11));
  nor2  gate5066(.a(gate1330inter11), .b(gate1330inter6), .O(gate1330inter12));
  nand2 gate5067(.a(gate1330inter12), .b(gate1330inter1), .O(N5290));
nand2 gate1331( .a(N3694), .b(N4619), .O(N5291) );
nand2 gate1332( .a(N3691), .b(N4620), .O(N5292) );
nand2 gate1333( .a(N3700), .b(N4621), .O(N5293) );
nand2 gate1334( .a(N3697), .b(N4622), .O(N5294) );
nand2 gate1335( .a(N3706), .b(N4623), .O(N5295) );
nand2 gate1336( .a(N3703), .b(N4624), .O(N5296) );
nand2 gate1337( .a(N3712), .b(N4625), .O(N5297) );
nand2 gate1338( .a(N3709), .b(N4626), .O(N5298) );
nand2 gate1339( .a(N3718), .b(N4627), .O(N5299) );
nand2 gate1340( .a(N3715), .b(N4628), .O(N5300) );
nand2 gate1341( .a(N3739), .b(N4643), .O(N5314) );
nand2 gate1342( .a(N3736), .b(N4644), .O(N5315) );
nand2 gate1343( .a(N3745), .b(N4645), .O(N5316) );
nand2 gate1344( .a(N3742), .b(N4646), .O(N5317) );
nand2 gate1345( .a(N3751), .b(N4647), .O(N5318) );
nand2 gate1346( .a(N3748), .b(N4648), .O(N5319) );

  xor2  gate4690(.a(N4649), .b(N3757), .O(gate1347inter0));
  nand2 gate4691(.a(gate1347inter0), .b(s_168), .O(gate1347inter1));
  and2  gate4692(.a(N4649), .b(N3757), .O(gate1347inter2));
  inv1  gate4693(.a(s_168), .O(gate1347inter3));
  inv1  gate4694(.a(s_169), .O(gate1347inter4));
  nand2 gate4695(.a(gate1347inter4), .b(gate1347inter3), .O(gate1347inter5));
  nor2  gate4696(.a(gate1347inter5), .b(gate1347inter2), .O(gate1347inter6));
  inv1  gate4697(.a(N3757), .O(gate1347inter7));
  inv1  gate4698(.a(N4649), .O(gate1347inter8));
  nand2 gate4699(.a(gate1347inter8), .b(gate1347inter7), .O(gate1347inter9));
  nand2 gate4700(.a(s_169), .b(gate1347inter3), .O(gate1347inter10));
  nor2  gate4701(.a(gate1347inter10), .b(gate1347inter9), .O(gate1347inter11));
  nor2  gate4702(.a(gate1347inter11), .b(gate1347inter6), .O(gate1347inter12));
  nand2 gate4703(.a(gate1347inter12), .b(gate1347inter1), .O(N5320));
nand2 gate1348( .a(N3754), .b(N4650), .O(N5321) );
nand2 gate1349( .a(N3763), .b(N4651), .O(N5322) );
nand2 gate1350( .a(N3760), .b(N4652), .O(N5323) );
inv1 gate1351( .a(N4193), .O(N5324) );
nand2 gate1352( .a(N2781), .b(N4693), .O(N5363) );
nand2 gate1353( .a(N3772), .b(N4695), .O(N5364) );
nand2 gate1354( .a(N3769), .b(N4696), .O(N5365) );
nand2 gate1355( .a(N3778), .b(N4697), .O(N5366) );

  xor2  gate4606(.a(N4698), .b(N3775), .O(gate1356inter0));
  nand2 gate4607(.a(gate1356inter0), .b(s_156), .O(gate1356inter1));
  and2  gate4608(.a(N4698), .b(N3775), .O(gate1356inter2));
  inv1  gate4609(.a(s_156), .O(gate1356inter3));
  inv1  gate4610(.a(s_157), .O(gate1356inter4));
  nand2 gate4611(.a(gate1356inter4), .b(gate1356inter3), .O(gate1356inter5));
  nor2  gate4612(.a(gate1356inter5), .b(gate1356inter2), .O(gate1356inter6));
  inv1  gate4613(.a(N3775), .O(gate1356inter7));
  inv1  gate4614(.a(N4698), .O(gate1356inter8));
  nand2 gate4615(.a(gate1356inter8), .b(gate1356inter7), .O(gate1356inter9));
  nand2 gate4616(.a(s_157), .b(gate1356inter3), .O(gate1356inter10));
  nor2  gate4617(.a(gate1356inter10), .b(gate1356inter9), .O(gate1356inter11));
  nor2  gate4618(.a(gate1356inter11), .b(gate1356inter6), .O(gate1356inter12));
  nand2 gate4619(.a(gate1356inter12), .b(gate1356inter1), .O(N5367));
nand2 gate1357( .a(N2790), .b(N4745), .O(N5425) );
nand2 gate1358( .a(N3813), .b(N4747), .O(N5426) );

  xor2  gate4564(.a(N4748), .b(N3810), .O(gate1359inter0));
  nand2 gate4565(.a(gate1359inter0), .b(s_150), .O(gate1359inter1));
  and2  gate4566(.a(N4748), .b(N3810), .O(gate1359inter2));
  inv1  gate4567(.a(s_150), .O(gate1359inter3));
  inv1  gate4568(.a(s_151), .O(gate1359inter4));
  nand2 gate4569(.a(gate1359inter4), .b(gate1359inter3), .O(gate1359inter5));
  nor2  gate4570(.a(gate1359inter5), .b(gate1359inter2), .O(gate1359inter6));
  inv1  gate4571(.a(N3810), .O(gate1359inter7));
  inv1  gate4572(.a(N4748), .O(gate1359inter8));
  nand2 gate4573(.a(gate1359inter8), .b(gate1359inter7), .O(gate1359inter9));
  nand2 gate4574(.a(s_151), .b(gate1359inter3), .O(gate1359inter10));
  nor2  gate4575(.a(gate1359inter10), .b(gate1359inter9), .O(gate1359inter11));
  nor2  gate4576(.a(gate1359inter11), .b(gate1359inter6), .O(gate1359inter12));
  nand2 gate4577(.a(gate1359inter12), .b(gate1359inter1), .O(N5427));
nand2 gate1360( .a(N2793), .b(N4750), .O(N5429) );
nand2 gate1361( .a(N3825), .b(N4752), .O(N5430) );

  xor2  gate4242(.a(N4753), .b(N3822), .O(gate1362inter0));
  nand2 gate4243(.a(gate1362inter0), .b(s_104), .O(gate1362inter1));
  and2  gate4244(.a(N4753), .b(N3822), .O(gate1362inter2));
  inv1  gate4245(.a(s_104), .O(gate1362inter3));
  inv1  gate4246(.a(s_105), .O(gate1362inter4));
  nand2 gate4247(.a(gate1362inter4), .b(gate1362inter3), .O(gate1362inter5));
  nor2  gate4248(.a(gate1362inter5), .b(gate1362inter2), .O(gate1362inter6));
  inv1  gate4249(.a(N3822), .O(gate1362inter7));
  inv1  gate4250(.a(N4753), .O(gate1362inter8));
  nand2 gate4251(.a(gate1362inter8), .b(gate1362inter7), .O(gate1362inter9));
  nand2 gate4252(.a(s_105), .b(gate1362inter3), .O(gate1362inter10));
  nor2  gate4253(.a(gate1362inter10), .b(gate1362inter9), .O(gate1362inter11));
  nor2  gate4254(.a(gate1362inter11), .b(gate1362inter6), .O(gate1362inter12));
  nand2 gate4255(.a(gate1362inter12), .b(gate1362inter1), .O(N5431));
nand2 gate1363( .a(N3831), .b(N4754), .O(N5432) );

  xor2  gate4872(.a(N4755), .b(N3828), .O(gate1364inter0));
  nand2 gate4873(.a(gate1364inter0), .b(s_194), .O(gate1364inter1));
  and2  gate4874(.a(N4755), .b(N3828), .O(gate1364inter2));
  inv1  gate4875(.a(s_194), .O(gate1364inter3));
  inv1  gate4876(.a(s_195), .O(gate1364inter4));
  nand2 gate4877(.a(gate1364inter4), .b(gate1364inter3), .O(gate1364inter5));
  nor2  gate4878(.a(gate1364inter5), .b(gate1364inter2), .O(gate1364inter6));
  inv1  gate4879(.a(N3828), .O(gate1364inter7));
  inv1  gate4880(.a(N4755), .O(gate1364inter8));
  nand2 gate4881(.a(gate1364inter8), .b(gate1364inter7), .O(gate1364inter9));
  nand2 gate4882(.a(s_195), .b(gate1364inter3), .O(gate1364inter10));
  nor2  gate4883(.a(gate1364inter10), .b(gate1364inter9), .O(gate1364inter11));
  nor2  gate4884(.a(gate1364inter11), .b(gate1364inter6), .O(gate1364inter12));
  nand2 gate4885(.a(gate1364inter12), .b(gate1364inter1), .O(N5433));
nand2 gate1365( .a(N2796), .b(N4775), .O(N5451) );
nand2 gate1366( .a(N3864), .b(N4777), .O(N5452) );

  xor2  gate4186(.a(N4778), .b(N3861), .O(gate1367inter0));
  nand2 gate4187(.a(gate1367inter0), .b(s_96), .O(gate1367inter1));
  and2  gate4188(.a(N4778), .b(N3861), .O(gate1367inter2));
  inv1  gate4189(.a(s_96), .O(gate1367inter3));
  inv1  gate4190(.a(s_97), .O(gate1367inter4));
  nand2 gate4191(.a(gate1367inter4), .b(gate1367inter3), .O(gate1367inter5));
  nor2  gate4192(.a(gate1367inter5), .b(gate1367inter2), .O(gate1367inter6));
  inv1  gate4193(.a(N3861), .O(gate1367inter7));
  inv1  gate4194(.a(N4778), .O(gate1367inter8));
  nand2 gate4195(.a(gate1367inter8), .b(gate1367inter7), .O(gate1367inter9));
  nand2 gate4196(.a(s_97), .b(gate1367inter3), .O(gate1367inter10));
  nor2  gate4197(.a(gate1367inter10), .b(gate1367inter9), .O(gate1367inter11));
  nor2  gate4198(.a(gate1367inter11), .b(gate1367inter6), .O(gate1367inter12));
  nand2 gate4199(.a(gate1367inter12), .b(gate1367inter1), .O(N5453));
nand2 gate1368( .a(N3870), .b(N4779), .O(N5454) );
nand2 gate1369( .a(N3867), .b(N4780), .O(N5455) );
nand2 gate1370( .a(N3888), .b(N4781), .O(N5456) );

  xor2  gate5012(.a(N4782), .b(N3885), .O(gate1371inter0));
  nand2 gate5013(.a(gate1371inter0), .b(s_214), .O(gate1371inter1));
  and2  gate5014(.a(N4782), .b(N3885), .O(gate1371inter2));
  inv1  gate5015(.a(s_214), .O(gate1371inter3));
  inv1  gate5016(.a(s_215), .O(gate1371inter4));
  nand2 gate5017(.a(gate1371inter4), .b(gate1371inter3), .O(gate1371inter5));
  nor2  gate5018(.a(gate1371inter5), .b(gate1371inter2), .O(gate1371inter6));
  inv1  gate5019(.a(N3885), .O(gate1371inter7));
  inv1  gate5020(.a(N4782), .O(gate1371inter8));
  nand2 gate5021(.a(gate1371inter8), .b(gate1371inter7), .O(gate1371inter9));
  nand2 gate5022(.a(s_215), .b(gate1371inter3), .O(gate1371inter10));
  nor2  gate5023(.a(gate1371inter10), .b(gate1371inter9), .O(gate1371inter11));
  nor2  gate5024(.a(gate1371inter11), .b(gate1371inter6), .O(gate1371inter12));
  nand2 gate5025(.a(gate1371inter12), .b(gate1371inter1), .O(N5457));
inv1 gate1372( .a(N4303), .O(N5469) );
nand2 gate1373( .a(N3589), .b(N4799), .O(N5474) );
nand2 gate1374( .a(N3586), .b(N4800), .O(N5475) );
nand2 gate1375( .a(N3595), .b(N4801), .O(N5476) );
nand2 gate1376( .a(N3592), .b(N4802), .O(N5477) );
nand2 gate1377( .a(N3798), .b(N5045), .O(N5571) );
nand2 gate1378( .a(N3795), .b(N5046), .O(N5572) );

  xor2  gate3850(.a(N5047), .b(N3804), .O(gate1379inter0));
  nand2 gate3851(.a(gate1379inter0), .b(s_48), .O(gate1379inter1));
  and2  gate3852(.a(N5047), .b(N3804), .O(gate1379inter2));
  inv1  gate3853(.a(s_48), .O(gate1379inter3));
  inv1  gate3854(.a(s_49), .O(gate1379inter4));
  nand2 gate3855(.a(gate1379inter4), .b(gate1379inter3), .O(gate1379inter5));
  nor2  gate3856(.a(gate1379inter5), .b(gate1379inter2), .O(gate1379inter6));
  inv1  gate3857(.a(N3804), .O(gate1379inter7));
  inv1  gate3858(.a(N5047), .O(gate1379inter8));
  nand2 gate3859(.a(gate1379inter8), .b(gate1379inter7), .O(gate1379inter9));
  nand2 gate3860(.a(s_49), .b(gate1379inter3), .O(gate1379inter10));
  nor2  gate3861(.a(gate1379inter10), .b(gate1379inter9), .O(gate1379inter11));
  nor2  gate3862(.a(gate1379inter11), .b(gate1379inter6), .O(gate1379inter12));
  nand2 gate3863(.a(gate1379inter12), .b(gate1379inter1), .O(N5573));
nand2 gate1380( .a(N3801), .b(N5048), .O(N5574) );
nand2 gate1381( .a(N3837), .b(N5064), .O(N5584) );
nand2 gate1382( .a(N3834), .b(N5065), .O(N5585) );
nand2 gate1383( .a(N3843), .b(N5066), .O(N5586) );
nand2 gate1384( .a(N3840), .b(N5067), .O(N5587) );
nand2 gate1385( .a(N3876), .b(N5110), .O(N5602) );
nand2 gate1386( .a(N3873), .b(N5111), .O(N5603) );
nand2 gate1387( .a(N3882), .b(N5112), .O(N5604) );
nand2 gate1388( .a(N3879), .b(N5113), .O(N5605) );
nand2 gate1389( .a(N5324), .b(N4653), .O(N5631) );
nand2 gate1390( .a(N4463), .b(N5167), .O(N5632) );

  xor2  gate4928(.a(N5168), .b(N4465), .O(gate1391inter0));
  nand2 gate4929(.a(gate1391inter0), .b(s_202), .O(gate1391inter1));
  and2  gate4930(.a(N5168), .b(N4465), .O(gate1391inter2));
  inv1  gate4931(.a(s_202), .O(gate1391inter3));
  inv1  gate4932(.a(s_203), .O(gate1391inter4));
  nand2 gate4933(.a(gate1391inter4), .b(gate1391inter3), .O(gate1391inter5));
  nor2  gate4934(.a(gate1391inter5), .b(gate1391inter2), .O(gate1391inter6));
  inv1  gate4935(.a(N4465), .O(gate1391inter7));
  inv1  gate4936(.a(N5168), .O(gate1391inter8));
  nand2 gate4937(.a(gate1391inter8), .b(gate1391inter7), .O(gate1391inter9));
  nand2 gate4938(.a(s_203), .b(gate1391inter3), .O(gate1391inter10));
  nor2  gate4939(.a(gate1391inter10), .b(gate1391inter9), .O(gate1391inter11));
  nor2  gate4940(.a(gate1391inter11), .b(gate1391inter6), .O(gate1391inter12));
  nand2 gate4941(.a(gate1391inter12), .b(gate1391inter1), .O(N5640));
nand2 gate1392( .a(N4467), .b(N5169), .O(N5654) );
nand2 gate1393( .a(N4469), .b(N5170), .O(N5670) );
nand2 gate1394( .a(N4471), .b(N5171), .O(N5683) );
nand2 gate1395( .a(N4475), .b(N5172), .O(N5690) );
nand2 gate1396( .a(N4477), .b(N5173), .O(N5697) );

  xor2  gate4676(.a(N5174), .b(N4479), .O(gate1397inter0));
  nand2 gate4677(.a(gate1397inter0), .b(s_166), .O(gate1397inter1));
  and2  gate4678(.a(N5174), .b(N4479), .O(gate1397inter2));
  inv1  gate4679(.a(s_166), .O(gate1397inter3));
  inv1  gate4680(.a(s_167), .O(gate1397inter4));
  nand2 gate4681(.a(gate1397inter4), .b(gate1397inter3), .O(gate1397inter5));
  nor2  gate4682(.a(gate1397inter5), .b(gate1397inter2), .O(gate1397inter6));
  inv1  gate4683(.a(N4479), .O(gate1397inter7));
  inv1  gate4684(.a(N5174), .O(gate1397inter8));
  nand2 gate4685(.a(gate1397inter8), .b(gate1397inter7), .O(gate1397inter9));
  nand2 gate4686(.a(s_167), .b(gate1397inter3), .O(gate1397inter10));
  nor2  gate4687(.a(gate1397inter10), .b(gate1397inter9), .O(gate1397inter11));
  nor2  gate4688(.a(gate1397inter11), .b(gate1397inter6), .O(gate1397inter12));
  nand2 gate4689(.a(gate1397inter12), .b(gate1397inter1), .O(N5707));
nand2 gate1398( .a(N4481), .b(N5175), .O(N5718) );
nand2 gate1399( .a(N4483), .b(N5176), .O(N5728) );
inv1 gate1400( .a(N5177), .O(N5735) );
nand2 gate1401( .a(N5179), .b(N4490), .O(N5736) );
nand2 gate1402( .a(N5180), .b(N5181), .O(N5740) );
nand2 gate1403( .a(N5182), .b(N5183), .O(N5744) );
nand2 gate1404( .a(N5184), .b(N4496), .O(N5747) );

  xor2  gate3640(.a(N5186), .b(N5185), .O(gate1405inter0));
  nand2 gate3641(.a(gate1405inter0), .b(s_18), .O(gate1405inter1));
  and2  gate3642(.a(N5186), .b(N5185), .O(gate1405inter2));
  inv1  gate3643(.a(s_18), .O(gate1405inter3));
  inv1  gate3644(.a(s_19), .O(gate1405inter4));
  nand2 gate3645(.a(gate1405inter4), .b(gate1405inter3), .O(gate1405inter5));
  nor2  gate3646(.a(gate1405inter5), .b(gate1405inter2), .O(gate1405inter6));
  inv1  gate3647(.a(N5185), .O(gate1405inter7));
  inv1  gate3648(.a(N5186), .O(gate1405inter8));
  nand2 gate3649(.a(gate1405inter8), .b(gate1405inter7), .O(gate1405inter9));
  nand2 gate3650(.a(s_19), .b(gate1405inter3), .O(gate1405inter10));
  nor2  gate3651(.a(gate1405inter10), .b(gate1405inter9), .O(gate1405inter11));
  nor2  gate3652(.a(gate1405inter11), .b(gate1405inter6), .O(gate1405inter12));
  nand2 gate3653(.a(gate1405inter12), .b(gate1405inter1), .O(N5751));
nand2 gate1406( .a(N5187), .b(N5188), .O(N5755) );
nand2 gate1407( .a(N5189), .b(N4502), .O(N5758) );
nand2 gate1408( .a(N5190), .b(N5191), .O(N5762) );
nand2 gate1409( .a(N5192), .b(N5193), .O(N5766) );
inv1 gate1410( .a(N4803), .O(N5769) );
inv1 gate1411( .a(N4806), .O(N5770) );

  xor2  gate3962(.a(N5196), .b(N4507), .O(gate1412inter0));
  nand2 gate3963(.a(gate1412inter0), .b(s_64), .O(gate1412inter1));
  and2  gate3964(.a(N5196), .b(N4507), .O(gate1412inter2));
  inv1  gate3965(.a(s_64), .O(gate1412inter3));
  inv1  gate3966(.a(s_65), .O(gate1412inter4));
  nand2 gate3967(.a(gate1412inter4), .b(gate1412inter3), .O(gate1412inter5));
  nor2  gate3968(.a(gate1412inter5), .b(gate1412inter2), .O(gate1412inter6));
  inv1  gate3969(.a(N4507), .O(gate1412inter7));
  inv1  gate3970(.a(N5196), .O(gate1412inter8));
  nand2 gate3971(.a(gate1412inter8), .b(gate1412inter7), .O(gate1412inter9));
  nand2 gate3972(.a(s_65), .b(gate1412inter3), .O(gate1412inter10));
  nor2  gate3973(.a(gate1412inter10), .b(gate1412inter9), .O(gate1412inter11));
  nor2  gate3974(.a(gate1412inter11), .b(gate1412inter6), .O(gate1412inter12));
  nand2 gate3975(.a(gate1412inter12), .b(gate1412inter1), .O(N5771));
nand2 gate1413( .a(N4509), .b(N5197), .O(N5778) );
nand2 gate1414( .a(N4511), .b(N5198), .O(N5789) );
nand2 gate1415( .a(N4513), .b(N5199), .O(N5799) );
nand2 gate1416( .a(N4515), .b(N5200), .O(N5807) );
nand2 gate1417( .a(N4517), .b(N5201), .O(N5821) );
nand2 gate1418( .a(N4519), .b(N5202), .O(N5837) );
nand2 gate1419( .a(N4521), .b(N5203), .O(N5850) );
nand2 gate1420( .a(N4523), .b(N5204), .O(N5856) );

  xor2  gate3598(.a(N5205), .b(N4525), .O(gate1421inter0));
  nand2 gate3599(.a(gate1421inter0), .b(s_12), .O(gate1421inter1));
  and2  gate3600(.a(N5205), .b(N4525), .O(gate1421inter2));
  inv1  gate3601(.a(s_12), .O(gate1421inter3));
  inv1  gate3602(.a(s_13), .O(gate1421inter4));
  nand2 gate3603(.a(gate1421inter4), .b(gate1421inter3), .O(gate1421inter5));
  nor2  gate3604(.a(gate1421inter5), .b(gate1421inter2), .O(gate1421inter6));
  inv1  gate3605(.a(N4525), .O(gate1421inter7));
  inv1  gate3606(.a(N5205), .O(gate1421inter8));
  nand2 gate3607(.a(gate1421inter8), .b(gate1421inter7), .O(gate1421inter9));
  nand2 gate3608(.a(s_13), .b(gate1421inter3), .O(gate1421inter10));
  nor2  gate3609(.a(gate1421inter10), .b(gate1421inter9), .O(gate1421inter11));
  nor2  gate3610(.a(gate1421inter11), .b(gate1421inter6), .O(gate1421inter12));
  nand2 gate3611(.a(gate1421inter12), .b(gate1421inter1), .O(N5863));
nand2 gate1422( .a(N4527), .b(N5206), .O(N5870) );
nand2 gate1423( .a(N4529), .b(N5207), .O(N5881) );
nand2 gate1424( .a(N4531), .b(N5208), .O(N5892) );
nand2 gate1425( .a(N4533), .b(N5209), .O(N5898) );
nand2 gate1426( .a(N4535), .b(N5210), .O(N5905) );
nand2 gate1427( .a(N4537), .b(N5211), .O(N5915) );
nand2 gate1428( .a(N4539), .b(N5212), .O(N5926) );
nand2 gate1429( .a(N4541), .b(N5213), .O(N5936) );
inv1 gate1430( .a(N4817), .O(N5943) );
nand2 gate1431( .a(N4820), .b(N1931), .O(N5944) );
inv1 gate1432( .a(N4820), .O(N5945) );
nand2 gate1433( .a(N4823), .b(N1932), .O(N5946) );
inv1 gate1434( .a(N4823), .O(N5947) );
nand2 gate1435( .a(N4826), .b(N1933), .O(N5948) );
inv1 gate1436( .a(N4826), .O(N5949) );
nand2 gate1437( .a(N4829), .b(N1934), .O(N5950) );
inv1 gate1438( .a(N4829), .O(N5951) );
nand2 gate1439( .a(N4832), .b(N1935), .O(N5952) );
inv1 gate1440( .a(N4832), .O(N5953) );
nand2 gate1441( .a(N4835), .b(N1936), .O(N5954) );
inv1 gate1442( .a(N4835), .O(N5955) );
nand2 gate1443( .a(N4838), .b(N1937), .O(N5956) );
inv1 gate1444( .a(N4838), .O(N5957) );
nand2 gate1445( .a(N4841), .b(N1938), .O(N5958) );
inv1 gate1446( .a(N4841), .O(N5959) );
and2 gate1447( .a(N2674), .b(N4769), .O(N5960) );
inv1 gate1448( .a(N4844), .O(N5966) );
nand2 gate1449( .a(N4847), .b(N1939), .O(N5967) );
inv1 gate1450( .a(N4847), .O(N5968) );
nand2 gate1451( .a(N4850), .b(N1940), .O(N5969) );
inv1 gate1452( .a(N4850), .O(N5970) );
nand2 gate1453( .a(N4853), .b(N1941), .O(N5971) );
inv1 gate1454( .a(N4853), .O(N5972) );
nand2 gate1455( .a(N4856), .b(N1942), .O(N5973) );
inv1 gate1456( .a(N4856), .O(N5974) );
nand2 gate1457( .a(N4859), .b(N1943), .O(N5975) );
inv1 gate1458( .a(N4859), .O(N5976) );
nand2 gate1459( .a(N4862), .b(N1944), .O(N5977) );
inv1 gate1460( .a(N4862), .O(N5978) );
nand2 gate1461( .a(N4865), .b(N1945), .O(N5979) );
inv1 gate1462( .a(N4865), .O(N5980) );
and2 gate1463( .a(N2674), .b(N4769), .O(N5981) );
nand2 gate1464( .a(N4868), .b(N1946), .O(N5989) );
inv1 gate1465( .a(N4868), .O(N5990) );

  xor2  gate4956(.a(N5284), .b(N5283), .O(gate1466inter0));
  nand2 gate4957(.a(gate1466inter0), .b(s_206), .O(gate1466inter1));
  and2  gate4958(.a(N5284), .b(N5283), .O(gate1466inter2));
  inv1  gate4959(.a(s_206), .O(gate1466inter3));
  inv1  gate4960(.a(s_207), .O(gate1466inter4));
  nand2 gate4961(.a(gate1466inter4), .b(gate1466inter3), .O(gate1466inter5));
  nor2  gate4962(.a(gate1466inter5), .b(gate1466inter2), .O(gate1466inter6));
  inv1  gate4963(.a(N5283), .O(gate1466inter7));
  inv1  gate4964(.a(N5284), .O(gate1466inter8));
  nand2 gate4965(.a(gate1466inter8), .b(gate1466inter7), .O(gate1466inter9));
  nand2 gate4966(.a(s_207), .b(gate1466inter3), .O(gate1466inter10));
  nor2  gate4967(.a(gate1466inter10), .b(gate1466inter9), .O(gate1466inter11));
  nor2  gate4968(.a(gate1466inter11), .b(gate1466inter6), .O(gate1466inter12));
  nand2 gate4969(.a(gate1466inter12), .b(gate1466inter1), .O(N5991));
nand2 gate1467( .a(N5285), .b(N5286), .O(N5996) );
nand2 gate1468( .a(N5287), .b(N5288), .O(N6000) );
nand2 gate1469( .a(N5289), .b(N5290), .O(N6003) );
nand2 gate1470( .a(N5291), .b(N5292), .O(N6009) );
nand2 gate1471( .a(N5293), .b(N5294), .O(N6014) );
nand2 gate1472( .a(N5295), .b(N5296), .O(N6018) );
nand2 gate1473( .a(N5297), .b(N5298), .O(N6021) );

  xor2  gate5320(.a(N5300), .b(N5299), .O(gate1474inter0));
  nand2 gate5321(.a(gate1474inter0), .b(s_258), .O(gate1474inter1));
  and2  gate5322(.a(N5300), .b(N5299), .O(gate1474inter2));
  inv1  gate5323(.a(s_258), .O(gate1474inter3));
  inv1  gate5324(.a(s_259), .O(gate1474inter4));
  nand2 gate5325(.a(gate1474inter4), .b(gate1474inter3), .O(gate1474inter5));
  nor2  gate5326(.a(gate1474inter5), .b(gate1474inter2), .O(gate1474inter6));
  inv1  gate5327(.a(N5299), .O(gate1474inter7));
  inv1  gate5328(.a(N5300), .O(gate1474inter8));
  nand2 gate5329(.a(gate1474inter8), .b(gate1474inter7), .O(gate1474inter9));
  nand2 gate5330(.a(s_259), .b(gate1474inter3), .O(gate1474inter10));
  nor2  gate5331(.a(gate1474inter10), .b(gate1474inter9), .O(gate1474inter11));
  nor2  gate5332(.a(gate1474inter11), .b(gate1474inter6), .O(gate1474inter12));
  nand2 gate5333(.a(gate1474inter12), .b(gate1474inter1), .O(N6022));
inv1 gate1475( .a(N4874), .O(N6023) );
nand2 gate1476( .a(N4874), .b(N4629), .O(N6024) );
inv1 gate1477( .a(N4877), .O(N6025) );

  xor2  gate4704(.a(N4631), .b(N4877), .O(gate1478inter0));
  nand2 gate4705(.a(gate1478inter0), .b(s_170), .O(gate1478inter1));
  and2  gate4706(.a(N4631), .b(N4877), .O(gate1478inter2));
  inv1  gate4707(.a(s_170), .O(gate1478inter3));
  inv1  gate4708(.a(s_171), .O(gate1478inter4));
  nand2 gate4709(.a(gate1478inter4), .b(gate1478inter3), .O(gate1478inter5));
  nor2  gate4710(.a(gate1478inter5), .b(gate1478inter2), .O(gate1478inter6));
  inv1  gate4711(.a(N4877), .O(gate1478inter7));
  inv1  gate4712(.a(N4631), .O(gate1478inter8));
  nand2 gate4713(.a(gate1478inter8), .b(gate1478inter7), .O(gate1478inter9));
  nand2 gate4714(.a(s_171), .b(gate1478inter3), .O(gate1478inter10));
  nor2  gate4715(.a(gate1478inter10), .b(gate1478inter9), .O(gate1478inter11));
  nor2  gate4716(.a(gate1478inter11), .b(gate1478inter6), .O(gate1478inter12));
  nand2 gate4717(.a(gate1478inter12), .b(gate1478inter1), .O(N6026));
inv1 gate1479( .a(N4880), .O(N6027) );
nand2 gate1480( .a(N4880), .b(N4633), .O(N6028) );
inv1 gate1481( .a(N4883), .O(N6029) );
nand2 gate1482( .a(N4883), .b(N4636), .O(N6030) );
inv1 gate1483( .a(N4886), .O(N6031) );
inv1 gate1484( .a(N4889), .O(N6032) );
inv1 gate1485( .a(N4892), .O(N6033) );
inv1 gate1486( .a(N4895), .O(N6034) );
inv1 gate1487( .a(N4898), .O(N6035) );
inv1 gate1488( .a(N4901), .O(N6036) );
inv1 gate1489( .a(N4904), .O(N6037) );
nand2 gate1490( .a(N4904), .b(N4642), .O(N6038) );
inv1 gate1491( .a(N4907), .O(N6039) );
inv1 gate1492( .a(N4910), .O(N6040) );
nand2 gate1493( .a(N5314), .b(N5315), .O(N6041) );
nand2 gate1494( .a(N5316), .b(N5317), .O(N6047) );

  xor2  gate3570(.a(N5319), .b(N5318), .O(gate1495inter0));
  nand2 gate3571(.a(gate1495inter0), .b(s_8), .O(gate1495inter1));
  and2  gate3572(.a(N5319), .b(N5318), .O(gate1495inter2));
  inv1  gate3573(.a(s_8), .O(gate1495inter3));
  inv1  gate3574(.a(s_9), .O(gate1495inter4));
  nand2 gate3575(.a(gate1495inter4), .b(gate1495inter3), .O(gate1495inter5));
  nor2  gate3576(.a(gate1495inter5), .b(gate1495inter2), .O(gate1495inter6));
  inv1  gate3577(.a(N5318), .O(gate1495inter7));
  inv1  gate3578(.a(N5319), .O(gate1495inter8));
  nand2 gate3579(.a(gate1495inter8), .b(gate1495inter7), .O(gate1495inter9));
  nand2 gate3580(.a(s_9), .b(gate1495inter3), .O(gate1495inter10));
  nor2  gate3581(.a(gate1495inter10), .b(gate1495inter9), .O(gate1495inter11));
  nor2  gate3582(.a(gate1495inter11), .b(gate1495inter6), .O(gate1495inter12));
  nand2 gate3583(.a(gate1495inter12), .b(gate1495inter1), .O(N6052));
nand2 gate1496( .a(N5320), .b(N5321), .O(N6056) );
nand2 gate1497( .a(N5322), .b(N5323), .O(N6059) );
nand2 gate1498( .a(N4913), .b(N1968), .O(N6060) );
inv1 gate1499( .a(N4913), .O(N6061) );
nand2 gate1500( .a(N4916), .b(N1969), .O(N6062) );
inv1 gate1501( .a(N4916), .O(N6063) );
nand2 gate1502( .a(N4919), .b(N1970), .O(N6064) );
inv1 gate1503( .a(N4919), .O(N6065) );
nand2 gate1504( .a(N4922), .b(N1971), .O(N6066) );
inv1 gate1505( .a(N4922), .O(N6067) );
nand2 gate1506( .a(N4925), .b(N1972), .O(N6068) );
inv1 gate1507( .a(N4925), .O(N6069) );
nand2 gate1508( .a(N4928), .b(N1973), .O(N6070) );
inv1 gate1509( .a(N4928), .O(N6071) );

  xor2  gate4130(.a(N1974), .b(N4931), .O(gate1510inter0));
  nand2 gate4131(.a(gate1510inter0), .b(s_88), .O(gate1510inter1));
  and2  gate4132(.a(N1974), .b(N4931), .O(gate1510inter2));
  inv1  gate4133(.a(s_88), .O(gate1510inter3));
  inv1  gate4134(.a(s_89), .O(gate1510inter4));
  nand2 gate4135(.a(gate1510inter4), .b(gate1510inter3), .O(gate1510inter5));
  nor2  gate4136(.a(gate1510inter5), .b(gate1510inter2), .O(gate1510inter6));
  inv1  gate4137(.a(N4931), .O(gate1510inter7));
  inv1  gate4138(.a(N1974), .O(gate1510inter8));
  nand2 gate4139(.a(gate1510inter8), .b(gate1510inter7), .O(gate1510inter9));
  nand2 gate4140(.a(s_89), .b(gate1510inter3), .O(gate1510inter10));
  nor2  gate4141(.a(gate1510inter10), .b(gate1510inter9), .O(gate1510inter11));
  nor2  gate4142(.a(gate1510inter11), .b(gate1510inter6), .O(gate1510inter12));
  nand2 gate4143(.a(gate1510inter12), .b(gate1510inter1), .O(N6072));
inv1 gate1511( .a(N4931), .O(N6073) );
nand2 gate1512( .a(N4934), .b(N1975), .O(N6074) );
inv1 gate1513( .a(N4934), .O(N6075) );
nand2 gate1514( .a(N4937), .b(N1976), .O(N6076) );
inv1 gate1515( .a(N4937), .O(N6077) );
inv1 gate1516( .a(N4940), .O(N6078) );
nand2 gate1517( .a(N5363), .b(N4694), .O(N6079) );
nand2 gate1518( .a(N5364), .b(N5365), .O(N6083) );
nand2 gate1519( .a(N5366), .b(N5367), .O(N6087) );
inv1 gate1520( .a(N4943), .O(N6090) );
nand2 gate1521( .a(N4943), .b(N4699), .O(N6091) );
inv1 gate1522( .a(N4946), .O(N6092) );
inv1 gate1523( .a(N4949), .O(N6093) );
inv1 gate1524( .a(N4952), .O(N6094) );
inv1 gate1525( .a(N4955), .O(N6095) );
inv1 gate1526( .a(N4970), .O(N6096) );
nand2 gate1527( .a(N4970), .b(N4700), .O(N6097) );
inv1 gate1528( .a(N4973), .O(N6098) );
inv1 gate1529( .a(N4976), .O(N6099) );
inv1 gate1530( .a(N4979), .O(N6100) );
inv1 gate1531( .a(N4982), .O(N6101) );
inv1 gate1532( .a(N4997), .O(N6102) );
nand2 gate1533( .a(N5000), .b(N2015), .O(N6103) );
inv1 gate1534( .a(N5000), .O(N6104) );

  xor2  gate4578(.a(N2016), .b(N5003), .O(gate1535inter0));
  nand2 gate4579(.a(gate1535inter0), .b(s_152), .O(gate1535inter1));
  and2  gate4580(.a(N2016), .b(N5003), .O(gate1535inter2));
  inv1  gate4581(.a(s_152), .O(gate1535inter3));
  inv1  gate4582(.a(s_153), .O(gate1535inter4));
  nand2 gate4583(.a(gate1535inter4), .b(gate1535inter3), .O(gate1535inter5));
  nor2  gate4584(.a(gate1535inter5), .b(gate1535inter2), .O(gate1535inter6));
  inv1  gate4585(.a(N5003), .O(gate1535inter7));
  inv1  gate4586(.a(N2016), .O(gate1535inter8));
  nand2 gate4587(.a(gate1535inter8), .b(gate1535inter7), .O(gate1535inter9));
  nand2 gate4588(.a(s_153), .b(gate1535inter3), .O(gate1535inter10));
  nor2  gate4589(.a(gate1535inter10), .b(gate1535inter9), .O(gate1535inter11));
  nor2  gate4590(.a(gate1535inter11), .b(gate1535inter6), .O(gate1535inter12));
  nand2 gate4591(.a(gate1535inter12), .b(gate1535inter1), .O(N6105));
inv1 gate1536( .a(N5003), .O(N6106) );

  xor2  gate4536(.a(N2017), .b(N5006), .O(gate1537inter0));
  nand2 gate4537(.a(gate1537inter0), .b(s_146), .O(gate1537inter1));
  and2  gate4538(.a(N2017), .b(N5006), .O(gate1537inter2));
  inv1  gate4539(.a(s_146), .O(gate1537inter3));
  inv1  gate4540(.a(s_147), .O(gate1537inter4));
  nand2 gate4541(.a(gate1537inter4), .b(gate1537inter3), .O(gate1537inter5));
  nor2  gate4542(.a(gate1537inter5), .b(gate1537inter2), .O(gate1537inter6));
  inv1  gate4543(.a(N5006), .O(gate1537inter7));
  inv1  gate4544(.a(N2017), .O(gate1537inter8));
  nand2 gate4545(.a(gate1537inter8), .b(gate1537inter7), .O(gate1537inter9));
  nand2 gate4546(.a(s_147), .b(gate1537inter3), .O(gate1537inter10));
  nor2  gate4547(.a(gate1537inter10), .b(gate1537inter9), .O(gate1537inter11));
  nor2  gate4548(.a(gate1537inter11), .b(gate1537inter6), .O(gate1537inter12));
  nand2 gate4549(.a(gate1537inter12), .b(gate1537inter1), .O(N6107));
inv1 gate1538( .a(N5006), .O(N6108) );
nand2 gate1539( .a(N5009), .b(N2018), .O(N6109) );
inv1 gate1540( .a(N5009), .O(N6110) );
nand2 gate1541( .a(N5012), .b(N2019), .O(N6111) );
inv1 gate1542( .a(N5012), .O(N6112) );
nand2 gate1543( .a(N5015), .b(N2020), .O(N6113) );
inv1 gate1544( .a(N5015), .O(N6114) );
nand2 gate1545( .a(N5018), .b(N2021), .O(N6115) );
inv1 gate1546( .a(N5018), .O(N6116) );
nand2 gate1547( .a(N5021), .b(N2022), .O(N6117) );
inv1 gate1548( .a(N5021), .O(N6118) );
nand2 gate1549( .a(N5024), .b(N2023), .O(N6119) );
inv1 gate1550( .a(N5024), .O(N6120) );
inv1 gate1551( .a(N5033), .O(N6121) );
nand2 gate1552( .a(N5033), .b(N4743), .O(N6122) );
inv1 gate1553( .a(N5036), .O(N6123) );
inv1 gate1554( .a(N5039), .O(N6124) );

  xor2  gate4620(.a(N4744), .b(N5042), .O(gate1555inter0));
  nand2 gate4621(.a(gate1555inter0), .b(s_158), .O(gate1555inter1));
  and2  gate4622(.a(N4744), .b(N5042), .O(gate1555inter2));
  inv1  gate4623(.a(s_158), .O(gate1555inter3));
  inv1  gate4624(.a(s_159), .O(gate1555inter4));
  nand2 gate4625(.a(gate1555inter4), .b(gate1555inter3), .O(gate1555inter5));
  nor2  gate4626(.a(gate1555inter5), .b(gate1555inter2), .O(gate1555inter6));
  inv1  gate4627(.a(N5042), .O(gate1555inter7));
  inv1  gate4628(.a(N4744), .O(gate1555inter8));
  nand2 gate4629(.a(gate1555inter8), .b(gate1555inter7), .O(gate1555inter9));
  nand2 gate4630(.a(s_159), .b(gate1555inter3), .O(gate1555inter10));
  nor2  gate4631(.a(gate1555inter10), .b(gate1555inter9), .O(gate1555inter11));
  nor2  gate4632(.a(gate1555inter11), .b(gate1555inter6), .O(gate1555inter12));
  nand2 gate4633(.a(gate1555inter12), .b(gate1555inter1), .O(N6125));
inv1 gate1556( .a(N5042), .O(N6126) );

  xor2  gate4060(.a(N4746), .b(N5425), .O(gate1557inter0));
  nand2 gate4061(.a(gate1557inter0), .b(s_78), .O(gate1557inter1));
  and2  gate4062(.a(N4746), .b(N5425), .O(gate1557inter2));
  inv1  gate4063(.a(s_78), .O(gate1557inter3));
  inv1  gate4064(.a(s_79), .O(gate1557inter4));
  nand2 gate4065(.a(gate1557inter4), .b(gate1557inter3), .O(gate1557inter5));
  nor2  gate4066(.a(gate1557inter5), .b(gate1557inter2), .O(gate1557inter6));
  inv1  gate4067(.a(N5425), .O(gate1557inter7));
  inv1  gate4068(.a(N4746), .O(gate1557inter8));
  nand2 gate4069(.a(gate1557inter8), .b(gate1557inter7), .O(gate1557inter9));
  nand2 gate4070(.a(s_79), .b(gate1557inter3), .O(gate1557inter10));
  nor2  gate4071(.a(gate1557inter10), .b(gate1557inter9), .O(gate1557inter11));
  nor2  gate4072(.a(gate1557inter11), .b(gate1557inter6), .O(gate1557inter12));
  nand2 gate4073(.a(gate1557inter12), .b(gate1557inter1), .O(N6127));

  xor2  gate5208(.a(N5427), .b(N5426), .O(gate1558inter0));
  nand2 gate5209(.a(gate1558inter0), .b(s_242), .O(gate1558inter1));
  and2  gate5210(.a(N5427), .b(N5426), .O(gate1558inter2));
  inv1  gate5211(.a(s_242), .O(gate1558inter3));
  inv1  gate5212(.a(s_243), .O(gate1558inter4));
  nand2 gate5213(.a(gate1558inter4), .b(gate1558inter3), .O(gate1558inter5));
  nor2  gate5214(.a(gate1558inter5), .b(gate1558inter2), .O(gate1558inter6));
  inv1  gate5215(.a(N5426), .O(gate1558inter7));
  inv1  gate5216(.a(N5427), .O(gate1558inter8));
  nand2 gate5217(.a(gate1558inter8), .b(gate1558inter7), .O(gate1558inter9));
  nand2 gate5218(.a(s_243), .b(gate1558inter3), .O(gate1558inter10));
  nor2  gate5219(.a(gate1558inter10), .b(gate1558inter9), .O(gate1558inter11));
  nor2  gate5220(.a(gate1558inter11), .b(gate1558inter6), .O(gate1558inter12));
  nand2 gate5221(.a(gate1558inter12), .b(gate1558inter1), .O(N6131));
inv1 gate1559( .a(N5049), .O(N6135) );
nand2 gate1560( .a(N5049), .b(N4749), .O(N6136) );
nand2 gate1561( .a(N5429), .b(N4751), .O(N6137) );
nand2 gate1562( .a(N5430), .b(N5431), .O(N6141) );
nand2 gate1563( .a(N5432), .b(N5433), .O(N6145) );
inv1 gate1564( .a(N5068), .O(N6148) );
inv1 gate1565( .a(N5071), .O(N6149) );
inv1 gate1566( .a(N5074), .O(N6150) );
inv1 gate1567( .a(N5077), .O(N6151) );
inv1 gate1568( .a(N5080), .O(N6152) );
inv1 gate1569( .a(N5083), .O(N6153) );
inv1 gate1570( .a(N5086), .O(N6154) );
inv1 gate1571( .a(N5089), .O(N6155) );
inv1 gate1572( .a(N5092), .O(N6156) );
nand2 gate1573( .a(N5092), .b(N4761), .O(N6157) );
inv1 gate1574( .a(N5095), .O(N6158) );
nand2 gate1575( .a(N5095), .b(N4763), .O(N6159) );
inv1 gate1576( .a(N5098), .O(N6160) );
nand2 gate1577( .a(N5098), .b(N4765), .O(N6161) );
inv1 gate1578( .a(N5101), .O(N6162) );
inv1 gate1579( .a(N5104), .O(N6163) );
nand2 gate1580( .a(N5107), .b(N4768), .O(N6164) );
inv1 gate1581( .a(N5107), .O(N6165) );
nand2 gate1582( .a(N5451), .b(N4776), .O(N6166) );
nand2 gate1583( .a(N5452), .b(N5453), .O(N6170) );
nand2 gate1584( .a(N5454), .b(N5455), .O(N6174) );
nand2 gate1585( .a(N5456), .b(N5457), .O(N6177) );
inv1 gate1586( .a(N5114), .O(N6181) );
inv1 gate1587( .a(N5117), .O(N6182) );
inv1 gate1588( .a(N5120), .O(N6183) );
inv1 gate1589( .a(N5123), .O(N6184) );
inv1 gate1590( .a(N5138), .O(N6185) );
nand2 gate1591( .a(N5138), .b(N4783), .O(N6186) );
inv1 gate1592( .a(N5141), .O(N6187) );
inv1 gate1593( .a(N5144), .O(N6188) );
inv1 gate1594( .a(N5147), .O(N6189) );
inv1 gate1595( .a(N5150), .O(N6190) );
inv1 gate1596( .a(N4784), .O(N6191) );
nand2 gate1597( .a(N4784), .b(N2230), .O(N6192) );
inv1 gate1598( .a(N4790), .O(N6193) );
nand2 gate1599( .a(N4790), .b(N2765), .O(N6194) );
inv1 gate1600( .a(N4796), .O(N6195) );
nand2 gate1601( .a(N5476), .b(N5477), .O(N6196) );
nand2 gate1602( .a(N5474), .b(N5475), .O(N6199) );
inv1 gate1603( .a(N4810), .O(N6202) );
inv1 gate1604( .a(N4814), .O(N6203) );
buf1 gate1605( .a(N4769), .O(N6204) );
buf1 gate1606( .a(N4555), .O(N6207) );
buf1 gate1607( .a(N4769), .O(N6210) );
inv1 gate1608( .a(N4871), .O(N6213) );
buf1 gate1609( .a(N4586), .O(N6214) );

  xor2  gate3948(.a(N4769), .b(N2674), .O(gate1610inter0));
  nand2 gate3949(.a(gate1610inter0), .b(s_62), .O(gate1610inter1));
  and2  gate3950(.a(N4769), .b(N2674), .O(gate1610inter2));
  inv1  gate3951(.a(s_62), .O(gate1610inter3));
  inv1  gate3952(.a(s_63), .O(gate1610inter4));
  nand2 gate3953(.a(gate1610inter4), .b(gate1610inter3), .O(gate1610inter5));
  nor2  gate3954(.a(gate1610inter5), .b(gate1610inter2), .O(gate1610inter6));
  inv1  gate3955(.a(N2674), .O(gate1610inter7));
  inv1  gate3956(.a(N4769), .O(gate1610inter8));
  nand2 gate3957(.a(gate1610inter8), .b(gate1610inter7), .O(gate1610inter9));
  nand2 gate3958(.a(s_63), .b(gate1610inter3), .O(gate1610inter10));
  nor2  gate3959(.a(gate1610inter10), .b(gate1610inter9), .O(gate1610inter11));
  nor2  gate3960(.a(gate1610inter11), .b(gate1610inter6), .O(gate1610inter12));
  nand2 gate3961(.a(gate1610inter12), .b(gate1610inter1), .O(N6217));
buf1 gate1611( .a(N4667), .O(N6220) );
inv1 gate1612( .a(N4958), .O(N6223) );
inv1 gate1613( .a(N4961), .O(N6224) );
inv1 gate1614( .a(N4964), .O(N6225) );
inv1 gate1615( .a(N4967), .O(N6226) );
inv1 gate1616( .a(N4985), .O(N6227) );
inv1 gate1617( .a(N4988), .O(N6228) );
inv1 gate1618( .a(N4991), .O(N6229) );
inv1 gate1619( .a(N4994), .O(N6230) );
inv1 gate1620( .a(N5027), .O(N6231) );
buf1 gate1621( .a(N4711), .O(N6232) );
inv1 gate1622( .a(N5030), .O(N6235) );
buf1 gate1623( .a(N4735), .O(N6236) );
inv1 gate1624( .a(N5052), .O(N6239) );
inv1 gate1625( .a(N5055), .O(N6240) );
inv1 gate1626( .a(N5058), .O(N6241) );
inv1 gate1627( .a(N5061), .O(N6242) );
nand2 gate1628( .a(N5573), .b(N5574), .O(N6243) );
nand2 gate1629( .a(N5571), .b(N5572), .O(N6246) );

  xor2  gate4830(.a(N5587), .b(N5586), .O(gate1630inter0));
  nand2 gate4831(.a(gate1630inter0), .b(s_188), .O(gate1630inter1));
  and2  gate4832(.a(N5587), .b(N5586), .O(gate1630inter2));
  inv1  gate4833(.a(s_188), .O(gate1630inter3));
  inv1  gate4834(.a(s_189), .O(gate1630inter4));
  nand2 gate4835(.a(gate1630inter4), .b(gate1630inter3), .O(gate1630inter5));
  nor2  gate4836(.a(gate1630inter5), .b(gate1630inter2), .O(gate1630inter6));
  inv1  gate4837(.a(N5586), .O(gate1630inter7));
  inv1  gate4838(.a(N5587), .O(gate1630inter8));
  nand2 gate4839(.a(gate1630inter8), .b(gate1630inter7), .O(gate1630inter9));
  nand2 gate4840(.a(s_189), .b(gate1630inter3), .O(gate1630inter10));
  nor2  gate4841(.a(gate1630inter10), .b(gate1630inter9), .O(gate1630inter11));
  nor2  gate4842(.a(gate1630inter11), .b(gate1630inter6), .O(gate1630inter12));
  nand2 gate4843(.a(gate1630inter12), .b(gate1630inter1), .O(N6249));
nand2 gate1631( .a(N5584), .b(N5585), .O(N6252) );
inv1 gate1632( .a(N5126), .O(N6255) );
inv1 gate1633( .a(N5129), .O(N6256) );
inv1 gate1634( .a(N5132), .O(N6257) );
inv1 gate1635( .a(N5135), .O(N6258) );
inv1 gate1636( .a(N5153), .O(N6259) );
inv1 gate1637( .a(N5156), .O(N6260) );
inv1 gate1638( .a(N5159), .O(N6261) );
inv1 gate1639( .a(N5162), .O(N6262) );
nand2 gate1640( .a(N5604), .b(N5605), .O(N6263) );
nand2 gate1641( .a(N5602), .b(N5603), .O(N6266) );
nand2 gate1642( .a(N1380), .b(N5945), .O(N6540) );

  xor2  gate4284(.a(N5947), .b(N1383), .O(gate1643inter0));
  nand2 gate4285(.a(gate1643inter0), .b(s_110), .O(gate1643inter1));
  and2  gate4286(.a(N5947), .b(N1383), .O(gate1643inter2));
  inv1  gate4287(.a(s_110), .O(gate1643inter3));
  inv1  gate4288(.a(s_111), .O(gate1643inter4));
  nand2 gate4289(.a(gate1643inter4), .b(gate1643inter3), .O(gate1643inter5));
  nor2  gate4290(.a(gate1643inter5), .b(gate1643inter2), .O(gate1643inter6));
  inv1  gate4291(.a(N1383), .O(gate1643inter7));
  inv1  gate4292(.a(N5947), .O(gate1643inter8));
  nand2 gate4293(.a(gate1643inter8), .b(gate1643inter7), .O(gate1643inter9));
  nand2 gate4294(.a(s_111), .b(gate1643inter3), .O(gate1643inter10));
  nor2  gate4295(.a(gate1643inter10), .b(gate1643inter9), .O(gate1643inter11));
  nor2  gate4296(.a(gate1643inter11), .b(gate1643inter6), .O(gate1643inter12));
  nand2 gate4297(.a(gate1643inter12), .b(gate1643inter1), .O(N6541));
nand2 gate1644( .a(N1386), .b(N5949), .O(N6542) );
nand2 gate1645( .a(N1389), .b(N5951), .O(N6543) );
nand2 gate1646( .a(N1392), .b(N5953), .O(N6544) );
nand2 gate1647( .a(N1395), .b(N5955), .O(N6545) );
nand2 gate1648( .a(N1398), .b(N5957), .O(N6546) );

  xor2  gate4662(.a(N5959), .b(N1401), .O(gate1649inter0));
  nand2 gate4663(.a(gate1649inter0), .b(s_164), .O(gate1649inter1));
  and2  gate4664(.a(N5959), .b(N1401), .O(gate1649inter2));
  inv1  gate4665(.a(s_164), .O(gate1649inter3));
  inv1  gate4666(.a(s_165), .O(gate1649inter4));
  nand2 gate4667(.a(gate1649inter4), .b(gate1649inter3), .O(gate1649inter5));
  nor2  gate4668(.a(gate1649inter5), .b(gate1649inter2), .O(gate1649inter6));
  inv1  gate4669(.a(N1401), .O(gate1649inter7));
  inv1  gate4670(.a(N5959), .O(gate1649inter8));
  nand2 gate4671(.a(gate1649inter8), .b(gate1649inter7), .O(gate1649inter9));
  nand2 gate4672(.a(s_165), .b(gate1649inter3), .O(gate1649inter10));
  nor2  gate4673(.a(gate1649inter10), .b(gate1649inter9), .O(gate1649inter11));
  nor2  gate4674(.a(gate1649inter11), .b(gate1649inter6), .O(gate1649inter12));
  nand2 gate4675(.a(gate1649inter12), .b(gate1649inter1), .O(N6547));
nand2 gate1650( .a(N1404), .b(N5968), .O(N6555) );
nand2 gate1651( .a(N1407), .b(N5970), .O(N6556) );

  xor2  gate4368(.a(N5972), .b(N1410), .O(gate1652inter0));
  nand2 gate4369(.a(gate1652inter0), .b(s_122), .O(gate1652inter1));
  and2  gate4370(.a(N5972), .b(N1410), .O(gate1652inter2));
  inv1  gate4371(.a(s_122), .O(gate1652inter3));
  inv1  gate4372(.a(s_123), .O(gate1652inter4));
  nand2 gate4373(.a(gate1652inter4), .b(gate1652inter3), .O(gate1652inter5));
  nor2  gate4374(.a(gate1652inter5), .b(gate1652inter2), .O(gate1652inter6));
  inv1  gate4375(.a(N1410), .O(gate1652inter7));
  inv1  gate4376(.a(N5972), .O(gate1652inter8));
  nand2 gate4377(.a(gate1652inter8), .b(gate1652inter7), .O(gate1652inter9));
  nand2 gate4378(.a(s_123), .b(gate1652inter3), .O(gate1652inter10));
  nor2  gate4379(.a(gate1652inter10), .b(gate1652inter9), .O(gate1652inter11));
  nor2  gate4380(.a(gate1652inter11), .b(gate1652inter6), .O(gate1652inter12));
  nand2 gate4381(.a(gate1652inter12), .b(gate1652inter1), .O(N6557));
nand2 gate1653( .a(N1413), .b(N5974), .O(N6558) );
nand2 gate1654( .a(N1416), .b(N5976), .O(N6559) );

  xor2  gate4788(.a(N5978), .b(N1419), .O(gate1655inter0));
  nand2 gate4789(.a(gate1655inter0), .b(s_182), .O(gate1655inter1));
  and2  gate4790(.a(N5978), .b(N1419), .O(gate1655inter2));
  inv1  gate4791(.a(s_182), .O(gate1655inter3));
  inv1  gate4792(.a(s_183), .O(gate1655inter4));
  nand2 gate4793(.a(gate1655inter4), .b(gate1655inter3), .O(gate1655inter5));
  nor2  gate4794(.a(gate1655inter5), .b(gate1655inter2), .O(gate1655inter6));
  inv1  gate4795(.a(N1419), .O(gate1655inter7));
  inv1  gate4796(.a(N5978), .O(gate1655inter8));
  nand2 gate4797(.a(gate1655inter8), .b(gate1655inter7), .O(gate1655inter9));
  nand2 gate4798(.a(s_183), .b(gate1655inter3), .O(gate1655inter10));
  nor2  gate4799(.a(gate1655inter10), .b(gate1655inter9), .O(gate1655inter11));
  nor2  gate4800(.a(gate1655inter11), .b(gate1655inter6), .O(gate1655inter12));
  nand2 gate4801(.a(gate1655inter12), .b(gate1655inter1), .O(N6560));
nand2 gate1656( .a(N1422), .b(N5980), .O(N6561) );
nand2 gate1657( .a(N1425), .b(N5990), .O(N6569) );
nand2 gate1658( .a(N3721), .b(N6023), .O(N6594) );
nand2 gate1659( .a(N3724), .b(N6025), .O(N6595) );
nand2 gate1660( .a(N3727), .b(N6027), .O(N6596) );
nand2 gate1661( .a(N3730), .b(N6029), .O(N6597) );
nand2 gate1662( .a(N4889), .b(N6031), .O(N6598) );
nand2 gate1663( .a(N4886), .b(N6032), .O(N6599) );
nand2 gate1664( .a(N4895), .b(N6033), .O(N6600) );
nand2 gate1665( .a(N4892), .b(N6034), .O(N6601) );
nand2 gate1666( .a(N4901), .b(N6035), .O(N6602) );
nand2 gate1667( .a(N4898), .b(N6036), .O(N6603) );
nand2 gate1668( .a(N3733), .b(N6037), .O(N6604) );

  xor2  gate3584(.a(N6039), .b(N4910), .O(gate1669inter0));
  nand2 gate3585(.a(gate1669inter0), .b(s_10), .O(gate1669inter1));
  and2  gate3586(.a(N6039), .b(N4910), .O(gate1669inter2));
  inv1  gate3587(.a(s_10), .O(gate1669inter3));
  inv1  gate3588(.a(s_11), .O(gate1669inter4));
  nand2 gate3589(.a(gate1669inter4), .b(gate1669inter3), .O(gate1669inter5));
  nor2  gate3590(.a(gate1669inter5), .b(gate1669inter2), .O(gate1669inter6));
  inv1  gate3591(.a(N4910), .O(gate1669inter7));
  inv1  gate3592(.a(N6039), .O(gate1669inter8));
  nand2 gate3593(.a(gate1669inter8), .b(gate1669inter7), .O(gate1669inter9));
  nand2 gate3594(.a(s_11), .b(gate1669inter3), .O(gate1669inter10));
  nor2  gate3595(.a(gate1669inter10), .b(gate1669inter9), .O(gate1669inter11));
  nor2  gate3596(.a(gate1669inter11), .b(gate1669inter6), .O(gate1669inter12));
  nand2 gate3597(.a(gate1669inter12), .b(gate1669inter1), .O(N6605));
nand2 gate1670( .a(N4907), .b(N6040), .O(N6606) );
nand2 gate1671( .a(N1434), .b(N6061), .O(N6621) );

  xor2  gate4144(.a(N6063), .b(N1437), .O(gate1672inter0));
  nand2 gate4145(.a(gate1672inter0), .b(s_90), .O(gate1672inter1));
  and2  gate4146(.a(N6063), .b(N1437), .O(gate1672inter2));
  inv1  gate4147(.a(s_90), .O(gate1672inter3));
  inv1  gate4148(.a(s_91), .O(gate1672inter4));
  nand2 gate4149(.a(gate1672inter4), .b(gate1672inter3), .O(gate1672inter5));
  nor2  gate4150(.a(gate1672inter5), .b(gate1672inter2), .O(gate1672inter6));
  inv1  gate4151(.a(N1437), .O(gate1672inter7));
  inv1  gate4152(.a(N6063), .O(gate1672inter8));
  nand2 gate4153(.a(gate1672inter8), .b(gate1672inter7), .O(gate1672inter9));
  nand2 gate4154(.a(s_91), .b(gate1672inter3), .O(gate1672inter10));
  nor2  gate4155(.a(gate1672inter10), .b(gate1672inter9), .O(gate1672inter11));
  nor2  gate4156(.a(gate1672inter11), .b(gate1672inter6), .O(gate1672inter12));
  nand2 gate4157(.a(gate1672inter12), .b(gate1672inter1), .O(N6622));
nand2 gate1673( .a(N1440), .b(N6065), .O(N6623) );

  xor2  gate4424(.a(N6067), .b(N1443), .O(gate1674inter0));
  nand2 gate4425(.a(gate1674inter0), .b(s_130), .O(gate1674inter1));
  and2  gate4426(.a(N6067), .b(N1443), .O(gate1674inter2));
  inv1  gate4427(.a(s_130), .O(gate1674inter3));
  inv1  gate4428(.a(s_131), .O(gate1674inter4));
  nand2 gate4429(.a(gate1674inter4), .b(gate1674inter3), .O(gate1674inter5));
  nor2  gate4430(.a(gate1674inter5), .b(gate1674inter2), .O(gate1674inter6));
  inv1  gate4431(.a(N1443), .O(gate1674inter7));
  inv1  gate4432(.a(N6067), .O(gate1674inter8));
  nand2 gate4433(.a(gate1674inter8), .b(gate1674inter7), .O(gate1674inter9));
  nand2 gate4434(.a(s_131), .b(gate1674inter3), .O(gate1674inter10));
  nor2  gate4435(.a(gate1674inter10), .b(gate1674inter9), .O(gate1674inter11));
  nor2  gate4436(.a(gate1674inter11), .b(gate1674inter6), .O(gate1674inter12));
  nand2 gate4437(.a(gate1674inter12), .b(gate1674inter1), .O(N6624));
nand2 gate1675( .a(N1446), .b(N6069), .O(N6625) );
nand2 gate1676( .a(N1449), .b(N6071), .O(N6626) );
nand2 gate1677( .a(N1452), .b(N6073), .O(N6627) );
nand2 gate1678( .a(N1455), .b(N6075), .O(N6628) );
nand2 gate1679( .a(N1458), .b(N6077), .O(N6629) );
nand2 gate1680( .a(N3783), .b(N6090), .O(N6639) );
nand2 gate1681( .a(N4949), .b(N6092), .O(N6640) );
nand2 gate1682( .a(N4946), .b(N6093), .O(N6641) );
nand2 gate1683( .a(N4955), .b(N6094), .O(N6642) );
nand2 gate1684( .a(N4952), .b(N6095), .O(N6643) );
nand2 gate1685( .a(N3786), .b(N6096), .O(N6644) );
nand2 gate1686( .a(N4976), .b(N6098), .O(N6645) );

  xor2  gate3696(.a(N6099), .b(N4973), .O(gate1687inter0));
  nand2 gate3697(.a(gate1687inter0), .b(s_26), .O(gate1687inter1));
  and2  gate3698(.a(N6099), .b(N4973), .O(gate1687inter2));
  inv1  gate3699(.a(s_26), .O(gate1687inter3));
  inv1  gate3700(.a(s_27), .O(gate1687inter4));
  nand2 gate3701(.a(gate1687inter4), .b(gate1687inter3), .O(gate1687inter5));
  nor2  gate3702(.a(gate1687inter5), .b(gate1687inter2), .O(gate1687inter6));
  inv1  gate3703(.a(N4973), .O(gate1687inter7));
  inv1  gate3704(.a(N6099), .O(gate1687inter8));
  nand2 gate3705(.a(gate1687inter8), .b(gate1687inter7), .O(gate1687inter9));
  nand2 gate3706(.a(s_27), .b(gate1687inter3), .O(gate1687inter10));
  nor2  gate3707(.a(gate1687inter10), .b(gate1687inter9), .O(gate1687inter11));
  nor2  gate3708(.a(gate1687inter11), .b(gate1687inter6), .O(gate1687inter12));
  nand2 gate3709(.a(gate1687inter12), .b(gate1687inter1), .O(N6646));
nand2 gate1688( .a(N4982), .b(N6100), .O(N6647) );
nand2 gate1689( .a(N4979), .b(N6101), .O(N6648) );

  xor2  gate4480(.a(N6104), .b(N1461), .O(gate1690inter0));
  nand2 gate4481(.a(gate1690inter0), .b(s_138), .O(gate1690inter1));
  and2  gate4482(.a(N6104), .b(N1461), .O(gate1690inter2));
  inv1  gate4483(.a(s_138), .O(gate1690inter3));
  inv1  gate4484(.a(s_139), .O(gate1690inter4));
  nand2 gate4485(.a(gate1690inter4), .b(gate1690inter3), .O(gate1690inter5));
  nor2  gate4486(.a(gate1690inter5), .b(gate1690inter2), .O(gate1690inter6));
  inv1  gate4487(.a(N1461), .O(gate1690inter7));
  inv1  gate4488(.a(N6104), .O(gate1690inter8));
  nand2 gate4489(.a(gate1690inter8), .b(gate1690inter7), .O(gate1690inter9));
  nand2 gate4490(.a(s_139), .b(gate1690inter3), .O(gate1690inter10));
  nor2  gate4491(.a(gate1690inter10), .b(gate1690inter9), .O(gate1690inter11));
  nor2  gate4492(.a(gate1690inter11), .b(gate1690inter6), .O(gate1690inter12));
  nand2 gate4493(.a(gate1690inter12), .b(gate1690inter1), .O(N6649));
nand2 gate1691( .a(N1464), .b(N6106), .O(N6650) );
nand2 gate1692( .a(N1467), .b(N6108), .O(N6651) );
nand2 gate1693( .a(N1470), .b(N6110), .O(N6652) );
nand2 gate1694( .a(N1473), .b(N6112), .O(N6653) );
nand2 gate1695( .a(N1476), .b(N6114), .O(N6654) );
nand2 gate1696( .a(N1479), .b(N6116), .O(N6655) );
nand2 gate1697( .a(N1482), .b(N6118), .O(N6656) );
nand2 gate1698( .a(N1485), .b(N6120), .O(N6657) );
nand2 gate1699( .a(N3789), .b(N6121), .O(N6658) );
nand2 gate1700( .a(N5039), .b(N6123), .O(N6659) );
nand2 gate1701( .a(N5036), .b(N6124), .O(N6660) );
nand2 gate1702( .a(N3792), .b(N6126), .O(N6661) );
nand2 gate1703( .a(N3816), .b(N6135), .O(N6668) );
nand2 gate1704( .a(N5071), .b(N6148), .O(N6677) );
nand2 gate1705( .a(N5068), .b(N6149), .O(N6678) );
nand2 gate1706( .a(N5077), .b(N6150), .O(N6679) );
nand2 gate1707( .a(N5074), .b(N6151), .O(N6680) );
nand2 gate1708( .a(N5083), .b(N6152), .O(N6681) );
nand2 gate1709( .a(N5080), .b(N6153), .O(N6682) );
nand2 gate1710( .a(N5089), .b(N6154), .O(N6683) );
nand2 gate1711( .a(N5086), .b(N6155), .O(N6684) );
nand2 gate1712( .a(N3846), .b(N6156), .O(N6685) );
nand2 gate1713( .a(N3849), .b(N6158), .O(N6686) );
nand2 gate1714( .a(N3852), .b(N6160), .O(N6687) );
nand2 gate1715( .a(N5104), .b(N6162), .O(N6688) );
nand2 gate1716( .a(N5101), .b(N6163), .O(N6689) );
nand2 gate1717( .a(N3855), .b(N6165), .O(N6690) );
nand2 gate1718( .a(N5117), .b(N6181), .O(N6702) );
nand2 gate1719( .a(N5114), .b(N6182), .O(N6703) );
nand2 gate1720( .a(N5123), .b(N6183), .O(N6704) );
nand2 gate1721( .a(N5120), .b(N6184), .O(N6705) );
nand2 gate1722( .a(N3891), .b(N6185), .O(N6706) );
nand2 gate1723( .a(N5144), .b(N6187), .O(N6707) );
nand2 gate1724( .a(N5141), .b(N6188), .O(N6708) );
nand2 gate1725( .a(N5150), .b(N6189), .O(N6709) );

  xor2  gate5264(.a(N6190), .b(N5147), .O(gate1726inter0));
  nand2 gate5265(.a(gate1726inter0), .b(s_250), .O(gate1726inter1));
  and2  gate5266(.a(N6190), .b(N5147), .O(gate1726inter2));
  inv1  gate5267(.a(s_250), .O(gate1726inter3));
  inv1  gate5268(.a(s_251), .O(gate1726inter4));
  nand2 gate5269(.a(gate1726inter4), .b(gate1726inter3), .O(gate1726inter5));
  nor2  gate5270(.a(gate1726inter5), .b(gate1726inter2), .O(gate1726inter6));
  inv1  gate5271(.a(N5147), .O(gate1726inter7));
  inv1  gate5272(.a(N6190), .O(gate1726inter8));
  nand2 gate5273(.a(gate1726inter8), .b(gate1726inter7), .O(gate1726inter9));
  nand2 gate5274(.a(s_251), .b(gate1726inter3), .O(gate1726inter10));
  nor2  gate5275(.a(gate1726inter10), .b(gate1726inter9), .O(gate1726inter11));
  nor2  gate5276(.a(gate1726inter11), .b(gate1726inter6), .O(gate1726inter12));
  nand2 gate5277(.a(gate1726inter12), .b(gate1726inter1), .O(N6710));

  xor2  gate5096(.a(N6191), .b(N1708), .O(gate1727inter0));
  nand2 gate5097(.a(gate1727inter0), .b(s_226), .O(gate1727inter1));
  and2  gate5098(.a(N6191), .b(N1708), .O(gate1727inter2));
  inv1  gate5099(.a(s_226), .O(gate1727inter3));
  inv1  gate5100(.a(s_227), .O(gate1727inter4));
  nand2 gate5101(.a(gate1727inter4), .b(gate1727inter3), .O(gate1727inter5));
  nor2  gate5102(.a(gate1727inter5), .b(gate1727inter2), .O(gate1727inter6));
  inv1  gate5103(.a(N1708), .O(gate1727inter7));
  inv1  gate5104(.a(N6191), .O(gate1727inter8));
  nand2 gate5105(.a(gate1727inter8), .b(gate1727inter7), .O(gate1727inter9));
  nand2 gate5106(.a(s_227), .b(gate1727inter3), .O(gate1727inter10));
  nor2  gate5107(.a(gate1727inter10), .b(gate1727inter9), .O(gate1727inter11));
  nor2  gate5108(.a(gate1727inter11), .b(gate1727inter6), .O(gate1727inter12));
  nand2 gate5109(.a(gate1727inter12), .b(gate1727inter1), .O(N6711));
nand2 gate1728( .a(N2231), .b(N6193), .O(N6712) );
nand2 gate1729( .a(N4961), .b(N6223), .O(N6729) );

  xor2  gate4172(.a(N6224), .b(N4958), .O(gate1730inter0));
  nand2 gate4173(.a(gate1730inter0), .b(s_94), .O(gate1730inter1));
  and2  gate4174(.a(N6224), .b(N4958), .O(gate1730inter2));
  inv1  gate4175(.a(s_94), .O(gate1730inter3));
  inv1  gate4176(.a(s_95), .O(gate1730inter4));
  nand2 gate4177(.a(gate1730inter4), .b(gate1730inter3), .O(gate1730inter5));
  nor2  gate4178(.a(gate1730inter5), .b(gate1730inter2), .O(gate1730inter6));
  inv1  gate4179(.a(N4958), .O(gate1730inter7));
  inv1  gate4180(.a(N6224), .O(gate1730inter8));
  nand2 gate4181(.a(gate1730inter8), .b(gate1730inter7), .O(gate1730inter9));
  nand2 gate4182(.a(s_95), .b(gate1730inter3), .O(gate1730inter10));
  nor2  gate4183(.a(gate1730inter10), .b(gate1730inter9), .O(gate1730inter11));
  nor2  gate4184(.a(gate1730inter11), .b(gate1730inter6), .O(gate1730inter12));
  nand2 gate4185(.a(gate1730inter12), .b(gate1730inter1), .O(N6730));
nand2 gate1731( .a(N4967), .b(N6225), .O(N6731) );
nand2 gate1732( .a(N4964), .b(N6226), .O(N6732) );
nand2 gate1733( .a(N4988), .b(N6227), .O(N6733) );
nand2 gate1734( .a(N4985), .b(N6228), .O(N6734) );
nand2 gate1735( .a(N4994), .b(N6229), .O(N6735) );
nand2 gate1736( .a(N4991), .b(N6230), .O(N6736) );
nand2 gate1737( .a(N5055), .b(N6239), .O(N6741) );
nand2 gate1738( .a(N5052), .b(N6240), .O(N6742) );
nand2 gate1739( .a(N5061), .b(N6241), .O(N6743) );

  xor2  gate4410(.a(N6242), .b(N5058), .O(gate1740inter0));
  nand2 gate4411(.a(gate1740inter0), .b(s_128), .O(gate1740inter1));
  and2  gate4412(.a(N6242), .b(N5058), .O(gate1740inter2));
  inv1  gate4413(.a(s_128), .O(gate1740inter3));
  inv1  gate4414(.a(s_129), .O(gate1740inter4));
  nand2 gate4415(.a(gate1740inter4), .b(gate1740inter3), .O(gate1740inter5));
  nor2  gate4416(.a(gate1740inter5), .b(gate1740inter2), .O(gate1740inter6));
  inv1  gate4417(.a(N5058), .O(gate1740inter7));
  inv1  gate4418(.a(N6242), .O(gate1740inter8));
  nand2 gate4419(.a(gate1740inter8), .b(gate1740inter7), .O(gate1740inter9));
  nand2 gate4420(.a(s_129), .b(gate1740inter3), .O(gate1740inter10));
  nor2  gate4421(.a(gate1740inter10), .b(gate1740inter9), .O(gate1740inter11));
  nor2  gate4422(.a(gate1740inter11), .b(gate1740inter6), .O(gate1740inter12));
  nand2 gate4423(.a(gate1740inter12), .b(gate1740inter1), .O(N6744));
nand2 gate1741( .a(N5129), .b(N6255), .O(N6751) );
nand2 gate1742( .a(N5126), .b(N6256), .O(N6752) );
nand2 gate1743( .a(N5135), .b(N6257), .O(N6753) );

  xor2  gate4018(.a(N6258), .b(N5132), .O(gate1744inter0));
  nand2 gate4019(.a(gate1744inter0), .b(s_72), .O(gate1744inter1));
  and2  gate4020(.a(N6258), .b(N5132), .O(gate1744inter2));
  inv1  gate4021(.a(s_72), .O(gate1744inter3));
  inv1  gate4022(.a(s_73), .O(gate1744inter4));
  nand2 gate4023(.a(gate1744inter4), .b(gate1744inter3), .O(gate1744inter5));
  nor2  gate4024(.a(gate1744inter5), .b(gate1744inter2), .O(gate1744inter6));
  inv1  gate4025(.a(N5132), .O(gate1744inter7));
  inv1  gate4026(.a(N6258), .O(gate1744inter8));
  nand2 gate4027(.a(gate1744inter8), .b(gate1744inter7), .O(gate1744inter9));
  nand2 gate4028(.a(s_73), .b(gate1744inter3), .O(gate1744inter10));
  nor2  gate4029(.a(gate1744inter10), .b(gate1744inter9), .O(gate1744inter11));
  nor2  gate4030(.a(gate1744inter11), .b(gate1744inter6), .O(gate1744inter12));
  nand2 gate4031(.a(gate1744inter12), .b(gate1744inter1), .O(N6754));
nand2 gate1745( .a(N5156), .b(N6259), .O(N6755) );
nand2 gate1746( .a(N5153), .b(N6260), .O(N6756) );
nand2 gate1747( .a(N5162), .b(N6261), .O(N6757) );
nand2 gate1748( .a(N5159), .b(N6262), .O(N6758) );
inv1 gate1749( .a(N5892), .O(N6761) );
and5 gate1750( .a(N5683), .b(N5670), .c(N5654), .d(N5640), .e(N5632), .O(N6762) );
and2 gate1751( .a(N5632), .b(N3097), .O(N6766) );
and3 gate1752( .a(N5640), .b(N5632), .c(N3101), .O(N6767) );
and4 gate1753( .a(N5654), .b(N5632), .c(N3107), .d(N5640), .O(N6768) );
and5 gate1754( .a(N5670), .b(N5654), .c(N5632), .d(N3114), .e(N5640), .O(N6769) );
and2 gate1755( .a(N5640), .b(N3101), .O(N6770) );
and3 gate1756( .a(N5654), .b(N3107), .c(N5640), .O(N6771) );
and4 gate1757( .a(N5670), .b(N5654), .c(N3114), .d(N5640), .O(N6772) );
and4 gate1758( .a(N5683), .b(N5654), .c(N5640), .d(N5670), .O(N6773) );
and2 gate1759( .a(N5640), .b(N3101), .O(N6774) );
and3 gate1760( .a(N5654), .b(N3107), .c(N5640), .O(N6775) );
and4 gate1761( .a(N5670), .b(N5654), .c(N3114), .d(N5640), .O(N6776) );
and2 gate1762( .a(N5654), .b(N3107), .O(N6777) );
and3 gate1763( .a(N5670), .b(N5654), .c(N3114), .O(N6778) );
and3 gate1764( .a(N5683), .b(N5654), .c(N5670), .O(N6779) );
and2 gate1765( .a(N5654), .b(N3107), .O(N6780) );
and3 gate1766( .a(N5670), .b(N5654), .c(N3114), .O(N6781) );
and2 gate1767( .a(N5670), .b(N3114), .O(N6782) );
and2 gate1768( .a(N5683), .b(N5670), .O(N6783) );
and5 gate1769( .a(N5697), .b(N5728), .c(N5707), .d(N5690), .e(N5718), .O(N6784) );
and2 gate1770( .a(N5690), .b(N3137), .O(N6787) );
and3 gate1771( .a(N5697), .b(N5690), .c(N3140), .O(N6788) );
and4 gate1772( .a(N5707), .b(N5690), .c(N3144), .d(N5697), .O(N6789) );
and5 gate1773( .a(N5718), .b(N5707), .c(N5690), .d(N3149), .e(N5697), .O(N6790) );
and2 gate1774( .a(N5697), .b(N3140), .O(N6791) );
and3 gate1775( .a(N5707), .b(N3144), .c(N5697), .O(N6792) );
and4 gate1776( .a(N5718), .b(N5707), .c(N3149), .d(N5697), .O(N6793) );
and2 gate1777( .a(N3144), .b(N5707), .O(N6794) );
and3 gate1778( .a(N5718), .b(N5707), .c(N3149), .O(N6795) );
and2 gate1779( .a(N5718), .b(N3149), .O(N6796) );
inv1 gate1780( .a(N5736), .O(N6797) );
inv1 gate1781( .a(N5740), .O(N6800) );
inv1 gate1782( .a(N5747), .O(N6803) );
inv1 gate1783( .a(N5751), .O(N6806) );
inv1 gate1784( .a(N5758), .O(N6809) );
inv1 gate1785( .a(N5762), .O(N6812) );
buf1 gate1786( .a(N5744), .O(N6815) );
buf1 gate1787( .a(N5744), .O(N6818) );
buf1 gate1788( .a(N5755), .O(N6821) );
buf1 gate1789( .a(N5755), .O(N6824) );
buf1 gate1790( .a(N5766), .O(N6827) );
buf1 gate1791( .a(N5766), .O(N6830) );
and4 gate1792( .a(N5850), .b(N5789), .c(N5778), .d(N5771), .O(N6833) );
and2 gate1793( .a(N5771), .b(N3169), .O(N6836) );
and3 gate1794( .a(N5778), .b(N5771), .c(N3173), .O(N6837) );
and4 gate1795( .a(N5789), .b(N5771), .c(N3178), .d(N5778), .O(N6838) );
and2 gate1796( .a(N5778), .b(N3173), .O(N6839) );
and3 gate1797( .a(N5789), .b(N3178), .c(N5778), .O(N6840) );
and3 gate1798( .a(N5850), .b(N5789), .c(N5778), .O(N6841) );
and2 gate1799( .a(N5778), .b(N3173), .O(N6842) );
and3 gate1800( .a(N5789), .b(N3178), .c(N5778), .O(N6843) );
and2 gate1801( .a(N5789), .b(N3178), .O(N6844) );
and5 gate1802( .a(N5856), .b(N5837), .c(N5821), .d(N5807), .e(N5799), .O(N6845) );
and2 gate1803( .a(N5799), .b(N3185), .O(N6848) );
and3 gate1804( .a(N5807), .b(N5799), .c(N3189), .O(N6849) );
and4 gate1805( .a(N5821), .b(N5799), .c(N3195), .d(N5807), .O(N6850) );
and5 gate1806( .a(N5837), .b(N5821), .c(N5799), .d(N3202), .e(N5807), .O(N6851) );
and2 gate1807( .a(N5807), .b(N3189), .O(N6852) );
and3 gate1808( .a(N5821), .b(N3195), .c(N5807), .O(N6853) );
and4 gate1809( .a(N5837), .b(N5821), .c(N3202), .d(N5807), .O(N6854) );
and4 gate1810( .a(N5856), .b(N5821), .c(N5807), .d(N5837), .O(N6855) );
and2 gate1811( .a(N5807), .b(N3189), .O(N6856) );
and3 gate1812( .a(N5821), .b(N3195), .c(N5807), .O(N6857) );
and4 gate1813( .a(N5837), .b(N5821), .c(N3202), .d(N5807), .O(N6858) );
and2 gate1814( .a(N5821), .b(N3195), .O(N6859) );
and3 gate1815( .a(N5837), .b(N5821), .c(N3202), .O(N6860) );
and3 gate1816( .a(N5856), .b(N5821), .c(N5837), .O(N6861) );
and2 gate1817( .a(N5821), .b(N3195), .O(N6862) );
and3 gate1818( .a(N5837), .b(N5821), .c(N3202), .O(N6863) );
and2 gate1819( .a(N5837), .b(N3202), .O(N6864) );
and2 gate1820( .a(N5850), .b(N5789), .O(N6865) );
and2 gate1821( .a(N5856), .b(N5837), .O(N6866) );
and4 gate1822( .a(N5870), .b(N5892), .c(N5881), .d(N5863), .O(N6867) );
and2 gate1823( .a(N5863), .b(N3211), .O(N6870) );
and3 gate1824( .a(N5870), .b(N5863), .c(N3215), .O(N6871) );
and4 gate1825( .a(N5881), .b(N5863), .c(N3221), .d(N5870), .O(N6872) );
and2 gate1826( .a(N5870), .b(N3215), .O(N6873) );
and3 gate1827( .a(N5881), .b(N3221), .c(N5870), .O(N6874) );
and3 gate1828( .a(N5892), .b(N5881), .c(N5870), .O(N6875) );
and2 gate1829( .a(N5870), .b(N3215), .O(N6876) );
and3 gate1830( .a(N3221), .b(N5881), .c(N5870), .O(N6877) );
and2 gate1831( .a(N5881), .b(N3221), .O(N6878) );
and2 gate1832( .a(N5892), .b(N5881), .O(N6879) );
and2 gate1833( .a(N5881), .b(N3221), .O(N6880) );
and5 gate1834( .a(N5905), .b(N5936), .c(N5915), .d(N5898), .e(N5926), .O(N6881) );
and2 gate1835( .a(N5898), .b(N3229), .O(N6884) );
and3 gate1836( .a(N5905), .b(N5898), .c(N3232), .O(N6885) );
and4 gate1837( .a(N5915), .b(N5898), .c(N3236), .d(N5905), .O(N6886) );
and5 gate1838( .a(N5926), .b(N5915), .c(N5898), .d(N3241), .e(N5905), .O(N6887) );
and2 gate1839( .a(N5905), .b(N3232), .O(N6888) );
and3 gate1840( .a(N5915), .b(N3236), .c(N5905), .O(N6889) );
and4 gate1841( .a(N5926), .b(N5915), .c(N3241), .d(N5905), .O(N6890) );
and2 gate1842( .a(N3236), .b(N5915), .O(N6891) );
and3 gate1843( .a(N5926), .b(N5915), .c(N3241), .O(N6892) );
and2 gate1844( .a(N5926), .b(N3241), .O(N6893) );
nand2 gate1845( .a(N5944), .b(N6540), .O(N6894) );

  xor2  gate4074(.a(N6541), .b(N5946), .O(gate1846inter0));
  nand2 gate4075(.a(gate1846inter0), .b(s_80), .O(gate1846inter1));
  and2  gate4076(.a(N6541), .b(N5946), .O(gate1846inter2));
  inv1  gate4077(.a(s_80), .O(gate1846inter3));
  inv1  gate4078(.a(s_81), .O(gate1846inter4));
  nand2 gate4079(.a(gate1846inter4), .b(gate1846inter3), .O(gate1846inter5));
  nor2  gate4080(.a(gate1846inter5), .b(gate1846inter2), .O(gate1846inter6));
  inv1  gate4081(.a(N5946), .O(gate1846inter7));
  inv1  gate4082(.a(N6541), .O(gate1846inter8));
  nand2 gate4083(.a(gate1846inter8), .b(gate1846inter7), .O(gate1846inter9));
  nand2 gate4084(.a(s_81), .b(gate1846inter3), .O(gate1846inter10));
  nor2  gate4085(.a(gate1846inter10), .b(gate1846inter9), .O(gate1846inter11));
  nor2  gate4086(.a(gate1846inter11), .b(gate1846inter6), .O(gate1846inter12));
  nand2 gate4087(.a(gate1846inter12), .b(gate1846inter1), .O(N6901));
nand2 gate1847( .a(N5948), .b(N6542), .O(N6912) );
nand2 gate1848( .a(N5950), .b(N6543), .O(N6923) );
nand2 gate1849( .a(N5952), .b(N6544), .O(N6929) );
nand2 gate1850( .a(N5954), .b(N6545), .O(N6936) );
nand2 gate1851( .a(N5956), .b(N6546), .O(N6946) );
nand2 gate1852( .a(N5958), .b(N6547), .O(N6957) );
nand2 gate1853( .a(N6204), .b(N4575), .O(N6967) );
inv1 gate1854( .a(N6204), .O(N6968) );
inv1 gate1855( .a(N6207), .O(N6969) );
nand2 gate1856( .a(N5967), .b(N6555), .O(N6970) );
nand2 gate1857( .a(N5969), .b(N6556), .O(N6977) );
nand2 gate1858( .a(N5971), .b(N6557), .O(N6988) );

  xor2  gate5068(.a(N6558), .b(N5973), .O(gate1859inter0));
  nand2 gate5069(.a(gate1859inter0), .b(s_222), .O(gate1859inter1));
  and2  gate5070(.a(N6558), .b(N5973), .O(gate1859inter2));
  inv1  gate5071(.a(s_222), .O(gate1859inter3));
  inv1  gate5072(.a(s_223), .O(gate1859inter4));
  nand2 gate5073(.a(gate1859inter4), .b(gate1859inter3), .O(gate1859inter5));
  nor2  gate5074(.a(gate1859inter5), .b(gate1859inter2), .O(gate1859inter6));
  inv1  gate5075(.a(N5973), .O(gate1859inter7));
  inv1  gate5076(.a(N6558), .O(gate1859inter8));
  nand2 gate5077(.a(gate1859inter8), .b(gate1859inter7), .O(gate1859inter9));
  nand2 gate5078(.a(s_223), .b(gate1859inter3), .O(gate1859inter10));
  nor2  gate5079(.a(gate1859inter10), .b(gate1859inter9), .O(gate1859inter11));
  nor2  gate5080(.a(gate1859inter11), .b(gate1859inter6), .O(gate1859inter12));
  nand2 gate5081(.a(gate1859inter12), .b(gate1859inter1), .O(N6998));
nand2 gate1860( .a(N5975), .b(N6559), .O(N7006) );

  xor2  gate4004(.a(N6560), .b(N5977), .O(gate1861inter0));
  nand2 gate4005(.a(gate1861inter0), .b(s_70), .O(gate1861inter1));
  and2  gate4006(.a(N6560), .b(N5977), .O(gate1861inter2));
  inv1  gate4007(.a(s_70), .O(gate1861inter3));
  inv1  gate4008(.a(s_71), .O(gate1861inter4));
  nand2 gate4009(.a(gate1861inter4), .b(gate1861inter3), .O(gate1861inter5));
  nor2  gate4010(.a(gate1861inter5), .b(gate1861inter2), .O(gate1861inter6));
  inv1  gate4011(.a(N5977), .O(gate1861inter7));
  inv1  gate4012(.a(N6560), .O(gate1861inter8));
  nand2 gate4013(.a(gate1861inter8), .b(gate1861inter7), .O(gate1861inter9));
  nand2 gate4014(.a(s_71), .b(gate1861inter3), .O(gate1861inter10));
  nor2  gate4015(.a(gate1861inter10), .b(gate1861inter9), .O(gate1861inter11));
  nor2  gate4016(.a(gate1861inter11), .b(gate1861inter6), .O(gate1861inter12));
  nand2 gate4017(.a(gate1861inter12), .b(gate1861inter1), .O(N7020));
nand2 gate1862( .a(N5979), .b(N6561), .O(N7036) );
nand2 gate1863( .a(N5989), .b(N6569), .O(N7049) );
nand2 gate1864( .a(N6210), .b(N4610), .O(N7055) );
inv1 gate1865( .a(N6210), .O(N7056) );
and4 gate1866( .a(N6021), .b(N6000), .c(N5996), .d(N5991), .O(N7057) );
and2 gate1867( .a(N5991), .b(N3362), .O(N7060) );
and3 gate1868( .a(N5996), .b(N5991), .c(N3363), .O(N7061) );
and4 gate1869( .a(N6000), .b(N5991), .c(N3364), .d(N5996), .O(N7062) );
and5 gate1870( .a(N6022), .b(N6018), .c(N6014), .d(N6009), .e(N6003), .O(N7063) );
and2 gate1871( .a(N6003), .b(N3366), .O(N7064) );
and3 gate1872( .a(N6009), .b(N6003), .c(N3367), .O(N7065) );
and4 gate1873( .a(N6014), .b(N6003), .c(N3368), .d(N6009), .O(N7066) );
and5 gate1874( .a(N6018), .b(N6014), .c(N6003), .d(N3369), .e(N6009), .O(N7067) );
nand2 gate1875( .a(N6594), .b(N6024), .O(N7068) );
nand2 gate1876( .a(N6595), .b(N6026), .O(N7073) );
nand2 gate1877( .a(N6596), .b(N6028), .O(N7077) );
nand2 gate1878( .a(N6597), .b(N6030), .O(N7080) );

  xor2  gate4914(.a(N6599), .b(N6598), .O(gate1879inter0));
  nand2 gate4915(.a(gate1879inter0), .b(s_200), .O(gate1879inter1));
  and2  gate4916(.a(N6599), .b(N6598), .O(gate1879inter2));
  inv1  gate4917(.a(s_200), .O(gate1879inter3));
  inv1  gate4918(.a(s_201), .O(gate1879inter4));
  nand2 gate4919(.a(gate1879inter4), .b(gate1879inter3), .O(gate1879inter5));
  nor2  gate4920(.a(gate1879inter5), .b(gate1879inter2), .O(gate1879inter6));
  inv1  gate4921(.a(N6598), .O(gate1879inter7));
  inv1  gate4922(.a(N6599), .O(gate1879inter8));
  nand2 gate4923(.a(gate1879inter8), .b(gate1879inter7), .O(gate1879inter9));
  nand2 gate4924(.a(s_201), .b(gate1879inter3), .O(gate1879inter10));
  nor2  gate4925(.a(gate1879inter10), .b(gate1879inter9), .O(gate1879inter11));
  nor2  gate4926(.a(gate1879inter11), .b(gate1879inter6), .O(gate1879inter12));
  nand2 gate4927(.a(gate1879inter12), .b(gate1879inter1), .O(N7086));
nand2 gate1880( .a(N6600), .b(N6601), .O(N7091) );
nand2 gate1881( .a(N6602), .b(N6603), .O(N7095) );
nand2 gate1882( .a(N6604), .b(N6038), .O(N7098) );
nand2 gate1883( .a(N6605), .b(N6606), .O(N7099) );
and5 gate1884( .a(N6059), .b(N6056), .c(N6052), .d(N6047), .e(N6041), .O(N7100) );
and2 gate1885( .a(N6041), .b(N3371), .O(N7103) );
and3 gate1886( .a(N6047), .b(N6041), .c(N3372), .O(N7104) );
and4 gate1887( .a(N6052), .b(N6041), .c(N3373), .d(N6047), .O(N7105) );
and5 gate1888( .a(N6056), .b(N6052), .c(N6041), .d(N3374), .e(N6047), .O(N7106) );
nand2 gate1889( .a(N6060), .b(N6621), .O(N7107) );

  xor2  gate4382(.a(N6622), .b(N6062), .O(gate1890inter0));
  nand2 gate4383(.a(gate1890inter0), .b(s_124), .O(gate1890inter1));
  and2  gate4384(.a(N6622), .b(N6062), .O(gate1890inter2));
  inv1  gate4385(.a(s_124), .O(gate1890inter3));
  inv1  gate4386(.a(s_125), .O(gate1890inter4));
  nand2 gate4387(.a(gate1890inter4), .b(gate1890inter3), .O(gate1890inter5));
  nor2  gate4388(.a(gate1890inter5), .b(gate1890inter2), .O(gate1890inter6));
  inv1  gate4389(.a(N6062), .O(gate1890inter7));
  inv1  gate4390(.a(N6622), .O(gate1890inter8));
  nand2 gate4391(.a(gate1890inter8), .b(gate1890inter7), .O(gate1890inter9));
  nand2 gate4392(.a(s_125), .b(gate1890inter3), .O(gate1890inter10));
  nor2  gate4393(.a(gate1890inter10), .b(gate1890inter9), .O(gate1890inter11));
  nor2  gate4394(.a(gate1890inter11), .b(gate1890inter6), .O(gate1890inter12));
  nand2 gate4395(.a(gate1890inter12), .b(gate1890inter1), .O(N7114));
nand2 gate1891( .a(N6064), .b(N6623), .O(N7125) );
nand2 gate1892( .a(N6066), .b(N6624), .O(N7136) );
nand2 gate1893( .a(N6068), .b(N6625), .O(N7142) );
nand2 gate1894( .a(N6070), .b(N6626), .O(N7149) );
nand2 gate1895( .a(N6072), .b(N6627), .O(N7159) );
nand2 gate1896( .a(N6074), .b(N6628), .O(N7170) );
nand2 gate1897( .a(N6076), .b(N6629), .O(N7180) );
inv1 gate1898( .a(N6220), .O(N7187) );
inv1 gate1899( .a(N6079), .O(N7188) );
inv1 gate1900( .a(N6083), .O(N7191) );
nand2 gate1901( .a(N6639), .b(N6091), .O(N7194) );
nand2 gate1902( .a(N6640), .b(N6641), .O(N7198) );
nand2 gate1903( .a(N6642), .b(N6643), .O(N7202) );
nand2 gate1904( .a(N6644), .b(N6097), .O(N7205) );
nand2 gate1905( .a(N6645), .b(N6646), .O(N7209) );
nand2 gate1906( .a(N6647), .b(N6648), .O(N7213) );
buf1 gate1907( .a(N6087), .O(N7216) );
buf1 gate1908( .a(N6087), .O(N7219) );
nand2 gate1909( .a(N6103), .b(N6649), .O(N7222) );
nand2 gate1910( .a(N6105), .b(N6650), .O(N7229) );
nand2 gate1911( .a(N6107), .b(N6651), .O(N7240) );
nand2 gate1912( .a(N6109), .b(N6652), .O(N7250) );

  xor2  gate4228(.a(N6653), .b(N6111), .O(gate1913inter0));
  nand2 gate4229(.a(gate1913inter0), .b(s_102), .O(gate1913inter1));
  and2  gate4230(.a(N6653), .b(N6111), .O(gate1913inter2));
  inv1  gate4231(.a(s_102), .O(gate1913inter3));
  inv1  gate4232(.a(s_103), .O(gate1913inter4));
  nand2 gate4233(.a(gate1913inter4), .b(gate1913inter3), .O(gate1913inter5));
  nor2  gate4234(.a(gate1913inter5), .b(gate1913inter2), .O(gate1913inter6));
  inv1  gate4235(.a(N6111), .O(gate1913inter7));
  inv1  gate4236(.a(N6653), .O(gate1913inter8));
  nand2 gate4237(.a(gate1913inter8), .b(gate1913inter7), .O(gate1913inter9));
  nand2 gate4238(.a(s_103), .b(gate1913inter3), .O(gate1913inter10));
  nor2  gate4239(.a(gate1913inter10), .b(gate1913inter9), .O(gate1913inter11));
  nor2  gate4240(.a(gate1913inter11), .b(gate1913inter6), .O(gate1913inter12));
  nand2 gate4241(.a(gate1913inter12), .b(gate1913inter1), .O(N7258));
nand2 gate1914( .a(N6113), .b(N6654), .O(N7272) );
nand2 gate1915( .a(N6115), .b(N6655), .O(N7288) );
nand2 gate1916( .a(N6117), .b(N6656), .O(N7301) );
nand2 gate1917( .a(N6119), .b(N6657), .O(N7307) );
nand2 gate1918( .a(N6658), .b(N6122), .O(N7314) );
nand2 gate1919( .a(N6659), .b(N6660), .O(N7318) );

  xor2  gate4718(.a(N6661), .b(N6125), .O(gate1920inter0));
  nand2 gate4719(.a(gate1920inter0), .b(s_172), .O(gate1920inter1));
  and2  gate4720(.a(N6661), .b(N6125), .O(gate1920inter2));
  inv1  gate4721(.a(s_172), .O(gate1920inter3));
  inv1  gate4722(.a(s_173), .O(gate1920inter4));
  nand2 gate4723(.a(gate1920inter4), .b(gate1920inter3), .O(gate1920inter5));
  nor2  gate4724(.a(gate1920inter5), .b(gate1920inter2), .O(gate1920inter6));
  inv1  gate4725(.a(N6125), .O(gate1920inter7));
  inv1  gate4726(.a(N6661), .O(gate1920inter8));
  nand2 gate4727(.a(gate1920inter8), .b(gate1920inter7), .O(gate1920inter9));
  nand2 gate4728(.a(s_173), .b(gate1920inter3), .O(gate1920inter10));
  nor2  gate4729(.a(gate1920inter10), .b(gate1920inter9), .O(gate1920inter11));
  nor2  gate4730(.a(gate1920inter11), .b(gate1920inter6), .O(gate1920inter12));
  nand2 gate4731(.a(gate1920inter12), .b(gate1920inter1), .O(N7322));
inv1 gate1921( .a(N6127), .O(N7325) );
inv1 gate1922( .a(N6131), .O(N7328) );
nand2 gate1923( .a(N6668), .b(N6136), .O(N7331) );
inv1 gate1924( .a(N6137), .O(N7334) );
inv1 gate1925( .a(N6141), .O(N7337) );
buf1 gate1926( .a(N6145), .O(N7340) );
buf1 gate1927( .a(N6145), .O(N7343) );
nand2 gate1928( .a(N6677), .b(N6678), .O(N7346) );
nand2 gate1929( .a(N6679), .b(N6680), .O(N7351) );

  xor2  gate4508(.a(N6682), .b(N6681), .O(gate1930inter0));
  nand2 gate4509(.a(gate1930inter0), .b(s_142), .O(gate1930inter1));
  and2  gate4510(.a(N6682), .b(N6681), .O(gate1930inter2));
  inv1  gate4511(.a(s_142), .O(gate1930inter3));
  inv1  gate4512(.a(s_143), .O(gate1930inter4));
  nand2 gate4513(.a(gate1930inter4), .b(gate1930inter3), .O(gate1930inter5));
  nor2  gate4514(.a(gate1930inter5), .b(gate1930inter2), .O(gate1930inter6));
  inv1  gate4515(.a(N6681), .O(gate1930inter7));
  inv1  gate4516(.a(N6682), .O(gate1930inter8));
  nand2 gate4517(.a(gate1930inter8), .b(gate1930inter7), .O(gate1930inter9));
  nand2 gate4518(.a(s_143), .b(gate1930inter3), .O(gate1930inter10));
  nor2  gate4519(.a(gate1930inter10), .b(gate1930inter9), .O(gate1930inter11));
  nor2  gate4520(.a(gate1930inter11), .b(gate1930inter6), .O(gate1930inter12));
  nand2 gate4521(.a(gate1930inter12), .b(gate1930inter1), .O(N7355));
nand2 gate1931( .a(N6683), .b(N6684), .O(N7358) );
nand2 gate1932( .a(N6685), .b(N6157), .O(N7364) );
nand2 gate1933( .a(N6686), .b(N6159), .O(N7369) );
nand2 gate1934( .a(N6687), .b(N6161), .O(N7373) );
nand2 gate1935( .a(N6688), .b(N6689), .O(N7376) );
nand2 gate1936( .a(N6164), .b(N6690), .O(N7377) );
inv1 gate1937( .a(N6166), .O(N7378) );
inv1 gate1938( .a(N6170), .O(N7381) );
inv1 gate1939( .a(N6177), .O(N7384) );
nand2 gate1940( .a(N6702), .b(N6703), .O(N7387) );
nand2 gate1941( .a(N6704), .b(N6705), .O(N7391) );
nand2 gate1942( .a(N6706), .b(N6186), .O(N7394) );
nand2 gate1943( .a(N6707), .b(N6708), .O(N7398) );
nand2 gate1944( .a(N6709), .b(N6710), .O(N7402) );
buf1 gate1945( .a(N6174), .O(N7405) );
buf1 gate1946( .a(N6174), .O(N7408) );
buf1 gate1947( .a(N5936), .O(N7411) );
buf1 gate1948( .a(N5898), .O(N7414) );
buf1 gate1949( .a(N5905), .O(N7417) );
buf1 gate1950( .a(N5915), .O(N7420) );
buf1 gate1951( .a(N5926), .O(N7423) );
buf1 gate1952( .a(N5728), .O(N7426) );
buf1 gate1953( .a(N5690), .O(N7429) );
buf1 gate1954( .a(N5697), .O(N7432) );
buf1 gate1955( .a(N5707), .O(N7435) );
buf1 gate1956( .a(N5718), .O(N7438) );
nand2 gate1957( .a(N6192), .b(N6711), .O(N7441) );
nand2 gate1958( .a(N6194), .b(N6712), .O(N7444) );
buf1 gate1959( .a(N5683), .O(N7447) );
buf1 gate1960( .a(N5670), .O(N7450) );
buf1 gate1961( .a(N5632), .O(N7453) );
buf1 gate1962( .a(N5654), .O(N7456) );
buf1 gate1963( .a(N5640), .O(N7459) );
buf1 gate1964( .a(N5640), .O(N7462) );
buf1 gate1965( .a(N5683), .O(N7465) );
buf1 gate1966( .a(N5670), .O(N7468) );
buf1 gate1967( .a(N5632), .O(N7471) );
buf1 gate1968( .a(N5654), .O(N7474) );
inv1 gate1969( .a(N6196), .O(N7477) );
inv1 gate1970( .a(N6199), .O(N7478) );
buf1 gate1971( .a(N5850), .O(N7479) );
buf1 gate1972( .a(N5789), .O(N7482) );
buf1 gate1973( .a(N5771), .O(N7485) );
buf1 gate1974( .a(N5778), .O(N7488) );
buf1 gate1975( .a(N5850), .O(N7491) );
buf1 gate1976( .a(N5789), .O(N7494) );
buf1 gate1977( .a(N5771), .O(N7497) );
buf1 gate1978( .a(N5778), .O(N7500) );
buf1 gate1979( .a(N5856), .O(N7503) );
buf1 gate1980( .a(N5837), .O(N7506) );
buf1 gate1981( .a(N5799), .O(N7509) );
buf1 gate1982( .a(N5821), .O(N7512) );
buf1 gate1983( .a(N5807), .O(N7515) );
buf1 gate1984( .a(N5807), .O(N7518) );
buf1 gate1985( .a(N5856), .O(N7521) );
buf1 gate1986( .a(N5837), .O(N7524) );
buf1 gate1987( .a(N5799), .O(N7527) );
buf1 gate1988( .a(N5821), .O(N7530) );
buf1 gate1989( .a(N5863), .O(N7533) );
buf1 gate1990( .a(N5863), .O(N7536) );
buf1 gate1991( .a(N5870), .O(N7539) );
buf1 gate1992( .a(N5870), .O(N7542) );
buf1 gate1993( .a(N5881), .O(N7545) );
buf1 gate1994( .a(N5881), .O(N7548) );
inv1 gate1995( .a(N6214), .O(N7551) );
inv1 gate1996( .a(N6217), .O(N7552) );
buf1 gate1997( .a(N5981), .O(N7553) );
inv1 gate1998( .a(N6249), .O(N7556) );
inv1 gate1999( .a(N6252), .O(N7557) );
inv1 gate2000( .a(N6243), .O(N7558) );
inv1 gate2001( .a(N6246), .O(N7559) );
nand2 gate2002( .a(N6731), .b(N6732), .O(N7560) );
nand2 gate2003( .a(N6729), .b(N6730), .O(N7563) );
nand2 gate2004( .a(N6735), .b(N6736), .O(N7566) );
nand2 gate2005( .a(N6733), .b(N6734), .O(N7569) );
inv1 gate2006( .a(N6232), .O(N7572) );
inv1 gate2007( .a(N6236), .O(N7573) );
nand2 gate2008( .a(N6743), .b(N6744), .O(N7574) );
nand2 gate2009( .a(N6741), .b(N6742), .O(N7577) );
inv1 gate2010( .a(N6263), .O(N7580) );
inv1 gate2011( .a(N6266), .O(N7581) );
nand2 gate2012( .a(N6753), .b(N6754), .O(N7582) );
nand2 gate2013( .a(N6751), .b(N6752), .O(N7585) );
nand2 gate2014( .a(N6757), .b(N6758), .O(N7588) );
nand2 gate2015( .a(N6755), .b(N6756), .O(N7591) );
or5 gate2016( .a(N3096), .b(N6766), .c(N6767), .d(N6768), .e(N6769), .O(N7609) );
or2 gate2017( .a(N3107), .b(N6782), .O(N7613) );
or5 gate2018( .a(N3136), .b(N6787), .c(N6788), .d(N6789), .e(N6790), .O(N7620) );
or4 gate2019( .a(N3168), .b(N6836), .c(N6837), .d(N6838), .O(N7649) );
or2 gate2020( .a(N3173), .b(N6844), .O(N7650) );
or5 gate2021( .a(N3184), .b(N6848), .c(N6849), .d(N6850), .e(N6851), .O(N7655) );
or2 gate2022( .a(N3195), .b(N6864), .O(N7659) );
or4 gate2023( .a(N3210), .b(N6870), .c(N6871), .d(N6872), .O(N7668) );
or5 gate2024( .a(N3228), .b(N6884), .c(N6885), .d(N6886), .e(N6887), .O(N7671) );
nand2 gate2025( .a(N3661), .b(N6968), .O(N7744) );
nand2 gate2026( .a(N3664), .b(N7056), .O(N7822) );
or4 gate2027( .a(N3361), .b(N7060), .c(N7061), .d(N7062), .O(N7825) );
or5 gate2028( .a(N3365), .b(N7064), .c(N7065), .d(N7066), .e(N7067), .O(N7826) );
or5 gate2029( .a(N3370), .b(N7103), .c(N7104), .d(N7105), .e(N7106), .O(N7852) );
or4 gate2030( .a(N3101), .b(N6777), .c(N6778), .d(N6779), .O(N8114) );
or5 gate2031( .a(N3097), .b(N6770), .c(N6771), .d(N6772), .e(N6773), .O(N8117) );
nor3 gate2032( .a(N3101), .b(N6780), .c(N6781), .O(N8131) );
nor4 gate2033( .a(N3097), .b(N6774), .c(N6775), .d(N6776), .O(N8134) );
nand2 gate2034( .a(N6199), .b(N7477), .O(N8144) );
nand2 gate2035( .a(N6196), .b(N7478), .O(N8145) );
or4 gate2036( .a(N3169), .b(N6839), .c(N6840), .d(N6841), .O(N8146) );
nor3 gate2037( .a(N3169), .b(N6842), .c(N6843), .O(N8156) );
or4 gate2038( .a(N3189), .b(N6859), .c(N6860), .d(N6861), .O(N8166) );
or5 gate2039( .a(N3185), .b(N6852), .c(N6853), .d(N6854), .e(N6855), .O(N8169) );
nor3 gate2040( .a(N3189), .b(N6862), .c(N6863), .O(N8183) );
nor4 gate2041( .a(N3185), .b(N6856), .c(N6857), .d(N6858), .O(N8186) );
or4 gate2042( .a(N3211), .b(N6873), .c(N6874), .d(N6875), .O(N8196) );
nor3 gate2043( .a(N3211), .b(N6876), .c(N6877), .O(N8200) );
or3 gate2044( .a(N3215), .b(N6878), .c(N6879), .O(N8204) );
nor2 gate2045( .a(N3215), .b(N6880), .O(N8208) );
nand2 gate2046( .a(N6252), .b(N7556), .O(N8216) );

  xor2  gate4270(.a(N7557), .b(N6249), .O(gate2047inter0));
  nand2 gate4271(.a(gate2047inter0), .b(s_108), .O(gate2047inter1));
  and2  gate4272(.a(N7557), .b(N6249), .O(gate2047inter2));
  inv1  gate4273(.a(s_108), .O(gate2047inter3));
  inv1  gate4274(.a(s_109), .O(gate2047inter4));
  nand2 gate4275(.a(gate2047inter4), .b(gate2047inter3), .O(gate2047inter5));
  nor2  gate4276(.a(gate2047inter5), .b(gate2047inter2), .O(gate2047inter6));
  inv1  gate4277(.a(N6249), .O(gate2047inter7));
  inv1  gate4278(.a(N7557), .O(gate2047inter8));
  nand2 gate4279(.a(gate2047inter8), .b(gate2047inter7), .O(gate2047inter9));
  nand2 gate4280(.a(s_109), .b(gate2047inter3), .O(gate2047inter10));
  nor2  gate4281(.a(gate2047inter10), .b(gate2047inter9), .O(gate2047inter11));
  nor2  gate4282(.a(gate2047inter11), .b(gate2047inter6), .O(gate2047inter12));
  nand2 gate4283(.a(gate2047inter12), .b(gate2047inter1), .O(N8217));
nand2 gate2048( .a(N6246), .b(N7558), .O(N8218) );
nand2 gate2049( .a(N6243), .b(N7559), .O(N8219) );

  xor2  gate4760(.a(N7580), .b(N6266), .O(gate2050inter0));
  nand2 gate4761(.a(gate2050inter0), .b(s_178), .O(gate2050inter1));
  and2  gate4762(.a(N7580), .b(N6266), .O(gate2050inter2));
  inv1  gate4763(.a(s_178), .O(gate2050inter3));
  inv1  gate4764(.a(s_179), .O(gate2050inter4));
  nand2 gate4765(.a(gate2050inter4), .b(gate2050inter3), .O(gate2050inter5));
  nor2  gate4766(.a(gate2050inter5), .b(gate2050inter2), .O(gate2050inter6));
  inv1  gate4767(.a(N6266), .O(gate2050inter7));
  inv1  gate4768(.a(N7580), .O(gate2050inter8));
  nand2 gate4769(.a(gate2050inter8), .b(gate2050inter7), .O(gate2050inter9));
  nand2 gate4770(.a(s_179), .b(gate2050inter3), .O(gate2050inter10));
  nor2  gate4771(.a(gate2050inter10), .b(gate2050inter9), .O(gate2050inter11));
  nor2  gate4772(.a(gate2050inter11), .b(gate2050inter6), .O(gate2050inter12));
  nand2 gate4773(.a(gate2050inter12), .b(gate2050inter1), .O(N8232));
nand2 gate2051( .a(N6263), .b(N7581), .O(N8233) );
inv1 gate2052( .a(N7411), .O(N8242) );
inv1 gate2053( .a(N7414), .O(N8243) );
inv1 gate2054( .a(N7417), .O(N8244) );
inv1 gate2055( .a(N7420), .O(N8245) );
inv1 gate2056( .a(N7423), .O(N8246) );
inv1 gate2057( .a(N7426), .O(N8247) );
inv1 gate2058( .a(N7429), .O(N8248) );
inv1 gate2059( .a(N7432), .O(N8249) );
inv1 gate2060( .a(N7435), .O(N8250) );
inv1 gate2061( .a(N7438), .O(N8251) );
inv1 gate2062( .a(N7136), .O(N8252) );
inv1 gate2063( .a(N6923), .O(N8253) );
inv1 gate2064( .a(N6762), .O(N8254) );
inv1 gate2065( .a(N7459), .O(N8260) );
inv1 gate2066( .a(N7462), .O(N8261) );
and2 gate2067( .a(N3122), .b(N6762), .O(N8262) );
and2 gate2068( .a(N3155), .b(N6784), .O(N8269) );
inv1 gate2069( .a(N6815), .O(N8274) );
inv1 gate2070( .a(N6818), .O(N8275) );
inv1 gate2071( .a(N6821), .O(N8276) );
inv1 gate2072( .a(N6824), .O(N8277) );
inv1 gate2073( .a(N6827), .O(N8278) );
inv1 gate2074( .a(N6830), .O(N8279) );
and3 gate2075( .a(N5740), .b(N5736), .c(N6815), .O(N8280) );
and3 gate2076( .a(N6800), .b(N6797), .c(N6818), .O(N8281) );
and3 gate2077( .a(N5751), .b(N5747), .c(N6821), .O(N8282) );
and3 gate2078( .a(N6806), .b(N6803), .c(N6824), .O(N8283) );
and3 gate2079( .a(N5762), .b(N5758), .c(N6827), .O(N8284) );
and3 gate2080( .a(N6812), .b(N6809), .c(N6830), .O(N8285) );
inv1 gate2081( .a(N6845), .O(N8288) );
inv1 gate2082( .a(N7488), .O(N8294) );
inv1 gate2083( .a(N7500), .O(N8295) );
inv1 gate2084( .a(N7515), .O(N8296) );
inv1 gate2085( .a(N7518), .O(N8297) );
and2 gate2086( .a(N6833), .b(N6845), .O(N8298) );
and2 gate2087( .a(N6867), .b(N6881), .O(N8307) );
inv1 gate2088( .a(N7533), .O(N8315) );
inv1 gate2089( .a(N7536), .O(N8317) );
inv1 gate2090( .a(N7539), .O(N8319) );
inv1 gate2091( .a(N7542), .O(N8321) );
nand2 gate2092( .a(N7545), .b(N4543), .O(N8322) );
inv1 gate2093( .a(N7545), .O(N8323) );
nand2 gate2094( .a(N7548), .b(N5943), .O(N8324) );
inv1 gate2095( .a(N7548), .O(N8325) );
nand2 gate2096( .a(N6967), .b(N7744), .O(N8326) );
and4 gate2097( .a(N6901), .b(N6923), .c(N6912), .d(N6894), .O(N8333) );
and2 gate2098( .a(N6894), .b(N4545), .O(N8337) );
and3 gate2099( .a(N6901), .b(N6894), .c(N4549), .O(N8338) );
and4 gate2100( .a(N6912), .b(N6894), .c(N4555), .d(N6901), .O(N8339) );
and2 gate2101( .a(N6901), .b(N4549), .O(N8340) );
and3 gate2102( .a(N6912), .b(N4555), .c(N6901), .O(N8341) );
and3 gate2103( .a(N6923), .b(N6912), .c(N6901), .O(N8342) );
and2 gate2104( .a(N6901), .b(N4549), .O(N8343) );
and3 gate2105( .a(N4555), .b(N6912), .c(N6901), .O(N8344) );
and2 gate2106( .a(N6912), .b(N4555), .O(N8345) );
and2 gate2107( .a(N6923), .b(N6912), .O(N8346) );
and2 gate2108( .a(N6912), .b(N4555), .O(N8347) );
and2 gate2109( .a(N6929), .b(N4563), .O(N8348) );
and3 gate2110( .a(N6936), .b(N6929), .c(N4566), .O(N8349) );
and4 gate2111( .a(N6946), .b(N6929), .c(N4570), .d(N6936), .O(N8350) );
and5 gate2112( .a(N6957), .b(N6946), .c(N6929), .d(N5960), .e(N6936), .O(N8351) );
and2 gate2113( .a(N6936), .b(N4566), .O(N8352) );
and3 gate2114( .a(N6946), .b(N4570), .c(N6936), .O(N8353) );
and4 gate2115( .a(N6957), .b(N6946), .c(N5960), .d(N6936), .O(N8354) );
and2 gate2116( .a(N4570), .b(N6946), .O(N8355) );
and3 gate2117( .a(N6957), .b(N6946), .c(N5960), .O(N8356) );
and2 gate2118( .a(N6957), .b(N5960), .O(N8357) );
nand2 gate2119( .a(N7055), .b(N7822), .O(N8358) );
and4 gate2120( .a(N7049), .b(N6988), .c(N6977), .d(N6970), .O(N8365) );
and2 gate2121( .a(N6970), .b(N4577), .O(N8369) );
and3 gate2122( .a(N6977), .b(N6970), .c(N4581), .O(N8370) );
and4 gate2123( .a(N6988), .b(N6970), .c(N4586), .d(N6977), .O(N8371) );
and2 gate2124( .a(N6977), .b(N4581), .O(N8372) );
and3 gate2125( .a(N6988), .b(N4586), .c(N6977), .O(N8373) );
and3 gate2126( .a(N7049), .b(N6988), .c(N6977), .O(N8374) );
and2 gate2127( .a(N6977), .b(N4581), .O(N8375) );
and3 gate2128( .a(N6988), .b(N4586), .c(N6977), .O(N8376) );
and2 gate2129( .a(N6988), .b(N4586), .O(N8377) );
and2 gate2130( .a(N6998), .b(N4593), .O(N8378) );
and3 gate2131( .a(N7006), .b(N6998), .c(N4597), .O(N8379) );
and4 gate2132( .a(N7020), .b(N6998), .c(N4603), .d(N7006), .O(N8380) );
and5 gate2133( .a(N7036), .b(N7020), .c(N6998), .d(N5981), .e(N7006), .O(N8381) );
and2 gate2134( .a(N7006), .b(N4597), .O(N8382) );
and3 gate2135( .a(N7020), .b(N4603), .c(N7006), .O(N8383) );
and4 gate2136( .a(N7036), .b(N7020), .c(N5981), .d(N7006), .O(N8384) );
and2 gate2137( .a(N7006), .b(N4597), .O(N8385) );
and3 gate2138( .a(N7020), .b(N4603), .c(N7006), .O(N8386) );
and4 gate2139( .a(N7036), .b(N7020), .c(N5981), .d(N7006), .O(N8387) );
and2 gate2140( .a(N7020), .b(N4603), .O(N8388) );
and3 gate2141( .a(N7036), .b(N7020), .c(N5981), .O(N8389) );
and2 gate2142( .a(N7020), .b(N4603), .O(N8390) );
and3 gate2143( .a(N7036), .b(N7020), .c(N5981), .O(N8391) );
and2 gate2144( .a(N7036), .b(N5981), .O(N8392) );
and2 gate2145( .a(N7049), .b(N6988), .O(N8393) );
and2 gate2146( .a(N7057), .b(N7063), .O(N8394) );
and2 gate2147( .a(N7057), .b(N7826), .O(N8404) );
and4 gate2148( .a(N7098), .b(N7077), .c(N7073), .d(N7068), .O(N8405) );
and2 gate2149( .a(N7068), .b(N4632), .O(N8409) );
and3 gate2150( .a(N7073), .b(N7068), .c(N4634), .O(N8410) );
and4 gate2151( .a(N7077), .b(N7068), .c(N4635), .d(N7073), .O(N8411) );
and5 gate2152( .a(N7099), .b(N7095), .c(N7091), .d(N7086), .e(N7080), .O(N8412) );
and2 gate2153( .a(N7080), .b(N4638), .O(N8415) );
and3 gate2154( .a(N7086), .b(N7080), .c(N4639), .O(N8416) );
and4 gate2155( .a(N7091), .b(N7080), .c(N4640), .d(N7086), .O(N8417) );
and5 gate2156( .a(N7095), .b(N7091), .c(N7080), .d(N4641), .e(N7086), .O(N8418) );
and2 gate2157( .a(N3375), .b(N7100), .O(N8421) );
and4 gate2158( .a(N7114), .b(N7136), .c(N7125), .d(N7107), .O(N8430) );
and2 gate2159( .a(N7107), .b(N4657), .O(N8433) );
and3 gate2160( .a(N7114), .b(N7107), .c(N4661), .O(N8434) );
and4 gate2161( .a(N7125), .b(N7107), .c(N4667), .d(N7114), .O(N8435) );
and2 gate2162( .a(N7114), .b(N4661), .O(N8436) );
and3 gate2163( .a(N7125), .b(N4667), .c(N7114), .O(N8437) );
and3 gate2164( .a(N7136), .b(N7125), .c(N7114), .O(N8438) );
and2 gate2165( .a(N7114), .b(N4661), .O(N8439) );
and3 gate2166( .a(N4667), .b(N7125), .c(N7114), .O(N8440) );
and2 gate2167( .a(N7125), .b(N4667), .O(N8441) );
and2 gate2168( .a(N7136), .b(N7125), .O(N8442) );
and2 gate2169( .a(N7125), .b(N4667), .O(N8443) );
and5 gate2170( .a(N7149), .b(N7180), .c(N7159), .d(N7142), .e(N7170), .O(N8444) );
and2 gate2171( .a(N7142), .b(N4675), .O(N8447) );
and3 gate2172( .a(N7149), .b(N7142), .c(N4678), .O(N8448) );
and4 gate2173( .a(N7159), .b(N7142), .c(N4682), .d(N7149), .O(N8449) );
and5 gate2174( .a(N7170), .b(N7159), .c(N7142), .d(N4687), .e(N7149), .O(N8450) );
and2 gate2175( .a(N7149), .b(N4678), .O(N8451) );
and3 gate2176( .a(N7159), .b(N4682), .c(N7149), .O(N8452) );
and4 gate2177( .a(N7170), .b(N7159), .c(N4687), .d(N7149), .O(N8453) );
and2 gate2178( .a(N4682), .b(N7159), .O(N8454) );
and3 gate2179( .a(N7170), .b(N7159), .c(N4687), .O(N8455) );
and2 gate2180( .a(N7170), .b(N4687), .O(N8456) );
inv1 gate2181( .a(N7194), .O(N8457) );
inv1 gate2182( .a(N7198), .O(N8460) );
inv1 gate2183( .a(N7205), .O(N8463) );
inv1 gate2184( .a(N7209), .O(N8466) );
inv1 gate2185( .a(N7216), .O(N8469) );
inv1 gate2186( .a(N7219), .O(N8470) );
buf1 gate2187( .a(N7202), .O(N8471) );
buf1 gate2188( .a(N7202), .O(N8474) );
buf1 gate2189( .a(N7213), .O(N8477) );
buf1 gate2190( .a(N7213), .O(N8480) );
and3 gate2191( .a(N6083), .b(N6079), .c(N7216), .O(N8483) );
and3 gate2192( .a(N7191), .b(N7188), .c(N7219), .O(N8484) );
and4 gate2193( .a(N7301), .b(N7240), .c(N7229), .d(N7222), .O(N8485) );
and2 gate2194( .a(N7222), .b(N4702), .O(N8488) );
and3 gate2195( .a(N7229), .b(N7222), .c(N4706), .O(N8489) );
and4 gate2196( .a(N7240), .b(N7222), .c(N4711), .d(N7229), .O(N8490) );
and2 gate2197( .a(N7229), .b(N4706), .O(N8491) );
and3 gate2198( .a(N7240), .b(N4711), .c(N7229), .O(N8492) );
and3 gate2199( .a(N7301), .b(N7240), .c(N7229), .O(N8493) );
and2 gate2200( .a(N7229), .b(N4706), .O(N8494) );
and3 gate2201( .a(N7240), .b(N4711), .c(N7229), .O(N8495) );
and2 gate2202( .a(N7240), .b(N4711), .O(N8496) );
and5 gate2203( .a(N7307), .b(N7288), .c(N7272), .d(N7258), .e(N7250), .O(N8497) );
and2 gate2204( .a(N7250), .b(N4718), .O(N8500) );
and3 gate2205( .a(N7258), .b(N7250), .c(N4722), .O(N8501) );
and4 gate2206( .a(N7272), .b(N7250), .c(N4728), .d(N7258), .O(N8502) );
and5 gate2207( .a(N7288), .b(N7272), .c(N7250), .d(N4735), .e(N7258), .O(N8503) );
and2 gate2208( .a(N7258), .b(N4722), .O(N8504) );
and3 gate2209( .a(N7272), .b(N4728), .c(N7258), .O(N8505) );
and4 gate2210( .a(N7288), .b(N7272), .c(N4735), .d(N7258), .O(N8506) );
and4 gate2211( .a(N7307), .b(N7272), .c(N7258), .d(N7288), .O(N8507) );
and2 gate2212( .a(N7258), .b(N4722), .O(N8508) );
and3 gate2213( .a(N7272), .b(N4728), .c(N7258), .O(N8509) );
and4 gate2214( .a(N7288), .b(N7272), .c(N4735), .d(N7258), .O(N8510) );
and2 gate2215( .a(N7272), .b(N4728), .O(N8511) );
and3 gate2216( .a(N7288), .b(N7272), .c(N4735), .O(N8512) );
and3 gate2217( .a(N7307), .b(N7272), .c(N7288), .O(N8513) );
and2 gate2218( .a(N7272), .b(N4728), .O(N8514) );
and3 gate2219( .a(N7288), .b(N7272), .c(N4735), .O(N8515) );
and2 gate2220( .a(N7288), .b(N4735), .O(N8516) );
and2 gate2221( .a(N7301), .b(N7240), .O(N8517) );
and2 gate2222( .a(N7307), .b(N7288), .O(N8518) );
inv1 gate2223( .a(N7314), .O(N8519) );
inv1 gate2224( .a(N7318), .O(N8522) );
buf1 gate2225( .a(N7322), .O(N8525) );
buf1 gate2226( .a(N7322), .O(N8528) );
buf1 gate2227( .a(N7331), .O(N8531) );
buf1 gate2228( .a(N7331), .O(N8534) );
inv1 gate2229( .a(N7340), .O(N8537) );
inv1 gate2230( .a(N7343), .O(N8538) );
and3 gate2231( .a(N6141), .b(N6137), .c(N7340), .O(N8539) );
and3 gate2232( .a(N7337), .b(N7334), .c(N7343), .O(N8540) );
and4 gate2233( .a(N7376), .b(N7355), .c(N7351), .d(N7346), .O(N8541) );
and2 gate2234( .a(N7346), .b(N4757), .O(N8545) );
and3 gate2235( .a(N7351), .b(N7346), .c(N4758), .O(N8546) );
and4 gate2236( .a(N7355), .b(N7346), .c(N4759), .d(N7351), .O(N8547) );
and5 gate2237( .a(N7377), .b(N7373), .c(N7369), .d(N7364), .e(N7358), .O(N8548) );
and2 gate2238( .a(N7358), .b(N4762), .O(N8551) );
and3 gate2239( .a(N7364), .b(N7358), .c(N4764), .O(N8552) );
and4 gate2240( .a(N7369), .b(N7358), .c(N4766), .d(N7364), .O(N8553) );
and5 gate2241( .a(N7373), .b(N7369), .c(N7358), .d(N4767), .e(N7364), .O(N8554) );
inv1 gate2242( .a(N7387), .O(N8555) );
inv1 gate2243( .a(N7394), .O(N8558) );
inv1 gate2244( .a(N7398), .O(N8561) );
inv1 gate2245( .a(N7405), .O(N8564) );
inv1 gate2246( .a(N7408), .O(N8565) );
buf1 gate2247( .a(N7391), .O(N8566) );
buf1 gate2248( .a(N7391), .O(N8569) );
buf1 gate2249( .a(N7402), .O(N8572) );
buf1 gate2250( .a(N7402), .O(N8575) );
and3 gate2251( .a(N6170), .b(N6166), .c(N7405), .O(N8578) );
and3 gate2252( .a(N7381), .b(N7378), .c(N7408), .O(N8579) );
buf1 gate2253( .a(N7180), .O(N8580) );
buf1 gate2254( .a(N7142), .O(N8583) );
buf1 gate2255( .a(N7149), .O(N8586) );
buf1 gate2256( .a(N7159), .O(N8589) );
buf1 gate2257( .a(N7170), .O(N8592) );
buf1 gate2258( .a(N6929), .O(N8595) );
buf1 gate2259( .a(N6936), .O(N8598) );
buf1 gate2260( .a(N6946), .O(N8601) );
buf1 gate2261( .a(N6957), .O(N8604) );
inv1 gate2262( .a(N7441), .O(N8607) );

  xor2  gate3542(.a(N5469), .b(N7441), .O(gate2263inter0));
  nand2 gate3543(.a(gate2263inter0), .b(s_4), .O(gate2263inter1));
  and2  gate3544(.a(N5469), .b(N7441), .O(gate2263inter2));
  inv1  gate3545(.a(s_4), .O(gate2263inter3));
  inv1  gate3546(.a(s_5), .O(gate2263inter4));
  nand2 gate3547(.a(gate2263inter4), .b(gate2263inter3), .O(gate2263inter5));
  nor2  gate3548(.a(gate2263inter5), .b(gate2263inter2), .O(gate2263inter6));
  inv1  gate3549(.a(N7441), .O(gate2263inter7));
  inv1  gate3550(.a(N5469), .O(gate2263inter8));
  nand2 gate3551(.a(gate2263inter8), .b(gate2263inter7), .O(gate2263inter9));
  nand2 gate3552(.a(s_5), .b(gate2263inter3), .O(gate2263inter10));
  nor2  gate3553(.a(gate2263inter10), .b(gate2263inter9), .O(gate2263inter11));
  nor2  gate3554(.a(gate2263inter11), .b(gate2263inter6), .O(gate2263inter12));
  nand2 gate3555(.a(gate2263inter12), .b(gate2263inter1), .O(N8608));
inv1 gate2264( .a(N7444), .O(N8609) );
nand2 gate2265( .a(N7444), .b(N4793), .O(N8610) );
inv1 gate2266( .a(N7447), .O(N8615) );
inv1 gate2267( .a(N7450), .O(N8616) );
inv1 gate2268( .a(N7453), .O(N8617) );
inv1 gate2269( .a(N7456), .O(N8618) );
inv1 gate2270( .a(N7474), .O(N8619) );
inv1 gate2271( .a(N7465), .O(N8624) );
inv1 gate2272( .a(N7468), .O(N8625) );
inv1 gate2273( .a(N7471), .O(N8626) );
nand2 gate2274( .a(N8144), .b(N8145), .O(N8627) );
inv1 gate2275( .a(N7479), .O(N8632) );
inv1 gate2276( .a(N7482), .O(N8633) );
inv1 gate2277( .a(N7485), .O(N8634) );
inv1 gate2278( .a(N7491), .O(N8637) );
inv1 gate2279( .a(N7494), .O(N8638) );
inv1 gate2280( .a(N7497), .O(N8639) );
inv1 gate2281( .a(N7503), .O(N8644) );
inv1 gate2282( .a(N7506), .O(N8645) );
inv1 gate2283( .a(N7509), .O(N8646) );
inv1 gate2284( .a(N7512), .O(N8647) );
inv1 gate2285( .a(N7530), .O(N8648) );
inv1 gate2286( .a(N7521), .O(N8653) );
inv1 gate2287( .a(N7524), .O(N8654) );
inv1 gate2288( .a(N7527), .O(N8655) );
buf1 gate2289( .a(N6894), .O(N8660) );
buf1 gate2290( .a(N6894), .O(N8663) );
buf1 gate2291( .a(N6901), .O(N8666) );
buf1 gate2292( .a(N6901), .O(N8669) );
buf1 gate2293( .a(N6912), .O(N8672) );
buf1 gate2294( .a(N6912), .O(N8675) );
buf1 gate2295( .a(N7049), .O(N8678) );
buf1 gate2296( .a(N6988), .O(N8681) );
buf1 gate2297( .a(N6970), .O(N8684) );
buf1 gate2298( .a(N6977), .O(N8687) );
buf1 gate2299( .a(N7049), .O(N8690) );
buf1 gate2300( .a(N6988), .O(N8693) );
buf1 gate2301( .a(N6970), .O(N8696) );
buf1 gate2302( .a(N6977), .O(N8699) );
buf1 gate2303( .a(N7036), .O(N8702) );
buf1 gate2304( .a(N6998), .O(N8705) );
buf1 gate2305( .a(N7020), .O(N8708) );
buf1 gate2306( .a(N7006), .O(N8711) );
buf1 gate2307( .a(N7006), .O(N8714) );
inv1 gate2308( .a(N7553), .O(N8717) );
buf1 gate2309( .a(N7036), .O(N8718) );
buf1 gate2310( .a(N6998), .O(N8721) );
buf1 gate2311( .a(N7020), .O(N8724) );

  xor2  gate4634(.a(N8217), .b(N8216), .O(gate2312inter0));
  nand2 gate4635(.a(gate2312inter0), .b(s_160), .O(gate2312inter1));
  and2  gate4636(.a(N8217), .b(N8216), .O(gate2312inter2));
  inv1  gate4637(.a(s_160), .O(gate2312inter3));
  inv1  gate4638(.a(s_161), .O(gate2312inter4));
  nand2 gate4639(.a(gate2312inter4), .b(gate2312inter3), .O(gate2312inter5));
  nor2  gate4640(.a(gate2312inter5), .b(gate2312inter2), .O(gate2312inter6));
  inv1  gate4641(.a(N8216), .O(gate2312inter7));
  inv1  gate4642(.a(N8217), .O(gate2312inter8));
  nand2 gate4643(.a(gate2312inter8), .b(gate2312inter7), .O(gate2312inter9));
  nand2 gate4644(.a(s_161), .b(gate2312inter3), .O(gate2312inter10));
  nor2  gate4645(.a(gate2312inter10), .b(gate2312inter9), .O(gate2312inter11));
  nor2  gate4646(.a(gate2312inter11), .b(gate2312inter6), .O(gate2312inter12));
  nand2 gate4647(.a(gate2312inter12), .b(gate2312inter1), .O(N8727));
nand2 gate2313( .a(N8218), .b(N8219), .O(N8730) );
inv1 gate2314( .a(N7574), .O(N8733) );
inv1 gate2315( .a(N7577), .O(N8734) );
buf1 gate2316( .a(N7107), .O(N8735) );
buf1 gate2317( .a(N7107), .O(N8738) );
buf1 gate2318( .a(N7114), .O(N8741) );
buf1 gate2319( .a(N7114), .O(N8744) );
buf1 gate2320( .a(N7125), .O(N8747) );
buf1 gate2321( .a(N7125), .O(N8750) );
inv1 gate2322( .a(N7560), .O(N8753) );
inv1 gate2323( .a(N7563), .O(N8754) );
inv1 gate2324( .a(N7566), .O(N8755) );
inv1 gate2325( .a(N7569), .O(N8756) );
buf1 gate2326( .a(N7301), .O(N8757) );
buf1 gate2327( .a(N7240), .O(N8760) );
buf1 gate2328( .a(N7222), .O(N8763) );
buf1 gate2329( .a(N7229), .O(N8766) );
buf1 gate2330( .a(N7301), .O(N8769) );
buf1 gate2331( .a(N7240), .O(N8772) );
buf1 gate2332( .a(N7222), .O(N8775) );
buf1 gate2333( .a(N7229), .O(N8778) );
buf1 gate2334( .a(N7307), .O(N8781) );
buf1 gate2335( .a(N7288), .O(N8784) );
buf1 gate2336( .a(N7250), .O(N8787) );
buf1 gate2337( .a(N7272), .O(N8790) );
buf1 gate2338( .a(N7258), .O(N8793) );
buf1 gate2339( .a(N7258), .O(N8796) );
buf1 gate2340( .a(N7307), .O(N8799) );
buf1 gate2341( .a(N7288), .O(N8802) );
buf1 gate2342( .a(N7250), .O(N8805) );
buf1 gate2343( .a(N7272), .O(N8808) );
nand2 gate2344( .a(N8232), .b(N8233), .O(N8811) );
inv1 gate2345( .a(N7588), .O(N8814) );
inv1 gate2346( .a(N7591), .O(N8815) );
inv1 gate2347( .a(N7582), .O(N8816) );
inv1 gate2348( .a(N7585), .O(N8817) );
and2 gate2349( .a(N7620), .b(N3155), .O(N8818) );
and2 gate2350( .a(N3122), .b(N7609), .O(N8840) );
inv1 gate2351( .a(N7609), .O(N8857) );
and3 gate2352( .a(N6797), .b(N5740), .c(N8274), .O(N8861) );
and3 gate2353( .a(N5736), .b(N6800), .c(N8275), .O(N8862) );
and3 gate2354( .a(N6803), .b(N5751), .c(N8276), .O(N8863) );
and3 gate2355( .a(N5747), .b(N6806), .c(N8277), .O(N8864) );
and3 gate2356( .a(N6809), .b(N5762), .c(N8278), .O(N8865) );
and3 gate2357( .a(N5758), .b(N6812), .c(N8279), .O(N8866) );
inv1 gate2358( .a(N7655), .O(N8871) );
and2 gate2359( .a(N6833), .b(N7655), .O(N8874) );
and2 gate2360( .a(N7671), .b(N6867), .O(N8878) );
inv1 gate2361( .a(N8196), .O(N8879) );
nand2 gate2362( .a(N8196), .b(N8315), .O(N8880) );
inv1 gate2363( .a(N8200), .O(N8881) );
nand2 gate2364( .a(N8200), .b(N8317), .O(N8882) );
inv1 gate2365( .a(N8204), .O(N8883) );
nand2 gate2366( .a(N8204), .b(N8319), .O(N8884) );
inv1 gate2367( .a(N8208), .O(N8885) );
nand2 gate2368( .a(N8208), .b(N8321), .O(N8886) );
nand2 gate2369( .a(N3658), .b(N8323), .O(N8887) );
nand2 gate2370( .a(N4817), .b(N8325), .O(N8888) );
or4 gate2371( .a(N4544), .b(N8337), .c(N8338), .d(N8339), .O(N8898) );
or5 gate2372( .a(N4562), .b(N8348), .c(N8349), .d(N8350), .e(N8351), .O(N8902) );
or4 gate2373( .a(N4576), .b(N8369), .c(N8370), .d(N8371), .O(N8920) );
or2 gate2374( .a(N4581), .b(N8377), .O(N8924) );
or5 gate2375( .a(N4592), .b(N8378), .c(N8379), .d(N8380), .e(N8381), .O(N8927) );
or2 gate2376( .a(N4603), .b(N8392), .O(N8931) );
or2 gate2377( .a(N7825), .b(N8404), .O(N8943) );
or4 gate2378( .a(N4630), .b(N8409), .c(N8410), .d(N8411), .O(N8950) );
or5 gate2379( .a(N4637), .b(N8415), .c(N8416), .d(N8417), .e(N8418), .O(N8956) );
inv1 gate2380( .a(N7852), .O(N8959) );
and2 gate2381( .a(N3375), .b(N7852), .O(N8960) );
or4 gate2382( .a(N4656), .b(N8433), .c(N8434), .d(N8435), .O(N8963) );
or5 gate2383( .a(N4674), .b(N8447), .c(N8448), .d(N8449), .e(N8450), .O(N8966) );
and3 gate2384( .a(N7188), .b(N6083), .c(N8469), .O(N8991) );
and3 gate2385( .a(N6079), .b(N7191), .c(N8470), .O(N8992) );
or4 gate2386( .a(N4701), .b(N8488), .c(N8489), .d(N8490), .O(N8995) );
or2 gate2387( .a(N4706), .b(N8496), .O(N8996) );
or5 gate2388( .a(N4717), .b(N8500), .c(N8501), .d(N8502), .e(N8503), .O(N9001) );
or2 gate2389( .a(N4728), .b(N8516), .O(N9005) );
and3 gate2390( .a(N7334), .b(N6141), .c(N8537), .O(N9024) );
and3 gate2391( .a(N6137), .b(N7337), .c(N8538), .O(N9025) );
or4 gate2392( .a(N4756), .b(N8545), .c(N8546), .d(N8547), .O(N9029) );
or5 gate2393( .a(N4760), .b(N8551), .c(N8552), .d(N8553), .e(N8554), .O(N9035) );
and3 gate2394( .a(N7378), .b(N6170), .c(N8564), .O(N9053) );
and3 gate2395( .a(N6166), .b(N7381), .c(N8565), .O(N9054) );
nand2 gate2396( .a(N4303), .b(N8607), .O(N9064) );
nand2 gate2397( .a(N3507), .b(N8609), .O(N9065) );
inv1 gate2398( .a(N8114), .O(N9066) );
nand2 gate2399( .a(N8114), .b(N4795), .O(N9067) );
or2 gate2400( .a(N7613), .b(N6783), .O(N9068) );
inv1 gate2401( .a(N8117), .O(N9071) );
inv1 gate2402( .a(N8131), .O(N9072) );
nand2 gate2403( .a(N8131), .b(N6195), .O(N9073) );
inv1 gate2404( .a(N7613), .O(N9074) );
inv1 gate2405( .a(N8134), .O(N9077) );
or2 gate2406( .a(N7650), .b(N6865), .O(N9079) );
inv1 gate2407( .a(N8146), .O(N9082) );
inv1 gate2408( .a(N7650), .O(N9083) );
inv1 gate2409( .a(N8156), .O(N9086) );
inv1 gate2410( .a(N8166), .O(N9087) );

  xor2  gate4998(.a(N4813), .b(N8166), .O(gate2411inter0));
  nand2 gate4999(.a(gate2411inter0), .b(s_212), .O(gate2411inter1));
  and2  gate5000(.a(N4813), .b(N8166), .O(gate2411inter2));
  inv1  gate5001(.a(s_212), .O(gate2411inter3));
  inv1  gate5002(.a(s_213), .O(gate2411inter4));
  nand2 gate5003(.a(gate2411inter4), .b(gate2411inter3), .O(gate2411inter5));
  nor2  gate5004(.a(gate2411inter5), .b(gate2411inter2), .O(gate2411inter6));
  inv1  gate5005(.a(N8166), .O(gate2411inter7));
  inv1  gate5006(.a(N4813), .O(gate2411inter8));
  nand2 gate5007(.a(gate2411inter8), .b(gate2411inter7), .O(gate2411inter9));
  nand2 gate5008(.a(s_213), .b(gate2411inter3), .O(gate2411inter10));
  nor2  gate5009(.a(gate2411inter10), .b(gate2411inter9), .O(gate2411inter11));
  nor2  gate5010(.a(gate2411inter11), .b(gate2411inter6), .O(gate2411inter12));
  nand2 gate5011(.a(gate2411inter12), .b(gate2411inter1), .O(N9088));
or2 gate2412( .a(N7659), .b(N6866), .O(N9089) );
inv1 gate2413( .a(N8169), .O(N9092) );
inv1 gate2414( .a(N8183), .O(N9093) );
nand2 gate2415( .a(N8183), .b(N6203), .O(N9094) );
inv1 gate2416( .a(N7659), .O(N9095) );
inv1 gate2417( .a(N8186), .O(N9098) );
or4 gate2418( .a(N4545), .b(N8340), .c(N8341), .d(N8342), .O(N9099) );
nor3 gate2419( .a(N4545), .b(N8343), .c(N8344), .O(N9103) );
or3 gate2420( .a(N4549), .b(N8345), .c(N8346), .O(N9107) );
nor2 gate2421( .a(N4549), .b(N8347), .O(N9111) );
or4 gate2422( .a(N4577), .b(N8372), .c(N8373), .d(N8374), .O(N9117) );
nor3 gate2423( .a(N4577), .b(N8375), .c(N8376), .O(N9127) );
nor3 gate2424( .a(N4597), .b(N8390), .c(N8391), .O(N9146) );
nor4 gate2425( .a(N4593), .b(N8385), .c(N8386), .d(N8387), .O(N9149) );

  xor2  gate4844(.a(N8733), .b(N7577), .O(gate2426inter0));
  nand2 gate4845(.a(gate2426inter0), .b(s_190), .O(gate2426inter1));
  and2  gate4846(.a(N8733), .b(N7577), .O(gate2426inter2));
  inv1  gate4847(.a(s_190), .O(gate2426inter3));
  inv1  gate4848(.a(s_191), .O(gate2426inter4));
  nand2 gate4849(.a(gate2426inter4), .b(gate2426inter3), .O(gate2426inter5));
  nor2  gate4850(.a(gate2426inter5), .b(gate2426inter2), .O(gate2426inter6));
  inv1  gate4851(.a(N7577), .O(gate2426inter7));
  inv1  gate4852(.a(N8733), .O(gate2426inter8));
  nand2 gate4853(.a(gate2426inter8), .b(gate2426inter7), .O(gate2426inter9));
  nand2 gate4854(.a(s_191), .b(gate2426inter3), .O(gate2426inter10));
  nor2  gate4855(.a(gate2426inter10), .b(gate2426inter9), .O(gate2426inter11));
  nor2  gate4856(.a(gate2426inter11), .b(gate2426inter6), .O(gate2426inter12));
  nand2 gate4857(.a(gate2426inter12), .b(gate2426inter1), .O(N9159));
nand2 gate2427( .a(N7574), .b(N8734), .O(N9160) );
or4 gate2428( .a(N4657), .b(N8436), .c(N8437), .d(N8438), .O(N9161) );
nor3 gate2429( .a(N4657), .b(N8439), .c(N8440), .O(N9165) );
or3 gate2430( .a(N4661), .b(N8441), .c(N8442), .O(N9169) );
nor2 gate2431( .a(N4661), .b(N8443), .O(N9173) );
nand2 gate2432( .a(N7563), .b(N8753), .O(N9179) );
nand2 gate2433( .a(N7560), .b(N8754), .O(N9180) );
nand2 gate2434( .a(N7569), .b(N8755), .O(N9181) );
nand2 gate2435( .a(N7566), .b(N8756), .O(N9182) );
or4 gate2436( .a(N4702), .b(N8491), .c(N8492), .d(N8493), .O(N9183) );
nor3 gate2437( .a(N4702), .b(N8494), .c(N8495), .O(N9193) );
or4 gate2438( .a(N4722), .b(N8511), .c(N8512), .d(N8513), .O(N9203) );
or5 gate2439( .a(N4718), .b(N8504), .c(N8505), .d(N8506), .e(N8507), .O(N9206) );
nor3 gate2440( .a(N4722), .b(N8514), .c(N8515), .O(N9220) );
nor4 gate2441( .a(N4718), .b(N8508), .c(N8509), .d(N8510), .O(N9223) );
nand2 gate2442( .a(N7591), .b(N8814), .O(N9234) );

  xor2  gate5306(.a(N8815), .b(N7588), .O(gate2443inter0));
  nand2 gate5307(.a(gate2443inter0), .b(s_256), .O(gate2443inter1));
  and2  gate5308(.a(N8815), .b(N7588), .O(gate2443inter2));
  inv1  gate5309(.a(s_256), .O(gate2443inter3));
  inv1  gate5310(.a(s_257), .O(gate2443inter4));
  nand2 gate5311(.a(gate2443inter4), .b(gate2443inter3), .O(gate2443inter5));
  nor2  gate5312(.a(gate2443inter5), .b(gate2443inter2), .O(gate2443inter6));
  inv1  gate5313(.a(N7588), .O(gate2443inter7));
  inv1  gate5314(.a(N8815), .O(gate2443inter8));
  nand2 gate5315(.a(gate2443inter8), .b(gate2443inter7), .O(gate2443inter9));
  nand2 gate5316(.a(s_257), .b(gate2443inter3), .O(gate2443inter10));
  nor2  gate5317(.a(gate2443inter10), .b(gate2443inter9), .O(gate2443inter11));
  nor2  gate5318(.a(gate2443inter11), .b(gate2443inter6), .O(gate2443inter12));
  nand2 gate5319(.a(gate2443inter12), .b(gate2443inter1), .O(N9235));
nand2 gate2444( .a(N7585), .b(N8816), .O(N9236) );
nand2 gate2445( .a(N7582), .b(N8817), .O(N9237) );
or2 gate2446( .a(N3159), .b(N8818), .O(N9238) );
or2 gate2447( .a(N3126), .b(N8840), .O(N9242) );
nand2 gate2448( .a(N8324), .b(N8888), .O(N9243) );
inv1 gate2449( .a(N8580), .O(N9244) );
inv1 gate2450( .a(N8583), .O(N9245) );
inv1 gate2451( .a(N8586), .O(N9246) );
inv1 gate2452( .a(N8589), .O(N9247) );
inv1 gate2453( .a(N8592), .O(N9248) );
inv1 gate2454( .a(N8595), .O(N9249) );
inv1 gate2455( .a(N8598), .O(N9250) );
inv1 gate2456( .a(N8601), .O(N9251) );
inv1 gate2457( .a(N8604), .O(N9252) );
nor2 gate2458( .a(N8861), .b(N8280), .O(N9256) );

  xor2  gate3654(.a(N8281), .b(N8862), .O(gate2459inter0));
  nand2 gate3655(.a(gate2459inter0), .b(s_20), .O(gate2459inter1));
  and2  gate3656(.a(N8281), .b(N8862), .O(gate2459inter2));
  inv1  gate3657(.a(s_20), .O(gate2459inter3));
  inv1  gate3658(.a(s_21), .O(gate2459inter4));
  nand2 gate3659(.a(gate2459inter4), .b(gate2459inter3), .O(gate2459inter5));
  nor2  gate3660(.a(gate2459inter5), .b(gate2459inter2), .O(gate2459inter6));
  inv1  gate3661(.a(N8862), .O(gate2459inter7));
  inv1  gate3662(.a(N8281), .O(gate2459inter8));
  nand2 gate3663(.a(gate2459inter8), .b(gate2459inter7), .O(gate2459inter9));
  nand2 gate3664(.a(s_21), .b(gate2459inter3), .O(gate2459inter10));
  nor2  gate3665(.a(gate2459inter10), .b(gate2459inter9), .O(gate2459inter11));
  nor2  gate3666(.a(gate2459inter11), .b(gate2459inter6), .O(gate2459inter12));
  nand2 gate3667(.a(gate2459inter12), .b(gate2459inter1), .O(N9257));
nor2 gate2460( .a(N8863), .b(N8282), .O(N9258) );
nor2 gate2461( .a(N8864), .b(N8283), .O(N9259) );
nor2 gate2462( .a(N8865), .b(N8284), .O(N9260) );
nor2 gate2463( .a(N8866), .b(N8285), .O(N9261) );
inv1 gate2464( .a(N8627), .O(N9262) );
or2 gate2465( .a(N7649), .b(N8874), .O(N9265) );
or2 gate2466( .a(N7668), .b(N8878), .O(N9268) );
nand2 gate2467( .a(N7533), .b(N8879), .O(N9271) );
nand2 gate2468( .a(N7536), .b(N8881), .O(N9272) );
nand2 gate2469( .a(N7539), .b(N8883), .O(N9273) );
nand2 gate2470( .a(N7542), .b(N8885), .O(N9274) );
nand2 gate2471( .a(N8322), .b(N8887), .O(N9275) );
inv1 gate2472( .a(N8333), .O(N9276) );
and5 gate2473( .a(N6936), .b(N8326), .c(N6946), .d(N6929), .e(N6957), .O(N9280) );
and5 gate2474( .a(N367), .b(N8326), .c(N6946), .d(N6957), .e(N6936), .O(N9285) );
and4 gate2475( .a(N367), .b(N8326), .c(N6946), .d(N6957), .O(N9286) );
and3 gate2476( .a(N367), .b(N8326), .c(N6957), .O(N9287) );
and2 gate2477( .a(N367), .b(N8326), .O(N9288) );
inv1 gate2478( .a(N8660), .O(N9290) );
inv1 gate2479( .a(N8663), .O(N9292) );
inv1 gate2480( .a(N8666), .O(N9294) );
inv1 gate2481( .a(N8669), .O(N9296) );
nand2 gate2482( .a(N8672), .b(N5966), .O(N9297) );
inv1 gate2483( .a(N8672), .O(N9298) );
nand2 gate2484( .a(N8675), .b(N6969), .O(N9299) );
inv1 gate2485( .a(N8675), .O(N9300) );
inv1 gate2486( .a(N8365), .O(N9301) );
and5 gate2487( .a(N8358), .b(N7036), .c(N7020), .d(N7006), .e(N6998), .O(N9307) );
and4 gate2488( .a(N8358), .b(N7020), .c(N7006), .d(N7036), .O(N9314) );
and3 gate2489( .a(N8358), .b(N7020), .c(N7036), .O(N9315) );
and2 gate2490( .a(N8358), .b(N7036), .O(N9318) );
inv1 gate2491( .a(N8687), .O(N9319) );
inv1 gate2492( .a(N8699), .O(N9320) );
inv1 gate2493( .a(N8711), .O(N9321) );
inv1 gate2494( .a(N8714), .O(N9322) );
inv1 gate2495( .a(N8727), .O(N9323) );
inv1 gate2496( .a(N8730), .O(N9324) );
inv1 gate2497( .a(N8405), .O(N9326) );
and2 gate2498( .a(N8405), .b(N8412), .O(N9332) );
or2 gate2499( .a(N4193), .b(N8960), .O(N9339) );
and2 gate2500( .a(N8430), .b(N8444), .O(N9344) );
inv1 gate2501( .a(N8735), .O(N9352) );
inv1 gate2502( .a(N8738), .O(N9354) );
inv1 gate2503( .a(N8741), .O(N9356) );
inv1 gate2504( .a(N8744), .O(N9358) );
nand2 gate2505( .a(N8747), .b(N6078), .O(N9359) );
inv1 gate2506( .a(N8747), .O(N9360) );
nand2 gate2507( .a(N8750), .b(N7187), .O(N9361) );
inv1 gate2508( .a(N8750), .O(N9362) );
inv1 gate2509( .a(N8471), .O(N9363) );
inv1 gate2510( .a(N8474), .O(N9364) );
inv1 gate2511( .a(N8477), .O(N9365) );
inv1 gate2512( .a(N8480), .O(N9366) );
nor2 gate2513( .a(N8991), .b(N8483), .O(N9367) );
nor2 gate2514( .a(N8992), .b(N8484), .O(N9368) );
and3 gate2515( .a(N7198), .b(N7194), .c(N8471), .O(N9369) );
and3 gate2516( .a(N8460), .b(N8457), .c(N8474), .O(N9370) );
and3 gate2517( .a(N7209), .b(N7205), .c(N8477), .O(N9371) );
and3 gate2518( .a(N8466), .b(N8463), .c(N8480), .O(N9372) );
inv1 gate2519( .a(N8497), .O(N9375) );
inv1 gate2520( .a(N8766), .O(N9381) );
inv1 gate2521( .a(N8778), .O(N9382) );
inv1 gate2522( .a(N8793), .O(N9383) );
inv1 gate2523( .a(N8796), .O(N9384) );
and2 gate2524( .a(N8485), .b(N8497), .O(N9385) );
inv1 gate2525( .a(N8525), .O(N9392) );
inv1 gate2526( .a(N8528), .O(N9393) );
inv1 gate2527( .a(N8531), .O(N9394) );
inv1 gate2528( .a(N8534), .O(N9395) );
and3 gate2529( .a(N7318), .b(N7314), .c(N8525), .O(N9396) );
and3 gate2530( .a(N8522), .b(N8519), .c(N8528), .O(N9397) );
and3 gate2531( .a(N6131), .b(N6127), .c(N8531), .O(N9398) );
and3 gate2532( .a(N7328), .b(N7325), .c(N8534), .O(N9399) );
nor2 gate2533( .a(N9024), .b(N8539), .O(N9400) );
nor2 gate2534( .a(N9025), .b(N8540), .O(N9401) );
inv1 gate2535( .a(N8541), .O(N9402) );
nand2 gate2536( .a(N8548), .b(N89), .O(N9407) );
and2 gate2537( .a(N8541), .b(N8548), .O(N9408) );
inv1 gate2538( .a(N8811), .O(N9412) );
inv1 gate2539( .a(N8566), .O(N9413) );
inv1 gate2540( .a(N8569), .O(N9414) );
inv1 gate2541( .a(N8572), .O(N9415) );
inv1 gate2542( .a(N8575), .O(N9416) );
nor2 gate2543( .a(N9053), .b(N8578), .O(N9417) );
nor2 gate2544( .a(N9054), .b(N8579), .O(N9418) );
and3 gate2545( .a(N7387), .b(N6177), .c(N8566), .O(N9419) );
and3 gate2546( .a(N8555), .b(N7384), .c(N8569), .O(N9420) );
and3 gate2547( .a(N7398), .b(N7394), .c(N8572), .O(N9421) );
and3 gate2548( .a(N8561), .b(N8558), .c(N8575), .O(N9422) );
buf1 gate2549( .a(N8326), .O(N9423) );
nand2 gate2550( .a(N9064), .b(N8608), .O(N9426) );
nand2 gate2551( .a(N9065), .b(N8610), .O(N9429) );
nand2 gate2552( .a(N3515), .b(N9066), .O(N9432) );
nand2 gate2553( .a(N4796), .b(N9072), .O(N9435) );
nand2 gate2554( .a(N3628), .b(N9087), .O(N9442) );
nand2 gate2555( .a(N4814), .b(N9093), .O(N9445) );
inv1 gate2556( .a(N8678), .O(N9454) );
inv1 gate2557( .a(N8681), .O(N9455) );
inv1 gate2558( .a(N8684), .O(N9456) );
inv1 gate2559( .a(N8690), .O(N9459) );
inv1 gate2560( .a(N8693), .O(N9460) );
inv1 gate2561( .a(N8696), .O(N9461) );
buf1 gate2562( .a(N8358), .O(N9462) );
inv1 gate2563( .a(N8702), .O(N9465) );
inv1 gate2564( .a(N8705), .O(N9466) );
inv1 gate2565( .a(N8708), .O(N9467) );
inv1 gate2566( .a(N8724), .O(N9468) );
buf1 gate2567( .a(N8358), .O(N9473) );
inv1 gate2568( .a(N8718), .O(N9476) );
inv1 gate2569( .a(N8721), .O(N9477) );
nand2 gate2570( .a(N9159), .b(N9160), .O(N9478) );

  xor2  gate3752(.a(N9180), .b(N9179), .O(gate2571inter0));
  nand2 gate3753(.a(gate2571inter0), .b(s_34), .O(gate2571inter1));
  and2  gate3754(.a(N9180), .b(N9179), .O(gate2571inter2));
  inv1  gate3755(.a(s_34), .O(gate2571inter3));
  inv1  gate3756(.a(s_35), .O(gate2571inter4));
  nand2 gate3757(.a(gate2571inter4), .b(gate2571inter3), .O(gate2571inter5));
  nor2  gate3758(.a(gate2571inter5), .b(gate2571inter2), .O(gate2571inter6));
  inv1  gate3759(.a(N9179), .O(gate2571inter7));
  inv1  gate3760(.a(N9180), .O(gate2571inter8));
  nand2 gate3761(.a(gate2571inter8), .b(gate2571inter7), .O(gate2571inter9));
  nand2 gate3762(.a(s_35), .b(gate2571inter3), .O(gate2571inter10));
  nor2  gate3763(.a(gate2571inter10), .b(gate2571inter9), .O(gate2571inter11));
  nor2  gate3764(.a(gate2571inter11), .b(gate2571inter6), .O(gate2571inter12));
  nand2 gate3765(.a(gate2571inter12), .b(gate2571inter1), .O(N9485));

  xor2  gate4046(.a(N9182), .b(N9181), .O(gate2572inter0));
  nand2 gate4047(.a(gate2572inter0), .b(s_76), .O(gate2572inter1));
  and2  gate4048(.a(N9182), .b(N9181), .O(gate2572inter2));
  inv1  gate4049(.a(s_76), .O(gate2572inter3));
  inv1  gate4050(.a(s_77), .O(gate2572inter4));
  nand2 gate4051(.a(gate2572inter4), .b(gate2572inter3), .O(gate2572inter5));
  nor2  gate4052(.a(gate2572inter5), .b(gate2572inter2), .O(gate2572inter6));
  inv1  gate4053(.a(N9181), .O(gate2572inter7));
  inv1  gate4054(.a(N9182), .O(gate2572inter8));
  nand2 gate4055(.a(gate2572inter8), .b(gate2572inter7), .O(gate2572inter9));
  nand2 gate4056(.a(s_77), .b(gate2572inter3), .O(gate2572inter10));
  nor2  gate4057(.a(gate2572inter10), .b(gate2572inter9), .O(gate2572inter11));
  nor2  gate4058(.a(gate2572inter11), .b(gate2572inter6), .O(gate2572inter12));
  nand2 gate4059(.a(gate2572inter12), .b(gate2572inter1), .O(N9488));
inv1 gate2573( .a(N8757), .O(N9493) );
inv1 gate2574( .a(N8760), .O(N9494) );
inv1 gate2575( .a(N8763), .O(N9495) );
inv1 gate2576( .a(N8769), .O(N9498) );
inv1 gate2577( .a(N8772), .O(N9499) );
inv1 gate2578( .a(N8775), .O(N9500) );
inv1 gate2579( .a(N8781), .O(N9505) );
inv1 gate2580( .a(N8784), .O(N9506) );
inv1 gate2581( .a(N8787), .O(N9507) );
inv1 gate2582( .a(N8790), .O(N9508) );
inv1 gate2583( .a(N8808), .O(N9509) );
inv1 gate2584( .a(N8799), .O(N9514) );
inv1 gate2585( .a(N8802), .O(N9515) );
inv1 gate2586( .a(N8805), .O(N9516) );
nand2 gate2587( .a(N9234), .b(N9235), .O(N9517) );
nand2 gate2588( .a(N9236), .b(N9237), .O(N9520) );
and2 gate2589( .a(N8943), .b(N8421), .O(N9526) );
and2 gate2590( .a(N8943), .b(N8421), .O(N9531) );
nand2 gate2591( .a(N9271), .b(N8880), .O(N9539) );
nand2 gate2592( .a(N9273), .b(N8884), .O(N9540) );
inv1 gate2593( .a(N9275), .O(N9541) );
and2 gate2594( .a(N8857), .b(N8254), .O(N9543) );
and2 gate2595( .a(N8871), .b(N8288), .O(N9551) );
nand2 gate2596( .a(N9272), .b(N8882), .O(N9555) );
nand2 gate2597( .a(N9274), .b(N8886), .O(N9556) );
inv1 gate2598( .a(N8898), .O(N9557) );
and2 gate2599( .a(N8902), .b(N8333), .O(N9560) );
inv1 gate2600( .a(N9099), .O(N9561) );
nand2 gate2601( .a(N9099), .b(N9290), .O(N9562) );
inv1 gate2602( .a(N9103), .O(N9563) );
nand2 gate2603( .a(N9103), .b(N9292), .O(N9564) );
inv1 gate2604( .a(N9107), .O(N9565) );
nand2 gate2605( .a(N9107), .b(N9294), .O(N9566) );
inv1 gate2606( .a(N9111), .O(N9567) );
nand2 gate2607( .a(N9111), .b(N9296), .O(N9568) );
nand2 gate2608( .a(N4844), .b(N9298), .O(N9569) );
nand2 gate2609( .a(N6207), .b(N9300), .O(N9570) );
inv1 gate2610( .a(N8920), .O(N9571) );
inv1 gate2611( .a(N8927), .O(N9575) );
and2 gate2612( .a(N8365), .b(N8927), .O(N9579) );
inv1 gate2613( .a(N8950), .O(N9581) );
inv1 gate2614( .a(N8956), .O(N9582) );
and2 gate2615( .a(N8405), .b(N8956), .O(N9585) );
and2 gate2616( .a(N8966), .b(N8430), .O(N9591) );
inv1 gate2617( .a(N9161), .O(N9592) );
nand2 gate2618( .a(N9161), .b(N9352), .O(N9593) );
inv1 gate2619( .a(N9165), .O(N9594) );

  xor2  gate4354(.a(N9354), .b(N9165), .O(gate2620inter0));
  nand2 gate4355(.a(gate2620inter0), .b(s_120), .O(gate2620inter1));
  and2  gate4356(.a(N9354), .b(N9165), .O(gate2620inter2));
  inv1  gate4357(.a(s_120), .O(gate2620inter3));
  inv1  gate4358(.a(s_121), .O(gate2620inter4));
  nand2 gate4359(.a(gate2620inter4), .b(gate2620inter3), .O(gate2620inter5));
  nor2  gate4360(.a(gate2620inter5), .b(gate2620inter2), .O(gate2620inter6));
  inv1  gate4361(.a(N9165), .O(gate2620inter7));
  inv1  gate4362(.a(N9354), .O(gate2620inter8));
  nand2 gate4363(.a(gate2620inter8), .b(gate2620inter7), .O(gate2620inter9));
  nand2 gate4364(.a(s_121), .b(gate2620inter3), .O(gate2620inter10));
  nor2  gate4365(.a(gate2620inter10), .b(gate2620inter9), .O(gate2620inter11));
  nor2  gate4366(.a(gate2620inter11), .b(gate2620inter6), .O(gate2620inter12));
  nand2 gate4367(.a(gate2620inter12), .b(gate2620inter1), .O(N9595));
inv1 gate2621( .a(N9169), .O(N9596) );
nand2 gate2622( .a(N9169), .b(N9356), .O(N9597) );
inv1 gate2623( .a(N9173), .O(N9598) );
nand2 gate2624( .a(N9173), .b(N9358), .O(N9599) );
nand2 gate2625( .a(N4940), .b(N9360), .O(N9600) );
nand2 gate2626( .a(N6220), .b(N9362), .O(N9601) );
and3 gate2627( .a(N8457), .b(N7198), .c(N9363), .O(N9602) );
and3 gate2628( .a(N7194), .b(N8460), .c(N9364), .O(N9603) );
and3 gate2629( .a(N8463), .b(N7209), .c(N9365), .O(N9604) );
and3 gate2630( .a(N7205), .b(N8466), .c(N9366), .O(N9605) );
inv1 gate2631( .a(N9001), .O(N9608) );
and2 gate2632( .a(N8485), .b(N9001), .O(N9611) );
and3 gate2633( .a(N8519), .b(N7318), .c(N9392), .O(N9612) );
and3 gate2634( .a(N7314), .b(N8522), .c(N9393), .O(N9613) );
and3 gate2635( .a(N7325), .b(N6131), .c(N9394), .O(N9614) );
and3 gate2636( .a(N6127), .b(N7328), .c(N9395), .O(N9615) );
inv1 gate2637( .a(N9029), .O(N9616) );
inv1 gate2638( .a(N9035), .O(N9617) );
and2 gate2639( .a(N8541), .b(N9035), .O(N9618) );
and3 gate2640( .a(N7384), .b(N7387), .c(N9413), .O(N9621) );
and3 gate2641( .a(N6177), .b(N8555), .c(N9414), .O(N9622) );
and3 gate2642( .a(N8558), .b(N7398), .c(N9415), .O(N9623) );
and3 gate2643( .a(N7394), .b(N8561), .c(N9416), .O(N9624) );
or5 gate2644( .a(N4563), .b(N8352), .c(N8353), .d(N8354), .e(N9285), .O(N9626) );
or4 gate2645( .a(N4566), .b(N8355), .c(N8356), .d(N9286), .O(N9629) );
or3 gate2646( .a(N4570), .b(N8357), .c(N9287), .O(N9632) );
or2 gate2647( .a(N5960), .b(N9288), .O(N9635) );
nand2 gate2648( .a(N9067), .b(N9432), .O(N9642) );
inv1 gate2649( .a(N9068), .O(N9645) );
nand2 gate2650( .a(N9073), .b(N9435), .O(N9646) );
inv1 gate2651( .a(N9074), .O(N9649) );
nand2 gate2652( .a(N9257), .b(N9256), .O(N9650) );

  xor2  gate3864(.a(N9258), .b(N9259), .O(gate2653inter0));
  nand2 gate3865(.a(gate2653inter0), .b(s_50), .O(gate2653inter1));
  and2  gate3866(.a(N9258), .b(N9259), .O(gate2653inter2));
  inv1  gate3867(.a(s_50), .O(gate2653inter3));
  inv1  gate3868(.a(s_51), .O(gate2653inter4));
  nand2 gate3869(.a(gate2653inter4), .b(gate2653inter3), .O(gate2653inter5));
  nor2  gate3870(.a(gate2653inter5), .b(gate2653inter2), .O(gate2653inter6));
  inv1  gate3871(.a(N9259), .O(gate2653inter7));
  inv1  gate3872(.a(N9258), .O(gate2653inter8));
  nand2 gate3873(.a(gate2653inter8), .b(gate2653inter7), .O(gate2653inter9));
  nand2 gate3874(.a(s_51), .b(gate2653inter3), .O(gate2653inter10));
  nor2  gate3875(.a(gate2653inter10), .b(gate2653inter9), .O(gate2653inter11));
  nor2  gate3876(.a(gate2653inter11), .b(gate2653inter6), .O(gate2653inter12));
  nand2 gate3877(.a(gate2653inter12), .b(gate2653inter1), .O(N9653));
nand2 gate2654( .a(N9261), .b(N9260), .O(N9656) );
inv1 gate2655( .a(N9079), .O(N9659) );

  xor2  gate4900(.a(N4809), .b(N9079), .O(gate2656inter0));
  nand2 gate4901(.a(gate2656inter0), .b(s_198), .O(gate2656inter1));
  and2  gate4902(.a(N4809), .b(N9079), .O(gate2656inter2));
  inv1  gate4903(.a(s_198), .O(gate2656inter3));
  inv1  gate4904(.a(s_199), .O(gate2656inter4));
  nand2 gate4905(.a(gate2656inter4), .b(gate2656inter3), .O(gate2656inter5));
  nor2  gate4906(.a(gate2656inter5), .b(gate2656inter2), .O(gate2656inter6));
  inv1  gate4907(.a(N9079), .O(gate2656inter7));
  inv1  gate4908(.a(N4809), .O(gate2656inter8));
  nand2 gate4909(.a(gate2656inter8), .b(gate2656inter7), .O(gate2656inter9));
  nand2 gate4910(.a(s_199), .b(gate2656inter3), .O(gate2656inter10));
  nor2  gate4911(.a(gate2656inter10), .b(gate2656inter9), .O(gate2656inter11));
  nor2  gate4912(.a(gate2656inter11), .b(gate2656inter6), .O(gate2656inter12));
  nand2 gate4913(.a(gate2656inter12), .b(gate2656inter1), .O(N9660));
inv1 gate2657( .a(N9083), .O(N9661) );
nand2 gate2658( .a(N9083), .b(N6202), .O(N9662) );
nand2 gate2659( .a(N9088), .b(N9442), .O(N9663) );
inv1 gate2660( .a(N9089), .O(N9666) );

  xor2  gate4312(.a(N9445), .b(N9094), .O(gate2661inter0));
  nand2 gate4313(.a(gate2661inter0), .b(s_114), .O(gate2661inter1));
  and2  gate4314(.a(N9445), .b(N9094), .O(gate2661inter2));
  inv1  gate4315(.a(s_114), .O(gate2661inter3));
  inv1  gate4316(.a(s_115), .O(gate2661inter4));
  nand2 gate4317(.a(gate2661inter4), .b(gate2661inter3), .O(gate2661inter5));
  nor2  gate4318(.a(gate2661inter5), .b(gate2661inter2), .O(gate2661inter6));
  inv1  gate4319(.a(N9094), .O(gate2661inter7));
  inv1  gate4320(.a(N9445), .O(gate2661inter8));
  nand2 gate4321(.a(gate2661inter8), .b(gate2661inter7), .O(gate2661inter9));
  nand2 gate4322(.a(s_115), .b(gate2661inter3), .O(gate2661inter10));
  nor2  gate4323(.a(gate2661inter10), .b(gate2661inter9), .O(gate2661inter11));
  nor2  gate4324(.a(gate2661inter11), .b(gate2661inter6), .O(gate2661inter12));
  nand2 gate4325(.a(gate2661inter12), .b(gate2661inter1), .O(N9667));
inv1 gate2662( .a(N9095), .O(N9670) );
or2 gate2663( .a(N8924), .b(N8393), .O(N9671) );
inv1 gate2664( .a(N9117), .O(N9674) );
inv1 gate2665( .a(N8924), .O(N9675) );
inv1 gate2666( .a(N9127), .O(N9678) );
or4 gate2667( .a(N4597), .b(N8388), .c(N8389), .d(N9315), .O(N9679) );
or2 gate2668( .a(N8931), .b(N9318), .O(N9682) );
or5 gate2669( .a(N4593), .b(N8382), .c(N8383), .d(N8384), .e(N9314), .O(N9685) );
inv1 gate2670( .a(N9146), .O(N9690) );
nand2 gate2671( .a(N9146), .b(N8717), .O(N9691) );
inv1 gate2672( .a(N8931), .O(N9692) );
inv1 gate2673( .a(N9149), .O(N9695) );
nand2 gate2674( .a(N9401), .b(N9400), .O(N9698) );
nand2 gate2675( .a(N9368), .b(N9367), .O(N9702) );
or2 gate2676( .a(N8996), .b(N8517), .O(N9707) );
inv1 gate2677( .a(N9183), .O(N9710) );
inv1 gate2678( .a(N8996), .O(N9711) );
inv1 gate2679( .a(N9193), .O(N9714) );
inv1 gate2680( .a(N9203), .O(N9715) );
nand2 gate2681( .a(N9203), .b(N6235), .O(N9716) );
or2 gate2682( .a(N9005), .b(N8518), .O(N9717) );
inv1 gate2683( .a(N9206), .O(N9720) );
inv1 gate2684( .a(N9220), .O(N9721) );
nand2 gate2685( .a(N9220), .b(N7573), .O(N9722) );
inv1 gate2686( .a(N9005), .O(N9723) );
inv1 gate2687( .a(N9223), .O(N9726) );
nand2 gate2688( .a(N9418), .b(N9417), .O(N9727) );
and2 gate2689( .a(N9268), .b(N8269), .O(N9732) );
nand2 gate2690( .a(N9581), .b(N9326), .O(N9733) );
and5 gate2691( .a(N89), .b(N9408), .c(N9332), .d(N8394), .e(N8421), .O(N9734) );
and5 gate2692( .a(N89), .b(N9408), .c(N9332), .d(N8394), .e(N8421), .O(N9735) );
and2 gate2693( .a(N9265), .b(N8262), .O(N9736) );
inv1 gate2694( .a(N9555), .O(N9737) );
inv1 gate2695( .a(N9556), .O(N9738) );

  xor2  gate4214(.a(N9601), .b(N9361), .O(gate2696inter0));
  nand2 gate4215(.a(gate2696inter0), .b(s_100), .O(gate2696inter1));
  and2  gate4216(.a(N9601), .b(N9361), .O(gate2696inter2));
  inv1  gate4217(.a(s_100), .O(gate2696inter3));
  inv1  gate4218(.a(s_101), .O(gate2696inter4));
  nand2 gate4219(.a(gate2696inter4), .b(gate2696inter3), .O(gate2696inter5));
  nor2  gate4220(.a(gate2696inter5), .b(gate2696inter2), .O(gate2696inter6));
  inv1  gate4221(.a(N9361), .O(gate2696inter7));
  inv1  gate4222(.a(N9601), .O(gate2696inter8));
  nand2 gate4223(.a(gate2696inter8), .b(gate2696inter7), .O(gate2696inter9));
  nand2 gate4224(.a(s_101), .b(gate2696inter3), .O(gate2696inter10));
  nor2  gate4225(.a(gate2696inter10), .b(gate2696inter9), .O(gate2696inter11));
  nor2  gate4226(.a(gate2696inter11), .b(gate2696inter6), .O(gate2696inter12));
  nand2 gate4227(.a(gate2696inter12), .b(gate2696inter1), .O(N9739));
nand2 gate2697( .a(N9423), .b(N1115), .O(N9740) );
inv1 gate2698( .a(N9423), .O(N9741) );
nand2 gate2699( .a(N9299), .b(N9570), .O(N9742) );
and2 gate2700( .a(N8333), .b(N9280), .O(N9754) );
or2 gate2701( .a(N8898), .b(N9560), .O(N9758) );
nand2 gate2702( .a(N8660), .b(N9561), .O(N9762) );
nand2 gate2703( .a(N8663), .b(N9563), .O(N9763) );
nand2 gate2704( .a(N8666), .b(N9565), .O(N9764) );
nand2 gate2705( .a(N8669), .b(N9567), .O(N9765) );
nand2 gate2706( .a(N9297), .b(N9569), .O(N9766) );
and2 gate2707( .a(N9280), .b(N367), .O(N9767) );
nand2 gate2708( .a(N9557), .b(N9276), .O(N9768) );
inv1 gate2709( .a(N9307), .O(N9769) );
nand2 gate2710( .a(N9307), .b(N367), .O(N9773) );
nand2 gate2711( .a(N9571), .b(N9301), .O(N9774) );
and2 gate2712( .a(N8365), .b(N9307), .O(N9775) );
or2 gate2713( .a(N8920), .b(N9579), .O(N9779) );
inv1 gate2714( .a(N9478), .O(N9784) );

  xor2  gate4298(.a(N9402), .b(N9616), .O(gate2715inter0));
  nand2 gate4299(.a(gate2715inter0), .b(s_112), .O(gate2715inter1));
  and2  gate4300(.a(N9402), .b(N9616), .O(gate2715inter2));
  inv1  gate4301(.a(s_112), .O(gate2715inter3));
  inv1  gate4302(.a(s_113), .O(gate2715inter4));
  nand2 gate4303(.a(gate2715inter4), .b(gate2715inter3), .O(gate2715inter5));
  nor2  gate4304(.a(gate2715inter5), .b(gate2715inter2), .O(gate2715inter6));
  inv1  gate4305(.a(N9616), .O(gate2715inter7));
  inv1  gate4306(.a(N9402), .O(gate2715inter8));
  nand2 gate4307(.a(gate2715inter8), .b(gate2715inter7), .O(gate2715inter9));
  nand2 gate4308(.a(s_113), .b(gate2715inter3), .O(gate2715inter10));
  nor2  gate4309(.a(gate2715inter10), .b(gate2715inter9), .O(gate2715inter11));
  nor2  gate4310(.a(gate2715inter11), .b(gate2715inter6), .O(gate2715inter12));
  nand2 gate4311(.a(gate2715inter12), .b(gate2715inter1), .O(N9785));
or2 gate2716( .a(N8950), .b(N9585), .O(N9786) );
and4 gate2717( .a(N89), .b(N9408), .c(N9332), .d(N8394), .O(N9790) );
or2 gate2718( .a(N8963), .b(N9591), .O(N9791) );
nand2 gate2719( .a(N8735), .b(N9592), .O(N9795) );
nand2 gate2720( .a(N8738), .b(N9594), .O(N9796) );
nand2 gate2721( .a(N8741), .b(N9596), .O(N9797) );
nand2 gate2722( .a(N8744), .b(N9598), .O(N9798) );
nand2 gate2723( .a(N9359), .b(N9600), .O(N9799) );
nor2 gate2724( .a(N9602), .b(N9369), .O(N9800) );
nor2 gate2725( .a(N9603), .b(N9370), .O(N9801) );
nor2 gate2726( .a(N9604), .b(N9371), .O(N9802) );
nor2 gate2727( .a(N9605), .b(N9372), .O(N9803) );
inv1 gate2728( .a(N9485), .O(N9805) );
inv1 gate2729( .a(N9488), .O(N9806) );
or2 gate2730( .a(N8995), .b(N9611), .O(N9809) );
nor2 gate2731( .a(N9612), .b(N9396), .O(N9813) );
nor2 gate2732( .a(N9613), .b(N9397), .O(N9814) );
nor2 gate2733( .a(N9614), .b(N9398), .O(N9815) );
nor2 gate2734( .a(N9615), .b(N9399), .O(N9816) );
and2 gate2735( .a(N9617), .b(N9407), .O(N9817) );
or2 gate2736( .a(N9029), .b(N9618), .O(N9820) );
inv1 gate2737( .a(N9517), .O(N9825) );
inv1 gate2738( .a(N9520), .O(N9826) );
nor2 gate2739( .a(N9621), .b(N9419), .O(N9827) );
nor2 gate2740( .a(N9622), .b(N9420), .O(N9828) );
nor2 gate2741( .a(N9623), .b(N9421), .O(N9829) );
nor2 gate2742( .a(N9624), .b(N9422), .O(N9830) );
inv1 gate2743( .a(N9426), .O(N9835) );
nand2 gate2744( .a(N9426), .b(N4789), .O(N9836) );
inv1 gate2745( .a(N9429), .O(N9837) );
nand2 gate2746( .a(N9429), .b(N4794), .O(N9838) );

  xor2  gate3920(.a(N9659), .b(N3625), .O(gate2747inter0));
  nand2 gate3921(.a(gate2747inter0), .b(s_58), .O(gate2747inter1));
  and2  gate3922(.a(N9659), .b(N3625), .O(gate2747inter2));
  inv1  gate3923(.a(s_58), .O(gate2747inter3));
  inv1  gate3924(.a(s_59), .O(gate2747inter4));
  nand2 gate3925(.a(gate2747inter4), .b(gate2747inter3), .O(gate2747inter5));
  nor2  gate3926(.a(gate2747inter5), .b(gate2747inter2), .O(gate2747inter6));
  inv1  gate3927(.a(N3625), .O(gate2747inter7));
  inv1  gate3928(.a(N9659), .O(gate2747inter8));
  nand2 gate3929(.a(gate2747inter8), .b(gate2747inter7), .O(gate2747inter9));
  nand2 gate3930(.a(s_59), .b(gate2747inter3), .O(gate2747inter10));
  nor2  gate3931(.a(gate2747inter10), .b(gate2747inter9), .O(gate2747inter11));
  nor2  gate3932(.a(gate2747inter11), .b(gate2747inter6), .O(gate2747inter12));
  nand2 gate3933(.a(gate2747inter12), .b(gate2747inter1), .O(N9846));
nand2 gate2748( .a(N4810), .b(N9661), .O(N9847) );
inv1 gate2749( .a(N9462), .O(N9862) );
nand2 gate2750( .a(N7553), .b(N9690), .O(N9863) );
inv1 gate2751( .a(N9473), .O(N9866) );
nand2 gate2752( .a(N5030), .b(N9715), .O(N9873) );
nand2 gate2753( .a(N6236), .b(N9721), .O(N9876) );
nand2 gate2754( .a(N9795), .b(N9593), .O(N9890) );
nand2 gate2755( .a(N9797), .b(N9597), .O(N9891) );
inv1 gate2756( .a(N9799), .O(N9892) );

  xor2  gate4088(.a(N9741), .b(N871), .O(gate2757inter0));
  nand2 gate4089(.a(gate2757inter0), .b(s_82), .O(gate2757inter1));
  and2  gate4090(.a(N9741), .b(N871), .O(gate2757inter2));
  inv1  gate4091(.a(s_82), .O(gate2757inter3));
  inv1  gate4092(.a(s_83), .O(gate2757inter4));
  nand2 gate4093(.a(gate2757inter4), .b(gate2757inter3), .O(gate2757inter5));
  nor2  gate4094(.a(gate2757inter5), .b(gate2757inter2), .O(gate2757inter6));
  inv1  gate4095(.a(N871), .O(gate2757inter7));
  inv1  gate4096(.a(N9741), .O(gate2757inter8));
  nand2 gate4097(.a(gate2757inter8), .b(gate2757inter7), .O(gate2757inter9));
  nand2 gate4098(.a(s_83), .b(gate2757inter3), .O(gate2757inter10));
  nor2  gate4099(.a(gate2757inter10), .b(gate2757inter9), .O(gate2757inter11));
  nor2  gate4100(.a(gate2757inter11), .b(gate2757inter6), .O(gate2757inter12));
  nand2 gate4101(.a(gate2757inter12), .b(gate2757inter1), .O(N9893));
nand2 gate2758( .a(N9762), .b(N9562), .O(N9894) );
nand2 gate2759( .a(N9764), .b(N9566), .O(N9895) );
inv1 gate2760( .a(N9766), .O(N9896) );
inv1 gate2761( .a(N9626), .O(N9897) );
nand2 gate2762( .a(N9626), .b(N9249), .O(N9898) );
inv1 gate2763( .a(N9629), .O(N9899) );
nand2 gate2764( .a(N9629), .b(N9250), .O(N9900) );
inv1 gate2765( .a(N9632), .O(N9901) );
nand2 gate2766( .a(N9632), .b(N9251), .O(N9902) );
inv1 gate2767( .a(N9635), .O(N9903) );
nand2 gate2768( .a(N9635), .b(N9252), .O(N9904) );
inv1 gate2769( .a(N9543), .O(N9905) );
inv1 gate2770( .a(N9650), .O(N9906) );
nand2 gate2771( .a(N9650), .b(N5769), .O(N9907) );
inv1 gate2772( .a(N9653), .O(N9908) );
nand2 gate2773( .a(N9653), .b(N5770), .O(N9909) );
inv1 gate2774( .a(N9656), .O(N9910) );
nand2 gate2775( .a(N9656), .b(N9262), .O(N9911) );
inv1 gate2776( .a(N9551), .O(N9917) );
nand2 gate2777( .a(N9763), .b(N9564), .O(N9923) );
nand2 gate2778( .a(N9765), .b(N9568), .O(N9924) );
or2 gate2779( .a(N8902), .b(N9767), .O(N9925) );
and2 gate2780( .a(N9575), .b(N9773), .O(N9932) );
and2 gate2781( .a(N9575), .b(N9769), .O(N9935) );
inv1 gate2782( .a(N9698), .O(N9938) );
nand2 gate2783( .a(N9698), .b(N9323), .O(N9939) );
nand2 gate2784( .a(N9796), .b(N9595), .O(N9945) );
nand2 gate2785( .a(N9798), .b(N9599), .O(N9946) );
inv1 gate2786( .a(N9702), .O(N9947) );
nand2 gate2787( .a(N9702), .b(N6102), .O(N9948) );
and2 gate2788( .a(N9608), .b(N9375), .O(N9949) );
inv1 gate2789( .a(N9727), .O(N9953) );
nand2 gate2790( .a(N9727), .b(N9412), .O(N9954) );
nand2 gate2791( .a(N3502), .b(N9835), .O(N9955) );
nand2 gate2792( .a(N3510), .b(N9837), .O(N9956) );
inv1 gate2793( .a(N9642), .O(N9957) );
nand2 gate2794( .a(N9642), .b(N9645), .O(N9958) );
inv1 gate2795( .a(N9646), .O(N9959) );

  xor2  gate4648(.a(N9649), .b(N9646), .O(gate2796inter0));
  nand2 gate4649(.a(gate2796inter0), .b(s_162), .O(gate2796inter1));
  and2  gate4650(.a(N9649), .b(N9646), .O(gate2796inter2));
  inv1  gate4651(.a(s_162), .O(gate2796inter3));
  inv1  gate4652(.a(s_163), .O(gate2796inter4));
  nand2 gate4653(.a(gate2796inter4), .b(gate2796inter3), .O(gate2796inter5));
  nor2  gate4654(.a(gate2796inter5), .b(gate2796inter2), .O(gate2796inter6));
  inv1  gate4655(.a(N9646), .O(gate2796inter7));
  inv1  gate4656(.a(N9649), .O(gate2796inter8));
  nand2 gate4657(.a(gate2796inter8), .b(gate2796inter7), .O(gate2796inter9));
  nand2 gate4658(.a(s_163), .b(gate2796inter3), .O(gate2796inter10));
  nor2  gate4659(.a(gate2796inter10), .b(gate2796inter9), .O(gate2796inter11));
  nor2  gate4660(.a(gate2796inter11), .b(gate2796inter6), .O(gate2796inter12));
  nand2 gate4661(.a(gate2796inter12), .b(gate2796inter1), .O(N9960));

  xor2  gate5334(.a(N9846), .b(N9660), .O(gate2797inter0));
  nand2 gate5335(.a(gate2797inter0), .b(s_260), .O(gate2797inter1));
  and2  gate5336(.a(N9846), .b(N9660), .O(gate2797inter2));
  inv1  gate5337(.a(s_260), .O(gate2797inter3));
  inv1  gate5338(.a(s_261), .O(gate2797inter4));
  nand2 gate5339(.a(gate2797inter4), .b(gate2797inter3), .O(gate2797inter5));
  nor2  gate5340(.a(gate2797inter5), .b(gate2797inter2), .O(gate2797inter6));
  inv1  gate5341(.a(N9660), .O(gate2797inter7));
  inv1  gate5342(.a(N9846), .O(gate2797inter8));
  nand2 gate5343(.a(gate2797inter8), .b(gate2797inter7), .O(gate2797inter9));
  nand2 gate5344(.a(s_261), .b(gate2797inter3), .O(gate2797inter10));
  nor2  gate5345(.a(gate2797inter10), .b(gate2797inter9), .O(gate2797inter11));
  nor2  gate5346(.a(gate2797inter11), .b(gate2797inter6), .O(gate2797inter12));
  nand2 gate5347(.a(gate2797inter12), .b(gate2797inter1), .O(N9961));
nand2 gate2798( .a(N9662), .b(N9847), .O(N9964) );
inv1 gate2799( .a(N9663), .O(N9967) );
nand2 gate2800( .a(N9663), .b(N9666), .O(N9968) );
inv1 gate2801( .a(N9667), .O(N9969) );

  xor2  gate4550(.a(N9670), .b(N9667), .O(gate2802inter0));
  nand2 gate4551(.a(gate2802inter0), .b(s_148), .O(gate2802inter1));
  and2  gate4552(.a(N9670), .b(N9667), .O(gate2802inter2));
  inv1  gate4553(.a(s_148), .O(gate2802inter3));
  inv1  gate4554(.a(s_149), .O(gate2802inter4));
  nand2 gate4555(.a(gate2802inter4), .b(gate2802inter3), .O(gate2802inter5));
  nor2  gate4556(.a(gate2802inter5), .b(gate2802inter2), .O(gate2802inter6));
  inv1  gate4557(.a(N9667), .O(gate2802inter7));
  inv1  gate4558(.a(N9670), .O(gate2802inter8));
  nand2 gate4559(.a(gate2802inter8), .b(gate2802inter7), .O(gate2802inter9));
  nand2 gate4560(.a(s_149), .b(gate2802inter3), .O(gate2802inter10));
  nor2  gate4561(.a(gate2802inter10), .b(gate2802inter9), .O(gate2802inter11));
  nor2  gate4562(.a(gate2802inter11), .b(gate2802inter6), .O(gate2802inter12));
  nand2 gate4563(.a(gate2802inter12), .b(gate2802inter1), .O(N9970));
inv1 gate2803( .a(N9671), .O(N9971) );
nand2 gate2804( .a(N9671), .b(N6213), .O(N9972) );
inv1 gate2805( .a(N9675), .O(N9973) );
nand2 gate2806( .a(N9675), .b(N7551), .O(N9974) );
inv1 gate2807( .a(N9679), .O(N9975) );
nand2 gate2808( .a(N9679), .b(N7552), .O(N9976) );
inv1 gate2809( .a(N9682), .O(N9977) );
inv1 gate2810( .a(N9685), .O(N9978) );
nand2 gate2811( .a(N9691), .b(N9863), .O(N9979) );
inv1 gate2812( .a(N9692), .O(N9982) );
nand2 gate2813( .a(N9814), .b(N9813), .O(N9983) );
nand2 gate2814( .a(N9816), .b(N9815), .O(N9986) );
nand2 gate2815( .a(N9801), .b(N9800), .O(N9989) );
nand2 gate2816( .a(N9803), .b(N9802), .O(N9992) );
inv1 gate2817( .a(N9707), .O(N9995) );
nand2 gate2818( .a(N9707), .b(N6231), .O(N9996) );
inv1 gate2819( .a(N9711), .O(N9997) );
nand2 gate2820( .a(N9711), .b(N7572), .O(N9998) );
nand2 gate2821( .a(N9716), .b(N9873), .O(N9999) );
inv1 gate2822( .a(N9717), .O(N10002) );

  xor2  gate5236(.a(N9876), .b(N9722), .O(gate2823inter0));
  nand2 gate5237(.a(gate2823inter0), .b(s_246), .O(gate2823inter1));
  and2  gate5238(.a(N9876), .b(N9722), .O(gate2823inter2));
  inv1  gate5239(.a(s_246), .O(gate2823inter3));
  inv1  gate5240(.a(s_247), .O(gate2823inter4));
  nand2 gate5241(.a(gate2823inter4), .b(gate2823inter3), .O(gate2823inter5));
  nor2  gate5242(.a(gate2823inter5), .b(gate2823inter2), .O(gate2823inter6));
  inv1  gate5243(.a(N9722), .O(gate2823inter7));
  inv1  gate5244(.a(N9876), .O(gate2823inter8));
  nand2 gate5245(.a(gate2823inter8), .b(gate2823inter7), .O(gate2823inter9));
  nand2 gate5246(.a(s_247), .b(gate2823inter3), .O(gate2823inter10));
  nor2  gate5247(.a(gate2823inter10), .b(gate2823inter9), .O(gate2823inter11));
  nor2  gate5248(.a(gate2823inter11), .b(gate2823inter6), .O(gate2823inter12));
  nand2 gate5249(.a(gate2823inter12), .b(gate2823inter1), .O(N10003));
inv1 gate2824( .a(N9723), .O(N10006) );
nand2 gate2825( .a(N9830), .b(N9829), .O(N10007) );
nand2 gate2826( .a(N9828), .b(N9827), .O(N10010) );
and3 gate2827( .a(N9791), .b(N8307), .c(N8269), .O(N10013) );
and4 gate2828( .a(N9758), .b(N9344), .c(N8307), .d(N8269), .O(N10014) );
and5 gate2829( .a(N367), .b(N9754), .c(N9344), .d(N8307), .e(N8269), .O(N10015) );
and3 gate2830( .a(N9786), .b(N8394), .c(N8421), .O(N10016) );
and4 gate2831( .a(N9820), .b(N9332), .c(N8394), .d(N8421), .O(N10017) );
and3 gate2832( .a(N9786), .b(N8394), .c(N8421), .O(N10018) );
and4 gate2833( .a(N9820), .b(N9332), .c(N8394), .d(N8421), .O(N10019) );
and3 gate2834( .a(N9809), .b(N8298), .c(N8262), .O(N10020) );
and4 gate2835( .a(N9779), .b(N9385), .c(N8298), .d(N8262), .O(N10021) );
and5 gate2836( .a(N367), .b(N9775), .c(N9385), .d(N8298), .e(N8262), .O(N10022) );
inv1 gate2837( .a(N9945), .O(N10023) );
inv1 gate2838( .a(N9946), .O(N10024) );
nand2 gate2839( .a(N9740), .b(N9893), .O(N10025) );
inv1 gate2840( .a(N9923), .O(N10026) );
inv1 gate2841( .a(N9924), .O(N10028) );
nand2 gate2842( .a(N8595), .b(N9897), .O(N10032) );
nand2 gate2843( .a(N8598), .b(N9899), .O(N10033) );
nand2 gate2844( .a(N8601), .b(N9901), .O(N10034) );
nand2 gate2845( .a(N8604), .b(N9903), .O(N10035) );
nand2 gate2846( .a(N4803), .b(N9906), .O(N10036) );
nand2 gate2847( .a(N4806), .b(N9908), .O(N10037) );
nand2 gate2848( .a(N8627), .b(N9910), .O(N10038) );
and2 gate2849( .a(N9809), .b(N8298), .O(N10039) );
and3 gate2850( .a(N9779), .b(N9385), .c(N8298), .O(N10040) );
and4 gate2851( .a(N367), .b(N9775), .c(N9385), .d(N8298), .O(N10041) );
and2 gate2852( .a(N9779), .b(N9385), .O(N10042) );
and3 gate2853( .a(N367), .b(N9775), .c(N9385), .O(N10043) );
nand2 gate2854( .a(N8727), .b(N9938), .O(N10050) );
inv1 gate2855( .a(N9817), .O(N10053) );
and2 gate2856( .a(N9817), .b(N9029), .O(N10054) );
and2 gate2857( .a(N9786), .b(N8394), .O(N10055) );
and3 gate2858( .a(N9820), .b(N9332), .c(N8394), .O(N10056) );
and2 gate2859( .a(N9791), .b(N8307), .O(N10057) );
and3 gate2860( .a(N9758), .b(N9344), .c(N8307), .O(N10058) );
and4 gate2861( .a(N367), .b(N9754), .c(N9344), .d(N8307), .O(N10059) );
and2 gate2862( .a(N9758), .b(N9344), .O(N10060) );
and3 gate2863( .a(N367), .b(N9754), .c(N9344), .O(N10061) );
nand2 gate2864( .a(N4997), .b(N9947), .O(N10062) );
nand2 gate2865( .a(N8811), .b(N9953), .O(N10067) );
nand2 gate2866( .a(N9955), .b(N9836), .O(N10070) );
nand2 gate2867( .a(N9956), .b(N9838), .O(N10073) );
nand2 gate2868( .a(N9068), .b(N9957), .O(N10076) );
nand2 gate2869( .a(N9074), .b(N9959), .O(N10077) );

  xor2  gate3822(.a(N9967), .b(N9089), .O(gate2870inter0));
  nand2 gate3823(.a(gate2870inter0), .b(s_44), .O(gate2870inter1));
  and2  gate3824(.a(N9967), .b(N9089), .O(gate2870inter2));
  inv1  gate3825(.a(s_44), .O(gate2870inter3));
  inv1  gate3826(.a(s_45), .O(gate2870inter4));
  nand2 gate3827(.a(gate2870inter4), .b(gate2870inter3), .O(gate2870inter5));
  nor2  gate3828(.a(gate2870inter5), .b(gate2870inter2), .O(gate2870inter6));
  inv1  gate3829(.a(N9089), .O(gate2870inter7));
  inv1  gate3830(.a(N9967), .O(gate2870inter8));
  nand2 gate3831(.a(gate2870inter8), .b(gate2870inter7), .O(gate2870inter9));
  nand2 gate3832(.a(s_45), .b(gate2870inter3), .O(gate2870inter10));
  nor2  gate3833(.a(gate2870inter10), .b(gate2870inter9), .O(gate2870inter11));
  nor2  gate3834(.a(gate2870inter11), .b(gate2870inter6), .O(gate2870inter12));
  nand2 gate3835(.a(gate2870inter12), .b(gate2870inter1), .O(N10082));
nand2 gate2871( .a(N9095), .b(N9969), .O(N10083) );
nand2 gate2872( .a(N4871), .b(N9971), .O(N10084) );
nand2 gate2873( .a(N6214), .b(N9973), .O(N10085) );
nand2 gate2874( .a(N6217), .b(N9975), .O(N10086) );
nand2 gate2875( .a(N5027), .b(N9995), .O(N10093) );
nand2 gate2876( .a(N6232), .b(N9997), .O(N10094) );
or5 gate2877( .a(N9238), .b(N9732), .c(N10013), .d(N10014), .e(N10015), .O(N10101) );
or5 gate2878( .a(N9339), .b(N9526), .c(N10016), .d(N10017), .e(N9734), .O(N10102) );
or5 gate2879( .a(N9339), .b(N9531), .c(N10018), .d(N10019), .e(N9735), .O(N10103) );
or5 gate2880( .a(N9242), .b(N9736), .c(N10020), .d(N10021), .e(N10022), .O(N10104) );
and2 gate2881( .a(N9925), .b(N9894), .O(N10105) );
and2 gate2882( .a(N9925), .b(N9895), .O(N10106) );
and2 gate2883( .a(N9925), .b(N9896), .O(N10107) );
and2 gate2884( .a(N9925), .b(N8253), .O(N10108) );

  xor2  gate3668(.a(N9898), .b(N10032), .O(gate2885inter0));
  nand2 gate3669(.a(gate2885inter0), .b(s_22), .O(gate2885inter1));
  and2  gate3670(.a(N9898), .b(N10032), .O(gate2885inter2));
  inv1  gate3671(.a(s_22), .O(gate2885inter3));
  inv1  gate3672(.a(s_23), .O(gate2885inter4));
  nand2 gate3673(.a(gate2885inter4), .b(gate2885inter3), .O(gate2885inter5));
  nor2  gate3674(.a(gate2885inter5), .b(gate2885inter2), .O(gate2885inter6));
  inv1  gate3675(.a(N10032), .O(gate2885inter7));
  inv1  gate3676(.a(N9898), .O(gate2885inter8));
  nand2 gate3677(.a(gate2885inter8), .b(gate2885inter7), .O(gate2885inter9));
  nand2 gate3678(.a(s_23), .b(gate2885inter3), .O(gate2885inter10));
  nor2  gate3679(.a(gate2885inter10), .b(gate2885inter9), .O(gate2885inter11));
  nor2  gate3680(.a(gate2885inter11), .b(gate2885inter6), .O(gate2885inter12));
  nand2 gate3681(.a(gate2885inter12), .b(gate2885inter1), .O(N10109));
nand2 gate2886( .a(N10033), .b(N9900), .O(N10110) );
nand2 gate2887( .a(N10034), .b(N9902), .O(N10111) );
nand2 gate2888( .a(N10035), .b(N9904), .O(N10112) );
nand2 gate2889( .a(N10036), .b(N9907), .O(N10113) );
nand2 gate2890( .a(N10037), .b(N9909), .O(N10114) );

  xor2  gate4522(.a(N9911), .b(N10038), .O(gate2891inter0));
  nand2 gate4523(.a(gate2891inter0), .b(s_144), .O(gate2891inter1));
  and2  gate4524(.a(N9911), .b(N10038), .O(gate2891inter2));
  inv1  gate4525(.a(s_144), .O(gate2891inter3));
  inv1  gate4526(.a(s_145), .O(gate2891inter4));
  nand2 gate4527(.a(gate2891inter4), .b(gate2891inter3), .O(gate2891inter5));
  nor2  gate4528(.a(gate2891inter5), .b(gate2891inter2), .O(gate2891inter6));
  inv1  gate4529(.a(N10038), .O(gate2891inter7));
  inv1  gate4530(.a(N9911), .O(gate2891inter8));
  nand2 gate4531(.a(gate2891inter8), .b(gate2891inter7), .O(gate2891inter9));
  nand2 gate4532(.a(s_145), .b(gate2891inter3), .O(gate2891inter10));
  nor2  gate4533(.a(gate2891inter10), .b(gate2891inter9), .O(gate2891inter11));
  nor2  gate4534(.a(gate2891inter11), .b(gate2891inter6), .O(gate2891inter12));
  nand2 gate4535(.a(gate2891inter12), .b(gate2891inter1), .O(N10115));
or4 gate2892( .a(N9265), .b(N10039), .c(N10040), .d(N10041), .O(N10116) );
or3 gate2893( .a(N9809), .b(N10042), .c(N10043), .O(N10119) );
inv1 gate2894( .a(N9925), .O(N10124) );
and2 gate2895( .a(N9768), .b(N9925), .O(N10130) );
inv1 gate2896( .a(N9932), .O(N10131) );
inv1 gate2897( .a(N9935), .O(N10132) );
and2 gate2898( .a(N9932), .b(N8920), .O(N10133) );
nand2 gate2899( .a(N10050), .b(N9939), .O(N10134) );
inv1 gate2900( .a(N9983), .O(N10135) );
nand2 gate2901( .a(N9983), .b(N9324), .O(N10136) );
inv1 gate2902( .a(N9986), .O(N10137) );
nand2 gate2903( .a(N9986), .b(N9784), .O(N10138) );
and2 gate2904( .a(N9785), .b(N10053), .O(N10139) );
or4 gate2905( .a(N8943), .b(N10055), .c(N10056), .d(N9790), .O(N10140) );
or4 gate2906( .a(N9268), .b(N10057), .c(N10058), .d(N10059), .O(N10141) );
or3 gate2907( .a(N9791), .b(N10060), .c(N10061), .O(N10148) );
nand2 gate2908( .a(N10062), .b(N9948), .O(N10155) );
inv1 gate2909( .a(N9989), .O(N10156) );
nand2 gate2910( .a(N9989), .b(N9805), .O(N10157) );
inv1 gate2911( .a(N9992), .O(N10158) );
nand2 gate2912( .a(N9992), .b(N9806), .O(N10159) );
inv1 gate2913( .a(N9949), .O(N10160) );
nand2 gate2914( .a(N10067), .b(N9954), .O(N10161) );
inv1 gate2915( .a(N10007), .O(N10162) );
nand2 gate2916( .a(N10007), .b(N9825), .O(N10163) );
inv1 gate2917( .a(N10010), .O(N10164) );
nand2 gate2918( .a(N10010), .b(N9826), .O(N10165) );
nand2 gate2919( .a(N10076), .b(N9958), .O(N10170) );

  xor2  gate3724(.a(N9960), .b(N10077), .O(gate2920inter0));
  nand2 gate3725(.a(gate2920inter0), .b(s_30), .O(gate2920inter1));
  and2  gate3726(.a(N9960), .b(N10077), .O(gate2920inter2));
  inv1  gate3727(.a(s_30), .O(gate2920inter3));
  inv1  gate3728(.a(s_31), .O(gate2920inter4));
  nand2 gate3729(.a(gate2920inter4), .b(gate2920inter3), .O(gate2920inter5));
  nor2  gate3730(.a(gate2920inter5), .b(gate2920inter2), .O(gate2920inter6));
  inv1  gate3731(.a(N10077), .O(gate2920inter7));
  inv1  gate3732(.a(N9960), .O(gate2920inter8));
  nand2 gate3733(.a(gate2920inter8), .b(gate2920inter7), .O(gate2920inter9));
  nand2 gate3734(.a(s_31), .b(gate2920inter3), .O(gate2920inter10));
  nor2  gate3735(.a(gate2920inter10), .b(gate2920inter9), .O(gate2920inter11));
  nor2  gate3736(.a(gate2920inter11), .b(gate2920inter6), .O(gate2920inter12));
  nand2 gate3737(.a(gate2920inter12), .b(gate2920inter1), .O(N10173));
inv1 gate2921( .a(N9961), .O(N10176) );
nand2 gate2922( .a(N9961), .b(N9082), .O(N10177) );
inv1 gate2923( .a(N9964), .O(N10178) );
nand2 gate2924( .a(N9964), .b(N9086), .O(N10179) );
nand2 gate2925( .a(N10082), .b(N9968), .O(N10180) );
nand2 gate2926( .a(N10083), .b(N9970), .O(N10183) );
nand2 gate2927( .a(N9972), .b(N10084), .O(N10186) );
nand2 gate2928( .a(N9974), .b(N10085), .O(N10189) );
nand2 gate2929( .a(N9976), .b(N10086), .O(N10192) );
inv1 gate2930( .a(N9979), .O(N10195) );
nand2 gate2931( .a(N9979), .b(N9982), .O(N10196) );

  xor2  gate4886(.a(N10093), .b(N9996), .O(gate2932inter0));
  nand2 gate4887(.a(gate2932inter0), .b(s_196), .O(gate2932inter1));
  and2  gate4888(.a(N10093), .b(N9996), .O(gate2932inter2));
  inv1  gate4889(.a(s_196), .O(gate2932inter3));
  inv1  gate4890(.a(s_197), .O(gate2932inter4));
  nand2 gate4891(.a(gate2932inter4), .b(gate2932inter3), .O(gate2932inter5));
  nor2  gate4892(.a(gate2932inter5), .b(gate2932inter2), .O(gate2932inter6));
  inv1  gate4893(.a(N9996), .O(gate2932inter7));
  inv1  gate4894(.a(N10093), .O(gate2932inter8));
  nand2 gate4895(.a(gate2932inter8), .b(gate2932inter7), .O(gate2932inter9));
  nand2 gate4896(.a(s_197), .b(gate2932inter3), .O(gate2932inter10));
  nor2  gate4897(.a(gate2932inter10), .b(gate2932inter9), .O(gate2932inter11));
  nor2  gate4898(.a(gate2932inter11), .b(gate2932inter6), .O(gate2932inter12));
  nand2 gate4899(.a(gate2932inter12), .b(gate2932inter1), .O(N10197));
nand2 gate2933( .a(N9998), .b(N10094), .O(N10200) );
inv1 gate2934( .a(N9999), .O(N10203) );
nand2 gate2935( .a(N9999), .b(N10002), .O(N10204) );
inv1 gate2936( .a(N10003), .O(N10205) );
nand2 gate2937( .a(N10003), .b(N10006), .O(N10206) );
nand2 gate2938( .a(N10070), .b(N4308), .O(N10212) );
nand2 gate2939( .a(N10073), .b(N4313), .O(N10213) );
and2 gate2940( .a(N9774), .b(N10131), .O(N10230) );
nand2 gate2941( .a(N8730), .b(N10135), .O(N10231) );
nand2 gate2942( .a(N9478), .b(N10137), .O(N10232) );
or2 gate2943( .a(N10139), .b(N10054), .O(N10233) );
nand2 gate2944( .a(N7100), .b(N10140), .O(N10234) );
nand2 gate2945( .a(N9485), .b(N10156), .O(N10237) );

  xor2  gate4256(.a(N10158), .b(N9488), .O(gate2946inter0));
  nand2 gate4257(.a(gate2946inter0), .b(s_106), .O(gate2946inter1));
  and2  gate4258(.a(N10158), .b(N9488), .O(gate2946inter2));
  inv1  gate4259(.a(s_106), .O(gate2946inter3));
  inv1  gate4260(.a(s_107), .O(gate2946inter4));
  nand2 gate4261(.a(gate2946inter4), .b(gate2946inter3), .O(gate2946inter5));
  nor2  gate4262(.a(gate2946inter5), .b(gate2946inter2), .O(gate2946inter6));
  inv1  gate4263(.a(N9488), .O(gate2946inter7));
  inv1  gate4264(.a(N10158), .O(gate2946inter8));
  nand2 gate4265(.a(gate2946inter8), .b(gate2946inter7), .O(gate2946inter9));
  nand2 gate4266(.a(s_107), .b(gate2946inter3), .O(gate2946inter10));
  nor2  gate4267(.a(gate2946inter10), .b(gate2946inter9), .O(gate2946inter11));
  nor2  gate4268(.a(gate2946inter11), .b(gate2946inter6), .O(gate2946inter12));
  nand2 gate4269(.a(gate2946inter12), .b(gate2946inter1), .O(N10238));

  xor2  gate4466(.a(N10162), .b(N9517), .O(gate2947inter0));
  nand2 gate4467(.a(gate2947inter0), .b(s_136), .O(gate2947inter1));
  and2  gate4468(.a(N10162), .b(N9517), .O(gate2947inter2));
  inv1  gate4469(.a(s_136), .O(gate2947inter3));
  inv1  gate4470(.a(s_137), .O(gate2947inter4));
  nand2 gate4471(.a(gate2947inter4), .b(gate2947inter3), .O(gate2947inter5));
  nor2  gate4472(.a(gate2947inter5), .b(gate2947inter2), .O(gate2947inter6));
  inv1  gate4473(.a(N9517), .O(gate2947inter7));
  inv1  gate4474(.a(N10162), .O(gate2947inter8));
  nand2 gate4475(.a(gate2947inter8), .b(gate2947inter7), .O(gate2947inter9));
  nand2 gate4476(.a(s_137), .b(gate2947inter3), .O(gate2947inter10));
  nor2  gate4477(.a(gate2947inter10), .b(gate2947inter9), .O(gate2947inter11));
  nor2  gate4478(.a(gate2947inter11), .b(gate2947inter6), .O(gate2947inter12));
  nand2 gate4479(.a(gate2947inter12), .b(gate2947inter1), .O(N10239));
nand2 gate2948( .a(N9520), .b(N10164), .O(N10240) );
inv1 gate2949( .a(N10070), .O(N10241) );
inv1 gate2950( .a(N10073), .O(N10242) );
nand2 gate2951( .a(N8146), .b(N10176), .O(N10247) );
nand2 gate2952( .a(N8156), .b(N10178), .O(N10248) );
nand2 gate2953( .a(N9692), .b(N10195), .O(N10259) );
nand2 gate2954( .a(N9717), .b(N10203), .O(N10264) );
nand2 gate2955( .a(N9723), .b(N10205), .O(N10265) );
and2 gate2956( .a(N10026), .b(N10124), .O(N10266) );
and2 gate2957( .a(N10028), .b(N10124), .O(N10267) );
and2 gate2958( .a(N9742), .b(N10124), .O(N10268) );
and2 gate2959( .a(N6923), .b(N10124), .O(N10269) );
nand2 gate2960( .a(N6762), .b(N10116), .O(N10270) );
nand2 gate2961( .a(N3061), .b(N10241), .O(N10271) );
nand2 gate2962( .a(N3064), .b(N10242), .O(N10272) );
buf1 gate2963( .a(N10116), .O(N10273) );
and5 gate2964( .a(N10141), .b(N5728), .c(N5707), .d(N5718), .e(N5697), .O(N10278) );
and4 gate2965( .a(N10141), .b(N5728), .c(N5707), .d(N5718), .O(N10279) );
and3 gate2966( .a(N10141), .b(N5728), .c(N5718), .O(N10280) );
and2 gate2967( .a(N10141), .b(N5728), .O(N10281) );
and2 gate2968( .a(N6784), .b(N10141), .O(N10282) );
inv1 gate2969( .a(N10119), .O(N10283) );
and5 gate2970( .a(N10148), .b(N5936), .c(N5915), .d(N5926), .e(N5905), .O(N10287) );
and4 gate2971( .a(N10148), .b(N5936), .c(N5915), .d(N5926), .O(N10288) );
and3 gate2972( .a(N10148), .b(N5936), .c(N5926), .O(N10289) );
and2 gate2973( .a(N10148), .b(N5936), .O(N10290) );
and2 gate2974( .a(N6881), .b(N10148), .O(N10291) );
and2 gate2975( .a(N8898), .b(N10124), .O(N10292) );

  xor2  gate3794(.a(N10136), .b(N10231), .O(gate2976inter0));
  nand2 gate3795(.a(gate2976inter0), .b(s_40), .O(gate2976inter1));
  and2  gate3796(.a(N10136), .b(N10231), .O(gate2976inter2));
  inv1  gate3797(.a(s_40), .O(gate2976inter3));
  inv1  gate3798(.a(s_41), .O(gate2976inter4));
  nand2 gate3799(.a(gate2976inter4), .b(gate2976inter3), .O(gate2976inter5));
  nor2  gate3800(.a(gate2976inter5), .b(gate2976inter2), .O(gate2976inter6));
  inv1  gate3801(.a(N10231), .O(gate2976inter7));
  inv1  gate3802(.a(N10136), .O(gate2976inter8));
  nand2 gate3803(.a(gate2976inter8), .b(gate2976inter7), .O(gate2976inter9));
  nand2 gate3804(.a(s_41), .b(gate2976inter3), .O(gate2976inter10));
  nor2  gate3805(.a(gate2976inter10), .b(gate2976inter9), .O(gate2976inter11));
  nor2  gate3806(.a(gate2976inter11), .b(gate2976inter6), .O(gate2976inter12));
  nand2 gate3807(.a(gate2976inter12), .b(gate2976inter1), .O(N10293));
nand2 gate2977( .a(N10232), .b(N10138), .O(N10294) );
nand2 gate2978( .a(N8412), .b(N10233), .O(N10295) );
and2 gate2979( .a(N8959), .b(N10234), .O(N10296) );
nand2 gate2980( .a(N10237), .b(N10157), .O(N10299) );
nand2 gate2981( .a(N10238), .b(N10159), .O(N10300) );
or2 gate2982( .a(N10230), .b(N10133), .O(N10301) );
nand2 gate2983( .a(N10239), .b(N10163), .O(N10306) );
nand2 gate2984( .a(N10240), .b(N10165), .O(N10307) );
buf1 gate2985( .a(N10148), .O(N10308) );
buf1 gate2986( .a(N10141), .O(N10311) );
inv1 gate2987( .a(N10170), .O(N10314) );
nand2 gate2988( .a(N10170), .b(N9071), .O(N10315) );
inv1 gate2989( .a(N10173), .O(N10316) );
nand2 gate2990( .a(N10173), .b(N9077), .O(N10317) );
nand2 gate2991( .a(N10247), .b(N10177), .O(N10318) );
nand2 gate2992( .a(N10248), .b(N10179), .O(N10321) );
inv1 gate2993( .a(N10180), .O(N10324) );
nand2 gate2994( .a(N10180), .b(N9092), .O(N10325) );
inv1 gate2995( .a(N10183), .O(N10326) );
nand2 gate2996( .a(N10183), .b(N9098), .O(N10327) );
inv1 gate2997( .a(N10186), .O(N10328) );
nand2 gate2998( .a(N10186), .b(N9674), .O(N10329) );
inv1 gate2999( .a(N10189), .O(N10330) );
nand2 gate3000( .a(N10189), .b(N9678), .O(N10331) );
inv1 gate3001( .a(N10192), .O(N10332) );
nand2 gate3002( .a(N10192), .b(N9977), .O(N10333) );

  xor2  gate3780(.a(N10196), .b(N10259), .O(gate3003inter0));
  nand2 gate3781(.a(gate3003inter0), .b(s_38), .O(gate3003inter1));
  and2  gate3782(.a(N10196), .b(N10259), .O(gate3003inter2));
  inv1  gate3783(.a(s_38), .O(gate3003inter3));
  inv1  gate3784(.a(s_39), .O(gate3003inter4));
  nand2 gate3785(.a(gate3003inter4), .b(gate3003inter3), .O(gate3003inter5));
  nor2  gate3786(.a(gate3003inter5), .b(gate3003inter2), .O(gate3003inter6));
  inv1  gate3787(.a(N10259), .O(gate3003inter7));
  inv1  gate3788(.a(N10196), .O(gate3003inter8));
  nand2 gate3789(.a(gate3003inter8), .b(gate3003inter7), .O(gate3003inter9));
  nand2 gate3790(.a(s_39), .b(gate3003inter3), .O(gate3003inter10));
  nor2  gate3791(.a(gate3003inter10), .b(gate3003inter9), .O(gate3003inter11));
  nor2  gate3792(.a(gate3003inter11), .b(gate3003inter6), .O(gate3003inter12));
  nand2 gate3793(.a(gate3003inter12), .b(gate3003inter1), .O(N10334));
inv1 gate3004( .a(N10197), .O(N10337) );
nand2 gate3005( .a(N10197), .b(N9710), .O(N10338) );
inv1 gate3006( .a(N10200), .O(N10339) );
nand2 gate3007( .a(N10200), .b(N9714), .O(N10340) );
nand2 gate3008( .a(N10264), .b(N10204), .O(N10341) );
nand2 gate3009( .a(N10265), .b(N10206), .O(N10344) );
or2 gate3010( .a(N10266), .b(N10105), .O(N10350) );
or2 gate3011( .a(N10267), .b(N10106), .O(N10351) );
or2 gate3012( .a(N10268), .b(N10107), .O(N10352) );
or2 gate3013( .a(N10269), .b(N10108), .O(N10353) );
and2 gate3014( .a(N8857), .b(N10270), .O(N10354) );
nand2 gate3015( .a(N10271), .b(N10212), .O(N10357) );
nand2 gate3016( .a(N10272), .b(N10213), .O(N10360) );
or2 gate3017( .a(N7620), .b(N10282), .O(N10367) );
or2 gate3018( .a(N7671), .b(N10291), .O(N10375) );
or2 gate3019( .a(N10292), .b(N10130), .O(N10381) );
and4 gate3020( .a(N10114), .b(N10134), .c(N10293), .d(N10294), .O(N10388) );
and2 gate3021( .a(N9582), .b(N10295), .O(N10391) );
and4 gate3022( .a(N10113), .b(N10115), .c(N10299), .d(N10300), .O(N10399) );
and4 gate3023( .a(N10155), .b(N10161), .c(N10306), .d(N10307), .O(N10402) );
or5 gate3024( .a(N3229), .b(N6888), .c(N6889), .d(N6890), .e(N10287), .O(N10406) );
or4 gate3025( .a(N3232), .b(N6891), .c(N6892), .d(N10288), .O(N10409) );
or3 gate3026( .a(N3236), .b(N6893), .c(N10289), .O(N10412) );
or2 gate3027( .a(N3241), .b(N10290), .O(N10415) );
or5 gate3028( .a(N3137), .b(N6791), .c(N6792), .d(N6793), .e(N10278), .O(N10419) );
or4 gate3029( .a(N3140), .b(N6794), .c(N6795), .d(N10279), .O(N10422) );
or3 gate3030( .a(N3144), .b(N6796), .c(N10280), .O(N10425) );
or2 gate3031( .a(N3149), .b(N10281), .O(N10428) );
nand2 gate3032( .a(N8117), .b(N10314), .O(N10431) );
nand2 gate3033( .a(N8134), .b(N10316), .O(N10432) );
nand2 gate3034( .a(N8169), .b(N10324), .O(N10437) );
nand2 gate3035( .a(N8186), .b(N10326), .O(N10438) );
nand2 gate3036( .a(N9117), .b(N10328), .O(N10439) );
nand2 gate3037( .a(N9127), .b(N10330), .O(N10440) );

  xor2  gate4858(.a(N10332), .b(N9682), .O(gate3038inter0));
  nand2 gate4859(.a(gate3038inter0), .b(s_192), .O(gate3038inter1));
  and2  gate4860(.a(N10332), .b(N9682), .O(gate3038inter2));
  inv1  gate4861(.a(s_192), .O(gate3038inter3));
  inv1  gate4862(.a(s_193), .O(gate3038inter4));
  nand2 gate4863(.a(gate3038inter4), .b(gate3038inter3), .O(gate3038inter5));
  nor2  gate4864(.a(gate3038inter5), .b(gate3038inter2), .O(gate3038inter6));
  inv1  gate4865(.a(N9682), .O(gate3038inter7));
  inv1  gate4866(.a(N10332), .O(gate3038inter8));
  nand2 gate4867(.a(gate3038inter8), .b(gate3038inter7), .O(gate3038inter9));
  nand2 gate4868(.a(s_193), .b(gate3038inter3), .O(gate3038inter10));
  nor2  gate4869(.a(gate3038inter10), .b(gate3038inter9), .O(gate3038inter11));
  nor2  gate4870(.a(gate3038inter11), .b(gate3038inter6), .O(gate3038inter12));
  nand2 gate4871(.a(gate3038inter12), .b(gate3038inter1), .O(N10441));
nand2 gate3039( .a(N9183), .b(N10337), .O(N10444) );
nand2 gate3040( .a(N9193), .b(N10339), .O(N10445) );
inv1 gate3041( .a(N10296), .O(N10450) );
and2 gate3042( .a(N10296), .b(N4193), .O(N10451) );
inv1 gate3043( .a(N10308), .O(N10455) );
nand2 gate3044( .a(N10308), .b(N8242), .O(N10456) );
inv1 gate3045( .a(N10311), .O(N10465) );

  xor2  gate4942(.a(N8247), .b(N10311), .O(gate3046inter0));
  nand2 gate4943(.a(gate3046inter0), .b(s_204), .O(gate3046inter1));
  and2  gate4944(.a(N8247), .b(N10311), .O(gate3046inter2));
  inv1  gate4945(.a(s_204), .O(gate3046inter3));
  inv1  gate4946(.a(s_205), .O(gate3046inter4));
  nand2 gate4947(.a(gate3046inter4), .b(gate3046inter3), .O(gate3046inter5));
  nor2  gate4948(.a(gate3046inter5), .b(gate3046inter2), .O(gate3046inter6));
  inv1  gate4949(.a(N10311), .O(gate3046inter7));
  inv1  gate4950(.a(N8247), .O(gate3046inter8));
  nand2 gate4951(.a(gate3046inter8), .b(gate3046inter7), .O(gate3046inter9));
  nand2 gate4952(.a(s_205), .b(gate3046inter3), .O(gate3046inter10));
  nor2  gate4953(.a(gate3046inter10), .b(gate3046inter9), .O(gate3046inter11));
  nor2  gate4954(.a(gate3046inter11), .b(gate3046inter6), .O(gate3046inter12));
  nand2 gate4955(.a(gate3046inter12), .b(gate3046inter1), .O(N10466));
inv1 gate3047( .a(N10273), .O(N10479) );
inv1 gate3048( .a(N10301), .O(N10497) );
nand2 gate3049( .a(N10431), .b(N10315), .O(N10509) );

  xor2  gate4592(.a(N10317), .b(N10432), .O(gate3050inter0));
  nand2 gate4593(.a(gate3050inter0), .b(s_154), .O(gate3050inter1));
  and2  gate4594(.a(N10317), .b(N10432), .O(gate3050inter2));
  inv1  gate4595(.a(s_154), .O(gate3050inter3));
  inv1  gate4596(.a(s_155), .O(gate3050inter4));
  nand2 gate4597(.a(gate3050inter4), .b(gate3050inter3), .O(gate3050inter5));
  nor2  gate4598(.a(gate3050inter5), .b(gate3050inter2), .O(gate3050inter6));
  inv1  gate4599(.a(N10432), .O(gate3050inter7));
  inv1  gate4600(.a(N10317), .O(gate3050inter8));
  nand2 gate4601(.a(gate3050inter8), .b(gate3050inter7), .O(gate3050inter9));
  nand2 gate4602(.a(s_155), .b(gate3050inter3), .O(gate3050inter10));
  nor2  gate4603(.a(gate3050inter10), .b(gate3050inter9), .O(gate3050inter11));
  nor2  gate4604(.a(gate3050inter11), .b(gate3050inter6), .O(gate3050inter12));
  nand2 gate4605(.a(gate3050inter12), .b(gate3050inter1), .O(N10512));
inv1 gate3051( .a(N10318), .O(N10515) );
nand2 gate3052( .a(N10318), .b(N8632), .O(N10516) );
inv1 gate3053( .a(N10321), .O(N10517) );

  xor2  gate4340(.a(N8637), .b(N10321), .O(gate3054inter0));
  nand2 gate4341(.a(gate3054inter0), .b(s_118), .O(gate3054inter1));
  and2  gate4342(.a(N8637), .b(N10321), .O(gate3054inter2));
  inv1  gate4343(.a(s_118), .O(gate3054inter3));
  inv1  gate4344(.a(s_119), .O(gate3054inter4));
  nand2 gate4345(.a(gate3054inter4), .b(gate3054inter3), .O(gate3054inter5));
  nor2  gate4346(.a(gate3054inter5), .b(gate3054inter2), .O(gate3054inter6));
  inv1  gate4347(.a(N10321), .O(gate3054inter7));
  inv1  gate4348(.a(N8637), .O(gate3054inter8));
  nand2 gate4349(.a(gate3054inter8), .b(gate3054inter7), .O(gate3054inter9));
  nand2 gate4350(.a(s_119), .b(gate3054inter3), .O(gate3054inter10));
  nor2  gate4351(.a(gate3054inter10), .b(gate3054inter9), .O(gate3054inter11));
  nor2  gate4352(.a(gate3054inter11), .b(gate3054inter6), .O(gate3054inter12));
  nand2 gate4353(.a(gate3054inter12), .b(gate3054inter1), .O(N10518));
nand2 gate3055( .a(N10437), .b(N10325), .O(N10519) );
nand2 gate3056( .a(N10438), .b(N10327), .O(N10522) );
nand2 gate3057( .a(N10439), .b(N10329), .O(N10525) );
nand2 gate3058( .a(N10440), .b(N10331), .O(N10528) );
nand2 gate3059( .a(N10441), .b(N10333), .O(N10531) );
inv1 gate3060( .a(N10334), .O(N10534) );
nand2 gate3061( .a(N10334), .b(N9695), .O(N10535) );
nand2 gate3062( .a(N10444), .b(N10338), .O(N10536) );
nand2 gate3063( .a(N10445), .b(N10340), .O(N10539) );
inv1 gate3064( .a(N10341), .O(N10542) );
nand2 gate3065( .a(N10341), .b(N9720), .O(N10543) );
inv1 gate3066( .a(N10344), .O(N10544) );
nand2 gate3067( .a(N10344), .b(N9726), .O(N10545) );
and2 gate3068( .a(N5631), .b(N10450), .O(N10546) );
inv1 gate3069( .a(N10391), .O(N10547) );
and2 gate3070( .a(N10391), .b(N8950), .O(N10548) );
and2 gate3071( .a(N5165), .b(N10367), .O(N10549) );
inv1 gate3072( .a(N10354), .O(N10550) );
and2 gate3073( .a(N10354), .b(N3126), .O(N10551) );
nand2 gate3074( .a(N7411), .b(N10455), .O(N10552) );
and2 gate3075( .a(N10375), .b(N9539), .O(N10553) );
and2 gate3076( .a(N10375), .b(N9540), .O(N10554) );
and2 gate3077( .a(N10375), .b(N9541), .O(N10555) );
and2 gate3078( .a(N10375), .b(N6761), .O(N10556) );
inv1 gate3079( .a(N10406), .O(N10557) );
nand2 gate3080( .a(N10406), .b(N8243), .O(N10558) );
inv1 gate3081( .a(N10409), .O(N10559) );

  xor2  gate3626(.a(N8244), .b(N10409), .O(gate3082inter0));
  nand2 gate3627(.a(gate3082inter0), .b(s_16), .O(gate3082inter1));
  and2  gate3628(.a(N8244), .b(N10409), .O(gate3082inter2));
  inv1  gate3629(.a(s_16), .O(gate3082inter3));
  inv1  gate3630(.a(s_17), .O(gate3082inter4));
  nand2 gate3631(.a(gate3082inter4), .b(gate3082inter3), .O(gate3082inter5));
  nor2  gate3632(.a(gate3082inter5), .b(gate3082inter2), .O(gate3082inter6));
  inv1  gate3633(.a(N10409), .O(gate3082inter7));
  inv1  gate3634(.a(N8244), .O(gate3082inter8));
  nand2 gate3635(.a(gate3082inter8), .b(gate3082inter7), .O(gate3082inter9));
  nand2 gate3636(.a(s_17), .b(gate3082inter3), .O(gate3082inter10));
  nor2  gate3637(.a(gate3082inter10), .b(gate3082inter9), .O(gate3082inter11));
  nor2  gate3638(.a(gate3082inter11), .b(gate3082inter6), .O(gate3082inter12));
  nand2 gate3639(.a(gate3082inter12), .b(gate3082inter1), .O(N10560));
inv1 gate3083( .a(N10412), .O(N10561) );

  xor2  gate5110(.a(N8245), .b(N10412), .O(gate3084inter0));
  nand2 gate5111(.a(gate3084inter0), .b(s_228), .O(gate3084inter1));
  and2  gate5112(.a(N8245), .b(N10412), .O(gate3084inter2));
  inv1  gate5113(.a(s_228), .O(gate3084inter3));
  inv1  gate5114(.a(s_229), .O(gate3084inter4));
  nand2 gate5115(.a(gate3084inter4), .b(gate3084inter3), .O(gate3084inter5));
  nor2  gate5116(.a(gate3084inter5), .b(gate3084inter2), .O(gate3084inter6));
  inv1  gate5117(.a(N10412), .O(gate3084inter7));
  inv1  gate5118(.a(N8245), .O(gate3084inter8));
  nand2 gate5119(.a(gate3084inter8), .b(gate3084inter7), .O(gate3084inter9));
  nand2 gate5120(.a(s_229), .b(gate3084inter3), .O(gate3084inter10));
  nor2  gate5121(.a(gate3084inter10), .b(gate3084inter9), .O(gate3084inter11));
  nor2  gate5122(.a(gate3084inter11), .b(gate3084inter6), .O(gate3084inter12));
  nand2 gate5123(.a(gate3084inter12), .b(gate3084inter1), .O(N10562));
inv1 gate3085( .a(N10415), .O(N10563) );
nand2 gate3086( .a(N10415), .b(N8246), .O(N10564) );
nand2 gate3087( .a(N7426), .b(N10465), .O(N10565) );
inv1 gate3088( .a(N10419), .O(N10566) );
nand2 gate3089( .a(N10419), .b(N8248), .O(N10567) );
inv1 gate3090( .a(N10422), .O(N10568) );
nand2 gate3091( .a(N10422), .b(N8249), .O(N10569) );
inv1 gate3092( .a(N10425), .O(N10570) );
nand2 gate3093( .a(N10425), .b(N8250), .O(N10571) );
inv1 gate3094( .a(N10428), .O(N10572) );
nand2 gate3095( .a(N10428), .b(N8251), .O(N10573) );
inv1 gate3096( .a(N10399), .O(N10574) );
inv1 gate3097( .a(N10402), .O(N10575) );
inv1 gate3098( .a(N10388), .O(N10576) );
and3 gate3099( .a(N10399), .b(N10402), .c(N10388), .O(N10577) );
and3 gate3100( .a(N10360), .b(N9543), .c(N10273), .O(N10581) );
and3 gate3101( .a(N10357), .b(N9905), .c(N10273), .O(N10582) );
inv1 gate3102( .a(N10367), .O(N10583) );
and2 gate3103( .a(N10367), .b(N5735), .O(N10587) );
and2 gate3104( .a(N10367), .b(N3135), .O(N10588) );
inv1 gate3105( .a(N10375), .O(N10589) );
and5 gate3106( .a(N10381), .b(N7180), .c(N7159), .d(N7170), .e(N7149), .O(N10594) );
and4 gate3107( .a(N10381), .b(N7180), .c(N7159), .d(N7170), .O(N10595) );
and3 gate3108( .a(N10381), .b(N7180), .c(N7170), .O(N10596) );
and2 gate3109( .a(N10381), .b(N7180), .O(N10597) );
and2 gate3110( .a(N8444), .b(N10381), .O(N10598) );
buf1 gate3111( .a(N10381), .O(N10602) );
nand2 gate3112( .a(N7479), .b(N10515), .O(N10609) );
nand2 gate3113( .a(N7491), .b(N10517), .O(N10610) );
nand2 gate3114( .a(N9149), .b(N10534), .O(N10621) );
nand2 gate3115( .a(N9206), .b(N10542), .O(N10626) );
nand2 gate3116( .a(N9223), .b(N10544), .O(N10627) );
or2 gate3117( .a(N10546), .b(N10451), .O(N10628) );
and2 gate3118( .a(N9733), .b(N10547), .O(N10629) );
and2 gate3119( .a(N5166), .b(N10550), .O(N10631) );

  xor2  gate5194(.a(N10456), .b(N10552), .O(gate3120inter0));
  nand2 gate5195(.a(gate3120inter0), .b(s_240), .O(gate3120inter1));
  and2  gate5196(.a(N10456), .b(N10552), .O(gate3120inter2));
  inv1  gate5197(.a(s_240), .O(gate3120inter3));
  inv1  gate5198(.a(s_241), .O(gate3120inter4));
  nand2 gate5199(.a(gate3120inter4), .b(gate3120inter3), .O(gate3120inter5));
  nor2  gate5200(.a(gate3120inter5), .b(gate3120inter2), .O(gate3120inter6));
  inv1  gate5201(.a(N10552), .O(gate3120inter7));
  inv1  gate5202(.a(N10456), .O(gate3120inter8));
  nand2 gate5203(.a(gate3120inter8), .b(gate3120inter7), .O(gate3120inter9));
  nand2 gate5204(.a(s_241), .b(gate3120inter3), .O(gate3120inter10));
  nor2  gate5205(.a(gate3120inter10), .b(gate3120inter9), .O(gate3120inter11));
  nor2  gate5206(.a(gate3120inter11), .b(gate3120inter6), .O(gate3120inter12));
  nand2 gate5207(.a(gate3120inter12), .b(gate3120inter1), .O(N10632));
nand2 gate3121( .a(N7414), .b(N10557), .O(N10637) );

  xor2  gate4970(.a(N10559), .b(N7417), .O(gate3122inter0));
  nand2 gate4971(.a(gate3122inter0), .b(s_208), .O(gate3122inter1));
  and2  gate4972(.a(N10559), .b(N7417), .O(gate3122inter2));
  inv1  gate4973(.a(s_208), .O(gate3122inter3));
  inv1  gate4974(.a(s_209), .O(gate3122inter4));
  nand2 gate4975(.a(gate3122inter4), .b(gate3122inter3), .O(gate3122inter5));
  nor2  gate4976(.a(gate3122inter5), .b(gate3122inter2), .O(gate3122inter6));
  inv1  gate4977(.a(N7417), .O(gate3122inter7));
  inv1  gate4978(.a(N10559), .O(gate3122inter8));
  nand2 gate4979(.a(gate3122inter8), .b(gate3122inter7), .O(gate3122inter9));
  nand2 gate4980(.a(s_209), .b(gate3122inter3), .O(gate3122inter10));
  nor2  gate4981(.a(gate3122inter10), .b(gate3122inter9), .O(gate3122inter11));
  nor2  gate4982(.a(gate3122inter11), .b(gate3122inter6), .O(gate3122inter12));
  nand2 gate4983(.a(gate3122inter12), .b(gate3122inter1), .O(N10638));
nand2 gate3123( .a(N7420), .b(N10561), .O(N10639) );
nand2 gate3124( .a(N7423), .b(N10563), .O(N10640) );
nand2 gate3125( .a(N10565), .b(N10466), .O(N10641) );
nand2 gate3126( .a(N7429), .b(N10566), .O(N10642) );
nand2 gate3127( .a(N7432), .b(N10568), .O(N10643) );
nand2 gate3128( .a(N7435), .b(N10570), .O(N10644) );
nand2 gate3129( .a(N7438), .b(N10572), .O(N10645) );
and3 gate3130( .a(N886), .b(N887), .c(N10577), .O(N10647) );
and3 gate3131( .a(N10360), .b(N8857), .c(N10479), .O(N10648) );
and3 gate3132( .a(N10357), .b(N7609), .c(N10479), .O(N10649) );
or2 gate3133( .a(N8966), .b(N10598), .O(N10652) );
or5 gate3134( .a(N4675), .b(N8451), .c(N8452), .d(N8453), .e(N10594), .O(N10659) );
or4 gate3135( .a(N4678), .b(N8454), .c(N8455), .d(N10595), .O(N10662) );
or3 gate3136( .a(N4682), .b(N8456), .c(N10596), .O(N10665) );
or2 gate3137( .a(N4687), .b(N10597), .O(N10668) );
inv1 gate3138( .a(N10509), .O(N10671) );
nand2 gate3139( .a(N10509), .b(N8615), .O(N10672) );
inv1 gate3140( .a(N10512), .O(N10673) );
nand2 gate3141( .a(N10512), .b(N8624), .O(N10674) );
nand2 gate3142( .a(N10609), .b(N10516), .O(N10675) );
nand2 gate3143( .a(N10610), .b(N10518), .O(N10678) );
inv1 gate3144( .a(N10519), .O(N10681) );

  xor2  gate4032(.a(N8644), .b(N10519), .O(gate3145inter0));
  nand2 gate4033(.a(gate3145inter0), .b(s_74), .O(gate3145inter1));
  and2  gate4034(.a(N8644), .b(N10519), .O(gate3145inter2));
  inv1  gate4035(.a(s_74), .O(gate3145inter3));
  inv1  gate4036(.a(s_75), .O(gate3145inter4));
  nand2 gate4037(.a(gate3145inter4), .b(gate3145inter3), .O(gate3145inter5));
  nor2  gate4038(.a(gate3145inter5), .b(gate3145inter2), .O(gate3145inter6));
  inv1  gate4039(.a(N10519), .O(gate3145inter7));
  inv1  gate4040(.a(N8644), .O(gate3145inter8));
  nand2 gate4041(.a(gate3145inter8), .b(gate3145inter7), .O(gate3145inter9));
  nand2 gate4042(.a(s_75), .b(gate3145inter3), .O(gate3145inter10));
  nor2  gate4043(.a(gate3145inter10), .b(gate3145inter9), .O(gate3145inter11));
  nor2  gate4044(.a(gate3145inter11), .b(gate3145inter6), .O(gate3145inter12));
  nand2 gate4045(.a(gate3145inter12), .b(gate3145inter1), .O(N10682));
inv1 gate3146( .a(N10522), .O(N10683) );

  xor2  gate3976(.a(N8653), .b(N10522), .O(gate3147inter0));
  nand2 gate3977(.a(gate3147inter0), .b(s_66), .O(gate3147inter1));
  and2  gate3978(.a(N8653), .b(N10522), .O(gate3147inter2));
  inv1  gate3979(.a(s_66), .O(gate3147inter3));
  inv1  gate3980(.a(s_67), .O(gate3147inter4));
  nand2 gate3981(.a(gate3147inter4), .b(gate3147inter3), .O(gate3147inter5));
  nor2  gate3982(.a(gate3147inter5), .b(gate3147inter2), .O(gate3147inter6));
  inv1  gate3983(.a(N10522), .O(gate3147inter7));
  inv1  gate3984(.a(N8653), .O(gate3147inter8));
  nand2 gate3985(.a(gate3147inter8), .b(gate3147inter7), .O(gate3147inter9));
  nand2 gate3986(.a(s_67), .b(gate3147inter3), .O(gate3147inter10));
  nor2  gate3987(.a(gate3147inter10), .b(gate3147inter9), .O(gate3147inter11));
  nor2  gate3988(.a(gate3147inter11), .b(gate3147inter6), .O(gate3147inter12));
  nand2 gate3989(.a(gate3147inter12), .b(gate3147inter1), .O(N10684));
inv1 gate3148( .a(N10525), .O(N10685) );
nand2 gate3149( .a(N10525), .b(N9454), .O(N10686) );
inv1 gate3150( .a(N10528), .O(N10687) );
nand2 gate3151( .a(N10528), .b(N9459), .O(N10688) );
inv1 gate3152( .a(N10531), .O(N10689) );
nand2 gate3153( .a(N10531), .b(N9978), .O(N10690) );

  xor2  gate3528(.a(N10535), .b(N10621), .O(gate3154inter0));
  nand2 gate3529(.a(gate3154inter0), .b(s_2), .O(gate3154inter1));
  and2  gate3530(.a(N10535), .b(N10621), .O(gate3154inter2));
  inv1  gate3531(.a(s_2), .O(gate3154inter3));
  inv1  gate3532(.a(s_3), .O(gate3154inter4));
  nand2 gate3533(.a(gate3154inter4), .b(gate3154inter3), .O(gate3154inter5));
  nor2  gate3534(.a(gate3154inter5), .b(gate3154inter2), .O(gate3154inter6));
  inv1  gate3535(.a(N10621), .O(gate3154inter7));
  inv1  gate3536(.a(N10535), .O(gate3154inter8));
  nand2 gate3537(.a(gate3154inter8), .b(gate3154inter7), .O(gate3154inter9));
  nand2 gate3538(.a(s_3), .b(gate3154inter3), .O(gate3154inter10));
  nor2  gate3539(.a(gate3154inter10), .b(gate3154inter9), .O(gate3154inter11));
  nor2  gate3540(.a(gate3154inter11), .b(gate3154inter6), .O(gate3154inter12));
  nand2 gate3541(.a(gate3154inter12), .b(gate3154inter1), .O(N10691));
inv1 gate3155( .a(N10536), .O(N10694) );
nand2 gate3156( .a(N10536), .b(N9493), .O(N10695) );
inv1 gate3157( .a(N10539), .O(N10696) );
nand2 gate3158( .a(N10539), .b(N9498), .O(N10697) );
nand2 gate3159( .a(N10626), .b(N10543), .O(N10698) );
nand2 gate3160( .a(N10627), .b(N10545), .O(N10701) );
or2 gate3161( .a(N10629), .b(N10548), .O(N10704) );
and2 gate3162( .a(N3159), .b(N10583), .O(N10705) );
or2 gate3163( .a(N10631), .b(N10551), .O(N10706) );
and2 gate3164( .a(N9737), .b(N10589), .O(N10707) );
and2 gate3165( .a(N9738), .b(N10589), .O(N10708) );
and2 gate3166( .a(N9243), .b(N10589), .O(N10709) );
and2 gate3167( .a(N5892), .b(N10589), .O(N10710) );
nand2 gate3168( .a(N10637), .b(N10558), .O(N10711) );
nand2 gate3169( .a(N10638), .b(N10560), .O(N10712) );
nand2 gate3170( .a(N10639), .b(N10562), .O(N10713) );
nand2 gate3171( .a(N10640), .b(N10564), .O(N10714) );
nand2 gate3172( .a(N10642), .b(N10567), .O(N10715) );
nand2 gate3173( .a(N10643), .b(N10569), .O(N10716) );
nand2 gate3174( .a(N10644), .b(N10571), .O(N10717) );

  xor2  gate3710(.a(N10573), .b(N10645), .O(gate3175inter0));
  nand2 gate3711(.a(gate3175inter0), .b(s_28), .O(gate3175inter1));
  and2  gate3712(.a(N10573), .b(N10645), .O(gate3175inter2));
  inv1  gate3713(.a(s_28), .O(gate3175inter3));
  inv1  gate3714(.a(s_29), .O(gate3175inter4));
  nand2 gate3715(.a(gate3175inter4), .b(gate3175inter3), .O(gate3175inter5));
  nor2  gate3716(.a(gate3175inter5), .b(gate3175inter2), .O(gate3175inter6));
  inv1  gate3717(.a(N10645), .O(gate3175inter7));
  inv1  gate3718(.a(N10573), .O(gate3175inter8));
  nand2 gate3719(.a(gate3175inter8), .b(gate3175inter7), .O(gate3175inter9));
  nand2 gate3720(.a(s_29), .b(gate3175inter3), .O(gate3175inter10));
  nor2  gate3721(.a(gate3175inter10), .b(gate3175inter9), .O(gate3175inter11));
  nor2  gate3722(.a(gate3175inter11), .b(gate3175inter6), .O(gate3175inter12));
  nand2 gate3723(.a(gate3175inter12), .b(gate3175inter1), .O(N10718));
inv1 gate3176( .a(N10602), .O(N10719) );
nand2 gate3177( .a(N10602), .b(N9244), .O(N10720) );
inv1 gate3178( .a(N10647), .O(N10729) );
and2 gate3179( .a(N5178), .b(N10583), .O(N10730) );
and2 gate3180( .a(N2533), .b(N10583), .O(N10731) );
nand2 gate3181( .a(N7447), .b(N10671), .O(N10737) );
nand2 gate3182( .a(N7465), .b(N10673), .O(N10738) );
or4 gate3183( .a(N10648), .b(N10649), .c(N10581), .d(N10582), .O(N10739) );

  xor2  gate3514(.a(N10681), .b(N7503), .O(gate3184inter0));
  nand2 gate3515(.a(gate3184inter0), .b(s_0), .O(gate3184inter1));
  and2  gate3516(.a(N10681), .b(N7503), .O(gate3184inter2));
  inv1  gate3517(.a(s_0), .O(gate3184inter3));
  inv1  gate3518(.a(s_1), .O(gate3184inter4));
  nand2 gate3519(.a(gate3184inter4), .b(gate3184inter3), .O(gate3184inter5));
  nor2  gate3520(.a(gate3184inter5), .b(gate3184inter2), .O(gate3184inter6));
  inv1  gate3521(.a(N7503), .O(gate3184inter7));
  inv1  gate3522(.a(N10681), .O(gate3184inter8));
  nand2 gate3523(.a(gate3184inter8), .b(gate3184inter7), .O(gate3184inter9));
  nand2 gate3524(.a(s_1), .b(gate3184inter3), .O(gate3184inter10));
  nor2  gate3525(.a(gate3184inter10), .b(gate3184inter9), .O(gate3184inter11));
  nor2  gate3526(.a(gate3184inter11), .b(gate3184inter6), .O(gate3184inter12));
  nand2 gate3527(.a(gate3184inter12), .b(gate3184inter1), .O(N10746));
nand2 gate3185( .a(N7521), .b(N10683), .O(N10747) );

  xor2  gate4452(.a(N10685), .b(N8678), .O(gate3186inter0));
  nand2 gate4453(.a(gate3186inter0), .b(s_134), .O(gate3186inter1));
  and2  gate4454(.a(N10685), .b(N8678), .O(gate3186inter2));
  inv1  gate4455(.a(s_134), .O(gate3186inter3));
  inv1  gate4456(.a(s_135), .O(gate3186inter4));
  nand2 gate4457(.a(gate3186inter4), .b(gate3186inter3), .O(gate3186inter5));
  nor2  gate4458(.a(gate3186inter5), .b(gate3186inter2), .O(gate3186inter6));
  inv1  gate4459(.a(N8678), .O(gate3186inter7));
  inv1  gate4460(.a(N10685), .O(gate3186inter8));
  nand2 gate4461(.a(gate3186inter8), .b(gate3186inter7), .O(gate3186inter9));
  nand2 gate4462(.a(s_135), .b(gate3186inter3), .O(gate3186inter10));
  nor2  gate4463(.a(gate3186inter10), .b(gate3186inter9), .O(gate3186inter11));
  nor2  gate4464(.a(gate3186inter11), .b(gate3186inter6), .O(gate3186inter12));
  nand2 gate4465(.a(gate3186inter12), .b(gate3186inter1), .O(N10748));
nand2 gate3187( .a(N8690), .b(N10687), .O(N10749) );
nand2 gate3188( .a(N9685), .b(N10689), .O(N10750) );
nand2 gate3189( .a(N8757), .b(N10694), .O(N10753) );
nand2 gate3190( .a(N8769), .b(N10696), .O(N10754) );
or2 gate3191( .a(N10705), .b(N10549), .O(N10759) );
or2 gate3192( .a(N10707), .b(N10553), .O(N10760) );
or2 gate3193( .a(N10708), .b(N10554), .O(N10761) );
or2 gate3194( .a(N10709), .b(N10555), .O(N10762) );
or2 gate3195( .a(N10710), .b(N10556), .O(N10763) );
nand2 gate3196( .a(N8580), .b(N10719), .O(N10764) );
and2 gate3197( .a(N10652), .b(N9890), .O(N10765) );
and2 gate3198( .a(N10652), .b(N9891), .O(N10766) );
and2 gate3199( .a(N10652), .b(N9892), .O(N10767) );
and2 gate3200( .a(N10652), .b(N8252), .O(N10768) );
inv1 gate3201( .a(N10659), .O(N10769) );
nand2 gate3202( .a(N10659), .b(N9245), .O(N10770) );
inv1 gate3203( .a(N10662), .O(N10771) );

  xor2  gate4774(.a(N9246), .b(N10662), .O(gate3204inter0));
  nand2 gate4775(.a(gate3204inter0), .b(s_180), .O(gate3204inter1));
  and2  gate4776(.a(N9246), .b(N10662), .O(gate3204inter2));
  inv1  gate4777(.a(s_180), .O(gate3204inter3));
  inv1  gate4778(.a(s_181), .O(gate3204inter4));
  nand2 gate4779(.a(gate3204inter4), .b(gate3204inter3), .O(gate3204inter5));
  nor2  gate4780(.a(gate3204inter5), .b(gate3204inter2), .O(gate3204inter6));
  inv1  gate4781(.a(N10662), .O(gate3204inter7));
  inv1  gate4782(.a(N9246), .O(gate3204inter8));
  nand2 gate4783(.a(gate3204inter8), .b(gate3204inter7), .O(gate3204inter9));
  nand2 gate4784(.a(s_181), .b(gate3204inter3), .O(gate3204inter10));
  nor2  gate4785(.a(gate3204inter10), .b(gate3204inter9), .O(gate3204inter11));
  nor2  gate4786(.a(gate3204inter11), .b(gate3204inter6), .O(gate3204inter12));
  nand2 gate4787(.a(gate3204inter12), .b(gate3204inter1), .O(N10772));
inv1 gate3205( .a(N10665), .O(N10773) );
nand2 gate3206( .a(N10665), .b(N9247), .O(N10774) );
inv1 gate3207( .a(N10668), .O(N10775) );
nand2 gate3208( .a(N10668), .b(N9248), .O(N10776) );
or2 gate3209( .a(N10730), .b(N10587), .O(N10778) );
or2 gate3210( .a(N10731), .b(N10588), .O(N10781) );
inv1 gate3211( .a(N10652), .O(N10784) );

  xor2  gate5166(.a(N10672), .b(N10737), .O(gate3212inter0));
  nand2 gate5167(.a(gate3212inter0), .b(s_236), .O(gate3212inter1));
  and2  gate5168(.a(N10672), .b(N10737), .O(gate3212inter2));
  inv1  gate5169(.a(s_236), .O(gate3212inter3));
  inv1  gate5170(.a(s_237), .O(gate3212inter4));
  nand2 gate5171(.a(gate3212inter4), .b(gate3212inter3), .O(gate3212inter5));
  nor2  gate5172(.a(gate3212inter5), .b(gate3212inter2), .O(gate3212inter6));
  inv1  gate5173(.a(N10737), .O(gate3212inter7));
  inv1  gate5174(.a(N10672), .O(gate3212inter8));
  nand2 gate5175(.a(gate3212inter8), .b(gate3212inter7), .O(gate3212inter9));
  nand2 gate5176(.a(s_237), .b(gate3212inter3), .O(gate3212inter10));
  nor2  gate5177(.a(gate3212inter10), .b(gate3212inter9), .O(gate3212inter11));
  nor2  gate5178(.a(gate3212inter11), .b(gate3212inter6), .O(gate3212inter12));
  nand2 gate5179(.a(gate3212inter12), .b(gate3212inter1), .O(N10789));
nand2 gate3213( .a(N10738), .b(N10674), .O(N10792) );
inv1 gate3214( .a(N10675), .O(N10796) );

  xor2  gate5124(.a(N8633), .b(N10675), .O(gate3215inter0));
  nand2 gate5125(.a(gate3215inter0), .b(s_230), .O(gate3215inter1));
  and2  gate5126(.a(N8633), .b(N10675), .O(gate3215inter2));
  inv1  gate5127(.a(s_230), .O(gate3215inter3));
  inv1  gate5128(.a(s_231), .O(gate3215inter4));
  nand2 gate5129(.a(gate3215inter4), .b(gate3215inter3), .O(gate3215inter5));
  nor2  gate5130(.a(gate3215inter5), .b(gate3215inter2), .O(gate3215inter6));
  inv1  gate5131(.a(N10675), .O(gate3215inter7));
  inv1  gate5132(.a(N8633), .O(gate3215inter8));
  nand2 gate5133(.a(gate3215inter8), .b(gate3215inter7), .O(gate3215inter9));
  nand2 gate5134(.a(s_231), .b(gate3215inter3), .O(gate3215inter10));
  nor2  gate5135(.a(gate3215inter10), .b(gate3215inter9), .O(gate3215inter11));
  nor2  gate5136(.a(gate3215inter11), .b(gate3215inter6), .O(gate3215inter12));
  nand2 gate5137(.a(gate3215inter12), .b(gate3215inter1), .O(N10797));
inv1 gate3216( .a(N10678), .O(N10798) );

  xor2  gate4802(.a(N8638), .b(N10678), .O(gate3217inter0));
  nand2 gate4803(.a(gate3217inter0), .b(s_184), .O(gate3217inter1));
  and2  gate4804(.a(N8638), .b(N10678), .O(gate3217inter2));
  inv1  gate4805(.a(s_184), .O(gate3217inter3));
  inv1  gate4806(.a(s_185), .O(gate3217inter4));
  nand2 gate4807(.a(gate3217inter4), .b(gate3217inter3), .O(gate3217inter5));
  nor2  gate4808(.a(gate3217inter5), .b(gate3217inter2), .O(gate3217inter6));
  inv1  gate4809(.a(N10678), .O(gate3217inter7));
  inv1  gate4810(.a(N8638), .O(gate3217inter8));
  nand2 gate4811(.a(gate3217inter8), .b(gate3217inter7), .O(gate3217inter9));
  nand2 gate4812(.a(s_185), .b(gate3217inter3), .O(gate3217inter10));
  nor2  gate4813(.a(gate3217inter10), .b(gate3217inter9), .O(gate3217inter11));
  nor2  gate4814(.a(gate3217inter11), .b(gate3217inter6), .O(gate3217inter12));
  nand2 gate4815(.a(gate3217inter12), .b(gate3217inter1), .O(N10799));
nand2 gate3218( .a(N10746), .b(N10682), .O(N10800) );
nand2 gate3219( .a(N10747), .b(N10684), .O(N10803) );
nand2 gate3220( .a(N10748), .b(N10686), .O(N10806) );
nand2 gate3221( .a(N10749), .b(N10688), .O(N10809) );
nand2 gate3222( .a(N10750), .b(N10690), .O(N10812) );
inv1 gate3223( .a(N10691), .O(N10815) );
nand2 gate3224( .a(N10691), .b(N9866), .O(N10816) );
nand2 gate3225( .a(N10753), .b(N10695), .O(N10817) );
nand2 gate3226( .a(N10754), .b(N10697), .O(N10820) );
inv1 gate3227( .a(N10698), .O(N10823) );
nand2 gate3228( .a(N10698), .b(N9505), .O(N10824) );
inv1 gate3229( .a(N10701), .O(N10825) );
nand2 gate3230( .a(N10701), .b(N9514), .O(N10826) );
nand2 gate3231( .a(N10764), .b(N10720), .O(N10827) );
nand2 gate3232( .a(N8583), .b(N10769), .O(N10832) );
nand2 gate3233( .a(N8586), .b(N10771), .O(N10833) );
nand2 gate3234( .a(N8589), .b(N10773), .O(N10834) );
nand2 gate3235( .a(N8592), .b(N10775), .O(N10835) );
inv1 gate3236( .a(N10739), .O(N10836) );
buf1 gate3237( .a(N10778), .O(N10837) );
buf1 gate3238( .a(N10778), .O(N10838) );
buf1 gate3239( .a(N10781), .O(N10839) );
buf1 gate3240( .a(N10781), .O(N10840) );
nand2 gate3241( .a(N7482), .b(N10796), .O(N10845) );
nand2 gate3242( .a(N7494), .b(N10798), .O(N10846) );

  xor2  gate3934(.a(N10815), .b(N9473), .O(gate3243inter0));
  nand2 gate3935(.a(gate3243inter0), .b(s_60), .O(gate3243inter1));
  and2  gate3936(.a(N10815), .b(N9473), .O(gate3243inter2));
  inv1  gate3937(.a(s_60), .O(gate3243inter3));
  inv1  gate3938(.a(s_61), .O(gate3243inter4));
  nand2 gate3939(.a(gate3243inter4), .b(gate3243inter3), .O(gate3243inter5));
  nor2  gate3940(.a(gate3243inter5), .b(gate3243inter2), .O(gate3243inter6));
  inv1  gate3941(.a(N9473), .O(gate3243inter7));
  inv1  gate3942(.a(N10815), .O(gate3243inter8));
  nand2 gate3943(.a(gate3243inter8), .b(gate3243inter7), .O(gate3243inter9));
  nand2 gate3944(.a(s_61), .b(gate3243inter3), .O(gate3243inter10));
  nor2  gate3945(.a(gate3243inter10), .b(gate3243inter9), .O(gate3243inter11));
  nor2  gate3946(.a(gate3243inter11), .b(gate3243inter6), .O(gate3243inter12));
  nand2 gate3947(.a(gate3243inter12), .b(gate3243inter1), .O(N10857));

  xor2  gate4158(.a(N10823), .b(N8781), .O(gate3244inter0));
  nand2 gate4159(.a(gate3244inter0), .b(s_92), .O(gate3244inter1));
  and2  gate4160(.a(N10823), .b(N8781), .O(gate3244inter2));
  inv1  gate4161(.a(s_92), .O(gate3244inter3));
  inv1  gate4162(.a(s_93), .O(gate3244inter4));
  nand2 gate4163(.a(gate3244inter4), .b(gate3244inter3), .O(gate3244inter5));
  nor2  gate4164(.a(gate3244inter5), .b(gate3244inter2), .O(gate3244inter6));
  inv1  gate4165(.a(N8781), .O(gate3244inter7));
  inv1  gate4166(.a(N10823), .O(gate3244inter8));
  nand2 gate4167(.a(gate3244inter8), .b(gate3244inter7), .O(gate3244inter9));
  nand2 gate4168(.a(s_93), .b(gate3244inter3), .O(gate3244inter10));
  nor2  gate4169(.a(gate3244inter10), .b(gate3244inter9), .O(gate3244inter11));
  nor2  gate4170(.a(gate3244inter11), .b(gate3244inter6), .O(gate3244inter12));
  nand2 gate4171(.a(gate3244inter12), .b(gate3244inter1), .O(N10862));
nand2 gate3245( .a(N8799), .b(N10825), .O(N10863) );
and2 gate3246( .a(N10023), .b(N10784), .O(N10864) );
and2 gate3247( .a(N10024), .b(N10784), .O(N10865) );
and2 gate3248( .a(N9739), .b(N10784), .O(N10866) );
and2 gate3249( .a(N7136), .b(N10784), .O(N10867) );
nand2 gate3250( .a(N10832), .b(N10770), .O(N10868) );
nand2 gate3251( .a(N10833), .b(N10772), .O(N10869) );
nand2 gate3252( .a(N10834), .b(N10774), .O(N10870) );
nand2 gate3253( .a(N10835), .b(N10776), .O(N10871) );
inv1 gate3254( .a(N10789), .O(N10872) );
nand2 gate3255( .a(N10789), .b(N8616), .O(N10873) );
inv1 gate3256( .a(N10792), .O(N10874) );
nand2 gate3257( .a(N10792), .b(N8625), .O(N10875) );
nand2 gate3258( .a(N10845), .b(N10797), .O(N10876) );
nand2 gate3259( .a(N10846), .b(N10799), .O(N10879) );
inv1 gate3260( .a(N10800), .O(N10882) );
nand2 gate3261( .a(N10800), .b(N8645), .O(N10883) );
inv1 gate3262( .a(N10803), .O(N10884) );
nand2 gate3263( .a(N10803), .b(N8654), .O(N10885) );
inv1 gate3264( .a(N10806), .O(N10886) );
nand2 gate3265( .a(N10806), .b(N9455), .O(N10887) );
inv1 gate3266( .a(N10809), .O(N10888) );
nand2 gate3267( .a(N10809), .b(N9460), .O(N10889) );
inv1 gate3268( .a(N10812), .O(N10890) );
nand2 gate3269( .a(N10812), .b(N9862), .O(N10891) );
nand2 gate3270( .a(N10857), .b(N10816), .O(N10892) );
inv1 gate3271( .a(N10817), .O(N10895) );
nand2 gate3272( .a(N10817), .b(N9494), .O(N10896) );
inv1 gate3273( .a(N10820), .O(N10897) );
nand2 gate3274( .a(N10820), .b(N9499), .O(N10898) );
nand2 gate3275( .a(N10862), .b(N10824), .O(N10899) );
nand2 gate3276( .a(N10863), .b(N10826), .O(N10902) );
or2 gate3277( .a(N10864), .b(N10765), .O(N10905) );
or2 gate3278( .a(N10865), .b(N10766), .O(N10906) );
or2 gate3279( .a(N10866), .b(N10767), .O(N10907) );
or2 gate3280( .a(N10867), .b(N10768), .O(N10908) );
nand2 gate3281( .a(N7450), .b(N10872), .O(N10909) );
nand2 gate3282( .a(N7468), .b(N10874), .O(N10910) );
nand2 gate3283( .a(N7506), .b(N10882), .O(N10915) );
nand2 gate3284( .a(N7524), .b(N10884), .O(N10916) );
nand2 gate3285( .a(N8681), .b(N10886), .O(N10917) );
nand2 gate3286( .a(N8693), .b(N10888), .O(N10918) );
nand2 gate3287( .a(N9462), .b(N10890), .O(N10919) );
nand2 gate3288( .a(N8760), .b(N10895), .O(N10922) );
nand2 gate3289( .a(N8772), .b(N10897), .O(N10923) );
nand2 gate3290( .a(N10909), .b(N10873), .O(N10928) );
nand2 gate3291( .a(N10910), .b(N10875), .O(N10931) );
inv1 gate3292( .a(N10876), .O(N10934) );
nand2 gate3293( .a(N10876), .b(N8634), .O(N10935) );
inv1 gate3294( .a(N10879), .O(N10936) );
nand2 gate3295( .a(N10879), .b(N8639), .O(N10937) );

  xor2  gate5040(.a(N10883), .b(N10915), .O(gate3296inter0));
  nand2 gate5041(.a(gate3296inter0), .b(s_218), .O(gate3296inter1));
  and2  gate5042(.a(N10883), .b(N10915), .O(gate3296inter2));
  inv1  gate5043(.a(s_218), .O(gate3296inter3));
  inv1  gate5044(.a(s_219), .O(gate3296inter4));
  nand2 gate5045(.a(gate3296inter4), .b(gate3296inter3), .O(gate3296inter5));
  nor2  gate5046(.a(gate3296inter5), .b(gate3296inter2), .O(gate3296inter6));
  inv1  gate5047(.a(N10915), .O(gate3296inter7));
  inv1  gate5048(.a(N10883), .O(gate3296inter8));
  nand2 gate5049(.a(gate3296inter8), .b(gate3296inter7), .O(gate3296inter9));
  nand2 gate5050(.a(s_219), .b(gate3296inter3), .O(gate3296inter10));
  nor2  gate5051(.a(gate3296inter10), .b(gate3296inter9), .O(gate3296inter11));
  nor2  gate5052(.a(gate3296inter11), .b(gate3296inter6), .O(gate3296inter12));
  nand2 gate5053(.a(gate3296inter12), .b(gate3296inter1), .O(N10938));
nand2 gate3297( .a(N10916), .b(N10885), .O(N10941) );

  xor2  gate5222(.a(N10887), .b(N10917), .O(gate3298inter0));
  nand2 gate5223(.a(gate3298inter0), .b(s_244), .O(gate3298inter1));
  and2  gate5224(.a(N10887), .b(N10917), .O(gate3298inter2));
  inv1  gate5225(.a(s_244), .O(gate3298inter3));
  inv1  gate5226(.a(s_245), .O(gate3298inter4));
  nand2 gate5227(.a(gate3298inter4), .b(gate3298inter3), .O(gate3298inter5));
  nor2  gate5228(.a(gate3298inter5), .b(gate3298inter2), .O(gate3298inter6));
  inv1  gate5229(.a(N10917), .O(gate3298inter7));
  inv1  gate5230(.a(N10887), .O(gate3298inter8));
  nand2 gate5231(.a(gate3298inter8), .b(gate3298inter7), .O(gate3298inter9));
  nand2 gate5232(.a(s_245), .b(gate3298inter3), .O(gate3298inter10));
  nor2  gate5233(.a(gate3298inter10), .b(gate3298inter9), .O(gate3298inter11));
  nor2  gate5234(.a(gate3298inter11), .b(gate3298inter6), .O(gate3298inter12));
  nand2 gate5235(.a(gate3298inter12), .b(gate3298inter1), .O(N10944));
nand2 gate3299( .a(N10918), .b(N10889), .O(N10947) );
nand2 gate3300( .a(N10919), .b(N10891), .O(N10950) );
inv1 gate3301( .a(N10892), .O(N10953) );
nand2 gate3302( .a(N10892), .b(N9476), .O(N10954) );
nand2 gate3303( .a(N10922), .b(N10896), .O(N10955) );

  xor2  gate4984(.a(N10898), .b(N10923), .O(gate3304inter0));
  nand2 gate4985(.a(gate3304inter0), .b(s_210), .O(gate3304inter1));
  and2  gate4986(.a(N10898), .b(N10923), .O(gate3304inter2));
  inv1  gate4987(.a(s_210), .O(gate3304inter3));
  inv1  gate4988(.a(s_211), .O(gate3304inter4));
  nand2 gate4989(.a(gate3304inter4), .b(gate3304inter3), .O(gate3304inter5));
  nor2  gate4990(.a(gate3304inter5), .b(gate3304inter2), .O(gate3304inter6));
  inv1  gate4991(.a(N10923), .O(gate3304inter7));
  inv1  gate4992(.a(N10898), .O(gate3304inter8));
  nand2 gate4993(.a(gate3304inter8), .b(gate3304inter7), .O(gate3304inter9));
  nand2 gate4994(.a(s_211), .b(gate3304inter3), .O(gate3304inter10));
  nor2  gate4995(.a(gate3304inter10), .b(gate3304inter9), .O(gate3304inter11));
  nor2  gate4996(.a(gate3304inter11), .b(gate3304inter6), .O(gate3304inter12));
  nand2 gate4997(.a(gate3304inter12), .b(gate3304inter1), .O(N10958));
inv1 gate3305( .a(N10899), .O(N10961) );
nand2 gate3306( .a(N10899), .b(N9506), .O(N10962) );
inv1 gate3307( .a(N10902), .O(N10963) );
nand2 gate3308( .a(N10902), .b(N9515), .O(N10964) );
nand2 gate3309( .a(N7485), .b(N10934), .O(N10969) );
nand2 gate3310( .a(N7497), .b(N10936), .O(N10970) );
nand2 gate3311( .a(N8718), .b(N10953), .O(N10981) );
nand2 gate3312( .a(N8784), .b(N10961), .O(N10986) );
nand2 gate3313( .a(N8802), .b(N10963), .O(N10987) );
inv1 gate3314( .a(N10928), .O(N10988) );
nand2 gate3315( .a(N10928), .b(N8617), .O(N10989) );
inv1 gate3316( .a(N10931), .O(N10990) );
nand2 gate3317( .a(N10931), .b(N8626), .O(N10991) );
nand2 gate3318( .a(N10969), .b(N10935), .O(N10992) );
nand2 gate3319( .a(N10970), .b(N10937), .O(N10995) );
inv1 gate3320( .a(N10938), .O(N10998) );
nand2 gate3321( .a(N10938), .b(N8646), .O(N10999) );
inv1 gate3322( .a(N10941), .O(N11000) );
nand2 gate3323( .a(N10941), .b(N8655), .O(N11001) );
inv1 gate3324( .a(N10944), .O(N11002) );
nand2 gate3325( .a(N10944), .b(N9456), .O(N11003) );
inv1 gate3326( .a(N10947), .O(N11004) );
nand2 gate3327( .a(N10947), .b(N9461), .O(N11005) );
inv1 gate3328( .a(N10950), .O(N11006) );

  xor2  gate4732(.a(N9465), .b(N10950), .O(gate3329inter0));
  nand2 gate4733(.a(gate3329inter0), .b(s_174), .O(gate3329inter1));
  and2  gate4734(.a(N9465), .b(N10950), .O(gate3329inter2));
  inv1  gate4735(.a(s_174), .O(gate3329inter3));
  inv1  gate4736(.a(s_175), .O(gate3329inter4));
  nand2 gate4737(.a(gate3329inter4), .b(gate3329inter3), .O(gate3329inter5));
  nor2  gate4738(.a(gate3329inter5), .b(gate3329inter2), .O(gate3329inter6));
  inv1  gate4739(.a(N10950), .O(gate3329inter7));
  inv1  gate4740(.a(N9465), .O(gate3329inter8));
  nand2 gate4741(.a(gate3329inter8), .b(gate3329inter7), .O(gate3329inter9));
  nand2 gate4742(.a(s_175), .b(gate3329inter3), .O(gate3329inter10));
  nor2  gate4743(.a(gate3329inter10), .b(gate3329inter9), .O(gate3329inter11));
  nor2  gate4744(.a(gate3329inter11), .b(gate3329inter6), .O(gate3329inter12));
  nand2 gate4745(.a(gate3329inter12), .b(gate3329inter1), .O(N11007));
nand2 gate3330( .a(N10981), .b(N10954), .O(N11008) );
inv1 gate3331( .a(N10955), .O(N11011) );
nand2 gate3332( .a(N10955), .b(N9495), .O(N11012) );
inv1 gate3333( .a(N10958), .O(N11013) );
nand2 gate3334( .a(N10958), .b(N9500), .O(N11014) );
nand2 gate3335( .a(N10986), .b(N10962), .O(N11015) );

  xor2  gate3990(.a(N10964), .b(N10987), .O(gate3336inter0));
  nand2 gate3991(.a(gate3336inter0), .b(s_68), .O(gate3336inter1));
  and2  gate3992(.a(N10964), .b(N10987), .O(gate3336inter2));
  inv1  gate3993(.a(s_68), .O(gate3336inter3));
  inv1  gate3994(.a(s_69), .O(gate3336inter4));
  nand2 gate3995(.a(gate3336inter4), .b(gate3336inter3), .O(gate3336inter5));
  nor2  gate3996(.a(gate3336inter5), .b(gate3336inter2), .O(gate3336inter6));
  inv1  gate3997(.a(N10987), .O(gate3336inter7));
  inv1  gate3998(.a(N10964), .O(gate3336inter8));
  nand2 gate3999(.a(gate3336inter8), .b(gate3336inter7), .O(gate3336inter9));
  nand2 gate4000(.a(s_69), .b(gate3336inter3), .O(gate3336inter10));
  nor2  gate4001(.a(gate3336inter10), .b(gate3336inter9), .O(gate3336inter11));
  nor2  gate4002(.a(gate3336inter11), .b(gate3336inter6), .O(gate3336inter12));
  nand2 gate4003(.a(gate3336inter12), .b(gate3336inter1), .O(N11018));
nand2 gate3337( .a(N7453), .b(N10988), .O(N11023) );
nand2 gate3338( .a(N7471), .b(N10990), .O(N11024) );
nand2 gate3339( .a(N7509), .b(N10998), .O(N11027) );
nand2 gate3340( .a(N7527), .b(N11000), .O(N11028) );
nand2 gate3341( .a(N8684), .b(N11002), .O(N11029) );
nand2 gate3342( .a(N8696), .b(N11004), .O(N11030) );
nand2 gate3343( .a(N8702), .b(N11006), .O(N11031) );
nand2 gate3344( .a(N8763), .b(N11011), .O(N11034) );
nand2 gate3345( .a(N8775), .b(N11013), .O(N11035) );
inv1 gate3346( .a(N10992), .O(N11040) );
nand2 gate3347( .a(N10992), .b(N8294), .O(N11041) );
inv1 gate3348( .a(N10995), .O(N11042) );
nand2 gate3349( .a(N10995), .b(N8295), .O(N11043) );
nand2 gate3350( .a(N11023), .b(N10989), .O(N11044) );
nand2 gate3351( .a(N11024), .b(N10991), .O(N11047) );
nand2 gate3352( .a(N11027), .b(N10999), .O(N11050) );
nand2 gate3353( .a(N11028), .b(N11001), .O(N11053) );
nand2 gate3354( .a(N11029), .b(N11003), .O(N11056) );
nand2 gate3355( .a(N11030), .b(N11005), .O(N11059) );
nand2 gate3356( .a(N11031), .b(N11007), .O(N11062) );
inv1 gate3357( .a(N11008), .O(N11065) );
nand2 gate3358( .a(N11008), .b(N9477), .O(N11066) );
nand2 gate3359( .a(N11034), .b(N11012), .O(N11067) );
nand2 gate3360( .a(N11035), .b(N11014), .O(N11070) );
inv1 gate3361( .a(N11015), .O(N11073) );
nand2 gate3362( .a(N11015), .b(N9507), .O(N11074) );
inv1 gate3363( .a(N11018), .O(N11075) );
nand2 gate3364( .a(N11018), .b(N9516), .O(N11076) );
nand2 gate3365( .a(N7488), .b(N11040), .O(N11077) );
nand2 gate3366( .a(N7500), .b(N11042), .O(N11078) );

  xor2  gate4396(.a(N11065), .b(N8721), .O(gate3367inter0));
  nand2 gate4397(.a(gate3367inter0), .b(s_126), .O(gate3367inter1));
  and2  gate4398(.a(N11065), .b(N8721), .O(gate3367inter2));
  inv1  gate4399(.a(s_126), .O(gate3367inter3));
  inv1  gate4400(.a(s_127), .O(gate3367inter4));
  nand2 gate4401(.a(gate3367inter4), .b(gate3367inter3), .O(gate3367inter5));
  nor2  gate4402(.a(gate3367inter5), .b(gate3367inter2), .O(gate3367inter6));
  inv1  gate4403(.a(N8721), .O(gate3367inter7));
  inv1  gate4404(.a(N11065), .O(gate3367inter8));
  nand2 gate4405(.a(gate3367inter8), .b(gate3367inter7), .O(gate3367inter9));
  nand2 gate4406(.a(s_127), .b(gate3367inter3), .O(gate3367inter10));
  nor2  gate4407(.a(gate3367inter10), .b(gate3367inter9), .O(gate3367inter11));
  nor2  gate4408(.a(gate3367inter11), .b(gate3367inter6), .O(gate3367inter12));
  nand2 gate4409(.a(gate3367inter12), .b(gate3367inter1), .O(N11095));
nand2 gate3368( .a(N8787), .b(N11073), .O(N11098) );
nand2 gate3369( .a(N8805), .b(N11075), .O(N11099) );
nand2 gate3370( .a(N11077), .b(N11041), .O(N11100) );
nand2 gate3371( .a(N11078), .b(N11043), .O(N11103) );
inv1 gate3372( .a(N11056), .O(N11106) );
nand2 gate3373( .a(N11056), .b(N9319), .O(N11107) );
inv1 gate3374( .a(N11059), .O(N11108) );
nand2 gate3375( .a(N11059), .b(N9320), .O(N11109) );
inv1 gate3376( .a(N11067), .O(N11110) );

  xor2  gate3808(.a(N9381), .b(N11067), .O(gate3377inter0));
  nand2 gate3809(.a(gate3377inter0), .b(s_42), .O(gate3377inter1));
  and2  gate3810(.a(N9381), .b(N11067), .O(gate3377inter2));
  inv1  gate3811(.a(s_42), .O(gate3377inter3));
  inv1  gate3812(.a(s_43), .O(gate3377inter4));
  nand2 gate3813(.a(gate3377inter4), .b(gate3377inter3), .O(gate3377inter5));
  nor2  gate3814(.a(gate3377inter5), .b(gate3377inter2), .O(gate3377inter6));
  inv1  gate3815(.a(N11067), .O(gate3377inter7));
  inv1  gate3816(.a(N9381), .O(gate3377inter8));
  nand2 gate3817(.a(gate3377inter8), .b(gate3377inter7), .O(gate3377inter9));
  nand2 gate3818(.a(s_43), .b(gate3377inter3), .O(gate3377inter10));
  nor2  gate3819(.a(gate3377inter10), .b(gate3377inter9), .O(gate3377inter11));
  nor2  gate3820(.a(gate3377inter11), .b(gate3377inter6), .O(gate3377inter12));
  nand2 gate3821(.a(gate3377inter12), .b(gate3377inter1), .O(N11111));
inv1 gate3378( .a(N11070), .O(N11112) );
nand2 gate3379( .a(N11070), .b(N9382), .O(N11113) );
inv1 gate3380( .a(N11044), .O(N11114) );

  xor2  gate4494(.a(N8618), .b(N11044), .O(gate3381inter0));
  nand2 gate4495(.a(gate3381inter0), .b(s_140), .O(gate3381inter1));
  and2  gate4496(.a(N8618), .b(N11044), .O(gate3381inter2));
  inv1  gate4497(.a(s_140), .O(gate3381inter3));
  inv1  gate4498(.a(s_141), .O(gate3381inter4));
  nand2 gate4499(.a(gate3381inter4), .b(gate3381inter3), .O(gate3381inter5));
  nor2  gate4500(.a(gate3381inter5), .b(gate3381inter2), .O(gate3381inter6));
  inv1  gate4501(.a(N11044), .O(gate3381inter7));
  inv1  gate4502(.a(N8618), .O(gate3381inter8));
  nand2 gate4503(.a(gate3381inter8), .b(gate3381inter7), .O(gate3381inter9));
  nand2 gate4504(.a(s_141), .b(gate3381inter3), .O(gate3381inter10));
  nor2  gate4505(.a(gate3381inter10), .b(gate3381inter9), .O(gate3381inter11));
  nor2  gate4506(.a(gate3381inter11), .b(gate3381inter6), .O(gate3381inter12));
  nand2 gate4507(.a(gate3381inter12), .b(gate3381inter1), .O(N11115));
inv1 gate3382( .a(N11047), .O(N11116) );
nand2 gate3383( .a(N11047), .b(N8619), .O(N11117) );
inv1 gate3384( .a(N11050), .O(N11118) );
nand2 gate3385( .a(N11050), .b(N8647), .O(N11119) );
inv1 gate3386( .a(N11053), .O(N11120) );
nand2 gate3387( .a(N11053), .b(N8648), .O(N11121) );
inv1 gate3388( .a(N11062), .O(N11122) );
nand2 gate3389( .a(N11062), .b(N9466), .O(N11123) );
nand2 gate3390( .a(N11095), .b(N11066), .O(N11124) );
nand2 gate3391( .a(N11098), .b(N11074), .O(N11127) );
nand2 gate3392( .a(N11099), .b(N11076), .O(N11130) );
nand2 gate3393( .a(N8687), .b(N11106), .O(N11137) );
nand2 gate3394( .a(N8699), .b(N11108), .O(N11138) );
nand2 gate3395( .a(N8766), .b(N11110), .O(N11139) );

  xor2  gate5250(.a(N11112), .b(N8778), .O(gate3396inter0));
  nand2 gate5251(.a(gate3396inter0), .b(s_248), .O(gate3396inter1));
  and2  gate5252(.a(N11112), .b(N8778), .O(gate3396inter2));
  inv1  gate5253(.a(s_248), .O(gate3396inter3));
  inv1  gate5254(.a(s_249), .O(gate3396inter4));
  nand2 gate5255(.a(gate3396inter4), .b(gate3396inter3), .O(gate3396inter5));
  nor2  gate5256(.a(gate3396inter5), .b(gate3396inter2), .O(gate3396inter6));
  inv1  gate5257(.a(N8778), .O(gate3396inter7));
  inv1  gate5258(.a(N11112), .O(gate3396inter8));
  nand2 gate5259(.a(gate3396inter8), .b(gate3396inter7), .O(gate3396inter9));
  nand2 gate5260(.a(s_249), .b(gate3396inter3), .O(gate3396inter10));
  nor2  gate5261(.a(gate3396inter10), .b(gate3396inter9), .O(gate3396inter11));
  nor2  gate5262(.a(gate3396inter11), .b(gate3396inter6), .O(gate3396inter12));
  nand2 gate5263(.a(gate3396inter12), .b(gate3396inter1), .O(N11140));
nand2 gate3397( .a(N7456), .b(N11114), .O(N11141) );
nand2 gate3398( .a(N7474), .b(N11116), .O(N11142) );
nand2 gate3399( .a(N7512), .b(N11118), .O(N11143) );
nand2 gate3400( .a(N7530), .b(N11120), .O(N11144) );
nand2 gate3401( .a(N8705), .b(N11122), .O(N11145) );
and3 gate3402( .a(N11103), .b(N8871), .c(N10283), .O(N11152) );
and3 gate3403( .a(N11100), .b(N7655), .c(N10283), .O(N11153) );
and3 gate3404( .a(N11103), .b(N9551), .c(N10119), .O(N11154) );
and3 gate3405( .a(N11100), .b(N9917), .c(N10119), .O(N11155) );
nand2 gate3406( .a(N11137), .b(N11107), .O(N11156) );
nand2 gate3407( .a(N11138), .b(N11109), .O(N11159) );
nand2 gate3408( .a(N11139), .b(N11111), .O(N11162) );
nand2 gate3409( .a(N11140), .b(N11113), .O(N11165) );
nand2 gate3410( .a(N11141), .b(N11115), .O(N11168) );
nand2 gate3411( .a(N11142), .b(N11117), .O(N11171) );
nand2 gate3412( .a(N11143), .b(N11119), .O(N11174) );

  xor2  gate3612(.a(N11121), .b(N11144), .O(gate3413inter0));
  nand2 gate3613(.a(gate3413inter0), .b(s_14), .O(gate3413inter1));
  and2  gate3614(.a(N11121), .b(N11144), .O(gate3413inter2));
  inv1  gate3615(.a(s_14), .O(gate3413inter3));
  inv1  gate3616(.a(s_15), .O(gate3413inter4));
  nand2 gate3617(.a(gate3413inter4), .b(gate3413inter3), .O(gate3413inter5));
  nor2  gate3618(.a(gate3413inter5), .b(gate3413inter2), .O(gate3413inter6));
  inv1  gate3619(.a(N11144), .O(gate3413inter7));
  inv1  gate3620(.a(N11121), .O(gate3413inter8));
  nand2 gate3621(.a(gate3413inter8), .b(gate3413inter7), .O(gate3413inter9));
  nand2 gate3622(.a(s_15), .b(gate3413inter3), .O(gate3413inter10));
  nor2  gate3623(.a(gate3413inter10), .b(gate3413inter9), .O(gate3413inter11));
  nor2  gate3624(.a(gate3413inter11), .b(gate3413inter6), .O(gate3413inter12));
  nand2 gate3625(.a(gate3413inter12), .b(gate3413inter1), .O(N11177));
nand2 gate3414( .a(N11145), .b(N11123), .O(N11180) );
inv1 gate3415( .a(N11124), .O(N11183) );
nand2 gate3416( .a(N11124), .b(N9468), .O(N11184) );
inv1 gate3417( .a(N11127), .O(N11185) );
nand2 gate3418( .a(N11127), .b(N9508), .O(N11186) );
inv1 gate3419( .a(N11130), .O(N11187) );
nand2 gate3420( .a(N11130), .b(N9509), .O(N11188) );
or4 gate3421( .a(N11152), .b(N11153), .c(N11154), .d(N11155), .O(N11205) );
nand2 gate3422( .a(N8724), .b(N11183), .O(N11210) );
nand2 gate3423( .a(N8790), .b(N11185), .O(N11211) );
nand2 gate3424( .a(N8808), .b(N11187), .O(N11212) );
inv1 gate3425( .a(N11168), .O(N11213) );
nand2 gate3426( .a(N11168), .b(N8260), .O(N11214) );
inv1 gate3427( .a(N11171), .O(N11215) );
nand2 gate3428( .a(N11171), .b(N8261), .O(N11216) );
inv1 gate3429( .a(N11174), .O(N11217) );
nand2 gate3430( .a(N11174), .b(N8296), .O(N11218) );
inv1 gate3431( .a(N11177), .O(N11219) );
nand2 gate3432( .a(N11177), .b(N8297), .O(N11220) );
and3 gate3433( .a(N11159), .b(N9575), .c(N1218), .O(N11222) );
and3 gate3434( .a(N11156), .b(N8927), .c(N1218), .O(N11223) );
and3 gate3435( .a(N11159), .b(N9935), .c(N750), .O(N11224) );
and3 gate3436( .a(N11156), .b(N10132), .c(N750), .O(N11225) );
and3 gate3437( .a(N11165), .b(N9608), .c(N10497), .O(N11226) );
and3 gate3438( .a(N11162), .b(N9001), .c(N10497), .O(N11227) );
and3 gate3439( .a(N11165), .b(N9949), .c(N10301), .O(N11228) );
and3 gate3440( .a(N11162), .b(N10160), .c(N10301), .O(N11229) );
inv1 gate3441( .a(N11180), .O(N11231) );
nand2 gate3442( .a(N11180), .b(N9467), .O(N11232) );
nand2 gate3443( .a(N11210), .b(N11184), .O(N11233) );
nand2 gate3444( .a(N11211), .b(N11186), .O(N11236) );
nand2 gate3445( .a(N11212), .b(N11188), .O(N11239) );
nand2 gate3446( .a(N7459), .b(N11213), .O(N11242) );
nand2 gate3447( .a(N7462), .b(N11215), .O(N11243) );
nand2 gate3448( .a(N7515), .b(N11217), .O(N11244) );
nand2 gate3449( .a(N7518), .b(N11219), .O(N11245) );
inv1 gate3450( .a(N11205), .O(N11246) );
nand2 gate3451( .a(N8708), .b(N11231), .O(N11250) );
or4 gate3452( .a(N11222), .b(N11223), .c(N11224), .d(N11225), .O(N11252) );
or4 gate3453( .a(N11226), .b(N11227), .c(N11228), .d(N11229), .O(N11257) );
nand2 gate3454( .a(N11242), .b(N11214), .O(N11260) );

  xor2  gate4200(.a(N11216), .b(N11243), .O(gate3455inter0));
  nand2 gate4201(.a(gate3455inter0), .b(s_98), .O(gate3455inter1));
  and2  gate4202(.a(N11216), .b(N11243), .O(gate3455inter2));
  inv1  gate4203(.a(s_98), .O(gate3455inter3));
  inv1  gate4204(.a(s_99), .O(gate3455inter4));
  nand2 gate4205(.a(gate3455inter4), .b(gate3455inter3), .O(gate3455inter5));
  nor2  gate4206(.a(gate3455inter5), .b(gate3455inter2), .O(gate3455inter6));
  inv1  gate4207(.a(N11243), .O(gate3455inter7));
  inv1  gate4208(.a(N11216), .O(gate3455inter8));
  nand2 gate4209(.a(gate3455inter8), .b(gate3455inter7), .O(gate3455inter9));
  nand2 gate4210(.a(s_99), .b(gate3455inter3), .O(gate3455inter10));
  nor2  gate4211(.a(gate3455inter10), .b(gate3455inter9), .O(gate3455inter11));
  nor2  gate4212(.a(gate3455inter11), .b(gate3455inter6), .O(gate3455inter12));
  nand2 gate4213(.a(gate3455inter12), .b(gate3455inter1), .O(N11261));
nand2 gate3456( .a(N11244), .b(N11218), .O(N11262) );
nand2 gate3457( .a(N11245), .b(N11220), .O(N11263) );
inv1 gate3458( .a(N11233), .O(N11264) );
nand2 gate3459( .a(N11233), .b(N9322), .O(N11265) );
inv1 gate3460( .a(N11236), .O(N11267) );

  xor2  gate4438(.a(N9383), .b(N11236), .O(gate3461inter0));
  nand2 gate4439(.a(gate3461inter0), .b(s_132), .O(gate3461inter1));
  and2  gate4440(.a(N9383), .b(N11236), .O(gate3461inter2));
  inv1  gate4441(.a(s_132), .O(gate3461inter3));
  inv1  gate4442(.a(s_133), .O(gate3461inter4));
  nand2 gate4443(.a(gate3461inter4), .b(gate3461inter3), .O(gate3461inter5));
  nor2  gate4444(.a(gate3461inter5), .b(gate3461inter2), .O(gate3461inter6));
  inv1  gate4445(.a(N11236), .O(gate3461inter7));
  inv1  gate4446(.a(N9383), .O(gate3461inter8));
  nand2 gate4447(.a(gate3461inter8), .b(gate3461inter7), .O(gate3461inter9));
  nand2 gate4448(.a(s_133), .b(gate3461inter3), .O(gate3461inter10));
  nor2  gate4449(.a(gate3461inter10), .b(gate3461inter9), .O(gate3461inter11));
  nor2  gate4450(.a(gate3461inter11), .b(gate3461inter6), .O(gate3461inter12));
  nand2 gate4451(.a(gate3461inter12), .b(gate3461inter1), .O(N11268));
inv1 gate3462( .a(N11239), .O(N11269) );
nand2 gate3463( .a(N11239), .b(N9384), .O(N11270) );

  xor2  gate3906(.a(N11232), .b(N11250), .O(gate3464inter0));
  nand2 gate3907(.a(gate3464inter0), .b(s_56), .O(gate3464inter1));
  and2  gate3908(.a(N11232), .b(N11250), .O(gate3464inter2));
  inv1  gate3909(.a(s_56), .O(gate3464inter3));
  inv1  gate3910(.a(s_57), .O(gate3464inter4));
  nand2 gate3911(.a(gate3464inter4), .b(gate3464inter3), .O(gate3464inter5));
  nor2  gate3912(.a(gate3464inter5), .b(gate3464inter2), .O(gate3464inter6));
  inv1  gate3913(.a(N11250), .O(gate3464inter7));
  inv1  gate3914(.a(N11232), .O(gate3464inter8));
  nand2 gate3915(.a(gate3464inter8), .b(gate3464inter7), .O(gate3464inter9));
  nand2 gate3916(.a(s_57), .b(gate3464inter3), .O(gate3464inter10));
  nor2  gate3917(.a(gate3464inter10), .b(gate3464inter9), .O(gate3464inter11));
  nor2  gate3918(.a(gate3464inter11), .b(gate3464inter6), .O(gate3464inter12));
  nand2 gate3919(.a(gate3464inter12), .b(gate3464inter1), .O(N11272));
inv1 gate3465( .a(N11261), .O(N11277) );
and2 gate3466( .a(N10273), .b(N11260), .O(N11278) );
inv1 gate3467( .a(N11263), .O(N11279) );
and2 gate3468( .a(N10119), .b(N11262), .O(N11280) );
nand2 gate3469( .a(N8714), .b(N11264), .O(N11282) );
inv1 gate3470( .a(N11252), .O(N11283) );
nand2 gate3471( .a(N8793), .b(N11267), .O(N11284) );
nand2 gate3472( .a(N8796), .b(N11269), .O(N11285) );
inv1 gate3473( .a(N11257), .O(N11286) );
and2 gate3474( .a(N11277), .b(N10479), .O(N11288) );
and2 gate3475( .a(N11279), .b(N10283), .O(N11289) );
inv1 gate3476( .a(N11272), .O(N11290) );
nand2 gate3477( .a(N11272), .b(N9321), .O(N11291) );
nand2 gate3478( .a(N11282), .b(N11265), .O(N11292) );
nand2 gate3479( .a(N11284), .b(N11268), .O(N11293) );
nand2 gate3480( .a(N11285), .b(N11270), .O(N11294) );
nand2 gate3481( .a(N8711), .b(N11290), .O(N11295) );
inv1 gate3482( .a(N11292), .O(N11296) );
inv1 gate3483( .a(N11294), .O(N11297) );
and2 gate3484( .a(N10301), .b(N11293), .O(N11298) );
or2 gate3485( .a(N11288), .b(N11278), .O(N11299) );
or2 gate3486( .a(N11289), .b(N11280), .O(N11302) );
nand2 gate3487( .a(N11295), .b(N11291), .O(N11307) );
and2 gate3488( .a(N11296), .b(N1218), .O(N11308) );
and2 gate3489( .a(N11297), .b(N10497), .O(N11309) );
nand2 gate3490( .a(N11302), .b(N11246), .O(N11312) );
nand2 gate3491( .a(N11299), .b(N10836), .O(N11313) );
inv1 gate3492( .a(N11299), .O(N11314) );
inv1 gate3493( .a(N11302), .O(N11315) );
and2 gate3494( .a(N750), .b(N11307), .O(N11316) );
or2 gate3495( .a(N11309), .b(N11298), .O(N11317) );
nand2 gate3496( .a(N11205), .b(N11315), .O(N11320) );

  xor2  gate3892(.a(N11314), .b(N10739), .O(gate3497inter0));
  nand2 gate3893(.a(gate3497inter0), .b(s_54), .O(gate3497inter1));
  and2  gate3894(.a(N11314), .b(N10739), .O(gate3497inter2));
  inv1  gate3895(.a(s_54), .O(gate3497inter3));
  inv1  gate3896(.a(s_55), .O(gate3497inter4));
  nand2 gate3897(.a(gate3497inter4), .b(gate3497inter3), .O(gate3497inter5));
  nor2  gate3898(.a(gate3497inter5), .b(gate3497inter2), .O(gate3497inter6));
  inv1  gate3899(.a(N10739), .O(gate3497inter7));
  inv1  gate3900(.a(N11314), .O(gate3497inter8));
  nand2 gate3901(.a(gate3497inter8), .b(gate3497inter7), .O(gate3497inter9));
  nand2 gate3902(.a(s_55), .b(gate3497inter3), .O(gate3497inter10));
  nor2  gate3903(.a(gate3497inter10), .b(gate3497inter9), .O(gate3497inter11));
  nor2  gate3904(.a(gate3497inter11), .b(gate3497inter6), .O(gate3497inter12));
  nand2 gate3905(.a(gate3497inter12), .b(gate3497inter1), .O(N11321));
or2 gate3498( .a(N11308), .b(N11316), .O(N11323) );
nand2 gate3499( .a(N11312), .b(N11320), .O(N11327) );

  xor2  gate5180(.a(N11321), .b(N11313), .O(gate3500inter0));
  nand2 gate5181(.a(gate3500inter0), .b(s_238), .O(gate3500inter1));
  and2  gate5182(.a(N11321), .b(N11313), .O(gate3500inter2));
  inv1  gate5183(.a(s_238), .O(gate3500inter3));
  inv1  gate5184(.a(s_239), .O(gate3500inter4));
  nand2 gate5185(.a(gate3500inter4), .b(gate3500inter3), .O(gate3500inter5));
  nor2  gate5186(.a(gate3500inter5), .b(gate3500inter2), .O(gate3500inter6));
  inv1  gate5187(.a(N11313), .O(gate3500inter7));
  inv1  gate5188(.a(N11321), .O(gate3500inter8));
  nand2 gate5189(.a(gate3500inter8), .b(gate3500inter7), .O(gate3500inter9));
  nand2 gate5190(.a(s_239), .b(gate3500inter3), .O(gate3500inter10));
  nor2  gate5191(.a(gate3500inter10), .b(gate3500inter9), .O(gate3500inter11));
  nor2  gate5192(.a(gate3500inter11), .b(gate3500inter6), .O(gate3500inter12));
  nand2 gate5193(.a(gate3500inter12), .b(gate3500inter1), .O(N11328));
nand2 gate3501( .a(N11317), .b(N11286), .O(N11329) );
inv1 gate3502( .a(N11317), .O(N11331) );
inv1 gate3503( .a(N11327), .O(N11333) );
inv1 gate3504( .a(N11328), .O(N11334) );
nand2 gate3505( .a(N11257), .b(N11331), .O(N11335) );
nand2 gate3506( .a(N11323), .b(N11283), .O(N11336) );
inv1 gate3507( .a(N11323), .O(N11337) );
nand2 gate3508( .a(N11329), .b(N11335), .O(N11338) );
nand2 gate3509( .a(N11252), .b(N11337), .O(N11339) );
inv1 gate3510( .a(N11338), .O(N11340) );
nand2 gate3511( .a(N11336), .b(N11339), .O(N11341) );
inv1 gate3512( .a(N11341), .O(N11342) );
buf1 gate3513( .a(N241_I), .O(N241_O) );

endmodule