module c1908 (N1,N4,N7,N10,N13,N16,N19,N22,N25,N28,
              N31,N34,N37,N40,N43,N46,N49,N53,N56,N60,
              N63,N66,N69,N72,N76,N79,N82,N85,N88,N91,
              N94,N99,N104,N2753,N2754,N2755,N2756,N2762,N2767,N2768,
              N2779,N2780,N2781,N2782,N2783,N2784,N2785,N2786,N2787,N2811,
              N2886,N2887,N2888,N2889,N2890,N2891,N2892,N2899);
input N1,N4,N7,N10,N13,N16,N19,N22,N25,N28,
      N31,N34,N37,N40,N43,N46,N49,N53,N56,N60,
      N63,N66,N69,N72,N76,N79,N82,N85,N88,N91,
      N94,N99,N104;
  input s_0, s_1, s_2, s_3, s_4, s_5, s_6, s_7, s_8, s_9, s_10, s_11, s_12, s_13, s_14, s_15, s_16, s_17, s_18, s_19, s_20, s_21, s_22, s_23, s_24, s_25, s_26, s_27, s_28, s_29, s_30, s_31, s_32, s_33, s_34, s_35, s_36, s_37, s_38, s_39, s_40, s_41, s_42, s_43, s_44, s_45, s_46, s_47, s_48, s_49, s_50, s_51, s_52, s_53, s_54, s_55, s_56, s_57, s_58, s_59, s_60, s_61, s_62, s_63, s_64, s_65, s_66, s_67, s_68, s_69, s_70, s_71, s_72, s_73, s_74, s_75, s_76, s_77, s_78, s_79, s_80, s_81, s_82, s_83, s_84, s_85, s_86, s_87, s_88, s_89, s_90, s_91, s_92, s_93, s_94, s_95, s_96, s_97, s_98, s_99, s_100, s_101, s_102, s_103, s_104, s_105, s_106, s_107, s_108, s_109, s_110, s_111, s_112, s_113, s_114, s_115, s_116, s_117, s_118, s_119, s_120, s_121, s_122, s_123, s_124, s_125, s_126, s_127, s_128, s_129, s_130, s_131, s_132, s_133, s_134, s_135, s_136, s_137, s_138, s_139, s_140, s_141, s_142, s_143, s_144, s_145, s_146, s_147, s_148, s_149, s_150, s_151, s_152, s_153, s_154, s_155, s_156, s_157, s_158, s_159, s_160, s_161, s_162, s_163, s_164, s_165, s_166, s_167, s_168, s_169, s_170, s_171, s_172, s_173, s_174, s_175, s_176, s_177, s_178, s_179, s_180, s_181;
output N2753,N2754,N2755,N2756,N2762,N2767,N2768,N2779,N2780,N2781,
       N2782,N2783,N2784,N2785,N2786,N2787,N2811,N2886,N2887,N2888,
       N2889,N2890,N2891,N2892,N2899;
wire N190,N194,N197,N201,N206,N209,N212,N216,N220,N225,
     N229,N232,N235,N239,N243,N247,N251,N252,N253,N256,
     N257,N260,N263,N266,N269,N272,N275,N276,N277,N280,
     N283,N290,N297,N300,N303,N306,N313,N316,N319,N326,
     N331,N338,N343,N346,N349,N352,N355,N358,N361,N364,
     N367,N370,N373,N376,N379,N382,N385,N388,N534,N535,
     N536,N537,N538,N539,N540,N541,N542,N543,N544,N545,
     N546,N547,N548,N549,N550,N551,N552,N553,N554,N555,
     N556,N559,N562,N565,N568,N571,N574,N577,N580,N583,
     N586,N589,N592,N595,N598,N601,N602,N603,N608,N612,
     N616,N619,N622,N625,N628,N631,N634,N637,N640,N643,
     N646,N649,N652,N655,N658,N661,N664,N667,N670,N673,
     N676,N679,N682,N685,N688,N691,N694,N697,N700,N703,
     N706,N709,N712,N715,N718,N721,N724,N727,N730,N733,
     N736,N739,N742,N745,N748,N751,N886,N887,N888,N889,
     N890,N891,N892,N893,N894,N895,N896,N897,N898,N899,
     N903,N907,N910,N913,N914,N915,N916,N917,N918,N919,
     N920,N921,N922,N923,N926,N935,N938,N939,N942,N943,
     N946,N947,N950,N951,N954,N955,N958,N959,N962,N965,
     N968,N969,N972,N973,N976,N977,N980,N981,N984,N985,
     N988,N989,N990,N991,N992,N993,N994,N997,N998,N1001,
     N1002,N1003,N1004,N1005,N1006,N1007,N1008,N1009,N1010,N1013,
     N1016,N1019,N1022,N1025,N1028,N1031,N1034,N1037,N1040,N1043,
     N1046,N1049,N1054,N1055,N1063,N1064,N1067,N1068,N1119,N1120,
     N1121,N1122,N1128,N1129,N1130,N1131,N1132,N1133,N1148,N1149,
     N1150,N1151,N1152,N1153,N1154,N1155,N1156,N1157,N1158,N1159,
     N1160,N1161,N1162,N1163,N1164,N1167,N1168,N1171,N1188,N1205,
     N1206,N1207,N1208,N1209,N1210,N1211,N1212,N1213,N1214,N1215,
     N1216,N1217,N1218,N1219,N1220,N1221,N1222,N1223,N1224,N1225,
     N1226,N1227,N1228,N1229,N1230,N1231,N1232,N1235,N1238,N1239,
     N1240,N1241,N1242,N1243,N1246,N1249,N1252,N1255,N1258,N1261,
     N1264,N1267,N1309,N1310,N1311,N1312,N1313,N1314,N1315,N1316,
     N1317,N1318,N1319,N1322,N1327,N1328,N1334,N1344,N1345,N1346,
     N1348,N1349,N1350,N1351,N1352,N1355,N1358,N1361,N1364,N1367,
     N1370,N1373,N1376,N1379,N1383,N1386,N1387,N1388,N1389,N1390,
     N1393,N1396,N1397,N1398,N1399,N1409,N1412,N1413,N1416,N1419,
     N1433,N1434,N1438,N1439,N1440,N1443,N1444,N1445,N1446,N1447,
     N1448,N1451,N1452,N1453,N1454,N1455,N1456,N1457,N1458,N1459,
     N1460,N1461,N1462,N1463,N1464,N1468,N1469,N1470,N1471,N1472,
     N1475,N1476,N1478,N1481,N1484,N1487,N1488,N1489,N1490,N1491,
     N1492,N1493,N1494,N1495,N1496,N1498,N1499,N1500,N1501,N1504,
     N1510,N1513,N1514,N1517,N1520,N1521,N1522,N1526,N1527,N1528,
     N1529,N1530,N1531,N1532,N1534,N1537,N1540,N1546,N1554,N1557,
     N1561,N1567,N1568,N1569,N1571,N1576,N1588,N1591,N1593,N1594,
     N1595,N1596,N1600,N1603,N1606,N1609,N1612,N1615,N1620,N1623,
     N1635,N1636,N1638,N1639,N1640,N1643,N1647,N1651,N1658,N1661,
     N1664,N1671,N1672,N1675,N1677,N1678,N1679,N1680,N1681,N1682,
     N1683,N1685,N1688,N1697,N1701,N1706,N1707,N1708,N1709,N1710,
     N1711,N1712,N1713,N1714,N1717,N1720,N1721,N1723,N1727,N1728,
     N1730,N1731,N1734,N1740,N1741,N1742,N1746,N1747,N1748,N1751,
     N1759,N1761,N1762,N1763,N1764,N1768,N1769,N1772,N1773,N1774,
     N1777,N1783,N1784,N1785,N1786,N1787,N1788,N1791,N1792,N1795,
     N1796,N1798,N1801,N1802,N1807,N1808,N1809,N1810,N1812,N1815,
     N1818,N1821,N1822,N1823,N1824,N1825,N1826,N1827,N1830,N1837,
     N1838,N1841,N1848,N1849,N1850,N1852,N1855,N1856,N1857,N1858,
     N1864,N1865,N1866,N1869,N1872,N1875,N1878,N1879,N1882,N1883,
     N1884,N1885,N1889,N1895,N1896,N1897,N1898,N1902,N1910,N1911,
     N1912,N1913,N1915,N1919,N1920,N1921,N1922,N1923,N1924,N1927,
     N1930,N1933,N1936,N1937,N1938,N1941,N1942,N1944,N1947,N1950,
     N1953,N1958,N1961,N1965,N1968,N1975,N1976,N1977,N1978,N1979,
     N1980,N1985,N1987,N1999,N2000,N2002,N2003,N2004,N2005,N2006,
     N2007,N2008,N2009,N2012,N2013,N2014,N2015,N2016,N2018,N2019,
     N2020,N2021,N2022,N2023,N2024,N2025,N2026,N2027,N2030,N2033,
     N2036,N2037,N2038,N2039,N2040,N2041,N2042,N2047,N2052,N2055,
     N2060,N2061,N2062,N2067,N2068,N2071,N2076,N2077,N2078,N2081,
     N2086,N2089,N2104,N2119,N2129,N2143,N2148,N2151,N2196,N2199,
     N2202,N2205,N2214,N2215,N2216,N2217,N2222,N2223,N2224,N2225,
     N2226,N2227,N2228,N2229,N2230,N2231,N2232,N2233,N2234,N2235,
     N2236,N2237,N2240,N2241,N2244,N2245,N2250,N2253,N2256,N2257,
     N2260,N2263,N2266,N2269,N2272,N2279,N2286,N2297,N2315,N2326,
     N2340,N2353,N2361,N2375,N2384,N2385,N2386,N2426,N2427,N2537,
     N2540,N2543,N2546,N2549,N2552,N2555,N2558,N2561,N2564,N2567,
     N2570,N2573,N2576,N2594,N2597,N2600,N2603,N2606,N2611,N2614,
     N2617,N2620,N2627,N2628,N2629,N2630,N2631,N2632,N2633,N2634,
     N2639,N2642,N2645,N2648,N2651,N2655,N2658,N2661,N2664,N2669,
     N2670,N2671,N2672,N2673,N2674,N2675,N2676,N2682,N2683,N2688,
     N2689,N2690,N2691,N2710,N2720,N2721,N2722,N2723,N2724,N2725,
     N2726,N2727,N2728,N2729,N2730,N2731,N2732,N2733,N2734,N2735,
     N2736,N2737,N2738,N2739,N2740,N2741,N2742,N2743,N2744,N2745,
     N2746,N2747,N2750,N2757,N2758,N2759,N2760,N2761,N2763,N2764,
     N2765,N2766,N2773,N2776,N2788,N2789,N2800,N2807,N2808,N2809,
     N2810,N2812,N2815,N2818,N2821,N2824,N2827,N2828,N2829,N2843,
     N2846,N2850,N2851,N2852,N2853,N2854,N2857,N2858,N2859,N2860,
     N2861,N2862,N2863,N2866,N2867,N2868,N2869,N2870,N2871,N2872,
     N2873,N2874,N2875,N2876,N2877,N2878,N2879,N2880,N2881,N2882,
     N2883,N2895,N2896,N2897,N2898, gate319inter0, gate319inter1, gate319inter2, gate319inter3, gate319inter4, gate319inter5, gate319inter6, gate319inter7, gate319inter8, gate319inter9, gate319inter10, gate319inter11, gate319inter12, gate839inter0, gate839inter1, gate839inter2, gate839inter3, gate839inter4, gate839inter5, gate839inter6, gate839inter7, gate839inter8, gate839inter9, gate839inter10, gate839inter11, gate839inter12, gate522inter0, gate522inter1, gate522inter2, gate522inter3, gate522inter4, gate522inter5, gate522inter6, gate522inter7, gate522inter8, gate522inter9, gate522inter10, gate522inter11, gate522inter12, gate281inter0, gate281inter1, gate281inter2, gate281inter3, gate281inter4, gate281inter5, gate281inter6, gate281inter7, gate281inter8, gate281inter9, gate281inter10, gate281inter11, gate281inter12, gate527inter0, gate527inter1, gate527inter2, gate527inter3, gate527inter4, gate527inter5, gate527inter6, gate527inter7, gate527inter8, gate527inter9, gate527inter10, gate527inter11, gate527inter12, gate243inter0, gate243inter1, gate243inter2, gate243inter3, gate243inter4, gate243inter5, gate243inter6, gate243inter7, gate243inter8, gate243inter9, gate243inter10, gate243inter11, gate243inter12, gate247inter0, gate247inter1, gate247inter2, gate247inter3, gate247inter4, gate247inter5, gate247inter6, gate247inter7, gate247inter8, gate247inter9, gate247inter10, gate247inter11, gate247inter12, gate279inter0, gate279inter1, gate279inter2, gate279inter3, gate279inter4, gate279inter5, gate279inter6, gate279inter7, gate279inter8, gate279inter9, gate279inter10, gate279inter11, gate279inter12, gate814inter0, gate814inter1, gate814inter2, gate814inter3, gate814inter4, gate814inter5, gate814inter6, gate814inter7, gate814inter8, gate814inter9, gate814inter10, gate814inter11, gate814inter12, gate613inter0, gate613inter1, gate613inter2, gate613inter3, gate613inter4, gate613inter5, gate613inter6, gate613inter7, gate613inter8, gate613inter9, gate613inter10, gate613inter11, gate613inter12, gate570inter0, gate570inter1, gate570inter2, gate570inter3, gate570inter4, gate570inter5, gate570inter6, gate570inter7, gate570inter8, gate570inter9, gate570inter10, gate570inter11, gate570inter12, gate634inter0, gate634inter1, gate634inter2, gate634inter3, gate634inter4, gate634inter5, gate634inter6, gate634inter7, gate634inter8, gate634inter9, gate634inter10, gate634inter11, gate634inter12, gate798inter0, gate798inter1, gate798inter2, gate798inter3, gate798inter4, gate798inter5, gate798inter6, gate798inter7, gate798inter8, gate798inter9, gate798inter10, gate798inter11, gate798inter12, gate248inter0, gate248inter1, gate248inter2, gate248inter3, gate248inter4, gate248inter5, gate248inter6, gate248inter7, gate248inter8, gate248inter9, gate248inter10, gate248inter11, gate248inter12, gate840inter0, gate840inter1, gate840inter2, gate840inter3, gate840inter4, gate840inter5, gate840inter6, gate840inter7, gate840inter8, gate840inter9, gate840inter10, gate840inter11, gate840inter12, gate681inter0, gate681inter1, gate681inter2, gate681inter3, gate681inter4, gate681inter5, gate681inter6, gate681inter7, gate681inter8, gate681inter9, gate681inter10, gate681inter11, gate681inter12, gate271inter0, gate271inter1, gate271inter2, gate271inter3, gate271inter4, gate271inter5, gate271inter6, gate271inter7, gate271inter8, gate271inter9, gate271inter10, gate271inter11, gate271inter12, gate856inter0, gate856inter1, gate856inter2, gate856inter3, gate856inter4, gate856inter5, gate856inter6, gate856inter7, gate856inter8, gate856inter9, gate856inter10, gate856inter11, gate856inter12, gate494inter0, gate494inter1, gate494inter2, gate494inter3, gate494inter4, gate494inter5, gate494inter6, gate494inter7, gate494inter8, gate494inter9, gate494inter10, gate494inter11, gate494inter12, gate312inter0, gate312inter1, gate312inter2, gate312inter3, gate312inter4, gate312inter5, gate312inter6, gate312inter7, gate312inter8, gate312inter9, gate312inter10, gate312inter11, gate312inter12, gate511inter0, gate511inter1, gate511inter2, gate511inter3, gate511inter4, gate511inter5, gate511inter6, gate511inter7, gate511inter8, gate511inter9, gate511inter10, gate511inter11, gate511inter12, gate99inter0, gate99inter1, gate99inter2, gate99inter3, gate99inter4, gate99inter5, gate99inter6, gate99inter7, gate99inter8, gate99inter9, gate99inter10, gate99inter11, gate99inter12, gate453inter0, gate453inter1, gate453inter2, gate453inter3, gate453inter4, gate453inter5, gate453inter6, gate453inter7, gate453inter8, gate453inter9, gate453inter10, gate453inter11, gate453inter12, gate261inter0, gate261inter1, gate261inter2, gate261inter3, gate261inter4, gate261inter5, gate261inter6, gate261inter7, gate261inter8, gate261inter9, gate261inter10, gate261inter11, gate261inter12, gate402inter0, gate402inter1, gate402inter2, gate402inter3, gate402inter4, gate402inter5, gate402inter6, gate402inter7, gate402inter8, gate402inter9, gate402inter10, gate402inter11, gate402inter12, gate385inter0, gate385inter1, gate385inter2, gate385inter3, gate385inter4, gate385inter5, gate385inter6, gate385inter7, gate385inter8, gate385inter9, gate385inter10, gate385inter11, gate385inter12, gate242inter0, gate242inter1, gate242inter2, gate242inter3, gate242inter4, gate242inter5, gate242inter6, gate242inter7, gate242inter8, gate242inter9, gate242inter10, gate242inter11, gate242inter12, gate800inter0, gate800inter1, gate800inter2, gate800inter3, gate800inter4, gate800inter5, gate800inter6, gate800inter7, gate800inter8, gate800inter9, gate800inter10, gate800inter11, gate800inter12, gate478inter0, gate478inter1, gate478inter2, gate478inter3, gate478inter4, gate478inter5, gate478inter6, gate478inter7, gate478inter8, gate478inter9, gate478inter10, gate478inter11, gate478inter12, gate854inter0, gate854inter1, gate854inter2, gate854inter3, gate854inter4, gate854inter5, gate854inter6, gate854inter7, gate854inter8, gate854inter9, gate854inter10, gate854inter11, gate854inter12, gate754inter0, gate754inter1, gate754inter2, gate754inter3, gate754inter4, gate754inter5, gate754inter6, gate754inter7, gate754inter8, gate754inter9, gate754inter10, gate754inter11, gate754inter12, gate370inter0, gate370inter1, gate370inter2, gate370inter3, gate370inter4, gate370inter5, gate370inter6, gate370inter7, gate370inter8, gate370inter9, gate370inter10, gate370inter11, gate370inter12, gate336inter0, gate336inter1, gate336inter2, gate336inter3, gate336inter4, gate336inter5, gate336inter6, gate336inter7, gate336inter8, gate336inter9, gate336inter10, gate336inter11, gate336inter12, gate315inter0, gate315inter1, gate315inter2, gate315inter3, gate315inter4, gate315inter5, gate315inter6, gate315inter7, gate315inter8, gate315inter9, gate315inter10, gate315inter11, gate315inter12, gate404inter0, gate404inter1, gate404inter2, gate404inter3, gate404inter4, gate404inter5, gate404inter6, gate404inter7, gate404inter8, gate404inter9, gate404inter10, gate404inter11, gate404inter12, gate342inter0, gate342inter1, gate342inter2, gate342inter3, gate342inter4, gate342inter5, gate342inter6, gate342inter7, gate342inter8, gate342inter9, gate342inter10, gate342inter11, gate342inter12, gate752inter0, gate752inter1, gate752inter2, gate752inter3, gate752inter4, gate752inter5, gate752inter6, gate752inter7, gate752inter8, gate752inter9, gate752inter10, gate752inter11, gate752inter12, gate796inter0, gate796inter1, gate796inter2, gate796inter3, gate796inter4, gate796inter5, gate796inter6, gate796inter7, gate796inter8, gate796inter9, gate796inter10, gate796inter11, gate796inter12, gate621inter0, gate621inter1, gate621inter2, gate621inter3, gate621inter4, gate621inter5, gate621inter6, gate621inter7, gate621inter8, gate621inter9, gate621inter10, gate621inter11, gate621inter12, gate286inter0, gate286inter1, gate286inter2, gate286inter3, gate286inter4, gate286inter5, gate286inter6, gate286inter7, gate286inter8, gate286inter9, gate286inter10, gate286inter11, gate286inter12, gate353inter0, gate353inter1, gate353inter2, gate353inter3, gate353inter4, gate353inter5, gate353inter6, gate353inter7, gate353inter8, gate353inter9, gate353inter10, gate353inter11, gate353inter12, gate488inter0, gate488inter1, gate488inter2, gate488inter3, gate488inter4, gate488inter5, gate488inter6, gate488inter7, gate488inter8, gate488inter9, gate488inter10, gate488inter11, gate488inter12, gate878inter0, gate878inter1, gate878inter2, gate878inter3, gate878inter4, gate878inter5, gate878inter6, gate878inter7, gate878inter8, gate878inter9, gate878inter10, gate878inter11, gate878inter12, gate596inter0, gate596inter1, gate596inter2, gate596inter3, gate596inter4, gate596inter5, gate596inter6, gate596inter7, gate596inter8, gate596inter9, gate596inter10, gate596inter11, gate596inter12, gate524inter0, gate524inter1, gate524inter2, gate524inter3, gate524inter4, gate524inter5, gate524inter6, gate524inter7, gate524inter8, gate524inter9, gate524inter10, gate524inter11, gate524inter12, gate300inter0, gate300inter1, gate300inter2, gate300inter3, gate300inter4, gate300inter5, gate300inter6, gate300inter7, gate300inter8, gate300inter9, gate300inter10, gate300inter11, gate300inter12, gate17inter0, gate17inter1, gate17inter2, gate17inter3, gate17inter4, gate17inter5, gate17inter6, gate17inter7, gate17inter8, gate17inter9, gate17inter10, gate17inter11, gate17inter12, gate756inter0, gate756inter1, gate756inter2, gate756inter3, gate756inter4, gate756inter5, gate756inter6, gate756inter7, gate756inter8, gate756inter9, gate756inter10, gate756inter11, gate756inter12, gate818inter0, gate818inter1, gate818inter2, gate818inter3, gate818inter4, gate818inter5, gate818inter6, gate818inter7, gate818inter8, gate818inter9, gate818inter10, gate818inter11, gate818inter12, gate618inter0, gate618inter1, gate618inter2, gate618inter3, gate618inter4, gate618inter5, gate618inter6, gate618inter7, gate618inter8, gate618inter9, gate618inter10, gate618inter11, gate618inter12, gate628inter0, gate628inter1, gate628inter2, gate628inter3, gate628inter4, gate628inter5, gate628inter6, gate628inter7, gate628inter8, gate628inter9, gate628inter10, gate628inter11, gate628inter12, gate773inter0, gate773inter1, gate773inter2, gate773inter3, gate773inter4, gate773inter5, gate773inter6, gate773inter7, gate773inter8, gate773inter9, gate773inter10, gate773inter11, gate773inter12, gate235inter0, gate235inter1, gate235inter2, gate235inter3, gate235inter4, gate235inter5, gate235inter6, gate235inter7, gate235inter8, gate235inter9, gate235inter10, gate235inter11, gate235inter12, gate390inter0, gate390inter1, gate390inter2, gate390inter3, gate390inter4, gate390inter5, gate390inter6, gate390inter7, gate390inter8, gate390inter9, gate390inter10, gate390inter11, gate390inter12, gate826inter0, gate826inter1, gate826inter2, gate826inter3, gate826inter4, gate826inter5, gate826inter6, gate826inter7, gate826inter8, gate826inter9, gate826inter10, gate826inter11, gate826inter12, gate631inter0, gate631inter1, gate631inter2, gate631inter3, gate631inter4, gate631inter5, gate631inter6, gate631inter7, gate631inter8, gate631inter9, gate631inter10, gate631inter11, gate631inter12, gate245inter0, gate245inter1, gate245inter2, gate245inter3, gate245inter4, gate245inter5, gate245inter6, gate245inter7, gate245inter8, gate245inter9, gate245inter10, gate245inter11, gate245inter12, gate427inter0, gate427inter1, gate427inter2, gate427inter3, gate427inter4, gate427inter5, gate427inter6, gate427inter7, gate427inter8, gate427inter9, gate427inter10, gate427inter11, gate427inter12, gate518inter0, gate518inter1, gate518inter2, gate518inter3, gate518inter4, gate518inter5, gate518inter6, gate518inter7, gate518inter8, gate518inter9, gate518inter10, gate518inter11, gate518inter12, gate812inter0, gate812inter1, gate812inter2, gate812inter3, gate812inter4, gate812inter5, gate812inter6, gate812inter7, gate812inter8, gate812inter9, gate812inter10, gate812inter11, gate812inter12, gate393inter0, gate393inter1, gate393inter2, gate393inter3, gate393inter4, gate393inter5, gate393inter6, gate393inter7, gate393inter8, gate393inter9, gate393inter10, gate393inter11, gate393inter12, gate876inter0, gate876inter1, gate876inter2, gate876inter3, gate876inter4, gate876inter5, gate876inter6, gate876inter7, gate876inter8, gate876inter9, gate876inter10, gate876inter11, gate876inter12, gate607inter0, gate607inter1, gate607inter2, gate607inter3, gate607inter4, gate607inter5, gate607inter6, gate607inter7, gate607inter8, gate607inter9, gate607inter10, gate607inter11, gate607inter12, gate505inter0, gate505inter1, gate505inter2, gate505inter3, gate505inter4, gate505inter5, gate505inter6, gate505inter7, gate505inter8, gate505inter9, gate505inter10, gate505inter11, gate505inter12, gate415inter0, gate415inter1, gate415inter2, gate415inter3, gate415inter4, gate415inter5, gate415inter6, gate415inter7, gate415inter8, gate415inter9, gate415inter10, gate415inter11, gate415inter12, gate78inter0, gate78inter1, gate78inter2, gate78inter3, gate78inter4, gate78inter5, gate78inter6, gate78inter7, gate78inter8, gate78inter9, gate78inter10, gate78inter11, gate78inter12, gate529inter0, gate529inter1, gate529inter2, gate529inter3, gate529inter4, gate529inter5, gate529inter6, gate529inter7, gate529inter8, gate529inter9, gate529inter10, gate529inter11, gate529inter12, gate582inter0, gate582inter1, gate582inter2, gate582inter3, gate582inter4, gate582inter5, gate582inter6, gate582inter7, gate582inter8, gate582inter9, gate582inter10, gate582inter11, gate582inter12, gate79inter0, gate79inter1, gate79inter2, gate79inter3, gate79inter4, gate79inter5, gate79inter6, gate79inter7, gate79inter8, gate79inter9, gate79inter10, gate79inter11, gate79inter12, gate760inter0, gate760inter1, gate760inter2, gate760inter3, gate760inter4, gate760inter5, gate760inter6, gate760inter7, gate760inter8, gate760inter9, gate760inter10, gate760inter11, gate760inter12, gate676inter0, gate676inter1, gate676inter2, gate676inter3, gate676inter4, gate676inter5, gate676inter6, gate676inter7, gate676inter8, gate676inter9, gate676inter10, gate676inter11, gate676inter12, gate540inter0, gate540inter1, gate540inter2, gate540inter3, gate540inter4, gate540inter5, gate540inter6, gate540inter7, gate540inter8, gate540inter9, gate540inter10, gate540inter11, gate540inter12, gate852inter0, gate852inter1, gate852inter2, gate852inter3, gate852inter4, gate852inter5, gate852inter6, gate852inter7, gate852inter8, gate852inter9, gate852inter10, gate852inter11, gate852inter12, gate864inter0, gate864inter1, gate864inter2, gate864inter3, gate864inter4, gate864inter5, gate864inter6, gate864inter7, gate864inter8, gate864inter9, gate864inter10, gate864inter11, gate864inter12, gate344inter0, gate344inter1, gate344inter2, gate344inter3, gate344inter4, gate344inter5, gate344inter6, gate344inter7, gate344inter8, gate344inter9, gate344inter10, gate344inter11, gate344inter12, gate236inter0, gate236inter1, gate236inter2, gate236inter3, gate236inter4, gate236inter5, gate236inter6, gate236inter7, gate236inter8, gate236inter9, gate236inter10, gate236inter11, gate236inter12, gate640inter0, gate640inter1, gate640inter2, gate640inter3, gate640inter4, gate640inter5, gate640inter6, gate640inter7, gate640inter8, gate640inter9, gate640inter10, gate640inter11, gate640inter12, gate547inter0, gate547inter1, gate547inter2, gate547inter3, gate547inter4, gate547inter5, gate547inter6, gate547inter7, gate547inter8, gate547inter9, gate547inter10, gate547inter11, gate547inter12, gate806inter0, gate806inter1, gate806inter2, gate806inter3, gate806inter4, gate806inter5, gate806inter6, gate806inter7, gate806inter8, gate806inter9, gate806inter10, gate806inter11, gate806inter12, gate801inter0, gate801inter1, gate801inter2, gate801inter3, gate801inter4, gate801inter5, gate801inter6, gate801inter7, gate801inter8, gate801inter9, gate801inter10, gate801inter11, gate801inter12, gate537inter0, gate537inter1, gate537inter2, gate537inter3, gate537inter4, gate537inter5, gate537inter6, gate537inter7, gate537inter8, gate537inter9, gate537inter10, gate537inter11, gate537inter12, gate269inter0, gate269inter1, gate269inter2, gate269inter3, gate269inter4, gate269inter5, gate269inter6, gate269inter7, gate269inter8, gate269inter9, gate269inter10, gate269inter11, gate269inter12, gate347inter0, gate347inter1, gate347inter2, gate347inter3, gate347inter4, gate347inter5, gate347inter6, gate347inter7, gate347inter8, gate347inter9, gate347inter10, gate347inter11, gate347inter12, gate364inter0, gate364inter1, gate364inter2, gate364inter3, gate364inter4, gate364inter5, gate364inter6, gate364inter7, gate364inter8, gate364inter9, gate364inter10, gate364inter11, gate364inter12, gate161inter0, gate161inter1, gate161inter2, gate161inter3, gate161inter4, gate161inter5, gate161inter6, gate161inter7, gate161inter8, gate161inter9, gate161inter10, gate161inter11, gate161inter12, gate395inter0, gate395inter1, gate395inter2, gate395inter3, gate395inter4, gate395inter5, gate395inter6, gate395inter7, gate395inter8, gate395inter9, gate395inter10, gate395inter11, gate395inter12, gate601inter0, gate601inter1, gate601inter2, gate601inter3, gate601inter4, gate601inter5, gate601inter6, gate601inter7, gate601inter8, gate601inter9, gate601inter10, gate601inter11, gate601inter12, gate544inter0, gate544inter1, gate544inter2, gate544inter3, gate544inter4, gate544inter5, gate544inter6, gate544inter7, gate544inter8, gate544inter9, gate544inter10, gate544inter11, gate544inter12, gate780inter0, gate780inter1, gate780inter2, gate780inter3, gate780inter4, gate780inter5, gate780inter6, gate780inter7, gate780inter8, gate780inter9, gate780inter10, gate780inter11, gate780inter12, gate675inter0, gate675inter1, gate675inter2, gate675inter3, gate675inter4, gate675inter5, gate675inter6, gate675inter7, gate675inter8, gate675inter9, gate675inter10, gate675inter11, gate675inter12, gate339inter0, gate339inter1, gate339inter2, gate339inter3, gate339inter4, gate339inter5, gate339inter6, gate339inter7, gate339inter8, gate339inter9, gate339inter10, gate339inter11, gate339inter12;


inv1 gate1( .a(N1), .O(N190) );
inv1 gate2( .a(N4), .O(N194) );
inv1 gate3( .a(N7), .O(N197) );
inv1 gate4( .a(N10), .O(N201) );
inv1 gate5( .a(N13), .O(N206) );
inv1 gate6( .a(N16), .O(N209) );
inv1 gate7( .a(N19), .O(N212) );
inv1 gate8( .a(N22), .O(N216) );
inv1 gate9( .a(N25), .O(N220) );
inv1 gate10( .a(N28), .O(N225) );
inv1 gate11( .a(N31), .O(N229) );
inv1 gate12( .a(N34), .O(N232) );
inv1 gate13( .a(N37), .O(N235) );
inv1 gate14( .a(N40), .O(N239) );
inv1 gate15( .a(N43), .O(N243) );
inv1 gate16( .a(N46), .O(N247) );

  xor2  gate1525(.a(N88), .b(N63), .O(gate17inter0));
  nand2 gate1526(.a(gate17inter0), .b(s_92), .O(gate17inter1));
  and2  gate1527(.a(N88), .b(N63), .O(gate17inter2));
  inv1  gate1528(.a(s_92), .O(gate17inter3));
  inv1  gate1529(.a(s_93), .O(gate17inter4));
  nand2 gate1530(.a(gate17inter4), .b(gate17inter3), .O(gate17inter5));
  nor2  gate1531(.a(gate17inter5), .b(gate17inter2), .O(gate17inter6));
  inv1  gate1532(.a(N63), .O(gate17inter7));
  inv1  gate1533(.a(N88), .O(gate17inter8));
  nand2 gate1534(.a(gate17inter8), .b(gate17inter7), .O(gate17inter9));
  nand2 gate1535(.a(s_93), .b(gate17inter3), .O(gate17inter10));
  nor2  gate1536(.a(gate17inter10), .b(gate17inter9), .O(gate17inter11));
  nor2  gate1537(.a(gate17inter11), .b(gate17inter6), .O(gate17inter12));
  nand2 gate1538(.a(gate17inter12), .b(gate17inter1), .O(N251));
nand2 gate18( .a(N66), .b(N91), .O(N252) );
inv1 gate19( .a(N72), .O(N253) );
inv1 gate20( .a(N72), .O(N256) );
buf1 gate21( .a(N69), .O(N257) );
buf1 gate22( .a(N69), .O(N260) );
inv1 gate23( .a(N76), .O(N263) );
inv1 gate24( .a(N79), .O(N266) );
inv1 gate25( .a(N82), .O(N269) );
inv1 gate26( .a(N85), .O(N272) );
inv1 gate27( .a(N104), .O(N275) );
inv1 gate28( .a(N104), .O(N276) );
inv1 gate29( .a(N88), .O(N277) );
inv1 gate30( .a(N91), .O(N280) );
buf1 gate31( .a(N94), .O(N283) );
inv1 gate32( .a(N94), .O(N290) );
buf1 gate33( .a(N94), .O(N297) );
inv1 gate34( .a(N94), .O(N300) );
buf1 gate35( .a(N99), .O(N303) );
inv1 gate36( .a(N99), .O(N306) );
inv1 gate37( .a(N99), .O(N313) );
buf1 gate38( .a(N104), .O(N316) );
inv1 gate39( .a(N104), .O(N319) );
buf1 gate40( .a(N104), .O(N326) );
buf1 gate41( .a(N104), .O(N331) );
inv1 gate42( .a(N104), .O(N338) );
buf1 gate43( .a(N1), .O(N343) );
buf1 gate44( .a(N4), .O(N346) );
buf1 gate45( .a(N7), .O(N349) );
buf1 gate46( .a(N10), .O(N352) );
buf1 gate47( .a(N13), .O(N355) );
buf1 gate48( .a(N16), .O(N358) );
buf1 gate49( .a(N19), .O(N361) );
buf1 gate50( .a(N22), .O(N364) );
buf1 gate51( .a(N25), .O(N367) );
buf1 gate52( .a(N28), .O(N370) );
buf1 gate53( .a(N31), .O(N373) );
buf1 gate54( .a(N34), .O(N376) );
buf1 gate55( .a(N37), .O(N379) );
buf1 gate56( .a(N40), .O(N382) );
buf1 gate57( .a(N43), .O(N385) );
buf1 gate58( .a(N46), .O(N388) );
inv1 gate59( .a(N343), .O(N534) );
inv1 gate60( .a(N346), .O(N535) );
inv1 gate61( .a(N349), .O(N536) );
inv1 gate62( .a(N352), .O(N537) );
inv1 gate63( .a(N355), .O(N538) );
inv1 gate64( .a(N358), .O(N539) );
inv1 gate65( .a(N361), .O(N540) );
inv1 gate66( .a(N364), .O(N541) );
inv1 gate67( .a(N367), .O(N542) );
inv1 gate68( .a(N370), .O(N543) );
inv1 gate69( .a(N373), .O(N544) );
inv1 gate70( .a(N376), .O(N545) );
inv1 gate71( .a(N379), .O(N546) );
inv1 gate72( .a(N382), .O(N547) );
inv1 gate73( .a(N385), .O(N548) );
inv1 gate74( .a(N388), .O(N549) );
nand2 gate75( .a(N306), .b(N331), .O(N550) );
nand2 gate76( .a(N306), .b(N331), .O(N551) );
nand2 gate77( .a(N306), .b(N331), .O(N552) );

  xor2  gate1791(.a(N331), .b(N306), .O(gate78inter0));
  nand2 gate1792(.a(gate78inter0), .b(s_130), .O(gate78inter1));
  and2  gate1793(.a(N331), .b(N306), .O(gate78inter2));
  inv1  gate1794(.a(s_130), .O(gate78inter3));
  inv1  gate1795(.a(s_131), .O(gate78inter4));
  nand2 gate1796(.a(gate78inter4), .b(gate78inter3), .O(gate78inter5));
  nor2  gate1797(.a(gate78inter5), .b(gate78inter2), .O(gate78inter6));
  inv1  gate1798(.a(N306), .O(gate78inter7));
  inv1  gate1799(.a(N331), .O(gate78inter8));
  nand2 gate1800(.a(gate78inter8), .b(gate78inter7), .O(gate78inter9));
  nand2 gate1801(.a(s_131), .b(gate78inter3), .O(gate78inter10));
  nor2  gate1802(.a(gate78inter10), .b(gate78inter9), .O(gate78inter11));
  nor2  gate1803(.a(gate78inter11), .b(gate78inter6), .O(gate78inter12));
  nand2 gate1804(.a(gate78inter12), .b(gate78inter1), .O(N553));

  xor2  gate1833(.a(N331), .b(N306), .O(gate79inter0));
  nand2 gate1834(.a(gate79inter0), .b(s_136), .O(gate79inter1));
  and2  gate1835(.a(N331), .b(N306), .O(gate79inter2));
  inv1  gate1836(.a(s_136), .O(gate79inter3));
  inv1  gate1837(.a(s_137), .O(gate79inter4));
  nand2 gate1838(.a(gate79inter4), .b(gate79inter3), .O(gate79inter5));
  nor2  gate1839(.a(gate79inter5), .b(gate79inter2), .O(gate79inter6));
  inv1  gate1840(.a(N306), .O(gate79inter7));
  inv1  gate1841(.a(N331), .O(gate79inter8));
  nand2 gate1842(.a(gate79inter8), .b(gate79inter7), .O(gate79inter9));
  nand2 gate1843(.a(s_137), .b(gate79inter3), .O(gate79inter10));
  nor2  gate1844(.a(gate79inter10), .b(gate79inter9), .O(gate79inter11));
  nor2  gate1845(.a(gate79inter11), .b(gate79inter6), .O(gate79inter12));
  nand2 gate1846(.a(gate79inter12), .b(gate79inter1), .O(N554));
nand2 gate80( .a(N306), .b(N331), .O(N555) );
buf1 gate81( .a(N190), .O(N556) );
buf1 gate82( .a(N194), .O(N559) );
buf1 gate83( .a(N206), .O(N562) );
buf1 gate84( .a(N209), .O(N565) );
buf1 gate85( .a(N225), .O(N568) );
buf1 gate86( .a(N243), .O(N571) );
and2 gate87( .a(N63), .b(N319), .O(N574) );
buf1 gate88( .a(N220), .O(N577) );
buf1 gate89( .a(N229), .O(N580) );
buf1 gate90( .a(N232), .O(N583) );
and2 gate91( .a(N66), .b(N319), .O(N586) );
buf1 gate92( .a(N239), .O(N589) );
and3 gate93( .a(N49), .b(N253), .c(N319), .O(N592) );
buf1 gate94( .a(N247), .O(N595) );
buf1 gate95( .a(N239), .O(N598) );
nand2 gate96( .a(N326), .b(N277), .O(N601) );
nand2 gate97( .a(N326), .b(N280), .O(N602) );
nand2 gate98( .a(N260), .b(N72), .O(N603) );

  xor2  gate1175(.a(N300), .b(N260), .O(gate99inter0));
  nand2 gate1176(.a(gate99inter0), .b(s_42), .O(gate99inter1));
  and2  gate1177(.a(N300), .b(N260), .O(gate99inter2));
  inv1  gate1178(.a(s_42), .O(gate99inter3));
  inv1  gate1179(.a(s_43), .O(gate99inter4));
  nand2 gate1180(.a(gate99inter4), .b(gate99inter3), .O(gate99inter5));
  nor2  gate1181(.a(gate99inter5), .b(gate99inter2), .O(gate99inter6));
  inv1  gate1182(.a(N260), .O(gate99inter7));
  inv1  gate1183(.a(N300), .O(gate99inter8));
  nand2 gate1184(.a(gate99inter8), .b(gate99inter7), .O(gate99inter9));
  nand2 gate1185(.a(s_43), .b(gate99inter3), .O(gate99inter10));
  nor2  gate1186(.a(gate99inter10), .b(gate99inter9), .O(gate99inter11));
  nor2  gate1187(.a(gate99inter11), .b(gate99inter6), .O(gate99inter12));
  nand2 gate1188(.a(gate99inter12), .b(gate99inter1), .O(N608));
nand2 gate100( .a(N256), .b(N300), .O(N612) );
buf1 gate101( .a(N201), .O(N616) );
buf1 gate102( .a(N216), .O(N619) );
buf1 gate103( .a(N220), .O(N622) );
buf1 gate104( .a(N239), .O(N625) );
buf1 gate105( .a(N190), .O(N628) );
buf1 gate106( .a(N190), .O(N631) );
buf1 gate107( .a(N194), .O(N634) );
buf1 gate108( .a(N229), .O(N637) );
buf1 gate109( .a(N197), .O(N640) );
and3 gate110( .a(N56), .b(N257), .c(N319), .O(N643) );
buf1 gate111( .a(N232), .O(N646) );
buf1 gate112( .a(N201), .O(N649) );
buf1 gate113( .a(N235), .O(N652) );
and3 gate114( .a(N60), .b(N257), .c(N319), .O(N655) );
buf1 gate115( .a(N263), .O(N658) );
buf1 gate116( .a(N263), .O(N661) );
buf1 gate117( .a(N266), .O(N664) );
buf1 gate118( .a(N266), .O(N667) );
buf1 gate119( .a(N269), .O(N670) );
buf1 gate120( .a(N269), .O(N673) );
buf1 gate121( .a(N272), .O(N676) );
buf1 gate122( .a(N272), .O(N679) );
and2 gate123( .a(N251), .b(N316), .O(N682) );
and2 gate124( .a(N252), .b(N316), .O(N685) );
buf1 gate125( .a(N197), .O(N688) );
buf1 gate126( .a(N197), .O(N691) );
buf1 gate127( .a(N212), .O(N694) );
buf1 gate128( .a(N212), .O(N697) );
buf1 gate129( .a(N247), .O(N700) );
buf1 gate130( .a(N247), .O(N703) );
buf1 gate131( .a(N235), .O(N706) );
buf1 gate132( .a(N235), .O(N709) );
buf1 gate133( .a(N201), .O(N712) );
buf1 gate134( .a(N201), .O(N715) );
buf1 gate135( .a(N206), .O(N718) );
buf1 gate136( .a(N216), .O(N721) );
and3 gate137( .a(N53), .b(N253), .c(N319), .O(N724) );
buf1 gate138( .a(N243), .O(N727) );
buf1 gate139( .a(N220), .O(N730) );
buf1 gate140( .a(N220), .O(N733) );
buf1 gate141( .a(N209), .O(N736) );
buf1 gate142( .a(N216), .O(N739) );
buf1 gate143( .a(N225), .O(N742) );
buf1 gate144( .a(N243), .O(N745) );
buf1 gate145( .a(N212), .O(N748) );
buf1 gate146( .a(N225), .O(N751) );
inv1 gate147( .a(N682), .O(N886) );
inv1 gate148( .a(N685), .O(N887) );
inv1 gate149( .a(N616), .O(N888) );
inv1 gate150( .a(N619), .O(N889) );
inv1 gate151( .a(N622), .O(N890) );
inv1 gate152( .a(N625), .O(N891) );
inv1 gate153( .a(N631), .O(N892) );
inv1 gate154( .a(N643), .O(N893) );
inv1 gate155( .a(N649), .O(N894) );
inv1 gate156( .a(N652), .O(N895) );
inv1 gate157( .a(N655), .O(N896) );
and2 gate158( .a(N49), .b(N612), .O(N897) );
and2 gate159( .a(N56), .b(N608), .O(N898) );
nand2 gate160( .a(N53), .b(N612), .O(N899) );

  xor2  gate2057(.a(N608), .b(N60), .O(gate161inter0));
  nand2 gate2058(.a(gate161inter0), .b(s_168), .O(gate161inter1));
  and2  gate2059(.a(N608), .b(N60), .O(gate161inter2));
  inv1  gate2060(.a(s_168), .O(gate161inter3));
  inv1  gate2061(.a(s_169), .O(gate161inter4));
  nand2 gate2062(.a(gate161inter4), .b(gate161inter3), .O(gate161inter5));
  nor2  gate2063(.a(gate161inter5), .b(gate161inter2), .O(gate161inter6));
  inv1  gate2064(.a(N60), .O(gate161inter7));
  inv1  gate2065(.a(N608), .O(gate161inter8));
  nand2 gate2066(.a(gate161inter8), .b(gate161inter7), .O(gate161inter9));
  nand2 gate2067(.a(s_169), .b(gate161inter3), .O(gate161inter10));
  nor2  gate2068(.a(gate161inter10), .b(gate161inter9), .O(gate161inter11));
  nor2  gate2069(.a(gate161inter11), .b(gate161inter6), .O(gate161inter12));
  nand2 gate2070(.a(gate161inter12), .b(gate161inter1), .O(N903));
nand2 gate162( .a(N49), .b(N612), .O(N907) );
nand2 gate163( .a(N56), .b(N608), .O(N910) );
inv1 gate164( .a(N661), .O(N913) );
inv1 gate165( .a(N658), .O(N914) );
inv1 gate166( .a(N667), .O(N915) );
inv1 gate167( .a(N664), .O(N916) );
inv1 gate168( .a(N673), .O(N917) );
inv1 gate169( .a(N670), .O(N918) );
inv1 gate170( .a(N679), .O(N919) );
inv1 gate171( .a(N676), .O(N920) );
nand4 gate172( .a(N277), .b(N297), .c(N326), .d(N603), .O(N921) );
nand4 gate173( .a(N280), .b(N297), .c(N326), .d(N603), .O(N922) );
nand3 gate174( .a(N303), .b(N338), .c(N603), .O(N923) );
and3 gate175( .a(N303), .b(N338), .c(N603), .O(N926) );
buf1 gate176( .a(N556), .O(N935) );
inv1 gate177( .a(N688), .O(N938) );
buf1 gate178( .a(N556), .O(N939) );
inv1 gate179( .a(N691), .O(N942) );
buf1 gate180( .a(N562), .O(N943) );
inv1 gate181( .a(N694), .O(N946) );
buf1 gate182( .a(N562), .O(N947) );
inv1 gate183( .a(N697), .O(N950) );
buf1 gate184( .a(N568), .O(N951) );
inv1 gate185( .a(N700), .O(N954) );
buf1 gate186( .a(N568), .O(N955) );
inv1 gate187( .a(N703), .O(N958) );
buf1 gate188( .a(N574), .O(N959) );
buf1 gate189( .a(N574), .O(N962) );
buf1 gate190( .a(N580), .O(N965) );
inv1 gate191( .a(N706), .O(N968) );
buf1 gate192( .a(N580), .O(N969) );
inv1 gate193( .a(N709), .O(N972) );
buf1 gate194( .a(N586), .O(N973) );
inv1 gate195( .a(N712), .O(N976) );
buf1 gate196( .a(N586), .O(N977) );
inv1 gate197( .a(N715), .O(N980) );
buf1 gate198( .a(N592), .O(N981) );
inv1 gate199( .a(N628), .O(N984) );
buf1 gate200( .a(N592), .O(N985) );
inv1 gate201( .a(N718), .O(N988) );
inv1 gate202( .a(N721), .O(N989) );
inv1 gate203( .a(N634), .O(N990) );
inv1 gate204( .a(N724), .O(N991) );
inv1 gate205( .a(N727), .O(N992) );
inv1 gate206( .a(N637), .O(N993) );
buf1 gate207( .a(N595), .O(N994) );
inv1 gate208( .a(N730), .O(N997) );
buf1 gate209( .a(N595), .O(N998) );
inv1 gate210( .a(N733), .O(N1001) );
inv1 gate211( .a(N736), .O(N1002) );
inv1 gate212( .a(N739), .O(N1003) );
inv1 gate213( .a(N640), .O(N1004) );
inv1 gate214( .a(N742), .O(N1005) );
inv1 gate215( .a(N745), .O(N1006) );
inv1 gate216( .a(N646), .O(N1007) );
inv1 gate217( .a(N748), .O(N1008) );
inv1 gate218( .a(N751), .O(N1009) );
buf1 gate219( .a(N559), .O(N1010) );
buf1 gate220( .a(N559), .O(N1013) );
buf1 gate221( .a(N565), .O(N1016) );
buf1 gate222( .a(N565), .O(N1019) );
buf1 gate223( .a(N571), .O(N1022) );
buf1 gate224( .a(N571), .O(N1025) );
buf1 gate225( .a(N577), .O(N1028) );
buf1 gate226( .a(N577), .O(N1031) );
buf1 gate227( .a(N583), .O(N1034) );
buf1 gate228( .a(N583), .O(N1037) );
buf1 gate229( .a(N589), .O(N1040) );
buf1 gate230( .a(N589), .O(N1043) );
buf1 gate231( .a(N598), .O(N1046) );
buf1 gate232( .a(N598), .O(N1049) );
nand2 gate233( .a(N619), .b(N888), .O(N1054) );
nand2 gate234( .a(N616), .b(N889), .O(N1055) );

  xor2  gate1609(.a(N890), .b(N625), .O(gate235inter0));
  nand2 gate1610(.a(gate235inter0), .b(s_104), .O(gate235inter1));
  and2  gate1611(.a(N890), .b(N625), .O(gate235inter2));
  inv1  gate1612(.a(s_104), .O(gate235inter3));
  inv1  gate1613(.a(s_105), .O(gate235inter4));
  nand2 gate1614(.a(gate235inter4), .b(gate235inter3), .O(gate235inter5));
  nor2  gate1615(.a(gate235inter5), .b(gate235inter2), .O(gate235inter6));
  inv1  gate1616(.a(N625), .O(gate235inter7));
  inv1  gate1617(.a(N890), .O(gate235inter8));
  nand2 gate1618(.a(gate235inter8), .b(gate235inter7), .O(gate235inter9));
  nand2 gate1619(.a(s_105), .b(gate235inter3), .O(gate235inter10));
  nor2  gate1620(.a(gate235inter10), .b(gate235inter9), .O(gate235inter11));
  nor2  gate1621(.a(gate235inter11), .b(gate235inter6), .O(gate235inter12));
  nand2 gate1622(.a(gate235inter12), .b(gate235inter1), .O(N1063));

  xor2  gate1931(.a(N891), .b(N622), .O(gate236inter0));
  nand2 gate1932(.a(gate236inter0), .b(s_150), .O(gate236inter1));
  and2  gate1933(.a(N891), .b(N622), .O(gate236inter2));
  inv1  gate1934(.a(s_150), .O(gate236inter3));
  inv1  gate1935(.a(s_151), .O(gate236inter4));
  nand2 gate1936(.a(gate236inter4), .b(gate236inter3), .O(gate236inter5));
  nor2  gate1937(.a(gate236inter5), .b(gate236inter2), .O(gate236inter6));
  inv1  gate1938(.a(N622), .O(gate236inter7));
  inv1  gate1939(.a(N891), .O(gate236inter8));
  nand2 gate1940(.a(gate236inter8), .b(gate236inter7), .O(gate236inter9));
  nand2 gate1941(.a(s_151), .b(gate236inter3), .O(gate236inter10));
  nor2  gate1942(.a(gate236inter10), .b(gate236inter9), .O(gate236inter11));
  nor2  gate1943(.a(gate236inter11), .b(gate236inter6), .O(gate236inter12));
  nand2 gate1944(.a(gate236inter12), .b(gate236inter1), .O(N1064));
nand2 gate237( .a(N655), .b(N895), .O(N1067) );
nand2 gate238( .a(N652), .b(N896), .O(N1068) );
nand2 gate239( .a(N721), .b(N988), .O(N1119) );
nand2 gate240( .a(N718), .b(N989), .O(N1120) );
nand2 gate241( .a(N727), .b(N991), .O(N1121) );

  xor2  gate1245(.a(N992), .b(N724), .O(gate242inter0));
  nand2 gate1246(.a(gate242inter0), .b(s_52), .O(gate242inter1));
  and2  gate1247(.a(N992), .b(N724), .O(gate242inter2));
  inv1  gate1248(.a(s_52), .O(gate242inter3));
  inv1  gate1249(.a(s_53), .O(gate242inter4));
  nand2 gate1250(.a(gate242inter4), .b(gate242inter3), .O(gate242inter5));
  nor2  gate1251(.a(gate242inter5), .b(gate242inter2), .O(gate242inter6));
  inv1  gate1252(.a(N724), .O(gate242inter7));
  inv1  gate1253(.a(N992), .O(gate242inter8));
  nand2 gate1254(.a(gate242inter8), .b(gate242inter7), .O(gate242inter9));
  nand2 gate1255(.a(s_53), .b(gate242inter3), .O(gate242inter10));
  nor2  gate1256(.a(gate242inter10), .b(gate242inter9), .O(gate242inter11));
  nor2  gate1257(.a(gate242inter11), .b(gate242inter6), .O(gate242inter12));
  nand2 gate1258(.a(gate242inter12), .b(gate242inter1), .O(N1122));

  xor2  gate951(.a(N1002), .b(N739), .O(gate243inter0));
  nand2 gate952(.a(gate243inter0), .b(s_10), .O(gate243inter1));
  and2  gate953(.a(N1002), .b(N739), .O(gate243inter2));
  inv1  gate954(.a(s_10), .O(gate243inter3));
  inv1  gate955(.a(s_11), .O(gate243inter4));
  nand2 gate956(.a(gate243inter4), .b(gate243inter3), .O(gate243inter5));
  nor2  gate957(.a(gate243inter5), .b(gate243inter2), .O(gate243inter6));
  inv1  gate958(.a(N739), .O(gate243inter7));
  inv1  gate959(.a(N1002), .O(gate243inter8));
  nand2 gate960(.a(gate243inter8), .b(gate243inter7), .O(gate243inter9));
  nand2 gate961(.a(s_11), .b(gate243inter3), .O(gate243inter10));
  nor2  gate962(.a(gate243inter10), .b(gate243inter9), .O(gate243inter11));
  nor2  gate963(.a(gate243inter11), .b(gate243inter6), .O(gate243inter12));
  nand2 gate964(.a(gate243inter12), .b(gate243inter1), .O(N1128));
nand2 gate244( .a(N736), .b(N1003), .O(N1129) );

  xor2  gate1665(.a(N1005), .b(N745), .O(gate245inter0));
  nand2 gate1666(.a(gate245inter0), .b(s_112), .O(gate245inter1));
  and2  gate1667(.a(N1005), .b(N745), .O(gate245inter2));
  inv1  gate1668(.a(s_112), .O(gate245inter3));
  inv1  gate1669(.a(s_113), .O(gate245inter4));
  nand2 gate1670(.a(gate245inter4), .b(gate245inter3), .O(gate245inter5));
  nor2  gate1671(.a(gate245inter5), .b(gate245inter2), .O(gate245inter6));
  inv1  gate1672(.a(N745), .O(gate245inter7));
  inv1  gate1673(.a(N1005), .O(gate245inter8));
  nand2 gate1674(.a(gate245inter8), .b(gate245inter7), .O(gate245inter9));
  nand2 gate1675(.a(s_113), .b(gate245inter3), .O(gate245inter10));
  nor2  gate1676(.a(gate245inter10), .b(gate245inter9), .O(gate245inter11));
  nor2  gate1677(.a(gate245inter11), .b(gate245inter6), .O(gate245inter12));
  nand2 gate1678(.a(gate245inter12), .b(gate245inter1), .O(N1130));
nand2 gate246( .a(N742), .b(N1006), .O(N1131) );

  xor2  gate965(.a(N1008), .b(N751), .O(gate247inter0));
  nand2 gate966(.a(gate247inter0), .b(s_12), .O(gate247inter1));
  and2  gate967(.a(N1008), .b(N751), .O(gate247inter2));
  inv1  gate968(.a(s_12), .O(gate247inter3));
  inv1  gate969(.a(s_13), .O(gate247inter4));
  nand2 gate970(.a(gate247inter4), .b(gate247inter3), .O(gate247inter5));
  nor2  gate971(.a(gate247inter5), .b(gate247inter2), .O(gate247inter6));
  inv1  gate972(.a(N751), .O(gate247inter7));
  inv1  gate973(.a(N1008), .O(gate247inter8));
  nand2 gate974(.a(gate247inter8), .b(gate247inter7), .O(gate247inter9));
  nand2 gate975(.a(s_13), .b(gate247inter3), .O(gate247inter10));
  nor2  gate976(.a(gate247inter10), .b(gate247inter9), .O(gate247inter11));
  nor2  gate977(.a(gate247inter11), .b(gate247inter6), .O(gate247inter12));
  nand2 gate978(.a(gate247inter12), .b(gate247inter1), .O(N1132));

  xor2  gate1063(.a(N1009), .b(N748), .O(gate248inter0));
  nand2 gate1064(.a(gate248inter0), .b(s_26), .O(gate248inter1));
  and2  gate1065(.a(N1009), .b(N748), .O(gate248inter2));
  inv1  gate1066(.a(s_26), .O(gate248inter3));
  inv1  gate1067(.a(s_27), .O(gate248inter4));
  nand2 gate1068(.a(gate248inter4), .b(gate248inter3), .O(gate248inter5));
  nor2  gate1069(.a(gate248inter5), .b(gate248inter2), .O(gate248inter6));
  inv1  gate1070(.a(N748), .O(gate248inter7));
  inv1  gate1071(.a(N1009), .O(gate248inter8));
  nand2 gate1072(.a(gate248inter8), .b(gate248inter7), .O(gate248inter9));
  nand2 gate1073(.a(s_27), .b(gate248inter3), .O(gate248inter10));
  nor2  gate1074(.a(gate248inter10), .b(gate248inter9), .O(gate248inter11));
  nor2  gate1075(.a(gate248inter11), .b(gate248inter6), .O(gate248inter12));
  nand2 gate1076(.a(gate248inter12), .b(gate248inter1), .O(N1133));
inv1 gate249( .a(N939), .O(N1148) );
inv1 gate250( .a(N935), .O(N1149) );
nand2 gate251( .a(N1054), .b(N1055), .O(N1150) );
inv1 gate252( .a(N943), .O(N1151) );
inv1 gate253( .a(N947), .O(N1152) );
inv1 gate254( .a(N955), .O(N1153) );
inv1 gate255( .a(N951), .O(N1154) );
inv1 gate256( .a(N962), .O(N1155) );
inv1 gate257( .a(N969), .O(N1156) );
inv1 gate258( .a(N977), .O(N1157) );
nand2 gate259( .a(N1063), .b(N1064), .O(N1158) );
inv1 gate260( .a(N985), .O(N1159) );

  xor2  gate1203(.a(N892), .b(N985), .O(gate261inter0));
  nand2 gate1204(.a(gate261inter0), .b(s_46), .O(gate261inter1));
  and2  gate1205(.a(N892), .b(N985), .O(gate261inter2));
  inv1  gate1206(.a(s_46), .O(gate261inter3));
  inv1  gate1207(.a(s_47), .O(gate261inter4));
  nand2 gate1208(.a(gate261inter4), .b(gate261inter3), .O(gate261inter5));
  nor2  gate1209(.a(gate261inter5), .b(gate261inter2), .O(gate261inter6));
  inv1  gate1210(.a(N985), .O(gate261inter7));
  inv1  gate1211(.a(N892), .O(gate261inter8));
  nand2 gate1212(.a(gate261inter8), .b(gate261inter7), .O(gate261inter9));
  nand2 gate1213(.a(s_47), .b(gate261inter3), .O(gate261inter10));
  nor2  gate1214(.a(gate261inter10), .b(gate261inter9), .O(gate261inter11));
  nor2  gate1215(.a(gate261inter11), .b(gate261inter6), .O(gate261inter12));
  nand2 gate1216(.a(gate261inter12), .b(gate261inter1), .O(N1160));
inv1 gate262( .a(N998), .O(N1161) );
nand2 gate263( .a(N1067), .b(N1068), .O(N1162) );
inv1 gate264( .a(N899), .O(N1163) );
buf1 gate265( .a(N899), .O(N1164) );
inv1 gate266( .a(N903), .O(N1167) );
buf1 gate267( .a(N903), .O(N1168) );
nand2 gate268( .a(N921), .b(N923), .O(N1171) );

  xor2  gate2015(.a(N923), .b(N922), .O(gate269inter0));
  nand2 gate2016(.a(gate269inter0), .b(s_162), .O(gate269inter1));
  and2  gate2017(.a(N923), .b(N922), .O(gate269inter2));
  inv1  gate2018(.a(s_162), .O(gate269inter3));
  inv1  gate2019(.a(s_163), .O(gate269inter4));
  nand2 gate2020(.a(gate269inter4), .b(gate269inter3), .O(gate269inter5));
  nor2  gate2021(.a(gate269inter5), .b(gate269inter2), .O(gate269inter6));
  inv1  gate2022(.a(N922), .O(gate269inter7));
  inv1  gate2023(.a(N923), .O(gate269inter8));
  nand2 gate2024(.a(gate269inter8), .b(gate269inter7), .O(gate269inter9));
  nand2 gate2025(.a(s_163), .b(gate269inter3), .O(gate269inter10));
  nor2  gate2026(.a(gate269inter10), .b(gate269inter9), .O(gate269inter11));
  nor2  gate2027(.a(gate269inter11), .b(gate269inter6), .O(gate269inter12));
  nand2 gate2028(.a(gate269inter12), .b(gate269inter1), .O(N1188));
inv1 gate270( .a(N1010), .O(N1205) );

  xor2  gate1105(.a(N938), .b(N1010), .O(gate271inter0));
  nand2 gate1106(.a(gate271inter0), .b(s_32), .O(gate271inter1));
  and2  gate1107(.a(N938), .b(N1010), .O(gate271inter2));
  inv1  gate1108(.a(s_32), .O(gate271inter3));
  inv1  gate1109(.a(s_33), .O(gate271inter4));
  nand2 gate1110(.a(gate271inter4), .b(gate271inter3), .O(gate271inter5));
  nor2  gate1111(.a(gate271inter5), .b(gate271inter2), .O(gate271inter6));
  inv1  gate1112(.a(N1010), .O(gate271inter7));
  inv1  gate1113(.a(N938), .O(gate271inter8));
  nand2 gate1114(.a(gate271inter8), .b(gate271inter7), .O(gate271inter9));
  nand2 gate1115(.a(s_33), .b(gate271inter3), .O(gate271inter10));
  nor2  gate1116(.a(gate271inter10), .b(gate271inter9), .O(gate271inter11));
  nor2  gate1117(.a(gate271inter11), .b(gate271inter6), .O(gate271inter12));
  nand2 gate1118(.a(gate271inter12), .b(gate271inter1), .O(N1206));
inv1 gate272( .a(N1013), .O(N1207) );
nand2 gate273( .a(N1013), .b(N942), .O(N1208) );
inv1 gate274( .a(N1016), .O(N1209) );
nand2 gate275( .a(N1016), .b(N946), .O(N1210) );
inv1 gate276( .a(N1019), .O(N1211) );
nand2 gate277( .a(N1019), .b(N950), .O(N1212) );
inv1 gate278( .a(N1022), .O(N1213) );

  xor2  gate979(.a(N954), .b(N1022), .O(gate279inter0));
  nand2 gate980(.a(gate279inter0), .b(s_14), .O(gate279inter1));
  and2  gate981(.a(N954), .b(N1022), .O(gate279inter2));
  inv1  gate982(.a(s_14), .O(gate279inter3));
  inv1  gate983(.a(s_15), .O(gate279inter4));
  nand2 gate984(.a(gate279inter4), .b(gate279inter3), .O(gate279inter5));
  nor2  gate985(.a(gate279inter5), .b(gate279inter2), .O(gate279inter6));
  inv1  gate986(.a(N1022), .O(gate279inter7));
  inv1  gate987(.a(N954), .O(gate279inter8));
  nand2 gate988(.a(gate279inter8), .b(gate279inter7), .O(gate279inter9));
  nand2 gate989(.a(s_15), .b(gate279inter3), .O(gate279inter10));
  nor2  gate990(.a(gate279inter10), .b(gate279inter9), .O(gate279inter11));
  nor2  gate991(.a(gate279inter11), .b(gate279inter6), .O(gate279inter12));
  nand2 gate992(.a(gate279inter12), .b(gate279inter1), .O(N1214));
inv1 gate280( .a(N1025), .O(N1215) );

  xor2  gate923(.a(N958), .b(N1025), .O(gate281inter0));
  nand2 gate924(.a(gate281inter0), .b(s_6), .O(gate281inter1));
  and2  gate925(.a(N958), .b(N1025), .O(gate281inter2));
  inv1  gate926(.a(s_6), .O(gate281inter3));
  inv1  gate927(.a(s_7), .O(gate281inter4));
  nand2 gate928(.a(gate281inter4), .b(gate281inter3), .O(gate281inter5));
  nor2  gate929(.a(gate281inter5), .b(gate281inter2), .O(gate281inter6));
  inv1  gate930(.a(N1025), .O(gate281inter7));
  inv1  gate931(.a(N958), .O(gate281inter8));
  nand2 gate932(.a(gate281inter8), .b(gate281inter7), .O(gate281inter9));
  nand2 gate933(.a(s_7), .b(gate281inter3), .O(gate281inter10));
  nor2  gate934(.a(gate281inter10), .b(gate281inter9), .O(gate281inter11));
  nor2  gate935(.a(gate281inter11), .b(gate281inter6), .O(gate281inter12));
  nand2 gate936(.a(gate281inter12), .b(gate281inter1), .O(N1216));
inv1 gate282( .a(N1028), .O(N1217) );
inv1 gate283( .a(N959), .O(N1218) );
inv1 gate284( .a(N1031), .O(N1219) );
inv1 gate285( .a(N1034), .O(N1220) );

  xor2  gate1427(.a(N968), .b(N1034), .O(gate286inter0));
  nand2 gate1428(.a(gate286inter0), .b(s_78), .O(gate286inter1));
  and2  gate1429(.a(N968), .b(N1034), .O(gate286inter2));
  inv1  gate1430(.a(s_78), .O(gate286inter3));
  inv1  gate1431(.a(s_79), .O(gate286inter4));
  nand2 gate1432(.a(gate286inter4), .b(gate286inter3), .O(gate286inter5));
  nor2  gate1433(.a(gate286inter5), .b(gate286inter2), .O(gate286inter6));
  inv1  gate1434(.a(N1034), .O(gate286inter7));
  inv1  gate1435(.a(N968), .O(gate286inter8));
  nand2 gate1436(.a(gate286inter8), .b(gate286inter7), .O(gate286inter9));
  nand2 gate1437(.a(s_79), .b(gate286inter3), .O(gate286inter10));
  nor2  gate1438(.a(gate286inter10), .b(gate286inter9), .O(gate286inter11));
  nor2  gate1439(.a(gate286inter11), .b(gate286inter6), .O(gate286inter12));
  nand2 gate1440(.a(gate286inter12), .b(gate286inter1), .O(N1221));
inv1 gate287( .a(N965), .O(N1222) );
inv1 gate288( .a(N1037), .O(N1223) );
nand2 gate289( .a(N1037), .b(N972), .O(N1224) );
inv1 gate290( .a(N1040), .O(N1225) );
nand2 gate291( .a(N1040), .b(N976), .O(N1226) );
inv1 gate292( .a(N973), .O(N1227) );
inv1 gate293( .a(N1043), .O(N1228) );
nand2 gate294( .a(N1043), .b(N980), .O(N1229) );
inv1 gate295( .a(N981), .O(N1230) );
nand2 gate296( .a(N981), .b(N984), .O(N1231) );
nand2 gate297( .a(N1119), .b(N1120), .O(N1232) );
nand2 gate298( .a(N1121), .b(N1122), .O(N1235) );
inv1 gate299( .a(N1046), .O(N1238) );

  xor2  gate1511(.a(N997), .b(N1046), .O(gate300inter0));
  nand2 gate1512(.a(gate300inter0), .b(s_90), .O(gate300inter1));
  and2  gate1513(.a(N997), .b(N1046), .O(gate300inter2));
  inv1  gate1514(.a(s_90), .O(gate300inter3));
  inv1  gate1515(.a(s_91), .O(gate300inter4));
  nand2 gate1516(.a(gate300inter4), .b(gate300inter3), .O(gate300inter5));
  nor2  gate1517(.a(gate300inter5), .b(gate300inter2), .O(gate300inter6));
  inv1  gate1518(.a(N1046), .O(gate300inter7));
  inv1  gate1519(.a(N997), .O(gate300inter8));
  nand2 gate1520(.a(gate300inter8), .b(gate300inter7), .O(gate300inter9));
  nand2 gate1521(.a(s_91), .b(gate300inter3), .O(gate300inter10));
  nor2  gate1522(.a(gate300inter10), .b(gate300inter9), .O(gate300inter11));
  nor2  gate1523(.a(gate300inter11), .b(gate300inter6), .O(gate300inter12));
  nand2 gate1524(.a(gate300inter12), .b(gate300inter1), .O(N1239));
inv1 gate301( .a(N994), .O(N1240) );
inv1 gate302( .a(N1049), .O(N1241) );
nand2 gate303( .a(N1049), .b(N1001), .O(N1242) );
nand2 gate304( .a(N1128), .b(N1129), .O(N1243) );
nand2 gate305( .a(N1130), .b(N1131), .O(N1246) );
nand2 gate306( .a(N1132), .b(N1133), .O(N1249) );
buf1 gate307( .a(N907), .O(N1252) );
buf1 gate308( .a(N907), .O(N1255) );
buf1 gate309( .a(N910), .O(N1258) );
buf1 gate310( .a(N910), .O(N1261) );
inv1 gate311( .a(N1150), .O(N1264) );

  xor2  gate1147(.a(N1159), .b(N631), .O(gate312inter0));
  nand2 gate1148(.a(gate312inter0), .b(s_38), .O(gate312inter1));
  and2  gate1149(.a(N1159), .b(N631), .O(gate312inter2));
  inv1  gate1150(.a(s_38), .O(gate312inter3));
  inv1  gate1151(.a(s_39), .O(gate312inter4));
  nand2 gate1152(.a(gate312inter4), .b(gate312inter3), .O(gate312inter5));
  nor2  gate1153(.a(gate312inter5), .b(gate312inter2), .O(gate312inter6));
  inv1  gate1154(.a(N631), .O(gate312inter7));
  inv1  gate1155(.a(N1159), .O(gate312inter8));
  nand2 gate1156(.a(gate312inter8), .b(gate312inter7), .O(gate312inter9));
  nand2 gate1157(.a(s_39), .b(gate312inter3), .O(gate312inter10));
  nor2  gate1158(.a(gate312inter10), .b(gate312inter9), .O(gate312inter11));
  nor2  gate1159(.a(gate312inter11), .b(gate312inter6), .O(gate312inter12));
  nand2 gate1160(.a(gate312inter12), .b(gate312inter1), .O(N1267));
nand2 gate313( .a(N688), .b(N1205), .O(N1309) );
nand2 gate314( .a(N691), .b(N1207), .O(N1310) );

  xor2  gate1343(.a(N1209), .b(N694), .O(gate315inter0));
  nand2 gate1344(.a(gate315inter0), .b(s_66), .O(gate315inter1));
  and2  gate1345(.a(N1209), .b(N694), .O(gate315inter2));
  inv1  gate1346(.a(s_66), .O(gate315inter3));
  inv1  gate1347(.a(s_67), .O(gate315inter4));
  nand2 gate1348(.a(gate315inter4), .b(gate315inter3), .O(gate315inter5));
  nor2  gate1349(.a(gate315inter5), .b(gate315inter2), .O(gate315inter6));
  inv1  gate1350(.a(N694), .O(gate315inter7));
  inv1  gate1351(.a(N1209), .O(gate315inter8));
  nand2 gate1352(.a(gate315inter8), .b(gate315inter7), .O(gate315inter9));
  nand2 gate1353(.a(s_67), .b(gate315inter3), .O(gate315inter10));
  nor2  gate1354(.a(gate315inter10), .b(gate315inter9), .O(gate315inter11));
  nor2  gate1355(.a(gate315inter11), .b(gate315inter6), .O(gate315inter12));
  nand2 gate1356(.a(gate315inter12), .b(gate315inter1), .O(N1311));
nand2 gate316( .a(N697), .b(N1211), .O(N1312) );
nand2 gate317( .a(N700), .b(N1213), .O(N1313) );
nand2 gate318( .a(N703), .b(N1215), .O(N1314) );

  xor2  gate881(.a(N1220), .b(N706), .O(gate319inter0));
  nand2 gate882(.a(gate319inter0), .b(s_0), .O(gate319inter1));
  and2  gate883(.a(N1220), .b(N706), .O(gate319inter2));
  inv1  gate884(.a(s_0), .O(gate319inter3));
  inv1  gate885(.a(s_1), .O(gate319inter4));
  nand2 gate886(.a(gate319inter4), .b(gate319inter3), .O(gate319inter5));
  nor2  gate887(.a(gate319inter5), .b(gate319inter2), .O(gate319inter6));
  inv1  gate888(.a(N706), .O(gate319inter7));
  inv1  gate889(.a(N1220), .O(gate319inter8));
  nand2 gate890(.a(gate319inter8), .b(gate319inter7), .O(gate319inter9));
  nand2 gate891(.a(s_1), .b(gate319inter3), .O(gate319inter10));
  nor2  gate892(.a(gate319inter10), .b(gate319inter9), .O(gate319inter11));
  nor2  gate893(.a(gate319inter11), .b(gate319inter6), .O(gate319inter12));
  nand2 gate894(.a(gate319inter12), .b(gate319inter1), .O(N1315));
nand2 gate320( .a(N709), .b(N1223), .O(N1316) );
nand2 gate321( .a(N712), .b(N1225), .O(N1317) );
nand2 gate322( .a(N715), .b(N1228), .O(N1318) );
inv1 gate323( .a(N1158), .O(N1319) );
nand2 gate324( .a(N628), .b(N1230), .O(N1322) );
nand2 gate325( .a(N730), .b(N1238), .O(N1327) );
nand2 gate326( .a(N733), .b(N1241), .O(N1328) );
inv1 gate327( .a(N1162), .O(N1334) );
nand2 gate328( .a(N1267), .b(N1160), .O(N1344) );
nand2 gate329( .a(N1249), .b(N894), .O(N1345) );
inv1 gate330( .a(N1249), .O(N1346) );
inv1 gate331( .a(N1255), .O(N1348) );
inv1 gate332( .a(N1252), .O(N1349) );
inv1 gate333( .a(N1261), .O(N1350) );
inv1 gate334( .a(N1258), .O(N1351) );
nand2 gate335( .a(N1309), .b(N1206), .O(N1352) );

  xor2  gate1329(.a(N1208), .b(N1310), .O(gate336inter0));
  nand2 gate1330(.a(gate336inter0), .b(s_64), .O(gate336inter1));
  and2  gate1331(.a(N1208), .b(N1310), .O(gate336inter2));
  inv1  gate1332(.a(s_64), .O(gate336inter3));
  inv1  gate1333(.a(s_65), .O(gate336inter4));
  nand2 gate1334(.a(gate336inter4), .b(gate336inter3), .O(gate336inter5));
  nor2  gate1335(.a(gate336inter5), .b(gate336inter2), .O(gate336inter6));
  inv1  gate1336(.a(N1310), .O(gate336inter7));
  inv1  gate1337(.a(N1208), .O(gate336inter8));
  nand2 gate1338(.a(gate336inter8), .b(gate336inter7), .O(gate336inter9));
  nand2 gate1339(.a(s_65), .b(gate336inter3), .O(gate336inter10));
  nor2  gate1340(.a(gate336inter10), .b(gate336inter9), .O(gate336inter11));
  nor2  gate1341(.a(gate336inter11), .b(gate336inter6), .O(gate336inter12));
  nand2 gate1342(.a(gate336inter12), .b(gate336inter1), .O(N1355));
nand2 gate337( .a(N1311), .b(N1210), .O(N1358) );
nand2 gate338( .a(N1312), .b(N1212), .O(N1361) );

  xor2  gate2141(.a(N1214), .b(N1313), .O(gate339inter0));
  nand2 gate2142(.a(gate339inter0), .b(s_180), .O(gate339inter1));
  and2  gate2143(.a(N1214), .b(N1313), .O(gate339inter2));
  inv1  gate2144(.a(s_180), .O(gate339inter3));
  inv1  gate2145(.a(s_181), .O(gate339inter4));
  nand2 gate2146(.a(gate339inter4), .b(gate339inter3), .O(gate339inter5));
  nor2  gate2147(.a(gate339inter5), .b(gate339inter2), .O(gate339inter6));
  inv1  gate2148(.a(N1313), .O(gate339inter7));
  inv1  gate2149(.a(N1214), .O(gate339inter8));
  nand2 gate2150(.a(gate339inter8), .b(gate339inter7), .O(gate339inter9));
  nand2 gate2151(.a(s_181), .b(gate339inter3), .O(gate339inter10));
  nor2  gate2152(.a(gate339inter10), .b(gate339inter9), .O(gate339inter11));
  nor2  gate2153(.a(gate339inter11), .b(gate339inter6), .O(gate339inter12));
  nand2 gate2154(.a(gate339inter12), .b(gate339inter1), .O(N1364));
nand2 gate340( .a(N1314), .b(N1216), .O(N1367) );
nand2 gate341( .a(N1315), .b(N1221), .O(N1370) );

  xor2  gate1371(.a(N1224), .b(N1316), .O(gate342inter0));
  nand2 gate1372(.a(gate342inter0), .b(s_70), .O(gate342inter1));
  and2  gate1373(.a(N1224), .b(N1316), .O(gate342inter2));
  inv1  gate1374(.a(s_70), .O(gate342inter3));
  inv1  gate1375(.a(s_71), .O(gate342inter4));
  nand2 gate1376(.a(gate342inter4), .b(gate342inter3), .O(gate342inter5));
  nor2  gate1377(.a(gate342inter5), .b(gate342inter2), .O(gate342inter6));
  inv1  gate1378(.a(N1316), .O(gate342inter7));
  inv1  gate1379(.a(N1224), .O(gate342inter8));
  nand2 gate1380(.a(gate342inter8), .b(gate342inter7), .O(gate342inter9));
  nand2 gate1381(.a(s_71), .b(gate342inter3), .O(gate342inter10));
  nor2  gate1382(.a(gate342inter10), .b(gate342inter9), .O(gate342inter11));
  nor2  gate1383(.a(gate342inter11), .b(gate342inter6), .O(gate342inter12));
  nand2 gate1384(.a(gate342inter12), .b(gate342inter1), .O(N1373));
nand2 gate343( .a(N1317), .b(N1226), .O(N1376) );

  xor2  gate1917(.a(N1229), .b(N1318), .O(gate344inter0));
  nand2 gate1918(.a(gate344inter0), .b(s_148), .O(gate344inter1));
  and2  gate1919(.a(N1229), .b(N1318), .O(gate344inter2));
  inv1  gate1920(.a(s_148), .O(gate344inter3));
  inv1  gate1921(.a(s_149), .O(gate344inter4));
  nand2 gate1922(.a(gate344inter4), .b(gate344inter3), .O(gate344inter5));
  nor2  gate1923(.a(gate344inter5), .b(gate344inter2), .O(gate344inter6));
  inv1  gate1924(.a(N1318), .O(gate344inter7));
  inv1  gate1925(.a(N1229), .O(gate344inter8));
  nand2 gate1926(.a(gate344inter8), .b(gate344inter7), .O(gate344inter9));
  nand2 gate1927(.a(s_149), .b(gate344inter3), .O(gate344inter10));
  nor2  gate1928(.a(gate344inter10), .b(gate344inter9), .O(gate344inter11));
  nor2  gate1929(.a(gate344inter11), .b(gate344inter6), .O(gate344inter12));
  nand2 gate1930(.a(gate344inter12), .b(gate344inter1), .O(N1379));
nand2 gate345( .a(N1322), .b(N1231), .O(N1383) );
inv1 gate346( .a(N1232), .O(N1386) );

  xor2  gate2029(.a(N990), .b(N1232), .O(gate347inter0));
  nand2 gate2030(.a(gate347inter0), .b(s_164), .O(gate347inter1));
  and2  gate2031(.a(N990), .b(N1232), .O(gate347inter2));
  inv1  gate2032(.a(s_164), .O(gate347inter3));
  inv1  gate2033(.a(s_165), .O(gate347inter4));
  nand2 gate2034(.a(gate347inter4), .b(gate347inter3), .O(gate347inter5));
  nor2  gate2035(.a(gate347inter5), .b(gate347inter2), .O(gate347inter6));
  inv1  gate2036(.a(N1232), .O(gate347inter7));
  inv1  gate2037(.a(N990), .O(gate347inter8));
  nand2 gate2038(.a(gate347inter8), .b(gate347inter7), .O(gate347inter9));
  nand2 gate2039(.a(s_165), .b(gate347inter3), .O(gate347inter10));
  nor2  gate2040(.a(gate347inter10), .b(gate347inter9), .O(gate347inter11));
  nor2  gate2041(.a(gate347inter11), .b(gate347inter6), .O(gate347inter12));
  nand2 gate2042(.a(gate347inter12), .b(gate347inter1), .O(N1387));
inv1 gate348( .a(N1235), .O(N1388) );
nand2 gate349( .a(N1235), .b(N993), .O(N1389) );
nand2 gate350( .a(N1327), .b(N1239), .O(N1390) );
nand2 gate351( .a(N1328), .b(N1242), .O(N1393) );
inv1 gate352( .a(N1243), .O(N1396) );

  xor2  gate1441(.a(N1004), .b(N1243), .O(gate353inter0));
  nand2 gate1442(.a(gate353inter0), .b(s_80), .O(gate353inter1));
  and2  gate1443(.a(N1004), .b(N1243), .O(gate353inter2));
  inv1  gate1444(.a(s_80), .O(gate353inter3));
  inv1  gate1445(.a(s_81), .O(gate353inter4));
  nand2 gate1446(.a(gate353inter4), .b(gate353inter3), .O(gate353inter5));
  nor2  gate1447(.a(gate353inter5), .b(gate353inter2), .O(gate353inter6));
  inv1  gate1448(.a(N1243), .O(gate353inter7));
  inv1  gate1449(.a(N1004), .O(gate353inter8));
  nand2 gate1450(.a(gate353inter8), .b(gate353inter7), .O(gate353inter9));
  nand2 gate1451(.a(s_81), .b(gate353inter3), .O(gate353inter10));
  nor2  gate1452(.a(gate353inter10), .b(gate353inter9), .O(gate353inter11));
  nor2  gate1453(.a(gate353inter11), .b(gate353inter6), .O(gate353inter12));
  nand2 gate1454(.a(gate353inter12), .b(gate353inter1), .O(N1397));
inv1 gate354( .a(N1246), .O(N1398) );
nand2 gate355( .a(N1246), .b(N1007), .O(N1399) );
inv1 gate356( .a(N1319), .O(N1409) );
nand2 gate357( .a(N649), .b(N1346), .O(N1412) );
inv1 gate358( .a(N1334), .O(N1413) );
buf1 gate359( .a(N1264), .O(N1416) );
buf1 gate360( .a(N1264), .O(N1419) );
nand2 gate361( .a(N634), .b(N1386), .O(N1433) );
nand2 gate362( .a(N637), .b(N1388), .O(N1434) );
nand2 gate363( .a(N640), .b(N1396), .O(N1438) );

  xor2  gate2043(.a(N1398), .b(N646), .O(gate364inter0));
  nand2 gate2044(.a(gate364inter0), .b(s_166), .O(gate364inter1));
  and2  gate2045(.a(N1398), .b(N646), .O(gate364inter2));
  inv1  gate2046(.a(s_166), .O(gate364inter3));
  inv1  gate2047(.a(s_167), .O(gate364inter4));
  nand2 gate2048(.a(gate364inter4), .b(gate364inter3), .O(gate364inter5));
  nor2  gate2049(.a(gate364inter5), .b(gate364inter2), .O(gate364inter6));
  inv1  gate2050(.a(N646), .O(gate364inter7));
  inv1  gate2051(.a(N1398), .O(gate364inter8));
  nand2 gate2052(.a(gate364inter8), .b(gate364inter7), .O(gate364inter9));
  nand2 gate2053(.a(s_167), .b(gate364inter3), .O(gate364inter10));
  nor2  gate2054(.a(gate364inter10), .b(gate364inter9), .O(gate364inter11));
  nor2  gate2055(.a(gate364inter11), .b(gate364inter6), .O(gate364inter12));
  nand2 gate2056(.a(gate364inter12), .b(gate364inter1), .O(N1439));
inv1 gate365( .a(N1344), .O(N1440) );
nand2 gate366( .a(N1355), .b(N1148), .O(N1443) );
inv1 gate367( .a(N1355), .O(N1444) );
nand2 gate368( .a(N1352), .b(N1149), .O(N1445) );
inv1 gate369( .a(N1352), .O(N1446) );

  xor2  gate1315(.a(N1151), .b(N1358), .O(gate370inter0));
  nand2 gate1316(.a(gate370inter0), .b(s_62), .O(gate370inter1));
  and2  gate1317(.a(N1151), .b(N1358), .O(gate370inter2));
  inv1  gate1318(.a(s_62), .O(gate370inter3));
  inv1  gate1319(.a(s_63), .O(gate370inter4));
  nand2 gate1320(.a(gate370inter4), .b(gate370inter3), .O(gate370inter5));
  nor2  gate1321(.a(gate370inter5), .b(gate370inter2), .O(gate370inter6));
  inv1  gate1322(.a(N1358), .O(gate370inter7));
  inv1  gate1323(.a(N1151), .O(gate370inter8));
  nand2 gate1324(.a(gate370inter8), .b(gate370inter7), .O(gate370inter9));
  nand2 gate1325(.a(s_63), .b(gate370inter3), .O(gate370inter10));
  nor2  gate1326(.a(gate370inter10), .b(gate370inter9), .O(gate370inter11));
  nor2  gate1327(.a(gate370inter11), .b(gate370inter6), .O(gate370inter12));
  nand2 gate1328(.a(gate370inter12), .b(gate370inter1), .O(N1447));
inv1 gate371( .a(N1358), .O(N1448) );
nand2 gate372( .a(N1361), .b(N1152), .O(N1451) );
inv1 gate373( .a(N1361), .O(N1452) );
nand2 gate374( .a(N1367), .b(N1153), .O(N1453) );
inv1 gate375( .a(N1367), .O(N1454) );
nand2 gate376( .a(N1364), .b(N1154), .O(N1455) );
inv1 gate377( .a(N1364), .O(N1456) );
nand2 gate378( .a(N1373), .b(N1156), .O(N1457) );
inv1 gate379( .a(N1373), .O(N1458) );
nand2 gate380( .a(N1379), .b(N1157), .O(N1459) );
inv1 gate381( .a(N1379), .O(N1460) );
inv1 gate382( .a(N1383), .O(N1461) );
nand2 gate383( .a(N1393), .b(N1161), .O(N1462) );
inv1 gate384( .a(N1393), .O(N1463) );

  xor2  gate1231(.a(N1412), .b(N1345), .O(gate385inter0));
  nand2 gate1232(.a(gate385inter0), .b(s_50), .O(gate385inter1));
  and2  gate1233(.a(N1412), .b(N1345), .O(gate385inter2));
  inv1  gate1234(.a(s_50), .O(gate385inter3));
  inv1  gate1235(.a(s_51), .O(gate385inter4));
  nand2 gate1236(.a(gate385inter4), .b(gate385inter3), .O(gate385inter5));
  nor2  gate1237(.a(gate385inter5), .b(gate385inter2), .O(gate385inter6));
  inv1  gate1238(.a(N1345), .O(gate385inter7));
  inv1  gate1239(.a(N1412), .O(gate385inter8));
  nand2 gate1240(.a(gate385inter8), .b(gate385inter7), .O(gate385inter9));
  nand2 gate1241(.a(s_51), .b(gate385inter3), .O(gate385inter10));
  nor2  gate1242(.a(gate385inter10), .b(gate385inter9), .O(gate385inter11));
  nor2  gate1243(.a(gate385inter11), .b(gate385inter6), .O(gate385inter12));
  nand2 gate1244(.a(gate385inter12), .b(gate385inter1), .O(N1464));
inv1 gate386( .a(N1370), .O(N1468) );
nand2 gate387( .a(N1370), .b(N1222), .O(N1469) );
inv1 gate388( .a(N1376), .O(N1470) );
nand2 gate389( .a(N1376), .b(N1227), .O(N1471) );

  xor2  gate1623(.a(N1433), .b(N1387), .O(gate390inter0));
  nand2 gate1624(.a(gate390inter0), .b(s_106), .O(gate390inter1));
  and2  gate1625(.a(N1433), .b(N1387), .O(gate390inter2));
  inv1  gate1626(.a(s_106), .O(gate390inter3));
  inv1  gate1627(.a(s_107), .O(gate390inter4));
  nand2 gate1628(.a(gate390inter4), .b(gate390inter3), .O(gate390inter5));
  nor2  gate1629(.a(gate390inter5), .b(gate390inter2), .O(gate390inter6));
  inv1  gate1630(.a(N1387), .O(gate390inter7));
  inv1  gate1631(.a(N1433), .O(gate390inter8));
  nand2 gate1632(.a(gate390inter8), .b(gate390inter7), .O(gate390inter9));
  nand2 gate1633(.a(s_107), .b(gate390inter3), .O(gate390inter10));
  nor2  gate1634(.a(gate390inter10), .b(gate390inter9), .O(gate390inter11));
  nor2  gate1635(.a(gate390inter11), .b(gate390inter6), .O(gate390inter12));
  nand2 gate1636(.a(gate390inter12), .b(gate390inter1), .O(N1472));
inv1 gate391( .a(N1390), .O(N1475) );
nand2 gate392( .a(N1390), .b(N1240), .O(N1476) );

  xor2  gate1721(.a(N1434), .b(N1389), .O(gate393inter0));
  nand2 gate1722(.a(gate393inter0), .b(s_120), .O(gate393inter1));
  and2  gate1723(.a(N1434), .b(N1389), .O(gate393inter2));
  inv1  gate1724(.a(s_120), .O(gate393inter3));
  inv1  gate1725(.a(s_121), .O(gate393inter4));
  nand2 gate1726(.a(gate393inter4), .b(gate393inter3), .O(gate393inter5));
  nor2  gate1727(.a(gate393inter5), .b(gate393inter2), .O(gate393inter6));
  inv1  gate1728(.a(N1389), .O(gate393inter7));
  inv1  gate1729(.a(N1434), .O(gate393inter8));
  nand2 gate1730(.a(gate393inter8), .b(gate393inter7), .O(gate393inter9));
  nand2 gate1731(.a(s_121), .b(gate393inter3), .O(gate393inter10));
  nor2  gate1732(.a(gate393inter10), .b(gate393inter9), .O(gate393inter11));
  nor2  gate1733(.a(gate393inter11), .b(gate393inter6), .O(gate393inter12));
  nand2 gate1734(.a(gate393inter12), .b(gate393inter1), .O(N1478));
nand2 gate394( .a(N1399), .b(N1439), .O(N1481) );

  xor2  gate2071(.a(N1438), .b(N1397), .O(gate395inter0));
  nand2 gate2072(.a(gate395inter0), .b(s_170), .O(gate395inter1));
  and2  gate2073(.a(N1438), .b(N1397), .O(gate395inter2));
  inv1  gate2074(.a(s_170), .O(gate395inter3));
  inv1  gate2075(.a(s_171), .O(gate395inter4));
  nand2 gate2076(.a(gate395inter4), .b(gate395inter3), .O(gate395inter5));
  nor2  gate2077(.a(gate395inter5), .b(gate395inter2), .O(gate395inter6));
  inv1  gate2078(.a(N1397), .O(gate395inter7));
  inv1  gate2079(.a(N1438), .O(gate395inter8));
  nand2 gate2080(.a(gate395inter8), .b(gate395inter7), .O(gate395inter9));
  nand2 gate2081(.a(s_171), .b(gate395inter3), .O(gate395inter10));
  nor2  gate2082(.a(gate395inter10), .b(gate395inter9), .O(gate395inter11));
  nor2  gate2083(.a(gate395inter11), .b(gate395inter6), .O(gate395inter12));
  nand2 gate2084(.a(gate395inter12), .b(gate395inter1), .O(N1484));
nand2 gate396( .a(N939), .b(N1444), .O(N1487) );
nand2 gate397( .a(N935), .b(N1446), .O(N1488) );
nand2 gate398( .a(N943), .b(N1448), .O(N1489) );
inv1 gate399( .a(N1419), .O(N1490) );
inv1 gate400( .a(N1416), .O(N1491) );
nand2 gate401( .a(N947), .b(N1452), .O(N1492) );

  xor2  gate1217(.a(N1454), .b(N955), .O(gate402inter0));
  nand2 gate1218(.a(gate402inter0), .b(s_48), .O(gate402inter1));
  and2  gate1219(.a(N1454), .b(N955), .O(gate402inter2));
  inv1  gate1220(.a(s_48), .O(gate402inter3));
  inv1  gate1221(.a(s_49), .O(gate402inter4));
  nand2 gate1222(.a(gate402inter4), .b(gate402inter3), .O(gate402inter5));
  nor2  gate1223(.a(gate402inter5), .b(gate402inter2), .O(gate402inter6));
  inv1  gate1224(.a(N955), .O(gate402inter7));
  inv1  gate1225(.a(N1454), .O(gate402inter8));
  nand2 gate1226(.a(gate402inter8), .b(gate402inter7), .O(gate402inter9));
  nand2 gate1227(.a(s_49), .b(gate402inter3), .O(gate402inter10));
  nor2  gate1228(.a(gate402inter10), .b(gate402inter9), .O(gate402inter11));
  nor2  gate1229(.a(gate402inter11), .b(gate402inter6), .O(gate402inter12));
  nand2 gate1230(.a(gate402inter12), .b(gate402inter1), .O(N1493));
nand2 gate403( .a(N951), .b(N1456), .O(N1494) );

  xor2  gate1357(.a(N1458), .b(N969), .O(gate404inter0));
  nand2 gate1358(.a(gate404inter0), .b(s_68), .O(gate404inter1));
  and2  gate1359(.a(N1458), .b(N969), .O(gate404inter2));
  inv1  gate1360(.a(s_68), .O(gate404inter3));
  inv1  gate1361(.a(s_69), .O(gate404inter4));
  nand2 gate1362(.a(gate404inter4), .b(gate404inter3), .O(gate404inter5));
  nor2  gate1363(.a(gate404inter5), .b(gate404inter2), .O(gate404inter6));
  inv1  gate1364(.a(N969), .O(gate404inter7));
  inv1  gate1365(.a(N1458), .O(gate404inter8));
  nand2 gate1366(.a(gate404inter8), .b(gate404inter7), .O(gate404inter9));
  nand2 gate1367(.a(s_69), .b(gate404inter3), .O(gate404inter10));
  nor2  gate1368(.a(gate404inter10), .b(gate404inter9), .O(gate404inter11));
  nor2  gate1369(.a(gate404inter11), .b(gate404inter6), .O(gate404inter12));
  nand2 gate1370(.a(gate404inter12), .b(gate404inter1), .O(N1495));
nand2 gate405( .a(N977), .b(N1460), .O(N1496) );
nand2 gate406( .a(N998), .b(N1463), .O(N1498) );
inv1 gate407( .a(N1440), .O(N1499) );
nand2 gate408( .a(N965), .b(N1468), .O(N1500) );
nand2 gate409( .a(N973), .b(N1470), .O(N1501) );
nand2 gate410( .a(N994), .b(N1475), .O(N1504) );
inv1 gate411( .a(N1464), .O(N1510) );
nand2 gate412( .a(N1443), .b(N1487), .O(N1513) );
nand2 gate413( .a(N1445), .b(N1488), .O(N1514) );
nand2 gate414( .a(N1447), .b(N1489), .O(N1517) );

  xor2  gate1777(.a(N1492), .b(N1451), .O(gate415inter0));
  nand2 gate1778(.a(gate415inter0), .b(s_128), .O(gate415inter1));
  and2  gate1779(.a(N1492), .b(N1451), .O(gate415inter2));
  inv1  gate1780(.a(s_128), .O(gate415inter3));
  inv1  gate1781(.a(s_129), .O(gate415inter4));
  nand2 gate1782(.a(gate415inter4), .b(gate415inter3), .O(gate415inter5));
  nor2  gate1783(.a(gate415inter5), .b(gate415inter2), .O(gate415inter6));
  inv1  gate1784(.a(N1451), .O(gate415inter7));
  inv1  gate1785(.a(N1492), .O(gate415inter8));
  nand2 gate1786(.a(gate415inter8), .b(gate415inter7), .O(gate415inter9));
  nand2 gate1787(.a(s_129), .b(gate415inter3), .O(gate415inter10));
  nor2  gate1788(.a(gate415inter10), .b(gate415inter9), .O(gate415inter11));
  nor2  gate1789(.a(gate415inter11), .b(gate415inter6), .O(gate415inter12));
  nand2 gate1790(.a(gate415inter12), .b(gate415inter1), .O(N1520));
nand2 gate416( .a(N1453), .b(N1493), .O(N1521) );
nand2 gate417( .a(N1455), .b(N1494), .O(N1522) );
nand2 gate418( .a(N1457), .b(N1495), .O(N1526) );
nand2 gate419( .a(N1459), .b(N1496), .O(N1527) );
inv1 gate420( .a(N1472), .O(N1528) );
nand2 gate421( .a(N1462), .b(N1498), .O(N1529) );
inv1 gate422( .a(N1478), .O(N1530) );
inv1 gate423( .a(N1481), .O(N1531) );
inv1 gate424( .a(N1484), .O(N1532) );
nand2 gate425( .a(N1471), .b(N1501), .O(N1534) );
nand2 gate426( .a(N1469), .b(N1500), .O(N1537) );

  xor2  gate1679(.a(N1504), .b(N1476), .O(gate427inter0));
  nand2 gate1680(.a(gate427inter0), .b(s_114), .O(gate427inter1));
  and2  gate1681(.a(N1504), .b(N1476), .O(gate427inter2));
  inv1  gate1682(.a(s_114), .O(gate427inter3));
  inv1  gate1683(.a(s_115), .O(gate427inter4));
  nand2 gate1684(.a(gate427inter4), .b(gate427inter3), .O(gate427inter5));
  nor2  gate1685(.a(gate427inter5), .b(gate427inter2), .O(gate427inter6));
  inv1  gate1686(.a(N1476), .O(gate427inter7));
  inv1  gate1687(.a(N1504), .O(gate427inter8));
  nand2 gate1688(.a(gate427inter8), .b(gate427inter7), .O(gate427inter9));
  nand2 gate1689(.a(s_115), .b(gate427inter3), .O(gate427inter10));
  nor2  gate1690(.a(gate427inter10), .b(gate427inter9), .O(gate427inter11));
  nor2  gate1691(.a(gate427inter11), .b(gate427inter6), .O(gate427inter12));
  nand2 gate1692(.a(gate427inter12), .b(gate427inter1), .O(N1540));
inv1 gate428( .a(N1513), .O(N1546) );
inv1 gate429( .a(N1521), .O(N1554) );
inv1 gate430( .a(N1526), .O(N1557) );
inv1 gate431( .a(N1520), .O(N1561) );
nand2 gate432( .a(N1484), .b(N1531), .O(N1567) );
nand2 gate433( .a(N1481), .b(N1532), .O(N1568) );
inv1 gate434( .a(N1510), .O(N1569) );
inv1 gate435( .a(N1527), .O(N1571) );
inv1 gate436( .a(N1529), .O(N1576) );
buf1 gate437( .a(N1522), .O(N1588) );
inv1 gate438( .a(N1534), .O(N1591) );
inv1 gate439( .a(N1537), .O(N1593) );
nand2 gate440( .a(N1540), .b(N1530), .O(N1594) );
inv1 gate441( .a(N1540), .O(N1595) );
nand2 gate442( .a(N1567), .b(N1568), .O(N1596) );
buf1 gate443( .a(N1517), .O(N1600) );
buf1 gate444( .a(N1517), .O(N1603) );
buf1 gate445( .a(N1522), .O(N1606) );
buf1 gate446( .a(N1522), .O(N1609) );
buf1 gate447( .a(N1514), .O(N1612) );
buf1 gate448( .a(N1514), .O(N1615) );
buf1 gate449( .a(N1557), .O(N1620) );
buf1 gate450( .a(N1554), .O(N1623) );
inv1 gate451( .a(N1571), .O(N1635) );
nand2 gate452( .a(N1478), .b(N1595), .O(N1636) );

  xor2  gate1189(.a(N1569), .b(N1576), .O(gate453inter0));
  nand2 gate1190(.a(gate453inter0), .b(s_44), .O(gate453inter1));
  and2  gate1191(.a(N1569), .b(N1576), .O(gate453inter2));
  inv1  gate1192(.a(s_44), .O(gate453inter3));
  inv1  gate1193(.a(s_45), .O(gate453inter4));
  nand2 gate1194(.a(gate453inter4), .b(gate453inter3), .O(gate453inter5));
  nor2  gate1195(.a(gate453inter5), .b(gate453inter2), .O(gate453inter6));
  inv1  gate1196(.a(N1576), .O(gate453inter7));
  inv1  gate1197(.a(N1569), .O(gate453inter8));
  nand2 gate1198(.a(gate453inter8), .b(gate453inter7), .O(gate453inter9));
  nand2 gate1199(.a(s_45), .b(gate453inter3), .O(gate453inter10));
  nor2  gate1200(.a(gate453inter10), .b(gate453inter9), .O(gate453inter11));
  nor2  gate1201(.a(gate453inter11), .b(gate453inter6), .O(gate453inter12));
  nand2 gate1202(.a(gate453inter12), .b(gate453inter1), .O(N1638));
inv1 gate454( .a(N1576), .O(N1639) );
buf1 gate455( .a(N1561), .O(N1640) );
buf1 gate456( .a(N1561), .O(N1643) );
buf1 gate457( .a(N1546), .O(N1647) );
buf1 gate458( .a(N1546), .O(N1651) );
buf1 gate459( .a(N1554), .O(N1658) );
buf1 gate460( .a(N1557), .O(N1661) );
buf1 gate461( .a(N1557), .O(N1664) );
nand2 gate462( .a(N1596), .b(N893), .O(N1671) );
inv1 gate463( .a(N1596), .O(N1672) );
inv1 gate464( .a(N1600), .O(N1675) );
inv1 gate465( .a(N1603), .O(N1677) );
nand2 gate466( .a(N1606), .b(N1217), .O(N1678) );
inv1 gate467( .a(N1606), .O(N1679) );
nand2 gate468( .a(N1609), .b(N1219), .O(N1680) );
inv1 gate469( .a(N1609), .O(N1681) );
inv1 gate470( .a(N1612), .O(N1682) );
inv1 gate471( .a(N1615), .O(N1683) );
nand2 gate472( .a(N1594), .b(N1636), .O(N1685) );
nand2 gate473( .a(N1510), .b(N1639), .O(N1688) );
buf1 gate474( .a(N1588), .O(N1697) );
buf1 gate475( .a(N1588), .O(N1701) );
nand2 gate476( .a(N643), .b(N1672), .O(N1706) );
inv1 gate477( .a(N1643), .O(N1707) );

  xor2  gate1273(.a(N1675), .b(N1647), .O(gate478inter0));
  nand2 gate1274(.a(gate478inter0), .b(s_56), .O(gate478inter1));
  and2  gate1275(.a(N1675), .b(N1647), .O(gate478inter2));
  inv1  gate1276(.a(s_56), .O(gate478inter3));
  inv1  gate1277(.a(s_57), .O(gate478inter4));
  nand2 gate1278(.a(gate478inter4), .b(gate478inter3), .O(gate478inter5));
  nor2  gate1279(.a(gate478inter5), .b(gate478inter2), .O(gate478inter6));
  inv1  gate1280(.a(N1647), .O(gate478inter7));
  inv1  gate1281(.a(N1675), .O(gate478inter8));
  nand2 gate1282(.a(gate478inter8), .b(gate478inter7), .O(gate478inter9));
  nand2 gate1283(.a(s_57), .b(gate478inter3), .O(gate478inter10));
  nor2  gate1284(.a(gate478inter10), .b(gate478inter9), .O(gate478inter11));
  nor2  gate1285(.a(gate478inter11), .b(gate478inter6), .O(gate478inter12));
  nand2 gate1286(.a(gate478inter12), .b(gate478inter1), .O(N1708));
inv1 gate479( .a(N1647), .O(N1709) );
nand2 gate480( .a(N1651), .b(N1677), .O(N1710) );
inv1 gate481( .a(N1651), .O(N1711) );
nand2 gate482( .a(N1028), .b(N1679), .O(N1712) );
nand2 gate483( .a(N1031), .b(N1681), .O(N1713) );
buf1 gate484( .a(N1620), .O(N1714) );
buf1 gate485( .a(N1620), .O(N1717) );
nand2 gate486( .a(N1658), .b(N1593), .O(N1720) );
inv1 gate487( .a(N1658), .O(N1721) );

  xor2  gate1455(.a(N1688), .b(N1638), .O(gate488inter0));
  nand2 gate1456(.a(gate488inter0), .b(s_82), .O(gate488inter1));
  and2  gate1457(.a(N1688), .b(N1638), .O(gate488inter2));
  inv1  gate1458(.a(s_82), .O(gate488inter3));
  inv1  gate1459(.a(s_83), .O(gate488inter4));
  nand2 gate1460(.a(gate488inter4), .b(gate488inter3), .O(gate488inter5));
  nor2  gate1461(.a(gate488inter5), .b(gate488inter2), .O(gate488inter6));
  inv1  gate1462(.a(N1638), .O(gate488inter7));
  inv1  gate1463(.a(N1688), .O(gate488inter8));
  nand2 gate1464(.a(gate488inter8), .b(gate488inter7), .O(gate488inter9));
  nand2 gate1465(.a(s_83), .b(gate488inter3), .O(gate488inter10));
  nor2  gate1466(.a(gate488inter10), .b(gate488inter9), .O(gate488inter11));
  nor2  gate1467(.a(gate488inter11), .b(gate488inter6), .O(gate488inter12));
  nand2 gate1468(.a(gate488inter12), .b(gate488inter1), .O(N1723));
inv1 gate489( .a(N1661), .O(N1727) );
inv1 gate490( .a(N1640), .O(N1728) );
inv1 gate491( .a(N1664), .O(N1730) );
buf1 gate492( .a(N1623), .O(N1731) );
buf1 gate493( .a(N1623), .O(N1734) );

  xor2  gate1133(.a(N1528), .b(N1685), .O(gate494inter0));
  nand2 gate1134(.a(gate494inter0), .b(s_36), .O(gate494inter1));
  and2  gate1135(.a(N1528), .b(N1685), .O(gate494inter2));
  inv1  gate1136(.a(s_36), .O(gate494inter3));
  inv1  gate1137(.a(s_37), .O(gate494inter4));
  nand2 gate1138(.a(gate494inter4), .b(gate494inter3), .O(gate494inter5));
  nor2  gate1139(.a(gate494inter5), .b(gate494inter2), .O(gate494inter6));
  inv1  gate1140(.a(N1685), .O(gate494inter7));
  inv1  gate1141(.a(N1528), .O(gate494inter8));
  nand2 gate1142(.a(gate494inter8), .b(gate494inter7), .O(gate494inter9));
  nand2 gate1143(.a(s_37), .b(gate494inter3), .O(gate494inter10));
  nor2  gate1144(.a(gate494inter10), .b(gate494inter9), .O(gate494inter11));
  nor2  gate1145(.a(gate494inter11), .b(gate494inter6), .O(gate494inter12));
  nand2 gate1146(.a(gate494inter12), .b(gate494inter1), .O(N1740));
inv1 gate495( .a(N1685), .O(N1741) );
nand2 gate496( .a(N1671), .b(N1706), .O(N1742) );
nand2 gate497( .a(N1600), .b(N1709), .O(N1746) );
nand2 gate498( .a(N1603), .b(N1711), .O(N1747) );
nand2 gate499( .a(N1678), .b(N1712), .O(N1748) );
nand2 gate500( .a(N1680), .b(N1713), .O(N1751) );
nand2 gate501( .a(N1537), .b(N1721), .O(N1759) );
inv1 gate502( .a(N1697), .O(N1761) );
nand2 gate503( .a(N1697), .b(N1727), .O(N1762) );
inv1 gate504( .a(N1701), .O(N1763) );

  xor2  gate1763(.a(N1730), .b(N1701), .O(gate505inter0));
  nand2 gate1764(.a(gate505inter0), .b(s_126), .O(gate505inter1));
  and2  gate1765(.a(N1730), .b(N1701), .O(gate505inter2));
  inv1  gate1766(.a(s_126), .O(gate505inter3));
  inv1  gate1767(.a(s_127), .O(gate505inter4));
  nand2 gate1768(.a(gate505inter4), .b(gate505inter3), .O(gate505inter5));
  nor2  gate1769(.a(gate505inter5), .b(gate505inter2), .O(gate505inter6));
  inv1  gate1770(.a(N1701), .O(gate505inter7));
  inv1  gate1771(.a(N1730), .O(gate505inter8));
  nand2 gate1772(.a(gate505inter8), .b(gate505inter7), .O(gate505inter9));
  nand2 gate1773(.a(s_127), .b(gate505inter3), .O(gate505inter10));
  nor2  gate1774(.a(gate505inter10), .b(gate505inter9), .O(gate505inter11));
  nor2  gate1775(.a(gate505inter11), .b(gate505inter6), .O(gate505inter12));
  nand2 gate1776(.a(gate505inter12), .b(gate505inter1), .O(N1764));
inv1 gate506( .a(N1717), .O(N1768) );
nand2 gate507( .a(N1472), .b(N1741), .O(N1769) );
nand2 gate508( .a(N1723), .b(N1413), .O(N1772) );
inv1 gate509( .a(N1723), .O(N1773) );
nand2 gate510( .a(N1708), .b(N1746), .O(N1774) );

  xor2  gate1161(.a(N1747), .b(N1710), .O(gate511inter0));
  nand2 gate1162(.a(gate511inter0), .b(s_40), .O(gate511inter1));
  and2  gate1163(.a(N1747), .b(N1710), .O(gate511inter2));
  inv1  gate1164(.a(s_40), .O(gate511inter3));
  inv1  gate1165(.a(s_41), .O(gate511inter4));
  nand2 gate1166(.a(gate511inter4), .b(gate511inter3), .O(gate511inter5));
  nor2  gate1167(.a(gate511inter5), .b(gate511inter2), .O(gate511inter6));
  inv1  gate1168(.a(N1710), .O(gate511inter7));
  inv1  gate1169(.a(N1747), .O(gate511inter8));
  nand2 gate1170(.a(gate511inter8), .b(gate511inter7), .O(gate511inter9));
  nand2 gate1171(.a(s_41), .b(gate511inter3), .O(gate511inter10));
  nor2  gate1172(.a(gate511inter10), .b(gate511inter9), .O(gate511inter11));
  nor2  gate1173(.a(gate511inter11), .b(gate511inter6), .O(gate511inter12));
  nand2 gate1174(.a(gate511inter12), .b(gate511inter1), .O(N1777));
inv1 gate512( .a(N1731), .O(N1783) );
nand2 gate513( .a(N1731), .b(N1682), .O(N1784) );
inv1 gate514( .a(N1714), .O(N1785) );
inv1 gate515( .a(N1734), .O(N1786) );
nand2 gate516( .a(N1734), .b(N1683), .O(N1787) );
nand2 gate517( .a(N1720), .b(N1759), .O(N1788) );

  xor2  gate1693(.a(N1761), .b(N1661), .O(gate518inter0));
  nand2 gate1694(.a(gate518inter0), .b(s_116), .O(gate518inter1));
  and2  gate1695(.a(N1761), .b(N1661), .O(gate518inter2));
  inv1  gate1696(.a(s_116), .O(gate518inter3));
  inv1  gate1697(.a(s_117), .O(gate518inter4));
  nand2 gate1698(.a(gate518inter4), .b(gate518inter3), .O(gate518inter5));
  nor2  gate1699(.a(gate518inter5), .b(gate518inter2), .O(gate518inter6));
  inv1  gate1700(.a(N1661), .O(gate518inter7));
  inv1  gate1701(.a(N1761), .O(gate518inter8));
  nand2 gate1702(.a(gate518inter8), .b(gate518inter7), .O(gate518inter9));
  nand2 gate1703(.a(s_117), .b(gate518inter3), .O(gate518inter10));
  nor2  gate1704(.a(gate518inter10), .b(gate518inter9), .O(gate518inter11));
  nor2  gate1705(.a(gate518inter11), .b(gate518inter6), .O(gate518inter12));
  nand2 gate1706(.a(gate518inter12), .b(gate518inter1), .O(N1791));
nand2 gate519( .a(N1664), .b(N1763), .O(N1792) );
nand2 gate520( .a(N1751), .b(N1155), .O(N1795) );
inv1 gate521( .a(N1751), .O(N1796) );

  xor2  gate909(.a(N1769), .b(N1740), .O(gate522inter0));
  nand2 gate910(.a(gate522inter0), .b(s_4), .O(gate522inter1));
  and2  gate911(.a(N1769), .b(N1740), .O(gate522inter2));
  inv1  gate912(.a(s_4), .O(gate522inter3));
  inv1  gate913(.a(s_5), .O(gate522inter4));
  nand2 gate914(.a(gate522inter4), .b(gate522inter3), .O(gate522inter5));
  nor2  gate915(.a(gate522inter5), .b(gate522inter2), .O(gate522inter6));
  inv1  gate916(.a(N1740), .O(gate522inter7));
  inv1  gate917(.a(N1769), .O(gate522inter8));
  nand2 gate918(.a(gate522inter8), .b(gate522inter7), .O(gate522inter9));
  nand2 gate919(.a(s_5), .b(gate522inter3), .O(gate522inter10));
  nor2  gate920(.a(gate522inter10), .b(gate522inter9), .O(gate522inter11));
  nor2  gate921(.a(gate522inter11), .b(gate522inter6), .O(gate522inter12));
  nand2 gate922(.a(gate522inter12), .b(gate522inter1), .O(N1798));
nand2 gate523( .a(N1334), .b(N1773), .O(N1801) );

  xor2  gate1497(.a(N290), .b(N1742), .O(gate524inter0));
  nand2 gate1498(.a(gate524inter0), .b(s_88), .O(gate524inter1));
  and2  gate1499(.a(N290), .b(N1742), .O(gate524inter2));
  inv1  gate1500(.a(s_88), .O(gate524inter3));
  inv1  gate1501(.a(s_89), .O(gate524inter4));
  nand2 gate1502(.a(gate524inter4), .b(gate524inter3), .O(gate524inter5));
  nor2  gate1503(.a(gate524inter5), .b(gate524inter2), .O(gate524inter6));
  inv1  gate1504(.a(N1742), .O(gate524inter7));
  inv1  gate1505(.a(N290), .O(gate524inter8));
  nand2 gate1506(.a(gate524inter8), .b(gate524inter7), .O(gate524inter9));
  nand2 gate1507(.a(s_89), .b(gate524inter3), .O(gate524inter10));
  nor2  gate1508(.a(gate524inter10), .b(gate524inter9), .O(gate524inter11));
  nor2  gate1509(.a(gate524inter11), .b(gate524inter6), .O(gate524inter12));
  nand2 gate1510(.a(gate524inter12), .b(gate524inter1), .O(N1802));
inv1 gate525( .a(N1748), .O(N1807) );
nand2 gate526( .a(N1748), .b(N1218), .O(N1808) );

  xor2  gate937(.a(N1783), .b(N1612), .O(gate527inter0));
  nand2 gate938(.a(gate527inter0), .b(s_8), .O(gate527inter1));
  and2  gate939(.a(N1783), .b(N1612), .O(gate527inter2));
  inv1  gate940(.a(s_8), .O(gate527inter3));
  inv1  gate941(.a(s_9), .O(gate527inter4));
  nand2 gate942(.a(gate527inter4), .b(gate527inter3), .O(gate527inter5));
  nor2  gate943(.a(gate527inter5), .b(gate527inter2), .O(gate527inter6));
  inv1  gate944(.a(N1612), .O(gate527inter7));
  inv1  gate945(.a(N1783), .O(gate527inter8));
  nand2 gate946(.a(gate527inter8), .b(gate527inter7), .O(gate527inter9));
  nand2 gate947(.a(s_9), .b(gate527inter3), .O(gate527inter10));
  nor2  gate948(.a(gate527inter10), .b(gate527inter9), .O(gate527inter11));
  nor2  gate949(.a(gate527inter11), .b(gate527inter6), .O(gate527inter12));
  nand2 gate950(.a(gate527inter12), .b(gate527inter1), .O(N1809));
nand2 gate528( .a(N1615), .b(N1786), .O(N1810) );

  xor2  gate1805(.a(N1762), .b(N1791), .O(gate529inter0));
  nand2 gate1806(.a(gate529inter0), .b(s_132), .O(gate529inter1));
  and2  gate1807(.a(N1762), .b(N1791), .O(gate529inter2));
  inv1  gate1808(.a(s_132), .O(gate529inter3));
  inv1  gate1809(.a(s_133), .O(gate529inter4));
  nand2 gate1810(.a(gate529inter4), .b(gate529inter3), .O(gate529inter5));
  nor2  gate1811(.a(gate529inter5), .b(gate529inter2), .O(gate529inter6));
  inv1  gate1812(.a(N1791), .O(gate529inter7));
  inv1  gate1813(.a(N1762), .O(gate529inter8));
  nand2 gate1814(.a(gate529inter8), .b(gate529inter7), .O(gate529inter9));
  nand2 gate1815(.a(s_133), .b(gate529inter3), .O(gate529inter10));
  nor2  gate1816(.a(gate529inter10), .b(gate529inter9), .O(gate529inter11));
  nor2  gate1817(.a(gate529inter11), .b(gate529inter6), .O(gate529inter12));
  nand2 gate1818(.a(gate529inter12), .b(gate529inter1), .O(N1812));
nand2 gate530( .a(N1792), .b(N1764), .O(N1815) );
buf1 gate531( .a(N1742), .O(N1818) );
nand2 gate532( .a(N1777), .b(N1490), .O(N1821) );
inv1 gate533( .a(N1777), .O(N1822) );
nand2 gate534( .a(N1774), .b(N1491), .O(N1823) );
inv1 gate535( .a(N1774), .O(N1824) );
nand2 gate536( .a(N962), .b(N1796), .O(N1825) );

  xor2  gate2001(.a(N1409), .b(N1788), .O(gate537inter0));
  nand2 gate2002(.a(gate537inter0), .b(s_160), .O(gate537inter1));
  and2  gate2003(.a(N1409), .b(N1788), .O(gate537inter2));
  inv1  gate2004(.a(s_160), .O(gate537inter3));
  inv1  gate2005(.a(s_161), .O(gate537inter4));
  nand2 gate2006(.a(gate537inter4), .b(gate537inter3), .O(gate537inter5));
  nor2  gate2007(.a(gate537inter5), .b(gate537inter2), .O(gate537inter6));
  inv1  gate2008(.a(N1788), .O(gate537inter7));
  inv1  gate2009(.a(N1409), .O(gate537inter8));
  nand2 gate2010(.a(gate537inter8), .b(gate537inter7), .O(gate537inter9));
  nand2 gate2011(.a(s_161), .b(gate537inter3), .O(gate537inter10));
  nor2  gate2012(.a(gate537inter10), .b(gate537inter9), .O(gate537inter11));
  nor2  gate2013(.a(gate537inter11), .b(gate537inter6), .O(gate537inter12));
  nand2 gate2014(.a(gate537inter12), .b(gate537inter1), .O(N1826));
inv1 gate538( .a(N1788), .O(N1827) );
nand2 gate539( .a(N1772), .b(N1801), .O(N1830) );

  xor2  gate1875(.a(N1807), .b(N959), .O(gate540inter0));
  nand2 gate1876(.a(gate540inter0), .b(s_142), .O(gate540inter1));
  and2  gate1877(.a(N1807), .b(N959), .O(gate540inter2));
  inv1  gate1878(.a(s_142), .O(gate540inter3));
  inv1  gate1879(.a(s_143), .O(gate540inter4));
  nand2 gate1880(.a(gate540inter4), .b(gate540inter3), .O(gate540inter5));
  nor2  gate1881(.a(gate540inter5), .b(gate540inter2), .O(gate540inter6));
  inv1  gate1882(.a(N959), .O(gate540inter7));
  inv1  gate1883(.a(N1807), .O(gate540inter8));
  nand2 gate1884(.a(gate540inter8), .b(gate540inter7), .O(gate540inter9));
  nand2 gate1885(.a(s_143), .b(gate540inter3), .O(gate540inter10));
  nor2  gate1886(.a(gate540inter10), .b(gate540inter9), .O(gate540inter11));
  nor2  gate1887(.a(gate540inter11), .b(gate540inter6), .O(gate540inter12));
  nand2 gate1888(.a(gate540inter12), .b(gate540inter1), .O(N1837));
nand2 gate541( .a(N1809), .b(N1784), .O(N1838) );
nand2 gate542( .a(N1810), .b(N1787), .O(N1841) );
nand2 gate543( .a(N1419), .b(N1822), .O(N1848) );

  xor2  gate2099(.a(N1824), .b(N1416), .O(gate544inter0));
  nand2 gate2100(.a(gate544inter0), .b(s_174), .O(gate544inter1));
  and2  gate2101(.a(N1824), .b(N1416), .O(gate544inter2));
  inv1  gate2102(.a(s_174), .O(gate544inter3));
  inv1  gate2103(.a(s_175), .O(gate544inter4));
  nand2 gate2104(.a(gate544inter4), .b(gate544inter3), .O(gate544inter5));
  nor2  gate2105(.a(gate544inter5), .b(gate544inter2), .O(gate544inter6));
  inv1  gate2106(.a(N1416), .O(gate544inter7));
  inv1  gate2107(.a(N1824), .O(gate544inter8));
  nand2 gate2108(.a(gate544inter8), .b(gate544inter7), .O(gate544inter9));
  nand2 gate2109(.a(s_175), .b(gate544inter3), .O(gate544inter10));
  nor2  gate2110(.a(gate544inter10), .b(gate544inter9), .O(gate544inter11));
  nor2  gate2111(.a(gate544inter11), .b(gate544inter6), .O(gate544inter12));
  nand2 gate2112(.a(gate544inter12), .b(gate544inter1), .O(N1849));
nand2 gate545( .a(N1795), .b(N1825), .O(N1850) );
nand2 gate546( .a(N1319), .b(N1827), .O(N1852) );

  xor2  gate1959(.a(N1707), .b(N1815), .O(gate547inter0));
  nand2 gate1960(.a(gate547inter0), .b(s_154), .O(gate547inter1));
  and2  gate1961(.a(N1707), .b(N1815), .O(gate547inter2));
  inv1  gate1962(.a(s_154), .O(gate547inter3));
  inv1  gate1963(.a(s_155), .O(gate547inter4));
  nand2 gate1964(.a(gate547inter4), .b(gate547inter3), .O(gate547inter5));
  nor2  gate1965(.a(gate547inter5), .b(gate547inter2), .O(gate547inter6));
  inv1  gate1966(.a(N1815), .O(gate547inter7));
  inv1  gate1967(.a(N1707), .O(gate547inter8));
  nand2 gate1968(.a(gate547inter8), .b(gate547inter7), .O(gate547inter9));
  nand2 gate1969(.a(s_155), .b(gate547inter3), .O(gate547inter10));
  nor2  gate1970(.a(gate547inter10), .b(gate547inter9), .O(gate547inter11));
  nor2  gate1971(.a(gate547inter11), .b(gate547inter6), .O(gate547inter12));
  nand2 gate1972(.a(gate547inter12), .b(gate547inter1), .O(N1855));
inv1 gate548( .a(N1815), .O(N1856) );
inv1 gate549( .a(N1818), .O(N1857) );
nand2 gate550( .a(N1798), .b(N290), .O(N1858) );
inv1 gate551( .a(N1812), .O(N1864) );
nand2 gate552( .a(N1812), .b(N1728), .O(N1865) );
buf1 gate553( .a(N1798), .O(N1866) );
buf1 gate554( .a(N1802), .O(N1869) );
buf1 gate555( .a(N1802), .O(N1872) );
nand2 gate556( .a(N1808), .b(N1837), .O(N1875) );
nand2 gate557( .a(N1821), .b(N1848), .O(N1878) );
nand2 gate558( .a(N1823), .b(N1849), .O(N1879) );
nand2 gate559( .a(N1841), .b(N1768), .O(N1882) );
inv1 gate560( .a(N1841), .O(N1883) );
nand2 gate561( .a(N1826), .b(N1852), .O(N1884) );
nand2 gate562( .a(N1643), .b(N1856), .O(N1885) );
nand2 gate563( .a(N1830), .b(N290), .O(N1889) );
inv1 gate564( .a(N1838), .O(N1895) );
nand2 gate565( .a(N1838), .b(N1785), .O(N1896) );
nand2 gate566( .a(N1640), .b(N1864), .O(N1897) );
inv1 gate567( .a(N1850), .O(N1898) );
buf1 gate568( .a(N1830), .O(N1902) );
inv1 gate569( .a(N1878), .O(N1910) );

  xor2  gate1021(.a(N1883), .b(N1717), .O(gate570inter0));
  nand2 gate1022(.a(gate570inter0), .b(s_20), .O(gate570inter1));
  and2  gate1023(.a(N1883), .b(N1717), .O(gate570inter2));
  inv1  gate1024(.a(s_20), .O(gate570inter3));
  inv1  gate1025(.a(s_21), .O(gate570inter4));
  nand2 gate1026(.a(gate570inter4), .b(gate570inter3), .O(gate570inter5));
  nor2  gate1027(.a(gate570inter5), .b(gate570inter2), .O(gate570inter6));
  inv1  gate1028(.a(N1717), .O(gate570inter7));
  inv1  gate1029(.a(N1883), .O(gate570inter8));
  nand2 gate1030(.a(gate570inter8), .b(gate570inter7), .O(gate570inter9));
  nand2 gate1031(.a(s_21), .b(gate570inter3), .O(gate570inter10));
  nor2  gate1032(.a(gate570inter10), .b(gate570inter9), .O(gate570inter11));
  nor2  gate1033(.a(gate570inter11), .b(gate570inter6), .O(gate570inter12));
  nand2 gate1034(.a(gate570inter12), .b(gate570inter1), .O(N1911));
inv1 gate571( .a(N1884), .O(N1912) );
nand2 gate572( .a(N1855), .b(N1885), .O(N1913) );
inv1 gate573( .a(N1866), .O(N1915) );
nand2 gate574( .a(N1872), .b(N919), .O(N1919) );
inv1 gate575( .a(N1872), .O(N1920) );
nand2 gate576( .a(N1869), .b(N920), .O(N1921) );
inv1 gate577( .a(N1869), .O(N1922) );
inv1 gate578( .a(N1875), .O(N1923) );
nand2 gate579( .a(N1714), .b(N1895), .O(N1924) );
buf1 gate580( .a(N1858), .O(N1927) );
buf1 gate581( .a(N1858), .O(N1930) );

  xor2  gate1819(.a(N1897), .b(N1865), .O(gate582inter0));
  nand2 gate1820(.a(gate582inter0), .b(s_134), .O(gate582inter1));
  and2  gate1821(.a(N1897), .b(N1865), .O(gate582inter2));
  inv1  gate1822(.a(s_134), .O(gate582inter3));
  inv1  gate1823(.a(s_135), .O(gate582inter4));
  nand2 gate1824(.a(gate582inter4), .b(gate582inter3), .O(gate582inter5));
  nor2  gate1825(.a(gate582inter5), .b(gate582inter2), .O(gate582inter6));
  inv1  gate1826(.a(N1865), .O(gate582inter7));
  inv1  gate1827(.a(N1897), .O(gate582inter8));
  nand2 gate1828(.a(gate582inter8), .b(gate582inter7), .O(gate582inter9));
  nand2 gate1829(.a(s_135), .b(gate582inter3), .O(gate582inter10));
  nor2  gate1830(.a(gate582inter10), .b(gate582inter9), .O(gate582inter11));
  nor2  gate1831(.a(gate582inter11), .b(gate582inter6), .O(gate582inter12));
  nand2 gate1832(.a(gate582inter12), .b(gate582inter1), .O(N1933));
nand2 gate583( .a(N1882), .b(N1911), .O(N1936) );
inv1 gate584( .a(N1898), .O(N1937) );
inv1 gate585( .a(N1902), .O(N1938) );
nand2 gate586( .a(N679), .b(N1920), .O(N1941) );
nand2 gate587( .a(N676), .b(N1922), .O(N1942) );
buf1 gate588( .a(N1879), .O(N1944) );
inv1 gate589( .a(N1913), .O(N1947) );
buf1 gate590( .a(N1889), .O(N1950) );
buf1 gate591( .a(N1889), .O(N1953) );
buf1 gate592( .a(N1879), .O(N1958) );
nand2 gate593( .a(N1896), .b(N1924), .O(N1961) );
and2 gate594( .a(N1910), .b(N601), .O(N1965) );
and2 gate595( .a(N602), .b(N1912), .O(N1968) );

  xor2  gate1483(.a(N917), .b(N1930), .O(gate596inter0));
  nand2 gate1484(.a(gate596inter0), .b(s_86), .O(gate596inter1));
  and2  gate1485(.a(N917), .b(N1930), .O(gate596inter2));
  inv1  gate1486(.a(s_86), .O(gate596inter3));
  inv1  gate1487(.a(s_87), .O(gate596inter4));
  nand2 gate1488(.a(gate596inter4), .b(gate596inter3), .O(gate596inter5));
  nor2  gate1489(.a(gate596inter5), .b(gate596inter2), .O(gate596inter6));
  inv1  gate1490(.a(N1930), .O(gate596inter7));
  inv1  gate1491(.a(N917), .O(gate596inter8));
  nand2 gate1492(.a(gate596inter8), .b(gate596inter7), .O(gate596inter9));
  nand2 gate1493(.a(s_87), .b(gate596inter3), .O(gate596inter10));
  nor2  gate1494(.a(gate596inter10), .b(gate596inter9), .O(gate596inter11));
  nor2  gate1495(.a(gate596inter11), .b(gate596inter6), .O(gate596inter12));
  nand2 gate1496(.a(gate596inter12), .b(gate596inter1), .O(N1975));
inv1 gate597( .a(N1930), .O(N1976) );
nand2 gate598( .a(N1927), .b(N918), .O(N1977) );
inv1 gate599( .a(N1927), .O(N1978) );
nand2 gate600( .a(N1919), .b(N1941), .O(N1979) );

  xor2  gate2085(.a(N1942), .b(N1921), .O(gate601inter0));
  nand2 gate2086(.a(gate601inter0), .b(s_172), .O(gate601inter1));
  and2  gate2087(.a(N1942), .b(N1921), .O(gate601inter2));
  inv1  gate2088(.a(s_172), .O(gate601inter3));
  inv1  gate2089(.a(s_173), .O(gate601inter4));
  nand2 gate2090(.a(gate601inter4), .b(gate601inter3), .O(gate601inter5));
  nor2  gate2091(.a(gate601inter5), .b(gate601inter2), .O(gate601inter6));
  inv1  gate2092(.a(N1921), .O(gate601inter7));
  inv1  gate2093(.a(N1942), .O(gate601inter8));
  nand2 gate2094(.a(gate601inter8), .b(gate601inter7), .O(gate601inter9));
  nand2 gate2095(.a(s_173), .b(gate601inter3), .O(gate601inter10));
  nor2  gate2096(.a(gate601inter10), .b(gate601inter9), .O(gate601inter11));
  nor2  gate2097(.a(gate601inter11), .b(gate601inter6), .O(gate601inter12));
  nand2 gate2098(.a(gate601inter12), .b(gate601inter1), .O(N1980));
inv1 gate602( .a(N1933), .O(N1985) );
inv1 gate603( .a(N1936), .O(N1987) );
inv1 gate604( .a(N1944), .O(N1999) );
nand2 gate605( .a(N1944), .b(N1937), .O(N2000) );
inv1 gate606( .a(N1947), .O(N2002) );

  xor2  gate1749(.a(N1499), .b(N1947), .O(gate607inter0));
  nand2 gate1750(.a(gate607inter0), .b(s_124), .O(gate607inter1));
  and2  gate1751(.a(N1499), .b(N1947), .O(gate607inter2));
  inv1  gate1752(.a(s_124), .O(gate607inter3));
  inv1  gate1753(.a(s_125), .O(gate607inter4));
  nand2 gate1754(.a(gate607inter4), .b(gate607inter3), .O(gate607inter5));
  nor2  gate1755(.a(gate607inter5), .b(gate607inter2), .O(gate607inter6));
  inv1  gate1756(.a(N1947), .O(gate607inter7));
  inv1  gate1757(.a(N1499), .O(gate607inter8));
  nand2 gate1758(.a(gate607inter8), .b(gate607inter7), .O(gate607inter9));
  nand2 gate1759(.a(s_125), .b(gate607inter3), .O(gate607inter10));
  nor2  gate1760(.a(gate607inter10), .b(gate607inter9), .O(gate607inter11));
  nor2  gate1761(.a(gate607inter11), .b(gate607inter6), .O(gate607inter12));
  nand2 gate1762(.a(gate607inter12), .b(gate607inter1), .O(N2003));
nand2 gate608( .a(N1953), .b(N1350), .O(N2004) );
inv1 gate609( .a(N1953), .O(N2005) );
nand2 gate610( .a(N1950), .b(N1351), .O(N2006) );
inv1 gate611( .a(N1950), .O(N2007) );
nand2 gate612( .a(N673), .b(N1976), .O(N2008) );

  xor2  gate1007(.a(N1978), .b(N670), .O(gate613inter0));
  nand2 gate1008(.a(gate613inter0), .b(s_18), .O(gate613inter1));
  and2  gate1009(.a(N1978), .b(N670), .O(gate613inter2));
  inv1  gate1010(.a(s_18), .O(gate613inter3));
  inv1  gate1011(.a(s_19), .O(gate613inter4));
  nand2 gate1012(.a(gate613inter4), .b(gate613inter3), .O(gate613inter5));
  nor2  gate1013(.a(gate613inter5), .b(gate613inter2), .O(gate613inter6));
  inv1  gate1014(.a(N670), .O(gate613inter7));
  inv1  gate1015(.a(N1978), .O(gate613inter8));
  nand2 gate1016(.a(gate613inter8), .b(gate613inter7), .O(gate613inter9));
  nand2 gate1017(.a(s_19), .b(gate613inter3), .O(gate613inter10));
  nor2  gate1018(.a(gate613inter10), .b(gate613inter9), .O(gate613inter11));
  nor2  gate1019(.a(gate613inter11), .b(gate613inter6), .O(gate613inter12));
  nand2 gate1020(.a(gate613inter12), .b(gate613inter1), .O(N2009));
inv1 gate614( .a(N1979), .O(N2012) );
inv1 gate615( .a(N1958), .O(N2013) );
nand2 gate616( .a(N1958), .b(N1923), .O(N2014) );
inv1 gate617( .a(N1961), .O(N2015) );

  xor2  gate1567(.a(N1635), .b(N1961), .O(gate618inter0));
  nand2 gate1568(.a(gate618inter0), .b(s_98), .O(gate618inter1));
  and2  gate1569(.a(N1635), .b(N1961), .O(gate618inter2));
  inv1  gate1570(.a(s_98), .O(gate618inter3));
  inv1  gate1571(.a(s_99), .O(gate618inter4));
  nand2 gate1572(.a(gate618inter4), .b(gate618inter3), .O(gate618inter5));
  nor2  gate1573(.a(gate618inter5), .b(gate618inter2), .O(gate618inter6));
  inv1  gate1574(.a(N1961), .O(gate618inter7));
  inv1  gate1575(.a(N1635), .O(gate618inter8));
  nand2 gate1576(.a(gate618inter8), .b(gate618inter7), .O(gate618inter9));
  nand2 gate1577(.a(s_99), .b(gate618inter3), .O(gate618inter10));
  nor2  gate1578(.a(gate618inter10), .b(gate618inter9), .O(gate618inter11));
  nor2  gate1579(.a(gate618inter11), .b(gate618inter6), .O(gate618inter12));
  nand2 gate1580(.a(gate618inter12), .b(gate618inter1), .O(N2016));
inv1 gate619( .a(N1965), .O(N2018) );
inv1 gate620( .a(N1968), .O(N2019) );

  xor2  gate1413(.a(N1999), .b(N1898), .O(gate621inter0));
  nand2 gate1414(.a(gate621inter0), .b(s_76), .O(gate621inter1));
  and2  gate1415(.a(N1999), .b(N1898), .O(gate621inter2));
  inv1  gate1416(.a(s_76), .O(gate621inter3));
  inv1  gate1417(.a(s_77), .O(gate621inter4));
  nand2 gate1418(.a(gate621inter4), .b(gate621inter3), .O(gate621inter5));
  nor2  gate1419(.a(gate621inter5), .b(gate621inter2), .O(gate621inter6));
  inv1  gate1420(.a(N1898), .O(gate621inter7));
  inv1  gate1421(.a(N1999), .O(gate621inter8));
  nand2 gate1422(.a(gate621inter8), .b(gate621inter7), .O(gate621inter9));
  nand2 gate1423(.a(s_77), .b(gate621inter3), .O(gate621inter10));
  nor2  gate1424(.a(gate621inter10), .b(gate621inter9), .O(gate621inter11));
  nor2  gate1425(.a(gate621inter11), .b(gate621inter6), .O(gate621inter12));
  nand2 gate1426(.a(gate621inter12), .b(gate621inter1), .O(N2020));
inv1 gate622( .a(N1987), .O(N2021) );
nand2 gate623( .a(N1987), .b(N1591), .O(N2022) );
nand2 gate624( .a(N1440), .b(N2002), .O(N2023) );
nand2 gate625( .a(N1261), .b(N2005), .O(N2024) );
nand2 gate626( .a(N1258), .b(N2007), .O(N2025) );
nand2 gate627( .a(N1975), .b(N2008), .O(N2026) );

  xor2  gate1581(.a(N2009), .b(N1977), .O(gate628inter0));
  nand2 gate1582(.a(gate628inter0), .b(s_100), .O(gate628inter1));
  and2  gate1583(.a(N2009), .b(N1977), .O(gate628inter2));
  inv1  gate1584(.a(s_100), .O(gate628inter3));
  inv1  gate1585(.a(s_101), .O(gate628inter4));
  nand2 gate1586(.a(gate628inter4), .b(gate628inter3), .O(gate628inter5));
  nor2  gate1587(.a(gate628inter5), .b(gate628inter2), .O(gate628inter6));
  inv1  gate1588(.a(N1977), .O(gate628inter7));
  inv1  gate1589(.a(N2009), .O(gate628inter8));
  nand2 gate1590(.a(gate628inter8), .b(gate628inter7), .O(gate628inter9));
  nand2 gate1591(.a(s_101), .b(gate628inter3), .O(gate628inter10));
  nor2  gate1592(.a(gate628inter10), .b(gate628inter9), .O(gate628inter11));
  nor2  gate1593(.a(gate628inter11), .b(gate628inter6), .O(gate628inter12));
  nand2 gate1594(.a(gate628inter12), .b(gate628inter1), .O(N2027));
inv1 gate629( .a(N1980), .O(N2030) );
buf1 gate630( .a(N1980), .O(N2033) );

  xor2  gate1651(.a(N2013), .b(N1875), .O(gate631inter0));
  nand2 gate1652(.a(gate631inter0), .b(s_110), .O(gate631inter1));
  and2  gate1653(.a(N2013), .b(N1875), .O(gate631inter2));
  inv1  gate1654(.a(s_110), .O(gate631inter3));
  inv1  gate1655(.a(s_111), .O(gate631inter4));
  nand2 gate1656(.a(gate631inter4), .b(gate631inter3), .O(gate631inter5));
  nor2  gate1657(.a(gate631inter5), .b(gate631inter2), .O(gate631inter6));
  inv1  gate1658(.a(N1875), .O(gate631inter7));
  inv1  gate1659(.a(N2013), .O(gate631inter8));
  nand2 gate1660(.a(gate631inter8), .b(gate631inter7), .O(gate631inter9));
  nand2 gate1661(.a(s_111), .b(gate631inter3), .O(gate631inter10));
  nor2  gate1662(.a(gate631inter10), .b(gate631inter9), .O(gate631inter11));
  nor2  gate1663(.a(gate631inter11), .b(gate631inter6), .O(gate631inter12));
  nand2 gate1664(.a(gate631inter12), .b(gate631inter1), .O(N2036));
nand2 gate632( .a(N1571), .b(N2015), .O(N2037) );
nand2 gate633( .a(N2020), .b(N2000), .O(N2038) );

  xor2  gate1035(.a(N2021), .b(N1534), .O(gate634inter0));
  nand2 gate1036(.a(gate634inter0), .b(s_22), .O(gate634inter1));
  and2  gate1037(.a(N2021), .b(N1534), .O(gate634inter2));
  inv1  gate1038(.a(s_22), .O(gate634inter3));
  inv1  gate1039(.a(s_23), .O(gate634inter4));
  nand2 gate1040(.a(gate634inter4), .b(gate634inter3), .O(gate634inter5));
  nor2  gate1041(.a(gate634inter5), .b(gate634inter2), .O(gate634inter6));
  inv1  gate1042(.a(N1534), .O(gate634inter7));
  inv1  gate1043(.a(N2021), .O(gate634inter8));
  nand2 gate1044(.a(gate634inter8), .b(gate634inter7), .O(gate634inter9));
  nand2 gate1045(.a(s_23), .b(gate634inter3), .O(gate634inter10));
  nor2  gate1046(.a(gate634inter10), .b(gate634inter9), .O(gate634inter11));
  nor2  gate1047(.a(gate634inter11), .b(gate634inter6), .O(gate634inter12));
  nand2 gate1048(.a(gate634inter12), .b(gate634inter1), .O(N2039));
nand2 gate635( .a(N2023), .b(N2003), .O(N2040) );
nand2 gate636( .a(N2004), .b(N2024), .O(N2041) );
nand2 gate637( .a(N2006), .b(N2025), .O(N2042) );
inv1 gate638( .a(N2026), .O(N2047) );
nand2 gate639( .a(N2036), .b(N2014), .O(N2052) );

  xor2  gate1945(.a(N2016), .b(N2037), .O(gate640inter0));
  nand2 gate1946(.a(gate640inter0), .b(s_152), .O(gate640inter1));
  and2  gate1947(.a(N2016), .b(N2037), .O(gate640inter2));
  inv1  gate1948(.a(s_152), .O(gate640inter3));
  inv1  gate1949(.a(s_153), .O(gate640inter4));
  nand2 gate1950(.a(gate640inter4), .b(gate640inter3), .O(gate640inter5));
  nor2  gate1951(.a(gate640inter5), .b(gate640inter2), .O(gate640inter6));
  inv1  gate1952(.a(N2037), .O(gate640inter7));
  inv1  gate1953(.a(N2016), .O(gate640inter8));
  nand2 gate1954(.a(gate640inter8), .b(gate640inter7), .O(gate640inter9));
  nand2 gate1955(.a(s_153), .b(gate640inter3), .O(gate640inter10));
  nor2  gate1956(.a(gate640inter10), .b(gate640inter9), .O(gate640inter11));
  nor2  gate1957(.a(gate640inter11), .b(gate640inter6), .O(gate640inter12));
  nand2 gate1958(.a(gate640inter12), .b(gate640inter1), .O(N2055));
inv1 gate641( .a(N2038), .O(N2060) );
nand2 gate642( .a(N2039), .b(N2022), .O(N2061) );
nand2 gate643( .a(N2040), .b(N290), .O(N2062) );
inv1 gate644( .a(N2041), .O(N2067) );
inv1 gate645( .a(N2027), .O(N2068) );
buf1 gate646( .a(N2027), .O(N2071) );
inv1 gate647( .a(N2052), .O(N2076) );
inv1 gate648( .a(N2055), .O(N2077) );
nand2 gate649( .a(N2060), .b(N290), .O(N2078) );
nand2 gate650( .a(N2061), .b(N290), .O(N2081) );
inv1 gate651( .a(N2042), .O(N2086) );
buf1 gate652( .a(N2042), .O(N2089) );
and2 gate653( .a(N2030), .b(N2068), .O(N2104) );
and2 gate654( .a(N2033), .b(N2068), .O(N2119) );
and2 gate655( .a(N2030), .b(N2071), .O(N2129) );
and2 gate656( .a(N2033), .b(N2071), .O(N2143) );
buf1 gate657( .a(N2062), .O(N2148) );
buf1 gate658( .a(N2062), .O(N2151) );
buf1 gate659( .a(N2078), .O(N2196) );
buf1 gate660( .a(N2078), .O(N2199) );
buf1 gate661( .a(N2081), .O(N2202) );
buf1 gate662( .a(N2081), .O(N2205) );
nand2 gate663( .a(N2151), .b(N915), .O(N2214) );
inv1 gate664( .a(N2151), .O(N2215) );
nand2 gate665( .a(N2148), .b(N916), .O(N2216) );
inv1 gate666( .a(N2148), .O(N2217) );
nand2 gate667( .a(N2199), .b(N1348), .O(N2222) );
inv1 gate668( .a(N2199), .O(N2223) );
nand2 gate669( .a(N2196), .b(N1349), .O(N2224) );
inv1 gate670( .a(N2196), .O(N2225) );
nand2 gate671( .a(N2205), .b(N913), .O(N2226) );
inv1 gate672( .a(N2205), .O(N2227) );
nand2 gate673( .a(N2202), .b(N914), .O(N2228) );
inv1 gate674( .a(N2202), .O(N2229) );

  xor2  gate2127(.a(N2215), .b(N667), .O(gate675inter0));
  nand2 gate2128(.a(gate675inter0), .b(s_178), .O(gate675inter1));
  and2  gate2129(.a(N2215), .b(N667), .O(gate675inter2));
  inv1  gate2130(.a(s_178), .O(gate675inter3));
  inv1  gate2131(.a(s_179), .O(gate675inter4));
  nand2 gate2132(.a(gate675inter4), .b(gate675inter3), .O(gate675inter5));
  nor2  gate2133(.a(gate675inter5), .b(gate675inter2), .O(gate675inter6));
  inv1  gate2134(.a(N667), .O(gate675inter7));
  inv1  gate2135(.a(N2215), .O(gate675inter8));
  nand2 gate2136(.a(gate675inter8), .b(gate675inter7), .O(gate675inter9));
  nand2 gate2137(.a(s_179), .b(gate675inter3), .O(gate675inter10));
  nor2  gate2138(.a(gate675inter10), .b(gate675inter9), .O(gate675inter11));
  nor2  gate2139(.a(gate675inter11), .b(gate675inter6), .O(gate675inter12));
  nand2 gate2140(.a(gate675inter12), .b(gate675inter1), .O(N2230));

  xor2  gate1861(.a(N2217), .b(N664), .O(gate676inter0));
  nand2 gate1862(.a(gate676inter0), .b(s_140), .O(gate676inter1));
  and2  gate1863(.a(N2217), .b(N664), .O(gate676inter2));
  inv1  gate1864(.a(s_140), .O(gate676inter3));
  inv1  gate1865(.a(s_141), .O(gate676inter4));
  nand2 gate1866(.a(gate676inter4), .b(gate676inter3), .O(gate676inter5));
  nor2  gate1867(.a(gate676inter5), .b(gate676inter2), .O(gate676inter6));
  inv1  gate1868(.a(N664), .O(gate676inter7));
  inv1  gate1869(.a(N2217), .O(gate676inter8));
  nand2 gate1870(.a(gate676inter8), .b(gate676inter7), .O(gate676inter9));
  nand2 gate1871(.a(s_141), .b(gate676inter3), .O(gate676inter10));
  nor2  gate1872(.a(gate676inter10), .b(gate676inter9), .O(gate676inter11));
  nor2  gate1873(.a(gate676inter11), .b(gate676inter6), .O(gate676inter12));
  nand2 gate1874(.a(gate676inter12), .b(gate676inter1), .O(N2231));
nand2 gate677( .a(N1255), .b(N2223), .O(N2232) );
nand2 gate678( .a(N1252), .b(N2225), .O(N2233) );
nand2 gate679( .a(N661), .b(N2227), .O(N2234) );
nand2 gate680( .a(N658), .b(N2229), .O(N2235) );

  xor2  gate1091(.a(N2230), .b(N2214), .O(gate681inter0));
  nand2 gate1092(.a(gate681inter0), .b(s_30), .O(gate681inter1));
  and2  gate1093(.a(N2230), .b(N2214), .O(gate681inter2));
  inv1  gate1094(.a(s_30), .O(gate681inter3));
  inv1  gate1095(.a(s_31), .O(gate681inter4));
  nand2 gate1096(.a(gate681inter4), .b(gate681inter3), .O(gate681inter5));
  nor2  gate1097(.a(gate681inter5), .b(gate681inter2), .O(gate681inter6));
  inv1  gate1098(.a(N2214), .O(gate681inter7));
  inv1  gate1099(.a(N2230), .O(gate681inter8));
  nand2 gate1100(.a(gate681inter8), .b(gate681inter7), .O(gate681inter9));
  nand2 gate1101(.a(s_31), .b(gate681inter3), .O(gate681inter10));
  nor2  gate1102(.a(gate681inter10), .b(gate681inter9), .O(gate681inter11));
  nor2  gate1103(.a(gate681inter11), .b(gate681inter6), .O(gate681inter12));
  nand2 gate1104(.a(gate681inter12), .b(gate681inter1), .O(N2236));
nand2 gate682( .a(N2216), .b(N2231), .O(N2237) );
nand2 gate683( .a(N2222), .b(N2232), .O(N2240) );
nand2 gate684( .a(N2224), .b(N2233), .O(N2241) );
nand2 gate685( .a(N2226), .b(N2234), .O(N2244) );
nand2 gate686( .a(N2228), .b(N2235), .O(N2245) );
inv1 gate687( .a(N2236), .O(N2250) );
inv1 gate688( .a(N2240), .O(N2253) );
inv1 gate689( .a(N2244), .O(N2256) );
inv1 gate690( .a(N2237), .O(N2257) );
buf1 gate691( .a(N2237), .O(N2260) );
inv1 gate692( .a(N2241), .O(N2263) );
and2 gate693( .a(N1164), .b(N2241), .O(N2266) );
inv1 gate694( .a(N2245), .O(N2269) );
and2 gate695( .a(N1168), .b(N2245), .O(N2272) );
nand8 gate696( .a(N2067), .b(N2012), .c(N2047), .d(N2250), .e(N899), .f(N2256), .g(N2253), .h(N903), .O(N2279) );
buf1 gate697( .a(N2266), .O(N2286) );
buf1 gate698( .a(N2266), .O(N2297) );
buf1 gate699( .a(N2272), .O(N2315) );
buf1 gate700( .a(N2272), .O(N2326) );
and2 gate701( .a(N2086), .b(N2257), .O(N2340) );
and2 gate702( .a(N2089), .b(N2257), .O(N2353) );
and2 gate703( .a(N2086), .b(N2260), .O(N2361) );
and2 gate704( .a(N2089), .b(N2260), .O(N2375) );
and4 gate705( .a(N338), .b(N2279), .c(N313), .d(N313), .O(N2384) );
and2 gate706( .a(N1163), .b(N2263), .O(N2385) );
and2 gate707( .a(N1164), .b(N2263), .O(N2386) );
and2 gate708( .a(N1167), .b(N2269), .O(N2426) );
and2 gate709( .a(N1168), .b(N2269), .O(N2427) );
nand5 gate710( .a(N2286), .b(N2315), .c(N2361), .d(N2104), .e(N1171), .O(N2537) );
nand5 gate711( .a(N2286), .b(N2315), .c(N2340), .d(N2129), .e(N1171), .O(N2540) );
nand5 gate712( .a(N2286), .b(N2315), .c(N2340), .d(N2119), .e(N1171), .O(N2543) );
nand5 gate713( .a(N2286), .b(N2315), .c(N2353), .d(N2104), .e(N1171), .O(N2546) );
nand5 gate714( .a(N2297), .b(N2315), .c(N2375), .d(N2119), .e(N1188), .O(N2549) );
nand5 gate715( .a(N2297), .b(N2326), .c(N2361), .d(N2143), .e(N1188), .O(N2552) );
nand5 gate716( .a(N2297), .b(N2326), .c(N2375), .d(N2129), .e(N1188), .O(N2555) );
and5 gate717( .a(N2286), .b(N2315), .c(N2361), .d(N2104), .e(N1171), .O(N2558) );
and5 gate718( .a(N2286), .b(N2315), .c(N2340), .d(N2129), .e(N1171), .O(N2561) );
and5 gate719( .a(N2286), .b(N2315), .c(N2340), .d(N2119), .e(N1171), .O(N2564) );
and5 gate720( .a(N2286), .b(N2315), .c(N2353), .d(N2104), .e(N1171), .O(N2567) );
and5 gate721( .a(N2297), .b(N2315), .c(N2375), .d(N2119), .e(N1188), .O(N2570) );
and5 gate722( .a(N2297), .b(N2326), .c(N2361), .d(N2143), .e(N1188), .O(N2573) );
and5 gate723( .a(N2297), .b(N2326), .c(N2375), .d(N2129), .e(N1188), .O(N2576) );
nand5 gate724( .a(N2286), .b(N2427), .c(N2361), .d(N2129), .e(N1171), .O(N2594) );
nand5 gate725( .a(N2297), .b(N2427), .c(N2361), .d(N2119), .e(N1171), .O(N2597) );
nand5 gate726( .a(N2297), .b(N2427), .c(N2375), .d(N2104), .e(N1171), .O(N2600) );
nand5 gate727( .a(N2297), .b(N2427), .c(N2340), .d(N2143), .e(N1171), .O(N2603) );
nand5 gate728( .a(N2297), .b(N2427), .c(N2353), .d(N2129), .e(N1188), .O(N2606) );
nand5 gate729( .a(N2386), .b(N2326), .c(N2361), .d(N2129), .e(N1188), .O(N2611) );
nand5 gate730( .a(N2386), .b(N2326), .c(N2361), .d(N2119), .e(N1188), .O(N2614) );
nand5 gate731( .a(N2386), .b(N2326), .c(N2375), .d(N2104), .e(N1188), .O(N2617) );
nand5 gate732( .a(N2386), .b(N2326), .c(N2353), .d(N2129), .e(N1188), .O(N2620) );
nand5 gate733( .a(N2297), .b(N2427), .c(N2340), .d(N2104), .e(N926), .O(N2627) );
nand5 gate734( .a(N2386), .b(N2326), .c(N2340), .d(N2104), .e(N926), .O(N2628) );
nand5 gate735( .a(N2386), .b(N2427), .c(N2361), .d(N2104), .e(N926), .O(N2629) );
nand5 gate736( .a(N2386), .b(N2427), .c(N2340), .d(N2129), .e(N926), .O(N2630) );
nand5 gate737( .a(N2386), .b(N2427), .c(N2340), .d(N2119), .e(N926), .O(N2631) );
nand5 gate738( .a(N2386), .b(N2427), .c(N2353), .d(N2104), .e(N926), .O(N2632) );
nand5 gate739( .a(N2386), .b(N2426), .c(N2340), .d(N2104), .e(N926), .O(N2633) );
nand5 gate740( .a(N2385), .b(N2427), .c(N2340), .d(N2104), .e(N926), .O(N2634) );
and5 gate741( .a(N2286), .b(N2427), .c(N2361), .d(N2129), .e(N1171), .O(N2639) );
and5 gate742( .a(N2297), .b(N2427), .c(N2361), .d(N2119), .e(N1171), .O(N2642) );
and5 gate743( .a(N2297), .b(N2427), .c(N2375), .d(N2104), .e(N1171), .O(N2645) );
and5 gate744( .a(N2297), .b(N2427), .c(N2340), .d(N2143), .e(N1171), .O(N2648) );
and5 gate745( .a(N2297), .b(N2427), .c(N2353), .d(N2129), .e(N1188), .O(N2651) );
and5 gate746( .a(N2386), .b(N2326), .c(N2361), .d(N2129), .e(N1188), .O(N2655) );
and5 gate747( .a(N2386), .b(N2326), .c(N2361), .d(N2119), .e(N1188), .O(N2658) );
and5 gate748( .a(N2386), .b(N2326), .c(N2375), .d(N2104), .e(N1188), .O(N2661) );
and5 gate749( .a(N2386), .b(N2326), .c(N2353), .d(N2129), .e(N1188), .O(N2664) );
nand2 gate750( .a(N2558), .b(N534), .O(N2669) );
inv1 gate751( .a(N2558), .O(N2670) );

  xor2  gate1385(.a(N535), .b(N2561), .O(gate752inter0));
  nand2 gate1386(.a(gate752inter0), .b(s_72), .O(gate752inter1));
  and2  gate1387(.a(N535), .b(N2561), .O(gate752inter2));
  inv1  gate1388(.a(s_72), .O(gate752inter3));
  inv1  gate1389(.a(s_73), .O(gate752inter4));
  nand2 gate1390(.a(gate752inter4), .b(gate752inter3), .O(gate752inter5));
  nor2  gate1391(.a(gate752inter5), .b(gate752inter2), .O(gate752inter6));
  inv1  gate1392(.a(N2561), .O(gate752inter7));
  inv1  gate1393(.a(N535), .O(gate752inter8));
  nand2 gate1394(.a(gate752inter8), .b(gate752inter7), .O(gate752inter9));
  nand2 gate1395(.a(s_73), .b(gate752inter3), .O(gate752inter10));
  nor2  gate1396(.a(gate752inter10), .b(gate752inter9), .O(gate752inter11));
  nor2  gate1397(.a(gate752inter11), .b(gate752inter6), .O(gate752inter12));
  nand2 gate1398(.a(gate752inter12), .b(gate752inter1), .O(N2671));
inv1 gate753( .a(N2561), .O(N2672) );

  xor2  gate1301(.a(N536), .b(N2564), .O(gate754inter0));
  nand2 gate1302(.a(gate754inter0), .b(s_60), .O(gate754inter1));
  and2  gate1303(.a(N536), .b(N2564), .O(gate754inter2));
  inv1  gate1304(.a(s_60), .O(gate754inter3));
  inv1  gate1305(.a(s_61), .O(gate754inter4));
  nand2 gate1306(.a(gate754inter4), .b(gate754inter3), .O(gate754inter5));
  nor2  gate1307(.a(gate754inter5), .b(gate754inter2), .O(gate754inter6));
  inv1  gate1308(.a(N2564), .O(gate754inter7));
  inv1  gate1309(.a(N536), .O(gate754inter8));
  nand2 gate1310(.a(gate754inter8), .b(gate754inter7), .O(gate754inter9));
  nand2 gate1311(.a(s_61), .b(gate754inter3), .O(gate754inter10));
  nor2  gate1312(.a(gate754inter10), .b(gate754inter9), .O(gate754inter11));
  nor2  gate1313(.a(gate754inter11), .b(gate754inter6), .O(gate754inter12));
  nand2 gate1314(.a(gate754inter12), .b(gate754inter1), .O(N2673));
inv1 gate755( .a(N2564), .O(N2674) );

  xor2  gate1539(.a(N537), .b(N2567), .O(gate756inter0));
  nand2 gate1540(.a(gate756inter0), .b(s_94), .O(gate756inter1));
  and2  gate1541(.a(N537), .b(N2567), .O(gate756inter2));
  inv1  gate1542(.a(s_94), .O(gate756inter3));
  inv1  gate1543(.a(s_95), .O(gate756inter4));
  nand2 gate1544(.a(gate756inter4), .b(gate756inter3), .O(gate756inter5));
  nor2  gate1545(.a(gate756inter5), .b(gate756inter2), .O(gate756inter6));
  inv1  gate1546(.a(N2567), .O(gate756inter7));
  inv1  gate1547(.a(N537), .O(gate756inter8));
  nand2 gate1548(.a(gate756inter8), .b(gate756inter7), .O(gate756inter9));
  nand2 gate1549(.a(s_95), .b(gate756inter3), .O(gate756inter10));
  nor2  gate1550(.a(gate756inter10), .b(gate756inter9), .O(gate756inter11));
  nor2  gate1551(.a(gate756inter11), .b(gate756inter6), .O(gate756inter12));
  nand2 gate1552(.a(gate756inter12), .b(gate756inter1), .O(N2675));
inv1 gate757( .a(N2567), .O(N2676) );
nand2 gate758( .a(N2570), .b(N543), .O(N2682) );
inv1 gate759( .a(N2570), .O(N2683) );

  xor2  gate1847(.a(N548), .b(N2573), .O(gate760inter0));
  nand2 gate1848(.a(gate760inter0), .b(s_138), .O(gate760inter1));
  and2  gate1849(.a(N548), .b(N2573), .O(gate760inter2));
  inv1  gate1850(.a(s_138), .O(gate760inter3));
  inv1  gate1851(.a(s_139), .O(gate760inter4));
  nand2 gate1852(.a(gate760inter4), .b(gate760inter3), .O(gate760inter5));
  nor2  gate1853(.a(gate760inter5), .b(gate760inter2), .O(gate760inter6));
  inv1  gate1854(.a(N2573), .O(gate760inter7));
  inv1  gate1855(.a(N548), .O(gate760inter8));
  nand2 gate1856(.a(gate760inter8), .b(gate760inter7), .O(gate760inter9));
  nand2 gate1857(.a(s_139), .b(gate760inter3), .O(gate760inter10));
  nor2  gate1858(.a(gate760inter10), .b(gate760inter9), .O(gate760inter11));
  nor2  gate1859(.a(gate760inter11), .b(gate760inter6), .O(gate760inter12));
  nand2 gate1860(.a(gate760inter12), .b(gate760inter1), .O(N2688));
inv1 gate761( .a(N2573), .O(N2689) );
nand2 gate762( .a(N2576), .b(N549), .O(N2690) );
inv1 gate763( .a(N2576), .O(N2691) );
and8 gate764( .a(N2627), .b(N2628), .c(N2629), .d(N2630), .e(N2631), .f(N2632), .g(N2633), .h(N2634), .O(N2710) );
nand2 gate765( .a(N343), .b(N2670), .O(N2720) );
nand2 gate766( .a(N346), .b(N2672), .O(N2721) );
nand2 gate767( .a(N349), .b(N2674), .O(N2722) );
nand2 gate768( .a(N352), .b(N2676), .O(N2723) );
nand2 gate769( .a(N2639), .b(N538), .O(N2724) );
inv1 gate770( .a(N2639), .O(N2725) );
nand2 gate771( .a(N2642), .b(N539), .O(N2726) );
inv1 gate772( .a(N2642), .O(N2727) );

  xor2  gate1595(.a(N540), .b(N2645), .O(gate773inter0));
  nand2 gate1596(.a(gate773inter0), .b(s_102), .O(gate773inter1));
  and2  gate1597(.a(N540), .b(N2645), .O(gate773inter2));
  inv1  gate1598(.a(s_102), .O(gate773inter3));
  inv1  gate1599(.a(s_103), .O(gate773inter4));
  nand2 gate1600(.a(gate773inter4), .b(gate773inter3), .O(gate773inter5));
  nor2  gate1601(.a(gate773inter5), .b(gate773inter2), .O(gate773inter6));
  inv1  gate1602(.a(N2645), .O(gate773inter7));
  inv1  gate1603(.a(N540), .O(gate773inter8));
  nand2 gate1604(.a(gate773inter8), .b(gate773inter7), .O(gate773inter9));
  nand2 gate1605(.a(s_103), .b(gate773inter3), .O(gate773inter10));
  nor2  gate1606(.a(gate773inter10), .b(gate773inter9), .O(gate773inter11));
  nor2  gate1607(.a(gate773inter11), .b(gate773inter6), .O(gate773inter12));
  nand2 gate1608(.a(gate773inter12), .b(gate773inter1), .O(N2728));
inv1 gate774( .a(N2645), .O(N2729) );
nand2 gate775( .a(N2648), .b(N541), .O(N2730) );
inv1 gate776( .a(N2648), .O(N2731) );
nand2 gate777( .a(N2651), .b(N542), .O(N2732) );
inv1 gate778( .a(N2651), .O(N2733) );
nand2 gate779( .a(N370), .b(N2683), .O(N2734) );

  xor2  gate2113(.a(N544), .b(N2655), .O(gate780inter0));
  nand2 gate2114(.a(gate780inter0), .b(s_176), .O(gate780inter1));
  and2  gate2115(.a(N544), .b(N2655), .O(gate780inter2));
  inv1  gate2116(.a(s_176), .O(gate780inter3));
  inv1  gate2117(.a(s_177), .O(gate780inter4));
  nand2 gate2118(.a(gate780inter4), .b(gate780inter3), .O(gate780inter5));
  nor2  gate2119(.a(gate780inter5), .b(gate780inter2), .O(gate780inter6));
  inv1  gate2120(.a(N2655), .O(gate780inter7));
  inv1  gate2121(.a(N544), .O(gate780inter8));
  nand2 gate2122(.a(gate780inter8), .b(gate780inter7), .O(gate780inter9));
  nand2 gate2123(.a(s_177), .b(gate780inter3), .O(gate780inter10));
  nor2  gate2124(.a(gate780inter10), .b(gate780inter9), .O(gate780inter11));
  nor2  gate2125(.a(gate780inter11), .b(gate780inter6), .O(gate780inter12));
  nand2 gate2126(.a(gate780inter12), .b(gate780inter1), .O(N2735));
inv1 gate781( .a(N2655), .O(N2736) );
nand2 gate782( .a(N2658), .b(N545), .O(N2737) );
inv1 gate783( .a(N2658), .O(N2738) );
nand2 gate784( .a(N2661), .b(N546), .O(N2739) );
inv1 gate785( .a(N2661), .O(N2740) );
nand2 gate786( .a(N2664), .b(N547), .O(N2741) );
inv1 gate787( .a(N2664), .O(N2742) );
nand2 gate788( .a(N385), .b(N2689), .O(N2743) );
nand2 gate789( .a(N388), .b(N2691), .O(N2744) );
nand8 gate790( .a(N2537), .b(N2540), .c(N2543), .d(N2546), .e(N2594), .f(N2597), .g(N2600), .h(N2603), .O(N2745) );
nand8 gate791( .a(N2606), .b(N2549), .c(N2611), .d(N2614), .e(N2617), .f(N2620), .g(N2552), .h(N2555), .O(N2746) );
and8 gate792( .a(N2537), .b(N2540), .c(N2543), .d(N2546), .e(N2594), .f(N2597), .g(N2600), .h(N2603), .O(N2747) );
and8 gate793( .a(N2606), .b(N2549), .c(N2611), .d(N2614), .e(N2617), .f(N2620), .g(N2552), .h(N2555), .O(N2750) );
nand2 gate794( .a(N2669), .b(N2720), .O(N2753) );
nand2 gate795( .a(N2671), .b(N2721), .O(N2754) );

  xor2  gate1399(.a(N2722), .b(N2673), .O(gate796inter0));
  nand2 gate1400(.a(gate796inter0), .b(s_74), .O(gate796inter1));
  and2  gate1401(.a(N2722), .b(N2673), .O(gate796inter2));
  inv1  gate1402(.a(s_74), .O(gate796inter3));
  inv1  gate1403(.a(s_75), .O(gate796inter4));
  nand2 gate1404(.a(gate796inter4), .b(gate796inter3), .O(gate796inter5));
  nor2  gate1405(.a(gate796inter5), .b(gate796inter2), .O(gate796inter6));
  inv1  gate1406(.a(N2673), .O(gate796inter7));
  inv1  gate1407(.a(N2722), .O(gate796inter8));
  nand2 gate1408(.a(gate796inter8), .b(gate796inter7), .O(gate796inter9));
  nand2 gate1409(.a(s_75), .b(gate796inter3), .O(gate796inter10));
  nor2  gate1410(.a(gate796inter10), .b(gate796inter9), .O(gate796inter11));
  nor2  gate1411(.a(gate796inter11), .b(gate796inter6), .O(gate796inter12));
  nand2 gate1412(.a(gate796inter12), .b(gate796inter1), .O(N2755));
nand2 gate797( .a(N2675), .b(N2723), .O(N2756) );

  xor2  gate1049(.a(N2725), .b(N355), .O(gate798inter0));
  nand2 gate1050(.a(gate798inter0), .b(s_24), .O(gate798inter1));
  and2  gate1051(.a(N2725), .b(N355), .O(gate798inter2));
  inv1  gate1052(.a(s_24), .O(gate798inter3));
  inv1  gate1053(.a(s_25), .O(gate798inter4));
  nand2 gate1054(.a(gate798inter4), .b(gate798inter3), .O(gate798inter5));
  nor2  gate1055(.a(gate798inter5), .b(gate798inter2), .O(gate798inter6));
  inv1  gate1056(.a(N355), .O(gate798inter7));
  inv1  gate1057(.a(N2725), .O(gate798inter8));
  nand2 gate1058(.a(gate798inter8), .b(gate798inter7), .O(gate798inter9));
  nand2 gate1059(.a(s_25), .b(gate798inter3), .O(gate798inter10));
  nor2  gate1060(.a(gate798inter10), .b(gate798inter9), .O(gate798inter11));
  nor2  gate1061(.a(gate798inter11), .b(gate798inter6), .O(gate798inter12));
  nand2 gate1062(.a(gate798inter12), .b(gate798inter1), .O(N2757));
nand2 gate799( .a(N358), .b(N2727), .O(N2758) );

  xor2  gate1259(.a(N2729), .b(N361), .O(gate800inter0));
  nand2 gate1260(.a(gate800inter0), .b(s_54), .O(gate800inter1));
  and2  gate1261(.a(N2729), .b(N361), .O(gate800inter2));
  inv1  gate1262(.a(s_54), .O(gate800inter3));
  inv1  gate1263(.a(s_55), .O(gate800inter4));
  nand2 gate1264(.a(gate800inter4), .b(gate800inter3), .O(gate800inter5));
  nor2  gate1265(.a(gate800inter5), .b(gate800inter2), .O(gate800inter6));
  inv1  gate1266(.a(N361), .O(gate800inter7));
  inv1  gate1267(.a(N2729), .O(gate800inter8));
  nand2 gate1268(.a(gate800inter8), .b(gate800inter7), .O(gate800inter9));
  nand2 gate1269(.a(s_55), .b(gate800inter3), .O(gate800inter10));
  nor2  gate1270(.a(gate800inter10), .b(gate800inter9), .O(gate800inter11));
  nor2  gate1271(.a(gate800inter11), .b(gate800inter6), .O(gate800inter12));
  nand2 gate1272(.a(gate800inter12), .b(gate800inter1), .O(N2759));

  xor2  gate1987(.a(N2731), .b(N364), .O(gate801inter0));
  nand2 gate1988(.a(gate801inter0), .b(s_158), .O(gate801inter1));
  and2  gate1989(.a(N2731), .b(N364), .O(gate801inter2));
  inv1  gate1990(.a(s_158), .O(gate801inter3));
  inv1  gate1991(.a(s_159), .O(gate801inter4));
  nand2 gate1992(.a(gate801inter4), .b(gate801inter3), .O(gate801inter5));
  nor2  gate1993(.a(gate801inter5), .b(gate801inter2), .O(gate801inter6));
  inv1  gate1994(.a(N364), .O(gate801inter7));
  inv1  gate1995(.a(N2731), .O(gate801inter8));
  nand2 gate1996(.a(gate801inter8), .b(gate801inter7), .O(gate801inter9));
  nand2 gate1997(.a(s_159), .b(gate801inter3), .O(gate801inter10));
  nor2  gate1998(.a(gate801inter10), .b(gate801inter9), .O(gate801inter11));
  nor2  gate1999(.a(gate801inter11), .b(gate801inter6), .O(gate801inter12));
  nand2 gate2000(.a(gate801inter12), .b(gate801inter1), .O(N2760));
nand2 gate802( .a(N367), .b(N2733), .O(N2761) );
nand2 gate803( .a(N2682), .b(N2734), .O(N2762) );
nand2 gate804( .a(N373), .b(N2736), .O(N2763) );
nand2 gate805( .a(N376), .b(N2738), .O(N2764) );

  xor2  gate1973(.a(N2740), .b(N379), .O(gate806inter0));
  nand2 gate1974(.a(gate806inter0), .b(s_156), .O(gate806inter1));
  and2  gate1975(.a(N2740), .b(N379), .O(gate806inter2));
  inv1  gate1976(.a(s_156), .O(gate806inter3));
  inv1  gate1977(.a(s_157), .O(gate806inter4));
  nand2 gate1978(.a(gate806inter4), .b(gate806inter3), .O(gate806inter5));
  nor2  gate1979(.a(gate806inter5), .b(gate806inter2), .O(gate806inter6));
  inv1  gate1980(.a(N379), .O(gate806inter7));
  inv1  gate1981(.a(N2740), .O(gate806inter8));
  nand2 gate1982(.a(gate806inter8), .b(gate806inter7), .O(gate806inter9));
  nand2 gate1983(.a(s_157), .b(gate806inter3), .O(gate806inter10));
  nor2  gate1984(.a(gate806inter10), .b(gate806inter9), .O(gate806inter11));
  nor2  gate1985(.a(gate806inter11), .b(gate806inter6), .O(gate806inter12));
  nand2 gate1986(.a(gate806inter12), .b(gate806inter1), .O(N2765));
nand2 gate807( .a(N382), .b(N2742), .O(N2766) );
nand2 gate808( .a(N2688), .b(N2743), .O(N2767) );
nand2 gate809( .a(N2690), .b(N2744), .O(N2768) );
and2 gate810( .a(N2745), .b(N275), .O(N2773) );
and2 gate811( .a(N2746), .b(N276), .O(N2776) );

  xor2  gate1707(.a(N2757), .b(N2724), .O(gate812inter0));
  nand2 gate1708(.a(gate812inter0), .b(s_118), .O(gate812inter1));
  and2  gate1709(.a(N2757), .b(N2724), .O(gate812inter2));
  inv1  gate1710(.a(s_118), .O(gate812inter3));
  inv1  gate1711(.a(s_119), .O(gate812inter4));
  nand2 gate1712(.a(gate812inter4), .b(gate812inter3), .O(gate812inter5));
  nor2  gate1713(.a(gate812inter5), .b(gate812inter2), .O(gate812inter6));
  inv1  gate1714(.a(N2724), .O(gate812inter7));
  inv1  gate1715(.a(N2757), .O(gate812inter8));
  nand2 gate1716(.a(gate812inter8), .b(gate812inter7), .O(gate812inter9));
  nand2 gate1717(.a(s_119), .b(gate812inter3), .O(gate812inter10));
  nor2  gate1718(.a(gate812inter10), .b(gate812inter9), .O(gate812inter11));
  nor2  gate1719(.a(gate812inter11), .b(gate812inter6), .O(gate812inter12));
  nand2 gate1720(.a(gate812inter12), .b(gate812inter1), .O(N2779));
nand2 gate813( .a(N2726), .b(N2758), .O(N2780) );

  xor2  gate993(.a(N2759), .b(N2728), .O(gate814inter0));
  nand2 gate994(.a(gate814inter0), .b(s_16), .O(gate814inter1));
  and2  gate995(.a(N2759), .b(N2728), .O(gate814inter2));
  inv1  gate996(.a(s_16), .O(gate814inter3));
  inv1  gate997(.a(s_17), .O(gate814inter4));
  nand2 gate998(.a(gate814inter4), .b(gate814inter3), .O(gate814inter5));
  nor2  gate999(.a(gate814inter5), .b(gate814inter2), .O(gate814inter6));
  inv1  gate1000(.a(N2728), .O(gate814inter7));
  inv1  gate1001(.a(N2759), .O(gate814inter8));
  nand2 gate1002(.a(gate814inter8), .b(gate814inter7), .O(gate814inter9));
  nand2 gate1003(.a(s_17), .b(gate814inter3), .O(gate814inter10));
  nor2  gate1004(.a(gate814inter10), .b(gate814inter9), .O(gate814inter11));
  nor2  gate1005(.a(gate814inter11), .b(gate814inter6), .O(gate814inter12));
  nand2 gate1006(.a(gate814inter12), .b(gate814inter1), .O(N2781));
nand2 gate815( .a(N2730), .b(N2760), .O(N2782) );
nand2 gate816( .a(N2732), .b(N2761), .O(N2783) );
nand2 gate817( .a(N2735), .b(N2763), .O(N2784) );

  xor2  gate1553(.a(N2764), .b(N2737), .O(gate818inter0));
  nand2 gate1554(.a(gate818inter0), .b(s_96), .O(gate818inter1));
  and2  gate1555(.a(N2764), .b(N2737), .O(gate818inter2));
  inv1  gate1556(.a(s_96), .O(gate818inter3));
  inv1  gate1557(.a(s_97), .O(gate818inter4));
  nand2 gate1558(.a(gate818inter4), .b(gate818inter3), .O(gate818inter5));
  nor2  gate1559(.a(gate818inter5), .b(gate818inter2), .O(gate818inter6));
  inv1  gate1560(.a(N2737), .O(gate818inter7));
  inv1  gate1561(.a(N2764), .O(gate818inter8));
  nand2 gate1562(.a(gate818inter8), .b(gate818inter7), .O(gate818inter9));
  nand2 gate1563(.a(s_97), .b(gate818inter3), .O(gate818inter10));
  nor2  gate1564(.a(gate818inter10), .b(gate818inter9), .O(gate818inter11));
  nor2  gate1565(.a(gate818inter11), .b(gate818inter6), .O(gate818inter12));
  nand2 gate1566(.a(gate818inter12), .b(gate818inter1), .O(N2785));
nand2 gate819( .a(N2739), .b(N2765), .O(N2786) );
nand2 gate820( .a(N2741), .b(N2766), .O(N2787) );
and3 gate821( .a(N2747), .b(N2750), .c(N2710), .O(N2788) );
nand2 gate822( .a(N2747), .b(N2750), .O(N2789) );
and4 gate823( .a(N338), .b(N2279), .c(N99), .d(N2788), .O(N2800) );
nand2 gate824( .a(N2773), .b(N2018), .O(N2807) );
inv1 gate825( .a(N2773), .O(N2808) );

  xor2  gate1637(.a(N2019), .b(N2776), .O(gate826inter0));
  nand2 gate1638(.a(gate826inter0), .b(s_108), .O(gate826inter1));
  and2  gate1639(.a(N2019), .b(N2776), .O(gate826inter2));
  inv1  gate1640(.a(s_108), .O(gate826inter3));
  inv1  gate1641(.a(s_109), .O(gate826inter4));
  nand2 gate1642(.a(gate826inter4), .b(gate826inter3), .O(gate826inter5));
  nor2  gate1643(.a(gate826inter5), .b(gate826inter2), .O(gate826inter6));
  inv1  gate1644(.a(N2776), .O(gate826inter7));
  inv1  gate1645(.a(N2019), .O(gate826inter8));
  nand2 gate1646(.a(gate826inter8), .b(gate826inter7), .O(gate826inter9));
  nand2 gate1647(.a(s_109), .b(gate826inter3), .O(gate826inter10));
  nor2  gate1648(.a(gate826inter10), .b(gate826inter9), .O(gate826inter11));
  nor2  gate1649(.a(gate826inter11), .b(gate826inter6), .O(gate826inter12));
  nand2 gate1650(.a(gate826inter12), .b(gate826inter1), .O(N2809));
inv1 gate827( .a(N2776), .O(N2810) );
nor2 gate828( .a(N2384), .b(N2800), .O(N2811) );
and3 gate829( .a(N897), .b(N283), .c(N2789), .O(N2812) );
and3 gate830( .a(N76), .b(N283), .c(N2789), .O(N2815) );
and3 gate831( .a(N82), .b(N283), .c(N2789), .O(N2818) );
and3 gate832( .a(N85), .b(N283), .c(N2789), .O(N2821) );
and3 gate833( .a(N898), .b(N283), .c(N2789), .O(N2824) );
nand2 gate834( .a(N1965), .b(N2808), .O(N2827) );
nand2 gate835( .a(N1968), .b(N2810), .O(N2828) );
and3 gate836( .a(N79), .b(N283), .c(N2789), .O(N2829) );
nand2 gate837( .a(N2807), .b(N2827), .O(N2843) );
nand2 gate838( .a(N2809), .b(N2828), .O(N2846) );

  xor2  gate895(.a(N2076), .b(N2812), .O(gate839inter0));
  nand2 gate896(.a(gate839inter0), .b(s_2), .O(gate839inter1));
  and2  gate897(.a(N2076), .b(N2812), .O(gate839inter2));
  inv1  gate898(.a(s_2), .O(gate839inter3));
  inv1  gate899(.a(s_3), .O(gate839inter4));
  nand2 gate900(.a(gate839inter4), .b(gate839inter3), .O(gate839inter5));
  nor2  gate901(.a(gate839inter5), .b(gate839inter2), .O(gate839inter6));
  inv1  gate902(.a(N2812), .O(gate839inter7));
  inv1  gate903(.a(N2076), .O(gate839inter8));
  nand2 gate904(.a(gate839inter8), .b(gate839inter7), .O(gate839inter9));
  nand2 gate905(.a(s_3), .b(gate839inter3), .O(gate839inter10));
  nor2  gate906(.a(gate839inter10), .b(gate839inter9), .O(gate839inter11));
  nor2  gate907(.a(gate839inter11), .b(gate839inter6), .O(gate839inter12));
  nand2 gate908(.a(gate839inter12), .b(gate839inter1), .O(N2850));

  xor2  gate1077(.a(N2077), .b(N2815), .O(gate840inter0));
  nand2 gate1078(.a(gate840inter0), .b(s_28), .O(gate840inter1));
  and2  gate1079(.a(N2077), .b(N2815), .O(gate840inter2));
  inv1  gate1080(.a(s_28), .O(gate840inter3));
  inv1  gate1081(.a(s_29), .O(gate840inter4));
  nand2 gate1082(.a(gate840inter4), .b(gate840inter3), .O(gate840inter5));
  nor2  gate1083(.a(gate840inter5), .b(gate840inter2), .O(gate840inter6));
  inv1  gate1084(.a(N2815), .O(gate840inter7));
  inv1  gate1085(.a(N2077), .O(gate840inter8));
  nand2 gate1086(.a(gate840inter8), .b(gate840inter7), .O(gate840inter9));
  nand2 gate1087(.a(s_29), .b(gate840inter3), .O(gate840inter10));
  nor2  gate1088(.a(gate840inter10), .b(gate840inter9), .O(gate840inter11));
  nor2  gate1089(.a(gate840inter11), .b(gate840inter6), .O(gate840inter12));
  nand2 gate1090(.a(gate840inter12), .b(gate840inter1), .O(N2851));
nand2 gate841( .a(N2818), .b(N1915), .O(N2852) );
nand2 gate842( .a(N2821), .b(N1857), .O(N2853) );
nand2 gate843( .a(N2824), .b(N1938), .O(N2854) );
inv1 gate844( .a(N2812), .O(N2857) );
inv1 gate845( .a(N2815), .O(N2858) );
inv1 gate846( .a(N2818), .O(N2859) );
inv1 gate847( .a(N2821), .O(N2860) );
inv1 gate848( .a(N2824), .O(N2861) );
inv1 gate849( .a(N2829), .O(N2862) );
nand2 gate850( .a(N2829), .b(N1985), .O(N2863) );
nand2 gate851( .a(N2052), .b(N2857), .O(N2866) );

  xor2  gate1889(.a(N2858), .b(N2055), .O(gate852inter0));
  nand2 gate1890(.a(gate852inter0), .b(s_144), .O(gate852inter1));
  and2  gate1891(.a(N2858), .b(N2055), .O(gate852inter2));
  inv1  gate1892(.a(s_144), .O(gate852inter3));
  inv1  gate1893(.a(s_145), .O(gate852inter4));
  nand2 gate1894(.a(gate852inter4), .b(gate852inter3), .O(gate852inter5));
  nor2  gate1895(.a(gate852inter5), .b(gate852inter2), .O(gate852inter6));
  inv1  gate1896(.a(N2055), .O(gate852inter7));
  inv1  gate1897(.a(N2858), .O(gate852inter8));
  nand2 gate1898(.a(gate852inter8), .b(gate852inter7), .O(gate852inter9));
  nand2 gate1899(.a(s_145), .b(gate852inter3), .O(gate852inter10));
  nor2  gate1900(.a(gate852inter10), .b(gate852inter9), .O(gate852inter11));
  nor2  gate1901(.a(gate852inter11), .b(gate852inter6), .O(gate852inter12));
  nand2 gate1902(.a(gate852inter12), .b(gate852inter1), .O(N2867));
nand2 gate853( .a(N1866), .b(N2859), .O(N2868) );

  xor2  gate1287(.a(N2860), .b(N1818), .O(gate854inter0));
  nand2 gate1288(.a(gate854inter0), .b(s_58), .O(gate854inter1));
  and2  gate1289(.a(N2860), .b(N1818), .O(gate854inter2));
  inv1  gate1290(.a(s_58), .O(gate854inter3));
  inv1  gate1291(.a(s_59), .O(gate854inter4));
  nand2 gate1292(.a(gate854inter4), .b(gate854inter3), .O(gate854inter5));
  nor2  gate1293(.a(gate854inter5), .b(gate854inter2), .O(gate854inter6));
  inv1  gate1294(.a(N1818), .O(gate854inter7));
  inv1  gate1295(.a(N2860), .O(gate854inter8));
  nand2 gate1296(.a(gate854inter8), .b(gate854inter7), .O(gate854inter9));
  nand2 gate1297(.a(s_59), .b(gate854inter3), .O(gate854inter10));
  nor2  gate1298(.a(gate854inter10), .b(gate854inter9), .O(gate854inter11));
  nor2  gate1299(.a(gate854inter11), .b(gate854inter6), .O(gate854inter12));
  nand2 gate1300(.a(gate854inter12), .b(gate854inter1), .O(N2869));
nand2 gate855( .a(N1902), .b(N2861), .O(N2870) );

  xor2  gate1119(.a(N886), .b(N2843), .O(gate856inter0));
  nand2 gate1120(.a(gate856inter0), .b(s_34), .O(gate856inter1));
  and2  gate1121(.a(N886), .b(N2843), .O(gate856inter2));
  inv1  gate1122(.a(s_34), .O(gate856inter3));
  inv1  gate1123(.a(s_35), .O(gate856inter4));
  nand2 gate1124(.a(gate856inter4), .b(gate856inter3), .O(gate856inter5));
  nor2  gate1125(.a(gate856inter5), .b(gate856inter2), .O(gate856inter6));
  inv1  gate1126(.a(N2843), .O(gate856inter7));
  inv1  gate1127(.a(N886), .O(gate856inter8));
  nand2 gate1128(.a(gate856inter8), .b(gate856inter7), .O(gate856inter9));
  nand2 gate1129(.a(s_35), .b(gate856inter3), .O(gate856inter10));
  nor2  gate1130(.a(gate856inter10), .b(gate856inter9), .O(gate856inter11));
  nor2  gate1131(.a(gate856inter11), .b(gate856inter6), .O(gate856inter12));
  nand2 gate1132(.a(gate856inter12), .b(gate856inter1), .O(N2871));
inv1 gate857( .a(N2843), .O(N2872) );
nand2 gate858( .a(N2846), .b(N887), .O(N2873) );
inv1 gate859( .a(N2846), .O(N2874) );
nand2 gate860( .a(N1933), .b(N2862), .O(N2875) );
nand2 gate861( .a(N2866), .b(N2850), .O(N2876) );
nand2 gate862( .a(N2867), .b(N2851), .O(N2877) );
nand2 gate863( .a(N2868), .b(N2852), .O(N2878) );

  xor2  gate1903(.a(N2853), .b(N2869), .O(gate864inter0));
  nand2 gate1904(.a(gate864inter0), .b(s_146), .O(gate864inter1));
  and2  gate1905(.a(N2853), .b(N2869), .O(gate864inter2));
  inv1  gate1906(.a(s_146), .O(gate864inter3));
  inv1  gate1907(.a(s_147), .O(gate864inter4));
  nand2 gate1908(.a(gate864inter4), .b(gate864inter3), .O(gate864inter5));
  nor2  gate1909(.a(gate864inter5), .b(gate864inter2), .O(gate864inter6));
  inv1  gate1910(.a(N2869), .O(gate864inter7));
  inv1  gate1911(.a(N2853), .O(gate864inter8));
  nand2 gate1912(.a(gate864inter8), .b(gate864inter7), .O(gate864inter9));
  nand2 gate1913(.a(s_147), .b(gate864inter3), .O(gate864inter10));
  nor2  gate1914(.a(gate864inter10), .b(gate864inter9), .O(gate864inter11));
  nor2  gate1915(.a(gate864inter11), .b(gate864inter6), .O(gate864inter12));
  nand2 gate1916(.a(gate864inter12), .b(gate864inter1), .O(N2879));
nand2 gate865( .a(N2870), .b(N2854), .O(N2880) );
nand2 gate866( .a(N682), .b(N2872), .O(N2881) );
nand2 gate867( .a(N685), .b(N2874), .O(N2882) );
nand2 gate868( .a(N2875), .b(N2863), .O(N2883) );
and2 gate869( .a(N2876), .b(N550), .O(N2886) );
and2 gate870( .a(N551), .b(N2877), .O(N2887) );
and2 gate871( .a(N553), .b(N2878), .O(N2888) );
and2 gate872( .a(N2879), .b(N554), .O(N2889) );
and2 gate873( .a(N555), .b(N2880), .O(N2890) );
nand2 gate874( .a(N2871), .b(N2881), .O(N2891) );
nand2 gate875( .a(N2873), .b(N2882), .O(N2892) );

  xor2  gate1735(.a(N1461), .b(N2883), .O(gate876inter0));
  nand2 gate1736(.a(gate876inter0), .b(s_122), .O(gate876inter1));
  and2  gate1737(.a(N1461), .b(N2883), .O(gate876inter2));
  inv1  gate1738(.a(s_122), .O(gate876inter3));
  inv1  gate1739(.a(s_123), .O(gate876inter4));
  nand2 gate1740(.a(gate876inter4), .b(gate876inter3), .O(gate876inter5));
  nor2  gate1741(.a(gate876inter5), .b(gate876inter2), .O(gate876inter6));
  inv1  gate1742(.a(N2883), .O(gate876inter7));
  inv1  gate1743(.a(N1461), .O(gate876inter8));
  nand2 gate1744(.a(gate876inter8), .b(gate876inter7), .O(gate876inter9));
  nand2 gate1745(.a(s_123), .b(gate876inter3), .O(gate876inter10));
  nor2  gate1746(.a(gate876inter10), .b(gate876inter9), .O(gate876inter11));
  nor2  gate1747(.a(gate876inter11), .b(gate876inter6), .O(gate876inter12));
  nand2 gate1748(.a(gate876inter12), .b(gate876inter1), .O(N2895));
inv1 gate877( .a(N2883), .O(N2896) );

  xor2  gate1469(.a(N2896), .b(N1383), .O(gate878inter0));
  nand2 gate1470(.a(gate878inter0), .b(s_84), .O(gate878inter1));
  and2  gate1471(.a(N2896), .b(N1383), .O(gate878inter2));
  inv1  gate1472(.a(s_84), .O(gate878inter3));
  inv1  gate1473(.a(s_85), .O(gate878inter4));
  nand2 gate1474(.a(gate878inter4), .b(gate878inter3), .O(gate878inter5));
  nor2  gate1475(.a(gate878inter5), .b(gate878inter2), .O(gate878inter6));
  inv1  gate1476(.a(N1383), .O(gate878inter7));
  inv1  gate1477(.a(N2896), .O(gate878inter8));
  nand2 gate1478(.a(gate878inter8), .b(gate878inter7), .O(gate878inter9));
  nand2 gate1479(.a(s_85), .b(gate878inter3), .O(gate878inter10));
  nor2  gate1480(.a(gate878inter10), .b(gate878inter9), .O(gate878inter11));
  nor2  gate1481(.a(gate878inter11), .b(gate878inter6), .O(gate878inter12));
  nand2 gate1482(.a(gate878inter12), .b(gate878inter1), .O(N2897));
nand2 gate879( .a(N2895), .b(N2897), .O(N2898) );
and2 gate880( .a(N2898), .b(N552), .O(N2899) );

endmodule