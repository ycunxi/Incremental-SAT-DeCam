module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);

input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;//RE__PI;

input s_0,s_1;//RE__ALLOW(00,01,10,11);
input s_2,s_3;//RE__ALLOW(00,01,10,11);
input s_4,s_5;//RE__ALLOW(00,01,10,11);
input s_6,s_7;//RE__ALLOW(00,01,10,11);
input s_8,s_9;//RE__ALLOW(00,01,10,11);
input s_10,s_11;//RE__ALLOW(00,01,10,11);
input s_12,s_13;//RE__ALLOW(00,01,10,11);
input s_14,s_15;//RE__ALLOW(00,01,10,11);
input s_16,s_17;//RE__ALLOW(00,01,10,11);
input s_18,s_19;//RE__ALLOW(00,01,10,11);
input s_20,s_21;//RE__ALLOW(00,01,10,11);
input s_22,s_23;//RE__ALLOW(00,01,10,11);
input s_24,s_25;//RE__ALLOW(00,01,10,11);
input s_26,s_27;//RE__ALLOW(00,01,10,11);
input s_28,s_29;//RE__ALLOW(00,01,10,11);
input s_30,s_31;//RE__ALLOW(00,01,10,11);
input s_32,s_33;//RE__ALLOW(00,01,10,11);
input s_34,s_35;//RE__ALLOW(00,01,10,11);
input s_36,s_37;//RE__ALLOW(00,01,10,11);
input s_38,s_39;//RE__ALLOW(00,01,10,11);
input s_40,s_41;//RE__ALLOW(00,01,10,11);
input s_42,s_43;//RE__ALLOW(00,01,10,11);
input s_44,s_45;//RE__ALLOW(00,01,10,11);
input s_46,s_47;//RE__ALLOW(00,01,10,11);
input s_48,s_49;//RE__ALLOW(00,01,10,11);
input s_50,s_51;//RE__ALLOW(00,01,10,11);
input s_52,s_53;//RE__ALLOW(00,01,10,11);
input s_54,s_55;//RE__ALLOW(00,01,10,11);
input s_56,s_57;//RE__ALLOW(00,01,10,11);
input s_58,s_59;//RE__ALLOW(00,01,10,11);
input s_60,s_61;//RE__ALLOW(00,01,10,11);
input s_62,s_63;//RE__ALLOW(00,01,10,11);
input s_64,s_65;//RE__ALLOW(00,01,10,11);
input s_66,s_67;//RE__ALLOW(00,01,10,11);
input s_68,s_69;//RE__ALLOW(00,01,10,11);
input s_70,s_71;//RE__ALLOW(00,01,10,11);
input s_72,s_73;//RE__ALLOW(00,01,10,11);
input s_74,s_75;//RE__ALLOW(00,01,10,11);
input s_76,s_77;//RE__ALLOW(00,01,10,11);
input s_78,s_79;//RE__ALLOW(00,01,10,11);
input s_80,s_81;//RE__ALLOW(00,01,10,11);
input s_82,s_83;//RE__ALLOW(00,01,10,11);
input s_84,s_85;//RE__ALLOW(00,01,10,11);
input s_86,s_87;//RE__ALLOW(00,01,10,11);
input s_88,s_89;//RE__ALLOW(00,01,10,11);
input s_90,s_91;//RE__ALLOW(00,01,10,11);
input s_92,s_93;//RE__ALLOW(00,01,10,11);
input s_94,s_95;//RE__ALLOW(00,01,10,11);
input s_96,s_97;//RE__ALLOW(00,01,10,11);
input s_98,s_99;//RE__ALLOW(00,01,10,11);
input s_100,s_101;//RE__ALLOW(00,01,10,11);
input s_102,s_103;//RE__ALLOW(00,01,10,11);
input s_104,s_105;//RE__ALLOW(00,01,10,11);
input s_106,s_107;//RE__ALLOW(00,01,10,11);
input s_108,s_109;//RE__ALLOW(00,01,10,11);
input s_110,s_111;//RE__ALLOW(00,01,10,11);
input s_112,s_113;//RE__ALLOW(00,01,10,11);
input s_114,s_115;//RE__ALLOW(00,01,10,11);
input s_116,s_117;//RE__ALLOW(00,01,10,11);
input s_118,s_119;//RE__ALLOW(00,01,10,11);
input s_120,s_121;//RE__ALLOW(00,01,10,11);
input s_122,s_123;//RE__ALLOW(00,01,10,11);
input s_124,s_125;//RE__ALLOW(00,01,10,11);
input s_126,s_127;//RE__ALLOW(00,01,10,11);
input s_128,s_129;//RE__ALLOW(00,01,10,11);
input s_130,s_131;//RE__ALLOW(00,01,10,11);
input s_132,s_133;//RE__ALLOW(00,01,10,11);
input s_134,s_135;//RE__ALLOW(00,01,10,11);
input s_136,s_137;//RE__ALLOW(00,01,10,11);
input s_138,s_139;//RE__ALLOW(00,01,10,11);
input s_140,s_141;//RE__ALLOW(00,01,10,11);
input s_142,s_143;//RE__ALLOW(00,01,10,11);
input s_144,s_145;//RE__ALLOW(00,01,10,11);
input s_146,s_147;//RE__ALLOW(00,01,10,11);
input s_148,s_149;//RE__ALLOW(00,01,10,11);
input s_150,s_151;//RE__ALLOW(00,01,10,11);
input s_152,s_153;//RE__ALLOW(00,01,10,11);
input s_154,s_155;//RE__ALLOW(00,01,10,11);
input s_156,s_157;//RE__ALLOW(00,01,10,11);
input s_158,s_159;//RE__ALLOW(00,01,10,11);
input s_160,s_161;//RE__ALLOW(00,01,10,11);
input s_162,s_163;//RE__ALLOW(00,01,10,11);
input s_164,s_165;//RE__ALLOW(00,01,10,11);
input s_166,s_167;//RE__ALLOW(00,01,10,11);
input s_168,s_169;//RE__ALLOW(00,01,10,11);
input s_170,s_171;//RE__ALLOW(00,01,10,11);
input s_172,s_173;//RE__ALLOW(00,01,10,11);
input s_174,s_175;//RE__ALLOW(00,01,10,11);
input s_176,s_177;//RE__ALLOW(00,01,10,11);
input s_178,s_179;//RE__ALLOW(00,01,10,11);
input s_180,s_181;//RE__ALLOW(00,01,10,11);
input s_182,s_183;//RE__ALLOW(00,01,10,11);
input s_184,s_185;//RE__ALLOW(00,01,10,11);
input s_186,s_187;//RE__ALLOW(00,01,10,11);
input s_188,s_189;//RE__ALLOW(00,01,10,11);
input s_190,s_191;//RE__ALLOW(00,01,10,11);
input s_192,s_193;//RE__ALLOW(00,01,10,11);
input s_194,s_195;//RE__ALLOW(00,01,10,11);
input s_196,s_197;//RE__ALLOW(00,01,10,11);
input s_198,s_199;//RE__ALLOW(00,01,10,11);
input s_200,s_201;//RE__ALLOW(00,01,10,11);
input s_202,s_203;//RE__ALLOW(00,01,10,11);
input s_204,s_205;//RE__ALLOW(00,01,10,11);
input s_206,s_207;//RE__ALLOW(00,01,10,11);
input s_208,s_209;//RE__ALLOW(00,01,10,11);
input s_210,s_211;//RE__ALLOW(00,01,10,11);
input s_212,s_213;//RE__ALLOW(00,01,10,11);
input s_214,s_215;//RE__ALLOW(00,01,10,11);
input s_216,s_217;//RE__ALLOW(00,01,10,11);
input s_218,s_219;//RE__ALLOW(00,01,10,11);
input s_220,s_221;//RE__ALLOW(00,01,10,11);
input s_222,s_223;//RE__ALLOW(00,01,10,11);
input s_224,s_225;//RE__ALLOW(00,01,10,11);
input s_226,s_227;//RE__ALLOW(00,01,10,11);
input s_228,s_229;//RE__ALLOW(00,01,10,11);
input s_230,s_231;//RE__ALLOW(00,01,10,11);
input s_232,s_233;//RE__ALLOW(00,01,10,11);
input s_234,s_235;//RE__ALLOW(00,01,10,11);
input s_236,s_237;//RE__ALLOW(00,01,10,11);
input s_238,s_239;//RE__ALLOW(00,01,10,11);
input s_240,s_241;//RE__ALLOW(00,01,10,11);
input s_242,s_243;//RE__ALLOW(00,01,10,11);
input s_244,s_245;//RE__ALLOW(00,01,10,11);
input s_246,s_247;//RE__ALLOW(00,01,10,11);
input s_248,s_249;//RE__ALLOW(00,01,10,11);
input s_250,s_251;//RE__ALLOW(00,01,10,11);
input s_252,s_253;//RE__ALLOW(00,01,10,11);
input s_254,s_255;//RE__ALLOW(00,01,10,11);
input s_256,s_257;//RE__ALLOW(00,01,10,11);
input s_258,s_259;//RE__ALLOW(00,01,10,11);
input s_260,s_261;//RE__ALLOW(00,01,10,11);
input s_262,s_263;//RE__ALLOW(00,01,10,11);
input s_264,s_265;//RE__ALLOW(00,01,10,11);
input s_266,s_267;//RE__ALLOW(00,01,10,11);
input s_268,s_269;//RE__ALLOW(00,01,10,11);
input s_270,s_271;//RE__ALLOW(00,01,10,11);
input s_272,s_273;//RE__ALLOW(00,01,10,11);
input s_274,s_275;//RE__ALLOW(00,01,10,11);
input s_276,s_277;//RE__ALLOW(00,01,10,11);
input s_278,s_279;//RE__ALLOW(00,01,10,11);
input s_280,s_281;//RE__ALLOW(00,01,10,11);
input s_282,s_283;//RE__ALLOW(00,01,10,11);
input s_284,s_285;//RE__ALLOW(00,01,10,11);
input s_286,s_287;//RE__ALLOW(00,01,10,11);
input s_288,s_289;//RE__ALLOW(00,01,10,11);
input s_290,s_291;//RE__ALLOW(00,01,10,11);
input s_292,s_293;//RE__ALLOW(00,01,10,11);
input s_294,s_295;//RE__ALLOW(00,01,10,11);
input s_296,s_297;//RE__ALLOW(00,01,10,11);
input s_298,s_299;//RE__ALLOW(00,01,10,11);
input s_300,s_301;//RE__ALLOW(00,01,10,11);
input s_302,s_303;//RE__ALLOW(00,01,10,11);
input s_304,s_305;//RE__ALLOW(00,01,10,11);
input s_306,s_307;//RE__ALLOW(00,01,10,11);
input s_308,s_309;//RE__ALLOW(00,01,10,11);
input s_310,s_311;//RE__ALLOW(00,01,10,11);
input s_312,s_313;//RE__ALLOW(00,01,10,11);
input s_314,s_315;//RE__ALLOW(00,01,10,11);
input s_316,s_317;//RE__ALLOW(00,01,10,11);
input s_318,s_319;//RE__ALLOW(00,01,10,11);
input s_320,s_321;//RE__ALLOW(00,01,10,11);
input s_322,s_323;//RE__ALLOW(00,01,10,11);
input s_324,s_325;//RE__ALLOW(00,01,10,11);
input s_326,s_327;//RE__ALLOW(00,01,10,11);
input s_328,s_329;//RE__ALLOW(00,01,10,11);
input s_330,s_331;//RE__ALLOW(00,01,10,11);
input s_332,s_333;//RE__ALLOW(00,01,10,11);
input s_334,s_335;//RE__ALLOW(00,01,10,11);
input s_336,s_337;//RE__ALLOW(00,01,10,11);
input s_338,s_339;//RE__ALLOW(00,01,10,11);
input s_340,s_341;//RE__ALLOW(00,01,10,11);
input s_342,s_343;//RE__ALLOW(00,01,10,11);
input s_344,s_345;//RE__ALLOW(00,01,10,11);
input s_346,s_347;//RE__ALLOW(00,01,10,11);
input s_348,s_349;//RE__ALLOW(00,01,10,11);
input s_350,s_351;//RE__ALLOW(00,01,10,11);
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;

  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate125inter0, gate125inter1, gate125inter2, gate125inter3, gate125inter4, gate125inter5, gate125inter6, gate125inter7, gate125inter8, gate125inter9, gate125inter10, gate125inter11, gate125inter12, gate210inter0, gate210inter1, gate210inter2, gate210inter3, gate210inter4, gate210inter5, gate210inter6, gate210inter7, gate210inter8, gate210inter9, gate210inter10, gate210inter11, gate210inter12, gate294inter0, gate294inter1, gate294inter2, gate294inter3, gate294inter4, gate294inter5, gate294inter6, gate294inter7, gate294inter8, gate294inter9, gate294inter10, gate294inter11, gate294inter12, gate127inter0, gate127inter1, gate127inter2, gate127inter3, gate127inter4, gate127inter5, gate127inter6, gate127inter7, gate127inter8, gate127inter9, gate127inter10, gate127inter11, gate127inter12, gate292inter0, gate292inter1, gate292inter2, gate292inter3, gate292inter4, gate292inter5, gate292inter6, gate292inter7, gate292inter8, gate292inter9, gate292inter10, gate292inter11, gate292inter12, gate231inter0, gate231inter1, gate231inter2, gate231inter3, gate231inter4, gate231inter5, gate231inter6, gate231inter7, gate231inter8, gate231inter9, gate231inter10, gate231inter11, gate231inter12, gate284inter0, gate284inter1, gate284inter2, gate284inter3, gate284inter4, gate284inter5, gate284inter6, gate284inter7, gate284inter8, gate284inter9, gate284inter10, gate284inter11, gate284inter12, gate196inter0, gate196inter1, gate196inter2, gate196inter3, gate196inter4, gate196inter5, gate196inter6, gate196inter7, gate196inter8, gate196inter9, gate196inter10, gate196inter11, gate196inter12, gate400inter0, gate400inter1, gate400inter2, gate400inter3, gate400inter4, gate400inter5, gate400inter6, gate400inter7, gate400inter8, gate400inter9, gate400inter10, gate400inter11, gate400inter12, gate514inter0, gate514inter1, gate514inter2, gate514inter3, gate514inter4, gate514inter5, gate514inter6, gate514inter7, gate514inter8, gate514inter9, gate514inter10, gate514inter11, gate514inter12, gate413inter0, gate413inter1, gate413inter2, gate413inter3, gate413inter4, gate413inter5, gate413inter6, gate413inter7, gate413inter8, gate413inter9, gate413inter10, gate413inter11, gate413inter12, gate266inter0, gate266inter1, gate266inter2, gate266inter3, gate266inter4, gate266inter5, gate266inter6, gate266inter7, gate266inter8, gate266inter9, gate266inter10, gate266inter11, gate266inter12, gate296inter0, gate296inter1, gate296inter2, gate296inter3, gate296inter4, gate296inter5, gate296inter6, gate296inter7, gate296inter8, gate296inter9, gate296inter10, gate296inter11, gate296inter12, gate147inter0, gate147inter1, gate147inter2, gate147inter3, gate147inter4, gate147inter5, gate147inter6, gate147inter7, gate147inter8, gate147inter9, gate147inter10, gate147inter11, gate147inter12, gate457inter0, gate457inter1, gate457inter2, gate457inter3, gate457inter4, gate457inter5, gate457inter6, gate457inter7, gate457inter8, gate457inter9, gate457inter10, gate457inter11, gate457inter12, gate280inter0, gate280inter1, gate280inter2, gate280inter3, gate280inter4, gate280inter5, gate280inter6, gate280inter7, gate280inter8, gate280inter9, gate280inter10, gate280inter11, gate280inter12, gate408inter0, gate408inter1, gate408inter2, gate408inter3, gate408inter4, gate408inter5, gate408inter6, gate408inter7, gate408inter8, gate408inter9, gate408inter10, gate408inter11, gate408inter12, gate53inter0, gate53inter1, gate53inter2, gate53inter3, gate53inter4, gate53inter5, gate53inter6, gate53inter7, gate53inter8, gate53inter9, gate53inter10, gate53inter11, gate53inter12, gate174inter0, gate174inter1, gate174inter2, gate174inter3, gate174inter4, gate174inter5, gate174inter6, gate174inter7, gate174inter8, gate174inter9, gate174inter10, gate174inter11, gate174inter12, gate387inter0, gate387inter1, gate387inter2, gate387inter3, gate387inter4, gate387inter5, gate387inter6, gate387inter7, gate387inter8, gate387inter9, gate387inter10, gate387inter11, gate387inter12, gate162inter0, gate162inter1, gate162inter2, gate162inter3, gate162inter4, gate162inter5, gate162inter6, gate162inter7, gate162inter8, gate162inter9, gate162inter10, gate162inter11, gate162inter12, gate209inter0, gate209inter1, gate209inter2, gate209inter3, gate209inter4, gate209inter5, gate209inter6, gate209inter7, gate209inter8, gate209inter9, gate209inter10, gate209inter11, gate209inter12, gate405inter0, gate405inter1, gate405inter2, gate405inter3, gate405inter4, gate405inter5, gate405inter6, gate405inter7, gate405inter8, gate405inter9, gate405inter10, gate405inter11, gate405inter12, gate410inter0, gate410inter1, gate410inter2, gate410inter3, gate410inter4, gate410inter5, gate410inter6, gate410inter7, gate410inter8, gate410inter9, gate410inter10, gate410inter11, gate410inter12, gate155inter0, gate155inter1, gate155inter2, gate155inter3, gate155inter4, gate155inter5, gate155inter6, gate155inter7, gate155inter8, gate155inter9, gate155inter10, gate155inter11, gate155inter12, gate16inter0, gate16inter1, gate16inter2, gate16inter3, gate16inter4, gate16inter5, gate16inter6, gate16inter7, gate16inter8, gate16inter9, gate16inter10, gate16inter11, gate16inter12, gate97inter0, gate97inter1, gate97inter2, gate97inter3, gate97inter4, gate97inter5, gate97inter6, gate97inter7, gate97inter8, gate97inter9, gate97inter10, gate97inter11, gate97inter12, gate260inter0, gate260inter1, gate260inter2, gate260inter3, gate260inter4, gate260inter5, gate260inter6, gate260inter7, gate260inter8, gate260inter9, gate260inter10, gate260inter11, gate260inter12, gate197inter0, gate197inter1, gate197inter2, gate197inter3, gate197inter4, gate197inter5, gate197inter6, gate197inter7, gate197inter8, gate197inter9, gate197inter10, gate197inter11, gate197inter12, gate443inter0, gate443inter1, gate443inter2, gate443inter3, gate443inter4, gate443inter5, gate443inter6, gate443inter7, gate443inter8, gate443inter9, gate443inter10, gate443inter11, gate443inter12, gate129inter0, gate129inter1, gate129inter2, gate129inter3, gate129inter4, gate129inter5, gate129inter6, gate129inter7, gate129inter8, gate129inter9, gate129inter10, gate129inter11, gate129inter12, gate78inter0, gate78inter1, gate78inter2, gate78inter3, gate78inter4, gate78inter5, gate78inter6, gate78inter7, gate78inter8, gate78inter9, gate78inter10, gate78inter11, gate78inter12, gate180inter0, gate180inter1, gate180inter2, gate180inter3, gate180inter4, gate180inter5, gate180inter6, gate180inter7, gate180inter8, gate180inter9, gate180inter10, gate180inter11, gate180inter12, gate32inter0, gate32inter1, gate32inter2, gate32inter3, gate32inter4, gate32inter5, gate32inter6, gate32inter7, gate32inter8, gate32inter9, gate32inter10, gate32inter11, gate32inter12, gate109inter0, gate109inter1, gate109inter2, gate109inter3, gate109inter4, gate109inter5, gate109inter6, gate109inter7, gate109inter8, gate109inter9, gate109inter10, gate109inter11, gate109inter12, gate248inter0, gate248inter1, gate248inter2, gate248inter3, gate248inter4, gate248inter5, gate248inter6, gate248inter7, gate248inter8, gate248inter9, gate248inter10, gate248inter11, gate248inter12, gate490inter0, gate490inter1, gate490inter2, gate490inter3, gate490inter4, gate490inter5, gate490inter6, gate490inter7, gate490inter8, gate490inter9, gate490inter10, gate490inter11, gate490inter12, gate224inter0, gate224inter1, gate224inter2, gate224inter3, gate224inter4, gate224inter5, gate224inter6, gate224inter7, gate224inter8, gate224inter9, gate224inter10, gate224inter11, gate224inter12, gate240inter0, gate240inter1, gate240inter2, gate240inter3, gate240inter4, gate240inter5, gate240inter6, gate240inter7, gate240inter8, gate240inter9, gate240inter10, gate240inter11, gate240inter12, gate499inter0, gate499inter1, gate499inter2, gate499inter3, gate499inter4, gate499inter5, gate499inter6, gate499inter7, gate499inter8, gate499inter9, gate499inter10, gate499inter11, gate499inter12, gate214inter0, gate214inter1, gate214inter2, gate214inter3, gate214inter4, gate214inter5, gate214inter6, gate214inter7, gate214inter8, gate214inter9, gate214inter10, gate214inter11, gate214inter12, gate115inter0, gate115inter1, gate115inter2, gate115inter3, gate115inter4, gate115inter5, gate115inter6, gate115inter7, gate115inter8, gate115inter9, gate115inter10, gate115inter11, gate115inter12, gate116inter0, gate116inter1, gate116inter2, gate116inter3, gate116inter4, gate116inter5, gate116inter6, gate116inter7, gate116inter8, gate116inter9, gate116inter10, gate116inter11, gate116inter12, gate92inter0, gate92inter1, gate92inter2, gate92inter3, gate92inter4, gate92inter5, gate92inter6, gate92inter7, gate92inter8, gate92inter9, gate92inter10, gate92inter11, gate92inter12, gate235inter0, gate235inter1, gate235inter2, gate235inter3, gate235inter4, gate235inter5, gate235inter6, gate235inter7, gate235inter8, gate235inter9, gate235inter10, gate235inter11, gate235inter12, gate29inter0, gate29inter1, gate29inter2, gate29inter3, gate29inter4, gate29inter5, gate29inter6, gate29inter7, gate29inter8, gate29inter9, gate29inter10, gate29inter11, gate29inter12, gate154inter0, gate154inter1, gate154inter2, gate154inter3, gate154inter4, gate154inter5, gate154inter6, gate154inter7, gate154inter8, gate154inter9, gate154inter10, gate154inter11, gate154inter12, gate422inter0, gate422inter1, gate422inter2, gate422inter3, gate422inter4, gate422inter5, gate422inter6, gate422inter7, gate422inter8, gate422inter9, gate422inter10, gate422inter11, gate422inter12, gate399inter0, gate399inter1, gate399inter2, gate399inter3, gate399inter4, gate399inter5, gate399inter6, gate399inter7, gate399inter8, gate399inter9, gate399inter10, gate399inter11, gate399inter12, gate51inter0, gate51inter1, gate51inter2, gate51inter3, gate51inter4, gate51inter5, gate51inter6, gate51inter7, gate51inter8, gate51inter9, gate51inter10, gate51inter11, gate51inter12, gate440inter0, gate440inter1, gate440inter2, gate440inter3, gate440inter4, gate440inter5, gate440inter6, gate440inter7, gate440inter8, gate440inter9, gate440inter10, gate440inter11, gate440inter12, gate221inter0, gate221inter1, gate221inter2, gate221inter3, gate221inter4, gate221inter5, gate221inter6, gate221inter7, gate221inter8, gate221inter9, gate221inter10, gate221inter11, gate221inter12, gate123inter0, gate123inter1, gate123inter2, gate123inter3, gate123inter4, gate123inter5, gate123inter6, gate123inter7, gate123inter8, gate123inter9, gate123inter10, gate123inter11, gate123inter12, gate114inter0, gate114inter1, gate114inter2, gate114inter3, gate114inter4, gate114inter5, gate114inter6, gate114inter7, gate114inter8, gate114inter9, gate114inter10, gate114inter11, gate114inter12, gate460inter0, gate460inter1, gate460inter2, gate460inter3, gate460inter4, gate460inter5, gate460inter6, gate460inter7, gate460inter8, gate460inter9, gate460inter10, gate460inter11, gate460inter12, gate436inter0, gate436inter1, gate436inter2, gate436inter3, gate436inter4, gate436inter5, gate436inter6, gate436inter7, gate436inter8, gate436inter9, gate436inter10, gate436inter11, gate436inter12, gate204inter0, gate204inter1, gate204inter2, gate204inter3, gate204inter4, gate204inter5, gate204inter6, gate204inter7, gate204inter8, gate204inter9, gate204inter10, gate204inter11, gate204inter12, gate121inter0, gate121inter1, gate121inter2, gate121inter3, gate121inter4, gate121inter5, gate121inter6, gate121inter7, gate121inter8, gate121inter9, gate121inter10, gate121inter11, gate121inter12, gate478inter0, gate478inter1, gate478inter2, gate478inter3, gate478inter4, gate478inter5, gate478inter6, gate478inter7, gate478inter8, gate478inter9, gate478inter10, gate478inter11, gate478inter12, gate505inter0, gate505inter1, gate505inter2, gate505inter3, gate505inter4, gate505inter5, gate505inter6, gate505inter7, gate505inter8, gate505inter9, gate505inter10, gate505inter11, gate505inter12, gate220inter0, gate220inter1, gate220inter2, gate220inter3, gate220inter4, gate220inter5, gate220inter6, gate220inter7, gate220inter8, gate220inter9, gate220inter10, gate220inter11, gate220inter12, gate20inter0, gate20inter1, gate20inter2, gate20inter3, gate20inter4, gate20inter5, gate20inter6, gate20inter7, gate20inter8, gate20inter9, gate20inter10, gate20inter11, gate20inter12, gate459inter0, gate459inter1, gate459inter2, gate459inter3, gate459inter4, gate459inter5, gate459inter6, gate459inter7, gate459inter8, gate459inter9, gate459inter10, gate459inter11, gate459inter12, gate471inter0, gate471inter1, gate471inter2, gate471inter3, gate471inter4, gate471inter5, gate471inter6, gate471inter7, gate471inter8, gate471inter9, gate471inter10, gate471inter11, gate471inter12, gate278inter0, gate278inter1, gate278inter2, gate278inter3, gate278inter4, gate278inter5, gate278inter6, gate278inter7, gate278inter8, gate278inter9, gate278inter10, gate278inter11, gate278inter12, gate182inter0, gate182inter1, gate182inter2, gate182inter3, gate182inter4, gate182inter5, gate182inter6, gate182inter7, gate182inter8, gate182inter9, gate182inter10, gate182inter11, gate182inter12, gate11inter0, gate11inter1, gate11inter2, gate11inter3, gate11inter4, gate11inter5, gate11inter6, gate11inter7, gate11inter8, gate11inter9, gate11inter10, gate11inter11, gate11inter12, gate151inter0, gate151inter1, gate151inter2, gate151inter3, gate151inter4, gate151inter5, gate151inter6, gate151inter7, gate151inter8, gate151inter9, gate151inter10, gate151inter11, gate151inter12, gate251inter0, gate251inter1, gate251inter2, gate251inter3, gate251inter4, gate251inter5, gate251inter6, gate251inter7, gate251inter8, gate251inter9, gate251inter10, gate251inter11, gate251inter12, gate72inter0, gate72inter1, gate72inter2, gate72inter3, gate72inter4, gate72inter5, gate72inter6, gate72inter7, gate72inter8, gate72inter9, gate72inter10, gate72inter11, gate72inter12, gate12inter0, gate12inter1, gate12inter2, gate12inter3, gate12inter4, gate12inter5, gate12inter6, gate12inter7, gate12inter8, gate12inter9, gate12inter10, gate12inter11, gate12inter12, gate159inter0, gate159inter1, gate159inter2, gate159inter3, gate159inter4, gate159inter5, gate159inter6, gate159inter7, gate159inter8, gate159inter9, gate159inter10, gate159inter11, gate159inter12, gate285inter0, gate285inter1, gate285inter2, gate285inter3, gate285inter4, gate285inter5, gate285inter6, gate285inter7, gate285inter8, gate285inter9, gate285inter10, gate285inter11, gate285inter12, gate173inter0, gate173inter1, gate173inter2, gate173inter3, gate173inter4, gate173inter5, gate173inter6, gate173inter7, gate173inter8, gate173inter9, gate173inter10, gate173inter11, gate173inter12, gate136inter0, gate136inter1, gate136inter2, gate136inter3, gate136inter4, gate136inter5, gate136inter6, gate136inter7, gate136inter8, gate136inter9, gate136inter10, gate136inter11, gate136inter12, gate71inter0, gate71inter1, gate71inter2, gate71inter3, gate71inter4, gate71inter5, gate71inter6, gate71inter7, gate71inter8, gate71inter9, gate71inter10, gate71inter11, gate71inter12, gate419inter0, gate419inter1, gate419inter2, gate419inter3, gate419inter4, gate419inter5, gate419inter6, gate419inter7, gate419inter8, gate419inter9, gate419inter10, gate419inter11, gate419inter12, gate205inter0, gate205inter1, gate205inter2, gate205inter3, gate205inter4, gate205inter5, gate205inter6, gate205inter7, gate205inter8, gate205inter9, gate205inter10, gate205inter11, gate205inter12, gate463inter0, gate463inter1, gate463inter2, gate463inter3, gate463inter4, gate463inter5, gate463inter6, gate463inter7, gate463inter8, gate463inter9, gate463inter10, gate463inter11, gate463inter12, gate264inter0, gate264inter1, gate264inter2, gate264inter3, gate264inter4, gate264inter5, gate264inter6, gate264inter7, gate264inter8, gate264inter9, gate264inter10, gate264inter11, gate264inter12, gate420inter0, gate420inter1, gate420inter2, gate420inter3, gate420inter4, gate420inter5, gate420inter6, gate420inter7, gate420inter8, gate420inter9, gate420inter10, gate420inter11, gate420inter12, gate112inter0, gate112inter1, gate112inter2, gate112inter3, gate112inter4, gate112inter5, gate112inter6, gate112inter7, gate112inter8, gate112inter9, gate112inter10, gate112inter11, gate112inter12, gate80inter0, gate80inter1, gate80inter2, gate80inter3, gate80inter4, gate80inter5, gate80inter6, gate80inter7, gate80inter8, gate80inter9, gate80inter10, gate80inter11, gate80inter12, gate468inter0, gate468inter1, gate468inter2, gate468inter3, gate468inter4, gate468inter5, gate468inter6, gate468inter7, gate468inter8, gate468inter9, gate468inter10, gate468inter11, gate468inter12, gate26inter0, gate26inter1, gate26inter2, gate26inter3, gate26inter4, gate26inter5, gate26inter6, gate26inter7, gate26inter8, gate26inter9, gate26inter10, gate26inter11, gate26inter12, gate171inter0, gate171inter1, gate171inter2, gate171inter3, gate171inter4, gate171inter5, gate171inter6, gate171inter7, gate171inter8, gate171inter9, gate171inter10, gate171inter11, gate171inter12, gate431inter0, gate431inter1, gate431inter2, gate431inter3, gate431inter4, gate431inter5, gate431inter6, gate431inter7, gate431inter8, gate431inter9, gate431inter10, gate431inter11, gate431inter12, gate233inter0, gate233inter1, gate233inter2, gate233inter3, gate233inter4, gate233inter5, gate233inter6, gate233inter7, gate233inter8, gate233inter9, gate233inter10, gate233inter11, gate233inter12, gate194inter0, gate194inter1, gate194inter2, gate194inter3, gate194inter4, gate194inter5, gate194inter6, gate194inter7, gate194inter8, gate194inter9, gate194inter10, gate194inter11, gate194inter12, gate87inter0, gate87inter1, gate87inter2, gate87inter3, gate87inter4, gate87inter5, gate87inter6, gate87inter7, gate87inter8, gate87inter9, gate87inter10, gate87inter11, gate87inter12, gate492inter0, gate492inter1, gate492inter2, gate492inter3, gate492inter4, gate492inter5, gate492inter6, gate492inter7, gate492inter8, gate492inter9, gate492inter10, gate492inter11, gate492inter12, gate290inter0, gate290inter1, gate290inter2, gate290inter3, gate290inter4, gate290inter5, gate290inter6, gate290inter7, gate290inter8, gate290inter9, gate290inter10, gate290inter11, gate290inter12, gate56inter0, gate56inter1, gate56inter2, gate56inter3, gate56inter4, gate56inter5, gate56inter6, gate56inter7, gate56inter8, gate56inter9, gate56inter10, gate56inter11, gate56inter12, gate50inter0, gate50inter1, gate50inter2, gate50inter3, gate50inter4, gate50inter5, gate50inter6, gate50inter7, gate50inter8, gate50inter9, gate50inter10, gate50inter11, gate50inter12, gate433inter0, gate433inter1, gate433inter2, gate433inter3, gate433inter4, gate433inter5, gate433inter6, gate433inter7, gate433inter8, gate433inter9, gate433inter10, gate433inter11, gate433inter12, gate81inter0, gate81inter1, gate81inter2, gate81inter3, gate81inter4, gate81inter5, gate81inter6, gate81inter7, gate81inter8, gate81inter9, gate81inter10, gate81inter11, gate81inter12, gate504inter0, gate504inter1, gate504inter2, gate504inter3, gate504inter4, gate504inter5, gate504inter6, gate504inter7, gate504inter8, gate504inter9, gate504inter10, gate504inter11, gate504inter12, gate23inter0, gate23inter1, gate23inter2, gate23inter3, gate23inter4, gate23inter5, gate23inter6, gate23inter7, gate23inter8, gate23inter9, gate23inter10, gate23inter11, gate23inter12, gate418inter0, gate418inter1, gate418inter2, gate418inter3, gate418inter4, gate418inter5, gate418inter6, gate418inter7, gate418inter8, gate418inter9, gate418inter10, gate418inter11, gate418inter12, gate429inter0, gate429inter1, gate429inter2, gate429inter3, gate429inter4, gate429inter5, gate429inter6, gate429inter7, gate429inter8, gate429inter9, gate429inter10, gate429inter11, gate429inter12, gate60inter0, gate60inter1, gate60inter2, gate60inter3, gate60inter4, gate60inter5, gate60inter6, gate60inter7, gate60inter8, gate60inter9, gate60inter10, gate60inter11, gate60inter12, gate28inter0, gate28inter1, gate28inter2, gate28inter3, gate28inter4, gate28inter5, gate28inter6, gate28inter7, gate28inter8, gate28inter9, gate28inter10, gate28inter11, gate28inter12, gate101inter0, gate101inter1, gate101inter2, gate101inter3, gate101inter4, gate101inter5, gate101inter6, gate101inter7, gate101inter8, gate101inter9, gate101inter10, gate101inter11, gate101inter12, gate428inter0, gate428inter1, gate428inter2, gate428inter3, gate428inter4, gate428inter5, gate428inter6, gate428inter7, gate428inter8, gate428inter9, gate428inter10, gate428inter11, gate428inter12, gate445inter0, gate445inter1, gate445inter2, gate445inter3, gate445inter4, gate445inter5, gate445inter6, gate445inter7, gate445inter8, gate445inter9, gate445inter10, gate445inter11, gate445inter12, gate138inter0, gate138inter1, gate138inter2, gate138inter3, gate138inter4, gate138inter5, gate138inter6, gate138inter7, gate138inter8, gate138inter9, gate138inter10, gate138inter11, gate138inter12, gate100inter0, gate100inter1, gate100inter2, gate100inter3, gate100inter4, gate100inter5, gate100inter6, gate100inter7, gate100inter8, gate100inter9, gate100inter10, gate100inter11, gate100inter12, gate67inter0, gate67inter1, gate67inter2, gate67inter3, gate67inter4, gate67inter5, gate67inter6, gate67inter7, gate67inter8, gate67inter9, gate67inter10, gate67inter11, gate67inter12, gate55inter0, gate55inter1, gate55inter2, gate55inter3, gate55inter4, gate55inter5, gate55inter6, gate55inter7, gate55inter8, gate55inter9, gate55inter10, gate55inter11, gate55inter12, gate256inter0, gate256inter1, gate256inter2, gate256inter3, gate256inter4, gate256inter5, gate256inter6, gate256inter7, gate256inter8, gate256inter9, gate256inter10, gate256inter11, gate256inter12, gate249inter0, gate249inter1, gate249inter2, gate249inter3, gate249inter4, gate249inter5, gate249inter6, gate249inter7, gate249inter8, gate249inter9, gate249inter10, gate249inter11, gate249inter12, gate281inter0, gate281inter1, gate281inter2, gate281inter3, gate281inter4, gate281inter5, gate281inter6, gate281inter7, gate281inter8, gate281inter9, gate281inter10, gate281inter11, gate281inter12, gate132inter0, gate132inter1, gate132inter2, gate132inter3, gate132inter4, gate132inter5, gate132inter6, gate132inter7, gate132inter8, gate132inter9, gate132inter10, gate132inter11, gate132inter12, gate120inter0, gate120inter1, gate120inter2, gate120inter3, gate120inter4, gate120inter5, gate120inter6, gate120inter7, gate120inter8, gate120inter9, gate120inter10, gate120inter11, gate120inter12, gate437inter0, gate437inter1, gate437inter2, gate437inter3, gate437inter4, gate437inter5, gate437inter6, gate437inter7, gate437inter8, gate437inter9, gate437inter10, gate437inter11, gate437inter12, gate512inter0, gate512inter1, gate512inter2, gate512inter3, gate512inter4, gate512inter5, gate512inter6, gate512inter7, gate512inter8, gate512inter9, gate512inter10, gate512inter11, gate512inter12, gate203inter0, gate203inter1, gate203inter2, gate203inter3, gate203inter4, gate203inter5, gate203inter6, gate203inter7, gate203inter8, gate203inter9, gate203inter10, gate203inter11, gate203inter12, gate126inter0, gate126inter1, gate126inter2, gate126inter3, gate126inter4, gate126inter5, gate126inter6, gate126inter7, gate126inter8, gate126inter9, gate126inter10, gate126inter11, gate126inter12, gate191inter0, gate191inter1, gate191inter2, gate191inter3, gate191inter4, gate191inter5, gate191inter6, gate191inter7, gate191inter8, gate191inter9, gate191inter10, gate191inter11, gate191inter12, gate475inter0, gate475inter1, gate475inter2, gate475inter3, gate475inter4, gate475inter5, gate475inter6, gate475inter7, gate475inter8, gate475inter9, gate475inter10, gate475inter11, gate475inter12, gate283inter0, gate283inter1, gate283inter2, gate283inter3, gate283inter4, gate283inter5, gate283inter6, gate283inter7, gate283inter8, gate283inter9, gate283inter10, gate283inter11, gate283inter12, gate213inter0, gate213inter1, gate213inter2, gate213inter3, gate213inter4, gate213inter5, gate213inter6, gate213inter7, gate213inter8, gate213inter9, gate213inter10, gate213inter11, gate213inter12, gate498inter0, gate498inter1, gate498inter2, gate498inter3, gate498inter4, gate498inter5, gate498inter6, gate498inter7, gate498inter8, gate498inter9, gate498inter10, gate498inter11, gate498inter12, gate275inter0, gate275inter1, gate275inter2, gate275inter3, gate275inter4, gate275inter5, gate275inter6, gate275inter7, gate275inter8, gate275inter9, gate275inter10, gate275inter11, gate275inter12, gate74inter0, gate74inter1, gate74inter2, gate74inter3, gate74inter4, gate74inter5, gate74inter6, gate74inter7, gate74inter8, gate74inter9, gate74inter10, gate74inter11, gate74inter12, gate75inter0, gate75inter1, gate75inter2, gate75inter3, gate75inter4, gate75inter5, gate75inter6, gate75inter7, gate75inter8, gate75inter9, gate75inter10, gate75inter11, gate75inter12, gate450inter0, gate450inter1, gate450inter2, gate450inter3, gate450inter4, gate450inter5, gate450inter6, gate450inter7, gate450inter8, gate450inter9, gate450inter10, gate450inter11, gate450inter12, gate161inter0, gate161inter1, gate161inter2, gate161inter3, gate161inter4, gate161inter5, gate161inter6, gate161inter7, gate161inter8, gate161inter9, gate161inter10, gate161inter11, gate161inter12, gate36inter0, gate36inter1, gate36inter2, gate36inter3, gate36inter4, gate36inter5, gate36inter6, gate36inter7, gate36inter8, gate36inter9, gate36inter10, gate36inter11, gate36inter12, gate461inter0, gate461inter1, gate461inter2, gate461inter3, gate461inter4, gate461inter5, gate461inter6, gate461inter7, gate461inter8, gate461inter9, gate461inter10, gate461inter11, gate461inter12, gate389inter0, gate389inter1, gate389inter2, gate389inter3, gate389inter4, gate389inter5, gate389inter6, gate389inter7, gate389inter8, gate389inter9, gate389inter10, gate389inter11, gate389inter12, gate412inter0, gate412inter1, gate412inter2, gate412inter3, gate412inter4, gate412inter5, gate412inter6, gate412inter7, gate412inter8, gate412inter9, gate412inter10, gate412inter11, gate412inter12, gate239inter0, gate239inter1, gate239inter2, gate239inter3, gate239inter4, gate239inter5, gate239inter6, gate239inter7, gate239inter8, gate239inter9, gate239inter10, gate239inter11, gate239inter12, gate417inter0, gate417inter1, gate417inter2, gate417inter3, gate417inter4, gate417inter5, gate417inter6, gate417inter7, gate417inter8, gate417inter9, gate417inter10, gate417inter11, gate417inter12, gate502inter0, gate502inter1, gate502inter2, gate502inter3, gate502inter4, gate502inter5, gate502inter6, gate502inter7, gate502inter8, gate502inter9, gate502inter10, gate502inter11, gate502inter12, gate22inter0, gate22inter1, gate22inter2, gate22inter3, gate22inter4, gate22inter5, gate22inter6, gate22inter7, gate22inter8, gate22inter9, gate22inter10, gate22inter11, gate22inter12, gate207inter0, gate207inter1, gate207inter2, gate207inter3, gate207inter4, gate207inter5, gate207inter6, gate207inter7, gate207inter8, gate207inter9, gate207inter10, gate207inter11, gate207inter12, gate446inter0, gate446inter1, gate446inter2, gate446inter3, gate446inter4, gate446inter5, gate446inter6, gate446inter7, gate446inter8, gate446inter9, gate446inter10, gate446inter11, gate446inter12, gate476inter0, gate476inter1, gate476inter2, gate476inter3, gate476inter4, gate476inter5, gate476inter6, gate476inter7, gate476inter8, gate476inter9, gate476inter10, gate476inter11, gate476inter12, gate96inter0, gate96inter1, gate96inter2, gate96inter3, gate96inter4, gate96inter5, gate96inter6, gate96inter7, gate96inter8, gate96inter9, gate96inter10, gate96inter11, gate96inter12, gate258inter0, gate258inter1, gate258inter2, gate258inter3, gate258inter4, gate258inter5, gate258inter6, gate258inter7, gate258inter8, gate258inter9, gate258inter10, gate258inter11, gate258inter12, gate396inter0, gate396inter1, gate396inter2, gate396inter3, gate396inter4, gate396inter5, gate396inter6, gate396inter7, gate396inter8, gate396inter9, gate396inter10, gate396inter11, gate396inter12, gate106inter0, gate106inter1, gate106inter2, gate106inter3, gate106inter4, gate106inter5, gate106inter6, gate106inter7, gate106inter8, gate106inter9, gate106inter10, gate106inter11, gate106inter12, gate21inter0, gate21inter1, gate21inter2, gate21inter3, gate21inter4, gate21inter5, gate21inter6, gate21inter7, gate21inter8, gate21inter9, gate21inter10, gate21inter11, gate21inter12, gate265inter0, gate265inter1, gate265inter2, gate265inter3, gate265inter4, gate265inter5, gate265inter6, gate265inter7, gate265inter8, gate265inter9, gate265inter10, gate265inter11, gate265inter12, gate484inter0, gate484inter1, gate484inter2, gate484inter3, gate484inter4, gate484inter5, gate484inter6, gate484inter7, gate484inter8, gate484inter9, gate484inter10, gate484inter11, gate484inter12, gate17inter0, gate17inter1, gate17inter2, gate17inter3, gate17inter4, gate17inter5, gate17inter6, gate17inter7, gate17inter8, gate17inter9, gate17inter10, gate17inter11, gate17inter12, gate236inter0, gate236inter1, gate236inter2, gate236inter3, gate236inter4, gate236inter5, gate236inter6, gate236inter7, gate236inter8, gate236inter9, gate236inter10, gate236inter11, gate236inter12, gate467inter0, gate467inter1, gate467inter2, gate467inter3, gate467inter4, gate467inter5, gate467inter6, gate467inter7, gate467inter8, gate467inter9, gate467inter10, gate467inter11, gate467inter12, gate118inter0, gate118inter1, gate118inter2, gate118inter3, gate118inter4, gate118inter5, gate118inter6, gate118inter7, gate118inter8, gate118inter9, gate118inter10, gate118inter11, gate118inter12, gate145inter0, gate145inter1, gate145inter2, gate145inter3, gate145inter4, gate145inter5, gate145inter6, gate145inter7, gate145inter8, gate145inter9, gate145inter10, gate145inter11, gate145inter12, gate455inter0, gate455inter1, gate455inter2, gate455inter3, gate455inter4, gate455inter5, gate455inter6, gate455inter7, gate455inter8, gate455inter9, gate455inter10, gate455inter11, gate455inter12, gate494inter0, gate494inter1, gate494inter2, gate494inter3, gate494inter4, gate494inter5, gate494inter6, gate494inter7, gate494inter8, gate494inter9, gate494inter10, gate494inter11, gate494inter12, gate166inter0, gate166inter1, gate166inter2, gate166inter3, gate166inter4, gate166inter5, gate166inter6, gate166inter7, gate166inter8, gate166inter9, gate166inter10, gate166inter11, gate166inter12, gate510inter0, gate510inter1, gate510inter2, gate510inter3, gate510inter4, gate510inter5, gate510inter6, gate510inter7, gate510inter8, gate510inter9, gate510inter10, gate510inter11, gate510inter12, gate245inter0, gate245inter1, gate245inter2, gate245inter3, gate245inter4, gate245inter5, gate245inter6, gate245inter7, gate245inter8, gate245inter9, gate245inter10, gate245inter11, gate245inter12, gate454inter0, gate454inter1, gate454inter2, gate454inter3, gate454inter4, gate454inter5, gate454inter6, gate454inter7, gate454inter8, gate454inter9, gate454inter10, gate454inter11, gate454inter12, gate135inter0, gate135inter1, gate135inter2, gate135inter3, gate135inter4, gate135inter5, gate135inter6, gate135inter7, gate135inter8, gate135inter9, gate135inter10, gate135inter11, gate135inter12, gate223inter0, gate223inter1, gate223inter2, gate223inter3, gate223inter4, gate223inter5, gate223inter6, gate223inter7, gate223inter8, gate223inter9, gate223inter10, gate223inter11, gate223inter12, gate444inter0, gate444inter1, gate444inter2, gate444inter3, gate444inter4, gate444inter5, gate444inter6, gate444inter7, gate444inter8, gate444inter9, gate444inter10, gate444inter11, gate444inter12, gate44inter0, gate44inter1, gate44inter2, gate44inter3, gate44inter4, gate44inter5, gate44inter6, gate44inter7, gate44inter8, gate44inter9, gate44inter10, gate44inter11, gate44inter12, gate65inter0, gate65inter1, gate65inter2, gate65inter3, gate65inter4, gate65inter5, gate65inter6, gate65inter7, gate65inter8, gate65inter9, gate65inter10, gate65inter11, gate65inter12, gate416inter0, gate416inter1, gate416inter2, gate416inter3, gate416inter4, gate416inter5, gate416inter6, gate416inter7, gate416inter8, gate416inter9, gate416inter10, gate416inter11, gate416inter12, gate211inter0, gate211inter1, gate211inter2, gate211inter3, gate211inter4, gate211inter5, gate211inter6, gate211inter7, gate211inter8, gate211inter9, gate211inter10, gate211inter11, gate211inter12, gate134inter0, gate134inter1, gate134inter2, gate134inter3, gate134inter4, gate134inter5, gate134inter6, gate134inter7, gate134inter8, gate134inter9, gate134inter10, gate134inter11, gate134inter12, gate156inter0, gate156inter1, gate156inter2, gate156inter3, gate156inter4, gate156inter5, gate156inter6, gate156inter7, gate156inter8, gate156inter9, gate156inter10, gate156inter11, gate156inter12, gate509inter0, gate509inter1, gate509inter2, gate509inter3, gate509inter4, gate509inter5, gate509inter6, gate509inter7, gate509inter8, gate509inter9, gate509inter10, gate509inter11, gate509inter12, gate148inter0, gate148inter1, gate148inter2, gate148inter3, gate148inter4, gate148inter5, gate148inter6, gate148inter7, gate148inter8, gate148inter9, gate148inter10, gate148inter11, gate148inter12, gate404inter0, gate404inter1, gate404inter2, gate404inter3, gate404inter4, gate404inter5, gate404inter6, gate404inter7, gate404inter8, gate404inter9, gate404inter10, gate404inter11, gate404inter12, gate286inter0, gate286inter1, gate286inter2, gate286inter3, gate286inter4, gate286inter5, gate286inter6, gate286inter7, gate286inter8, gate286inter9, gate286inter10, gate286inter11, gate286inter12, gate212inter0, gate212inter1, gate212inter2, gate212inter3, gate212inter4, gate212inter5, gate212inter6, gate212inter7, gate212inter8, gate212inter9, gate212inter10, gate212inter11, gate212inter12, gate453inter0, gate453inter1, gate453inter2, gate453inter3, gate453inter4, gate453inter5, gate453inter6, gate453inter7, gate453inter8, gate453inter9, gate453inter10, gate453inter11, gate453inter12, gate289inter0, gate289inter1, gate289inter2, gate289inter3, gate289inter4, gate289inter5, gate289inter6, gate289inter7, gate289inter8, gate289inter9, gate289inter10, gate289inter11, gate289inter12, gate496inter0, gate496inter1, gate496inter2, gate496inter3, gate496inter4, gate496inter5, gate496inter6, gate496inter7, gate496inter8, gate496inter9, gate496inter10, gate496inter11, gate496inter12, gate77inter0, gate77inter1, gate77inter2, gate77inter3, gate77inter4, gate77inter5, gate77inter6, gate77inter7, gate77inter8, gate77inter9, gate77inter10, gate77inter11, gate77inter12, gate409inter0, gate409inter1, gate409inter2, gate409inter3, gate409inter4, gate409inter5, gate409inter6, gate409inter7, gate409inter8, gate409inter9, gate409inter10, gate409inter11, gate409inter12;



and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );
nand2 gate9( .a(G1), .b(G2), .O(G266) );
nand2 gate10( .a(G3), .b(G4), .O(G269) );

  xor2  gate1471(.a(G6), .b(G5), .O(gate11inter0));
  nand2 gate1472(.a(gate11inter0), .b(s_132), .O(gate11inter1));
  and2  gate1473(.a(G6), .b(G5), .O(gate11inter2));
  inv1  gate1474(.a(s_132), .O(gate11inter3));
  inv1  gate1475(.a(s_133), .O(gate11inter4));
  nand2 gate1476(.a(gate11inter4), .b(gate11inter3), .O(gate11inter5));
  nor2  gate1477(.a(gate11inter5), .b(gate11inter2), .O(gate11inter6));
  inv1  gate1478(.a(G5), .O(gate11inter7));
  inv1  gate1479(.a(G6), .O(gate11inter8));
  nand2 gate1480(.a(gate11inter8), .b(gate11inter7), .O(gate11inter9));
  nand2 gate1481(.a(s_133), .b(gate11inter3), .O(gate11inter10));
  nor2  gate1482(.a(gate11inter10), .b(gate11inter9), .O(gate11inter11));
  nor2  gate1483(.a(gate11inter11), .b(gate11inter6), .O(gate11inter12));
  nand2 gate1484(.a(gate11inter12), .b(gate11inter1), .O(G272));

  xor2  gate1527(.a(G8), .b(G7), .O(gate12inter0));
  nand2 gate1528(.a(gate12inter0), .b(s_140), .O(gate12inter1));
  and2  gate1529(.a(G8), .b(G7), .O(gate12inter2));
  inv1  gate1530(.a(s_140), .O(gate12inter3));
  inv1  gate1531(.a(s_141), .O(gate12inter4));
  nand2 gate1532(.a(gate12inter4), .b(gate12inter3), .O(gate12inter5));
  nor2  gate1533(.a(gate12inter5), .b(gate12inter2), .O(gate12inter6));
  inv1  gate1534(.a(G7), .O(gate12inter7));
  inv1  gate1535(.a(G8), .O(gate12inter8));
  nand2 gate1536(.a(gate12inter8), .b(gate12inter7), .O(gate12inter9));
  nand2 gate1537(.a(s_141), .b(gate12inter3), .O(gate12inter10));
  nor2  gate1538(.a(gate12inter10), .b(gate12inter9), .O(gate12inter11));
  nor2  gate1539(.a(gate12inter11), .b(gate12inter6), .O(gate12inter12));
  nand2 gate1540(.a(gate12inter12), .b(gate12inter1), .O(G275));
nand2 gate13( .a(G9), .b(G10), .O(G278) );
nand2 gate14( .a(G11), .b(G12), .O(G281) );
nand2 gate15( .a(G13), .b(G14), .O(G284) );

  xor2  gate897(.a(G16), .b(G15), .O(gate16inter0));
  nand2 gate898(.a(gate16inter0), .b(s_50), .O(gate16inter1));
  and2  gate899(.a(G16), .b(G15), .O(gate16inter2));
  inv1  gate900(.a(s_50), .O(gate16inter3));
  inv1  gate901(.a(s_51), .O(gate16inter4));
  nand2 gate902(.a(gate16inter4), .b(gate16inter3), .O(gate16inter5));
  nor2  gate903(.a(gate16inter5), .b(gate16inter2), .O(gate16inter6));
  inv1  gate904(.a(G15), .O(gate16inter7));
  inv1  gate905(.a(G16), .O(gate16inter8));
  nand2 gate906(.a(gate16inter8), .b(gate16inter7), .O(gate16inter9));
  nand2 gate907(.a(s_51), .b(gate16inter3), .O(gate16inter10));
  nor2  gate908(.a(gate16inter10), .b(gate16inter9), .O(gate16inter11));
  nor2  gate909(.a(gate16inter11), .b(gate16inter6), .O(gate16inter12));
  nand2 gate910(.a(gate16inter12), .b(gate16inter1), .O(G287));

  xor2  gate2591(.a(G18), .b(G17), .O(gate17inter0));
  nand2 gate2592(.a(gate17inter0), .b(s_292), .O(gate17inter1));
  and2  gate2593(.a(G18), .b(G17), .O(gate17inter2));
  inv1  gate2594(.a(s_292), .O(gate17inter3));
  inv1  gate2595(.a(s_293), .O(gate17inter4));
  nand2 gate2596(.a(gate17inter4), .b(gate17inter3), .O(gate17inter5));
  nor2  gate2597(.a(gate17inter5), .b(gate17inter2), .O(gate17inter6));
  inv1  gate2598(.a(G17), .O(gate17inter7));
  inv1  gate2599(.a(G18), .O(gate17inter8));
  nand2 gate2600(.a(gate17inter8), .b(gate17inter7), .O(gate17inter9));
  nand2 gate2601(.a(s_293), .b(gate17inter3), .O(gate17inter10));
  nor2  gate2602(.a(gate17inter10), .b(gate17inter9), .O(gate17inter11));
  nor2  gate2603(.a(gate17inter11), .b(gate17inter6), .O(gate17inter12));
  nand2 gate2604(.a(gate17inter12), .b(gate17inter1), .O(G290));
nand2 gate18( .a(G19), .b(G20), .O(G293) );
nand2 gate19( .a(G21), .b(G22), .O(G296) );

  xor2  gate1401(.a(G24), .b(G23), .O(gate20inter0));
  nand2 gate1402(.a(gate20inter0), .b(s_122), .O(gate20inter1));
  and2  gate1403(.a(G24), .b(G23), .O(gate20inter2));
  inv1  gate1404(.a(s_122), .O(gate20inter3));
  inv1  gate1405(.a(s_123), .O(gate20inter4));
  nand2 gate1406(.a(gate20inter4), .b(gate20inter3), .O(gate20inter5));
  nor2  gate1407(.a(gate20inter5), .b(gate20inter2), .O(gate20inter6));
  inv1  gate1408(.a(G23), .O(gate20inter7));
  inv1  gate1409(.a(G24), .O(gate20inter8));
  nand2 gate1410(.a(gate20inter8), .b(gate20inter7), .O(gate20inter9));
  nand2 gate1411(.a(s_123), .b(gate20inter3), .O(gate20inter10));
  nor2  gate1412(.a(gate20inter10), .b(gate20inter9), .O(gate20inter11));
  nor2  gate1413(.a(gate20inter11), .b(gate20inter6), .O(gate20inter12));
  nand2 gate1414(.a(gate20inter12), .b(gate20inter1), .O(G299));

  xor2  gate2549(.a(G26), .b(G25), .O(gate21inter0));
  nand2 gate2550(.a(gate21inter0), .b(s_286), .O(gate21inter1));
  and2  gate2551(.a(G26), .b(G25), .O(gate21inter2));
  inv1  gate2552(.a(s_286), .O(gate21inter3));
  inv1  gate2553(.a(s_287), .O(gate21inter4));
  nand2 gate2554(.a(gate21inter4), .b(gate21inter3), .O(gate21inter5));
  nor2  gate2555(.a(gate21inter5), .b(gate21inter2), .O(gate21inter6));
  inv1  gate2556(.a(G25), .O(gate21inter7));
  inv1  gate2557(.a(G26), .O(gate21inter8));
  nand2 gate2558(.a(gate21inter8), .b(gate21inter7), .O(gate21inter9));
  nand2 gate2559(.a(s_287), .b(gate21inter3), .O(gate21inter10));
  nor2  gate2560(.a(gate21inter10), .b(gate21inter9), .O(gate21inter11));
  nor2  gate2561(.a(gate21inter11), .b(gate21inter6), .O(gate21inter12));
  nand2 gate2562(.a(gate21inter12), .b(gate21inter1), .O(G302));

  xor2  gate2437(.a(G28), .b(G27), .O(gate22inter0));
  nand2 gate2438(.a(gate22inter0), .b(s_270), .O(gate22inter1));
  and2  gate2439(.a(G28), .b(G27), .O(gate22inter2));
  inv1  gate2440(.a(s_270), .O(gate22inter3));
  inv1  gate2441(.a(s_271), .O(gate22inter4));
  nand2 gate2442(.a(gate22inter4), .b(gate22inter3), .O(gate22inter5));
  nor2  gate2443(.a(gate22inter5), .b(gate22inter2), .O(gate22inter6));
  inv1  gate2444(.a(G27), .O(gate22inter7));
  inv1  gate2445(.a(G28), .O(gate22inter8));
  nand2 gate2446(.a(gate22inter8), .b(gate22inter7), .O(gate22inter9));
  nand2 gate2447(.a(s_271), .b(gate22inter3), .O(gate22inter10));
  nor2  gate2448(.a(gate22inter10), .b(gate22inter9), .O(gate22inter11));
  nor2  gate2449(.a(gate22inter11), .b(gate22inter6), .O(gate22inter12));
  nand2 gate2450(.a(gate22inter12), .b(gate22inter1), .O(G305));

  xor2  gate1905(.a(G30), .b(G29), .O(gate23inter0));
  nand2 gate1906(.a(gate23inter0), .b(s_194), .O(gate23inter1));
  and2  gate1907(.a(G30), .b(G29), .O(gate23inter2));
  inv1  gate1908(.a(s_194), .O(gate23inter3));
  inv1  gate1909(.a(s_195), .O(gate23inter4));
  nand2 gate1910(.a(gate23inter4), .b(gate23inter3), .O(gate23inter5));
  nor2  gate1911(.a(gate23inter5), .b(gate23inter2), .O(gate23inter6));
  inv1  gate1912(.a(G29), .O(gate23inter7));
  inv1  gate1913(.a(G30), .O(gate23inter8));
  nand2 gate1914(.a(gate23inter8), .b(gate23inter7), .O(gate23inter9));
  nand2 gate1915(.a(s_195), .b(gate23inter3), .O(gate23inter10));
  nor2  gate1916(.a(gate23inter10), .b(gate23inter9), .O(gate23inter11));
  nor2  gate1917(.a(gate23inter11), .b(gate23inter6), .O(gate23inter12));
  nand2 gate1918(.a(gate23inter12), .b(gate23inter1), .O(G308));
nand2 gate24( .a(G31), .b(G32), .O(G311) );
nand2 gate25( .a(G1), .b(G5), .O(G314) );

  xor2  gate1723(.a(G13), .b(G9), .O(gate26inter0));
  nand2 gate1724(.a(gate26inter0), .b(s_168), .O(gate26inter1));
  and2  gate1725(.a(G13), .b(G9), .O(gate26inter2));
  inv1  gate1726(.a(s_168), .O(gate26inter3));
  inv1  gate1727(.a(s_169), .O(gate26inter4));
  nand2 gate1728(.a(gate26inter4), .b(gate26inter3), .O(gate26inter5));
  nor2  gate1729(.a(gate26inter5), .b(gate26inter2), .O(gate26inter6));
  inv1  gate1730(.a(G9), .O(gate26inter7));
  inv1  gate1731(.a(G13), .O(gate26inter8));
  nand2 gate1732(.a(gate26inter8), .b(gate26inter7), .O(gate26inter9));
  nand2 gate1733(.a(s_169), .b(gate26inter3), .O(gate26inter10));
  nor2  gate1734(.a(gate26inter10), .b(gate26inter9), .O(gate26inter11));
  nor2  gate1735(.a(gate26inter11), .b(gate26inter6), .O(gate26inter12));
  nand2 gate1736(.a(gate26inter12), .b(gate26inter1), .O(G317));
nand2 gate27( .a(G2), .b(G6), .O(G320) );

  xor2  gate1961(.a(G14), .b(G10), .O(gate28inter0));
  nand2 gate1962(.a(gate28inter0), .b(s_202), .O(gate28inter1));
  and2  gate1963(.a(G14), .b(G10), .O(gate28inter2));
  inv1  gate1964(.a(s_202), .O(gate28inter3));
  inv1  gate1965(.a(s_203), .O(gate28inter4));
  nand2 gate1966(.a(gate28inter4), .b(gate28inter3), .O(gate28inter5));
  nor2  gate1967(.a(gate28inter5), .b(gate28inter2), .O(gate28inter6));
  inv1  gate1968(.a(G10), .O(gate28inter7));
  inv1  gate1969(.a(G14), .O(gate28inter8));
  nand2 gate1970(.a(gate28inter8), .b(gate28inter7), .O(gate28inter9));
  nand2 gate1971(.a(s_203), .b(gate28inter3), .O(gate28inter10));
  nor2  gate1972(.a(gate28inter10), .b(gate28inter9), .O(gate28inter11));
  nor2  gate1973(.a(gate28inter11), .b(gate28inter6), .O(gate28inter12));
  nand2 gate1974(.a(gate28inter12), .b(gate28inter1), .O(G323));

  xor2  gate1177(.a(G7), .b(G3), .O(gate29inter0));
  nand2 gate1178(.a(gate29inter0), .b(s_90), .O(gate29inter1));
  and2  gate1179(.a(G7), .b(G3), .O(gate29inter2));
  inv1  gate1180(.a(s_90), .O(gate29inter3));
  inv1  gate1181(.a(s_91), .O(gate29inter4));
  nand2 gate1182(.a(gate29inter4), .b(gate29inter3), .O(gate29inter5));
  nor2  gate1183(.a(gate29inter5), .b(gate29inter2), .O(gate29inter6));
  inv1  gate1184(.a(G3), .O(gate29inter7));
  inv1  gate1185(.a(G7), .O(gate29inter8));
  nand2 gate1186(.a(gate29inter8), .b(gate29inter7), .O(gate29inter9));
  nand2 gate1187(.a(s_91), .b(gate29inter3), .O(gate29inter10));
  nor2  gate1188(.a(gate29inter10), .b(gate29inter9), .O(gate29inter11));
  nor2  gate1189(.a(gate29inter11), .b(gate29inter6), .O(gate29inter12));
  nand2 gate1190(.a(gate29inter12), .b(gate29inter1), .O(G326));
nand2 gate30( .a(G11), .b(G15), .O(G329) );
nand2 gate31( .a(G4), .b(G8), .O(G332) );

  xor2  gate1009(.a(G16), .b(G12), .O(gate32inter0));
  nand2 gate1010(.a(gate32inter0), .b(s_66), .O(gate32inter1));
  and2  gate1011(.a(G16), .b(G12), .O(gate32inter2));
  inv1  gate1012(.a(s_66), .O(gate32inter3));
  inv1  gate1013(.a(s_67), .O(gate32inter4));
  nand2 gate1014(.a(gate32inter4), .b(gate32inter3), .O(gate32inter5));
  nor2  gate1015(.a(gate32inter5), .b(gate32inter2), .O(gate32inter6));
  inv1  gate1016(.a(G12), .O(gate32inter7));
  inv1  gate1017(.a(G16), .O(gate32inter8));
  nand2 gate1018(.a(gate32inter8), .b(gate32inter7), .O(gate32inter9));
  nand2 gate1019(.a(s_67), .b(gate32inter3), .O(gate32inter10));
  nor2  gate1020(.a(gate32inter10), .b(gate32inter9), .O(gate32inter11));
  nor2  gate1021(.a(gate32inter11), .b(gate32inter6), .O(gate32inter12));
  nand2 gate1022(.a(gate32inter12), .b(gate32inter1), .O(G335));
nand2 gate33( .a(G17), .b(G21), .O(G338) );
nand2 gate34( .a(G25), .b(G29), .O(G341) );
nand2 gate35( .a(G18), .b(G22), .O(G344) );

  xor2  gate2339(.a(G30), .b(G26), .O(gate36inter0));
  nand2 gate2340(.a(gate36inter0), .b(s_256), .O(gate36inter1));
  and2  gate2341(.a(G30), .b(G26), .O(gate36inter2));
  inv1  gate2342(.a(s_256), .O(gate36inter3));
  inv1  gate2343(.a(s_257), .O(gate36inter4));
  nand2 gate2344(.a(gate36inter4), .b(gate36inter3), .O(gate36inter5));
  nor2  gate2345(.a(gate36inter5), .b(gate36inter2), .O(gate36inter6));
  inv1  gate2346(.a(G26), .O(gate36inter7));
  inv1  gate2347(.a(G30), .O(gate36inter8));
  nand2 gate2348(.a(gate36inter8), .b(gate36inter7), .O(gate36inter9));
  nand2 gate2349(.a(s_257), .b(gate36inter3), .O(gate36inter10));
  nor2  gate2350(.a(gate36inter10), .b(gate36inter9), .O(gate36inter11));
  nor2  gate2351(.a(gate36inter11), .b(gate36inter6), .O(gate36inter12));
  nand2 gate2352(.a(gate36inter12), .b(gate36inter1), .O(G347));
nand2 gate37( .a(G19), .b(G23), .O(G350) );
nand2 gate38( .a(G27), .b(G31), .O(G353) );
nand2 gate39( .a(G20), .b(G24), .O(G356) );
nand2 gate40( .a(G28), .b(G32), .O(G359) );
nand2 gate41( .a(G1), .b(G266), .O(G362) );
nand2 gate42( .a(G2), .b(G266), .O(G363) );
nand2 gate43( .a(G3), .b(G269), .O(G364) );

  xor2  gate2787(.a(G269), .b(G4), .O(gate44inter0));
  nand2 gate2788(.a(gate44inter0), .b(s_320), .O(gate44inter1));
  and2  gate2789(.a(G269), .b(G4), .O(gate44inter2));
  inv1  gate2790(.a(s_320), .O(gate44inter3));
  inv1  gate2791(.a(s_321), .O(gate44inter4));
  nand2 gate2792(.a(gate44inter4), .b(gate44inter3), .O(gate44inter5));
  nor2  gate2793(.a(gate44inter5), .b(gate44inter2), .O(gate44inter6));
  inv1  gate2794(.a(G4), .O(gate44inter7));
  inv1  gate2795(.a(G269), .O(gate44inter8));
  nand2 gate2796(.a(gate44inter8), .b(gate44inter7), .O(gate44inter9));
  nand2 gate2797(.a(s_321), .b(gate44inter3), .O(gate44inter10));
  nor2  gate2798(.a(gate44inter10), .b(gate44inter9), .O(gate44inter11));
  nor2  gate2799(.a(gate44inter11), .b(gate44inter6), .O(gate44inter12));
  nand2 gate2800(.a(gate44inter12), .b(gate44inter1), .O(G365));
nand2 gate45( .a(G5), .b(G272), .O(G366) );
nand2 gate46( .a(G6), .b(G272), .O(G367) );
nand2 gate47( .a(G7), .b(G275), .O(G368) );
nand2 gate48( .a(G8), .b(G275), .O(G369) );
nand2 gate49( .a(G9), .b(G278), .O(G370) );

  xor2  gate1849(.a(G278), .b(G10), .O(gate50inter0));
  nand2 gate1850(.a(gate50inter0), .b(s_186), .O(gate50inter1));
  and2  gate1851(.a(G278), .b(G10), .O(gate50inter2));
  inv1  gate1852(.a(s_186), .O(gate50inter3));
  inv1  gate1853(.a(s_187), .O(gate50inter4));
  nand2 gate1854(.a(gate50inter4), .b(gate50inter3), .O(gate50inter5));
  nor2  gate1855(.a(gate50inter5), .b(gate50inter2), .O(gate50inter6));
  inv1  gate1856(.a(G10), .O(gate50inter7));
  inv1  gate1857(.a(G278), .O(gate50inter8));
  nand2 gate1858(.a(gate50inter8), .b(gate50inter7), .O(gate50inter9));
  nand2 gate1859(.a(s_187), .b(gate50inter3), .O(gate50inter10));
  nor2  gate1860(.a(gate50inter10), .b(gate50inter9), .O(gate50inter11));
  nor2  gate1861(.a(gate50inter11), .b(gate50inter6), .O(gate50inter12));
  nand2 gate1862(.a(gate50inter12), .b(gate50inter1), .O(G371));

  xor2  gate1233(.a(G281), .b(G11), .O(gate51inter0));
  nand2 gate1234(.a(gate51inter0), .b(s_98), .O(gate51inter1));
  and2  gate1235(.a(G281), .b(G11), .O(gate51inter2));
  inv1  gate1236(.a(s_98), .O(gate51inter3));
  inv1  gate1237(.a(s_99), .O(gate51inter4));
  nand2 gate1238(.a(gate51inter4), .b(gate51inter3), .O(gate51inter5));
  nor2  gate1239(.a(gate51inter5), .b(gate51inter2), .O(gate51inter6));
  inv1  gate1240(.a(G11), .O(gate51inter7));
  inv1  gate1241(.a(G281), .O(gate51inter8));
  nand2 gate1242(.a(gate51inter8), .b(gate51inter7), .O(gate51inter9));
  nand2 gate1243(.a(s_99), .b(gate51inter3), .O(gate51inter10));
  nor2  gate1244(.a(gate51inter10), .b(gate51inter9), .O(gate51inter11));
  nor2  gate1245(.a(gate51inter11), .b(gate51inter6), .O(gate51inter12));
  nand2 gate1246(.a(gate51inter12), .b(gate51inter1), .O(G372));
nand2 gate52( .a(G12), .b(G281), .O(G373) );

  xor2  gate785(.a(G284), .b(G13), .O(gate53inter0));
  nand2 gate786(.a(gate53inter0), .b(s_34), .O(gate53inter1));
  and2  gate787(.a(G284), .b(G13), .O(gate53inter2));
  inv1  gate788(.a(s_34), .O(gate53inter3));
  inv1  gate789(.a(s_35), .O(gate53inter4));
  nand2 gate790(.a(gate53inter4), .b(gate53inter3), .O(gate53inter5));
  nor2  gate791(.a(gate53inter5), .b(gate53inter2), .O(gate53inter6));
  inv1  gate792(.a(G13), .O(gate53inter7));
  inv1  gate793(.a(G284), .O(gate53inter8));
  nand2 gate794(.a(gate53inter8), .b(gate53inter7), .O(gate53inter9));
  nand2 gate795(.a(s_35), .b(gate53inter3), .O(gate53inter10));
  nor2  gate796(.a(gate53inter10), .b(gate53inter9), .O(gate53inter11));
  nor2  gate797(.a(gate53inter11), .b(gate53inter6), .O(gate53inter12));
  nand2 gate798(.a(gate53inter12), .b(gate53inter1), .O(G374));
nand2 gate54( .a(G14), .b(G284), .O(G375) );

  xor2  gate2059(.a(G287), .b(G15), .O(gate55inter0));
  nand2 gate2060(.a(gate55inter0), .b(s_216), .O(gate55inter1));
  and2  gate2061(.a(G287), .b(G15), .O(gate55inter2));
  inv1  gate2062(.a(s_216), .O(gate55inter3));
  inv1  gate2063(.a(s_217), .O(gate55inter4));
  nand2 gate2064(.a(gate55inter4), .b(gate55inter3), .O(gate55inter5));
  nor2  gate2065(.a(gate55inter5), .b(gate55inter2), .O(gate55inter6));
  inv1  gate2066(.a(G15), .O(gate55inter7));
  inv1  gate2067(.a(G287), .O(gate55inter8));
  nand2 gate2068(.a(gate55inter8), .b(gate55inter7), .O(gate55inter9));
  nand2 gate2069(.a(s_217), .b(gate55inter3), .O(gate55inter10));
  nor2  gate2070(.a(gate55inter10), .b(gate55inter9), .O(gate55inter11));
  nor2  gate2071(.a(gate55inter11), .b(gate55inter6), .O(gate55inter12));
  nand2 gate2072(.a(gate55inter12), .b(gate55inter1), .O(G376));

  xor2  gate1835(.a(G287), .b(G16), .O(gate56inter0));
  nand2 gate1836(.a(gate56inter0), .b(s_184), .O(gate56inter1));
  and2  gate1837(.a(G287), .b(G16), .O(gate56inter2));
  inv1  gate1838(.a(s_184), .O(gate56inter3));
  inv1  gate1839(.a(s_185), .O(gate56inter4));
  nand2 gate1840(.a(gate56inter4), .b(gate56inter3), .O(gate56inter5));
  nor2  gate1841(.a(gate56inter5), .b(gate56inter2), .O(gate56inter6));
  inv1  gate1842(.a(G16), .O(gate56inter7));
  inv1  gate1843(.a(G287), .O(gate56inter8));
  nand2 gate1844(.a(gate56inter8), .b(gate56inter7), .O(gate56inter9));
  nand2 gate1845(.a(s_185), .b(gate56inter3), .O(gate56inter10));
  nor2  gate1846(.a(gate56inter10), .b(gate56inter9), .O(gate56inter11));
  nor2  gate1847(.a(gate56inter11), .b(gate56inter6), .O(gate56inter12));
  nand2 gate1848(.a(gate56inter12), .b(gate56inter1), .O(G377));
nand2 gate57( .a(G17), .b(G290), .O(G378) );
nand2 gate58( .a(G18), .b(G290), .O(G379) );
nand2 gate59( .a(G19), .b(G293), .O(G380) );

  xor2  gate1947(.a(G293), .b(G20), .O(gate60inter0));
  nand2 gate1948(.a(gate60inter0), .b(s_200), .O(gate60inter1));
  and2  gate1949(.a(G293), .b(G20), .O(gate60inter2));
  inv1  gate1950(.a(s_200), .O(gate60inter3));
  inv1  gate1951(.a(s_201), .O(gate60inter4));
  nand2 gate1952(.a(gate60inter4), .b(gate60inter3), .O(gate60inter5));
  nor2  gate1953(.a(gate60inter5), .b(gate60inter2), .O(gate60inter6));
  inv1  gate1954(.a(G20), .O(gate60inter7));
  inv1  gate1955(.a(G293), .O(gate60inter8));
  nand2 gate1956(.a(gate60inter8), .b(gate60inter7), .O(gate60inter9));
  nand2 gate1957(.a(s_201), .b(gate60inter3), .O(gate60inter10));
  nor2  gate1958(.a(gate60inter10), .b(gate60inter9), .O(gate60inter11));
  nor2  gate1959(.a(gate60inter11), .b(gate60inter6), .O(gate60inter12));
  nand2 gate1960(.a(gate60inter12), .b(gate60inter1), .O(G381));
nand2 gate61( .a(G21), .b(G296), .O(G382) );
nand2 gate62( .a(G22), .b(G296), .O(G383) );
nand2 gate63( .a(G23), .b(G299), .O(G384) );
nand2 gate64( .a(G24), .b(G299), .O(G385) );

  xor2  gate2801(.a(G302), .b(G25), .O(gate65inter0));
  nand2 gate2802(.a(gate65inter0), .b(s_322), .O(gate65inter1));
  and2  gate2803(.a(G302), .b(G25), .O(gate65inter2));
  inv1  gate2804(.a(s_322), .O(gate65inter3));
  inv1  gate2805(.a(s_323), .O(gate65inter4));
  nand2 gate2806(.a(gate65inter4), .b(gate65inter3), .O(gate65inter5));
  nor2  gate2807(.a(gate65inter5), .b(gate65inter2), .O(gate65inter6));
  inv1  gate2808(.a(G25), .O(gate65inter7));
  inv1  gate2809(.a(G302), .O(gate65inter8));
  nand2 gate2810(.a(gate65inter8), .b(gate65inter7), .O(gate65inter9));
  nand2 gate2811(.a(s_323), .b(gate65inter3), .O(gate65inter10));
  nor2  gate2812(.a(gate65inter10), .b(gate65inter9), .O(gate65inter11));
  nor2  gate2813(.a(gate65inter11), .b(gate65inter6), .O(gate65inter12));
  nand2 gate2814(.a(gate65inter12), .b(gate65inter1), .O(G386));
nand2 gate66( .a(G26), .b(G302), .O(G387) );

  xor2  gate2045(.a(G305), .b(G27), .O(gate67inter0));
  nand2 gate2046(.a(gate67inter0), .b(s_214), .O(gate67inter1));
  and2  gate2047(.a(G305), .b(G27), .O(gate67inter2));
  inv1  gate2048(.a(s_214), .O(gate67inter3));
  inv1  gate2049(.a(s_215), .O(gate67inter4));
  nand2 gate2050(.a(gate67inter4), .b(gate67inter3), .O(gate67inter5));
  nor2  gate2051(.a(gate67inter5), .b(gate67inter2), .O(gate67inter6));
  inv1  gate2052(.a(G27), .O(gate67inter7));
  inv1  gate2053(.a(G305), .O(gate67inter8));
  nand2 gate2054(.a(gate67inter8), .b(gate67inter7), .O(gate67inter9));
  nand2 gate2055(.a(s_215), .b(gate67inter3), .O(gate67inter10));
  nor2  gate2056(.a(gate67inter10), .b(gate67inter9), .O(gate67inter11));
  nor2  gate2057(.a(gate67inter11), .b(gate67inter6), .O(gate67inter12));
  nand2 gate2058(.a(gate67inter12), .b(gate67inter1), .O(G388));
nand2 gate68( .a(G28), .b(G305), .O(G389) );
nand2 gate69( .a(G29), .b(G308), .O(G390) );
nand2 gate70( .a(G30), .b(G308), .O(G391) );

  xor2  gate1597(.a(G311), .b(G31), .O(gate71inter0));
  nand2 gate1598(.a(gate71inter0), .b(s_150), .O(gate71inter1));
  and2  gate1599(.a(G311), .b(G31), .O(gate71inter2));
  inv1  gate1600(.a(s_150), .O(gate71inter3));
  inv1  gate1601(.a(s_151), .O(gate71inter4));
  nand2 gate1602(.a(gate71inter4), .b(gate71inter3), .O(gate71inter5));
  nor2  gate1603(.a(gate71inter5), .b(gate71inter2), .O(gate71inter6));
  inv1  gate1604(.a(G31), .O(gate71inter7));
  inv1  gate1605(.a(G311), .O(gate71inter8));
  nand2 gate1606(.a(gate71inter8), .b(gate71inter7), .O(gate71inter9));
  nand2 gate1607(.a(s_151), .b(gate71inter3), .O(gate71inter10));
  nor2  gate1608(.a(gate71inter10), .b(gate71inter9), .O(gate71inter11));
  nor2  gate1609(.a(gate71inter11), .b(gate71inter6), .O(gate71inter12));
  nand2 gate1610(.a(gate71inter12), .b(gate71inter1), .O(G392));

  xor2  gate1513(.a(G311), .b(G32), .O(gate72inter0));
  nand2 gate1514(.a(gate72inter0), .b(s_138), .O(gate72inter1));
  and2  gate1515(.a(G311), .b(G32), .O(gate72inter2));
  inv1  gate1516(.a(s_138), .O(gate72inter3));
  inv1  gate1517(.a(s_139), .O(gate72inter4));
  nand2 gate1518(.a(gate72inter4), .b(gate72inter3), .O(gate72inter5));
  nor2  gate1519(.a(gate72inter5), .b(gate72inter2), .O(gate72inter6));
  inv1  gate1520(.a(G32), .O(gate72inter7));
  inv1  gate1521(.a(G311), .O(gate72inter8));
  nand2 gate1522(.a(gate72inter8), .b(gate72inter7), .O(gate72inter9));
  nand2 gate1523(.a(s_139), .b(gate72inter3), .O(gate72inter10));
  nor2  gate1524(.a(gate72inter10), .b(gate72inter9), .O(gate72inter11));
  nor2  gate1525(.a(gate72inter11), .b(gate72inter6), .O(gate72inter12));
  nand2 gate1526(.a(gate72inter12), .b(gate72inter1), .O(G393));
nand2 gate73( .a(G1), .b(G314), .O(G394) );

  xor2  gate2283(.a(G314), .b(G5), .O(gate74inter0));
  nand2 gate2284(.a(gate74inter0), .b(s_248), .O(gate74inter1));
  and2  gate2285(.a(G314), .b(G5), .O(gate74inter2));
  inv1  gate2286(.a(s_248), .O(gate74inter3));
  inv1  gate2287(.a(s_249), .O(gate74inter4));
  nand2 gate2288(.a(gate74inter4), .b(gate74inter3), .O(gate74inter5));
  nor2  gate2289(.a(gate74inter5), .b(gate74inter2), .O(gate74inter6));
  inv1  gate2290(.a(G5), .O(gate74inter7));
  inv1  gate2291(.a(G314), .O(gate74inter8));
  nand2 gate2292(.a(gate74inter8), .b(gate74inter7), .O(gate74inter9));
  nand2 gate2293(.a(s_249), .b(gate74inter3), .O(gate74inter10));
  nor2  gate2294(.a(gate74inter10), .b(gate74inter9), .O(gate74inter11));
  nor2  gate2295(.a(gate74inter11), .b(gate74inter6), .O(gate74inter12));
  nand2 gate2296(.a(gate74inter12), .b(gate74inter1), .O(G395));

  xor2  gate2297(.a(G317), .b(G9), .O(gate75inter0));
  nand2 gate2298(.a(gate75inter0), .b(s_250), .O(gate75inter1));
  and2  gate2299(.a(G317), .b(G9), .O(gate75inter2));
  inv1  gate2300(.a(s_250), .O(gate75inter3));
  inv1  gate2301(.a(s_251), .O(gate75inter4));
  nand2 gate2302(.a(gate75inter4), .b(gate75inter3), .O(gate75inter5));
  nor2  gate2303(.a(gate75inter5), .b(gate75inter2), .O(gate75inter6));
  inv1  gate2304(.a(G9), .O(gate75inter7));
  inv1  gate2305(.a(G317), .O(gate75inter8));
  nand2 gate2306(.a(gate75inter8), .b(gate75inter7), .O(gate75inter9));
  nand2 gate2307(.a(s_251), .b(gate75inter3), .O(gate75inter10));
  nor2  gate2308(.a(gate75inter10), .b(gate75inter9), .O(gate75inter11));
  nor2  gate2309(.a(gate75inter11), .b(gate75inter6), .O(gate75inter12));
  nand2 gate2310(.a(gate75inter12), .b(gate75inter1), .O(G396));
nand2 gate76( .a(G13), .b(G317), .O(G397) );

  xor2  gate2983(.a(G320), .b(G2), .O(gate77inter0));
  nand2 gate2984(.a(gate77inter0), .b(s_348), .O(gate77inter1));
  and2  gate2985(.a(G320), .b(G2), .O(gate77inter2));
  inv1  gate2986(.a(s_348), .O(gate77inter3));
  inv1  gate2987(.a(s_349), .O(gate77inter4));
  nand2 gate2988(.a(gate77inter4), .b(gate77inter3), .O(gate77inter5));
  nor2  gate2989(.a(gate77inter5), .b(gate77inter2), .O(gate77inter6));
  inv1  gate2990(.a(G2), .O(gate77inter7));
  inv1  gate2991(.a(G320), .O(gate77inter8));
  nand2 gate2992(.a(gate77inter8), .b(gate77inter7), .O(gate77inter9));
  nand2 gate2993(.a(s_349), .b(gate77inter3), .O(gate77inter10));
  nor2  gate2994(.a(gate77inter10), .b(gate77inter9), .O(gate77inter11));
  nor2  gate2995(.a(gate77inter11), .b(gate77inter6), .O(gate77inter12));
  nand2 gate2996(.a(gate77inter12), .b(gate77inter1), .O(G398));

  xor2  gate981(.a(G320), .b(G6), .O(gate78inter0));
  nand2 gate982(.a(gate78inter0), .b(s_62), .O(gate78inter1));
  and2  gate983(.a(G320), .b(G6), .O(gate78inter2));
  inv1  gate984(.a(s_62), .O(gate78inter3));
  inv1  gate985(.a(s_63), .O(gate78inter4));
  nand2 gate986(.a(gate78inter4), .b(gate78inter3), .O(gate78inter5));
  nor2  gate987(.a(gate78inter5), .b(gate78inter2), .O(gate78inter6));
  inv1  gate988(.a(G6), .O(gate78inter7));
  inv1  gate989(.a(G320), .O(gate78inter8));
  nand2 gate990(.a(gate78inter8), .b(gate78inter7), .O(gate78inter9));
  nand2 gate991(.a(s_63), .b(gate78inter3), .O(gate78inter10));
  nor2  gate992(.a(gate78inter10), .b(gate78inter9), .O(gate78inter11));
  nor2  gate993(.a(gate78inter11), .b(gate78inter6), .O(gate78inter12));
  nand2 gate994(.a(gate78inter12), .b(gate78inter1), .O(G399));
nand2 gate79( .a(G10), .b(G323), .O(G400) );

  xor2  gate1695(.a(G323), .b(G14), .O(gate80inter0));
  nand2 gate1696(.a(gate80inter0), .b(s_164), .O(gate80inter1));
  and2  gate1697(.a(G323), .b(G14), .O(gate80inter2));
  inv1  gate1698(.a(s_164), .O(gate80inter3));
  inv1  gate1699(.a(s_165), .O(gate80inter4));
  nand2 gate1700(.a(gate80inter4), .b(gate80inter3), .O(gate80inter5));
  nor2  gate1701(.a(gate80inter5), .b(gate80inter2), .O(gate80inter6));
  inv1  gate1702(.a(G14), .O(gate80inter7));
  inv1  gate1703(.a(G323), .O(gate80inter8));
  nand2 gate1704(.a(gate80inter8), .b(gate80inter7), .O(gate80inter9));
  nand2 gate1705(.a(s_165), .b(gate80inter3), .O(gate80inter10));
  nor2  gate1706(.a(gate80inter10), .b(gate80inter9), .O(gate80inter11));
  nor2  gate1707(.a(gate80inter11), .b(gate80inter6), .O(gate80inter12));
  nand2 gate1708(.a(gate80inter12), .b(gate80inter1), .O(G401));

  xor2  gate1877(.a(G326), .b(G3), .O(gate81inter0));
  nand2 gate1878(.a(gate81inter0), .b(s_190), .O(gate81inter1));
  and2  gate1879(.a(G326), .b(G3), .O(gate81inter2));
  inv1  gate1880(.a(s_190), .O(gate81inter3));
  inv1  gate1881(.a(s_191), .O(gate81inter4));
  nand2 gate1882(.a(gate81inter4), .b(gate81inter3), .O(gate81inter5));
  nor2  gate1883(.a(gate81inter5), .b(gate81inter2), .O(gate81inter6));
  inv1  gate1884(.a(G3), .O(gate81inter7));
  inv1  gate1885(.a(G326), .O(gate81inter8));
  nand2 gate1886(.a(gate81inter8), .b(gate81inter7), .O(gate81inter9));
  nand2 gate1887(.a(s_191), .b(gate81inter3), .O(gate81inter10));
  nor2  gate1888(.a(gate81inter10), .b(gate81inter9), .O(gate81inter11));
  nor2  gate1889(.a(gate81inter11), .b(gate81inter6), .O(gate81inter12));
  nand2 gate1890(.a(gate81inter12), .b(gate81inter1), .O(G402));
nand2 gate82( .a(G7), .b(G326), .O(G403) );
nand2 gate83( .a(G11), .b(G329), .O(G404) );
nand2 gate84( .a(G15), .b(G329), .O(G405) );
nand2 gate85( .a(G4), .b(G332), .O(G406) );
nand2 gate86( .a(G8), .b(G332), .O(G407) );

  xor2  gate1793(.a(G335), .b(G12), .O(gate87inter0));
  nand2 gate1794(.a(gate87inter0), .b(s_178), .O(gate87inter1));
  and2  gate1795(.a(G335), .b(G12), .O(gate87inter2));
  inv1  gate1796(.a(s_178), .O(gate87inter3));
  inv1  gate1797(.a(s_179), .O(gate87inter4));
  nand2 gate1798(.a(gate87inter4), .b(gate87inter3), .O(gate87inter5));
  nor2  gate1799(.a(gate87inter5), .b(gate87inter2), .O(gate87inter6));
  inv1  gate1800(.a(G12), .O(gate87inter7));
  inv1  gate1801(.a(G335), .O(gate87inter8));
  nand2 gate1802(.a(gate87inter8), .b(gate87inter7), .O(gate87inter9));
  nand2 gate1803(.a(s_179), .b(gate87inter3), .O(gate87inter10));
  nor2  gate1804(.a(gate87inter10), .b(gate87inter9), .O(gate87inter11));
  nor2  gate1805(.a(gate87inter11), .b(gate87inter6), .O(gate87inter12));
  nand2 gate1806(.a(gate87inter12), .b(gate87inter1), .O(G408));
nand2 gate88( .a(G16), .b(G335), .O(G409) );
nand2 gate89( .a(G17), .b(G338), .O(G410) );
nand2 gate90( .a(G21), .b(G338), .O(G411) );
nand2 gate91( .a(G25), .b(G341), .O(G412) );

  xor2  gate1149(.a(G341), .b(G29), .O(gate92inter0));
  nand2 gate1150(.a(gate92inter0), .b(s_86), .O(gate92inter1));
  and2  gate1151(.a(G341), .b(G29), .O(gate92inter2));
  inv1  gate1152(.a(s_86), .O(gate92inter3));
  inv1  gate1153(.a(s_87), .O(gate92inter4));
  nand2 gate1154(.a(gate92inter4), .b(gate92inter3), .O(gate92inter5));
  nor2  gate1155(.a(gate92inter5), .b(gate92inter2), .O(gate92inter6));
  inv1  gate1156(.a(G29), .O(gate92inter7));
  inv1  gate1157(.a(G341), .O(gate92inter8));
  nand2 gate1158(.a(gate92inter8), .b(gate92inter7), .O(gate92inter9));
  nand2 gate1159(.a(s_87), .b(gate92inter3), .O(gate92inter10));
  nor2  gate1160(.a(gate92inter10), .b(gate92inter9), .O(gate92inter11));
  nor2  gate1161(.a(gate92inter11), .b(gate92inter6), .O(gate92inter12));
  nand2 gate1162(.a(gate92inter12), .b(gate92inter1), .O(G413));
nand2 gate93( .a(G18), .b(G344), .O(G414) );
nand2 gate94( .a(G22), .b(G344), .O(G415) );
nand2 gate95( .a(G26), .b(G347), .O(G416) );

  xor2  gate2493(.a(G347), .b(G30), .O(gate96inter0));
  nand2 gate2494(.a(gate96inter0), .b(s_278), .O(gate96inter1));
  and2  gate2495(.a(G347), .b(G30), .O(gate96inter2));
  inv1  gate2496(.a(s_278), .O(gate96inter3));
  inv1  gate2497(.a(s_279), .O(gate96inter4));
  nand2 gate2498(.a(gate96inter4), .b(gate96inter3), .O(gate96inter5));
  nor2  gate2499(.a(gate96inter5), .b(gate96inter2), .O(gate96inter6));
  inv1  gate2500(.a(G30), .O(gate96inter7));
  inv1  gate2501(.a(G347), .O(gate96inter8));
  nand2 gate2502(.a(gate96inter8), .b(gate96inter7), .O(gate96inter9));
  nand2 gate2503(.a(s_279), .b(gate96inter3), .O(gate96inter10));
  nor2  gate2504(.a(gate96inter10), .b(gate96inter9), .O(gate96inter11));
  nor2  gate2505(.a(gate96inter11), .b(gate96inter6), .O(gate96inter12));
  nand2 gate2506(.a(gate96inter12), .b(gate96inter1), .O(G417));

  xor2  gate911(.a(G350), .b(G19), .O(gate97inter0));
  nand2 gate912(.a(gate97inter0), .b(s_52), .O(gate97inter1));
  and2  gate913(.a(G350), .b(G19), .O(gate97inter2));
  inv1  gate914(.a(s_52), .O(gate97inter3));
  inv1  gate915(.a(s_53), .O(gate97inter4));
  nand2 gate916(.a(gate97inter4), .b(gate97inter3), .O(gate97inter5));
  nor2  gate917(.a(gate97inter5), .b(gate97inter2), .O(gate97inter6));
  inv1  gate918(.a(G19), .O(gate97inter7));
  inv1  gate919(.a(G350), .O(gate97inter8));
  nand2 gate920(.a(gate97inter8), .b(gate97inter7), .O(gate97inter9));
  nand2 gate921(.a(s_53), .b(gate97inter3), .O(gate97inter10));
  nor2  gate922(.a(gate97inter10), .b(gate97inter9), .O(gate97inter11));
  nor2  gate923(.a(gate97inter11), .b(gate97inter6), .O(gate97inter12));
  nand2 gate924(.a(gate97inter12), .b(gate97inter1), .O(G418));
nand2 gate98( .a(G23), .b(G350), .O(G419) );
nand2 gate99( .a(G27), .b(G353), .O(G420) );

  xor2  gate2031(.a(G353), .b(G31), .O(gate100inter0));
  nand2 gate2032(.a(gate100inter0), .b(s_212), .O(gate100inter1));
  and2  gate2033(.a(G353), .b(G31), .O(gate100inter2));
  inv1  gate2034(.a(s_212), .O(gate100inter3));
  inv1  gate2035(.a(s_213), .O(gate100inter4));
  nand2 gate2036(.a(gate100inter4), .b(gate100inter3), .O(gate100inter5));
  nor2  gate2037(.a(gate100inter5), .b(gate100inter2), .O(gate100inter6));
  inv1  gate2038(.a(G31), .O(gate100inter7));
  inv1  gate2039(.a(G353), .O(gate100inter8));
  nand2 gate2040(.a(gate100inter8), .b(gate100inter7), .O(gate100inter9));
  nand2 gate2041(.a(s_213), .b(gate100inter3), .O(gate100inter10));
  nor2  gate2042(.a(gate100inter10), .b(gate100inter9), .O(gate100inter11));
  nor2  gate2043(.a(gate100inter11), .b(gate100inter6), .O(gate100inter12));
  nand2 gate2044(.a(gate100inter12), .b(gate100inter1), .O(G421));

  xor2  gate1975(.a(G356), .b(G20), .O(gate101inter0));
  nand2 gate1976(.a(gate101inter0), .b(s_204), .O(gate101inter1));
  and2  gate1977(.a(G356), .b(G20), .O(gate101inter2));
  inv1  gate1978(.a(s_204), .O(gate101inter3));
  inv1  gate1979(.a(s_205), .O(gate101inter4));
  nand2 gate1980(.a(gate101inter4), .b(gate101inter3), .O(gate101inter5));
  nor2  gate1981(.a(gate101inter5), .b(gate101inter2), .O(gate101inter6));
  inv1  gate1982(.a(G20), .O(gate101inter7));
  inv1  gate1983(.a(G356), .O(gate101inter8));
  nand2 gate1984(.a(gate101inter8), .b(gate101inter7), .O(gate101inter9));
  nand2 gate1985(.a(s_205), .b(gate101inter3), .O(gate101inter10));
  nor2  gate1986(.a(gate101inter10), .b(gate101inter9), .O(gate101inter11));
  nor2  gate1987(.a(gate101inter11), .b(gate101inter6), .O(gate101inter12));
  nand2 gate1988(.a(gate101inter12), .b(gate101inter1), .O(G422));
nand2 gate102( .a(G24), .b(G356), .O(G423) );
nand2 gate103( .a(G28), .b(G359), .O(G424) );
nand2 gate104( .a(G32), .b(G359), .O(G425) );
nand2 gate105( .a(G362), .b(G363), .O(G426) );

  xor2  gate2535(.a(G365), .b(G364), .O(gate106inter0));
  nand2 gate2536(.a(gate106inter0), .b(s_284), .O(gate106inter1));
  and2  gate2537(.a(G365), .b(G364), .O(gate106inter2));
  inv1  gate2538(.a(s_284), .O(gate106inter3));
  inv1  gate2539(.a(s_285), .O(gate106inter4));
  nand2 gate2540(.a(gate106inter4), .b(gate106inter3), .O(gate106inter5));
  nor2  gate2541(.a(gate106inter5), .b(gate106inter2), .O(gate106inter6));
  inv1  gate2542(.a(G364), .O(gate106inter7));
  inv1  gate2543(.a(G365), .O(gate106inter8));
  nand2 gate2544(.a(gate106inter8), .b(gate106inter7), .O(gate106inter9));
  nand2 gate2545(.a(s_285), .b(gate106inter3), .O(gate106inter10));
  nor2  gate2546(.a(gate106inter10), .b(gate106inter9), .O(gate106inter11));
  nor2  gate2547(.a(gate106inter11), .b(gate106inter6), .O(gate106inter12));
  nand2 gate2548(.a(gate106inter12), .b(gate106inter1), .O(G429));
nand2 gate107( .a(G366), .b(G367), .O(G432) );
nand2 gate108( .a(G368), .b(G369), .O(G435) );

  xor2  gate1023(.a(G371), .b(G370), .O(gate109inter0));
  nand2 gate1024(.a(gate109inter0), .b(s_68), .O(gate109inter1));
  and2  gate1025(.a(G371), .b(G370), .O(gate109inter2));
  inv1  gate1026(.a(s_68), .O(gate109inter3));
  inv1  gate1027(.a(s_69), .O(gate109inter4));
  nand2 gate1028(.a(gate109inter4), .b(gate109inter3), .O(gate109inter5));
  nor2  gate1029(.a(gate109inter5), .b(gate109inter2), .O(gate109inter6));
  inv1  gate1030(.a(G370), .O(gate109inter7));
  inv1  gate1031(.a(G371), .O(gate109inter8));
  nand2 gate1032(.a(gate109inter8), .b(gate109inter7), .O(gate109inter9));
  nand2 gate1033(.a(s_69), .b(gate109inter3), .O(gate109inter10));
  nor2  gate1034(.a(gate109inter10), .b(gate109inter9), .O(gate109inter11));
  nor2  gate1035(.a(gate109inter11), .b(gate109inter6), .O(gate109inter12));
  nand2 gate1036(.a(gate109inter12), .b(gate109inter1), .O(G438));
nand2 gate110( .a(G372), .b(G373), .O(G441) );
nand2 gate111( .a(G374), .b(G375), .O(G444) );

  xor2  gate1681(.a(G377), .b(G376), .O(gate112inter0));
  nand2 gate1682(.a(gate112inter0), .b(s_162), .O(gate112inter1));
  and2  gate1683(.a(G377), .b(G376), .O(gate112inter2));
  inv1  gate1684(.a(s_162), .O(gate112inter3));
  inv1  gate1685(.a(s_163), .O(gate112inter4));
  nand2 gate1686(.a(gate112inter4), .b(gate112inter3), .O(gate112inter5));
  nor2  gate1687(.a(gate112inter5), .b(gate112inter2), .O(gate112inter6));
  inv1  gate1688(.a(G376), .O(gate112inter7));
  inv1  gate1689(.a(G377), .O(gate112inter8));
  nand2 gate1690(.a(gate112inter8), .b(gate112inter7), .O(gate112inter9));
  nand2 gate1691(.a(s_163), .b(gate112inter3), .O(gate112inter10));
  nor2  gate1692(.a(gate112inter10), .b(gate112inter9), .O(gate112inter11));
  nor2  gate1693(.a(gate112inter11), .b(gate112inter6), .O(gate112inter12));
  nand2 gate1694(.a(gate112inter12), .b(gate112inter1), .O(G447));
nand2 gate113( .a(G378), .b(G379), .O(G450) );

  xor2  gate1289(.a(G381), .b(G380), .O(gate114inter0));
  nand2 gate1290(.a(gate114inter0), .b(s_106), .O(gate114inter1));
  and2  gate1291(.a(G381), .b(G380), .O(gate114inter2));
  inv1  gate1292(.a(s_106), .O(gate114inter3));
  inv1  gate1293(.a(s_107), .O(gate114inter4));
  nand2 gate1294(.a(gate114inter4), .b(gate114inter3), .O(gate114inter5));
  nor2  gate1295(.a(gate114inter5), .b(gate114inter2), .O(gate114inter6));
  inv1  gate1296(.a(G380), .O(gate114inter7));
  inv1  gate1297(.a(G381), .O(gate114inter8));
  nand2 gate1298(.a(gate114inter8), .b(gate114inter7), .O(gate114inter9));
  nand2 gate1299(.a(s_107), .b(gate114inter3), .O(gate114inter10));
  nor2  gate1300(.a(gate114inter10), .b(gate114inter9), .O(gate114inter11));
  nor2  gate1301(.a(gate114inter11), .b(gate114inter6), .O(gate114inter12));
  nand2 gate1302(.a(gate114inter12), .b(gate114inter1), .O(G453));

  xor2  gate1121(.a(G383), .b(G382), .O(gate115inter0));
  nand2 gate1122(.a(gate115inter0), .b(s_82), .O(gate115inter1));
  and2  gate1123(.a(G383), .b(G382), .O(gate115inter2));
  inv1  gate1124(.a(s_82), .O(gate115inter3));
  inv1  gate1125(.a(s_83), .O(gate115inter4));
  nand2 gate1126(.a(gate115inter4), .b(gate115inter3), .O(gate115inter5));
  nor2  gate1127(.a(gate115inter5), .b(gate115inter2), .O(gate115inter6));
  inv1  gate1128(.a(G382), .O(gate115inter7));
  inv1  gate1129(.a(G383), .O(gate115inter8));
  nand2 gate1130(.a(gate115inter8), .b(gate115inter7), .O(gate115inter9));
  nand2 gate1131(.a(s_83), .b(gate115inter3), .O(gate115inter10));
  nor2  gate1132(.a(gate115inter10), .b(gate115inter9), .O(gate115inter11));
  nor2  gate1133(.a(gate115inter11), .b(gate115inter6), .O(gate115inter12));
  nand2 gate1134(.a(gate115inter12), .b(gate115inter1), .O(G456));

  xor2  gate1135(.a(G385), .b(G384), .O(gate116inter0));
  nand2 gate1136(.a(gate116inter0), .b(s_84), .O(gate116inter1));
  and2  gate1137(.a(G385), .b(G384), .O(gate116inter2));
  inv1  gate1138(.a(s_84), .O(gate116inter3));
  inv1  gate1139(.a(s_85), .O(gate116inter4));
  nand2 gate1140(.a(gate116inter4), .b(gate116inter3), .O(gate116inter5));
  nor2  gate1141(.a(gate116inter5), .b(gate116inter2), .O(gate116inter6));
  inv1  gate1142(.a(G384), .O(gate116inter7));
  inv1  gate1143(.a(G385), .O(gate116inter8));
  nand2 gate1144(.a(gate116inter8), .b(gate116inter7), .O(gate116inter9));
  nand2 gate1145(.a(s_85), .b(gate116inter3), .O(gate116inter10));
  nor2  gate1146(.a(gate116inter10), .b(gate116inter9), .O(gate116inter11));
  nor2  gate1147(.a(gate116inter11), .b(gate116inter6), .O(gate116inter12));
  nand2 gate1148(.a(gate116inter12), .b(gate116inter1), .O(G459));
nand2 gate117( .a(G386), .b(G387), .O(G462) );

  xor2  gate2633(.a(G389), .b(G388), .O(gate118inter0));
  nand2 gate2634(.a(gate118inter0), .b(s_298), .O(gate118inter1));
  and2  gate2635(.a(G389), .b(G388), .O(gate118inter2));
  inv1  gate2636(.a(s_298), .O(gate118inter3));
  inv1  gate2637(.a(s_299), .O(gate118inter4));
  nand2 gate2638(.a(gate118inter4), .b(gate118inter3), .O(gate118inter5));
  nor2  gate2639(.a(gate118inter5), .b(gate118inter2), .O(gate118inter6));
  inv1  gate2640(.a(G388), .O(gate118inter7));
  inv1  gate2641(.a(G389), .O(gate118inter8));
  nand2 gate2642(.a(gate118inter8), .b(gate118inter7), .O(gate118inter9));
  nand2 gate2643(.a(s_299), .b(gate118inter3), .O(gate118inter10));
  nor2  gate2644(.a(gate118inter10), .b(gate118inter9), .O(gate118inter11));
  nor2  gate2645(.a(gate118inter11), .b(gate118inter6), .O(gate118inter12));
  nand2 gate2646(.a(gate118inter12), .b(gate118inter1), .O(G465));
nand2 gate119( .a(G390), .b(G391), .O(G468) );

  xor2  gate2129(.a(G393), .b(G392), .O(gate120inter0));
  nand2 gate2130(.a(gate120inter0), .b(s_226), .O(gate120inter1));
  and2  gate2131(.a(G393), .b(G392), .O(gate120inter2));
  inv1  gate2132(.a(s_226), .O(gate120inter3));
  inv1  gate2133(.a(s_227), .O(gate120inter4));
  nand2 gate2134(.a(gate120inter4), .b(gate120inter3), .O(gate120inter5));
  nor2  gate2135(.a(gate120inter5), .b(gate120inter2), .O(gate120inter6));
  inv1  gate2136(.a(G392), .O(gate120inter7));
  inv1  gate2137(.a(G393), .O(gate120inter8));
  nand2 gate2138(.a(gate120inter8), .b(gate120inter7), .O(gate120inter9));
  nand2 gate2139(.a(s_227), .b(gate120inter3), .O(gate120inter10));
  nor2  gate2140(.a(gate120inter10), .b(gate120inter9), .O(gate120inter11));
  nor2  gate2141(.a(gate120inter11), .b(gate120inter6), .O(gate120inter12));
  nand2 gate2142(.a(gate120inter12), .b(gate120inter1), .O(G471));

  xor2  gate1345(.a(G395), .b(G394), .O(gate121inter0));
  nand2 gate1346(.a(gate121inter0), .b(s_114), .O(gate121inter1));
  and2  gate1347(.a(G395), .b(G394), .O(gate121inter2));
  inv1  gate1348(.a(s_114), .O(gate121inter3));
  inv1  gate1349(.a(s_115), .O(gate121inter4));
  nand2 gate1350(.a(gate121inter4), .b(gate121inter3), .O(gate121inter5));
  nor2  gate1351(.a(gate121inter5), .b(gate121inter2), .O(gate121inter6));
  inv1  gate1352(.a(G394), .O(gate121inter7));
  inv1  gate1353(.a(G395), .O(gate121inter8));
  nand2 gate1354(.a(gate121inter8), .b(gate121inter7), .O(gate121inter9));
  nand2 gate1355(.a(s_115), .b(gate121inter3), .O(gate121inter10));
  nor2  gate1356(.a(gate121inter10), .b(gate121inter9), .O(gate121inter11));
  nor2  gate1357(.a(gate121inter11), .b(gate121inter6), .O(gate121inter12));
  nand2 gate1358(.a(gate121inter12), .b(gate121inter1), .O(G474));
nand2 gate122( .a(G396), .b(G397), .O(G477) );

  xor2  gate1275(.a(G399), .b(G398), .O(gate123inter0));
  nand2 gate1276(.a(gate123inter0), .b(s_104), .O(gate123inter1));
  and2  gate1277(.a(G399), .b(G398), .O(gate123inter2));
  inv1  gate1278(.a(s_104), .O(gate123inter3));
  inv1  gate1279(.a(s_105), .O(gate123inter4));
  nand2 gate1280(.a(gate123inter4), .b(gate123inter3), .O(gate123inter5));
  nor2  gate1281(.a(gate123inter5), .b(gate123inter2), .O(gate123inter6));
  inv1  gate1282(.a(G398), .O(gate123inter7));
  inv1  gate1283(.a(G399), .O(gate123inter8));
  nand2 gate1284(.a(gate123inter8), .b(gate123inter7), .O(gate123inter9));
  nand2 gate1285(.a(s_105), .b(gate123inter3), .O(gate123inter10));
  nor2  gate1286(.a(gate123inter10), .b(gate123inter9), .O(gate123inter11));
  nor2  gate1287(.a(gate123inter11), .b(gate123inter6), .O(gate123inter12));
  nand2 gate1288(.a(gate123inter12), .b(gate123inter1), .O(G480));
nand2 gate124( .a(G400), .b(G401), .O(G483) );

  xor2  gate547(.a(G403), .b(G402), .O(gate125inter0));
  nand2 gate548(.a(gate125inter0), .b(s_0), .O(gate125inter1));
  and2  gate549(.a(G403), .b(G402), .O(gate125inter2));
  inv1  gate550(.a(s_0), .O(gate125inter3));
  inv1  gate551(.a(s_1), .O(gate125inter4));
  nand2 gate552(.a(gate125inter4), .b(gate125inter3), .O(gate125inter5));
  nor2  gate553(.a(gate125inter5), .b(gate125inter2), .O(gate125inter6));
  inv1  gate554(.a(G402), .O(gate125inter7));
  inv1  gate555(.a(G403), .O(gate125inter8));
  nand2 gate556(.a(gate125inter8), .b(gate125inter7), .O(gate125inter9));
  nand2 gate557(.a(s_1), .b(gate125inter3), .O(gate125inter10));
  nor2  gate558(.a(gate125inter10), .b(gate125inter9), .O(gate125inter11));
  nor2  gate559(.a(gate125inter11), .b(gate125inter6), .O(gate125inter12));
  nand2 gate560(.a(gate125inter12), .b(gate125inter1), .O(G486));

  xor2  gate2185(.a(G405), .b(G404), .O(gate126inter0));
  nand2 gate2186(.a(gate126inter0), .b(s_234), .O(gate126inter1));
  and2  gate2187(.a(G405), .b(G404), .O(gate126inter2));
  inv1  gate2188(.a(s_234), .O(gate126inter3));
  inv1  gate2189(.a(s_235), .O(gate126inter4));
  nand2 gate2190(.a(gate126inter4), .b(gate126inter3), .O(gate126inter5));
  nor2  gate2191(.a(gate126inter5), .b(gate126inter2), .O(gate126inter6));
  inv1  gate2192(.a(G404), .O(gate126inter7));
  inv1  gate2193(.a(G405), .O(gate126inter8));
  nand2 gate2194(.a(gate126inter8), .b(gate126inter7), .O(gate126inter9));
  nand2 gate2195(.a(s_235), .b(gate126inter3), .O(gate126inter10));
  nor2  gate2196(.a(gate126inter10), .b(gate126inter9), .O(gate126inter11));
  nor2  gate2197(.a(gate126inter11), .b(gate126inter6), .O(gate126inter12));
  nand2 gate2198(.a(gate126inter12), .b(gate126inter1), .O(G489));

  xor2  gate589(.a(G407), .b(G406), .O(gate127inter0));
  nand2 gate590(.a(gate127inter0), .b(s_6), .O(gate127inter1));
  and2  gate591(.a(G407), .b(G406), .O(gate127inter2));
  inv1  gate592(.a(s_6), .O(gate127inter3));
  inv1  gate593(.a(s_7), .O(gate127inter4));
  nand2 gate594(.a(gate127inter4), .b(gate127inter3), .O(gate127inter5));
  nor2  gate595(.a(gate127inter5), .b(gate127inter2), .O(gate127inter6));
  inv1  gate596(.a(G406), .O(gate127inter7));
  inv1  gate597(.a(G407), .O(gate127inter8));
  nand2 gate598(.a(gate127inter8), .b(gate127inter7), .O(gate127inter9));
  nand2 gate599(.a(s_7), .b(gate127inter3), .O(gate127inter10));
  nor2  gate600(.a(gate127inter10), .b(gate127inter9), .O(gate127inter11));
  nor2  gate601(.a(gate127inter11), .b(gate127inter6), .O(gate127inter12));
  nand2 gate602(.a(gate127inter12), .b(gate127inter1), .O(G492));
nand2 gate128( .a(G408), .b(G409), .O(G495) );

  xor2  gate967(.a(G411), .b(G410), .O(gate129inter0));
  nand2 gate968(.a(gate129inter0), .b(s_60), .O(gate129inter1));
  and2  gate969(.a(G411), .b(G410), .O(gate129inter2));
  inv1  gate970(.a(s_60), .O(gate129inter3));
  inv1  gate971(.a(s_61), .O(gate129inter4));
  nand2 gate972(.a(gate129inter4), .b(gate129inter3), .O(gate129inter5));
  nor2  gate973(.a(gate129inter5), .b(gate129inter2), .O(gate129inter6));
  inv1  gate974(.a(G410), .O(gate129inter7));
  inv1  gate975(.a(G411), .O(gate129inter8));
  nand2 gate976(.a(gate129inter8), .b(gate129inter7), .O(gate129inter9));
  nand2 gate977(.a(s_61), .b(gate129inter3), .O(gate129inter10));
  nor2  gate978(.a(gate129inter10), .b(gate129inter9), .O(gate129inter11));
  nor2  gate979(.a(gate129inter11), .b(gate129inter6), .O(gate129inter12));
  nand2 gate980(.a(gate129inter12), .b(gate129inter1), .O(G498));
nand2 gate130( .a(G412), .b(G413), .O(G501) );
nand2 gate131( .a(G414), .b(G415), .O(G504) );

  xor2  gate2115(.a(G417), .b(G416), .O(gate132inter0));
  nand2 gate2116(.a(gate132inter0), .b(s_224), .O(gate132inter1));
  and2  gate2117(.a(G417), .b(G416), .O(gate132inter2));
  inv1  gate2118(.a(s_224), .O(gate132inter3));
  inv1  gate2119(.a(s_225), .O(gate132inter4));
  nand2 gate2120(.a(gate132inter4), .b(gate132inter3), .O(gate132inter5));
  nor2  gate2121(.a(gate132inter5), .b(gate132inter2), .O(gate132inter6));
  inv1  gate2122(.a(G416), .O(gate132inter7));
  inv1  gate2123(.a(G417), .O(gate132inter8));
  nand2 gate2124(.a(gate132inter8), .b(gate132inter7), .O(gate132inter9));
  nand2 gate2125(.a(s_225), .b(gate132inter3), .O(gate132inter10));
  nor2  gate2126(.a(gate132inter10), .b(gate132inter9), .O(gate132inter11));
  nor2  gate2127(.a(gate132inter11), .b(gate132inter6), .O(gate132inter12));
  nand2 gate2128(.a(gate132inter12), .b(gate132inter1), .O(G507));
nand2 gate133( .a(G418), .b(G419), .O(G510) );

  xor2  gate2843(.a(G421), .b(G420), .O(gate134inter0));
  nand2 gate2844(.a(gate134inter0), .b(s_328), .O(gate134inter1));
  and2  gate2845(.a(G421), .b(G420), .O(gate134inter2));
  inv1  gate2846(.a(s_328), .O(gate134inter3));
  inv1  gate2847(.a(s_329), .O(gate134inter4));
  nand2 gate2848(.a(gate134inter4), .b(gate134inter3), .O(gate134inter5));
  nor2  gate2849(.a(gate134inter5), .b(gate134inter2), .O(gate134inter6));
  inv1  gate2850(.a(G420), .O(gate134inter7));
  inv1  gate2851(.a(G421), .O(gate134inter8));
  nand2 gate2852(.a(gate134inter8), .b(gate134inter7), .O(gate134inter9));
  nand2 gate2853(.a(s_329), .b(gate134inter3), .O(gate134inter10));
  nor2  gate2854(.a(gate134inter10), .b(gate134inter9), .O(gate134inter11));
  nor2  gate2855(.a(gate134inter11), .b(gate134inter6), .O(gate134inter12));
  nand2 gate2856(.a(gate134inter12), .b(gate134inter1), .O(G513));

  xor2  gate2745(.a(G423), .b(G422), .O(gate135inter0));
  nand2 gate2746(.a(gate135inter0), .b(s_314), .O(gate135inter1));
  and2  gate2747(.a(G423), .b(G422), .O(gate135inter2));
  inv1  gate2748(.a(s_314), .O(gate135inter3));
  inv1  gate2749(.a(s_315), .O(gate135inter4));
  nand2 gate2750(.a(gate135inter4), .b(gate135inter3), .O(gate135inter5));
  nor2  gate2751(.a(gate135inter5), .b(gate135inter2), .O(gate135inter6));
  inv1  gate2752(.a(G422), .O(gate135inter7));
  inv1  gate2753(.a(G423), .O(gate135inter8));
  nand2 gate2754(.a(gate135inter8), .b(gate135inter7), .O(gate135inter9));
  nand2 gate2755(.a(s_315), .b(gate135inter3), .O(gate135inter10));
  nor2  gate2756(.a(gate135inter10), .b(gate135inter9), .O(gate135inter11));
  nor2  gate2757(.a(gate135inter11), .b(gate135inter6), .O(gate135inter12));
  nand2 gate2758(.a(gate135inter12), .b(gate135inter1), .O(G516));

  xor2  gate1583(.a(G425), .b(G424), .O(gate136inter0));
  nand2 gate1584(.a(gate136inter0), .b(s_148), .O(gate136inter1));
  and2  gate1585(.a(G425), .b(G424), .O(gate136inter2));
  inv1  gate1586(.a(s_148), .O(gate136inter3));
  inv1  gate1587(.a(s_149), .O(gate136inter4));
  nand2 gate1588(.a(gate136inter4), .b(gate136inter3), .O(gate136inter5));
  nor2  gate1589(.a(gate136inter5), .b(gate136inter2), .O(gate136inter6));
  inv1  gate1590(.a(G424), .O(gate136inter7));
  inv1  gate1591(.a(G425), .O(gate136inter8));
  nand2 gate1592(.a(gate136inter8), .b(gate136inter7), .O(gate136inter9));
  nand2 gate1593(.a(s_149), .b(gate136inter3), .O(gate136inter10));
  nor2  gate1594(.a(gate136inter10), .b(gate136inter9), .O(gate136inter11));
  nor2  gate1595(.a(gate136inter11), .b(gate136inter6), .O(gate136inter12));
  nand2 gate1596(.a(gate136inter12), .b(gate136inter1), .O(G519));
nand2 gate137( .a(G426), .b(G429), .O(G522) );

  xor2  gate2017(.a(G435), .b(G432), .O(gate138inter0));
  nand2 gate2018(.a(gate138inter0), .b(s_210), .O(gate138inter1));
  and2  gate2019(.a(G435), .b(G432), .O(gate138inter2));
  inv1  gate2020(.a(s_210), .O(gate138inter3));
  inv1  gate2021(.a(s_211), .O(gate138inter4));
  nand2 gate2022(.a(gate138inter4), .b(gate138inter3), .O(gate138inter5));
  nor2  gate2023(.a(gate138inter5), .b(gate138inter2), .O(gate138inter6));
  inv1  gate2024(.a(G432), .O(gate138inter7));
  inv1  gate2025(.a(G435), .O(gate138inter8));
  nand2 gate2026(.a(gate138inter8), .b(gate138inter7), .O(gate138inter9));
  nand2 gate2027(.a(s_211), .b(gate138inter3), .O(gate138inter10));
  nor2  gate2028(.a(gate138inter10), .b(gate138inter9), .O(gate138inter11));
  nor2  gate2029(.a(gate138inter11), .b(gate138inter6), .O(gate138inter12));
  nand2 gate2030(.a(gate138inter12), .b(gate138inter1), .O(G525));
nand2 gate139( .a(G438), .b(G441), .O(G528) );
nand2 gate140( .a(G444), .b(G447), .O(G531) );
nand2 gate141( .a(G450), .b(G453), .O(G534) );
nand2 gate142( .a(G456), .b(G459), .O(G537) );
nand2 gate143( .a(G462), .b(G465), .O(G540) );
nand2 gate144( .a(G468), .b(G471), .O(G543) );

  xor2  gate2647(.a(G477), .b(G474), .O(gate145inter0));
  nand2 gate2648(.a(gate145inter0), .b(s_300), .O(gate145inter1));
  and2  gate2649(.a(G477), .b(G474), .O(gate145inter2));
  inv1  gate2650(.a(s_300), .O(gate145inter3));
  inv1  gate2651(.a(s_301), .O(gate145inter4));
  nand2 gate2652(.a(gate145inter4), .b(gate145inter3), .O(gate145inter5));
  nor2  gate2653(.a(gate145inter5), .b(gate145inter2), .O(gate145inter6));
  inv1  gate2654(.a(G474), .O(gate145inter7));
  inv1  gate2655(.a(G477), .O(gate145inter8));
  nand2 gate2656(.a(gate145inter8), .b(gate145inter7), .O(gate145inter9));
  nand2 gate2657(.a(s_301), .b(gate145inter3), .O(gate145inter10));
  nor2  gate2658(.a(gate145inter10), .b(gate145inter9), .O(gate145inter11));
  nor2  gate2659(.a(gate145inter11), .b(gate145inter6), .O(gate145inter12));
  nand2 gate2660(.a(gate145inter12), .b(gate145inter1), .O(G546));
nand2 gate146( .a(G480), .b(G483), .O(G549) );

  xor2  gate729(.a(G489), .b(G486), .O(gate147inter0));
  nand2 gate730(.a(gate147inter0), .b(s_26), .O(gate147inter1));
  and2  gate731(.a(G489), .b(G486), .O(gate147inter2));
  inv1  gate732(.a(s_26), .O(gate147inter3));
  inv1  gate733(.a(s_27), .O(gate147inter4));
  nand2 gate734(.a(gate147inter4), .b(gate147inter3), .O(gate147inter5));
  nor2  gate735(.a(gate147inter5), .b(gate147inter2), .O(gate147inter6));
  inv1  gate736(.a(G486), .O(gate147inter7));
  inv1  gate737(.a(G489), .O(gate147inter8));
  nand2 gate738(.a(gate147inter8), .b(gate147inter7), .O(gate147inter9));
  nand2 gate739(.a(s_27), .b(gate147inter3), .O(gate147inter10));
  nor2  gate740(.a(gate147inter10), .b(gate147inter9), .O(gate147inter11));
  nor2  gate741(.a(gate147inter11), .b(gate147inter6), .O(gate147inter12));
  nand2 gate742(.a(gate147inter12), .b(gate147inter1), .O(G552));

  xor2  gate2885(.a(G495), .b(G492), .O(gate148inter0));
  nand2 gate2886(.a(gate148inter0), .b(s_334), .O(gate148inter1));
  and2  gate2887(.a(G495), .b(G492), .O(gate148inter2));
  inv1  gate2888(.a(s_334), .O(gate148inter3));
  inv1  gate2889(.a(s_335), .O(gate148inter4));
  nand2 gate2890(.a(gate148inter4), .b(gate148inter3), .O(gate148inter5));
  nor2  gate2891(.a(gate148inter5), .b(gate148inter2), .O(gate148inter6));
  inv1  gate2892(.a(G492), .O(gate148inter7));
  inv1  gate2893(.a(G495), .O(gate148inter8));
  nand2 gate2894(.a(gate148inter8), .b(gate148inter7), .O(gate148inter9));
  nand2 gate2895(.a(s_335), .b(gate148inter3), .O(gate148inter10));
  nor2  gate2896(.a(gate148inter10), .b(gate148inter9), .O(gate148inter11));
  nor2  gate2897(.a(gate148inter11), .b(gate148inter6), .O(gate148inter12));
  nand2 gate2898(.a(gate148inter12), .b(gate148inter1), .O(G555));
nand2 gate149( .a(G498), .b(G501), .O(G558) );
nand2 gate150( .a(G504), .b(G507), .O(G561) );

  xor2  gate1485(.a(G513), .b(G510), .O(gate151inter0));
  nand2 gate1486(.a(gate151inter0), .b(s_134), .O(gate151inter1));
  and2  gate1487(.a(G513), .b(G510), .O(gate151inter2));
  inv1  gate1488(.a(s_134), .O(gate151inter3));
  inv1  gate1489(.a(s_135), .O(gate151inter4));
  nand2 gate1490(.a(gate151inter4), .b(gate151inter3), .O(gate151inter5));
  nor2  gate1491(.a(gate151inter5), .b(gate151inter2), .O(gate151inter6));
  inv1  gate1492(.a(G510), .O(gate151inter7));
  inv1  gate1493(.a(G513), .O(gate151inter8));
  nand2 gate1494(.a(gate151inter8), .b(gate151inter7), .O(gate151inter9));
  nand2 gate1495(.a(s_135), .b(gate151inter3), .O(gate151inter10));
  nor2  gate1496(.a(gate151inter10), .b(gate151inter9), .O(gate151inter11));
  nor2  gate1497(.a(gate151inter11), .b(gate151inter6), .O(gate151inter12));
  nand2 gate1498(.a(gate151inter12), .b(gate151inter1), .O(G564));
nand2 gate152( .a(G516), .b(G519), .O(G567) );
nand2 gate153( .a(G426), .b(G522), .O(G570) );

  xor2  gate1191(.a(G522), .b(G429), .O(gate154inter0));
  nand2 gate1192(.a(gate154inter0), .b(s_92), .O(gate154inter1));
  and2  gate1193(.a(G522), .b(G429), .O(gate154inter2));
  inv1  gate1194(.a(s_92), .O(gate154inter3));
  inv1  gate1195(.a(s_93), .O(gate154inter4));
  nand2 gate1196(.a(gate154inter4), .b(gate154inter3), .O(gate154inter5));
  nor2  gate1197(.a(gate154inter5), .b(gate154inter2), .O(gate154inter6));
  inv1  gate1198(.a(G429), .O(gate154inter7));
  inv1  gate1199(.a(G522), .O(gate154inter8));
  nand2 gate1200(.a(gate154inter8), .b(gate154inter7), .O(gate154inter9));
  nand2 gate1201(.a(s_93), .b(gate154inter3), .O(gate154inter10));
  nor2  gate1202(.a(gate154inter10), .b(gate154inter9), .O(gate154inter11));
  nor2  gate1203(.a(gate154inter11), .b(gate154inter6), .O(gate154inter12));
  nand2 gate1204(.a(gate154inter12), .b(gate154inter1), .O(G571));

  xor2  gate883(.a(G525), .b(G432), .O(gate155inter0));
  nand2 gate884(.a(gate155inter0), .b(s_48), .O(gate155inter1));
  and2  gate885(.a(G525), .b(G432), .O(gate155inter2));
  inv1  gate886(.a(s_48), .O(gate155inter3));
  inv1  gate887(.a(s_49), .O(gate155inter4));
  nand2 gate888(.a(gate155inter4), .b(gate155inter3), .O(gate155inter5));
  nor2  gate889(.a(gate155inter5), .b(gate155inter2), .O(gate155inter6));
  inv1  gate890(.a(G432), .O(gate155inter7));
  inv1  gate891(.a(G525), .O(gate155inter8));
  nand2 gate892(.a(gate155inter8), .b(gate155inter7), .O(gate155inter9));
  nand2 gate893(.a(s_49), .b(gate155inter3), .O(gate155inter10));
  nor2  gate894(.a(gate155inter10), .b(gate155inter9), .O(gate155inter11));
  nor2  gate895(.a(gate155inter11), .b(gate155inter6), .O(gate155inter12));
  nand2 gate896(.a(gate155inter12), .b(gate155inter1), .O(G572));

  xor2  gate2857(.a(G525), .b(G435), .O(gate156inter0));
  nand2 gate2858(.a(gate156inter0), .b(s_330), .O(gate156inter1));
  and2  gate2859(.a(G525), .b(G435), .O(gate156inter2));
  inv1  gate2860(.a(s_330), .O(gate156inter3));
  inv1  gate2861(.a(s_331), .O(gate156inter4));
  nand2 gate2862(.a(gate156inter4), .b(gate156inter3), .O(gate156inter5));
  nor2  gate2863(.a(gate156inter5), .b(gate156inter2), .O(gate156inter6));
  inv1  gate2864(.a(G435), .O(gate156inter7));
  inv1  gate2865(.a(G525), .O(gate156inter8));
  nand2 gate2866(.a(gate156inter8), .b(gate156inter7), .O(gate156inter9));
  nand2 gate2867(.a(s_331), .b(gate156inter3), .O(gate156inter10));
  nor2  gate2868(.a(gate156inter10), .b(gate156inter9), .O(gate156inter11));
  nor2  gate2869(.a(gate156inter11), .b(gate156inter6), .O(gate156inter12));
  nand2 gate2870(.a(gate156inter12), .b(gate156inter1), .O(G573));
nand2 gate157( .a(G438), .b(G528), .O(G574) );
nand2 gate158( .a(G441), .b(G528), .O(G575) );

  xor2  gate1541(.a(G531), .b(G444), .O(gate159inter0));
  nand2 gate1542(.a(gate159inter0), .b(s_142), .O(gate159inter1));
  and2  gate1543(.a(G531), .b(G444), .O(gate159inter2));
  inv1  gate1544(.a(s_142), .O(gate159inter3));
  inv1  gate1545(.a(s_143), .O(gate159inter4));
  nand2 gate1546(.a(gate159inter4), .b(gate159inter3), .O(gate159inter5));
  nor2  gate1547(.a(gate159inter5), .b(gate159inter2), .O(gate159inter6));
  inv1  gate1548(.a(G444), .O(gate159inter7));
  inv1  gate1549(.a(G531), .O(gate159inter8));
  nand2 gate1550(.a(gate159inter8), .b(gate159inter7), .O(gate159inter9));
  nand2 gate1551(.a(s_143), .b(gate159inter3), .O(gate159inter10));
  nor2  gate1552(.a(gate159inter10), .b(gate159inter9), .O(gate159inter11));
  nor2  gate1553(.a(gate159inter11), .b(gate159inter6), .O(gate159inter12));
  nand2 gate1554(.a(gate159inter12), .b(gate159inter1), .O(G576));
nand2 gate160( .a(G447), .b(G531), .O(G577) );

  xor2  gate2325(.a(G534), .b(G450), .O(gate161inter0));
  nand2 gate2326(.a(gate161inter0), .b(s_254), .O(gate161inter1));
  and2  gate2327(.a(G534), .b(G450), .O(gate161inter2));
  inv1  gate2328(.a(s_254), .O(gate161inter3));
  inv1  gate2329(.a(s_255), .O(gate161inter4));
  nand2 gate2330(.a(gate161inter4), .b(gate161inter3), .O(gate161inter5));
  nor2  gate2331(.a(gate161inter5), .b(gate161inter2), .O(gate161inter6));
  inv1  gate2332(.a(G450), .O(gate161inter7));
  inv1  gate2333(.a(G534), .O(gate161inter8));
  nand2 gate2334(.a(gate161inter8), .b(gate161inter7), .O(gate161inter9));
  nand2 gate2335(.a(s_255), .b(gate161inter3), .O(gate161inter10));
  nor2  gate2336(.a(gate161inter10), .b(gate161inter9), .O(gate161inter11));
  nor2  gate2337(.a(gate161inter11), .b(gate161inter6), .O(gate161inter12));
  nand2 gate2338(.a(gate161inter12), .b(gate161inter1), .O(G578));

  xor2  gate827(.a(G534), .b(G453), .O(gate162inter0));
  nand2 gate828(.a(gate162inter0), .b(s_40), .O(gate162inter1));
  and2  gate829(.a(G534), .b(G453), .O(gate162inter2));
  inv1  gate830(.a(s_40), .O(gate162inter3));
  inv1  gate831(.a(s_41), .O(gate162inter4));
  nand2 gate832(.a(gate162inter4), .b(gate162inter3), .O(gate162inter5));
  nor2  gate833(.a(gate162inter5), .b(gate162inter2), .O(gate162inter6));
  inv1  gate834(.a(G453), .O(gate162inter7));
  inv1  gate835(.a(G534), .O(gate162inter8));
  nand2 gate836(.a(gate162inter8), .b(gate162inter7), .O(gate162inter9));
  nand2 gate837(.a(s_41), .b(gate162inter3), .O(gate162inter10));
  nor2  gate838(.a(gate162inter10), .b(gate162inter9), .O(gate162inter11));
  nor2  gate839(.a(gate162inter11), .b(gate162inter6), .O(gate162inter12));
  nand2 gate840(.a(gate162inter12), .b(gate162inter1), .O(G579));
nand2 gate163( .a(G456), .b(G537), .O(G580) );
nand2 gate164( .a(G459), .b(G537), .O(G581) );
nand2 gate165( .a(G462), .b(G540), .O(G582) );

  xor2  gate2689(.a(G540), .b(G465), .O(gate166inter0));
  nand2 gate2690(.a(gate166inter0), .b(s_306), .O(gate166inter1));
  and2  gate2691(.a(G540), .b(G465), .O(gate166inter2));
  inv1  gate2692(.a(s_306), .O(gate166inter3));
  inv1  gate2693(.a(s_307), .O(gate166inter4));
  nand2 gate2694(.a(gate166inter4), .b(gate166inter3), .O(gate166inter5));
  nor2  gate2695(.a(gate166inter5), .b(gate166inter2), .O(gate166inter6));
  inv1  gate2696(.a(G465), .O(gate166inter7));
  inv1  gate2697(.a(G540), .O(gate166inter8));
  nand2 gate2698(.a(gate166inter8), .b(gate166inter7), .O(gate166inter9));
  nand2 gate2699(.a(s_307), .b(gate166inter3), .O(gate166inter10));
  nor2  gate2700(.a(gate166inter10), .b(gate166inter9), .O(gate166inter11));
  nor2  gate2701(.a(gate166inter11), .b(gate166inter6), .O(gate166inter12));
  nand2 gate2702(.a(gate166inter12), .b(gate166inter1), .O(G583));
nand2 gate167( .a(G468), .b(G543), .O(G584) );
nand2 gate168( .a(G471), .b(G543), .O(G585) );
nand2 gate169( .a(G474), .b(G546), .O(G586) );
nand2 gate170( .a(G477), .b(G546), .O(G587) );

  xor2  gate1737(.a(G549), .b(G480), .O(gate171inter0));
  nand2 gate1738(.a(gate171inter0), .b(s_170), .O(gate171inter1));
  and2  gate1739(.a(G549), .b(G480), .O(gate171inter2));
  inv1  gate1740(.a(s_170), .O(gate171inter3));
  inv1  gate1741(.a(s_171), .O(gate171inter4));
  nand2 gate1742(.a(gate171inter4), .b(gate171inter3), .O(gate171inter5));
  nor2  gate1743(.a(gate171inter5), .b(gate171inter2), .O(gate171inter6));
  inv1  gate1744(.a(G480), .O(gate171inter7));
  inv1  gate1745(.a(G549), .O(gate171inter8));
  nand2 gate1746(.a(gate171inter8), .b(gate171inter7), .O(gate171inter9));
  nand2 gate1747(.a(s_171), .b(gate171inter3), .O(gate171inter10));
  nor2  gate1748(.a(gate171inter10), .b(gate171inter9), .O(gate171inter11));
  nor2  gate1749(.a(gate171inter11), .b(gate171inter6), .O(gate171inter12));
  nand2 gate1750(.a(gate171inter12), .b(gate171inter1), .O(G588));
nand2 gate172( .a(G483), .b(G549), .O(G589) );

  xor2  gate1569(.a(G552), .b(G486), .O(gate173inter0));
  nand2 gate1570(.a(gate173inter0), .b(s_146), .O(gate173inter1));
  and2  gate1571(.a(G552), .b(G486), .O(gate173inter2));
  inv1  gate1572(.a(s_146), .O(gate173inter3));
  inv1  gate1573(.a(s_147), .O(gate173inter4));
  nand2 gate1574(.a(gate173inter4), .b(gate173inter3), .O(gate173inter5));
  nor2  gate1575(.a(gate173inter5), .b(gate173inter2), .O(gate173inter6));
  inv1  gate1576(.a(G486), .O(gate173inter7));
  inv1  gate1577(.a(G552), .O(gate173inter8));
  nand2 gate1578(.a(gate173inter8), .b(gate173inter7), .O(gate173inter9));
  nand2 gate1579(.a(s_147), .b(gate173inter3), .O(gate173inter10));
  nor2  gate1580(.a(gate173inter10), .b(gate173inter9), .O(gate173inter11));
  nor2  gate1581(.a(gate173inter11), .b(gate173inter6), .O(gate173inter12));
  nand2 gate1582(.a(gate173inter12), .b(gate173inter1), .O(G590));

  xor2  gate799(.a(G552), .b(G489), .O(gate174inter0));
  nand2 gate800(.a(gate174inter0), .b(s_36), .O(gate174inter1));
  and2  gate801(.a(G552), .b(G489), .O(gate174inter2));
  inv1  gate802(.a(s_36), .O(gate174inter3));
  inv1  gate803(.a(s_37), .O(gate174inter4));
  nand2 gate804(.a(gate174inter4), .b(gate174inter3), .O(gate174inter5));
  nor2  gate805(.a(gate174inter5), .b(gate174inter2), .O(gate174inter6));
  inv1  gate806(.a(G489), .O(gate174inter7));
  inv1  gate807(.a(G552), .O(gate174inter8));
  nand2 gate808(.a(gate174inter8), .b(gate174inter7), .O(gate174inter9));
  nand2 gate809(.a(s_37), .b(gate174inter3), .O(gate174inter10));
  nor2  gate810(.a(gate174inter10), .b(gate174inter9), .O(gate174inter11));
  nor2  gate811(.a(gate174inter11), .b(gate174inter6), .O(gate174inter12));
  nand2 gate812(.a(gate174inter12), .b(gate174inter1), .O(G591));
nand2 gate175( .a(G492), .b(G555), .O(G592) );
nand2 gate176( .a(G495), .b(G555), .O(G593) );
nand2 gate177( .a(G498), .b(G558), .O(G594) );
nand2 gate178( .a(G501), .b(G558), .O(G595) );
nand2 gate179( .a(G504), .b(G561), .O(G596) );

  xor2  gate995(.a(G561), .b(G507), .O(gate180inter0));
  nand2 gate996(.a(gate180inter0), .b(s_64), .O(gate180inter1));
  and2  gate997(.a(G561), .b(G507), .O(gate180inter2));
  inv1  gate998(.a(s_64), .O(gate180inter3));
  inv1  gate999(.a(s_65), .O(gate180inter4));
  nand2 gate1000(.a(gate180inter4), .b(gate180inter3), .O(gate180inter5));
  nor2  gate1001(.a(gate180inter5), .b(gate180inter2), .O(gate180inter6));
  inv1  gate1002(.a(G507), .O(gate180inter7));
  inv1  gate1003(.a(G561), .O(gate180inter8));
  nand2 gate1004(.a(gate180inter8), .b(gate180inter7), .O(gate180inter9));
  nand2 gate1005(.a(s_65), .b(gate180inter3), .O(gate180inter10));
  nor2  gate1006(.a(gate180inter10), .b(gate180inter9), .O(gate180inter11));
  nor2  gate1007(.a(gate180inter11), .b(gate180inter6), .O(gate180inter12));
  nand2 gate1008(.a(gate180inter12), .b(gate180inter1), .O(G597));
nand2 gate181( .a(G510), .b(G564), .O(G598) );

  xor2  gate1457(.a(G564), .b(G513), .O(gate182inter0));
  nand2 gate1458(.a(gate182inter0), .b(s_130), .O(gate182inter1));
  and2  gate1459(.a(G564), .b(G513), .O(gate182inter2));
  inv1  gate1460(.a(s_130), .O(gate182inter3));
  inv1  gate1461(.a(s_131), .O(gate182inter4));
  nand2 gate1462(.a(gate182inter4), .b(gate182inter3), .O(gate182inter5));
  nor2  gate1463(.a(gate182inter5), .b(gate182inter2), .O(gate182inter6));
  inv1  gate1464(.a(G513), .O(gate182inter7));
  inv1  gate1465(.a(G564), .O(gate182inter8));
  nand2 gate1466(.a(gate182inter8), .b(gate182inter7), .O(gate182inter9));
  nand2 gate1467(.a(s_131), .b(gate182inter3), .O(gate182inter10));
  nor2  gate1468(.a(gate182inter10), .b(gate182inter9), .O(gate182inter11));
  nor2  gate1469(.a(gate182inter11), .b(gate182inter6), .O(gate182inter12));
  nand2 gate1470(.a(gate182inter12), .b(gate182inter1), .O(G599));
nand2 gate183( .a(G516), .b(G567), .O(G600) );
nand2 gate184( .a(G519), .b(G567), .O(G601) );
nand2 gate185( .a(G570), .b(G571), .O(G602) );
nand2 gate186( .a(G572), .b(G573), .O(G607) );
nand2 gate187( .a(G574), .b(G575), .O(G612) );
nand2 gate188( .a(G576), .b(G577), .O(G617) );
nand2 gate189( .a(G578), .b(G579), .O(G622) );
nand2 gate190( .a(G580), .b(G581), .O(G627) );

  xor2  gate2199(.a(G583), .b(G582), .O(gate191inter0));
  nand2 gate2200(.a(gate191inter0), .b(s_236), .O(gate191inter1));
  and2  gate2201(.a(G583), .b(G582), .O(gate191inter2));
  inv1  gate2202(.a(s_236), .O(gate191inter3));
  inv1  gate2203(.a(s_237), .O(gate191inter4));
  nand2 gate2204(.a(gate191inter4), .b(gate191inter3), .O(gate191inter5));
  nor2  gate2205(.a(gate191inter5), .b(gate191inter2), .O(gate191inter6));
  inv1  gate2206(.a(G582), .O(gate191inter7));
  inv1  gate2207(.a(G583), .O(gate191inter8));
  nand2 gate2208(.a(gate191inter8), .b(gate191inter7), .O(gate191inter9));
  nand2 gate2209(.a(s_237), .b(gate191inter3), .O(gate191inter10));
  nor2  gate2210(.a(gate191inter10), .b(gate191inter9), .O(gate191inter11));
  nor2  gate2211(.a(gate191inter11), .b(gate191inter6), .O(gate191inter12));
  nand2 gate2212(.a(gate191inter12), .b(gate191inter1), .O(G632));
nand2 gate192( .a(G584), .b(G585), .O(G637) );
nand2 gate193( .a(G586), .b(G587), .O(G642) );

  xor2  gate1779(.a(G589), .b(G588), .O(gate194inter0));
  nand2 gate1780(.a(gate194inter0), .b(s_176), .O(gate194inter1));
  and2  gate1781(.a(G589), .b(G588), .O(gate194inter2));
  inv1  gate1782(.a(s_176), .O(gate194inter3));
  inv1  gate1783(.a(s_177), .O(gate194inter4));
  nand2 gate1784(.a(gate194inter4), .b(gate194inter3), .O(gate194inter5));
  nor2  gate1785(.a(gate194inter5), .b(gate194inter2), .O(gate194inter6));
  inv1  gate1786(.a(G588), .O(gate194inter7));
  inv1  gate1787(.a(G589), .O(gate194inter8));
  nand2 gate1788(.a(gate194inter8), .b(gate194inter7), .O(gate194inter9));
  nand2 gate1789(.a(s_177), .b(gate194inter3), .O(gate194inter10));
  nor2  gate1790(.a(gate194inter10), .b(gate194inter9), .O(gate194inter11));
  nor2  gate1791(.a(gate194inter11), .b(gate194inter6), .O(gate194inter12));
  nand2 gate1792(.a(gate194inter12), .b(gate194inter1), .O(G645));
nand2 gate195( .a(G590), .b(G591), .O(G648) );

  xor2  gate645(.a(G593), .b(G592), .O(gate196inter0));
  nand2 gate646(.a(gate196inter0), .b(s_14), .O(gate196inter1));
  and2  gate647(.a(G593), .b(G592), .O(gate196inter2));
  inv1  gate648(.a(s_14), .O(gate196inter3));
  inv1  gate649(.a(s_15), .O(gate196inter4));
  nand2 gate650(.a(gate196inter4), .b(gate196inter3), .O(gate196inter5));
  nor2  gate651(.a(gate196inter5), .b(gate196inter2), .O(gate196inter6));
  inv1  gate652(.a(G592), .O(gate196inter7));
  inv1  gate653(.a(G593), .O(gate196inter8));
  nand2 gate654(.a(gate196inter8), .b(gate196inter7), .O(gate196inter9));
  nand2 gate655(.a(s_15), .b(gate196inter3), .O(gate196inter10));
  nor2  gate656(.a(gate196inter10), .b(gate196inter9), .O(gate196inter11));
  nor2  gate657(.a(gate196inter11), .b(gate196inter6), .O(gate196inter12));
  nand2 gate658(.a(gate196inter12), .b(gate196inter1), .O(G651));

  xor2  gate939(.a(G595), .b(G594), .O(gate197inter0));
  nand2 gate940(.a(gate197inter0), .b(s_56), .O(gate197inter1));
  and2  gate941(.a(G595), .b(G594), .O(gate197inter2));
  inv1  gate942(.a(s_56), .O(gate197inter3));
  inv1  gate943(.a(s_57), .O(gate197inter4));
  nand2 gate944(.a(gate197inter4), .b(gate197inter3), .O(gate197inter5));
  nor2  gate945(.a(gate197inter5), .b(gate197inter2), .O(gate197inter6));
  inv1  gate946(.a(G594), .O(gate197inter7));
  inv1  gate947(.a(G595), .O(gate197inter8));
  nand2 gate948(.a(gate197inter8), .b(gate197inter7), .O(gate197inter9));
  nand2 gate949(.a(s_57), .b(gate197inter3), .O(gate197inter10));
  nor2  gate950(.a(gate197inter10), .b(gate197inter9), .O(gate197inter11));
  nor2  gate951(.a(gate197inter11), .b(gate197inter6), .O(gate197inter12));
  nand2 gate952(.a(gate197inter12), .b(gate197inter1), .O(G654));
nand2 gate198( .a(G596), .b(G597), .O(G657) );
nand2 gate199( .a(G598), .b(G599), .O(G660) );
nand2 gate200( .a(G600), .b(G601), .O(G663) );
nand2 gate201( .a(G602), .b(G607), .O(G666) );
nand2 gate202( .a(G612), .b(G617), .O(G669) );

  xor2  gate2171(.a(G612), .b(G602), .O(gate203inter0));
  nand2 gate2172(.a(gate203inter0), .b(s_232), .O(gate203inter1));
  and2  gate2173(.a(G612), .b(G602), .O(gate203inter2));
  inv1  gate2174(.a(s_232), .O(gate203inter3));
  inv1  gate2175(.a(s_233), .O(gate203inter4));
  nand2 gate2176(.a(gate203inter4), .b(gate203inter3), .O(gate203inter5));
  nor2  gate2177(.a(gate203inter5), .b(gate203inter2), .O(gate203inter6));
  inv1  gate2178(.a(G602), .O(gate203inter7));
  inv1  gate2179(.a(G612), .O(gate203inter8));
  nand2 gate2180(.a(gate203inter8), .b(gate203inter7), .O(gate203inter9));
  nand2 gate2181(.a(s_233), .b(gate203inter3), .O(gate203inter10));
  nor2  gate2182(.a(gate203inter10), .b(gate203inter9), .O(gate203inter11));
  nor2  gate2183(.a(gate203inter11), .b(gate203inter6), .O(gate203inter12));
  nand2 gate2184(.a(gate203inter12), .b(gate203inter1), .O(G672));

  xor2  gate1331(.a(G617), .b(G607), .O(gate204inter0));
  nand2 gate1332(.a(gate204inter0), .b(s_112), .O(gate204inter1));
  and2  gate1333(.a(G617), .b(G607), .O(gate204inter2));
  inv1  gate1334(.a(s_112), .O(gate204inter3));
  inv1  gate1335(.a(s_113), .O(gate204inter4));
  nand2 gate1336(.a(gate204inter4), .b(gate204inter3), .O(gate204inter5));
  nor2  gate1337(.a(gate204inter5), .b(gate204inter2), .O(gate204inter6));
  inv1  gate1338(.a(G607), .O(gate204inter7));
  inv1  gate1339(.a(G617), .O(gate204inter8));
  nand2 gate1340(.a(gate204inter8), .b(gate204inter7), .O(gate204inter9));
  nand2 gate1341(.a(s_113), .b(gate204inter3), .O(gate204inter10));
  nor2  gate1342(.a(gate204inter10), .b(gate204inter9), .O(gate204inter11));
  nor2  gate1343(.a(gate204inter11), .b(gate204inter6), .O(gate204inter12));
  nand2 gate1344(.a(gate204inter12), .b(gate204inter1), .O(G675));

  xor2  gate1625(.a(G627), .b(G622), .O(gate205inter0));
  nand2 gate1626(.a(gate205inter0), .b(s_154), .O(gate205inter1));
  and2  gate1627(.a(G627), .b(G622), .O(gate205inter2));
  inv1  gate1628(.a(s_154), .O(gate205inter3));
  inv1  gate1629(.a(s_155), .O(gate205inter4));
  nand2 gate1630(.a(gate205inter4), .b(gate205inter3), .O(gate205inter5));
  nor2  gate1631(.a(gate205inter5), .b(gate205inter2), .O(gate205inter6));
  inv1  gate1632(.a(G622), .O(gate205inter7));
  inv1  gate1633(.a(G627), .O(gate205inter8));
  nand2 gate1634(.a(gate205inter8), .b(gate205inter7), .O(gate205inter9));
  nand2 gate1635(.a(s_155), .b(gate205inter3), .O(gate205inter10));
  nor2  gate1636(.a(gate205inter10), .b(gate205inter9), .O(gate205inter11));
  nor2  gate1637(.a(gate205inter11), .b(gate205inter6), .O(gate205inter12));
  nand2 gate1638(.a(gate205inter12), .b(gate205inter1), .O(G678));
nand2 gate206( .a(G632), .b(G637), .O(G681) );

  xor2  gate2451(.a(G632), .b(G622), .O(gate207inter0));
  nand2 gate2452(.a(gate207inter0), .b(s_272), .O(gate207inter1));
  and2  gate2453(.a(G632), .b(G622), .O(gate207inter2));
  inv1  gate2454(.a(s_272), .O(gate207inter3));
  inv1  gate2455(.a(s_273), .O(gate207inter4));
  nand2 gate2456(.a(gate207inter4), .b(gate207inter3), .O(gate207inter5));
  nor2  gate2457(.a(gate207inter5), .b(gate207inter2), .O(gate207inter6));
  inv1  gate2458(.a(G622), .O(gate207inter7));
  inv1  gate2459(.a(G632), .O(gate207inter8));
  nand2 gate2460(.a(gate207inter8), .b(gate207inter7), .O(gate207inter9));
  nand2 gate2461(.a(s_273), .b(gate207inter3), .O(gate207inter10));
  nor2  gate2462(.a(gate207inter10), .b(gate207inter9), .O(gate207inter11));
  nor2  gate2463(.a(gate207inter11), .b(gate207inter6), .O(gate207inter12));
  nand2 gate2464(.a(gate207inter12), .b(gate207inter1), .O(G684));
nand2 gate208( .a(G627), .b(G637), .O(G687) );

  xor2  gate841(.a(G666), .b(G602), .O(gate209inter0));
  nand2 gate842(.a(gate209inter0), .b(s_42), .O(gate209inter1));
  and2  gate843(.a(G666), .b(G602), .O(gate209inter2));
  inv1  gate844(.a(s_42), .O(gate209inter3));
  inv1  gate845(.a(s_43), .O(gate209inter4));
  nand2 gate846(.a(gate209inter4), .b(gate209inter3), .O(gate209inter5));
  nor2  gate847(.a(gate209inter5), .b(gate209inter2), .O(gate209inter6));
  inv1  gate848(.a(G602), .O(gate209inter7));
  inv1  gate849(.a(G666), .O(gate209inter8));
  nand2 gate850(.a(gate209inter8), .b(gate209inter7), .O(gate209inter9));
  nand2 gate851(.a(s_43), .b(gate209inter3), .O(gate209inter10));
  nor2  gate852(.a(gate209inter10), .b(gate209inter9), .O(gate209inter11));
  nor2  gate853(.a(gate209inter11), .b(gate209inter6), .O(gate209inter12));
  nand2 gate854(.a(gate209inter12), .b(gate209inter1), .O(G690));

  xor2  gate561(.a(G666), .b(G607), .O(gate210inter0));
  nand2 gate562(.a(gate210inter0), .b(s_2), .O(gate210inter1));
  and2  gate563(.a(G666), .b(G607), .O(gate210inter2));
  inv1  gate564(.a(s_2), .O(gate210inter3));
  inv1  gate565(.a(s_3), .O(gate210inter4));
  nand2 gate566(.a(gate210inter4), .b(gate210inter3), .O(gate210inter5));
  nor2  gate567(.a(gate210inter5), .b(gate210inter2), .O(gate210inter6));
  inv1  gate568(.a(G607), .O(gate210inter7));
  inv1  gate569(.a(G666), .O(gate210inter8));
  nand2 gate570(.a(gate210inter8), .b(gate210inter7), .O(gate210inter9));
  nand2 gate571(.a(s_3), .b(gate210inter3), .O(gate210inter10));
  nor2  gate572(.a(gate210inter10), .b(gate210inter9), .O(gate210inter11));
  nor2  gate573(.a(gate210inter11), .b(gate210inter6), .O(gate210inter12));
  nand2 gate574(.a(gate210inter12), .b(gate210inter1), .O(G691));

  xor2  gate2829(.a(G669), .b(G612), .O(gate211inter0));
  nand2 gate2830(.a(gate211inter0), .b(s_326), .O(gate211inter1));
  and2  gate2831(.a(G669), .b(G612), .O(gate211inter2));
  inv1  gate2832(.a(s_326), .O(gate211inter3));
  inv1  gate2833(.a(s_327), .O(gate211inter4));
  nand2 gate2834(.a(gate211inter4), .b(gate211inter3), .O(gate211inter5));
  nor2  gate2835(.a(gate211inter5), .b(gate211inter2), .O(gate211inter6));
  inv1  gate2836(.a(G612), .O(gate211inter7));
  inv1  gate2837(.a(G669), .O(gate211inter8));
  nand2 gate2838(.a(gate211inter8), .b(gate211inter7), .O(gate211inter9));
  nand2 gate2839(.a(s_327), .b(gate211inter3), .O(gate211inter10));
  nor2  gate2840(.a(gate211inter10), .b(gate211inter9), .O(gate211inter11));
  nor2  gate2841(.a(gate211inter11), .b(gate211inter6), .O(gate211inter12));
  nand2 gate2842(.a(gate211inter12), .b(gate211inter1), .O(G692));

  xor2  gate2927(.a(G669), .b(G617), .O(gate212inter0));
  nand2 gate2928(.a(gate212inter0), .b(s_340), .O(gate212inter1));
  and2  gate2929(.a(G669), .b(G617), .O(gate212inter2));
  inv1  gate2930(.a(s_340), .O(gate212inter3));
  inv1  gate2931(.a(s_341), .O(gate212inter4));
  nand2 gate2932(.a(gate212inter4), .b(gate212inter3), .O(gate212inter5));
  nor2  gate2933(.a(gate212inter5), .b(gate212inter2), .O(gate212inter6));
  inv1  gate2934(.a(G617), .O(gate212inter7));
  inv1  gate2935(.a(G669), .O(gate212inter8));
  nand2 gate2936(.a(gate212inter8), .b(gate212inter7), .O(gate212inter9));
  nand2 gate2937(.a(s_341), .b(gate212inter3), .O(gate212inter10));
  nor2  gate2938(.a(gate212inter10), .b(gate212inter9), .O(gate212inter11));
  nor2  gate2939(.a(gate212inter11), .b(gate212inter6), .O(gate212inter12));
  nand2 gate2940(.a(gate212inter12), .b(gate212inter1), .O(G693));

  xor2  gate2241(.a(G672), .b(G602), .O(gate213inter0));
  nand2 gate2242(.a(gate213inter0), .b(s_242), .O(gate213inter1));
  and2  gate2243(.a(G672), .b(G602), .O(gate213inter2));
  inv1  gate2244(.a(s_242), .O(gate213inter3));
  inv1  gate2245(.a(s_243), .O(gate213inter4));
  nand2 gate2246(.a(gate213inter4), .b(gate213inter3), .O(gate213inter5));
  nor2  gate2247(.a(gate213inter5), .b(gate213inter2), .O(gate213inter6));
  inv1  gate2248(.a(G602), .O(gate213inter7));
  inv1  gate2249(.a(G672), .O(gate213inter8));
  nand2 gate2250(.a(gate213inter8), .b(gate213inter7), .O(gate213inter9));
  nand2 gate2251(.a(s_243), .b(gate213inter3), .O(gate213inter10));
  nor2  gate2252(.a(gate213inter10), .b(gate213inter9), .O(gate213inter11));
  nor2  gate2253(.a(gate213inter11), .b(gate213inter6), .O(gate213inter12));
  nand2 gate2254(.a(gate213inter12), .b(gate213inter1), .O(G694));

  xor2  gate1107(.a(G672), .b(G612), .O(gate214inter0));
  nand2 gate1108(.a(gate214inter0), .b(s_80), .O(gate214inter1));
  and2  gate1109(.a(G672), .b(G612), .O(gate214inter2));
  inv1  gate1110(.a(s_80), .O(gate214inter3));
  inv1  gate1111(.a(s_81), .O(gate214inter4));
  nand2 gate1112(.a(gate214inter4), .b(gate214inter3), .O(gate214inter5));
  nor2  gate1113(.a(gate214inter5), .b(gate214inter2), .O(gate214inter6));
  inv1  gate1114(.a(G612), .O(gate214inter7));
  inv1  gate1115(.a(G672), .O(gate214inter8));
  nand2 gate1116(.a(gate214inter8), .b(gate214inter7), .O(gate214inter9));
  nand2 gate1117(.a(s_81), .b(gate214inter3), .O(gate214inter10));
  nor2  gate1118(.a(gate214inter10), .b(gate214inter9), .O(gate214inter11));
  nor2  gate1119(.a(gate214inter11), .b(gate214inter6), .O(gate214inter12));
  nand2 gate1120(.a(gate214inter12), .b(gate214inter1), .O(G695));
nand2 gate215( .a(G607), .b(G675), .O(G696) );
nand2 gate216( .a(G617), .b(G675), .O(G697) );
nand2 gate217( .a(G622), .b(G678), .O(G698) );
nand2 gate218( .a(G627), .b(G678), .O(G699) );
nand2 gate219( .a(G632), .b(G681), .O(G700) );

  xor2  gate1387(.a(G681), .b(G637), .O(gate220inter0));
  nand2 gate1388(.a(gate220inter0), .b(s_120), .O(gate220inter1));
  and2  gate1389(.a(G681), .b(G637), .O(gate220inter2));
  inv1  gate1390(.a(s_120), .O(gate220inter3));
  inv1  gate1391(.a(s_121), .O(gate220inter4));
  nand2 gate1392(.a(gate220inter4), .b(gate220inter3), .O(gate220inter5));
  nor2  gate1393(.a(gate220inter5), .b(gate220inter2), .O(gate220inter6));
  inv1  gate1394(.a(G637), .O(gate220inter7));
  inv1  gate1395(.a(G681), .O(gate220inter8));
  nand2 gate1396(.a(gate220inter8), .b(gate220inter7), .O(gate220inter9));
  nand2 gate1397(.a(s_121), .b(gate220inter3), .O(gate220inter10));
  nor2  gate1398(.a(gate220inter10), .b(gate220inter9), .O(gate220inter11));
  nor2  gate1399(.a(gate220inter11), .b(gate220inter6), .O(gate220inter12));
  nand2 gate1400(.a(gate220inter12), .b(gate220inter1), .O(G701));

  xor2  gate1261(.a(G684), .b(G622), .O(gate221inter0));
  nand2 gate1262(.a(gate221inter0), .b(s_102), .O(gate221inter1));
  and2  gate1263(.a(G684), .b(G622), .O(gate221inter2));
  inv1  gate1264(.a(s_102), .O(gate221inter3));
  inv1  gate1265(.a(s_103), .O(gate221inter4));
  nand2 gate1266(.a(gate221inter4), .b(gate221inter3), .O(gate221inter5));
  nor2  gate1267(.a(gate221inter5), .b(gate221inter2), .O(gate221inter6));
  inv1  gate1268(.a(G622), .O(gate221inter7));
  inv1  gate1269(.a(G684), .O(gate221inter8));
  nand2 gate1270(.a(gate221inter8), .b(gate221inter7), .O(gate221inter9));
  nand2 gate1271(.a(s_103), .b(gate221inter3), .O(gate221inter10));
  nor2  gate1272(.a(gate221inter10), .b(gate221inter9), .O(gate221inter11));
  nor2  gate1273(.a(gate221inter11), .b(gate221inter6), .O(gate221inter12));
  nand2 gate1274(.a(gate221inter12), .b(gate221inter1), .O(G702));
nand2 gate222( .a(G632), .b(G684), .O(G703) );

  xor2  gate2759(.a(G687), .b(G627), .O(gate223inter0));
  nand2 gate2760(.a(gate223inter0), .b(s_316), .O(gate223inter1));
  and2  gate2761(.a(G687), .b(G627), .O(gate223inter2));
  inv1  gate2762(.a(s_316), .O(gate223inter3));
  inv1  gate2763(.a(s_317), .O(gate223inter4));
  nand2 gate2764(.a(gate223inter4), .b(gate223inter3), .O(gate223inter5));
  nor2  gate2765(.a(gate223inter5), .b(gate223inter2), .O(gate223inter6));
  inv1  gate2766(.a(G627), .O(gate223inter7));
  inv1  gate2767(.a(G687), .O(gate223inter8));
  nand2 gate2768(.a(gate223inter8), .b(gate223inter7), .O(gate223inter9));
  nand2 gate2769(.a(s_317), .b(gate223inter3), .O(gate223inter10));
  nor2  gate2770(.a(gate223inter10), .b(gate223inter9), .O(gate223inter11));
  nor2  gate2771(.a(gate223inter11), .b(gate223inter6), .O(gate223inter12));
  nand2 gate2772(.a(gate223inter12), .b(gate223inter1), .O(G704));

  xor2  gate1065(.a(G687), .b(G637), .O(gate224inter0));
  nand2 gate1066(.a(gate224inter0), .b(s_74), .O(gate224inter1));
  and2  gate1067(.a(G687), .b(G637), .O(gate224inter2));
  inv1  gate1068(.a(s_74), .O(gate224inter3));
  inv1  gate1069(.a(s_75), .O(gate224inter4));
  nand2 gate1070(.a(gate224inter4), .b(gate224inter3), .O(gate224inter5));
  nor2  gate1071(.a(gate224inter5), .b(gate224inter2), .O(gate224inter6));
  inv1  gate1072(.a(G637), .O(gate224inter7));
  inv1  gate1073(.a(G687), .O(gate224inter8));
  nand2 gate1074(.a(gate224inter8), .b(gate224inter7), .O(gate224inter9));
  nand2 gate1075(.a(s_75), .b(gate224inter3), .O(gate224inter10));
  nor2  gate1076(.a(gate224inter10), .b(gate224inter9), .O(gate224inter11));
  nor2  gate1077(.a(gate224inter11), .b(gate224inter6), .O(gate224inter12));
  nand2 gate1078(.a(gate224inter12), .b(gate224inter1), .O(G705));
nand2 gate225( .a(G690), .b(G691), .O(G706) );
nand2 gate226( .a(G692), .b(G693), .O(G709) );
nand2 gate227( .a(G694), .b(G695), .O(G712) );
nand2 gate228( .a(G696), .b(G697), .O(G715) );
nand2 gate229( .a(G698), .b(G699), .O(G718) );
nand2 gate230( .a(G700), .b(G701), .O(G721) );

  xor2  gate617(.a(G703), .b(G702), .O(gate231inter0));
  nand2 gate618(.a(gate231inter0), .b(s_10), .O(gate231inter1));
  and2  gate619(.a(G703), .b(G702), .O(gate231inter2));
  inv1  gate620(.a(s_10), .O(gate231inter3));
  inv1  gate621(.a(s_11), .O(gate231inter4));
  nand2 gate622(.a(gate231inter4), .b(gate231inter3), .O(gate231inter5));
  nor2  gate623(.a(gate231inter5), .b(gate231inter2), .O(gate231inter6));
  inv1  gate624(.a(G702), .O(gate231inter7));
  inv1  gate625(.a(G703), .O(gate231inter8));
  nand2 gate626(.a(gate231inter8), .b(gate231inter7), .O(gate231inter9));
  nand2 gate627(.a(s_11), .b(gate231inter3), .O(gate231inter10));
  nor2  gate628(.a(gate231inter10), .b(gate231inter9), .O(gate231inter11));
  nor2  gate629(.a(gate231inter11), .b(gate231inter6), .O(gate231inter12));
  nand2 gate630(.a(gate231inter12), .b(gate231inter1), .O(G724));
nand2 gate232( .a(G704), .b(G705), .O(G727) );

  xor2  gate1765(.a(G718), .b(G242), .O(gate233inter0));
  nand2 gate1766(.a(gate233inter0), .b(s_174), .O(gate233inter1));
  and2  gate1767(.a(G718), .b(G242), .O(gate233inter2));
  inv1  gate1768(.a(s_174), .O(gate233inter3));
  inv1  gate1769(.a(s_175), .O(gate233inter4));
  nand2 gate1770(.a(gate233inter4), .b(gate233inter3), .O(gate233inter5));
  nor2  gate1771(.a(gate233inter5), .b(gate233inter2), .O(gate233inter6));
  inv1  gate1772(.a(G242), .O(gate233inter7));
  inv1  gate1773(.a(G718), .O(gate233inter8));
  nand2 gate1774(.a(gate233inter8), .b(gate233inter7), .O(gate233inter9));
  nand2 gate1775(.a(s_175), .b(gate233inter3), .O(gate233inter10));
  nor2  gate1776(.a(gate233inter10), .b(gate233inter9), .O(gate233inter11));
  nor2  gate1777(.a(gate233inter11), .b(gate233inter6), .O(gate233inter12));
  nand2 gate1778(.a(gate233inter12), .b(gate233inter1), .O(G730));
nand2 gate234( .a(G245), .b(G721), .O(G733) );

  xor2  gate1163(.a(G724), .b(G248), .O(gate235inter0));
  nand2 gate1164(.a(gate235inter0), .b(s_88), .O(gate235inter1));
  and2  gate1165(.a(G724), .b(G248), .O(gate235inter2));
  inv1  gate1166(.a(s_88), .O(gate235inter3));
  inv1  gate1167(.a(s_89), .O(gate235inter4));
  nand2 gate1168(.a(gate235inter4), .b(gate235inter3), .O(gate235inter5));
  nor2  gate1169(.a(gate235inter5), .b(gate235inter2), .O(gate235inter6));
  inv1  gate1170(.a(G248), .O(gate235inter7));
  inv1  gate1171(.a(G724), .O(gate235inter8));
  nand2 gate1172(.a(gate235inter8), .b(gate235inter7), .O(gate235inter9));
  nand2 gate1173(.a(s_89), .b(gate235inter3), .O(gate235inter10));
  nor2  gate1174(.a(gate235inter10), .b(gate235inter9), .O(gate235inter11));
  nor2  gate1175(.a(gate235inter11), .b(gate235inter6), .O(gate235inter12));
  nand2 gate1176(.a(gate235inter12), .b(gate235inter1), .O(G736));

  xor2  gate2605(.a(G727), .b(G251), .O(gate236inter0));
  nand2 gate2606(.a(gate236inter0), .b(s_294), .O(gate236inter1));
  and2  gate2607(.a(G727), .b(G251), .O(gate236inter2));
  inv1  gate2608(.a(s_294), .O(gate236inter3));
  inv1  gate2609(.a(s_295), .O(gate236inter4));
  nand2 gate2610(.a(gate236inter4), .b(gate236inter3), .O(gate236inter5));
  nor2  gate2611(.a(gate236inter5), .b(gate236inter2), .O(gate236inter6));
  inv1  gate2612(.a(G251), .O(gate236inter7));
  inv1  gate2613(.a(G727), .O(gate236inter8));
  nand2 gate2614(.a(gate236inter8), .b(gate236inter7), .O(gate236inter9));
  nand2 gate2615(.a(s_295), .b(gate236inter3), .O(gate236inter10));
  nor2  gate2616(.a(gate236inter10), .b(gate236inter9), .O(gate236inter11));
  nor2  gate2617(.a(gate236inter11), .b(gate236inter6), .O(gate236inter12));
  nand2 gate2618(.a(gate236inter12), .b(gate236inter1), .O(G739));
nand2 gate237( .a(G254), .b(G706), .O(G742) );
nand2 gate238( .a(G257), .b(G709), .O(G745) );

  xor2  gate2395(.a(G712), .b(G260), .O(gate239inter0));
  nand2 gate2396(.a(gate239inter0), .b(s_264), .O(gate239inter1));
  and2  gate2397(.a(G712), .b(G260), .O(gate239inter2));
  inv1  gate2398(.a(s_264), .O(gate239inter3));
  inv1  gate2399(.a(s_265), .O(gate239inter4));
  nand2 gate2400(.a(gate239inter4), .b(gate239inter3), .O(gate239inter5));
  nor2  gate2401(.a(gate239inter5), .b(gate239inter2), .O(gate239inter6));
  inv1  gate2402(.a(G260), .O(gate239inter7));
  inv1  gate2403(.a(G712), .O(gate239inter8));
  nand2 gate2404(.a(gate239inter8), .b(gate239inter7), .O(gate239inter9));
  nand2 gate2405(.a(s_265), .b(gate239inter3), .O(gate239inter10));
  nor2  gate2406(.a(gate239inter10), .b(gate239inter9), .O(gate239inter11));
  nor2  gate2407(.a(gate239inter11), .b(gate239inter6), .O(gate239inter12));
  nand2 gate2408(.a(gate239inter12), .b(gate239inter1), .O(G748));

  xor2  gate1079(.a(G715), .b(G263), .O(gate240inter0));
  nand2 gate1080(.a(gate240inter0), .b(s_76), .O(gate240inter1));
  and2  gate1081(.a(G715), .b(G263), .O(gate240inter2));
  inv1  gate1082(.a(s_76), .O(gate240inter3));
  inv1  gate1083(.a(s_77), .O(gate240inter4));
  nand2 gate1084(.a(gate240inter4), .b(gate240inter3), .O(gate240inter5));
  nor2  gate1085(.a(gate240inter5), .b(gate240inter2), .O(gate240inter6));
  inv1  gate1086(.a(G263), .O(gate240inter7));
  inv1  gate1087(.a(G715), .O(gate240inter8));
  nand2 gate1088(.a(gate240inter8), .b(gate240inter7), .O(gate240inter9));
  nand2 gate1089(.a(s_77), .b(gate240inter3), .O(gate240inter10));
  nor2  gate1090(.a(gate240inter10), .b(gate240inter9), .O(gate240inter11));
  nor2  gate1091(.a(gate240inter11), .b(gate240inter6), .O(gate240inter12));
  nand2 gate1092(.a(gate240inter12), .b(gate240inter1), .O(G751));
nand2 gate241( .a(G242), .b(G730), .O(G754) );
nand2 gate242( .a(G718), .b(G730), .O(G755) );
nand2 gate243( .a(G245), .b(G733), .O(G756) );
nand2 gate244( .a(G721), .b(G733), .O(G757) );

  xor2  gate2717(.a(G736), .b(G248), .O(gate245inter0));
  nand2 gate2718(.a(gate245inter0), .b(s_310), .O(gate245inter1));
  and2  gate2719(.a(G736), .b(G248), .O(gate245inter2));
  inv1  gate2720(.a(s_310), .O(gate245inter3));
  inv1  gate2721(.a(s_311), .O(gate245inter4));
  nand2 gate2722(.a(gate245inter4), .b(gate245inter3), .O(gate245inter5));
  nor2  gate2723(.a(gate245inter5), .b(gate245inter2), .O(gate245inter6));
  inv1  gate2724(.a(G248), .O(gate245inter7));
  inv1  gate2725(.a(G736), .O(gate245inter8));
  nand2 gate2726(.a(gate245inter8), .b(gate245inter7), .O(gate245inter9));
  nand2 gate2727(.a(s_311), .b(gate245inter3), .O(gate245inter10));
  nor2  gate2728(.a(gate245inter10), .b(gate245inter9), .O(gate245inter11));
  nor2  gate2729(.a(gate245inter11), .b(gate245inter6), .O(gate245inter12));
  nand2 gate2730(.a(gate245inter12), .b(gate245inter1), .O(G758));
nand2 gate246( .a(G724), .b(G736), .O(G759) );
nand2 gate247( .a(G251), .b(G739), .O(G760) );

  xor2  gate1037(.a(G739), .b(G727), .O(gate248inter0));
  nand2 gate1038(.a(gate248inter0), .b(s_70), .O(gate248inter1));
  and2  gate1039(.a(G739), .b(G727), .O(gate248inter2));
  inv1  gate1040(.a(s_70), .O(gate248inter3));
  inv1  gate1041(.a(s_71), .O(gate248inter4));
  nand2 gate1042(.a(gate248inter4), .b(gate248inter3), .O(gate248inter5));
  nor2  gate1043(.a(gate248inter5), .b(gate248inter2), .O(gate248inter6));
  inv1  gate1044(.a(G727), .O(gate248inter7));
  inv1  gate1045(.a(G739), .O(gate248inter8));
  nand2 gate1046(.a(gate248inter8), .b(gate248inter7), .O(gate248inter9));
  nand2 gate1047(.a(s_71), .b(gate248inter3), .O(gate248inter10));
  nor2  gate1048(.a(gate248inter10), .b(gate248inter9), .O(gate248inter11));
  nor2  gate1049(.a(gate248inter11), .b(gate248inter6), .O(gate248inter12));
  nand2 gate1050(.a(gate248inter12), .b(gate248inter1), .O(G761));

  xor2  gate2087(.a(G742), .b(G254), .O(gate249inter0));
  nand2 gate2088(.a(gate249inter0), .b(s_220), .O(gate249inter1));
  and2  gate2089(.a(G742), .b(G254), .O(gate249inter2));
  inv1  gate2090(.a(s_220), .O(gate249inter3));
  inv1  gate2091(.a(s_221), .O(gate249inter4));
  nand2 gate2092(.a(gate249inter4), .b(gate249inter3), .O(gate249inter5));
  nor2  gate2093(.a(gate249inter5), .b(gate249inter2), .O(gate249inter6));
  inv1  gate2094(.a(G254), .O(gate249inter7));
  inv1  gate2095(.a(G742), .O(gate249inter8));
  nand2 gate2096(.a(gate249inter8), .b(gate249inter7), .O(gate249inter9));
  nand2 gate2097(.a(s_221), .b(gate249inter3), .O(gate249inter10));
  nor2  gate2098(.a(gate249inter10), .b(gate249inter9), .O(gate249inter11));
  nor2  gate2099(.a(gate249inter11), .b(gate249inter6), .O(gate249inter12));
  nand2 gate2100(.a(gate249inter12), .b(gate249inter1), .O(G762));
nand2 gate250( .a(G706), .b(G742), .O(G763) );

  xor2  gate1499(.a(G745), .b(G257), .O(gate251inter0));
  nand2 gate1500(.a(gate251inter0), .b(s_136), .O(gate251inter1));
  and2  gate1501(.a(G745), .b(G257), .O(gate251inter2));
  inv1  gate1502(.a(s_136), .O(gate251inter3));
  inv1  gate1503(.a(s_137), .O(gate251inter4));
  nand2 gate1504(.a(gate251inter4), .b(gate251inter3), .O(gate251inter5));
  nor2  gate1505(.a(gate251inter5), .b(gate251inter2), .O(gate251inter6));
  inv1  gate1506(.a(G257), .O(gate251inter7));
  inv1  gate1507(.a(G745), .O(gate251inter8));
  nand2 gate1508(.a(gate251inter8), .b(gate251inter7), .O(gate251inter9));
  nand2 gate1509(.a(s_137), .b(gate251inter3), .O(gate251inter10));
  nor2  gate1510(.a(gate251inter10), .b(gate251inter9), .O(gate251inter11));
  nor2  gate1511(.a(gate251inter11), .b(gate251inter6), .O(gate251inter12));
  nand2 gate1512(.a(gate251inter12), .b(gate251inter1), .O(G764));
nand2 gate252( .a(G709), .b(G745), .O(G765) );
nand2 gate253( .a(G260), .b(G748), .O(G766) );
nand2 gate254( .a(G712), .b(G748), .O(G767) );
nand2 gate255( .a(G263), .b(G751), .O(G768) );

  xor2  gate2073(.a(G751), .b(G715), .O(gate256inter0));
  nand2 gate2074(.a(gate256inter0), .b(s_218), .O(gate256inter1));
  and2  gate2075(.a(G751), .b(G715), .O(gate256inter2));
  inv1  gate2076(.a(s_218), .O(gate256inter3));
  inv1  gate2077(.a(s_219), .O(gate256inter4));
  nand2 gate2078(.a(gate256inter4), .b(gate256inter3), .O(gate256inter5));
  nor2  gate2079(.a(gate256inter5), .b(gate256inter2), .O(gate256inter6));
  inv1  gate2080(.a(G715), .O(gate256inter7));
  inv1  gate2081(.a(G751), .O(gate256inter8));
  nand2 gate2082(.a(gate256inter8), .b(gate256inter7), .O(gate256inter9));
  nand2 gate2083(.a(s_219), .b(gate256inter3), .O(gate256inter10));
  nor2  gate2084(.a(gate256inter10), .b(gate256inter9), .O(gate256inter11));
  nor2  gate2085(.a(gate256inter11), .b(gate256inter6), .O(gate256inter12));
  nand2 gate2086(.a(gate256inter12), .b(gate256inter1), .O(G769));
nand2 gate257( .a(G754), .b(G755), .O(G770) );

  xor2  gate2507(.a(G757), .b(G756), .O(gate258inter0));
  nand2 gate2508(.a(gate258inter0), .b(s_280), .O(gate258inter1));
  and2  gate2509(.a(G757), .b(G756), .O(gate258inter2));
  inv1  gate2510(.a(s_280), .O(gate258inter3));
  inv1  gate2511(.a(s_281), .O(gate258inter4));
  nand2 gate2512(.a(gate258inter4), .b(gate258inter3), .O(gate258inter5));
  nor2  gate2513(.a(gate258inter5), .b(gate258inter2), .O(gate258inter6));
  inv1  gate2514(.a(G756), .O(gate258inter7));
  inv1  gate2515(.a(G757), .O(gate258inter8));
  nand2 gate2516(.a(gate258inter8), .b(gate258inter7), .O(gate258inter9));
  nand2 gate2517(.a(s_281), .b(gate258inter3), .O(gate258inter10));
  nor2  gate2518(.a(gate258inter10), .b(gate258inter9), .O(gate258inter11));
  nor2  gate2519(.a(gate258inter11), .b(gate258inter6), .O(gate258inter12));
  nand2 gate2520(.a(gate258inter12), .b(gate258inter1), .O(G773));
nand2 gate259( .a(G758), .b(G759), .O(G776) );

  xor2  gate925(.a(G761), .b(G760), .O(gate260inter0));
  nand2 gate926(.a(gate260inter0), .b(s_54), .O(gate260inter1));
  and2  gate927(.a(G761), .b(G760), .O(gate260inter2));
  inv1  gate928(.a(s_54), .O(gate260inter3));
  inv1  gate929(.a(s_55), .O(gate260inter4));
  nand2 gate930(.a(gate260inter4), .b(gate260inter3), .O(gate260inter5));
  nor2  gate931(.a(gate260inter5), .b(gate260inter2), .O(gate260inter6));
  inv1  gate932(.a(G760), .O(gate260inter7));
  inv1  gate933(.a(G761), .O(gate260inter8));
  nand2 gate934(.a(gate260inter8), .b(gate260inter7), .O(gate260inter9));
  nand2 gate935(.a(s_55), .b(gate260inter3), .O(gate260inter10));
  nor2  gate936(.a(gate260inter10), .b(gate260inter9), .O(gate260inter11));
  nor2  gate937(.a(gate260inter11), .b(gate260inter6), .O(gate260inter12));
  nand2 gate938(.a(gate260inter12), .b(gate260inter1), .O(G779));
nand2 gate261( .a(G762), .b(G763), .O(G782) );
nand2 gate262( .a(G764), .b(G765), .O(G785) );
nand2 gate263( .a(G766), .b(G767), .O(G788) );

  xor2  gate1653(.a(G769), .b(G768), .O(gate264inter0));
  nand2 gate1654(.a(gate264inter0), .b(s_158), .O(gate264inter1));
  and2  gate1655(.a(G769), .b(G768), .O(gate264inter2));
  inv1  gate1656(.a(s_158), .O(gate264inter3));
  inv1  gate1657(.a(s_159), .O(gate264inter4));
  nand2 gate1658(.a(gate264inter4), .b(gate264inter3), .O(gate264inter5));
  nor2  gate1659(.a(gate264inter5), .b(gate264inter2), .O(gate264inter6));
  inv1  gate1660(.a(G768), .O(gate264inter7));
  inv1  gate1661(.a(G769), .O(gate264inter8));
  nand2 gate1662(.a(gate264inter8), .b(gate264inter7), .O(gate264inter9));
  nand2 gate1663(.a(s_159), .b(gate264inter3), .O(gate264inter10));
  nor2  gate1664(.a(gate264inter10), .b(gate264inter9), .O(gate264inter11));
  nor2  gate1665(.a(gate264inter11), .b(gate264inter6), .O(gate264inter12));
  nand2 gate1666(.a(gate264inter12), .b(gate264inter1), .O(G791));

  xor2  gate2563(.a(G770), .b(G642), .O(gate265inter0));
  nand2 gate2564(.a(gate265inter0), .b(s_288), .O(gate265inter1));
  and2  gate2565(.a(G770), .b(G642), .O(gate265inter2));
  inv1  gate2566(.a(s_288), .O(gate265inter3));
  inv1  gate2567(.a(s_289), .O(gate265inter4));
  nand2 gate2568(.a(gate265inter4), .b(gate265inter3), .O(gate265inter5));
  nor2  gate2569(.a(gate265inter5), .b(gate265inter2), .O(gate265inter6));
  inv1  gate2570(.a(G642), .O(gate265inter7));
  inv1  gate2571(.a(G770), .O(gate265inter8));
  nand2 gate2572(.a(gate265inter8), .b(gate265inter7), .O(gate265inter9));
  nand2 gate2573(.a(s_289), .b(gate265inter3), .O(gate265inter10));
  nor2  gate2574(.a(gate265inter10), .b(gate265inter9), .O(gate265inter11));
  nor2  gate2575(.a(gate265inter11), .b(gate265inter6), .O(gate265inter12));
  nand2 gate2576(.a(gate265inter12), .b(gate265inter1), .O(G794));

  xor2  gate701(.a(G773), .b(G645), .O(gate266inter0));
  nand2 gate702(.a(gate266inter0), .b(s_22), .O(gate266inter1));
  and2  gate703(.a(G773), .b(G645), .O(gate266inter2));
  inv1  gate704(.a(s_22), .O(gate266inter3));
  inv1  gate705(.a(s_23), .O(gate266inter4));
  nand2 gate706(.a(gate266inter4), .b(gate266inter3), .O(gate266inter5));
  nor2  gate707(.a(gate266inter5), .b(gate266inter2), .O(gate266inter6));
  inv1  gate708(.a(G645), .O(gate266inter7));
  inv1  gate709(.a(G773), .O(gate266inter8));
  nand2 gate710(.a(gate266inter8), .b(gate266inter7), .O(gate266inter9));
  nand2 gate711(.a(s_23), .b(gate266inter3), .O(gate266inter10));
  nor2  gate712(.a(gate266inter10), .b(gate266inter9), .O(gate266inter11));
  nor2  gate713(.a(gate266inter11), .b(gate266inter6), .O(gate266inter12));
  nand2 gate714(.a(gate266inter12), .b(gate266inter1), .O(G797));
nand2 gate267( .a(G648), .b(G776), .O(G800) );
nand2 gate268( .a(G651), .b(G779), .O(G803) );
nand2 gate269( .a(G654), .b(G782), .O(G806) );
nand2 gate270( .a(G657), .b(G785), .O(G809) );
nand2 gate271( .a(G660), .b(G788), .O(G812) );
nand2 gate272( .a(G663), .b(G791), .O(G815) );
nand2 gate273( .a(G642), .b(G794), .O(G818) );
nand2 gate274( .a(G770), .b(G794), .O(G819) );

  xor2  gate2269(.a(G797), .b(G645), .O(gate275inter0));
  nand2 gate2270(.a(gate275inter0), .b(s_246), .O(gate275inter1));
  and2  gate2271(.a(G797), .b(G645), .O(gate275inter2));
  inv1  gate2272(.a(s_246), .O(gate275inter3));
  inv1  gate2273(.a(s_247), .O(gate275inter4));
  nand2 gate2274(.a(gate275inter4), .b(gate275inter3), .O(gate275inter5));
  nor2  gate2275(.a(gate275inter5), .b(gate275inter2), .O(gate275inter6));
  inv1  gate2276(.a(G645), .O(gate275inter7));
  inv1  gate2277(.a(G797), .O(gate275inter8));
  nand2 gate2278(.a(gate275inter8), .b(gate275inter7), .O(gate275inter9));
  nand2 gate2279(.a(s_247), .b(gate275inter3), .O(gate275inter10));
  nor2  gate2280(.a(gate275inter10), .b(gate275inter9), .O(gate275inter11));
  nor2  gate2281(.a(gate275inter11), .b(gate275inter6), .O(gate275inter12));
  nand2 gate2282(.a(gate275inter12), .b(gate275inter1), .O(G820));
nand2 gate276( .a(G773), .b(G797), .O(G821) );
nand2 gate277( .a(G648), .b(G800), .O(G822) );

  xor2  gate1443(.a(G800), .b(G776), .O(gate278inter0));
  nand2 gate1444(.a(gate278inter0), .b(s_128), .O(gate278inter1));
  and2  gate1445(.a(G800), .b(G776), .O(gate278inter2));
  inv1  gate1446(.a(s_128), .O(gate278inter3));
  inv1  gate1447(.a(s_129), .O(gate278inter4));
  nand2 gate1448(.a(gate278inter4), .b(gate278inter3), .O(gate278inter5));
  nor2  gate1449(.a(gate278inter5), .b(gate278inter2), .O(gate278inter6));
  inv1  gate1450(.a(G776), .O(gate278inter7));
  inv1  gate1451(.a(G800), .O(gate278inter8));
  nand2 gate1452(.a(gate278inter8), .b(gate278inter7), .O(gate278inter9));
  nand2 gate1453(.a(s_129), .b(gate278inter3), .O(gate278inter10));
  nor2  gate1454(.a(gate278inter10), .b(gate278inter9), .O(gate278inter11));
  nor2  gate1455(.a(gate278inter11), .b(gate278inter6), .O(gate278inter12));
  nand2 gate1456(.a(gate278inter12), .b(gate278inter1), .O(G823));
nand2 gate279( .a(G651), .b(G803), .O(G824) );

  xor2  gate757(.a(G803), .b(G779), .O(gate280inter0));
  nand2 gate758(.a(gate280inter0), .b(s_30), .O(gate280inter1));
  and2  gate759(.a(G803), .b(G779), .O(gate280inter2));
  inv1  gate760(.a(s_30), .O(gate280inter3));
  inv1  gate761(.a(s_31), .O(gate280inter4));
  nand2 gate762(.a(gate280inter4), .b(gate280inter3), .O(gate280inter5));
  nor2  gate763(.a(gate280inter5), .b(gate280inter2), .O(gate280inter6));
  inv1  gate764(.a(G779), .O(gate280inter7));
  inv1  gate765(.a(G803), .O(gate280inter8));
  nand2 gate766(.a(gate280inter8), .b(gate280inter7), .O(gate280inter9));
  nand2 gate767(.a(s_31), .b(gate280inter3), .O(gate280inter10));
  nor2  gate768(.a(gate280inter10), .b(gate280inter9), .O(gate280inter11));
  nor2  gate769(.a(gate280inter11), .b(gate280inter6), .O(gate280inter12));
  nand2 gate770(.a(gate280inter12), .b(gate280inter1), .O(G825));

  xor2  gate2101(.a(G806), .b(G654), .O(gate281inter0));
  nand2 gate2102(.a(gate281inter0), .b(s_222), .O(gate281inter1));
  and2  gate2103(.a(G806), .b(G654), .O(gate281inter2));
  inv1  gate2104(.a(s_222), .O(gate281inter3));
  inv1  gate2105(.a(s_223), .O(gate281inter4));
  nand2 gate2106(.a(gate281inter4), .b(gate281inter3), .O(gate281inter5));
  nor2  gate2107(.a(gate281inter5), .b(gate281inter2), .O(gate281inter6));
  inv1  gate2108(.a(G654), .O(gate281inter7));
  inv1  gate2109(.a(G806), .O(gate281inter8));
  nand2 gate2110(.a(gate281inter8), .b(gate281inter7), .O(gate281inter9));
  nand2 gate2111(.a(s_223), .b(gate281inter3), .O(gate281inter10));
  nor2  gate2112(.a(gate281inter10), .b(gate281inter9), .O(gate281inter11));
  nor2  gate2113(.a(gate281inter11), .b(gate281inter6), .O(gate281inter12));
  nand2 gate2114(.a(gate281inter12), .b(gate281inter1), .O(G826));
nand2 gate282( .a(G782), .b(G806), .O(G827) );

  xor2  gate2227(.a(G809), .b(G657), .O(gate283inter0));
  nand2 gate2228(.a(gate283inter0), .b(s_240), .O(gate283inter1));
  and2  gate2229(.a(G809), .b(G657), .O(gate283inter2));
  inv1  gate2230(.a(s_240), .O(gate283inter3));
  inv1  gate2231(.a(s_241), .O(gate283inter4));
  nand2 gate2232(.a(gate283inter4), .b(gate283inter3), .O(gate283inter5));
  nor2  gate2233(.a(gate283inter5), .b(gate283inter2), .O(gate283inter6));
  inv1  gate2234(.a(G657), .O(gate283inter7));
  inv1  gate2235(.a(G809), .O(gate283inter8));
  nand2 gate2236(.a(gate283inter8), .b(gate283inter7), .O(gate283inter9));
  nand2 gate2237(.a(s_241), .b(gate283inter3), .O(gate283inter10));
  nor2  gate2238(.a(gate283inter10), .b(gate283inter9), .O(gate283inter11));
  nor2  gate2239(.a(gate283inter11), .b(gate283inter6), .O(gate283inter12));
  nand2 gate2240(.a(gate283inter12), .b(gate283inter1), .O(G828));

  xor2  gate631(.a(G809), .b(G785), .O(gate284inter0));
  nand2 gate632(.a(gate284inter0), .b(s_12), .O(gate284inter1));
  and2  gate633(.a(G809), .b(G785), .O(gate284inter2));
  inv1  gate634(.a(s_12), .O(gate284inter3));
  inv1  gate635(.a(s_13), .O(gate284inter4));
  nand2 gate636(.a(gate284inter4), .b(gate284inter3), .O(gate284inter5));
  nor2  gate637(.a(gate284inter5), .b(gate284inter2), .O(gate284inter6));
  inv1  gate638(.a(G785), .O(gate284inter7));
  inv1  gate639(.a(G809), .O(gate284inter8));
  nand2 gate640(.a(gate284inter8), .b(gate284inter7), .O(gate284inter9));
  nand2 gate641(.a(s_13), .b(gate284inter3), .O(gate284inter10));
  nor2  gate642(.a(gate284inter10), .b(gate284inter9), .O(gate284inter11));
  nor2  gate643(.a(gate284inter11), .b(gate284inter6), .O(gate284inter12));
  nand2 gate644(.a(gate284inter12), .b(gate284inter1), .O(G829));

  xor2  gate1555(.a(G812), .b(G660), .O(gate285inter0));
  nand2 gate1556(.a(gate285inter0), .b(s_144), .O(gate285inter1));
  and2  gate1557(.a(G812), .b(G660), .O(gate285inter2));
  inv1  gate1558(.a(s_144), .O(gate285inter3));
  inv1  gate1559(.a(s_145), .O(gate285inter4));
  nand2 gate1560(.a(gate285inter4), .b(gate285inter3), .O(gate285inter5));
  nor2  gate1561(.a(gate285inter5), .b(gate285inter2), .O(gate285inter6));
  inv1  gate1562(.a(G660), .O(gate285inter7));
  inv1  gate1563(.a(G812), .O(gate285inter8));
  nand2 gate1564(.a(gate285inter8), .b(gate285inter7), .O(gate285inter9));
  nand2 gate1565(.a(s_145), .b(gate285inter3), .O(gate285inter10));
  nor2  gate1566(.a(gate285inter10), .b(gate285inter9), .O(gate285inter11));
  nor2  gate1567(.a(gate285inter11), .b(gate285inter6), .O(gate285inter12));
  nand2 gate1568(.a(gate285inter12), .b(gate285inter1), .O(G830));

  xor2  gate2913(.a(G812), .b(G788), .O(gate286inter0));
  nand2 gate2914(.a(gate286inter0), .b(s_338), .O(gate286inter1));
  and2  gate2915(.a(G812), .b(G788), .O(gate286inter2));
  inv1  gate2916(.a(s_338), .O(gate286inter3));
  inv1  gate2917(.a(s_339), .O(gate286inter4));
  nand2 gate2918(.a(gate286inter4), .b(gate286inter3), .O(gate286inter5));
  nor2  gate2919(.a(gate286inter5), .b(gate286inter2), .O(gate286inter6));
  inv1  gate2920(.a(G788), .O(gate286inter7));
  inv1  gate2921(.a(G812), .O(gate286inter8));
  nand2 gate2922(.a(gate286inter8), .b(gate286inter7), .O(gate286inter9));
  nand2 gate2923(.a(s_339), .b(gate286inter3), .O(gate286inter10));
  nor2  gate2924(.a(gate286inter10), .b(gate286inter9), .O(gate286inter11));
  nor2  gate2925(.a(gate286inter11), .b(gate286inter6), .O(gate286inter12));
  nand2 gate2926(.a(gate286inter12), .b(gate286inter1), .O(G831));
nand2 gate287( .a(G663), .b(G815), .O(G832) );
nand2 gate288( .a(G791), .b(G815), .O(G833) );

  xor2  gate2955(.a(G819), .b(G818), .O(gate289inter0));
  nand2 gate2956(.a(gate289inter0), .b(s_344), .O(gate289inter1));
  and2  gate2957(.a(G819), .b(G818), .O(gate289inter2));
  inv1  gate2958(.a(s_344), .O(gate289inter3));
  inv1  gate2959(.a(s_345), .O(gate289inter4));
  nand2 gate2960(.a(gate289inter4), .b(gate289inter3), .O(gate289inter5));
  nor2  gate2961(.a(gate289inter5), .b(gate289inter2), .O(gate289inter6));
  inv1  gate2962(.a(G818), .O(gate289inter7));
  inv1  gate2963(.a(G819), .O(gate289inter8));
  nand2 gate2964(.a(gate289inter8), .b(gate289inter7), .O(gate289inter9));
  nand2 gate2965(.a(s_345), .b(gate289inter3), .O(gate289inter10));
  nor2  gate2966(.a(gate289inter10), .b(gate289inter9), .O(gate289inter11));
  nor2  gate2967(.a(gate289inter11), .b(gate289inter6), .O(gate289inter12));
  nand2 gate2968(.a(gate289inter12), .b(gate289inter1), .O(G834));

  xor2  gate1821(.a(G821), .b(G820), .O(gate290inter0));
  nand2 gate1822(.a(gate290inter0), .b(s_182), .O(gate290inter1));
  and2  gate1823(.a(G821), .b(G820), .O(gate290inter2));
  inv1  gate1824(.a(s_182), .O(gate290inter3));
  inv1  gate1825(.a(s_183), .O(gate290inter4));
  nand2 gate1826(.a(gate290inter4), .b(gate290inter3), .O(gate290inter5));
  nor2  gate1827(.a(gate290inter5), .b(gate290inter2), .O(gate290inter6));
  inv1  gate1828(.a(G820), .O(gate290inter7));
  inv1  gate1829(.a(G821), .O(gate290inter8));
  nand2 gate1830(.a(gate290inter8), .b(gate290inter7), .O(gate290inter9));
  nand2 gate1831(.a(s_183), .b(gate290inter3), .O(gate290inter10));
  nor2  gate1832(.a(gate290inter10), .b(gate290inter9), .O(gate290inter11));
  nor2  gate1833(.a(gate290inter11), .b(gate290inter6), .O(gate290inter12));
  nand2 gate1834(.a(gate290inter12), .b(gate290inter1), .O(G847));
nand2 gate291( .a(G822), .b(G823), .O(G860) );

  xor2  gate603(.a(G825), .b(G824), .O(gate292inter0));
  nand2 gate604(.a(gate292inter0), .b(s_8), .O(gate292inter1));
  and2  gate605(.a(G825), .b(G824), .O(gate292inter2));
  inv1  gate606(.a(s_8), .O(gate292inter3));
  inv1  gate607(.a(s_9), .O(gate292inter4));
  nand2 gate608(.a(gate292inter4), .b(gate292inter3), .O(gate292inter5));
  nor2  gate609(.a(gate292inter5), .b(gate292inter2), .O(gate292inter6));
  inv1  gate610(.a(G824), .O(gate292inter7));
  inv1  gate611(.a(G825), .O(gate292inter8));
  nand2 gate612(.a(gate292inter8), .b(gate292inter7), .O(gate292inter9));
  nand2 gate613(.a(s_9), .b(gate292inter3), .O(gate292inter10));
  nor2  gate614(.a(gate292inter10), .b(gate292inter9), .O(gate292inter11));
  nor2  gate615(.a(gate292inter11), .b(gate292inter6), .O(gate292inter12));
  nand2 gate616(.a(gate292inter12), .b(gate292inter1), .O(G873));
nand2 gate293( .a(G828), .b(G829), .O(G886) );

  xor2  gate575(.a(G833), .b(G832), .O(gate294inter0));
  nand2 gate576(.a(gate294inter0), .b(s_4), .O(gate294inter1));
  and2  gate577(.a(G833), .b(G832), .O(gate294inter2));
  inv1  gate578(.a(s_4), .O(gate294inter3));
  inv1  gate579(.a(s_5), .O(gate294inter4));
  nand2 gate580(.a(gate294inter4), .b(gate294inter3), .O(gate294inter5));
  nor2  gate581(.a(gate294inter5), .b(gate294inter2), .O(gate294inter6));
  inv1  gate582(.a(G832), .O(gate294inter7));
  inv1  gate583(.a(G833), .O(gate294inter8));
  nand2 gate584(.a(gate294inter8), .b(gate294inter7), .O(gate294inter9));
  nand2 gate585(.a(s_5), .b(gate294inter3), .O(gate294inter10));
  nor2  gate586(.a(gate294inter10), .b(gate294inter9), .O(gate294inter11));
  nor2  gate587(.a(gate294inter11), .b(gate294inter6), .O(gate294inter12));
  nand2 gate588(.a(gate294inter12), .b(gate294inter1), .O(G899));
nand2 gate295( .a(G830), .b(G831), .O(G912) );

  xor2  gate715(.a(G827), .b(G826), .O(gate296inter0));
  nand2 gate716(.a(gate296inter0), .b(s_24), .O(gate296inter1));
  and2  gate717(.a(G827), .b(G826), .O(gate296inter2));
  inv1  gate718(.a(s_24), .O(gate296inter3));
  inv1  gate719(.a(s_25), .O(gate296inter4));
  nand2 gate720(.a(gate296inter4), .b(gate296inter3), .O(gate296inter5));
  nor2  gate721(.a(gate296inter5), .b(gate296inter2), .O(gate296inter6));
  inv1  gate722(.a(G826), .O(gate296inter7));
  inv1  gate723(.a(G827), .O(gate296inter8));
  nand2 gate724(.a(gate296inter8), .b(gate296inter7), .O(gate296inter9));
  nand2 gate725(.a(s_25), .b(gate296inter3), .O(gate296inter10));
  nor2  gate726(.a(gate296inter10), .b(gate296inter9), .O(gate296inter11));
  nor2  gate727(.a(gate296inter11), .b(gate296inter6), .O(gate296inter12));
  nand2 gate728(.a(gate296inter12), .b(gate296inter1), .O(G925));
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );

  xor2  gate813(.a(G1036), .b(G1), .O(gate387inter0));
  nand2 gate814(.a(gate387inter0), .b(s_38), .O(gate387inter1));
  and2  gate815(.a(G1036), .b(G1), .O(gate387inter2));
  inv1  gate816(.a(s_38), .O(gate387inter3));
  inv1  gate817(.a(s_39), .O(gate387inter4));
  nand2 gate818(.a(gate387inter4), .b(gate387inter3), .O(gate387inter5));
  nor2  gate819(.a(gate387inter5), .b(gate387inter2), .O(gate387inter6));
  inv1  gate820(.a(G1), .O(gate387inter7));
  inv1  gate821(.a(G1036), .O(gate387inter8));
  nand2 gate822(.a(gate387inter8), .b(gate387inter7), .O(gate387inter9));
  nand2 gate823(.a(s_39), .b(gate387inter3), .O(gate387inter10));
  nor2  gate824(.a(gate387inter10), .b(gate387inter9), .O(gate387inter11));
  nor2  gate825(.a(gate387inter11), .b(gate387inter6), .O(gate387inter12));
  nand2 gate826(.a(gate387inter12), .b(gate387inter1), .O(G1132));
nand2 gate388( .a(G2), .b(G1039), .O(G1135) );

  xor2  gate2367(.a(G1042), .b(G3), .O(gate389inter0));
  nand2 gate2368(.a(gate389inter0), .b(s_260), .O(gate389inter1));
  and2  gate2369(.a(G1042), .b(G3), .O(gate389inter2));
  inv1  gate2370(.a(s_260), .O(gate389inter3));
  inv1  gate2371(.a(s_261), .O(gate389inter4));
  nand2 gate2372(.a(gate389inter4), .b(gate389inter3), .O(gate389inter5));
  nor2  gate2373(.a(gate389inter5), .b(gate389inter2), .O(gate389inter6));
  inv1  gate2374(.a(G3), .O(gate389inter7));
  inv1  gate2375(.a(G1042), .O(gate389inter8));
  nand2 gate2376(.a(gate389inter8), .b(gate389inter7), .O(gate389inter9));
  nand2 gate2377(.a(s_261), .b(gate389inter3), .O(gate389inter10));
  nor2  gate2378(.a(gate389inter10), .b(gate389inter9), .O(gate389inter11));
  nor2  gate2379(.a(gate389inter11), .b(gate389inter6), .O(gate389inter12));
  nand2 gate2380(.a(gate389inter12), .b(gate389inter1), .O(G1138));
nand2 gate390( .a(G4), .b(G1045), .O(G1141) );
nand2 gate391( .a(G5), .b(G1048), .O(G1144) );
nand2 gate392( .a(G6), .b(G1051), .O(G1147) );
nand2 gate393( .a(G7), .b(G1054), .O(G1150) );
nand2 gate394( .a(G8), .b(G1057), .O(G1153) );
nand2 gate395( .a(G9), .b(G1060), .O(G1156) );

  xor2  gate2521(.a(G1063), .b(G10), .O(gate396inter0));
  nand2 gate2522(.a(gate396inter0), .b(s_282), .O(gate396inter1));
  and2  gate2523(.a(G1063), .b(G10), .O(gate396inter2));
  inv1  gate2524(.a(s_282), .O(gate396inter3));
  inv1  gate2525(.a(s_283), .O(gate396inter4));
  nand2 gate2526(.a(gate396inter4), .b(gate396inter3), .O(gate396inter5));
  nor2  gate2527(.a(gate396inter5), .b(gate396inter2), .O(gate396inter6));
  inv1  gate2528(.a(G10), .O(gate396inter7));
  inv1  gate2529(.a(G1063), .O(gate396inter8));
  nand2 gate2530(.a(gate396inter8), .b(gate396inter7), .O(gate396inter9));
  nand2 gate2531(.a(s_283), .b(gate396inter3), .O(gate396inter10));
  nor2  gate2532(.a(gate396inter10), .b(gate396inter9), .O(gate396inter11));
  nor2  gate2533(.a(gate396inter11), .b(gate396inter6), .O(gate396inter12));
  nand2 gate2534(.a(gate396inter12), .b(gate396inter1), .O(G1159));
nand2 gate397( .a(G11), .b(G1066), .O(G1162) );
nand2 gate398( .a(G12), .b(G1069), .O(G1165) );

  xor2  gate1219(.a(G1072), .b(G13), .O(gate399inter0));
  nand2 gate1220(.a(gate399inter0), .b(s_96), .O(gate399inter1));
  and2  gate1221(.a(G1072), .b(G13), .O(gate399inter2));
  inv1  gate1222(.a(s_96), .O(gate399inter3));
  inv1  gate1223(.a(s_97), .O(gate399inter4));
  nand2 gate1224(.a(gate399inter4), .b(gate399inter3), .O(gate399inter5));
  nor2  gate1225(.a(gate399inter5), .b(gate399inter2), .O(gate399inter6));
  inv1  gate1226(.a(G13), .O(gate399inter7));
  inv1  gate1227(.a(G1072), .O(gate399inter8));
  nand2 gate1228(.a(gate399inter8), .b(gate399inter7), .O(gate399inter9));
  nand2 gate1229(.a(s_97), .b(gate399inter3), .O(gate399inter10));
  nor2  gate1230(.a(gate399inter10), .b(gate399inter9), .O(gate399inter11));
  nor2  gate1231(.a(gate399inter11), .b(gate399inter6), .O(gate399inter12));
  nand2 gate1232(.a(gate399inter12), .b(gate399inter1), .O(G1168));

  xor2  gate659(.a(G1075), .b(G14), .O(gate400inter0));
  nand2 gate660(.a(gate400inter0), .b(s_16), .O(gate400inter1));
  and2  gate661(.a(G1075), .b(G14), .O(gate400inter2));
  inv1  gate662(.a(s_16), .O(gate400inter3));
  inv1  gate663(.a(s_17), .O(gate400inter4));
  nand2 gate664(.a(gate400inter4), .b(gate400inter3), .O(gate400inter5));
  nor2  gate665(.a(gate400inter5), .b(gate400inter2), .O(gate400inter6));
  inv1  gate666(.a(G14), .O(gate400inter7));
  inv1  gate667(.a(G1075), .O(gate400inter8));
  nand2 gate668(.a(gate400inter8), .b(gate400inter7), .O(gate400inter9));
  nand2 gate669(.a(s_17), .b(gate400inter3), .O(gate400inter10));
  nor2  gate670(.a(gate400inter10), .b(gate400inter9), .O(gate400inter11));
  nor2  gate671(.a(gate400inter11), .b(gate400inter6), .O(gate400inter12));
  nand2 gate672(.a(gate400inter12), .b(gate400inter1), .O(G1171));
nand2 gate401( .a(G15), .b(G1078), .O(G1174) );
nand2 gate402( .a(G16), .b(G1081), .O(G1177) );
nand2 gate403( .a(G17), .b(G1084), .O(G1180) );

  xor2  gate2899(.a(G1087), .b(G18), .O(gate404inter0));
  nand2 gate2900(.a(gate404inter0), .b(s_336), .O(gate404inter1));
  and2  gate2901(.a(G1087), .b(G18), .O(gate404inter2));
  inv1  gate2902(.a(s_336), .O(gate404inter3));
  inv1  gate2903(.a(s_337), .O(gate404inter4));
  nand2 gate2904(.a(gate404inter4), .b(gate404inter3), .O(gate404inter5));
  nor2  gate2905(.a(gate404inter5), .b(gate404inter2), .O(gate404inter6));
  inv1  gate2906(.a(G18), .O(gate404inter7));
  inv1  gate2907(.a(G1087), .O(gate404inter8));
  nand2 gate2908(.a(gate404inter8), .b(gate404inter7), .O(gate404inter9));
  nand2 gate2909(.a(s_337), .b(gate404inter3), .O(gate404inter10));
  nor2  gate2910(.a(gate404inter10), .b(gate404inter9), .O(gate404inter11));
  nor2  gate2911(.a(gate404inter11), .b(gate404inter6), .O(gate404inter12));
  nand2 gate2912(.a(gate404inter12), .b(gate404inter1), .O(G1183));

  xor2  gate855(.a(G1090), .b(G19), .O(gate405inter0));
  nand2 gate856(.a(gate405inter0), .b(s_44), .O(gate405inter1));
  and2  gate857(.a(G1090), .b(G19), .O(gate405inter2));
  inv1  gate858(.a(s_44), .O(gate405inter3));
  inv1  gate859(.a(s_45), .O(gate405inter4));
  nand2 gate860(.a(gate405inter4), .b(gate405inter3), .O(gate405inter5));
  nor2  gate861(.a(gate405inter5), .b(gate405inter2), .O(gate405inter6));
  inv1  gate862(.a(G19), .O(gate405inter7));
  inv1  gate863(.a(G1090), .O(gate405inter8));
  nand2 gate864(.a(gate405inter8), .b(gate405inter7), .O(gate405inter9));
  nand2 gate865(.a(s_45), .b(gate405inter3), .O(gate405inter10));
  nor2  gate866(.a(gate405inter10), .b(gate405inter9), .O(gate405inter11));
  nor2  gate867(.a(gate405inter11), .b(gate405inter6), .O(gate405inter12));
  nand2 gate868(.a(gate405inter12), .b(gate405inter1), .O(G1186));
nand2 gate406( .a(G20), .b(G1093), .O(G1189) );
nand2 gate407( .a(G21), .b(G1096), .O(G1192) );

  xor2  gate771(.a(G1099), .b(G22), .O(gate408inter0));
  nand2 gate772(.a(gate408inter0), .b(s_32), .O(gate408inter1));
  and2  gate773(.a(G1099), .b(G22), .O(gate408inter2));
  inv1  gate774(.a(s_32), .O(gate408inter3));
  inv1  gate775(.a(s_33), .O(gate408inter4));
  nand2 gate776(.a(gate408inter4), .b(gate408inter3), .O(gate408inter5));
  nor2  gate777(.a(gate408inter5), .b(gate408inter2), .O(gate408inter6));
  inv1  gate778(.a(G22), .O(gate408inter7));
  inv1  gate779(.a(G1099), .O(gate408inter8));
  nand2 gate780(.a(gate408inter8), .b(gate408inter7), .O(gate408inter9));
  nand2 gate781(.a(s_33), .b(gate408inter3), .O(gate408inter10));
  nor2  gate782(.a(gate408inter10), .b(gate408inter9), .O(gate408inter11));
  nor2  gate783(.a(gate408inter11), .b(gate408inter6), .O(gate408inter12));
  nand2 gate784(.a(gate408inter12), .b(gate408inter1), .O(G1195));

  xor2  gate2997(.a(G1102), .b(G23), .O(gate409inter0));
  nand2 gate2998(.a(gate409inter0), .b(s_350), .O(gate409inter1));
  and2  gate2999(.a(G1102), .b(G23), .O(gate409inter2));
  inv1  gate3000(.a(s_350), .O(gate409inter3));
  inv1  gate3001(.a(s_351), .O(gate409inter4));
  nand2 gate3002(.a(gate409inter4), .b(gate409inter3), .O(gate409inter5));
  nor2  gate3003(.a(gate409inter5), .b(gate409inter2), .O(gate409inter6));
  inv1  gate3004(.a(G23), .O(gate409inter7));
  inv1  gate3005(.a(G1102), .O(gate409inter8));
  nand2 gate3006(.a(gate409inter8), .b(gate409inter7), .O(gate409inter9));
  nand2 gate3007(.a(s_351), .b(gate409inter3), .O(gate409inter10));
  nor2  gate3008(.a(gate409inter10), .b(gate409inter9), .O(gate409inter11));
  nor2  gate3009(.a(gate409inter11), .b(gate409inter6), .O(gate409inter12));
  nand2 gate3010(.a(gate409inter12), .b(gate409inter1), .O(G1198));

  xor2  gate869(.a(G1105), .b(G24), .O(gate410inter0));
  nand2 gate870(.a(gate410inter0), .b(s_46), .O(gate410inter1));
  and2  gate871(.a(G1105), .b(G24), .O(gate410inter2));
  inv1  gate872(.a(s_46), .O(gate410inter3));
  inv1  gate873(.a(s_47), .O(gate410inter4));
  nand2 gate874(.a(gate410inter4), .b(gate410inter3), .O(gate410inter5));
  nor2  gate875(.a(gate410inter5), .b(gate410inter2), .O(gate410inter6));
  inv1  gate876(.a(G24), .O(gate410inter7));
  inv1  gate877(.a(G1105), .O(gate410inter8));
  nand2 gate878(.a(gate410inter8), .b(gate410inter7), .O(gate410inter9));
  nand2 gate879(.a(s_47), .b(gate410inter3), .O(gate410inter10));
  nor2  gate880(.a(gate410inter10), .b(gate410inter9), .O(gate410inter11));
  nor2  gate881(.a(gate410inter11), .b(gate410inter6), .O(gate410inter12));
  nand2 gate882(.a(gate410inter12), .b(gate410inter1), .O(G1201));
nand2 gate411( .a(G25), .b(G1108), .O(G1204) );

  xor2  gate2381(.a(G1111), .b(G26), .O(gate412inter0));
  nand2 gate2382(.a(gate412inter0), .b(s_262), .O(gate412inter1));
  and2  gate2383(.a(G1111), .b(G26), .O(gate412inter2));
  inv1  gate2384(.a(s_262), .O(gate412inter3));
  inv1  gate2385(.a(s_263), .O(gate412inter4));
  nand2 gate2386(.a(gate412inter4), .b(gate412inter3), .O(gate412inter5));
  nor2  gate2387(.a(gate412inter5), .b(gate412inter2), .O(gate412inter6));
  inv1  gate2388(.a(G26), .O(gate412inter7));
  inv1  gate2389(.a(G1111), .O(gate412inter8));
  nand2 gate2390(.a(gate412inter8), .b(gate412inter7), .O(gate412inter9));
  nand2 gate2391(.a(s_263), .b(gate412inter3), .O(gate412inter10));
  nor2  gate2392(.a(gate412inter10), .b(gate412inter9), .O(gate412inter11));
  nor2  gate2393(.a(gate412inter11), .b(gate412inter6), .O(gate412inter12));
  nand2 gate2394(.a(gate412inter12), .b(gate412inter1), .O(G1207));

  xor2  gate687(.a(G1114), .b(G27), .O(gate413inter0));
  nand2 gate688(.a(gate413inter0), .b(s_20), .O(gate413inter1));
  and2  gate689(.a(G1114), .b(G27), .O(gate413inter2));
  inv1  gate690(.a(s_20), .O(gate413inter3));
  inv1  gate691(.a(s_21), .O(gate413inter4));
  nand2 gate692(.a(gate413inter4), .b(gate413inter3), .O(gate413inter5));
  nor2  gate693(.a(gate413inter5), .b(gate413inter2), .O(gate413inter6));
  inv1  gate694(.a(G27), .O(gate413inter7));
  inv1  gate695(.a(G1114), .O(gate413inter8));
  nand2 gate696(.a(gate413inter8), .b(gate413inter7), .O(gate413inter9));
  nand2 gate697(.a(s_21), .b(gate413inter3), .O(gate413inter10));
  nor2  gate698(.a(gate413inter10), .b(gate413inter9), .O(gate413inter11));
  nor2  gate699(.a(gate413inter11), .b(gate413inter6), .O(gate413inter12));
  nand2 gate700(.a(gate413inter12), .b(gate413inter1), .O(G1210));
nand2 gate414( .a(G28), .b(G1117), .O(G1213) );
nand2 gate415( .a(G29), .b(G1120), .O(G1216) );

  xor2  gate2815(.a(G1123), .b(G30), .O(gate416inter0));
  nand2 gate2816(.a(gate416inter0), .b(s_324), .O(gate416inter1));
  and2  gate2817(.a(G1123), .b(G30), .O(gate416inter2));
  inv1  gate2818(.a(s_324), .O(gate416inter3));
  inv1  gate2819(.a(s_325), .O(gate416inter4));
  nand2 gate2820(.a(gate416inter4), .b(gate416inter3), .O(gate416inter5));
  nor2  gate2821(.a(gate416inter5), .b(gate416inter2), .O(gate416inter6));
  inv1  gate2822(.a(G30), .O(gate416inter7));
  inv1  gate2823(.a(G1123), .O(gate416inter8));
  nand2 gate2824(.a(gate416inter8), .b(gate416inter7), .O(gate416inter9));
  nand2 gate2825(.a(s_325), .b(gate416inter3), .O(gate416inter10));
  nor2  gate2826(.a(gate416inter10), .b(gate416inter9), .O(gate416inter11));
  nor2  gate2827(.a(gate416inter11), .b(gate416inter6), .O(gate416inter12));
  nand2 gate2828(.a(gate416inter12), .b(gate416inter1), .O(G1219));

  xor2  gate2409(.a(G1126), .b(G31), .O(gate417inter0));
  nand2 gate2410(.a(gate417inter0), .b(s_266), .O(gate417inter1));
  and2  gate2411(.a(G1126), .b(G31), .O(gate417inter2));
  inv1  gate2412(.a(s_266), .O(gate417inter3));
  inv1  gate2413(.a(s_267), .O(gate417inter4));
  nand2 gate2414(.a(gate417inter4), .b(gate417inter3), .O(gate417inter5));
  nor2  gate2415(.a(gate417inter5), .b(gate417inter2), .O(gate417inter6));
  inv1  gate2416(.a(G31), .O(gate417inter7));
  inv1  gate2417(.a(G1126), .O(gate417inter8));
  nand2 gate2418(.a(gate417inter8), .b(gate417inter7), .O(gate417inter9));
  nand2 gate2419(.a(s_267), .b(gate417inter3), .O(gate417inter10));
  nor2  gate2420(.a(gate417inter10), .b(gate417inter9), .O(gate417inter11));
  nor2  gate2421(.a(gate417inter11), .b(gate417inter6), .O(gate417inter12));
  nand2 gate2422(.a(gate417inter12), .b(gate417inter1), .O(G1222));

  xor2  gate1919(.a(G1129), .b(G32), .O(gate418inter0));
  nand2 gate1920(.a(gate418inter0), .b(s_196), .O(gate418inter1));
  and2  gate1921(.a(G1129), .b(G32), .O(gate418inter2));
  inv1  gate1922(.a(s_196), .O(gate418inter3));
  inv1  gate1923(.a(s_197), .O(gate418inter4));
  nand2 gate1924(.a(gate418inter4), .b(gate418inter3), .O(gate418inter5));
  nor2  gate1925(.a(gate418inter5), .b(gate418inter2), .O(gate418inter6));
  inv1  gate1926(.a(G32), .O(gate418inter7));
  inv1  gate1927(.a(G1129), .O(gate418inter8));
  nand2 gate1928(.a(gate418inter8), .b(gate418inter7), .O(gate418inter9));
  nand2 gate1929(.a(s_197), .b(gate418inter3), .O(gate418inter10));
  nor2  gate1930(.a(gate418inter10), .b(gate418inter9), .O(gate418inter11));
  nor2  gate1931(.a(gate418inter11), .b(gate418inter6), .O(gate418inter12));
  nand2 gate1932(.a(gate418inter12), .b(gate418inter1), .O(G1225));

  xor2  gate1611(.a(G1132), .b(G1), .O(gate419inter0));
  nand2 gate1612(.a(gate419inter0), .b(s_152), .O(gate419inter1));
  and2  gate1613(.a(G1132), .b(G1), .O(gate419inter2));
  inv1  gate1614(.a(s_152), .O(gate419inter3));
  inv1  gate1615(.a(s_153), .O(gate419inter4));
  nand2 gate1616(.a(gate419inter4), .b(gate419inter3), .O(gate419inter5));
  nor2  gate1617(.a(gate419inter5), .b(gate419inter2), .O(gate419inter6));
  inv1  gate1618(.a(G1), .O(gate419inter7));
  inv1  gate1619(.a(G1132), .O(gate419inter8));
  nand2 gate1620(.a(gate419inter8), .b(gate419inter7), .O(gate419inter9));
  nand2 gate1621(.a(s_153), .b(gate419inter3), .O(gate419inter10));
  nor2  gate1622(.a(gate419inter10), .b(gate419inter9), .O(gate419inter11));
  nor2  gate1623(.a(gate419inter11), .b(gate419inter6), .O(gate419inter12));
  nand2 gate1624(.a(gate419inter12), .b(gate419inter1), .O(G1228));

  xor2  gate1667(.a(G1132), .b(G1036), .O(gate420inter0));
  nand2 gate1668(.a(gate420inter0), .b(s_160), .O(gate420inter1));
  and2  gate1669(.a(G1132), .b(G1036), .O(gate420inter2));
  inv1  gate1670(.a(s_160), .O(gate420inter3));
  inv1  gate1671(.a(s_161), .O(gate420inter4));
  nand2 gate1672(.a(gate420inter4), .b(gate420inter3), .O(gate420inter5));
  nor2  gate1673(.a(gate420inter5), .b(gate420inter2), .O(gate420inter6));
  inv1  gate1674(.a(G1036), .O(gate420inter7));
  inv1  gate1675(.a(G1132), .O(gate420inter8));
  nand2 gate1676(.a(gate420inter8), .b(gate420inter7), .O(gate420inter9));
  nand2 gate1677(.a(s_161), .b(gate420inter3), .O(gate420inter10));
  nor2  gate1678(.a(gate420inter10), .b(gate420inter9), .O(gate420inter11));
  nor2  gate1679(.a(gate420inter11), .b(gate420inter6), .O(gate420inter12));
  nand2 gate1680(.a(gate420inter12), .b(gate420inter1), .O(G1229));
nand2 gate421( .a(G2), .b(G1135), .O(G1230) );

  xor2  gate1205(.a(G1135), .b(G1039), .O(gate422inter0));
  nand2 gate1206(.a(gate422inter0), .b(s_94), .O(gate422inter1));
  and2  gate1207(.a(G1135), .b(G1039), .O(gate422inter2));
  inv1  gate1208(.a(s_94), .O(gate422inter3));
  inv1  gate1209(.a(s_95), .O(gate422inter4));
  nand2 gate1210(.a(gate422inter4), .b(gate422inter3), .O(gate422inter5));
  nor2  gate1211(.a(gate422inter5), .b(gate422inter2), .O(gate422inter6));
  inv1  gate1212(.a(G1039), .O(gate422inter7));
  inv1  gate1213(.a(G1135), .O(gate422inter8));
  nand2 gate1214(.a(gate422inter8), .b(gate422inter7), .O(gate422inter9));
  nand2 gate1215(.a(s_95), .b(gate422inter3), .O(gate422inter10));
  nor2  gate1216(.a(gate422inter10), .b(gate422inter9), .O(gate422inter11));
  nor2  gate1217(.a(gate422inter11), .b(gate422inter6), .O(gate422inter12));
  nand2 gate1218(.a(gate422inter12), .b(gate422inter1), .O(G1231));
nand2 gate423( .a(G3), .b(G1138), .O(G1232) );
nand2 gate424( .a(G1042), .b(G1138), .O(G1233) );
nand2 gate425( .a(G4), .b(G1141), .O(G1234) );
nand2 gate426( .a(G1045), .b(G1141), .O(G1235) );
nand2 gate427( .a(G5), .b(G1144), .O(G1236) );

  xor2  gate1989(.a(G1144), .b(G1048), .O(gate428inter0));
  nand2 gate1990(.a(gate428inter0), .b(s_206), .O(gate428inter1));
  and2  gate1991(.a(G1144), .b(G1048), .O(gate428inter2));
  inv1  gate1992(.a(s_206), .O(gate428inter3));
  inv1  gate1993(.a(s_207), .O(gate428inter4));
  nand2 gate1994(.a(gate428inter4), .b(gate428inter3), .O(gate428inter5));
  nor2  gate1995(.a(gate428inter5), .b(gate428inter2), .O(gate428inter6));
  inv1  gate1996(.a(G1048), .O(gate428inter7));
  inv1  gate1997(.a(G1144), .O(gate428inter8));
  nand2 gate1998(.a(gate428inter8), .b(gate428inter7), .O(gate428inter9));
  nand2 gate1999(.a(s_207), .b(gate428inter3), .O(gate428inter10));
  nor2  gate2000(.a(gate428inter10), .b(gate428inter9), .O(gate428inter11));
  nor2  gate2001(.a(gate428inter11), .b(gate428inter6), .O(gate428inter12));
  nand2 gate2002(.a(gate428inter12), .b(gate428inter1), .O(G1237));

  xor2  gate1933(.a(G1147), .b(G6), .O(gate429inter0));
  nand2 gate1934(.a(gate429inter0), .b(s_198), .O(gate429inter1));
  and2  gate1935(.a(G1147), .b(G6), .O(gate429inter2));
  inv1  gate1936(.a(s_198), .O(gate429inter3));
  inv1  gate1937(.a(s_199), .O(gate429inter4));
  nand2 gate1938(.a(gate429inter4), .b(gate429inter3), .O(gate429inter5));
  nor2  gate1939(.a(gate429inter5), .b(gate429inter2), .O(gate429inter6));
  inv1  gate1940(.a(G6), .O(gate429inter7));
  inv1  gate1941(.a(G1147), .O(gate429inter8));
  nand2 gate1942(.a(gate429inter8), .b(gate429inter7), .O(gate429inter9));
  nand2 gate1943(.a(s_199), .b(gate429inter3), .O(gate429inter10));
  nor2  gate1944(.a(gate429inter10), .b(gate429inter9), .O(gate429inter11));
  nor2  gate1945(.a(gate429inter11), .b(gate429inter6), .O(gate429inter12));
  nand2 gate1946(.a(gate429inter12), .b(gate429inter1), .O(G1238));
nand2 gate430( .a(G1051), .b(G1147), .O(G1239) );

  xor2  gate1751(.a(G1150), .b(G7), .O(gate431inter0));
  nand2 gate1752(.a(gate431inter0), .b(s_172), .O(gate431inter1));
  and2  gate1753(.a(G1150), .b(G7), .O(gate431inter2));
  inv1  gate1754(.a(s_172), .O(gate431inter3));
  inv1  gate1755(.a(s_173), .O(gate431inter4));
  nand2 gate1756(.a(gate431inter4), .b(gate431inter3), .O(gate431inter5));
  nor2  gate1757(.a(gate431inter5), .b(gate431inter2), .O(gate431inter6));
  inv1  gate1758(.a(G7), .O(gate431inter7));
  inv1  gate1759(.a(G1150), .O(gate431inter8));
  nand2 gate1760(.a(gate431inter8), .b(gate431inter7), .O(gate431inter9));
  nand2 gate1761(.a(s_173), .b(gate431inter3), .O(gate431inter10));
  nor2  gate1762(.a(gate431inter10), .b(gate431inter9), .O(gate431inter11));
  nor2  gate1763(.a(gate431inter11), .b(gate431inter6), .O(gate431inter12));
  nand2 gate1764(.a(gate431inter12), .b(gate431inter1), .O(G1240));
nand2 gate432( .a(G1054), .b(G1150), .O(G1241) );

  xor2  gate1863(.a(G1153), .b(G8), .O(gate433inter0));
  nand2 gate1864(.a(gate433inter0), .b(s_188), .O(gate433inter1));
  and2  gate1865(.a(G1153), .b(G8), .O(gate433inter2));
  inv1  gate1866(.a(s_188), .O(gate433inter3));
  inv1  gate1867(.a(s_189), .O(gate433inter4));
  nand2 gate1868(.a(gate433inter4), .b(gate433inter3), .O(gate433inter5));
  nor2  gate1869(.a(gate433inter5), .b(gate433inter2), .O(gate433inter6));
  inv1  gate1870(.a(G8), .O(gate433inter7));
  inv1  gate1871(.a(G1153), .O(gate433inter8));
  nand2 gate1872(.a(gate433inter8), .b(gate433inter7), .O(gate433inter9));
  nand2 gate1873(.a(s_189), .b(gate433inter3), .O(gate433inter10));
  nor2  gate1874(.a(gate433inter10), .b(gate433inter9), .O(gate433inter11));
  nor2  gate1875(.a(gate433inter11), .b(gate433inter6), .O(gate433inter12));
  nand2 gate1876(.a(gate433inter12), .b(gate433inter1), .O(G1242));
nand2 gate434( .a(G1057), .b(G1153), .O(G1243) );
nand2 gate435( .a(G9), .b(G1156), .O(G1244) );

  xor2  gate1317(.a(G1156), .b(G1060), .O(gate436inter0));
  nand2 gate1318(.a(gate436inter0), .b(s_110), .O(gate436inter1));
  and2  gate1319(.a(G1156), .b(G1060), .O(gate436inter2));
  inv1  gate1320(.a(s_110), .O(gate436inter3));
  inv1  gate1321(.a(s_111), .O(gate436inter4));
  nand2 gate1322(.a(gate436inter4), .b(gate436inter3), .O(gate436inter5));
  nor2  gate1323(.a(gate436inter5), .b(gate436inter2), .O(gate436inter6));
  inv1  gate1324(.a(G1060), .O(gate436inter7));
  inv1  gate1325(.a(G1156), .O(gate436inter8));
  nand2 gate1326(.a(gate436inter8), .b(gate436inter7), .O(gate436inter9));
  nand2 gate1327(.a(s_111), .b(gate436inter3), .O(gate436inter10));
  nor2  gate1328(.a(gate436inter10), .b(gate436inter9), .O(gate436inter11));
  nor2  gate1329(.a(gate436inter11), .b(gate436inter6), .O(gate436inter12));
  nand2 gate1330(.a(gate436inter12), .b(gate436inter1), .O(G1245));

  xor2  gate2143(.a(G1159), .b(G10), .O(gate437inter0));
  nand2 gate2144(.a(gate437inter0), .b(s_228), .O(gate437inter1));
  and2  gate2145(.a(G1159), .b(G10), .O(gate437inter2));
  inv1  gate2146(.a(s_228), .O(gate437inter3));
  inv1  gate2147(.a(s_229), .O(gate437inter4));
  nand2 gate2148(.a(gate437inter4), .b(gate437inter3), .O(gate437inter5));
  nor2  gate2149(.a(gate437inter5), .b(gate437inter2), .O(gate437inter6));
  inv1  gate2150(.a(G10), .O(gate437inter7));
  inv1  gate2151(.a(G1159), .O(gate437inter8));
  nand2 gate2152(.a(gate437inter8), .b(gate437inter7), .O(gate437inter9));
  nand2 gate2153(.a(s_229), .b(gate437inter3), .O(gate437inter10));
  nor2  gate2154(.a(gate437inter10), .b(gate437inter9), .O(gate437inter11));
  nor2  gate2155(.a(gate437inter11), .b(gate437inter6), .O(gate437inter12));
  nand2 gate2156(.a(gate437inter12), .b(gate437inter1), .O(G1246));
nand2 gate438( .a(G1063), .b(G1159), .O(G1247) );
nand2 gate439( .a(G11), .b(G1162), .O(G1248) );

  xor2  gate1247(.a(G1162), .b(G1066), .O(gate440inter0));
  nand2 gate1248(.a(gate440inter0), .b(s_100), .O(gate440inter1));
  and2  gate1249(.a(G1162), .b(G1066), .O(gate440inter2));
  inv1  gate1250(.a(s_100), .O(gate440inter3));
  inv1  gate1251(.a(s_101), .O(gate440inter4));
  nand2 gate1252(.a(gate440inter4), .b(gate440inter3), .O(gate440inter5));
  nor2  gate1253(.a(gate440inter5), .b(gate440inter2), .O(gate440inter6));
  inv1  gate1254(.a(G1066), .O(gate440inter7));
  inv1  gate1255(.a(G1162), .O(gate440inter8));
  nand2 gate1256(.a(gate440inter8), .b(gate440inter7), .O(gate440inter9));
  nand2 gate1257(.a(s_101), .b(gate440inter3), .O(gate440inter10));
  nor2  gate1258(.a(gate440inter10), .b(gate440inter9), .O(gate440inter11));
  nor2  gate1259(.a(gate440inter11), .b(gate440inter6), .O(gate440inter12));
  nand2 gate1260(.a(gate440inter12), .b(gate440inter1), .O(G1249));
nand2 gate441( .a(G12), .b(G1165), .O(G1250) );
nand2 gate442( .a(G1069), .b(G1165), .O(G1251) );

  xor2  gate953(.a(G1168), .b(G13), .O(gate443inter0));
  nand2 gate954(.a(gate443inter0), .b(s_58), .O(gate443inter1));
  and2  gate955(.a(G1168), .b(G13), .O(gate443inter2));
  inv1  gate956(.a(s_58), .O(gate443inter3));
  inv1  gate957(.a(s_59), .O(gate443inter4));
  nand2 gate958(.a(gate443inter4), .b(gate443inter3), .O(gate443inter5));
  nor2  gate959(.a(gate443inter5), .b(gate443inter2), .O(gate443inter6));
  inv1  gate960(.a(G13), .O(gate443inter7));
  inv1  gate961(.a(G1168), .O(gate443inter8));
  nand2 gate962(.a(gate443inter8), .b(gate443inter7), .O(gate443inter9));
  nand2 gate963(.a(s_59), .b(gate443inter3), .O(gate443inter10));
  nor2  gate964(.a(gate443inter10), .b(gate443inter9), .O(gate443inter11));
  nor2  gate965(.a(gate443inter11), .b(gate443inter6), .O(gate443inter12));
  nand2 gate966(.a(gate443inter12), .b(gate443inter1), .O(G1252));

  xor2  gate2773(.a(G1168), .b(G1072), .O(gate444inter0));
  nand2 gate2774(.a(gate444inter0), .b(s_318), .O(gate444inter1));
  and2  gate2775(.a(G1168), .b(G1072), .O(gate444inter2));
  inv1  gate2776(.a(s_318), .O(gate444inter3));
  inv1  gate2777(.a(s_319), .O(gate444inter4));
  nand2 gate2778(.a(gate444inter4), .b(gate444inter3), .O(gate444inter5));
  nor2  gate2779(.a(gate444inter5), .b(gate444inter2), .O(gate444inter6));
  inv1  gate2780(.a(G1072), .O(gate444inter7));
  inv1  gate2781(.a(G1168), .O(gate444inter8));
  nand2 gate2782(.a(gate444inter8), .b(gate444inter7), .O(gate444inter9));
  nand2 gate2783(.a(s_319), .b(gate444inter3), .O(gate444inter10));
  nor2  gate2784(.a(gate444inter10), .b(gate444inter9), .O(gate444inter11));
  nor2  gate2785(.a(gate444inter11), .b(gate444inter6), .O(gate444inter12));
  nand2 gate2786(.a(gate444inter12), .b(gate444inter1), .O(G1253));

  xor2  gate2003(.a(G1171), .b(G14), .O(gate445inter0));
  nand2 gate2004(.a(gate445inter0), .b(s_208), .O(gate445inter1));
  and2  gate2005(.a(G1171), .b(G14), .O(gate445inter2));
  inv1  gate2006(.a(s_208), .O(gate445inter3));
  inv1  gate2007(.a(s_209), .O(gate445inter4));
  nand2 gate2008(.a(gate445inter4), .b(gate445inter3), .O(gate445inter5));
  nor2  gate2009(.a(gate445inter5), .b(gate445inter2), .O(gate445inter6));
  inv1  gate2010(.a(G14), .O(gate445inter7));
  inv1  gate2011(.a(G1171), .O(gate445inter8));
  nand2 gate2012(.a(gate445inter8), .b(gate445inter7), .O(gate445inter9));
  nand2 gate2013(.a(s_209), .b(gate445inter3), .O(gate445inter10));
  nor2  gate2014(.a(gate445inter10), .b(gate445inter9), .O(gate445inter11));
  nor2  gate2015(.a(gate445inter11), .b(gate445inter6), .O(gate445inter12));
  nand2 gate2016(.a(gate445inter12), .b(gate445inter1), .O(G1254));

  xor2  gate2465(.a(G1171), .b(G1075), .O(gate446inter0));
  nand2 gate2466(.a(gate446inter0), .b(s_274), .O(gate446inter1));
  and2  gate2467(.a(G1171), .b(G1075), .O(gate446inter2));
  inv1  gate2468(.a(s_274), .O(gate446inter3));
  inv1  gate2469(.a(s_275), .O(gate446inter4));
  nand2 gate2470(.a(gate446inter4), .b(gate446inter3), .O(gate446inter5));
  nor2  gate2471(.a(gate446inter5), .b(gate446inter2), .O(gate446inter6));
  inv1  gate2472(.a(G1075), .O(gate446inter7));
  inv1  gate2473(.a(G1171), .O(gate446inter8));
  nand2 gate2474(.a(gate446inter8), .b(gate446inter7), .O(gate446inter9));
  nand2 gate2475(.a(s_275), .b(gate446inter3), .O(gate446inter10));
  nor2  gate2476(.a(gate446inter10), .b(gate446inter9), .O(gate446inter11));
  nor2  gate2477(.a(gate446inter11), .b(gate446inter6), .O(gate446inter12));
  nand2 gate2478(.a(gate446inter12), .b(gate446inter1), .O(G1255));
nand2 gate447( .a(G15), .b(G1174), .O(G1256) );
nand2 gate448( .a(G1078), .b(G1174), .O(G1257) );
nand2 gate449( .a(G16), .b(G1177), .O(G1258) );

  xor2  gate2311(.a(G1177), .b(G1081), .O(gate450inter0));
  nand2 gate2312(.a(gate450inter0), .b(s_252), .O(gate450inter1));
  and2  gate2313(.a(G1177), .b(G1081), .O(gate450inter2));
  inv1  gate2314(.a(s_252), .O(gate450inter3));
  inv1  gate2315(.a(s_253), .O(gate450inter4));
  nand2 gate2316(.a(gate450inter4), .b(gate450inter3), .O(gate450inter5));
  nor2  gate2317(.a(gate450inter5), .b(gate450inter2), .O(gate450inter6));
  inv1  gate2318(.a(G1081), .O(gate450inter7));
  inv1  gate2319(.a(G1177), .O(gate450inter8));
  nand2 gate2320(.a(gate450inter8), .b(gate450inter7), .O(gate450inter9));
  nand2 gate2321(.a(s_253), .b(gate450inter3), .O(gate450inter10));
  nor2  gate2322(.a(gate450inter10), .b(gate450inter9), .O(gate450inter11));
  nor2  gate2323(.a(gate450inter11), .b(gate450inter6), .O(gate450inter12));
  nand2 gate2324(.a(gate450inter12), .b(gate450inter1), .O(G1259));
nand2 gate451( .a(G17), .b(G1180), .O(G1260) );
nand2 gate452( .a(G1084), .b(G1180), .O(G1261) );

  xor2  gate2941(.a(G1183), .b(G18), .O(gate453inter0));
  nand2 gate2942(.a(gate453inter0), .b(s_342), .O(gate453inter1));
  and2  gate2943(.a(G1183), .b(G18), .O(gate453inter2));
  inv1  gate2944(.a(s_342), .O(gate453inter3));
  inv1  gate2945(.a(s_343), .O(gate453inter4));
  nand2 gate2946(.a(gate453inter4), .b(gate453inter3), .O(gate453inter5));
  nor2  gate2947(.a(gate453inter5), .b(gate453inter2), .O(gate453inter6));
  inv1  gate2948(.a(G18), .O(gate453inter7));
  inv1  gate2949(.a(G1183), .O(gate453inter8));
  nand2 gate2950(.a(gate453inter8), .b(gate453inter7), .O(gate453inter9));
  nand2 gate2951(.a(s_343), .b(gate453inter3), .O(gate453inter10));
  nor2  gate2952(.a(gate453inter10), .b(gate453inter9), .O(gate453inter11));
  nor2  gate2953(.a(gate453inter11), .b(gate453inter6), .O(gate453inter12));
  nand2 gate2954(.a(gate453inter12), .b(gate453inter1), .O(G1262));

  xor2  gate2731(.a(G1183), .b(G1087), .O(gate454inter0));
  nand2 gate2732(.a(gate454inter0), .b(s_312), .O(gate454inter1));
  and2  gate2733(.a(G1183), .b(G1087), .O(gate454inter2));
  inv1  gate2734(.a(s_312), .O(gate454inter3));
  inv1  gate2735(.a(s_313), .O(gate454inter4));
  nand2 gate2736(.a(gate454inter4), .b(gate454inter3), .O(gate454inter5));
  nor2  gate2737(.a(gate454inter5), .b(gate454inter2), .O(gate454inter6));
  inv1  gate2738(.a(G1087), .O(gate454inter7));
  inv1  gate2739(.a(G1183), .O(gate454inter8));
  nand2 gate2740(.a(gate454inter8), .b(gate454inter7), .O(gate454inter9));
  nand2 gate2741(.a(s_313), .b(gate454inter3), .O(gate454inter10));
  nor2  gate2742(.a(gate454inter10), .b(gate454inter9), .O(gate454inter11));
  nor2  gate2743(.a(gate454inter11), .b(gate454inter6), .O(gate454inter12));
  nand2 gate2744(.a(gate454inter12), .b(gate454inter1), .O(G1263));

  xor2  gate2661(.a(G1186), .b(G19), .O(gate455inter0));
  nand2 gate2662(.a(gate455inter0), .b(s_302), .O(gate455inter1));
  and2  gate2663(.a(G1186), .b(G19), .O(gate455inter2));
  inv1  gate2664(.a(s_302), .O(gate455inter3));
  inv1  gate2665(.a(s_303), .O(gate455inter4));
  nand2 gate2666(.a(gate455inter4), .b(gate455inter3), .O(gate455inter5));
  nor2  gate2667(.a(gate455inter5), .b(gate455inter2), .O(gate455inter6));
  inv1  gate2668(.a(G19), .O(gate455inter7));
  inv1  gate2669(.a(G1186), .O(gate455inter8));
  nand2 gate2670(.a(gate455inter8), .b(gate455inter7), .O(gate455inter9));
  nand2 gate2671(.a(s_303), .b(gate455inter3), .O(gate455inter10));
  nor2  gate2672(.a(gate455inter10), .b(gate455inter9), .O(gate455inter11));
  nor2  gate2673(.a(gate455inter11), .b(gate455inter6), .O(gate455inter12));
  nand2 gate2674(.a(gate455inter12), .b(gate455inter1), .O(G1264));
nand2 gate456( .a(G1090), .b(G1186), .O(G1265) );

  xor2  gate743(.a(G1189), .b(G20), .O(gate457inter0));
  nand2 gate744(.a(gate457inter0), .b(s_28), .O(gate457inter1));
  and2  gate745(.a(G1189), .b(G20), .O(gate457inter2));
  inv1  gate746(.a(s_28), .O(gate457inter3));
  inv1  gate747(.a(s_29), .O(gate457inter4));
  nand2 gate748(.a(gate457inter4), .b(gate457inter3), .O(gate457inter5));
  nor2  gate749(.a(gate457inter5), .b(gate457inter2), .O(gate457inter6));
  inv1  gate750(.a(G20), .O(gate457inter7));
  inv1  gate751(.a(G1189), .O(gate457inter8));
  nand2 gate752(.a(gate457inter8), .b(gate457inter7), .O(gate457inter9));
  nand2 gate753(.a(s_29), .b(gate457inter3), .O(gate457inter10));
  nor2  gate754(.a(gate457inter10), .b(gate457inter9), .O(gate457inter11));
  nor2  gate755(.a(gate457inter11), .b(gate457inter6), .O(gate457inter12));
  nand2 gate756(.a(gate457inter12), .b(gate457inter1), .O(G1266));
nand2 gate458( .a(G1093), .b(G1189), .O(G1267) );

  xor2  gate1415(.a(G1192), .b(G21), .O(gate459inter0));
  nand2 gate1416(.a(gate459inter0), .b(s_124), .O(gate459inter1));
  and2  gate1417(.a(G1192), .b(G21), .O(gate459inter2));
  inv1  gate1418(.a(s_124), .O(gate459inter3));
  inv1  gate1419(.a(s_125), .O(gate459inter4));
  nand2 gate1420(.a(gate459inter4), .b(gate459inter3), .O(gate459inter5));
  nor2  gate1421(.a(gate459inter5), .b(gate459inter2), .O(gate459inter6));
  inv1  gate1422(.a(G21), .O(gate459inter7));
  inv1  gate1423(.a(G1192), .O(gate459inter8));
  nand2 gate1424(.a(gate459inter8), .b(gate459inter7), .O(gate459inter9));
  nand2 gate1425(.a(s_125), .b(gate459inter3), .O(gate459inter10));
  nor2  gate1426(.a(gate459inter10), .b(gate459inter9), .O(gate459inter11));
  nor2  gate1427(.a(gate459inter11), .b(gate459inter6), .O(gate459inter12));
  nand2 gate1428(.a(gate459inter12), .b(gate459inter1), .O(G1268));

  xor2  gate1303(.a(G1192), .b(G1096), .O(gate460inter0));
  nand2 gate1304(.a(gate460inter0), .b(s_108), .O(gate460inter1));
  and2  gate1305(.a(G1192), .b(G1096), .O(gate460inter2));
  inv1  gate1306(.a(s_108), .O(gate460inter3));
  inv1  gate1307(.a(s_109), .O(gate460inter4));
  nand2 gate1308(.a(gate460inter4), .b(gate460inter3), .O(gate460inter5));
  nor2  gate1309(.a(gate460inter5), .b(gate460inter2), .O(gate460inter6));
  inv1  gate1310(.a(G1096), .O(gate460inter7));
  inv1  gate1311(.a(G1192), .O(gate460inter8));
  nand2 gate1312(.a(gate460inter8), .b(gate460inter7), .O(gate460inter9));
  nand2 gate1313(.a(s_109), .b(gate460inter3), .O(gate460inter10));
  nor2  gate1314(.a(gate460inter10), .b(gate460inter9), .O(gate460inter11));
  nor2  gate1315(.a(gate460inter11), .b(gate460inter6), .O(gate460inter12));
  nand2 gate1316(.a(gate460inter12), .b(gate460inter1), .O(G1269));

  xor2  gate2353(.a(G1195), .b(G22), .O(gate461inter0));
  nand2 gate2354(.a(gate461inter0), .b(s_258), .O(gate461inter1));
  and2  gate2355(.a(G1195), .b(G22), .O(gate461inter2));
  inv1  gate2356(.a(s_258), .O(gate461inter3));
  inv1  gate2357(.a(s_259), .O(gate461inter4));
  nand2 gate2358(.a(gate461inter4), .b(gate461inter3), .O(gate461inter5));
  nor2  gate2359(.a(gate461inter5), .b(gate461inter2), .O(gate461inter6));
  inv1  gate2360(.a(G22), .O(gate461inter7));
  inv1  gate2361(.a(G1195), .O(gate461inter8));
  nand2 gate2362(.a(gate461inter8), .b(gate461inter7), .O(gate461inter9));
  nand2 gate2363(.a(s_259), .b(gate461inter3), .O(gate461inter10));
  nor2  gate2364(.a(gate461inter10), .b(gate461inter9), .O(gate461inter11));
  nor2  gate2365(.a(gate461inter11), .b(gate461inter6), .O(gate461inter12));
  nand2 gate2366(.a(gate461inter12), .b(gate461inter1), .O(G1270));
nand2 gate462( .a(G1099), .b(G1195), .O(G1271) );

  xor2  gate1639(.a(G1198), .b(G23), .O(gate463inter0));
  nand2 gate1640(.a(gate463inter0), .b(s_156), .O(gate463inter1));
  and2  gate1641(.a(G1198), .b(G23), .O(gate463inter2));
  inv1  gate1642(.a(s_156), .O(gate463inter3));
  inv1  gate1643(.a(s_157), .O(gate463inter4));
  nand2 gate1644(.a(gate463inter4), .b(gate463inter3), .O(gate463inter5));
  nor2  gate1645(.a(gate463inter5), .b(gate463inter2), .O(gate463inter6));
  inv1  gate1646(.a(G23), .O(gate463inter7));
  inv1  gate1647(.a(G1198), .O(gate463inter8));
  nand2 gate1648(.a(gate463inter8), .b(gate463inter7), .O(gate463inter9));
  nand2 gate1649(.a(s_157), .b(gate463inter3), .O(gate463inter10));
  nor2  gate1650(.a(gate463inter10), .b(gate463inter9), .O(gate463inter11));
  nor2  gate1651(.a(gate463inter11), .b(gate463inter6), .O(gate463inter12));
  nand2 gate1652(.a(gate463inter12), .b(gate463inter1), .O(G1272));
nand2 gate464( .a(G1102), .b(G1198), .O(G1273) );
nand2 gate465( .a(G24), .b(G1201), .O(G1274) );
nand2 gate466( .a(G1105), .b(G1201), .O(G1275) );

  xor2  gate2619(.a(G1204), .b(G25), .O(gate467inter0));
  nand2 gate2620(.a(gate467inter0), .b(s_296), .O(gate467inter1));
  and2  gate2621(.a(G1204), .b(G25), .O(gate467inter2));
  inv1  gate2622(.a(s_296), .O(gate467inter3));
  inv1  gate2623(.a(s_297), .O(gate467inter4));
  nand2 gate2624(.a(gate467inter4), .b(gate467inter3), .O(gate467inter5));
  nor2  gate2625(.a(gate467inter5), .b(gate467inter2), .O(gate467inter6));
  inv1  gate2626(.a(G25), .O(gate467inter7));
  inv1  gate2627(.a(G1204), .O(gate467inter8));
  nand2 gate2628(.a(gate467inter8), .b(gate467inter7), .O(gate467inter9));
  nand2 gate2629(.a(s_297), .b(gate467inter3), .O(gate467inter10));
  nor2  gate2630(.a(gate467inter10), .b(gate467inter9), .O(gate467inter11));
  nor2  gate2631(.a(gate467inter11), .b(gate467inter6), .O(gate467inter12));
  nand2 gate2632(.a(gate467inter12), .b(gate467inter1), .O(G1276));

  xor2  gate1709(.a(G1204), .b(G1108), .O(gate468inter0));
  nand2 gate1710(.a(gate468inter0), .b(s_166), .O(gate468inter1));
  and2  gate1711(.a(G1204), .b(G1108), .O(gate468inter2));
  inv1  gate1712(.a(s_166), .O(gate468inter3));
  inv1  gate1713(.a(s_167), .O(gate468inter4));
  nand2 gate1714(.a(gate468inter4), .b(gate468inter3), .O(gate468inter5));
  nor2  gate1715(.a(gate468inter5), .b(gate468inter2), .O(gate468inter6));
  inv1  gate1716(.a(G1108), .O(gate468inter7));
  inv1  gate1717(.a(G1204), .O(gate468inter8));
  nand2 gate1718(.a(gate468inter8), .b(gate468inter7), .O(gate468inter9));
  nand2 gate1719(.a(s_167), .b(gate468inter3), .O(gate468inter10));
  nor2  gate1720(.a(gate468inter10), .b(gate468inter9), .O(gate468inter11));
  nor2  gate1721(.a(gate468inter11), .b(gate468inter6), .O(gate468inter12));
  nand2 gate1722(.a(gate468inter12), .b(gate468inter1), .O(G1277));
nand2 gate469( .a(G26), .b(G1207), .O(G1278) );
nand2 gate470( .a(G1111), .b(G1207), .O(G1279) );

  xor2  gate1429(.a(G1210), .b(G27), .O(gate471inter0));
  nand2 gate1430(.a(gate471inter0), .b(s_126), .O(gate471inter1));
  and2  gate1431(.a(G1210), .b(G27), .O(gate471inter2));
  inv1  gate1432(.a(s_126), .O(gate471inter3));
  inv1  gate1433(.a(s_127), .O(gate471inter4));
  nand2 gate1434(.a(gate471inter4), .b(gate471inter3), .O(gate471inter5));
  nor2  gate1435(.a(gate471inter5), .b(gate471inter2), .O(gate471inter6));
  inv1  gate1436(.a(G27), .O(gate471inter7));
  inv1  gate1437(.a(G1210), .O(gate471inter8));
  nand2 gate1438(.a(gate471inter8), .b(gate471inter7), .O(gate471inter9));
  nand2 gate1439(.a(s_127), .b(gate471inter3), .O(gate471inter10));
  nor2  gate1440(.a(gate471inter10), .b(gate471inter9), .O(gate471inter11));
  nor2  gate1441(.a(gate471inter11), .b(gate471inter6), .O(gate471inter12));
  nand2 gate1442(.a(gate471inter12), .b(gate471inter1), .O(G1280));
nand2 gate472( .a(G1114), .b(G1210), .O(G1281) );
nand2 gate473( .a(G28), .b(G1213), .O(G1282) );
nand2 gate474( .a(G1117), .b(G1213), .O(G1283) );

  xor2  gate2213(.a(G1216), .b(G29), .O(gate475inter0));
  nand2 gate2214(.a(gate475inter0), .b(s_238), .O(gate475inter1));
  and2  gate2215(.a(G1216), .b(G29), .O(gate475inter2));
  inv1  gate2216(.a(s_238), .O(gate475inter3));
  inv1  gate2217(.a(s_239), .O(gate475inter4));
  nand2 gate2218(.a(gate475inter4), .b(gate475inter3), .O(gate475inter5));
  nor2  gate2219(.a(gate475inter5), .b(gate475inter2), .O(gate475inter6));
  inv1  gate2220(.a(G29), .O(gate475inter7));
  inv1  gate2221(.a(G1216), .O(gate475inter8));
  nand2 gate2222(.a(gate475inter8), .b(gate475inter7), .O(gate475inter9));
  nand2 gate2223(.a(s_239), .b(gate475inter3), .O(gate475inter10));
  nor2  gate2224(.a(gate475inter10), .b(gate475inter9), .O(gate475inter11));
  nor2  gate2225(.a(gate475inter11), .b(gate475inter6), .O(gate475inter12));
  nand2 gate2226(.a(gate475inter12), .b(gate475inter1), .O(G1284));

  xor2  gate2479(.a(G1216), .b(G1120), .O(gate476inter0));
  nand2 gate2480(.a(gate476inter0), .b(s_276), .O(gate476inter1));
  and2  gate2481(.a(G1216), .b(G1120), .O(gate476inter2));
  inv1  gate2482(.a(s_276), .O(gate476inter3));
  inv1  gate2483(.a(s_277), .O(gate476inter4));
  nand2 gate2484(.a(gate476inter4), .b(gate476inter3), .O(gate476inter5));
  nor2  gate2485(.a(gate476inter5), .b(gate476inter2), .O(gate476inter6));
  inv1  gate2486(.a(G1120), .O(gate476inter7));
  inv1  gate2487(.a(G1216), .O(gate476inter8));
  nand2 gate2488(.a(gate476inter8), .b(gate476inter7), .O(gate476inter9));
  nand2 gate2489(.a(s_277), .b(gate476inter3), .O(gate476inter10));
  nor2  gate2490(.a(gate476inter10), .b(gate476inter9), .O(gate476inter11));
  nor2  gate2491(.a(gate476inter11), .b(gate476inter6), .O(gate476inter12));
  nand2 gate2492(.a(gate476inter12), .b(gate476inter1), .O(G1285));
nand2 gate477( .a(G30), .b(G1219), .O(G1286) );

  xor2  gate1359(.a(G1219), .b(G1123), .O(gate478inter0));
  nand2 gate1360(.a(gate478inter0), .b(s_116), .O(gate478inter1));
  and2  gate1361(.a(G1219), .b(G1123), .O(gate478inter2));
  inv1  gate1362(.a(s_116), .O(gate478inter3));
  inv1  gate1363(.a(s_117), .O(gate478inter4));
  nand2 gate1364(.a(gate478inter4), .b(gate478inter3), .O(gate478inter5));
  nor2  gate1365(.a(gate478inter5), .b(gate478inter2), .O(gate478inter6));
  inv1  gate1366(.a(G1123), .O(gate478inter7));
  inv1  gate1367(.a(G1219), .O(gate478inter8));
  nand2 gate1368(.a(gate478inter8), .b(gate478inter7), .O(gate478inter9));
  nand2 gate1369(.a(s_117), .b(gate478inter3), .O(gate478inter10));
  nor2  gate1370(.a(gate478inter10), .b(gate478inter9), .O(gate478inter11));
  nor2  gate1371(.a(gate478inter11), .b(gate478inter6), .O(gate478inter12));
  nand2 gate1372(.a(gate478inter12), .b(gate478inter1), .O(G1287));
nand2 gate479( .a(G31), .b(G1222), .O(G1288) );
nand2 gate480( .a(G1126), .b(G1222), .O(G1289) );
nand2 gate481( .a(G32), .b(G1225), .O(G1290) );
nand2 gate482( .a(G1129), .b(G1225), .O(G1291) );
nand2 gate483( .a(G1228), .b(G1229), .O(G1292) );

  xor2  gate2577(.a(G1231), .b(G1230), .O(gate484inter0));
  nand2 gate2578(.a(gate484inter0), .b(s_290), .O(gate484inter1));
  and2  gate2579(.a(G1231), .b(G1230), .O(gate484inter2));
  inv1  gate2580(.a(s_290), .O(gate484inter3));
  inv1  gate2581(.a(s_291), .O(gate484inter4));
  nand2 gate2582(.a(gate484inter4), .b(gate484inter3), .O(gate484inter5));
  nor2  gate2583(.a(gate484inter5), .b(gate484inter2), .O(gate484inter6));
  inv1  gate2584(.a(G1230), .O(gate484inter7));
  inv1  gate2585(.a(G1231), .O(gate484inter8));
  nand2 gate2586(.a(gate484inter8), .b(gate484inter7), .O(gate484inter9));
  nand2 gate2587(.a(s_291), .b(gate484inter3), .O(gate484inter10));
  nor2  gate2588(.a(gate484inter10), .b(gate484inter9), .O(gate484inter11));
  nor2  gate2589(.a(gate484inter11), .b(gate484inter6), .O(gate484inter12));
  nand2 gate2590(.a(gate484inter12), .b(gate484inter1), .O(G1293));
nand2 gate485( .a(G1232), .b(G1233), .O(G1294) );
nand2 gate486( .a(G1234), .b(G1235), .O(G1295) );
nand2 gate487( .a(G1236), .b(G1237), .O(G1296) );
nand2 gate488( .a(G1238), .b(G1239), .O(G1297) );
nand2 gate489( .a(G1240), .b(G1241), .O(G1298) );

  xor2  gate1051(.a(G1243), .b(G1242), .O(gate490inter0));
  nand2 gate1052(.a(gate490inter0), .b(s_72), .O(gate490inter1));
  and2  gate1053(.a(G1243), .b(G1242), .O(gate490inter2));
  inv1  gate1054(.a(s_72), .O(gate490inter3));
  inv1  gate1055(.a(s_73), .O(gate490inter4));
  nand2 gate1056(.a(gate490inter4), .b(gate490inter3), .O(gate490inter5));
  nor2  gate1057(.a(gate490inter5), .b(gate490inter2), .O(gate490inter6));
  inv1  gate1058(.a(G1242), .O(gate490inter7));
  inv1  gate1059(.a(G1243), .O(gate490inter8));
  nand2 gate1060(.a(gate490inter8), .b(gate490inter7), .O(gate490inter9));
  nand2 gate1061(.a(s_73), .b(gate490inter3), .O(gate490inter10));
  nor2  gate1062(.a(gate490inter10), .b(gate490inter9), .O(gate490inter11));
  nor2  gate1063(.a(gate490inter11), .b(gate490inter6), .O(gate490inter12));
  nand2 gate1064(.a(gate490inter12), .b(gate490inter1), .O(G1299));
nand2 gate491( .a(G1244), .b(G1245), .O(G1300) );

  xor2  gate1807(.a(G1247), .b(G1246), .O(gate492inter0));
  nand2 gate1808(.a(gate492inter0), .b(s_180), .O(gate492inter1));
  and2  gate1809(.a(G1247), .b(G1246), .O(gate492inter2));
  inv1  gate1810(.a(s_180), .O(gate492inter3));
  inv1  gate1811(.a(s_181), .O(gate492inter4));
  nand2 gate1812(.a(gate492inter4), .b(gate492inter3), .O(gate492inter5));
  nor2  gate1813(.a(gate492inter5), .b(gate492inter2), .O(gate492inter6));
  inv1  gate1814(.a(G1246), .O(gate492inter7));
  inv1  gate1815(.a(G1247), .O(gate492inter8));
  nand2 gate1816(.a(gate492inter8), .b(gate492inter7), .O(gate492inter9));
  nand2 gate1817(.a(s_181), .b(gate492inter3), .O(gate492inter10));
  nor2  gate1818(.a(gate492inter10), .b(gate492inter9), .O(gate492inter11));
  nor2  gate1819(.a(gate492inter11), .b(gate492inter6), .O(gate492inter12));
  nand2 gate1820(.a(gate492inter12), .b(gate492inter1), .O(G1301));
nand2 gate493( .a(G1248), .b(G1249), .O(G1302) );

  xor2  gate2675(.a(G1251), .b(G1250), .O(gate494inter0));
  nand2 gate2676(.a(gate494inter0), .b(s_304), .O(gate494inter1));
  and2  gate2677(.a(G1251), .b(G1250), .O(gate494inter2));
  inv1  gate2678(.a(s_304), .O(gate494inter3));
  inv1  gate2679(.a(s_305), .O(gate494inter4));
  nand2 gate2680(.a(gate494inter4), .b(gate494inter3), .O(gate494inter5));
  nor2  gate2681(.a(gate494inter5), .b(gate494inter2), .O(gate494inter6));
  inv1  gate2682(.a(G1250), .O(gate494inter7));
  inv1  gate2683(.a(G1251), .O(gate494inter8));
  nand2 gate2684(.a(gate494inter8), .b(gate494inter7), .O(gate494inter9));
  nand2 gate2685(.a(s_305), .b(gate494inter3), .O(gate494inter10));
  nor2  gate2686(.a(gate494inter10), .b(gate494inter9), .O(gate494inter11));
  nor2  gate2687(.a(gate494inter11), .b(gate494inter6), .O(gate494inter12));
  nand2 gate2688(.a(gate494inter12), .b(gate494inter1), .O(G1303));
nand2 gate495( .a(G1252), .b(G1253), .O(G1304) );

  xor2  gate2969(.a(G1255), .b(G1254), .O(gate496inter0));
  nand2 gate2970(.a(gate496inter0), .b(s_346), .O(gate496inter1));
  and2  gate2971(.a(G1255), .b(G1254), .O(gate496inter2));
  inv1  gate2972(.a(s_346), .O(gate496inter3));
  inv1  gate2973(.a(s_347), .O(gate496inter4));
  nand2 gate2974(.a(gate496inter4), .b(gate496inter3), .O(gate496inter5));
  nor2  gate2975(.a(gate496inter5), .b(gate496inter2), .O(gate496inter6));
  inv1  gate2976(.a(G1254), .O(gate496inter7));
  inv1  gate2977(.a(G1255), .O(gate496inter8));
  nand2 gate2978(.a(gate496inter8), .b(gate496inter7), .O(gate496inter9));
  nand2 gate2979(.a(s_347), .b(gate496inter3), .O(gate496inter10));
  nor2  gate2980(.a(gate496inter10), .b(gate496inter9), .O(gate496inter11));
  nor2  gate2981(.a(gate496inter11), .b(gate496inter6), .O(gate496inter12));
  nand2 gate2982(.a(gate496inter12), .b(gate496inter1), .O(G1305));
nand2 gate497( .a(G1256), .b(G1257), .O(G1306) );

  xor2  gate2255(.a(G1259), .b(G1258), .O(gate498inter0));
  nand2 gate2256(.a(gate498inter0), .b(s_244), .O(gate498inter1));
  and2  gate2257(.a(G1259), .b(G1258), .O(gate498inter2));
  inv1  gate2258(.a(s_244), .O(gate498inter3));
  inv1  gate2259(.a(s_245), .O(gate498inter4));
  nand2 gate2260(.a(gate498inter4), .b(gate498inter3), .O(gate498inter5));
  nor2  gate2261(.a(gate498inter5), .b(gate498inter2), .O(gate498inter6));
  inv1  gate2262(.a(G1258), .O(gate498inter7));
  inv1  gate2263(.a(G1259), .O(gate498inter8));
  nand2 gate2264(.a(gate498inter8), .b(gate498inter7), .O(gate498inter9));
  nand2 gate2265(.a(s_245), .b(gate498inter3), .O(gate498inter10));
  nor2  gate2266(.a(gate498inter10), .b(gate498inter9), .O(gate498inter11));
  nor2  gate2267(.a(gate498inter11), .b(gate498inter6), .O(gate498inter12));
  nand2 gate2268(.a(gate498inter12), .b(gate498inter1), .O(G1307));

  xor2  gate1093(.a(G1261), .b(G1260), .O(gate499inter0));
  nand2 gate1094(.a(gate499inter0), .b(s_78), .O(gate499inter1));
  and2  gate1095(.a(G1261), .b(G1260), .O(gate499inter2));
  inv1  gate1096(.a(s_78), .O(gate499inter3));
  inv1  gate1097(.a(s_79), .O(gate499inter4));
  nand2 gate1098(.a(gate499inter4), .b(gate499inter3), .O(gate499inter5));
  nor2  gate1099(.a(gate499inter5), .b(gate499inter2), .O(gate499inter6));
  inv1  gate1100(.a(G1260), .O(gate499inter7));
  inv1  gate1101(.a(G1261), .O(gate499inter8));
  nand2 gate1102(.a(gate499inter8), .b(gate499inter7), .O(gate499inter9));
  nand2 gate1103(.a(s_79), .b(gate499inter3), .O(gate499inter10));
  nor2  gate1104(.a(gate499inter10), .b(gate499inter9), .O(gate499inter11));
  nor2  gate1105(.a(gate499inter11), .b(gate499inter6), .O(gate499inter12));
  nand2 gate1106(.a(gate499inter12), .b(gate499inter1), .O(G1308));
nand2 gate500( .a(G1262), .b(G1263), .O(G1309) );
nand2 gate501( .a(G1264), .b(G1265), .O(G1310) );

  xor2  gate2423(.a(G1267), .b(G1266), .O(gate502inter0));
  nand2 gate2424(.a(gate502inter0), .b(s_268), .O(gate502inter1));
  and2  gate2425(.a(G1267), .b(G1266), .O(gate502inter2));
  inv1  gate2426(.a(s_268), .O(gate502inter3));
  inv1  gate2427(.a(s_269), .O(gate502inter4));
  nand2 gate2428(.a(gate502inter4), .b(gate502inter3), .O(gate502inter5));
  nor2  gate2429(.a(gate502inter5), .b(gate502inter2), .O(gate502inter6));
  inv1  gate2430(.a(G1266), .O(gate502inter7));
  inv1  gate2431(.a(G1267), .O(gate502inter8));
  nand2 gate2432(.a(gate502inter8), .b(gate502inter7), .O(gate502inter9));
  nand2 gate2433(.a(s_269), .b(gate502inter3), .O(gate502inter10));
  nor2  gate2434(.a(gate502inter10), .b(gate502inter9), .O(gate502inter11));
  nor2  gate2435(.a(gate502inter11), .b(gate502inter6), .O(gate502inter12));
  nand2 gate2436(.a(gate502inter12), .b(gate502inter1), .O(G1311));
nand2 gate503( .a(G1268), .b(G1269), .O(G1312) );

  xor2  gate1891(.a(G1271), .b(G1270), .O(gate504inter0));
  nand2 gate1892(.a(gate504inter0), .b(s_192), .O(gate504inter1));
  and2  gate1893(.a(G1271), .b(G1270), .O(gate504inter2));
  inv1  gate1894(.a(s_192), .O(gate504inter3));
  inv1  gate1895(.a(s_193), .O(gate504inter4));
  nand2 gate1896(.a(gate504inter4), .b(gate504inter3), .O(gate504inter5));
  nor2  gate1897(.a(gate504inter5), .b(gate504inter2), .O(gate504inter6));
  inv1  gate1898(.a(G1270), .O(gate504inter7));
  inv1  gate1899(.a(G1271), .O(gate504inter8));
  nand2 gate1900(.a(gate504inter8), .b(gate504inter7), .O(gate504inter9));
  nand2 gate1901(.a(s_193), .b(gate504inter3), .O(gate504inter10));
  nor2  gate1902(.a(gate504inter10), .b(gate504inter9), .O(gate504inter11));
  nor2  gate1903(.a(gate504inter11), .b(gate504inter6), .O(gate504inter12));
  nand2 gate1904(.a(gate504inter12), .b(gate504inter1), .O(G1313));

  xor2  gate1373(.a(G1273), .b(G1272), .O(gate505inter0));
  nand2 gate1374(.a(gate505inter0), .b(s_118), .O(gate505inter1));
  and2  gate1375(.a(G1273), .b(G1272), .O(gate505inter2));
  inv1  gate1376(.a(s_118), .O(gate505inter3));
  inv1  gate1377(.a(s_119), .O(gate505inter4));
  nand2 gate1378(.a(gate505inter4), .b(gate505inter3), .O(gate505inter5));
  nor2  gate1379(.a(gate505inter5), .b(gate505inter2), .O(gate505inter6));
  inv1  gate1380(.a(G1272), .O(gate505inter7));
  inv1  gate1381(.a(G1273), .O(gate505inter8));
  nand2 gate1382(.a(gate505inter8), .b(gate505inter7), .O(gate505inter9));
  nand2 gate1383(.a(s_119), .b(gate505inter3), .O(gate505inter10));
  nor2  gate1384(.a(gate505inter10), .b(gate505inter9), .O(gate505inter11));
  nor2  gate1385(.a(gate505inter11), .b(gate505inter6), .O(gate505inter12));
  nand2 gate1386(.a(gate505inter12), .b(gate505inter1), .O(G1314));
nand2 gate506( .a(G1274), .b(G1275), .O(G1315) );
nand2 gate507( .a(G1276), .b(G1277), .O(G1316) );
nand2 gate508( .a(G1278), .b(G1279), .O(G1317) );

  xor2  gate2871(.a(G1281), .b(G1280), .O(gate509inter0));
  nand2 gate2872(.a(gate509inter0), .b(s_332), .O(gate509inter1));
  and2  gate2873(.a(G1281), .b(G1280), .O(gate509inter2));
  inv1  gate2874(.a(s_332), .O(gate509inter3));
  inv1  gate2875(.a(s_333), .O(gate509inter4));
  nand2 gate2876(.a(gate509inter4), .b(gate509inter3), .O(gate509inter5));
  nor2  gate2877(.a(gate509inter5), .b(gate509inter2), .O(gate509inter6));
  inv1  gate2878(.a(G1280), .O(gate509inter7));
  inv1  gate2879(.a(G1281), .O(gate509inter8));
  nand2 gate2880(.a(gate509inter8), .b(gate509inter7), .O(gate509inter9));
  nand2 gate2881(.a(s_333), .b(gate509inter3), .O(gate509inter10));
  nor2  gate2882(.a(gate509inter10), .b(gate509inter9), .O(gate509inter11));
  nor2  gate2883(.a(gate509inter11), .b(gate509inter6), .O(gate509inter12));
  nand2 gate2884(.a(gate509inter12), .b(gate509inter1), .O(G1318));

  xor2  gate2703(.a(G1283), .b(G1282), .O(gate510inter0));
  nand2 gate2704(.a(gate510inter0), .b(s_308), .O(gate510inter1));
  and2  gate2705(.a(G1283), .b(G1282), .O(gate510inter2));
  inv1  gate2706(.a(s_308), .O(gate510inter3));
  inv1  gate2707(.a(s_309), .O(gate510inter4));
  nand2 gate2708(.a(gate510inter4), .b(gate510inter3), .O(gate510inter5));
  nor2  gate2709(.a(gate510inter5), .b(gate510inter2), .O(gate510inter6));
  inv1  gate2710(.a(G1282), .O(gate510inter7));
  inv1  gate2711(.a(G1283), .O(gate510inter8));
  nand2 gate2712(.a(gate510inter8), .b(gate510inter7), .O(gate510inter9));
  nand2 gate2713(.a(s_309), .b(gate510inter3), .O(gate510inter10));
  nor2  gate2714(.a(gate510inter10), .b(gate510inter9), .O(gate510inter11));
  nor2  gate2715(.a(gate510inter11), .b(gate510inter6), .O(gate510inter12));
  nand2 gate2716(.a(gate510inter12), .b(gate510inter1), .O(G1319));
nand2 gate511( .a(G1284), .b(G1285), .O(G1320) );

  xor2  gate2157(.a(G1287), .b(G1286), .O(gate512inter0));
  nand2 gate2158(.a(gate512inter0), .b(s_230), .O(gate512inter1));
  and2  gate2159(.a(G1287), .b(G1286), .O(gate512inter2));
  inv1  gate2160(.a(s_230), .O(gate512inter3));
  inv1  gate2161(.a(s_231), .O(gate512inter4));
  nand2 gate2162(.a(gate512inter4), .b(gate512inter3), .O(gate512inter5));
  nor2  gate2163(.a(gate512inter5), .b(gate512inter2), .O(gate512inter6));
  inv1  gate2164(.a(G1286), .O(gate512inter7));
  inv1  gate2165(.a(G1287), .O(gate512inter8));
  nand2 gate2166(.a(gate512inter8), .b(gate512inter7), .O(gate512inter9));
  nand2 gate2167(.a(s_231), .b(gate512inter3), .O(gate512inter10));
  nor2  gate2168(.a(gate512inter10), .b(gate512inter9), .O(gate512inter11));
  nor2  gate2169(.a(gate512inter11), .b(gate512inter6), .O(gate512inter12));
  nand2 gate2170(.a(gate512inter12), .b(gate512inter1), .O(G1321));
nand2 gate513( .a(G1288), .b(G1289), .O(G1322) );

  xor2  gate673(.a(G1291), .b(G1290), .O(gate514inter0));
  nand2 gate674(.a(gate514inter0), .b(s_18), .O(gate514inter1));
  and2  gate675(.a(G1291), .b(G1290), .O(gate514inter2));
  inv1  gate676(.a(s_18), .O(gate514inter3));
  inv1  gate677(.a(s_19), .O(gate514inter4));
  nand2 gate678(.a(gate514inter4), .b(gate514inter3), .O(gate514inter5));
  nor2  gate679(.a(gate514inter5), .b(gate514inter2), .O(gate514inter6));
  inv1  gate680(.a(G1290), .O(gate514inter7));
  inv1  gate681(.a(G1291), .O(gate514inter8));
  nand2 gate682(.a(gate514inter8), .b(gate514inter7), .O(gate514inter9));
  nand2 gate683(.a(s_19), .b(gate514inter3), .O(gate514inter10));
  nor2  gate684(.a(gate514inter10), .b(gate514inter9), .O(gate514inter11));
  nor2  gate685(.a(gate514inter11), .b(gate514inter6), .O(gate514inter12));
  nand2 gate686(.a(gate514inter12), .b(gate514inter1), .O(G1323));
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule