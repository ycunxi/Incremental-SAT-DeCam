module c1908 (N1,N4,N7,N10,N13,N16,N19,N22,N25,N28,
              N31,N34,N37,N40,N43,N46,N49,N53,N56,N60,
              N63,N66,N69,N72,N76,N79,N82,N85,N88,N91,
              N94,N99,N104,N2753,N2754,N2755,N2756,N2762,N2767,N2768,
              N2779,N2780,N2781,N2782,N2783,N2784,N2785,N2786,N2787,N2811,
              N2886,N2887,N2888,N2889,N2890,N2891,N2892,N2899);
input N1,N4,N7,N10,N13,N16,N19,N22,N25,N28,
      N31,N34,N37,N40,N43,N46,N49,N53,N56,N60,
      N63,N66,N69,N72,N76,N79,N82,N85,N88,N91,
      N94,N99,N104;
  input s_0, s_1, s_2, s_3, s_4, s_5, s_6, s_7, s_8, s_9, s_10, s_11, s_12, s_13, s_14, s_15, s_16, s_17, s_18, s_19, s_20, s_21, s_22, s_23, s_24, s_25, s_26, s_27, s_28, s_29, s_30, s_31, s_32, s_33, s_34, s_35, s_36, s_37, s_38, s_39, s_40, s_41, s_42, s_43, s_44, s_45, s_46, s_47, s_48, s_49, s_50, s_51, s_52, s_53, s_54, s_55, s_56, s_57, s_58, s_59, s_60, s_61, s_62, s_63, s_64, s_65, s_66, s_67, s_68, s_69, s_70, s_71, s_72, s_73, s_74, s_75, s_76, s_77, s_78, s_79, s_80, s_81, s_82, s_83, s_84, s_85, s_86, s_87, s_88, s_89, s_90, s_91, s_92, s_93, s_94, s_95, s_96, s_97, s_98, s_99, s_100, s_101, s_102, s_103, s_104, s_105, s_106, s_107, s_108, s_109, s_110, s_111, s_112, s_113, s_114, s_115, s_116, s_117, s_118, s_119, s_120, s_121, s_122, s_123, s_124, s_125, s_126, s_127, s_128, s_129, s_130, s_131;
output N2753,N2754,N2755,N2756,N2762,N2767,N2768,N2779,N2780,N2781,
       N2782,N2783,N2784,N2785,N2786,N2787,N2811,N2886,N2887,N2888,
       N2889,N2890,N2891,N2892,N2899;
wire N190,N194,N197,N201,N206,N209,N212,N216,N220,N225,
     N229,N232,N235,N239,N243,N247,N251,N252,N253,N256,
     N257,N260,N263,N266,N269,N272,N275,N276,N277,N280,
     N283,N290,N297,N300,N303,N306,N313,N316,N319,N326,
     N331,N338,N343,N346,N349,N352,N355,N358,N361,N364,
     N367,N370,N373,N376,N379,N382,N385,N388,N534,N535,
     N536,N537,N538,N539,N540,N541,N542,N543,N544,N545,
     N546,N547,N548,N549,N550,N551,N552,N553,N554,N555,
     N556,N559,N562,N565,N568,N571,N574,N577,N580,N583,
     N586,N589,N592,N595,N598,N601,N602,N603,N608,N612,
     N616,N619,N622,N625,N628,N631,N634,N637,N640,N643,
     N646,N649,N652,N655,N658,N661,N664,N667,N670,N673,
     N676,N679,N682,N685,N688,N691,N694,N697,N700,N703,
     N706,N709,N712,N715,N718,N721,N724,N727,N730,N733,
     N736,N739,N742,N745,N748,N751,N886,N887,N888,N889,
     N890,N891,N892,N893,N894,N895,N896,N897,N898,N899,
     N903,N907,N910,N913,N914,N915,N916,N917,N918,N919,
     N920,N921,N922,N923,N926,N935,N938,N939,N942,N943,
     N946,N947,N950,N951,N954,N955,N958,N959,N962,N965,
     N968,N969,N972,N973,N976,N977,N980,N981,N984,N985,
     N988,N989,N990,N991,N992,N993,N994,N997,N998,N1001,
     N1002,N1003,N1004,N1005,N1006,N1007,N1008,N1009,N1010,N1013,
     N1016,N1019,N1022,N1025,N1028,N1031,N1034,N1037,N1040,N1043,
     N1046,N1049,N1054,N1055,N1063,N1064,N1067,N1068,N1119,N1120,
     N1121,N1122,N1128,N1129,N1130,N1131,N1132,N1133,N1148,N1149,
     N1150,N1151,N1152,N1153,N1154,N1155,N1156,N1157,N1158,N1159,
     N1160,N1161,N1162,N1163,N1164,N1167,N1168,N1171,N1188,N1205,
     N1206,N1207,N1208,N1209,N1210,N1211,N1212,N1213,N1214,N1215,
     N1216,N1217,N1218,N1219,N1220,N1221,N1222,N1223,N1224,N1225,
     N1226,N1227,N1228,N1229,N1230,N1231,N1232,N1235,N1238,N1239,
     N1240,N1241,N1242,N1243,N1246,N1249,N1252,N1255,N1258,N1261,
     N1264,N1267,N1309,N1310,N1311,N1312,N1313,N1314,N1315,N1316,
     N1317,N1318,N1319,N1322,N1327,N1328,N1334,N1344,N1345,N1346,
     N1348,N1349,N1350,N1351,N1352,N1355,N1358,N1361,N1364,N1367,
     N1370,N1373,N1376,N1379,N1383,N1386,N1387,N1388,N1389,N1390,
     N1393,N1396,N1397,N1398,N1399,N1409,N1412,N1413,N1416,N1419,
     N1433,N1434,N1438,N1439,N1440,N1443,N1444,N1445,N1446,N1447,
     N1448,N1451,N1452,N1453,N1454,N1455,N1456,N1457,N1458,N1459,
     N1460,N1461,N1462,N1463,N1464,N1468,N1469,N1470,N1471,N1472,
     N1475,N1476,N1478,N1481,N1484,N1487,N1488,N1489,N1490,N1491,
     N1492,N1493,N1494,N1495,N1496,N1498,N1499,N1500,N1501,N1504,
     N1510,N1513,N1514,N1517,N1520,N1521,N1522,N1526,N1527,N1528,
     N1529,N1530,N1531,N1532,N1534,N1537,N1540,N1546,N1554,N1557,
     N1561,N1567,N1568,N1569,N1571,N1576,N1588,N1591,N1593,N1594,
     N1595,N1596,N1600,N1603,N1606,N1609,N1612,N1615,N1620,N1623,
     N1635,N1636,N1638,N1639,N1640,N1643,N1647,N1651,N1658,N1661,
     N1664,N1671,N1672,N1675,N1677,N1678,N1679,N1680,N1681,N1682,
     N1683,N1685,N1688,N1697,N1701,N1706,N1707,N1708,N1709,N1710,
     N1711,N1712,N1713,N1714,N1717,N1720,N1721,N1723,N1727,N1728,
     N1730,N1731,N1734,N1740,N1741,N1742,N1746,N1747,N1748,N1751,
     N1759,N1761,N1762,N1763,N1764,N1768,N1769,N1772,N1773,N1774,
     N1777,N1783,N1784,N1785,N1786,N1787,N1788,N1791,N1792,N1795,
     N1796,N1798,N1801,N1802,N1807,N1808,N1809,N1810,N1812,N1815,
     N1818,N1821,N1822,N1823,N1824,N1825,N1826,N1827,N1830,N1837,
     N1838,N1841,N1848,N1849,N1850,N1852,N1855,N1856,N1857,N1858,
     N1864,N1865,N1866,N1869,N1872,N1875,N1878,N1879,N1882,N1883,
     N1884,N1885,N1889,N1895,N1896,N1897,N1898,N1902,N1910,N1911,
     N1912,N1913,N1915,N1919,N1920,N1921,N1922,N1923,N1924,N1927,
     N1930,N1933,N1936,N1937,N1938,N1941,N1942,N1944,N1947,N1950,
     N1953,N1958,N1961,N1965,N1968,N1975,N1976,N1977,N1978,N1979,
     N1980,N1985,N1987,N1999,N2000,N2002,N2003,N2004,N2005,N2006,
     N2007,N2008,N2009,N2012,N2013,N2014,N2015,N2016,N2018,N2019,
     N2020,N2021,N2022,N2023,N2024,N2025,N2026,N2027,N2030,N2033,
     N2036,N2037,N2038,N2039,N2040,N2041,N2042,N2047,N2052,N2055,
     N2060,N2061,N2062,N2067,N2068,N2071,N2076,N2077,N2078,N2081,
     N2086,N2089,N2104,N2119,N2129,N2143,N2148,N2151,N2196,N2199,
     N2202,N2205,N2214,N2215,N2216,N2217,N2222,N2223,N2224,N2225,
     N2226,N2227,N2228,N2229,N2230,N2231,N2232,N2233,N2234,N2235,
     N2236,N2237,N2240,N2241,N2244,N2245,N2250,N2253,N2256,N2257,
     N2260,N2263,N2266,N2269,N2272,N2279,N2286,N2297,N2315,N2326,
     N2340,N2353,N2361,N2375,N2384,N2385,N2386,N2426,N2427,N2537,
     N2540,N2543,N2546,N2549,N2552,N2555,N2558,N2561,N2564,N2567,
     N2570,N2573,N2576,N2594,N2597,N2600,N2603,N2606,N2611,N2614,
     N2617,N2620,N2627,N2628,N2629,N2630,N2631,N2632,N2633,N2634,
     N2639,N2642,N2645,N2648,N2651,N2655,N2658,N2661,N2664,N2669,
     N2670,N2671,N2672,N2673,N2674,N2675,N2676,N2682,N2683,N2688,
     N2689,N2690,N2691,N2710,N2720,N2721,N2722,N2723,N2724,N2725,
     N2726,N2727,N2728,N2729,N2730,N2731,N2732,N2733,N2734,N2735,
     N2736,N2737,N2738,N2739,N2740,N2741,N2742,N2743,N2744,N2745,
     N2746,N2747,N2750,N2757,N2758,N2759,N2760,N2761,N2763,N2764,
     N2765,N2766,N2773,N2776,N2788,N2789,N2800,N2807,N2808,N2809,
     N2810,N2812,N2815,N2818,N2821,N2824,N2827,N2828,N2829,N2843,
     N2846,N2850,N2851,N2852,N2853,N2854,N2857,N2858,N2859,N2860,
     N2861,N2862,N2863,N2866,N2867,N2868,N2869,N2870,N2871,N2872,
     N2873,N2874,N2875,N2876,N2877,N2878,N2879,N2880,N2881,N2882,
     N2883,N2895,N2896,N2897,N2898, gate773inter0, gate773inter1, gate773inter2, gate773inter3, gate773inter4, gate773inter5, gate773inter6, gate773inter7, gate773inter8, gate773inter9, gate773inter10, gate773inter11, gate773inter12, gate754inter0, gate754inter1, gate754inter2, gate754inter3, gate754inter4, gate754inter5, gate754inter6, gate754inter7, gate754inter8, gate754inter9, gate754inter10, gate754inter11, gate754inter12, gate854inter0, gate854inter1, gate854inter2, gate854inter3, gate854inter4, gate854inter5, gate854inter6, gate854inter7, gate854inter8, gate854inter9, gate854inter10, gate854inter11, gate854inter12, gate586inter0, gate586inter1, gate586inter2, gate586inter3, gate586inter4, gate586inter5, gate586inter6, gate586inter7, gate586inter8, gate586inter9, gate586inter10, gate586inter11, gate586inter12, gate321inter0, gate321inter1, gate321inter2, gate321inter3, gate321inter4, gate321inter5, gate321inter6, gate321inter7, gate321inter8, gate321inter9, gate321inter10, gate321inter11, gate321inter12, gate233inter0, gate233inter1, gate233inter2, gate233inter3, gate233inter4, gate233inter5, gate233inter6, gate233inter7, gate233inter8, gate233inter9, gate233inter10, gate233inter11, gate233inter12, gate527inter0, gate527inter1, gate527inter2, gate527inter3, gate527inter4, gate527inter5, gate527inter6, gate527inter7, gate527inter8, gate527inter9, gate527inter10, gate527inter11, gate527inter12, gate499inter0, gate499inter1, gate499inter2, gate499inter3, gate499inter4, gate499inter5, gate499inter6, gate499inter7, gate499inter8, gate499inter9, gate499inter10, gate499inter11, gate499inter12, gate294inter0, gate294inter1, gate294inter2, gate294inter3, gate294inter4, gate294inter5, gate294inter6, gate294inter7, gate294inter8, gate294inter9, gate294inter10, gate294inter11, gate294inter12, gate683inter0, gate683inter1, gate683inter2, gate683inter3, gate683inter4, gate683inter5, gate683inter6, gate683inter7, gate683inter8, gate683inter9, gate683inter10, gate683inter11, gate683inter12, gate809inter0, gate809inter1, gate809inter2, gate809inter3, gate809inter4, gate809inter5, gate809inter6, gate809inter7, gate809inter8, gate809inter9, gate809inter10, gate809inter11, gate809inter12, gate339inter0, gate339inter1, gate339inter2, gate339inter3, gate339inter4, gate339inter5, gate339inter6, gate339inter7, gate339inter8, gate339inter9, gate339inter10, gate339inter11, gate339inter12, gate338inter0, gate338inter1, gate338inter2, gate338inter3, gate338inter4, gate338inter5, gate338inter6, gate338inter7, gate338inter8, gate338inter9, gate338inter10, gate338inter11, gate338inter12, gate350inter0, gate350inter1, gate350inter2, gate350inter3, gate350inter4, gate350inter5, gate350inter6, gate350inter7, gate350inter8, gate350inter9, gate350inter10, gate350inter11, gate350inter12, gate805inter0, gate805inter1, gate805inter2, gate805inter3, gate805inter4, gate805inter5, gate805inter6, gate805inter7, gate805inter8, gate805inter9, gate805inter10, gate805inter11, gate805inter12, gate412inter0, gate412inter1, gate412inter2, gate412inter3, gate412inter4, gate412inter5, gate412inter6, gate412inter7, gate412inter8, gate412inter9, gate412inter10, gate412inter11, gate412inter12, gate376inter0, gate376inter1, gate376inter2, gate376inter3, gate376inter4, gate376inter5, gate376inter6, gate376inter7, gate376inter8, gate376inter9, gate376inter10, gate376inter11, gate376inter12, gate563inter0, gate563inter1, gate563inter2, gate563inter3, gate563inter4, gate563inter5, gate563inter6, gate563inter7, gate563inter8, gate563inter9, gate563inter10, gate563inter11, gate563inter12, gate478inter0, gate478inter1, gate478inter2, gate478inter3, gate478inter4, gate478inter5, gate478inter6, gate478inter7, gate478inter8, gate478inter9, gate478inter10, gate478inter11, gate478inter12, gate335inter0, gate335inter1, gate335inter2, gate335inter3, gate335inter4, gate335inter5, gate335inter6, gate335inter7, gate335inter8, gate335inter9, gate335inter10, gate335inter11, gate335inter12, gate600inter0, gate600inter1, gate600inter2, gate600inter3, gate600inter4, gate600inter5, gate600inter6, gate600inter7, gate600inter8, gate600inter9, gate600inter10, gate600inter11, gate600inter12, gate574inter0, gate574inter1, gate574inter2, gate574inter3, gate574inter4, gate574inter5, gate574inter6, gate574inter7, gate574inter8, gate574inter9, gate574inter10, gate574inter11, gate574inter12, gate529inter0, gate529inter1, gate529inter2, gate529inter3, gate529inter4, gate529inter5, gate529inter6, gate529inter7, gate529inter8, gate529inter9, gate529inter10, gate529inter11, gate529inter12, gate419inter0, gate419inter1, gate419inter2, gate419inter3, gate419inter4, gate419inter5, gate419inter6, gate419inter7, gate419inter8, gate419inter9, gate419inter10, gate419inter11, gate419inter12, gate496inter0, gate496inter1, gate496inter2, gate496inter3, gate496inter4, gate496inter5, gate496inter6, gate496inter7, gate496inter8, gate496inter9, gate496inter10, gate496inter11, gate496inter12, gate396inter0, gate396inter1, gate396inter2, gate396inter3, gate396inter4, gate396inter5, gate396inter6, gate396inter7, gate396inter8, gate396inter9, gate396inter10, gate396inter11, gate396inter12, gate824inter0, gate824inter1, gate824inter2, gate824inter3, gate824inter4, gate824inter5, gate824inter6, gate824inter7, gate824inter8, gate824inter9, gate824inter10, gate824inter11, gate824inter12, gate234inter0, gate234inter1, gate234inter2, gate234inter3, gate234inter4, gate234inter5, gate234inter6, gate234inter7, gate234inter8, gate234inter9, gate234inter10, gate234inter11, gate234inter12, gate862inter0, gate862inter1, gate862inter2, gate862inter3, gate862inter4, gate862inter5, gate862inter6, gate862inter7, gate862inter8, gate862inter9, gate862inter10, gate862inter11, gate862inter12, gate163inter0, gate163inter1, gate163inter2, gate163inter3, gate163inter4, gate163inter5, gate163inter6, gate163inter7, gate163inter8, gate163inter9, gate163inter10, gate163inter11, gate163inter12, gate418inter0, gate418inter1, gate418inter2, gate418inter3, gate418inter4, gate418inter5, gate418inter6, gate418inter7, gate418inter8, gate418inter9, gate418inter10, gate418inter11, gate418inter12, gate852inter0, gate852inter1, gate852inter2, gate852inter3, gate852inter4, gate852inter5, gate852inter6, gate852inter7, gate852inter8, gate852inter9, gate852inter10, gate852inter11, gate852inter12, gate503inter0, gate503inter1, gate503inter2, gate503inter3, gate503inter4, gate503inter5, gate503inter6, gate503inter7, gate503inter8, gate503inter9, gate503inter10, gate503inter11, gate503inter12, gate633inter0, gate633inter1, gate633inter2, gate633inter3, gate633inter4, gate633inter5, gate633inter6, gate633inter7, gate633inter8, gate633inter9, gate633inter10, gate633inter11, gate633inter12, gate240inter0, gate240inter1, gate240inter2, gate240inter3, gate240inter4, gate240inter5, gate240inter6, gate240inter7, gate240inter8, gate240inter9, gate240inter10, gate240inter11, gate240inter12, gate526inter0, gate526inter1, gate526inter2, gate526inter3, gate526inter4, gate526inter5, gate526inter6, gate526inter7, gate526inter8, gate526inter9, gate526inter10, gate526inter11, gate526inter12, gate243inter0, gate243inter1, gate243inter2, gate243inter3, gate243inter4, gate243inter5, gate243inter6, gate243inter7, gate243inter8, gate243inter9, gate243inter10, gate243inter11, gate243inter12, gate625inter0, gate625inter1, gate625inter2, gate625inter3, gate625inter4, gate625inter5, gate625inter6, gate625inter7, gate625inter8, gate625inter9, gate625inter10, gate625inter11, gate625inter12, gate623inter0, gate623inter1, gate623inter2, gate623inter3, gate623inter4, gate623inter5, gate623inter6, gate623inter7, gate623inter8, gate623inter9, gate623inter10, gate623inter11, gate623inter12, gate624inter0, gate624inter1, gate624inter2, gate624inter3, gate624inter4, gate624inter5, gate624inter6, gate624inter7, gate624inter8, gate624inter9, gate624inter10, gate624inter11, gate624inter12, gate851inter0, gate851inter1, gate851inter2, gate851inter3, gate851inter4, gate851inter5, gate851inter6, gate851inter7, gate851inter8, gate851inter9, gate851inter10, gate851inter11, gate851inter12, gate298inter0, gate298inter1, gate298inter2, gate298inter3, gate298inter4, gate298inter5, gate298inter6, gate298inter7, gate298inter8, gate298inter9, gate298inter10, gate298inter11, gate298inter12, gate237inter0, gate237inter1, gate237inter2, gate237inter3, gate237inter4, gate237inter5, gate237inter6, gate237inter7, gate237inter8, gate237inter9, gate237inter10, gate237inter11, gate237inter12, gate401inter0, gate401inter1, gate401inter2, gate401inter3, gate401inter4, gate401inter5, gate401inter6, gate401inter7, gate401inter8, gate401inter9, gate401inter10, gate401inter11, gate401inter12, gate612inter0, gate612inter1, gate612inter2, gate612inter3, gate612inter4, gate612inter5, gate612inter6, gate612inter7, gate612inter8, gate612inter9, gate612inter10, gate612inter11, gate612inter12, gate528inter0, gate528inter1, gate528inter2, gate528inter3, gate528inter4, gate528inter5, gate528inter6, gate528inter7, gate528inter8, gate528inter9, gate528inter10, gate528inter11, gate528inter12, gate406inter0, gate406inter1, gate406inter2, gate406inter3, gate406inter4, gate406inter5, gate406inter6, gate406inter7, gate406inter8, gate406inter9, gate406inter10, gate406inter11, gate406inter12, gate635inter0, gate635inter1, gate635inter2, gate635inter3, gate635inter4, gate635inter5, gate635inter6, gate635inter7, gate635inter8, gate635inter9, gate635inter10, gate635inter11, gate635inter12, gate387inter0, gate387inter1, gate387inter2, gate387inter3, gate387inter4, gate387inter5, gate387inter6, gate387inter7, gate387inter8, gate387inter9, gate387inter10, gate387inter11, gate387inter12, gate628inter0, gate628inter1, gate628inter2, gate628inter3, gate628inter4, gate628inter5, gate628inter6, gate628inter7, gate628inter8, gate628inter9, gate628inter10, gate628inter11, gate628inter12, gate261inter0, gate261inter1, gate261inter2, gate261inter3, gate261inter4, gate261inter5, gate261inter6, gate261inter7, gate261inter8, gate261inter9, gate261inter10, gate261inter11, gate261inter12, gate539inter0, gate539inter1, gate539inter2, gate539inter3, gate539inter4, gate539inter5, gate539inter6, gate539inter7, gate539inter8, gate539inter9, gate539inter10, gate539inter11, gate539inter12, gate616inter0, gate616inter1, gate616inter2, gate616inter3, gate616inter4, gate616inter5, gate616inter6, gate616inter7, gate616inter8, gate616inter9, gate616inter10, gate616inter11, gate616inter12, gate405inter0, gate405inter1, gate405inter2, gate405inter3, gate405inter4, gate405inter5, gate405inter6, gate405inter7, gate405inter8, gate405inter9, gate405inter10, gate405inter11, gate405inter12, gate839inter0, gate839inter1, gate839inter2, gate839inter3, gate839inter4, gate839inter5, gate839inter6, gate839inter7, gate839inter8, gate839inter9, gate839inter10, gate839inter11, gate839inter12, gate607inter0, gate607inter1, gate607inter2, gate607inter3, gate607inter4, gate607inter5, gate607inter6, gate607inter7, gate607inter8, gate607inter9, gate607inter10, gate607inter11, gate607inter12, gate814inter0, gate814inter1, gate814inter2, gate814inter3, gate814inter4, gate814inter5, gate814inter6, gate814inter7, gate814inter8, gate814inter9, gate814inter10, gate814inter11, gate814inter12, gate547inter0, gate547inter1, gate547inter2, gate547inter3, gate547inter4, gate547inter5, gate547inter6, gate547inter7, gate547inter8, gate547inter9, gate547inter10, gate547inter11, gate547inter12, gate385inter0, gate385inter1, gate385inter2, gate385inter3, gate385inter4, gate385inter5, gate385inter6, gate385inter7, gate385inter8, gate385inter9, gate385inter10, gate385inter11, gate385inter12, gate756inter0, gate756inter1, gate756inter2, gate756inter3, gate756inter4, gate756inter5, gate756inter6, gate756inter7, gate756inter8, gate756inter9, gate756inter10, gate756inter11, gate756inter12, gate76inter0, gate76inter1, gate76inter2, gate76inter3, gate76inter4, gate76inter5, gate76inter6, gate76inter7, gate76inter8, gate76inter9, gate76inter10, gate76inter11, gate76inter12, gate806inter0, gate806inter1, gate806inter2, gate806inter3, gate806inter4, gate806inter5, gate806inter6, gate806inter7, gate806inter8, gate806inter9, gate806inter10, gate806inter11, gate806inter12, gate780inter0, gate780inter1, gate780inter2, gate780inter3, gate780inter4, gate780inter5, gate780inter6, gate780inter7, gate780inter8, gate780inter9, gate780inter10, gate780inter11, gate780inter12, gate523inter0, gate523inter1, gate523inter2, gate523inter3, gate523inter4, gate523inter5, gate523inter6, gate523inter7, gate523inter8, gate523inter9, gate523inter10, gate523inter11, gate523inter12, gate343inter0, gate343inter1, gate343inter2, gate343inter3, gate343inter4, gate343inter5, gate343inter6, gate343inter7, gate343inter8, gate343inter9, gate343inter10, gate343inter11, gate343inter12, gate337inter0, gate337inter1, gate337inter2, gate337inter3, gate337inter4, gate337inter5, gate337inter6, gate337inter7, gate337inter8, gate337inter9, gate337inter10, gate337inter11, gate337inter12;


inv1 gate1( .a(N1), .O(N190) );
inv1 gate2( .a(N4), .O(N194) );
inv1 gate3( .a(N7), .O(N197) );
inv1 gate4( .a(N10), .O(N201) );
inv1 gate5( .a(N13), .O(N206) );
inv1 gate6( .a(N16), .O(N209) );
inv1 gate7( .a(N19), .O(N212) );
inv1 gate8( .a(N22), .O(N216) );
inv1 gate9( .a(N25), .O(N220) );
inv1 gate10( .a(N28), .O(N225) );
inv1 gate11( .a(N31), .O(N229) );
inv1 gate12( .a(N34), .O(N232) );
inv1 gate13( .a(N37), .O(N235) );
inv1 gate14( .a(N40), .O(N239) );
inv1 gate15( .a(N43), .O(N243) );
inv1 gate16( .a(N46), .O(N247) );
nand2 gate17( .a(N63), .b(N88), .O(N251) );
nand2 gate18( .a(N66), .b(N91), .O(N252) );
inv1 gate19( .a(N72), .O(N253) );
inv1 gate20( .a(N72), .O(N256) );
buf1 gate21( .a(N69), .O(N257) );
buf1 gate22( .a(N69), .O(N260) );
inv1 gate23( .a(N76), .O(N263) );
inv1 gate24( .a(N79), .O(N266) );
inv1 gate25( .a(N82), .O(N269) );
inv1 gate26( .a(N85), .O(N272) );
inv1 gate27( .a(N104), .O(N275) );
inv1 gate28( .a(N104), .O(N276) );
inv1 gate29( .a(N88), .O(N277) );
inv1 gate30( .a(N91), .O(N280) );
buf1 gate31( .a(N94), .O(N283) );
inv1 gate32( .a(N94), .O(N290) );
buf1 gate33( .a(N94), .O(N297) );
inv1 gate34( .a(N94), .O(N300) );
buf1 gate35( .a(N99), .O(N303) );
inv1 gate36( .a(N99), .O(N306) );
inv1 gate37( .a(N99), .O(N313) );
buf1 gate38( .a(N104), .O(N316) );
inv1 gate39( .a(N104), .O(N319) );
buf1 gate40( .a(N104), .O(N326) );
buf1 gate41( .a(N104), .O(N331) );
inv1 gate42( .a(N104), .O(N338) );
buf1 gate43( .a(N1), .O(N343) );
buf1 gate44( .a(N4), .O(N346) );
buf1 gate45( .a(N7), .O(N349) );
buf1 gate46( .a(N10), .O(N352) );
buf1 gate47( .a(N13), .O(N355) );
buf1 gate48( .a(N16), .O(N358) );
buf1 gate49( .a(N19), .O(N361) );
buf1 gate50( .a(N22), .O(N364) );
buf1 gate51( .a(N25), .O(N367) );
buf1 gate52( .a(N28), .O(N370) );
buf1 gate53( .a(N31), .O(N373) );
buf1 gate54( .a(N34), .O(N376) );
buf1 gate55( .a(N37), .O(N379) );
buf1 gate56( .a(N40), .O(N382) );
buf1 gate57( .a(N43), .O(N385) );
buf1 gate58( .a(N46), .O(N388) );
inv1 gate59( .a(N343), .O(N534) );
inv1 gate60( .a(N346), .O(N535) );
inv1 gate61( .a(N349), .O(N536) );
inv1 gate62( .a(N352), .O(N537) );
inv1 gate63( .a(N355), .O(N538) );
inv1 gate64( .a(N358), .O(N539) );
inv1 gate65( .a(N361), .O(N540) );
inv1 gate66( .a(N364), .O(N541) );
inv1 gate67( .a(N367), .O(N542) );
inv1 gate68( .a(N370), .O(N543) );
inv1 gate69( .a(N373), .O(N544) );
inv1 gate70( .a(N376), .O(N545) );
inv1 gate71( .a(N379), .O(N546) );
inv1 gate72( .a(N382), .O(N547) );
inv1 gate73( .a(N385), .O(N548) );
inv1 gate74( .a(N388), .O(N549) );
nand2 gate75( .a(N306), .b(N331), .O(N550) );

  xor2  gate1721(.a(N331), .b(N306), .O(gate76inter0));
  nand2 gate1722(.a(gate76inter0), .b(s_120), .O(gate76inter1));
  and2  gate1723(.a(N331), .b(N306), .O(gate76inter2));
  inv1  gate1724(.a(s_120), .O(gate76inter3));
  inv1  gate1725(.a(s_121), .O(gate76inter4));
  nand2 gate1726(.a(gate76inter4), .b(gate76inter3), .O(gate76inter5));
  nor2  gate1727(.a(gate76inter5), .b(gate76inter2), .O(gate76inter6));
  inv1  gate1728(.a(N306), .O(gate76inter7));
  inv1  gate1729(.a(N331), .O(gate76inter8));
  nand2 gate1730(.a(gate76inter8), .b(gate76inter7), .O(gate76inter9));
  nand2 gate1731(.a(s_121), .b(gate76inter3), .O(gate76inter10));
  nor2  gate1732(.a(gate76inter10), .b(gate76inter9), .O(gate76inter11));
  nor2  gate1733(.a(gate76inter11), .b(gate76inter6), .O(gate76inter12));
  nand2 gate1734(.a(gate76inter12), .b(gate76inter1), .O(N551));
nand2 gate77( .a(N306), .b(N331), .O(N552) );
nand2 gate78( .a(N306), .b(N331), .O(N553) );
nand2 gate79( .a(N306), .b(N331), .O(N554) );
nand2 gate80( .a(N306), .b(N331), .O(N555) );
buf1 gate81( .a(N190), .O(N556) );
buf1 gate82( .a(N194), .O(N559) );
buf1 gate83( .a(N206), .O(N562) );
buf1 gate84( .a(N209), .O(N565) );
buf1 gate85( .a(N225), .O(N568) );
buf1 gate86( .a(N243), .O(N571) );
and2 gate87( .a(N63), .b(N319), .O(N574) );
buf1 gate88( .a(N220), .O(N577) );
buf1 gate89( .a(N229), .O(N580) );
buf1 gate90( .a(N232), .O(N583) );
and2 gate91( .a(N66), .b(N319), .O(N586) );
buf1 gate92( .a(N239), .O(N589) );
and3 gate93( .a(N49), .b(N253), .c(N319), .O(N592) );
buf1 gate94( .a(N247), .O(N595) );
buf1 gate95( .a(N239), .O(N598) );
nand2 gate96( .a(N326), .b(N277), .O(N601) );
nand2 gate97( .a(N326), .b(N280), .O(N602) );
nand2 gate98( .a(N260), .b(N72), .O(N603) );
nand2 gate99( .a(N260), .b(N300), .O(N608) );
nand2 gate100( .a(N256), .b(N300), .O(N612) );
buf1 gate101( .a(N201), .O(N616) );
buf1 gate102( .a(N216), .O(N619) );
buf1 gate103( .a(N220), .O(N622) );
buf1 gate104( .a(N239), .O(N625) );
buf1 gate105( .a(N190), .O(N628) );
buf1 gate106( .a(N190), .O(N631) );
buf1 gate107( .a(N194), .O(N634) );
buf1 gate108( .a(N229), .O(N637) );
buf1 gate109( .a(N197), .O(N640) );
and3 gate110( .a(N56), .b(N257), .c(N319), .O(N643) );
buf1 gate111( .a(N232), .O(N646) );
buf1 gate112( .a(N201), .O(N649) );
buf1 gate113( .a(N235), .O(N652) );
and3 gate114( .a(N60), .b(N257), .c(N319), .O(N655) );
buf1 gate115( .a(N263), .O(N658) );
buf1 gate116( .a(N263), .O(N661) );
buf1 gate117( .a(N266), .O(N664) );
buf1 gate118( .a(N266), .O(N667) );
buf1 gate119( .a(N269), .O(N670) );
buf1 gate120( .a(N269), .O(N673) );
buf1 gate121( .a(N272), .O(N676) );
buf1 gate122( .a(N272), .O(N679) );
and2 gate123( .a(N251), .b(N316), .O(N682) );
and2 gate124( .a(N252), .b(N316), .O(N685) );
buf1 gate125( .a(N197), .O(N688) );
buf1 gate126( .a(N197), .O(N691) );
buf1 gate127( .a(N212), .O(N694) );
buf1 gate128( .a(N212), .O(N697) );
buf1 gate129( .a(N247), .O(N700) );
buf1 gate130( .a(N247), .O(N703) );
buf1 gate131( .a(N235), .O(N706) );
buf1 gate132( .a(N235), .O(N709) );
buf1 gate133( .a(N201), .O(N712) );
buf1 gate134( .a(N201), .O(N715) );
buf1 gate135( .a(N206), .O(N718) );
buf1 gate136( .a(N216), .O(N721) );
and3 gate137( .a(N53), .b(N253), .c(N319), .O(N724) );
buf1 gate138( .a(N243), .O(N727) );
buf1 gate139( .a(N220), .O(N730) );
buf1 gate140( .a(N220), .O(N733) );
buf1 gate141( .a(N209), .O(N736) );
buf1 gate142( .a(N216), .O(N739) );
buf1 gate143( .a(N225), .O(N742) );
buf1 gate144( .a(N243), .O(N745) );
buf1 gate145( .a(N212), .O(N748) );
buf1 gate146( .a(N225), .O(N751) );
inv1 gate147( .a(N682), .O(N886) );
inv1 gate148( .a(N685), .O(N887) );
inv1 gate149( .a(N616), .O(N888) );
inv1 gate150( .a(N619), .O(N889) );
inv1 gate151( .a(N622), .O(N890) );
inv1 gate152( .a(N625), .O(N891) );
inv1 gate153( .a(N631), .O(N892) );
inv1 gate154( .a(N643), .O(N893) );
inv1 gate155( .a(N649), .O(N894) );
inv1 gate156( .a(N652), .O(N895) );
inv1 gate157( .a(N655), .O(N896) );
and2 gate158( .a(N49), .b(N612), .O(N897) );
and2 gate159( .a(N56), .b(N608), .O(N898) );
nand2 gate160( .a(N53), .b(N612), .O(N899) );
nand2 gate161( .a(N60), .b(N608), .O(N903) );
nand2 gate162( .a(N49), .b(N612), .O(N907) );

  xor2  gate1287(.a(N608), .b(N56), .O(gate163inter0));
  nand2 gate1288(.a(gate163inter0), .b(s_58), .O(gate163inter1));
  and2  gate1289(.a(N608), .b(N56), .O(gate163inter2));
  inv1  gate1290(.a(s_58), .O(gate163inter3));
  inv1  gate1291(.a(s_59), .O(gate163inter4));
  nand2 gate1292(.a(gate163inter4), .b(gate163inter3), .O(gate163inter5));
  nor2  gate1293(.a(gate163inter5), .b(gate163inter2), .O(gate163inter6));
  inv1  gate1294(.a(N56), .O(gate163inter7));
  inv1  gate1295(.a(N608), .O(gate163inter8));
  nand2 gate1296(.a(gate163inter8), .b(gate163inter7), .O(gate163inter9));
  nand2 gate1297(.a(s_59), .b(gate163inter3), .O(gate163inter10));
  nor2  gate1298(.a(gate163inter10), .b(gate163inter9), .O(gate163inter11));
  nor2  gate1299(.a(gate163inter11), .b(gate163inter6), .O(gate163inter12));
  nand2 gate1300(.a(gate163inter12), .b(gate163inter1), .O(N910));
inv1 gate164( .a(N661), .O(N913) );
inv1 gate165( .a(N658), .O(N914) );
inv1 gate166( .a(N667), .O(N915) );
inv1 gate167( .a(N664), .O(N916) );
inv1 gate168( .a(N673), .O(N917) );
inv1 gate169( .a(N670), .O(N918) );
inv1 gate170( .a(N679), .O(N919) );
inv1 gate171( .a(N676), .O(N920) );
nand4 gate172( .a(N277), .b(N297), .c(N326), .d(N603), .O(N921) );
nand4 gate173( .a(N280), .b(N297), .c(N326), .d(N603), .O(N922) );
nand3 gate174( .a(N303), .b(N338), .c(N603), .O(N923) );
and3 gate175( .a(N303), .b(N338), .c(N603), .O(N926) );
buf1 gate176( .a(N556), .O(N935) );
inv1 gate177( .a(N688), .O(N938) );
buf1 gate178( .a(N556), .O(N939) );
inv1 gate179( .a(N691), .O(N942) );
buf1 gate180( .a(N562), .O(N943) );
inv1 gate181( .a(N694), .O(N946) );
buf1 gate182( .a(N562), .O(N947) );
inv1 gate183( .a(N697), .O(N950) );
buf1 gate184( .a(N568), .O(N951) );
inv1 gate185( .a(N700), .O(N954) );
buf1 gate186( .a(N568), .O(N955) );
inv1 gate187( .a(N703), .O(N958) );
buf1 gate188( .a(N574), .O(N959) );
buf1 gate189( .a(N574), .O(N962) );
buf1 gate190( .a(N580), .O(N965) );
inv1 gate191( .a(N706), .O(N968) );
buf1 gate192( .a(N580), .O(N969) );
inv1 gate193( .a(N709), .O(N972) );
buf1 gate194( .a(N586), .O(N973) );
inv1 gate195( .a(N712), .O(N976) );
buf1 gate196( .a(N586), .O(N977) );
inv1 gate197( .a(N715), .O(N980) );
buf1 gate198( .a(N592), .O(N981) );
inv1 gate199( .a(N628), .O(N984) );
buf1 gate200( .a(N592), .O(N985) );
inv1 gate201( .a(N718), .O(N988) );
inv1 gate202( .a(N721), .O(N989) );
inv1 gate203( .a(N634), .O(N990) );
inv1 gate204( .a(N724), .O(N991) );
inv1 gate205( .a(N727), .O(N992) );
inv1 gate206( .a(N637), .O(N993) );
buf1 gate207( .a(N595), .O(N994) );
inv1 gate208( .a(N730), .O(N997) );
buf1 gate209( .a(N595), .O(N998) );
inv1 gate210( .a(N733), .O(N1001) );
inv1 gate211( .a(N736), .O(N1002) );
inv1 gate212( .a(N739), .O(N1003) );
inv1 gate213( .a(N640), .O(N1004) );
inv1 gate214( .a(N742), .O(N1005) );
inv1 gate215( .a(N745), .O(N1006) );
inv1 gate216( .a(N646), .O(N1007) );
inv1 gate217( .a(N748), .O(N1008) );
inv1 gate218( .a(N751), .O(N1009) );
buf1 gate219( .a(N559), .O(N1010) );
buf1 gate220( .a(N559), .O(N1013) );
buf1 gate221( .a(N565), .O(N1016) );
buf1 gate222( .a(N565), .O(N1019) );
buf1 gate223( .a(N571), .O(N1022) );
buf1 gate224( .a(N571), .O(N1025) );
buf1 gate225( .a(N577), .O(N1028) );
buf1 gate226( .a(N577), .O(N1031) );
buf1 gate227( .a(N583), .O(N1034) );
buf1 gate228( .a(N583), .O(N1037) );
buf1 gate229( .a(N589), .O(N1040) );
buf1 gate230( .a(N589), .O(N1043) );
buf1 gate231( .a(N598), .O(N1046) );
buf1 gate232( .a(N598), .O(N1049) );

  xor2  gate951(.a(N888), .b(N619), .O(gate233inter0));
  nand2 gate952(.a(gate233inter0), .b(s_10), .O(gate233inter1));
  and2  gate953(.a(N888), .b(N619), .O(gate233inter2));
  inv1  gate954(.a(s_10), .O(gate233inter3));
  inv1  gate955(.a(s_11), .O(gate233inter4));
  nand2 gate956(.a(gate233inter4), .b(gate233inter3), .O(gate233inter5));
  nor2  gate957(.a(gate233inter5), .b(gate233inter2), .O(gate233inter6));
  inv1  gate958(.a(N619), .O(gate233inter7));
  inv1  gate959(.a(N888), .O(gate233inter8));
  nand2 gate960(.a(gate233inter8), .b(gate233inter7), .O(gate233inter9));
  nand2 gate961(.a(s_11), .b(gate233inter3), .O(gate233inter10));
  nor2  gate962(.a(gate233inter10), .b(gate233inter9), .O(gate233inter11));
  nor2  gate963(.a(gate233inter11), .b(gate233inter6), .O(gate233inter12));
  nand2 gate964(.a(gate233inter12), .b(gate233inter1), .O(N1054));

  xor2  gate1259(.a(N889), .b(N616), .O(gate234inter0));
  nand2 gate1260(.a(gate234inter0), .b(s_54), .O(gate234inter1));
  and2  gate1261(.a(N889), .b(N616), .O(gate234inter2));
  inv1  gate1262(.a(s_54), .O(gate234inter3));
  inv1  gate1263(.a(s_55), .O(gate234inter4));
  nand2 gate1264(.a(gate234inter4), .b(gate234inter3), .O(gate234inter5));
  nor2  gate1265(.a(gate234inter5), .b(gate234inter2), .O(gate234inter6));
  inv1  gate1266(.a(N616), .O(gate234inter7));
  inv1  gate1267(.a(N889), .O(gate234inter8));
  nand2 gate1268(.a(gate234inter8), .b(gate234inter7), .O(gate234inter9));
  nand2 gate1269(.a(s_55), .b(gate234inter3), .O(gate234inter10));
  nor2  gate1270(.a(gate234inter10), .b(gate234inter9), .O(gate234inter11));
  nor2  gate1271(.a(gate234inter11), .b(gate234inter6), .O(gate234inter12));
  nand2 gate1272(.a(gate234inter12), .b(gate234inter1), .O(N1055));
nand2 gate235( .a(N625), .b(N890), .O(N1063) );
nand2 gate236( .a(N622), .b(N891), .O(N1064) );

  xor2  gate1469(.a(N895), .b(N655), .O(gate237inter0));
  nand2 gate1470(.a(gate237inter0), .b(s_84), .O(gate237inter1));
  and2  gate1471(.a(N895), .b(N655), .O(gate237inter2));
  inv1  gate1472(.a(s_84), .O(gate237inter3));
  inv1  gate1473(.a(s_85), .O(gate237inter4));
  nand2 gate1474(.a(gate237inter4), .b(gate237inter3), .O(gate237inter5));
  nor2  gate1475(.a(gate237inter5), .b(gate237inter2), .O(gate237inter6));
  inv1  gate1476(.a(N655), .O(gate237inter7));
  inv1  gate1477(.a(N895), .O(gate237inter8));
  nand2 gate1478(.a(gate237inter8), .b(gate237inter7), .O(gate237inter9));
  nand2 gate1479(.a(s_85), .b(gate237inter3), .O(gate237inter10));
  nor2  gate1480(.a(gate237inter10), .b(gate237inter9), .O(gate237inter11));
  nor2  gate1481(.a(gate237inter11), .b(gate237inter6), .O(gate237inter12));
  nand2 gate1482(.a(gate237inter12), .b(gate237inter1), .O(N1067));
nand2 gate238( .a(N652), .b(N896), .O(N1068) );
nand2 gate239( .a(N721), .b(N988), .O(N1119) );

  xor2  gate1357(.a(N989), .b(N718), .O(gate240inter0));
  nand2 gate1358(.a(gate240inter0), .b(s_68), .O(gate240inter1));
  and2  gate1359(.a(N989), .b(N718), .O(gate240inter2));
  inv1  gate1360(.a(s_68), .O(gate240inter3));
  inv1  gate1361(.a(s_69), .O(gate240inter4));
  nand2 gate1362(.a(gate240inter4), .b(gate240inter3), .O(gate240inter5));
  nor2  gate1363(.a(gate240inter5), .b(gate240inter2), .O(gate240inter6));
  inv1  gate1364(.a(N718), .O(gate240inter7));
  inv1  gate1365(.a(N989), .O(gate240inter8));
  nand2 gate1366(.a(gate240inter8), .b(gate240inter7), .O(gate240inter9));
  nand2 gate1367(.a(s_69), .b(gate240inter3), .O(gate240inter10));
  nor2  gate1368(.a(gate240inter10), .b(gate240inter9), .O(gate240inter11));
  nor2  gate1369(.a(gate240inter11), .b(gate240inter6), .O(gate240inter12));
  nand2 gate1370(.a(gate240inter12), .b(gate240inter1), .O(N1120));
nand2 gate241( .a(N727), .b(N991), .O(N1121) );
nand2 gate242( .a(N724), .b(N992), .O(N1122) );

  xor2  gate1385(.a(N1002), .b(N739), .O(gate243inter0));
  nand2 gate1386(.a(gate243inter0), .b(s_72), .O(gate243inter1));
  and2  gate1387(.a(N1002), .b(N739), .O(gate243inter2));
  inv1  gate1388(.a(s_72), .O(gate243inter3));
  inv1  gate1389(.a(s_73), .O(gate243inter4));
  nand2 gate1390(.a(gate243inter4), .b(gate243inter3), .O(gate243inter5));
  nor2  gate1391(.a(gate243inter5), .b(gate243inter2), .O(gate243inter6));
  inv1  gate1392(.a(N739), .O(gate243inter7));
  inv1  gate1393(.a(N1002), .O(gate243inter8));
  nand2 gate1394(.a(gate243inter8), .b(gate243inter7), .O(gate243inter9));
  nand2 gate1395(.a(s_73), .b(gate243inter3), .O(gate243inter10));
  nor2  gate1396(.a(gate243inter10), .b(gate243inter9), .O(gate243inter11));
  nor2  gate1397(.a(gate243inter11), .b(gate243inter6), .O(gate243inter12));
  nand2 gate1398(.a(gate243inter12), .b(gate243inter1), .O(N1128));
nand2 gate244( .a(N736), .b(N1003), .O(N1129) );
nand2 gate245( .a(N745), .b(N1005), .O(N1130) );
nand2 gate246( .a(N742), .b(N1006), .O(N1131) );
nand2 gate247( .a(N751), .b(N1008), .O(N1132) );
nand2 gate248( .a(N748), .b(N1009), .O(N1133) );
inv1 gate249( .a(N939), .O(N1148) );
inv1 gate250( .a(N935), .O(N1149) );
nand2 gate251( .a(N1054), .b(N1055), .O(N1150) );
inv1 gate252( .a(N943), .O(N1151) );
inv1 gate253( .a(N947), .O(N1152) );
inv1 gate254( .a(N955), .O(N1153) );
inv1 gate255( .a(N951), .O(N1154) );
inv1 gate256( .a(N962), .O(N1155) );
inv1 gate257( .a(N969), .O(N1156) );
inv1 gate258( .a(N977), .O(N1157) );
nand2 gate259( .a(N1063), .b(N1064), .O(N1158) );
inv1 gate260( .a(N985), .O(N1159) );

  xor2  gate1581(.a(N892), .b(N985), .O(gate261inter0));
  nand2 gate1582(.a(gate261inter0), .b(s_100), .O(gate261inter1));
  and2  gate1583(.a(N892), .b(N985), .O(gate261inter2));
  inv1  gate1584(.a(s_100), .O(gate261inter3));
  inv1  gate1585(.a(s_101), .O(gate261inter4));
  nand2 gate1586(.a(gate261inter4), .b(gate261inter3), .O(gate261inter5));
  nor2  gate1587(.a(gate261inter5), .b(gate261inter2), .O(gate261inter6));
  inv1  gate1588(.a(N985), .O(gate261inter7));
  inv1  gate1589(.a(N892), .O(gate261inter8));
  nand2 gate1590(.a(gate261inter8), .b(gate261inter7), .O(gate261inter9));
  nand2 gate1591(.a(s_101), .b(gate261inter3), .O(gate261inter10));
  nor2  gate1592(.a(gate261inter10), .b(gate261inter9), .O(gate261inter11));
  nor2  gate1593(.a(gate261inter11), .b(gate261inter6), .O(gate261inter12));
  nand2 gate1594(.a(gate261inter12), .b(gate261inter1), .O(N1160));
inv1 gate262( .a(N998), .O(N1161) );
nand2 gate263( .a(N1067), .b(N1068), .O(N1162) );
inv1 gate264( .a(N899), .O(N1163) );
buf1 gate265( .a(N899), .O(N1164) );
inv1 gate266( .a(N903), .O(N1167) );
buf1 gate267( .a(N903), .O(N1168) );
nand2 gate268( .a(N921), .b(N923), .O(N1171) );
nand2 gate269( .a(N922), .b(N923), .O(N1188) );
inv1 gate270( .a(N1010), .O(N1205) );
nand2 gate271( .a(N1010), .b(N938), .O(N1206) );
inv1 gate272( .a(N1013), .O(N1207) );
nand2 gate273( .a(N1013), .b(N942), .O(N1208) );
inv1 gate274( .a(N1016), .O(N1209) );
nand2 gate275( .a(N1016), .b(N946), .O(N1210) );
inv1 gate276( .a(N1019), .O(N1211) );
nand2 gate277( .a(N1019), .b(N950), .O(N1212) );
inv1 gate278( .a(N1022), .O(N1213) );
nand2 gate279( .a(N1022), .b(N954), .O(N1214) );
inv1 gate280( .a(N1025), .O(N1215) );
nand2 gate281( .a(N1025), .b(N958), .O(N1216) );
inv1 gate282( .a(N1028), .O(N1217) );
inv1 gate283( .a(N959), .O(N1218) );
inv1 gate284( .a(N1031), .O(N1219) );
inv1 gate285( .a(N1034), .O(N1220) );
nand2 gate286( .a(N1034), .b(N968), .O(N1221) );
inv1 gate287( .a(N965), .O(N1222) );
inv1 gate288( .a(N1037), .O(N1223) );
nand2 gate289( .a(N1037), .b(N972), .O(N1224) );
inv1 gate290( .a(N1040), .O(N1225) );
nand2 gate291( .a(N1040), .b(N976), .O(N1226) );
inv1 gate292( .a(N973), .O(N1227) );
inv1 gate293( .a(N1043), .O(N1228) );

  xor2  gate993(.a(N980), .b(N1043), .O(gate294inter0));
  nand2 gate994(.a(gate294inter0), .b(s_16), .O(gate294inter1));
  and2  gate995(.a(N980), .b(N1043), .O(gate294inter2));
  inv1  gate996(.a(s_16), .O(gate294inter3));
  inv1  gate997(.a(s_17), .O(gate294inter4));
  nand2 gate998(.a(gate294inter4), .b(gate294inter3), .O(gate294inter5));
  nor2  gate999(.a(gate294inter5), .b(gate294inter2), .O(gate294inter6));
  inv1  gate1000(.a(N1043), .O(gate294inter7));
  inv1  gate1001(.a(N980), .O(gate294inter8));
  nand2 gate1002(.a(gate294inter8), .b(gate294inter7), .O(gate294inter9));
  nand2 gate1003(.a(s_17), .b(gate294inter3), .O(gate294inter10));
  nor2  gate1004(.a(gate294inter10), .b(gate294inter9), .O(gate294inter11));
  nor2  gate1005(.a(gate294inter11), .b(gate294inter6), .O(gate294inter12));
  nand2 gate1006(.a(gate294inter12), .b(gate294inter1), .O(N1229));
inv1 gate295( .a(N981), .O(N1230) );
nand2 gate296( .a(N981), .b(N984), .O(N1231) );
nand2 gate297( .a(N1119), .b(N1120), .O(N1232) );

  xor2  gate1455(.a(N1122), .b(N1121), .O(gate298inter0));
  nand2 gate1456(.a(gate298inter0), .b(s_82), .O(gate298inter1));
  and2  gate1457(.a(N1122), .b(N1121), .O(gate298inter2));
  inv1  gate1458(.a(s_82), .O(gate298inter3));
  inv1  gate1459(.a(s_83), .O(gate298inter4));
  nand2 gate1460(.a(gate298inter4), .b(gate298inter3), .O(gate298inter5));
  nor2  gate1461(.a(gate298inter5), .b(gate298inter2), .O(gate298inter6));
  inv1  gate1462(.a(N1121), .O(gate298inter7));
  inv1  gate1463(.a(N1122), .O(gate298inter8));
  nand2 gate1464(.a(gate298inter8), .b(gate298inter7), .O(gate298inter9));
  nand2 gate1465(.a(s_83), .b(gate298inter3), .O(gate298inter10));
  nor2  gate1466(.a(gate298inter10), .b(gate298inter9), .O(gate298inter11));
  nor2  gate1467(.a(gate298inter11), .b(gate298inter6), .O(gate298inter12));
  nand2 gate1468(.a(gate298inter12), .b(gate298inter1), .O(N1235));
inv1 gate299( .a(N1046), .O(N1238) );
nand2 gate300( .a(N1046), .b(N997), .O(N1239) );
inv1 gate301( .a(N994), .O(N1240) );
inv1 gate302( .a(N1049), .O(N1241) );
nand2 gate303( .a(N1049), .b(N1001), .O(N1242) );
nand2 gate304( .a(N1128), .b(N1129), .O(N1243) );
nand2 gate305( .a(N1130), .b(N1131), .O(N1246) );
nand2 gate306( .a(N1132), .b(N1133), .O(N1249) );
buf1 gate307( .a(N907), .O(N1252) );
buf1 gate308( .a(N907), .O(N1255) );
buf1 gate309( .a(N910), .O(N1258) );
buf1 gate310( .a(N910), .O(N1261) );
inv1 gate311( .a(N1150), .O(N1264) );
nand2 gate312( .a(N631), .b(N1159), .O(N1267) );
nand2 gate313( .a(N688), .b(N1205), .O(N1309) );
nand2 gate314( .a(N691), .b(N1207), .O(N1310) );
nand2 gate315( .a(N694), .b(N1209), .O(N1311) );
nand2 gate316( .a(N697), .b(N1211), .O(N1312) );
nand2 gate317( .a(N700), .b(N1213), .O(N1313) );
nand2 gate318( .a(N703), .b(N1215), .O(N1314) );
nand2 gate319( .a(N706), .b(N1220), .O(N1315) );
nand2 gate320( .a(N709), .b(N1223), .O(N1316) );

  xor2  gate937(.a(N1225), .b(N712), .O(gate321inter0));
  nand2 gate938(.a(gate321inter0), .b(s_8), .O(gate321inter1));
  and2  gate939(.a(N1225), .b(N712), .O(gate321inter2));
  inv1  gate940(.a(s_8), .O(gate321inter3));
  inv1  gate941(.a(s_9), .O(gate321inter4));
  nand2 gate942(.a(gate321inter4), .b(gate321inter3), .O(gate321inter5));
  nor2  gate943(.a(gate321inter5), .b(gate321inter2), .O(gate321inter6));
  inv1  gate944(.a(N712), .O(gate321inter7));
  inv1  gate945(.a(N1225), .O(gate321inter8));
  nand2 gate946(.a(gate321inter8), .b(gate321inter7), .O(gate321inter9));
  nand2 gate947(.a(s_9), .b(gate321inter3), .O(gate321inter10));
  nor2  gate948(.a(gate321inter10), .b(gate321inter9), .O(gate321inter11));
  nor2  gate949(.a(gate321inter11), .b(gate321inter6), .O(gate321inter12));
  nand2 gate950(.a(gate321inter12), .b(gate321inter1), .O(N1317));
nand2 gate322( .a(N715), .b(N1228), .O(N1318) );
inv1 gate323( .a(N1158), .O(N1319) );
nand2 gate324( .a(N628), .b(N1230), .O(N1322) );
nand2 gate325( .a(N730), .b(N1238), .O(N1327) );
nand2 gate326( .a(N733), .b(N1241), .O(N1328) );
inv1 gate327( .a(N1162), .O(N1334) );
nand2 gate328( .a(N1267), .b(N1160), .O(N1344) );
nand2 gate329( .a(N1249), .b(N894), .O(N1345) );
inv1 gate330( .a(N1249), .O(N1346) );
inv1 gate331( .a(N1255), .O(N1348) );
inv1 gate332( .a(N1252), .O(N1349) );
inv1 gate333( .a(N1261), .O(N1350) );
inv1 gate334( .a(N1258), .O(N1351) );

  xor2  gate1147(.a(N1206), .b(N1309), .O(gate335inter0));
  nand2 gate1148(.a(gate335inter0), .b(s_38), .O(gate335inter1));
  and2  gate1149(.a(N1206), .b(N1309), .O(gate335inter2));
  inv1  gate1150(.a(s_38), .O(gate335inter3));
  inv1  gate1151(.a(s_39), .O(gate335inter4));
  nand2 gate1152(.a(gate335inter4), .b(gate335inter3), .O(gate335inter5));
  nor2  gate1153(.a(gate335inter5), .b(gate335inter2), .O(gate335inter6));
  inv1  gate1154(.a(N1309), .O(gate335inter7));
  inv1  gate1155(.a(N1206), .O(gate335inter8));
  nand2 gate1156(.a(gate335inter8), .b(gate335inter7), .O(gate335inter9));
  nand2 gate1157(.a(s_39), .b(gate335inter3), .O(gate335inter10));
  nor2  gate1158(.a(gate335inter10), .b(gate335inter9), .O(gate335inter11));
  nor2  gate1159(.a(gate335inter11), .b(gate335inter6), .O(gate335inter12));
  nand2 gate1160(.a(gate335inter12), .b(gate335inter1), .O(N1352));
nand2 gate336( .a(N1310), .b(N1208), .O(N1355) );

  xor2  gate1791(.a(N1210), .b(N1311), .O(gate337inter0));
  nand2 gate1792(.a(gate337inter0), .b(s_130), .O(gate337inter1));
  and2  gate1793(.a(N1210), .b(N1311), .O(gate337inter2));
  inv1  gate1794(.a(s_130), .O(gate337inter3));
  inv1  gate1795(.a(s_131), .O(gate337inter4));
  nand2 gate1796(.a(gate337inter4), .b(gate337inter3), .O(gate337inter5));
  nor2  gate1797(.a(gate337inter5), .b(gate337inter2), .O(gate337inter6));
  inv1  gate1798(.a(N1311), .O(gate337inter7));
  inv1  gate1799(.a(N1210), .O(gate337inter8));
  nand2 gate1800(.a(gate337inter8), .b(gate337inter7), .O(gate337inter9));
  nand2 gate1801(.a(s_131), .b(gate337inter3), .O(gate337inter10));
  nor2  gate1802(.a(gate337inter10), .b(gate337inter9), .O(gate337inter11));
  nor2  gate1803(.a(gate337inter11), .b(gate337inter6), .O(gate337inter12));
  nand2 gate1804(.a(gate337inter12), .b(gate337inter1), .O(N1358));

  xor2  gate1049(.a(N1212), .b(N1312), .O(gate338inter0));
  nand2 gate1050(.a(gate338inter0), .b(s_24), .O(gate338inter1));
  and2  gate1051(.a(N1212), .b(N1312), .O(gate338inter2));
  inv1  gate1052(.a(s_24), .O(gate338inter3));
  inv1  gate1053(.a(s_25), .O(gate338inter4));
  nand2 gate1054(.a(gate338inter4), .b(gate338inter3), .O(gate338inter5));
  nor2  gate1055(.a(gate338inter5), .b(gate338inter2), .O(gate338inter6));
  inv1  gate1056(.a(N1312), .O(gate338inter7));
  inv1  gate1057(.a(N1212), .O(gate338inter8));
  nand2 gate1058(.a(gate338inter8), .b(gate338inter7), .O(gate338inter9));
  nand2 gate1059(.a(s_25), .b(gate338inter3), .O(gate338inter10));
  nor2  gate1060(.a(gate338inter10), .b(gate338inter9), .O(gate338inter11));
  nor2  gate1061(.a(gate338inter11), .b(gate338inter6), .O(gate338inter12));
  nand2 gate1062(.a(gate338inter12), .b(gate338inter1), .O(N1361));

  xor2  gate1035(.a(N1214), .b(N1313), .O(gate339inter0));
  nand2 gate1036(.a(gate339inter0), .b(s_22), .O(gate339inter1));
  and2  gate1037(.a(N1214), .b(N1313), .O(gate339inter2));
  inv1  gate1038(.a(s_22), .O(gate339inter3));
  inv1  gate1039(.a(s_23), .O(gate339inter4));
  nand2 gate1040(.a(gate339inter4), .b(gate339inter3), .O(gate339inter5));
  nor2  gate1041(.a(gate339inter5), .b(gate339inter2), .O(gate339inter6));
  inv1  gate1042(.a(N1313), .O(gate339inter7));
  inv1  gate1043(.a(N1214), .O(gate339inter8));
  nand2 gate1044(.a(gate339inter8), .b(gate339inter7), .O(gate339inter9));
  nand2 gate1045(.a(s_23), .b(gate339inter3), .O(gate339inter10));
  nor2  gate1046(.a(gate339inter10), .b(gate339inter9), .O(gate339inter11));
  nor2  gate1047(.a(gate339inter11), .b(gate339inter6), .O(gate339inter12));
  nand2 gate1048(.a(gate339inter12), .b(gate339inter1), .O(N1364));
nand2 gate340( .a(N1314), .b(N1216), .O(N1367) );
nand2 gate341( .a(N1315), .b(N1221), .O(N1370) );
nand2 gate342( .a(N1316), .b(N1224), .O(N1373) );

  xor2  gate1777(.a(N1226), .b(N1317), .O(gate343inter0));
  nand2 gate1778(.a(gate343inter0), .b(s_128), .O(gate343inter1));
  and2  gate1779(.a(N1226), .b(N1317), .O(gate343inter2));
  inv1  gate1780(.a(s_128), .O(gate343inter3));
  inv1  gate1781(.a(s_129), .O(gate343inter4));
  nand2 gate1782(.a(gate343inter4), .b(gate343inter3), .O(gate343inter5));
  nor2  gate1783(.a(gate343inter5), .b(gate343inter2), .O(gate343inter6));
  inv1  gate1784(.a(N1317), .O(gate343inter7));
  inv1  gate1785(.a(N1226), .O(gate343inter8));
  nand2 gate1786(.a(gate343inter8), .b(gate343inter7), .O(gate343inter9));
  nand2 gate1787(.a(s_129), .b(gate343inter3), .O(gate343inter10));
  nor2  gate1788(.a(gate343inter10), .b(gate343inter9), .O(gate343inter11));
  nor2  gate1789(.a(gate343inter11), .b(gate343inter6), .O(gate343inter12));
  nand2 gate1790(.a(gate343inter12), .b(gate343inter1), .O(N1376));
nand2 gate344( .a(N1318), .b(N1229), .O(N1379) );
nand2 gate345( .a(N1322), .b(N1231), .O(N1383) );
inv1 gate346( .a(N1232), .O(N1386) );
nand2 gate347( .a(N1232), .b(N990), .O(N1387) );
inv1 gate348( .a(N1235), .O(N1388) );
nand2 gate349( .a(N1235), .b(N993), .O(N1389) );

  xor2  gate1063(.a(N1239), .b(N1327), .O(gate350inter0));
  nand2 gate1064(.a(gate350inter0), .b(s_26), .O(gate350inter1));
  and2  gate1065(.a(N1239), .b(N1327), .O(gate350inter2));
  inv1  gate1066(.a(s_26), .O(gate350inter3));
  inv1  gate1067(.a(s_27), .O(gate350inter4));
  nand2 gate1068(.a(gate350inter4), .b(gate350inter3), .O(gate350inter5));
  nor2  gate1069(.a(gate350inter5), .b(gate350inter2), .O(gate350inter6));
  inv1  gate1070(.a(N1327), .O(gate350inter7));
  inv1  gate1071(.a(N1239), .O(gate350inter8));
  nand2 gate1072(.a(gate350inter8), .b(gate350inter7), .O(gate350inter9));
  nand2 gate1073(.a(s_27), .b(gate350inter3), .O(gate350inter10));
  nor2  gate1074(.a(gate350inter10), .b(gate350inter9), .O(gate350inter11));
  nor2  gate1075(.a(gate350inter11), .b(gate350inter6), .O(gate350inter12));
  nand2 gate1076(.a(gate350inter12), .b(gate350inter1), .O(N1390));
nand2 gate351( .a(N1328), .b(N1242), .O(N1393) );
inv1 gate352( .a(N1243), .O(N1396) );
nand2 gate353( .a(N1243), .b(N1004), .O(N1397) );
inv1 gate354( .a(N1246), .O(N1398) );
nand2 gate355( .a(N1246), .b(N1007), .O(N1399) );
inv1 gate356( .a(N1319), .O(N1409) );
nand2 gate357( .a(N649), .b(N1346), .O(N1412) );
inv1 gate358( .a(N1334), .O(N1413) );
buf1 gate359( .a(N1264), .O(N1416) );
buf1 gate360( .a(N1264), .O(N1419) );
nand2 gate361( .a(N634), .b(N1386), .O(N1433) );
nand2 gate362( .a(N637), .b(N1388), .O(N1434) );
nand2 gate363( .a(N640), .b(N1396), .O(N1438) );
nand2 gate364( .a(N646), .b(N1398), .O(N1439) );
inv1 gate365( .a(N1344), .O(N1440) );
nand2 gate366( .a(N1355), .b(N1148), .O(N1443) );
inv1 gate367( .a(N1355), .O(N1444) );
nand2 gate368( .a(N1352), .b(N1149), .O(N1445) );
inv1 gate369( .a(N1352), .O(N1446) );
nand2 gate370( .a(N1358), .b(N1151), .O(N1447) );
inv1 gate371( .a(N1358), .O(N1448) );
nand2 gate372( .a(N1361), .b(N1152), .O(N1451) );
inv1 gate373( .a(N1361), .O(N1452) );
nand2 gate374( .a(N1367), .b(N1153), .O(N1453) );
inv1 gate375( .a(N1367), .O(N1454) );

  xor2  gate1105(.a(N1154), .b(N1364), .O(gate376inter0));
  nand2 gate1106(.a(gate376inter0), .b(s_32), .O(gate376inter1));
  and2  gate1107(.a(N1154), .b(N1364), .O(gate376inter2));
  inv1  gate1108(.a(s_32), .O(gate376inter3));
  inv1  gate1109(.a(s_33), .O(gate376inter4));
  nand2 gate1110(.a(gate376inter4), .b(gate376inter3), .O(gate376inter5));
  nor2  gate1111(.a(gate376inter5), .b(gate376inter2), .O(gate376inter6));
  inv1  gate1112(.a(N1364), .O(gate376inter7));
  inv1  gate1113(.a(N1154), .O(gate376inter8));
  nand2 gate1114(.a(gate376inter8), .b(gate376inter7), .O(gate376inter9));
  nand2 gate1115(.a(s_33), .b(gate376inter3), .O(gate376inter10));
  nor2  gate1116(.a(gate376inter10), .b(gate376inter9), .O(gate376inter11));
  nor2  gate1117(.a(gate376inter11), .b(gate376inter6), .O(gate376inter12));
  nand2 gate1118(.a(gate376inter12), .b(gate376inter1), .O(N1455));
inv1 gate377( .a(N1364), .O(N1456) );
nand2 gate378( .a(N1373), .b(N1156), .O(N1457) );
inv1 gate379( .a(N1373), .O(N1458) );
nand2 gate380( .a(N1379), .b(N1157), .O(N1459) );
inv1 gate381( .a(N1379), .O(N1460) );
inv1 gate382( .a(N1383), .O(N1461) );
nand2 gate383( .a(N1393), .b(N1161), .O(N1462) );
inv1 gate384( .a(N1393), .O(N1463) );

  xor2  gate1693(.a(N1412), .b(N1345), .O(gate385inter0));
  nand2 gate1694(.a(gate385inter0), .b(s_116), .O(gate385inter1));
  and2  gate1695(.a(N1412), .b(N1345), .O(gate385inter2));
  inv1  gate1696(.a(s_116), .O(gate385inter3));
  inv1  gate1697(.a(s_117), .O(gate385inter4));
  nand2 gate1698(.a(gate385inter4), .b(gate385inter3), .O(gate385inter5));
  nor2  gate1699(.a(gate385inter5), .b(gate385inter2), .O(gate385inter6));
  inv1  gate1700(.a(N1345), .O(gate385inter7));
  inv1  gate1701(.a(N1412), .O(gate385inter8));
  nand2 gate1702(.a(gate385inter8), .b(gate385inter7), .O(gate385inter9));
  nand2 gate1703(.a(s_117), .b(gate385inter3), .O(gate385inter10));
  nor2  gate1704(.a(gate385inter10), .b(gate385inter9), .O(gate385inter11));
  nor2  gate1705(.a(gate385inter11), .b(gate385inter6), .O(gate385inter12));
  nand2 gate1706(.a(gate385inter12), .b(gate385inter1), .O(N1464));
inv1 gate386( .a(N1370), .O(N1468) );

  xor2  gate1553(.a(N1222), .b(N1370), .O(gate387inter0));
  nand2 gate1554(.a(gate387inter0), .b(s_96), .O(gate387inter1));
  and2  gate1555(.a(N1222), .b(N1370), .O(gate387inter2));
  inv1  gate1556(.a(s_96), .O(gate387inter3));
  inv1  gate1557(.a(s_97), .O(gate387inter4));
  nand2 gate1558(.a(gate387inter4), .b(gate387inter3), .O(gate387inter5));
  nor2  gate1559(.a(gate387inter5), .b(gate387inter2), .O(gate387inter6));
  inv1  gate1560(.a(N1370), .O(gate387inter7));
  inv1  gate1561(.a(N1222), .O(gate387inter8));
  nand2 gate1562(.a(gate387inter8), .b(gate387inter7), .O(gate387inter9));
  nand2 gate1563(.a(s_97), .b(gate387inter3), .O(gate387inter10));
  nor2  gate1564(.a(gate387inter10), .b(gate387inter9), .O(gate387inter11));
  nor2  gate1565(.a(gate387inter11), .b(gate387inter6), .O(gate387inter12));
  nand2 gate1566(.a(gate387inter12), .b(gate387inter1), .O(N1469));
inv1 gate388( .a(N1376), .O(N1470) );
nand2 gate389( .a(N1376), .b(N1227), .O(N1471) );
nand2 gate390( .a(N1387), .b(N1433), .O(N1472) );
inv1 gate391( .a(N1390), .O(N1475) );
nand2 gate392( .a(N1390), .b(N1240), .O(N1476) );
nand2 gate393( .a(N1389), .b(N1434), .O(N1478) );
nand2 gate394( .a(N1399), .b(N1439), .O(N1481) );
nand2 gate395( .a(N1397), .b(N1438), .O(N1484) );

  xor2  gate1231(.a(N1444), .b(N939), .O(gate396inter0));
  nand2 gate1232(.a(gate396inter0), .b(s_50), .O(gate396inter1));
  and2  gate1233(.a(N1444), .b(N939), .O(gate396inter2));
  inv1  gate1234(.a(s_50), .O(gate396inter3));
  inv1  gate1235(.a(s_51), .O(gate396inter4));
  nand2 gate1236(.a(gate396inter4), .b(gate396inter3), .O(gate396inter5));
  nor2  gate1237(.a(gate396inter5), .b(gate396inter2), .O(gate396inter6));
  inv1  gate1238(.a(N939), .O(gate396inter7));
  inv1  gate1239(.a(N1444), .O(gate396inter8));
  nand2 gate1240(.a(gate396inter8), .b(gate396inter7), .O(gate396inter9));
  nand2 gate1241(.a(s_51), .b(gate396inter3), .O(gate396inter10));
  nor2  gate1242(.a(gate396inter10), .b(gate396inter9), .O(gate396inter11));
  nor2  gate1243(.a(gate396inter11), .b(gate396inter6), .O(gate396inter12));
  nand2 gate1244(.a(gate396inter12), .b(gate396inter1), .O(N1487));
nand2 gate397( .a(N935), .b(N1446), .O(N1488) );
nand2 gate398( .a(N943), .b(N1448), .O(N1489) );
inv1 gate399( .a(N1419), .O(N1490) );
inv1 gate400( .a(N1416), .O(N1491) );

  xor2  gate1483(.a(N1452), .b(N947), .O(gate401inter0));
  nand2 gate1484(.a(gate401inter0), .b(s_86), .O(gate401inter1));
  and2  gate1485(.a(N1452), .b(N947), .O(gate401inter2));
  inv1  gate1486(.a(s_86), .O(gate401inter3));
  inv1  gate1487(.a(s_87), .O(gate401inter4));
  nand2 gate1488(.a(gate401inter4), .b(gate401inter3), .O(gate401inter5));
  nor2  gate1489(.a(gate401inter5), .b(gate401inter2), .O(gate401inter6));
  inv1  gate1490(.a(N947), .O(gate401inter7));
  inv1  gate1491(.a(N1452), .O(gate401inter8));
  nand2 gate1492(.a(gate401inter8), .b(gate401inter7), .O(gate401inter9));
  nand2 gate1493(.a(s_87), .b(gate401inter3), .O(gate401inter10));
  nor2  gate1494(.a(gate401inter10), .b(gate401inter9), .O(gate401inter11));
  nor2  gate1495(.a(gate401inter11), .b(gate401inter6), .O(gate401inter12));
  nand2 gate1496(.a(gate401inter12), .b(gate401inter1), .O(N1492));
nand2 gate402( .a(N955), .b(N1454), .O(N1493) );
nand2 gate403( .a(N951), .b(N1456), .O(N1494) );
nand2 gate404( .a(N969), .b(N1458), .O(N1495) );

  xor2  gate1623(.a(N1460), .b(N977), .O(gate405inter0));
  nand2 gate1624(.a(gate405inter0), .b(s_106), .O(gate405inter1));
  and2  gate1625(.a(N1460), .b(N977), .O(gate405inter2));
  inv1  gate1626(.a(s_106), .O(gate405inter3));
  inv1  gate1627(.a(s_107), .O(gate405inter4));
  nand2 gate1628(.a(gate405inter4), .b(gate405inter3), .O(gate405inter5));
  nor2  gate1629(.a(gate405inter5), .b(gate405inter2), .O(gate405inter6));
  inv1  gate1630(.a(N977), .O(gate405inter7));
  inv1  gate1631(.a(N1460), .O(gate405inter8));
  nand2 gate1632(.a(gate405inter8), .b(gate405inter7), .O(gate405inter9));
  nand2 gate1633(.a(s_107), .b(gate405inter3), .O(gate405inter10));
  nor2  gate1634(.a(gate405inter10), .b(gate405inter9), .O(gate405inter11));
  nor2  gate1635(.a(gate405inter11), .b(gate405inter6), .O(gate405inter12));
  nand2 gate1636(.a(gate405inter12), .b(gate405inter1), .O(N1496));

  xor2  gate1525(.a(N1463), .b(N998), .O(gate406inter0));
  nand2 gate1526(.a(gate406inter0), .b(s_92), .O(gate406inter1));
  and2  gate1527(.a(N1463), .b(N998), .O(gate406inter2));
  inv1  gate1528(.a(s_92), .O(gate406inter3));
  inv1  gate1529(.a(s_93), .O(gate406inter4));
  nand2 gate1530(.a(gate406inter4), .b(gate406inter3), .O(gate406inter5));
  nor2  gate1531(.a(gate406inter5), .b(gate406inter2), .O(gate406inter6));
  inv1  gate1532(.a(N998), .O(gate406inter7));
  inv1  gate1533(.a(N1463), .O(gate406inter8));
  nand2 gate1534(.a(gate406inter8), .b(gate406inter7), .O(gate406inter9));
  nand2 gate1535(.a(s_93), .b(gate406inter3), .O(gate406inter10));
  nor2  gate1536(.a(gate406inter10), .b(gate406inter9), .O(gate406inter11));
  nor2  gate1537(.a(gate406inter11), .b(gate406inter6), .O(gate406inter12));
  nand2 gate1538(.a(gate406inter12), .b(gate406inter1), .O(N1498));
inv1 gate407( .a(N1440), .O(N1499) );
nand2 gate408( .a(N965), .b(N1468), .O(N1500) );
nand2 gate409( .a(N973), .b(N1470), .O(N1501) );
nand2 gate410( .a(N994), .b(N1475), .O(N1504) );
inv1 gate411( .a(N1464), .O(N1510) );

  xor2  gate1091(.a(N1487), .b(N1443), .O(gate412inter0));
  nand2 gate1092(.a(gate412inter0), .b(s_30), .O(gate412inter1));
  and2  gate1093(.a(N1487), .b(N1443), .O(gate412inter2));
  inv1  gate1094(.a(s_30), .O(gate412inter3));
  inv1  gate1095(.a(s_31), .O(gate412inter4));
  nand2 gate1096(.a(gate412inter4), .b(gate412inter3), .O(gate412inter5));
  nor2  gate1097(.a(gate412inter5), .b(gate412inter2), .O(gate412inter6));
  inv1  gate1098(.a(N1443), .O(gate412inter7));
  inv1  gate1099(.a(N1487), .O(gate412inter8));
  nand2 gate1100(.a(gate412inter8), .b(gate412inter7), .O(gate412inter9));
  nand2 gate1101(.a(s_31), .b(gate412inter3), .O(gate412inter10));
  nor2  gate1102(.a(gate412inter10), .b(gate412inter9), .O(gate412inter11));
  nor2  gate1103(.a(gate412inter11), .b(gate412inter6), .O(gate412inter12));
  nand2 gate1104(.a(gate412inter12), .b(gate412inter1), .O(N1513));
nand2 gate413( .a(N1445), .b(N1488), .O(N1514) );
nand2 gate414( .a(N1447), .b(N1489), .O(N1517) );
nand2 gate415( .a(N1451), .b(N1492), .O(N1520) );
nand2 gate416( .a(N1453), .b(N1493), .O(N1521) );
nand2 gate417( .a(N1455), .b(N1494), .O(N1522) );

  xor2  gate1301(.a(N1495), .b(N1457), .O(gate418inter0));
  nand2 gate1302(.a(gate418inter0), .b(s_60), .O(gate418inter1));
  and2  gate1303(.a(N1495), .b(N1457), .O(gate418inter2));
  inv1  gate1304(.a(s_60), .O(gate418inter3));
  inv1  gate1305(.a(s_61), .O(gate418inter4));
  nand2 gate1306(.a(gate418inter4), .b(gate418inter3), .O(gate418inter5));
  nor2  gate1307(.a(gate418inter5), .b(gate418inter2), .O(gate418inter6));
  inv1  gate1308(.a(N1457), .O(gate418inter7));
  inv1  gate1309(.a(N1495), .O(gate418inter8));
  nand2 gate1310(.a(gate418inter8), .b(gate418inter7), .O(gate418inter9));
  nand2 gate1311(.a(s_61), .b(gate418inter3), .O(gate418inter10));
  nor2  gate1312(.a(gate418inter10), .b(gate418inter9), .O(gate418inter11));
  nor2  gate1313(.a(gate418inter11), .b(gate418inter6), .O(gate418inter12));
  nand2 gate1314(.a(gate418inter12), .b(gate418inter1), .O(N1526));

  xor2  gate1203(.a(N1496), .b(N1459), .O(gate419inter0));
  nand2 gate1204(.a(gate419inter0), .b(s_46), .O(gate419inter1));
  and2  gate1205(.a(N1496), .b(N1459), .O(gate419inter2));
  inv1  gate1206(.a(s_46), .O(gate419inter3));
  inv1  gate1207(.a(s_47), .O(gate419inter4));
  nand2 gate1208(.a(gate419inter4), .b(gate419inter3), .O(gate419inter5));
  nor2  gate1209(.a(gate419inter5), .b(gate419inter2), .O(gate419inter6));
  inv1  gate1210(.a(N1459), .O(gate419inter7));
  inv1  gate1211(.a(N1496), .O(gate419inter8));
  nand2 gate1212(.a(gate419inter8), .b(gate419inter7), .O(gate419inter9));
  nand2 gate1213(.a(s_47), .b(gate419inter3), .O(gate419inter10));
  nor2  gate1214(.a(gate419inter10), .b(gate419inter9), .O(gate419inter11));
  nor2  gate1215(.a(gate419inter11), .b(gate419inter6), .O(gate419inter12));
  nand2 gate1216(.a(gate419inter12), .b(gate419inter1), .O(N1527));
inv1 gate420( .a(N1472), .O(N1528) );
nand2 gate421( .a(N1462), .b(N1498), .O(N1529) );
inv1 gate422( .a(N1478), .O(N1530) );
inv1 gate423( .a(N1481), .O(N1531) );
inv1 gate424( .a(N1484), .O(N1532) );
nand2 gate425( .a(N1471), .b(N1501), .O(N1534) );
nand2 gate426( .a(N1469), .b(N1500), .O(N1537) );
nand2 gate427( .a(N1476), .b(N1504), .O(N1540) );
inv1 gate428( .a(N1513), .O(N1546) );
inv1 gate429( .a(N1521), .O(N1554) );
inv1 gate430( .a(N1526), .O(N1557) );
inv1 gate431( .a(N1520), .O(N1561) );
nand2 gate432( .a(N1484), .b(N1531), .O(N1567) );
nand2 gate433( .a(N1481), .b(N1532), .O(N1568) );
inv1 gate434( .a(N1510), .O(N1569) );
inv1 gate435( .a(N1527), .O(N1571) );
inv1 gate436( .a(N1529), .O(N1576) );
buf1 gate437( .a(N1522), .O(N1588) );
inv1 gate438( .a(N1534), .O(N1591) );
inv1 gate439( .a(N1537), .O(N1593) );
nand2 gate440( .a(N1540), .b(N1530), .O(N1594) );
inv1 gate441( .a(N1540), .O(N1595) );
nand2 gate442( .a(N1567), .b(N1568), .O(N1596) );
buf1 gate443( .a(N1517), .O(N1600) );
buf1 gate444( .a(N1517), .O(N1603) );
buf1 gate445( .a(N1522), .O(N1606) );
buf1 gate446( .a(N1522), .O(N1609) );
buf1 gate447( .a(N1514), .O(N1612) );
buf1 gate448( .a(N1514), .O(N1615) );
buf1 gate449( .a(N1557), .O(N1620) );
buf1 gate450( .a(N1554), .O(N1623) );
inv1 gate451( .a(N1571), .O(N1635) );
nand2 gate452( .a(N1478), .b(N1595), .O(N1636) );
nand2 gate453( .a(N1576), .b(N1569), .O(N1638) );
inv1 gate454( .a(N1576), .O(N1639) );
buf1 gate455( .a(N1561), .O(N1640) );
buf1 gate456( .a(N1561), .O(N1643) );
buf1 gate457( .a(N1546), .O(N1647) );
buf1 gate458( .a(N1546), .O(N1651) );
buf1 gate459( .a(N1554), .O(N1658) );
buf1 gate460( .a(N1557), .O(N1661) );
buf1 gate461( .a(N1557), .O(N1664) );
nand2 gate462( .a(N1596), .b(N893), .O(N1671) );
inv1 gate463( .a(N1596), .O(N1672) );
inv1 gate464( .a(N1600), .O(N1675) );
inv1 gate465( .a(N1603), .O(N1677) );
nand2 gate466( .a(N1606), .b(N1217), .O(N1678) );
inv1 gate467( .a(N1606), .O(N1679) );
nand2 gate468( .a(N1609), .b(N1219), .O(N1680) );
inv1 gate469( .a(N1609), .O(N1681) );
inv1 gate470( .a(N1612), .O(N1682) );
inv1 gate471( .a(N1615), .O(N1683) );
nand2 gate472( .a(N1594), .b(N1636), .O(N1685) );
nand2 gate473( .a(N1510), .b(N1639), .O(N1688) );
buf1 gate474( .a(N1588), .O(N1697) );
buf1 gate475( .a(N1588), .O(N1701) );
nand2 gate476( .a(N643), .b(N1672), .O(N1706) );
inv1 gate477( .a(N1643), .O(N1707) );

  xor2  gate1133(.a(N1675), .b(N1647), .O(gate478inter0));
  nand2 gate1134(.a(gate478inter0), .b(s_36), .O(gate478inter1));
  and2  gate1135(.a(N1675), .b(N1647), .O(gate478inter2));
  inv1  gate1136(.a(s_36), .O(gate478inter3));
  inv1  gate1137(.a(s_37), .O(gate478inter4));
  nand2 gate1138(.a(gate478inter4), .b(gate478inter3), .O(gate478inter5));
  nor2  gate1139(.a(gate478inter5), .b(gate478inter2), .O(gate478inter6));
  inv1  gate1140(.a(N1647), .O(gate478inter7));
  inv1  gate1141(.a(N1675), .O(gate478inter8));
  nand2 gate1142(.a(gate478inter8), .b(gate478inter7), .O(gate478inter9));
  nand2 gate1143(.a(s_37), .b(gate478inter3), .O(gate478inter10));
  nor2  gate1144(.a(gate478inter10), .b(gate478inter9), .O(gate478inter11));
  nor2  gate1145(.a(gate478inter11), .b(gate478inter6), .O(gate478inter12));
  nand2 gate1146(.a(gate478inter12), .b(gate478inter1), .O(N1708));
inv1 gate479( .a(N1647), .O(N1709) );
nand2 gate480( .a(N1651), .b(N1677), .O(N1710) );
inv1 gate481( .a(N1651), .O(N1711) );
nand2 gate482( .a(N1028), .b(N1679), .O(N1712) );
nand2 gate483( .a(N1031), .b(N1681), .O(N1713) );
buf1 gate484( .a(N1620), .O(N1714) );
buf1 gate485( .a(N1620), .O(N1717) );
nand2 gate486( .a(N1658), .b(N1593), .O(N1720) );
inv1 gate487( .a(N1658), .O(N1721) );
nand2 gate488( .a(N1638), .b(N1688), .O(N1723) );
inv1 gate489( .a(N1661), .O(N1727) );
inv1 gate490( .a(N1640), .O(N1728) );
inv1 gate491( .a(N1664), .O(N1730) );
buf1 gate492( .a(N1623), .O(N1731) );
buf1 gate493( .a(N1623), .O(N1734) );
nand2 gate494( .a(N1685), .b(N1528), .O(N1740) );
inv1 gate495( .a(N1685), .O(N1741) );

  xor2  gate1217(.a(N1706), .b(N1671), .O(gate496inter0));
  nand2 gate1218(.a(gate496inter0), .b(s_48), .O(gate496inter1));
  and2  gate1219(.a(N1706), .b(N1671), .O(gate496inter2));
  inv1  gate1220(.a(s_48), .O(gate496inter3));
  inv1  gate1221(.a(s_49), .O(gate496inter4));
  nand2 gate1222(.a(gate496inter4), .b(gate496inter3), .O(gate496inter5));
  nor2  gate1223(.a(gate496inter5), .b(gate496inter2), .O(gate496inter6));
  inv1  gate1224(.a(N1671), .O(gate496inter7));
  inv1  gate1225(.a(N1706), .O(gate496inter8));
  nand2 gate1226(.a(gate496inter8), .b(gate496inter7), .O(gate496inter9));
  nand2 gate1227(.a(s_49), .b(gate496inter3), .O(gate496inter10));
  nor2  gate1228(.a(gate496inter10), .b(gate496inter9), .O(gate496inter11));
  nor2  gate1229(.a(gate496inter11), .b(gate496inter6), .O(gate496inter12));
  nand2 gate1230(.a(gate496inter12), .b(gate496inter1), .O(N1742));
nand2 gate497( .a(N1600), .b(N1709), .O(N1746) );
nand2 gate498( .a(N1603), .b(N1711), .O(N1747) );

  xor2  gate979(.a(N1712), .b(N1678), .O(gate499inter0));
  nand2 gate980(.a(gate499inter0), .b(s_14), .O(gate499inter1));
  and2  gate981(.a(N1712), .b(N1678), .O(gate499inter2));
  inv1  gate982(.a(s_14), .O(gate499inter3));
  inv1  gate983(.a(s_15), .O(gate499inter4));
  nand2 gate984(.a(gate499inter4), .b(gate499inter3), .O(gate499inter5));
  nor2  gate985(.a(gate499inter5), .b(gate499inter2), .O(gate499inter6));
  inv1  gate986(.a(N1678), .O(gate499inter7));
  inv1  gate987(.a(N1712), .O(gate499inter8));
  nand2 gate988(.a(gate499inter8), .b(gate499inter7), .O(gate499inter9));
  nand2 gate989(.a(s_15), .b(gate499inter3), .O(gate499inter10));
  nor2  gate990(.a(gate499inter10), .b(gate499inter9), .O(gate499inter11));
  nor2  gate991(.a(gate499inter11), .b(gate499inter6), .O(gate499inter12));
  nand2 gate992(.a(gate499inter12), .b(gate499inter1), .O(N1748));
nand2 gate500( .a(N1680), .b(N1713), .O(N1751) );
nand2 gate501( .a(N1537), .b(N1721), .O(N1759) );
inv1 gate502( .a(N1697), .O(N1761) );

  xor2  gate1329(.a(N1727), .b(N1697), .O(gate503inter0));
  nand2 gate1330(.a(gate503inter0), .b(s_64), .O(gate503inter1));
  and2  gate1331(.a(N1727), .b(N1697), .O(gate503inter2));
  inv1  gate1332(.a(s_64), .O(gate503inter3));
  inv1  gate1333(.a(s_65), .O(gate503inter4));
  nand2 gate1334(.a(gate503inter4), .b(gate503inter3), .O(gate503inter5));
  nor2  gate1335(.a(gate503inter5), .b(gate503inter2), .O(gate503inter6));
  inv1  gate1336(.a(N1697), .O(gate503inter7));
  inv1  gate1337(.a(N1727), .O(gate503inter8));
  nand2 gate1338(.a(gate503inter8), .b(gate503inter7), .O(gate503inter9));
  nand2 gate1339(.a(s_65), .b(gate503inter3), .O(gate503inter10));
  nor2  gate1340(.a(gate503inter10), .b(gate503inter9), .O(gate503inter11));
  nor2  gate1341(.a(gate503inter11), .b(gate503inter6), .O(gate503inter12));
  nand2 gate1342(.a(gate503inter12), .b(gate503inter1), .O(N1762));
inv1 gate504( .a(N1701), .O(N1763) );
nand2 gate505( .a(N1701), .b(N1730), .O(N1764) );
inv1 gate506( .a(N1717), .O(N1768) );
nand2 gate507( .a(N1472), .b(N1741), .O(N1769) );
nand2 gate508( .a(N1723), .b(N1413), .O(N1772) );
inv1 gate509( .a(N1723), .O(N1773) );
nand2 gate510( .a(N1708), .b(N1746), .O(N1774) );
nand2 gate511( .a(N1710), .b(N1747), .O(N1777) );
inv1 gate512( .a(N1731), .O(N1783) );
nand2 gate513( .a(N1731), .b(N1682), .O(N1784) );
inv1 gate514( .a(N1714), .O(N1785) );
inv1 gate515( .a(N1734), .O(N1786) );
nand2 gate516( .a(N1734), .b(N1683), .O(N1787) );
nand2 gate517( .a(N1720), .b(N1759), .O(N1788) );
nand2 gate518( .a(N1661), .b(N1761), .O(N1791) );
nand2 gate519( .a(N1664), .b(N1763), .O(N1792) );
nand2 gate520( .a(N1751), .b(N1155), .O(N1795) );
inv1 gate521( .a(N1751), .O(N1796) );
nand2 gate522( .a(N1740), .b(N1769), .O(N1798) );

  xor2  gate1763(.a(N1773), .b(N1334), .O(gate523inter0));
  nand2 gate1764(.a(gate523inter0), .b(s_126), .O(gate523inter1));
  and2  gate1765(.a(N1773), .b(N1334), .O(gate523inter2));
  inv1  gate1766(.a(s_126), .O(gate523inter3));
  inv1  gate1767(.a(s_127), .O(gate523inter4));
  nand2 gate1768(.a(gate523inter4), .b(gate523inter3), .O(gate523inter5));
  nor2  gate1769(.a(gate523inter5), .b(gate523inter2), .O(gate523inter6));
  inv1  gate1770(.a(N1334), .O(gate523inter7));
  inv1  gate1771(.a(N1773), .O(gate523inter8));
  nand2 gate1772(.a(gate523inter8), .b(gate523inter7), .O(gate523inter9));
  nand2 gate1773(.a(s_127), .b(gate523inter3), .O(gate523inter10));
  nor2  gate1774(.a(gate523inter10), .b(gate523inter9), .O(gate523inter11));
  nor2  gate1775(.a(gate523inter11), .b(gate523inter6), .O(gate523inter12));
  nand2 gate1776(.a(gate523inter12), .b(gate523inter1), .O(N1801));
nand2 gate524( .a(N1742), .b(N290), .O(N1802) );
inv1 gate525( .a(N1748), .O(N1807) );

  xor2  gate1371(.a(N1218), .b(N1748), .O(gate526inter0));
  nand2 gate1372(.a(gate526inter0), .b(s_70), .O(gate526inter1));
  and2  gate1373(.a(N1218), .b(N1748), .O(gate526inter2));
  inv1  gate1374(.a(s_70), .O(gate526inter3));
  inv1  gate1375(.a(s_71), .O(gate526inter4));
  nand2 gate1376(.a(gate526inter4), .b(gate526inter3), .O(gate526inter5));
  nor2  gate1377(.a(gate526inter5), .b(gate526inter2), .O(gate526inter6));
  inv1  gate1378(.a(N1748), .O(gate526inter7));
  inv1  gate1379(.a(N1218), .O(gate526inter8));
  nand2 gate1380(.a(gate526inter8), .b(gate526inter7), .O(gate526inter9));
  nand2 gate1381(.a(s_71), .b(gate526inter3), .O(gate526inter10));
  nor2  gate1382(.a(gate526inter10), .b(gate526inter9), .O(gate526inter11));
  nor2  gate1383(.a(gate526inter11), .b(gate526inter6), .O(gate526inter12));
  nand2 gate1384(.a(gate526inter12), .b(gate526inter1), .O(N1808));

  xor2  gate965(.a(N1783), .b(N1612), .O(gate527inter0));
  nand2 gate966(.a(gate527inter0), .b(s_12), .O(gate527inter1));
  and2  gate967(.a(N1783), .b(N1612), .O(gate527inter2));
  inv1  gate968(.a(s_12), .O(gate527inter3));
  inv1  gate969(.a(s_13), .O(gate527inter4));
  nand2 gate970(.a(gate527inter4), .b(gate527inter3), .O(gate527inter5));
  nor2  gate971(.a(gate527inter5), .b(gate527inter2), .O(gate527inter6));
  inv1  gate972(.a(N1612), .O(gate527inter7));
  inv1  gate973(.a(N1783), .O(gate527inter8));
  nand2 gate974(.a(gate527inter8), .b(gate527inter7), .O(gate527inter9));
  nand2 gate975(.a(s_13), .b(gate527inter3), .O(gate527inter10));
  nor2  gate976(.a(gate527inter10), .b(gate527inter9), .O(gate527inter11));
  nor2  gate977(.a(gate527inter11), .b(gate527inter6), .O(gate527inter12));
  nand2 gate978(.a(gate527inter12), .b(gate527inter1), .O(N1809));

  xor2  gate1511(.a(N1786), .b(N1615), .O(gate528inter0));
  nand2 gate1512(.a(gate528inter0), .b(s_90), .O(gate528inter1));
  and2  gate1513(.a(N1786), .b(N1615), .O(gate528inter2));
  inv1  gate1514(.a(s_90), .O(gate528inter3));
  inv1  gate1515(.a(s_91), .O(gate528inter4));
  nand2 gate1516(.a(gate528inter4), .b(gate528inter3), .O(gate528inter5));
  nor2  gate1517(.a(gate528inter5), .b(gate528inter2), .O(gate528inter6));
  inv1  gate1518(.a(N1615), .O(gate528inter7));
  inv1  gate1519(.a(N1786), .O(gate528inter8));
  nand2 gate1520(.a(gate528inter8), .b(gate528inter7), .O(gate528inter9));
  nand2 gate1521(.a(s_91), .b(gate528inter3), .O(gate528inter10));
  nor2  gate1522(.a(gate528inter10), .b(gate528inter9), .O(gate528inter11));
  nor2  gate1523(.a(gate528inter11), .b(gate528inter6), .O(gate528inter12));
  nand2 gate1524(.a(gate528inter12), .b(gate528inter1), .O(N1810));

  xor2  gate1189(.a(N1762), .b(N1791), .O(gate529inter0));
  nand2 gate1190(.a(gate529inter0), .b(s_44), .O(gate529inter1));
  and2  gate1191(.a(N1762), .b(N1791), .O(gate529inter2));
  inv1  gate1192(.a(s_44), .O(gate529inter3));
  inv1  gate1193(.a(s_45), .O(gate529inter4));
  nand2 gate1194(.a(gate529inter4), .b(gate529inter3), .O(gate529inter5));
  nor2  gate1195(.a(gate529inter5), .b(gate529inter2), .O(gate529inter6));
  inv1  gate1196(.a(N1791), .O(gate529inter7));
  inv1  gate1197(.a(N1762), .O(gate529inter8));
  nand2 gate1198(.a(gate529inter8), .b(gate529inter7), .O(gate529inter9));
  nand2 gate1199(.a(s_45), .b(gate529inter3), .O(gate529inter10));
  nor2  gate1200(.a(gate529inter10), .b(gate529inter9), .O(gate529inter11));
  nor2  gate1201(.a(gate529inter11), .b(gate529inter6), .O(gate529inter12));
  nand2 gate1202(.a(gate529inter12), .b(gate529inter1), .O(N1812));
nand2 gate530( .a(N1792), .b(N1764), .O(N1815) );
buf1 gate531( .a(N1742), .O(N1818) );
nand2 gate532( .a(N1777), .b(N1490), .O(N1821) );
inv1 gate533( .a(N1777), .O(N1822) );
nand2 gate534( .a(N1774), .b(N1491), .O(N1823) );
inv1 gate535( .a(N1774), .O(N1824) );
nand2 gate536( .a(N962), .b(N1796), .O(N1825) );
nand2 gate537( .a(N1788), .b(N1409), .O(N1826) );
inv1 gate538( .a(N1788), .O(N1827) );

  xor2  gate1595(.a(N1801), .b(N1772), .O(gate539inter0));
  nand2 gate1596(.a(gate539inter0), .b(s_102), .O(gate539inter1));
  and2  gate1597(.a(N1801), .b(N1772), .O(gate539inter2));
  inv1  gate1598(.a(s_102), .O(gate539inter3));
  inv1  gate1599(.a(s_103), .O(gate539inter4));
  nand2 gate1600(.a(gate539inter4), .b(gate539inter3), .O(gate539inter5));
  nor2  gate1601(.a(gate539inter5), .b(gate539inter2), .O(gate539inter6));
  inv1  gate1602(.a(N1772), .O(gate539inter7));
  inv1  gate1603(.a(N1801), .O(gate539inter8));
  nand2 gate1604(.a(gate539inter8), .b(gate539inter7), .O(gate539inter9));
  nand2 gate1605(.a(s_103), .b(gate539inter3), .O(gate539inter10));
  nor2  gate1606(.a(gate539inter10), .b(gate539inter9), .O(gate539inter11));
  nor2  gate1607(.a(gate539inter11), .b(gate539inter6), .O(gate539inter12));
  nand2 gate1608(.a(gate539inter12), .b(gate539inter1), .O(N1830));
nand2 gate540( .a(N959), .b(N1807), .O(N1837) );
nand2 gate541( .a(N1809), .b(N1784), .O(N1838) );
nand2 gate542( .a(N1810), .b(N1787), .O(N1841) );
nand2 gate543( .a(N1419), .b(N1822), .O(N1848) );
nand2 gate544( .a(N1416), .b(N1824), .O(N1849) );
nand2 gate545( .a(N1795), .b(N1825), .O(N1850) );
nand2 gate546( .a(N1319), .b(N1827), .O(N1852) );

  xor2  gate1679(.a(N1707), .b(N1815), .O(gate547inter0));
  nand2 gate1680(.a(gate547inter0), .b(s_114), .O(gate547inter1));
  and2  gate1681(.a(N1707), .b(N1815), .O(gate547inter2));
  inv1  gate1682(.a(s_114), .O(gate547inter3));
  inv1  gate1683(.a(s_115), .O(gate547inter4));
  nand2 gate1684(.a(gate547inter4), .b(gate547inter3), .O(gate547inter5));
  nor2  gate1685(.a(gate547inter5), .b(gate547inter2), .O(gate547inter6));
  inv1  gate1686(.a(N1815), .O(gate547inter7));
  inv1  gate1687(.a(N1707), .O(gate547inter8));
  nand2 gate1688(.a(gate547inter8), .b(gate547inter7), .O(gate547inter9));
  nand2 gate1689(.a(s_115), .b(gate547inter3), .O(gate547inter10));
  nor2  gate1690(.a(gate547inter10), .b(gate547inter9), .O(gate547inter11));
  nor2  gate1691(.a(gate547inter11), .b(gate547inter6), .O(gate547inter12));
  nand2 gate1692(.a(gate547inter12), .b(gate547inter1), .O(N1855));
inv1 gate548( .a(N1815), .O(N1856) );
inv1 gate549( .a(N1818), .O(N1857) );
nand2 gate550( .a(N1798), .b(N290), .O(N1858) );
inv1 gate551( .a(N1812), .O(N1864) );
nand2 gate552( .a(N1812), .b(N1728), .O(N1865) );
buf1 gate553( .a(N1798), .O(N1866) );
buf1 gate554( .a(N1802), .O(N1869) );
buf1 gate555( .a(N1802), .O(N1872) );
nand2 gate556( .a(N1808), .b(N1837), .O(N1875) );
nand2 gate557( .a(N1821), .b(N1848), .O(N1878) );
nand2 gate558( .a(N1823), .b(N1849), .O(N1879) );
nand2 gate559( .a(N1841), .b(N1768), .O(N1882) );
inv1 gate560( .a(N1841), .O(N1883) );
nand2 gate561( .a(N1826), .b(N1852), .O(N1884) );
nand2 gate562( .a(N1643), .b(N1856), .O(N1885) );

  xor2  gate1119(.a(N290), .b(N1830), .O(gate563inter0));
  nand2 gate1120(.a(gate563inter0), .b(s_34), .O(gate563inter1));
  and2  gate1121(.a(N290), .b(N1830), .O(gate563inter2));
  inv1  gate1122(.a(s_34), .O(gate563inter3));
  inv1  gate1123(.a(s_35), .O(gate563inter4));
  nand2 gate1124(.a(gate563inter4), .b(gate563inter3), .O(gate563inter5));
  nor2  gate1125(.a(gate563inter5), .b(gate563inter2), .O(gate563inter6));
  inv1  gate1126(.a(N1830), .O(gate563inter7));
  inv1  gate1127(.a(N290), .O(gate563inter8));
  nand2 gate1128(.a(gate563inter8), .b(gate563inter7), .O(gate563inter9));
  nand2 gate1129(.a(s_35), .b(gate563inter3), .O(gate563inter10));
  nor2  gate1130(.a(gate563inter10), .b(gate563inter9), .O(gate563inter11));
  nor2  gate1131(.a(gate563inter11), .b(gate563inter6), .O(gate563inter12));
  nand2 gate1132(.a(gate563inter12), .b(gate563inter1), .O(N1889));
inv1 gate564( .a(N1838), .O(N1895) );
nand2 gate565( .a(N1838), .b(N1785), .O(N1896) );
nand2 gate566( .a(N1640), .b(N1864), .O(N1897) );
inv1 gate567( .a(N1850), .O(N1898) );
buf1 gate568( .a(N1830), .O(N1902) );
inv1 gate569( .a(N1878), .O(N1910) );
nand2 gate570( .a(N1717), .b(N1883), .O(N1911) );
inv1 gate571( .a(N1884), .O(N1912) );
nand2 gate572( .a(N1855), .b(N1885), .O(N1913) );
inv1 gate573( .a(N1866), .O(N1915) );

  xor2  gate1175(.a(N919), .b(N1872), .O(gate574inter0));
  nand2 gate1176(.a(gate574inter0), .b(s_42), .O(gate574inter1));
  and2  gate1177(.a(N919), .b(N1872), .O(gate574inter2));
  inv1  gate1178(.a(s_42), .O(gate574inter3));
  inv1  gate1179(.a(s_43), .O(gate574inter4));
  nand2 gate1180(.a(gate574inter4), .b(gate574inter3), .O(gate574inter5));
  nor2  gate1181(.a(gate574inter5), .b(gate574inter2), .O(gate574inter6));
  inv1  gate1182(.a(N1872), .O(gate574inter7));
  inv1  gate1183(.a(N919), .O(gate574inter8));
  nand2 gate1184(.a(gate574inter8), .b(gate574inter7), .O(gate574inter9));
  nand2 gate1185(.a(s_43), .b(gate574inter3), .O(gate574inter10));
  nor2  gate1186(.a(gate574inter10), .b(gate574inter9), .O(gate574inter11));
  nor2  gate1187(.a(gate574inter11), .b(gate574inter6), .O(gate574inter12));
  nand2 gate1188(.a(gate574inter12), .b(gate574inter1), .O(N1919));
inv1 gate575( .a(N1872), .O(N1920) );
nand2 gate576( .a(N1869), .b(N920), .O(N1921) );
inv1 gate577( .a(N1869), .O(N1922) );
inv1 gate578( .a(N1875), .O(N1923) );
nand2 gate579( .a(N1714), .b(N1895), .O(N1924) );
buf1 gate580( .a(N1858), .O(N1927) );
buf1 gate581( .a(N1858), .O(N1930) );
nand2 gate582( .a(N1865), .b(N1897), .O(N1933) );
nand2 gate583( .a(N1882), .b(N1911), .O(N1936) );
inv1 gate584( .a(N1898), .O(N1937) );
inv1 gate585( .a(N1902), .O(N1938) );

  xor2  gate923(.a(N1920), .b(N679), .O(gate586inter0));
  nand2 gate924(.a(gate586inter0), .b(s_6), .O(gate586inter1));
  and2  gate925(.a(N1920), .b(N679), .O(gate586inter2));
  inv1  gate926(.a(s_6), .O(gate586inter3));
  inv1  gate927(.a(s_7), .O(gate586inter4));
  nand2 gate928(.a(gate586inter4), .b(gate586inter3), .O(gate586inter5));
  nor2  gate929(.a(gate586inter5), .b(gate586inter2), .O(gate586inter6));
  inv1  gate930(.a(N679), .O(gate586inter7));
  inv1  gate931(.a(N1920), .O(gate586inter8));
  nand2 gate932(.a(gate586inter8), .b(gate586inter7), .O(gate586inter9));
  nand2 gate933(.a(s_7), .b(gate586inter3), .O(gate586inter10));
  nor2  gate934(.a(gate586inter10), .b(gate586inter9), .O(gate586inter11));
  nor2  gate935(.a(gate586inter11), .b(gate586inter6), .O(gate586inter12));
  nand2 gate936(.a(gate586inter12), .b(gate586inter1), .O(N1941));
nand2 gate587( .a(N676), .b(N1922), .O(N1942) );
buf1 gate588( .a(N1879), .O(N1944) );
inv1 gate589( .a(N1913), .O(N1947) );
buf1 gate590( .a(N1889), .O(N1950) );
buf1 gate591( .a(N1889), .O(N1953) );
buf1 gate592( .a(N1879), .O(N1958) );
nand2 gate593( .a(N1896), .b(N1924), .O(N1961) );
and2 gate594( .a(N1910), .b(N601), .O(N1965) );
and2 gate595( .a(N602), .b(N1912), .O(N1968) );
nand2 gate596( .a(N1930), .b(N917), .O(N1975) );
inv1 gate597( .a(N1930), .O(N1976) );
nand2 gate598( .a(N1927), .b(N918), .O(N1977) );
inv1 gate599( .a(N1927), .O(N1978) );

  xor2  gate1161(.a(N1941), .b(N1919), .O(gate600inter0));
  nand2 gate1162(.a(gate600inter0), .b(s_40), .O(gate600inter1));
  and2  gate1163(.a(N1941), .b(N1919), .O(gate600inter2));
  inv1  gate1164(.a(s_40), .O(gate600inter3));
  inv1  gate1165(.a(s_41), .O(gate600inter4));
  nand2 gate1166(.a(gate600inter4), .b(gate600inter3), .O(gate600inter5));
  nor2  gate1167(.a(gate600inter5), .b(gate600inter2), .O(gate600inter6));
  inv1  gate1168(.a(N1919), .O(gate600inter7));
  inv1  gate1169(.a(N1941), .O(gate600inter8));
  nand2 gate1170(.a(gate600inter8), .b(gate600inter7), .O(gate600inter9));
  nand2 gate1171(.a(s_41), .b(gate600inter3), .O(gate600inter10));
  nor2  gate1172(.a(gate600inter10), .b(gate600inter9), .O(gate600inter11));
  nor2  gate1173(.a(gate600inter11), .b(gate600inter6), .O(gate600inter12));
  nand2 gate1174(.a(gate600inter12), .b(gate600inter1), .O(N1979));
nand2 gate601( .a(N1921), .b(N1942), .O(N1980) );
inv1 gate602( .a(N1933), .O(N1985) );
inv1 gate603( .a(N1936), .O(N1987) );
inv1 gate604( .a(N1944), .O(N1999) );
nand2 gate605( .a(N1944), .b(N1937), .O(N2000) );
inv1 gate606( .a(N1947), .O(N2002) );

  xor2  gate1651(.a(N1499), .b(N1947), .O(gate607inter0));
  nand2 gate1652(.a(gate607inter0), .b(s_110), .O(gate607inter1));
  and2  gate1653(.a(N1499), .b(N1947), .O(gate607inter2));
  inv1  gate1654(.a(s_110), .O(gate607inter3));
  inv1  gate1655(.a(s_111), .O(gate607inter4));
  nand2 gate1656(.a(gate607inter4), .b(gate607inter3), .O(gate607inter5));
  nor2  gate1657(.a(gate607inter5), .b(gate607inter2), .O(gate607inter6));
  inv1  gate1658(.a(N1947), .O(gate607inter7));
  inv1  gate1659(.a(N1499), .O(gate607inter8));
  nand2 gate1660(.a(gate607inter8), .b(gate607inter7), .O(gate607inter9));
  nand2 gate1661(.a(s_111), .b(gate607inter3), .O(gate607inter10));
  nor2  gate1662(.a(gate607inter10), .b(gate607inter9), .O(gate607inter11));
  nor2  gate1663(.a(gate607inter11), .b(gate607inter6), .O(gate607inter12));
  nand2 gate1664(.a(gate607inter12), .b(gate607inter1), .O(N2003));
nand2 gate608( .a(N1953), .b(N1350), .O(N2004) );
inv1 gate609( .a(N1953), .O(N2005) );
nand2 gate610( .a(N1950), .b(N1351), .O(N2006) );
inv1 gate611( .a(N1950), .O(N2007) );

  xor2  gate1497(.a(N1976), .b(N673), .O(gate612inter0));
  nand2 gate1498(.a(gate612inter0), .b(s_88), .O(gate612inter1));
  and2  gate1499(.a(N1976), .b(N673), .O(gate612inter2));
  inv1  gate1500(.a(s_88), .O(gate612inter3));
  inv1  gate1501(.a(s_89), .O(gate612inter4));
  nand2 gate1502(.a(gate612inter4), .b(gate612inter3), .O(gate612inter5));
  nor2  gate1503(.a(gate612inter5), .b(gate612inter2), .O(gate612inter6));
  inv1  gate1504(.a(N673), .O(gate612inter7));
  inv1  gate1505(.a(N1976), .O(gate612inter8));
  nand2 gate1506(.a(gate612inter8), .b(gate612inter7), .O(gate612inter9));
  nand2 gate1507(.a(s_89), .b(gate612inter3), .O(gate612inter10));
  nor2  gate1508(.a(gate612inter10), .b(gate612inter9), .O(gate612inter11));
  nor2  gate1509(.a(gate612inter11), .b(gate612inter6), .O(gate612inter12));
  nand2 gate1510(.a(gate612inter12), .b(gate612inter1), .O(N2008));
nand2 gate613( .a(N670), .b(N1978), .O(N2009) );
inv1 gate614( .a(N1979), .O(N2012) );
inv1 gate615( .a(N1958), .O(N2013) );

  xor2  gate1609(.a(N1923), .b(N1958), .O(gate616inter0));
  nand2 gate1610(.a(gate616inter0), .b(s_104), .O(gate616inter1));
  and2  gate1611(.a(N1923), .b(N1958), .O(gate616inter2));
  inv1  gate1612(.a(s_104), .O(gate616inter3));
  inv1  gate1613(.a(s_105), .O(gate616inter4));
  nand2 gate1614(.a(gate616inter4), .b(gate616inter3), .O(gate616inter5));
  nor2  gate1615(.a(gate616inter5), .b(gate616inter2), .O(gate616inter6));
  inv1  gate1616(.a(N1958), .O(gate616inter7));
  inv1  gate1617(.a(N1923), .O(gate616inter8));
  nand2 gate1618(.a(gate616inter8), .b(gate616inter7), .O(gate616inter9));
  nand2 gate1619(.a(s_105), .b(gate616inter3), .O(gate616inter10));
  nor2  gate1620(.a(gate616inter10), .b(gate616inter9), .O(gate616inter11));
  nor2  gate1621(.a(gate616inter11), .b(gate616inter6), .O(gate616inter12));
  nand2 gate1622(.a(gate616inter12), .b(gate616inter1), .O(N2014));
inv1 gate617( .a(N1961), .O(N2015) );
nand2 gate618( .a(N1961), .b(N1635), .O(N2016) );
inv1 gate619( .a(N1965), .O(N2018) );
inv1 gate620( .a(N1968), .O(N2019) );
nand2 gate621( .a(N1898), .b(N1999), .O(N2020) );
inv1 gate622( .a(N1987), .O(N2021) );

  xor2  gate1413(.a(N1591), .b(N1987), .O(gate623inter0));
  nand2 gate1414(.a(gate623inter0), .b(s_76), .O(gate623inter1));
  and2  gate1415(.a(N1591), .b(N1987), .O(gate623inter2));
  inv1  gate1416(.a(s_76), .O(gate623inter3));
  inv1  gate1417(.a(s_77), .O(gate623inter4));
  nand2 gate1418(.a(gate623inter4), .b(gate623inter3), .O(gate623inter5));
  nor2  gate1419(.a(gate623inter5), .b(gate623inter2), .O(gate623inter6));
  inv1  gate1420(.a(N1987), .O(gate623inter7));
  inv1  gate1421(.a(N1591), .O(gate623inter8));
  nand2 gate1422(.a(gate623inter8), .b(gate623inter7), .O(gate623inter9));
  nand2 gate1423(.a(s_77), .b(gate623inter3), .O(gate623inter10));
  nor2  gate1424(.a(gate623inter10), .b(gate623inter9), .O(gate623inter11));
  nor2  gate1425(.a(gate623inter11), .b(gate623inter6), .O(gate623inter12));
  nand2 gate1426(.a(gate623inter12), .b(gate623inter1), .O(N2022));

  xor2  gate1427(.a(N2002), .b(N1440), .O(gate624inter0));
  nand2 gate1428(.a(gate624inter0), .b(s_78), .O(gate624inter1));
  and2  gate1429(.a(N2002), .b(N1440), .O(gate624inter2));
  inv1  gate1430(.a(s_78), .O(gate624inter3));
  inv1  gate1431(.a(s_79), .O(gate624inter4));
  nand2 gate1432(.a(gate624inter4), .b(gate624inter3), .O(gate624inter5));
  nor2  gate1433(.a(gate624inter5), .b(gate624inter2), .O(gate624inter6));
  inv1  gate1434(.a(N1440), .O(gate624inter7));
  inv1  gate1435(.a(N2002), .O(gate624inter8));
  nand2 gate1436(.a(gate624inter8), .b(gate624inter7), .O(gate624inter9));
  nand2 gate1437(.a(s_79), .b(gate624inter3), .O(gate624inter10));
  nor2  gate1438(.a(gate624inter10), .b(gate624inter9), .O(gate624inter11));
  nor2  gate1439(.a(gate624inter11), .b(gate624inter6), .O(gate624inter12));
  nand2 gate1440(.a(gate624inter12), .b(gate624inter1), .O(N2023));

  xor2  gate1399(.a(N2005), .b(N1261), .O(gate625inter0));
  nand2 gate1400(.a(gate625inter0), .b(s_74), .O(gate625inter1));
  and2  gate1401(.a(N2005), .b(N1261), .O(gate625inter2));
  inv1  gate1402(.a(s_74), .O(gate625inter3));
  inv1  gate1403(.a(s_75), .O(gate625inter4));
  nand2 gate1404(.a(gate625inter4), .b(gate625inter3), .O(gate625inter5));
  nor2  gate1405(.a(gate625inter5), .b(gate625inter2), .O(gate625inter6));
  inv1  gate1406(.a(N1261), .O(gate625inter7));
  inv1  gate1407(.a(N2005), .O(gate625inter8));
  nand2 gate1408(.a(gate625inter8), .b(gate625inter7), .O(gate625inter9));
  nand2 gate1409(.a(s_75), .b(gate625inter3), .O(gate625inter10));
  nor2  gate1410(.a(gate625inter10), .b(gate625inter9), .O(gate625inter11));
  nor2  gate1411(.a(gate625inter11), .b(gate625inter6), .O(gate625inter12));
  nand2 gate1412(.a(gate625inter12), .b(gate625inter1), .O(N2024));
nand2 gate626( .a(N1258), .b(N2007), .O(N2025) );
nand2 gate627( .a(N1975), .b(N2008), .O(N2026) );

  xor2  gate1567(.a(N2009), .b(N1977), .O(gate628inter0));
  nand2 gate1568(.a(gate628inter0), .b(s_98), .O(gate628inter1));
  and2  gate1569(.a(N2009), .b(N1977), .O(gate628inter2));
  inv1  gate1570(.a(s_98), .O(gate628inter3));
  inv1  gate1571(.a(s_99), .O(gate628inter4));
  nand2 gate1572(.a(gate628inter4), .b(gate628inter3), .O(gate628inter5));
  nor2  gate1573(.a(gate628inter5), .b(gate628inter2), .O(gate628inter6));
  inv1  gate1574(.a(N1977), .O(gate628inter7));
  inv1  gate1575(.a(N2009), .O(gate628inter8));
  nand2 gate1576(.a(gate628inter8), .b(gate628inter7), .O(gate628inter9));
  nand2 gate1577(.a(s_99), .b(gate628inter3), .O(gate628inter10));
  nor2  gate1578(.a(gate628inter10), .b(gate628inter9), .O(gate628inter11));
  nor2  gate1579(.a(gate628inter11), .b(gate628inter6), .O(gate628inter12));
  nand2 gate1580(.a(gate628inter12), .b(gate628inter1), .O(N2027));
inv1 gate629( .a(N1980), .O(N2030) );
buf1 gate630( .a(N1980), .O(N2033) );
nand2 gate631( .a(N1875), .b(N2013), .O(N2036) );
nand2 gate632( .a(N1571), .b(N2015), .O(N2037) );

  xor2  gate1343(.a(N2000), .b(N2020), .O(gate633inter0));
  nand2 gate1344(.a(gate633inter0), .b(s_66), .O(gate633inter1));
  and2  gate1345(.a(N2000), .b(N2020), .O(gate633inter2));
  inv1  gate1346(.a(s_66), .O(gate633inter3));
  inv1  gate1347(.a(s_67), .O(gate633inter4));
  nand2 gate1348(.a(gate633inter4), .b(gate633inter3), .O(gate633inter5));
  nor2  gate1349(.a(gate633inter5), .b(gate633inter2), .O(gate633inter6));
  inv1  gate1350(.a(N2020), .O(gate633inter7));
  inv1  gate1351(.a(N2000), .O(gate633inter8));
  nand2 gate1352(.a(gate633inter8), .b(gate633inter7), .O(gate633inter9));
  nand2 gate1353(.a(s_67), .b(gate633inter3), .O(gate633inter10));
  nor2  gate1354(.a(gate633inter10), .b(gate633inter9), .O(gate633inter11));
  nor2  gate1355(.a(gate633inter11), .b(gate633inter6), .O(gate633inter12));
  nand2 gate1356(.a(gate633inter12), .b(gate633inter1), .O(N2038));
nand2 gate634( .a(N1534), .b(N2021), .O(N2039) );

  xor2  gate1539(.a(N2003), .b(N2023), .O(gate635inter0));
  nand2 gate1540(.a(gate635inter0), .b(s_94), .O(gate635inter1));
  and2  gate1541(.a(N2003), .b(N2023), .O(gate635inter2));
  inv1  gate1542(.a(s_94), .O(gate635inter3));
  inv1  gate1543(.a(s_95), .O(gate635inter4));
  nand2 gate1544(.a(gate635inter4), .b(gate635inter3), .O(gate635inter5));
  nor2  gate1545(.a(gate635inter5), .b(gate635inter2), .O(gate635inter6));
  inv1  gate1546(.a(N2023), .O(gate635inter7));
  inv1  gate1547(.a(N2003), .O(gate635inter8));
  nand2 gate1548(.a(gate635inter8), .b(gate635inter7), .O(gate635inter9));
  nand2 gate1549(.a(s_95), .b(gate635inter3), .O(gate635inter10));
  nor2  gate1550(.a(gate635inter10), .b(gate635inter9), .O(gate635inter11));
  nor2  gate1551(.a(gate635inter11), .b(gate635inter6), .O(gate635inter12));
  nand2 gate1552(.a(gate635inter12), .b(gate635inter1), .O(N2040));
nand2 gate636( .a(N2004), .b(N2024), .O(N2041) );
nand2 gate637( .a(N2006), .b(N2025), .O(N2042) );
inv1 gate638( .a(N2026), .O(N2047) );
nand2 gate639( .a(N2036), .b(N2014), .O(N2052) );
nand2 gate640( .a(N2037), .b(N2016), .O(N2055) );
inv1 gate641( .a(N2038), .O(N2060) );
nand2 gate642( .a(N2039), .b(N2022), .O(N2061) );
nand2 gate643( .a(N2040), .b(N290), .O(N2062) );
inv1 gate644( .a(N2041), .O(N2067) );
inv1 gate645( .a(N2027), .O(N2068) );
buf1 gate646( .a(N2027), .O(N2071) );
inv1 gate647( .a(N2052), .O(N2076) );
inv1 gate648( .a(N2055), .O(N2077) );
nand2 gate649( .a(N2060), .b(N290), .O(N2078) );
nand2 gate650( .a(N2061), .b(N290), .O(N2081) );
inv1 gate651( .a(N2042), .O(N2086) );
buf1 gate652( .a(N2042), .O(N2089) );
and2 gate653( .a(N2030), .b(N2068), .O(N2104) );
and2 gate654( .a(N2033), .b(N2068), .O(N2119) );
and2 gate655( .a(N2030), .b(N2071), .O(N2129) );
and2 gate656( .a(N2033), .b(N2071), .O(N2143) );
buf1 gate657( .a(N2062), .O(N2148) );
buf1 gate658( .a(N2062), .O(N2151) );
buf1 gate659( .a(N2078), .O(N2196) );
buf1 gate660( .a(N2078), .O(N2199) );
buf1 gate661( .a(N2081), .O(N2202) );
buf1 gate662( .a(N2081), .O(N2205) );
nand2 gate663( .a(N2151), .b(N915), .O(N2214) );
inv1 gate664( .a(N2151), .O(N2215) );
nand2 gate665( .a(N2148), .b(N916), .O(N2216) );
inv1 gate666( .a(N2148), .O(N2217) );
nand2 gate667( .a(N2199), .b(N1348), .O(N2222) );
inv1 gate668( .a(N2199), .O(N2223) );
nand2 gate669( .a(N2196), .b(N1349), .O(N2224) );
inv1 gate670( .a(N2196), .O(N2225) );
nand2 gate671( .a(N2205), .b(N913), .O(N2226) );
inv1 gate672( .a(N2205), .O(N2227) );
nand2 gate673( .a(N2202), .b(N914), .O(N2228) );
inv1 gate674( .a(N2202), .O(N2229) );
nand2 gate675( .a(N667), .b(N2215), .O(N2230) );
nand2 gate676( .a(N664), .b(N2217), .O(N2231) );
nand2 gate677( .a(N1255), .b(N2223), .O(N2232) );
nand2 gate678( .a(N1252), .b(N2225), .O(N2233) );
nand2 gate679( .a(N661), .b(N2227), .O(N2234) );
nand2 gate680( .a(N658), .b(N2229), .O(N2235) );
nand2 gate681( .a(N2214), .b(N2230), .O(N2236) );
nand2 gate682( .a(N2216), .b(N2231), .O(N2237) );

  xor2  gate1007(.a(N2232), .b(N2222), .O(gate683inter0));
  nand2 gate1008(.a(gate683inter0), .b(s_18), .O(gate683inter1));
  and2  gate1009(.a(N2232), .b(N2222), .O(gate683inter2));
  inv1  gate1010(.a(s_18), .O(gate683inter3));
  inv1  gate1011(.a(s_19), .O(gate683inter4));
  nand2 gate1012(.a(gate683inter4), .b(gate683inter3), .O(gate683inter5));
  nor2  gate1013(.a(gate683inter5), .b(gate683inter2), .O(gate683inter6));
  inv1  gate1014(.a(N2222), .O(gate683inter7));
  inv1  gate1015(.a(N2232), .O(gate683inter8));
  nand2 gate1016(.a(gate683inter8), .b(gate683inter7), .O(gate683inter9));
  nand2 gate1017(.a(s_19), .b(gate683inter3), .O(gate683inter10));
  nor2  gate1018(.a(gate683inter10), .b(gate683inter9), .O(gate683inter11));
  nor2  gate1019(.a(gate683inter11), .b(gate683inter6), .O(gate683inter12));
  nand2 gate1020(.a(gate683inter12), .b(gate683inter1), .O(N2240));
nand2 gate684( .a(N2224), .b(N2233), .O(N2241) );
nand2 gate685( .a(N2226), .b(N2234), .O(N2244) );
nand2 gate686( .a(N2228), .b(N2235), .O(N2245) );
inv1 gate687( .a(N2236), .O(N2250) );
inv1 gate688( .a(N2240), .O(N2253) );
inv1 gate689( .a(N2244), .O(N2256) );
inv1 gate690( .a(N2237), .O(N2257) );
buf1 gate691( .a(N2237), .O(N2260) );
inv1 gate692( .a(N2241), .O(N2263) );
and2 gate693( .a(N1164), .b(N2241), .O(N2266) );
inv1 gate694( .a(N2245), .O(N2269) );
and2 gate695( .a(N1168), .b(N2245), .O(N2272) );
nand8 gate696( .a(N2067), .b(N2012), .c(N2047), .d(N2250), .e(N899), .f(N2256), .g(N2253), .h(N903), .O(N2279) );
buf1 gate697( .a(N2266), .O(N2286) );
buf1 gate698( .a(N2266), .O(N2297) );
buf1 gate699( .a(N2272), .O(N2315) );
buf1 gate700( .a(N2272), .O(N2326) );
and2 gate701( .a(N2086), .b(N2257), .O(N2340) );
and2 gate702( .a(N2089), .b(N2257), .O(N2353) );
and2 gate703( .a(N2086), .b(N2260), .O(N2361) );
and2 gate704( .a(N2089), .b(N2260), .O(N2375) );
and4 gate705( .a(N338), .b(N2279), .c(N313), .d(N313), .O(N2384) );
and2 gate706( .a(N1163), .b(N2263), .O(N2385) );
and2 gate707( .a(N1164), .b(N2263), .O(N2386) );
and2 gate708( .a(N1167), .b(N2269), .O(N2426) );
and2 gate709( .a(N1168), .b(N2269), .O(N2427) );
nand5 gate710( .a(N2286), .b(N2315), .c(N2361), .d(N2104), .e(N1171), .O(N2537) );
nand5 gate711( .a(N2286), .b(N2315), .c(N2340), .d(N2129), .e(N1171), .O(N2540) );
nand5 gate712( .a(N2286), .b(N2315), .c(N2340), .d(N2119), .e(N1171), .O(N2543) );
nand5 gate713( .a(N2286), .b(N2315), .c(N2353), .d(N2104), .e(N1171), .O(N2546) );
nand5 gate714( .a(N2297), .b(N2315), .c(N2375), .d(N2119), .e(N1188), .O(N2549) );
nand5 gate715( .a(N2297), .b(N2326), .c(N2361), .d(N2143), .e(N1188), .O(N2552) );
nand5 gate716( .a(N2297), .b(N2326), .c(N2375), .d(N2129), .e(N1188), .O(N2555) );
and5 gate717( .a(N2286), .b(N2315), .c(N2361), .d(N2104), .e(N1171), .O(N2558) );
and5 gate718( .a(N2286), .b(N2315), .c(N2340), .d(N2129), .e(N1171), .O(N2561) );
and5 gate719( .a(N2286), .b(N2315), .c(N2340), .d(N2119), .e(N1171), .O(N2564) );
and5 gate720( .a(N2286), .b(N2315), .c(N2353), .d(N2104), .e(N1171), .O(N2567) );
and5 gate721( .a(N2297), .b(N2315), .c(N2375), .d(N2119), .e(N1188), .O(N2570) );
and5 gate722( .a(N2297), .b(N2326), .c(N2361), .d(N2143), .e(N1188), .O(N2573) );
and5 gate723( .a(N2297), .b(N2326), .c(N2375), .d(N2129), .e(N1188), .O(N2576) );
nand5 gate724( .a(N2286), .b(N2427), .c(N2361), .d(N2129), .e(N1171), .O(N2594) );
nand5 gate725( .a(N2297), .b(N2427), .c(N2361), .d(N2119), .e(N1171), .O(N2597) );
nand5 gate726( .a(N2297), .b(N2427), .c(N2375), .d(N2104), .e(N1171), .O(N2600) );
nand5 gate727( .a(N2297), .b(N2427), .c(N2340), .d(N2143), .e(N1171), .O(N2603) );
nand5 gate728( .a(N2297), .b(N2427), .c(N2353), .d(N2129), .e(N1188), .O(N2606) );
nand5 gate729( .a(N2386), .b(N2326), .c(N2361), .d(N2129), .e(N1188), .O(N2611) );
nand5 gate730( .a(N2386), .b(N2326), .c(N2361), .d(N2119), .e(N1188), .O(N2614) );
nand5 gate731( .a(N2386), .b(N2326), .c(N2375), .d(N2104), .e(N1188), .O(N2617) );
nand5 gate732( .a(N2386), .b(N2326), .c(N2353), .d(N2129), .e(N1188), .O(N2620) );
nand5 gate733( .a(N2297), .b(N2427), .c(N2340), .d(N2104), .e(N926), .O(N2627) );
nand5 gate734( .a(N2386), .b(N2326), .c(N2340), .d(N2104), .e(N926), .O(N2628) );
nand5 gate735( .a(N2386), .b(N2427), .c(N2361), .d(N2104), .e(N926), .O(N2629) );
nand5 gate736( .a(N2386), .b(N2427), .c(N2340), .d(N2129), .e(N926), .O(N2630) );
nand5 gate737( .a(N2386), .b(N2427), .c(N2340), .d(N2119), .e(N926), .O(N2631) );
nand5 gate738( .a(N2386), .b(N2427), .c(N2353), .d(N2104), .e(N926), .O(N2632) );
nand5 gate739( .a(N2386), .b(N2426), .c(N2340), .d(N2104), .e(N926), .O(N2633) );
nand5 gate740( .a(N2385), .b(N2427), .c(N2340), .d(N2104), .e(N926), .O(N2634) );
and5 gate741( .a(N2286), .b(N2427), .c(N2361), .d(N2129), .e(N1171), .O(N2639) );
and5 gate742( .a(N2297), .b(N2427), .c(N2361), .d(N2119), .e(N1171), .O(N2642) );
and5 gate743( .a(N2297), .b(N2427), .c(N2375), .d(N2104), .e(N1171), .O(N2645) );
and5 gate744( .a(N2297), .b(N2427), .c(N2340), .d(N2143), .e(N1171), .O(N2648) );
and5 gate745( .a(N2297), .b(N2427), .c(N2353), .d(N2129), .e(N1188), .O(N2651) );
and5 gate746( .a(N2386), .b(N2326), .c(N2361), .d(N2129), .e(N1188), .O(N2655) );
and5 gate747( .a(N2386), .b(N2326), .c(N2361), .d(N2119), .e(N1188), .O(N2658) );
and5 gate748( .a(N2386), .b(N2326), .c(N2375), .d(N2104), .e(N1188), .O(N2661) );
and5 gate749( .a(N2386), .b(N2326), .c(N2353), .d(N2129), .e(N1188), .O(N2664) );
nand2 gate750( .a(N2558), .b(N534), .O(N2669) );
inv1 gate751( .a(N2558), .O(N2670) );
nand2 gate752( .a(N2561), .b(N535), .O(N2671) );
inv1 gate753( .a(N2561), .O(N2672) );

  xor2  gate895(.a(N536), .b(N2564), .O(gate754inter0));
  nand2 gate896(.a(gate754inter0), .b(s_2), .O(gate754inter1));
  and2  gate897(.a(N536), .b(N2564), .O(gate754inter2));
  inv1  gate898(.a(s_2), .O(gate754inter3));
  inv1  gate899(.a(s_3), .O(gate754inter4));
  nand2 gate900(.a(gate754inter4), .b(gate754inter3), .O(gate754inter5));
  nor2  gate901(.a(gate754inter5), .b(gate754inter2), .O(gate754inter6));
  inv1  gate902(.a(N2564), .O(gate754inter7));
  inv1  gate903(.a(N536), .O(gate754inter8));
  nand2 gate904(.a(gate754inter8), .b(gate754inter7), .O(gate754inter9));
  nand2 gate905(.a(s_3), .b(gate754inter3), .O(gate754inter10));
  nor2  gate906(.a(gate754inter10), .b(gate754inter9), .O(gate754inter11));
  nor2  gate907(.a(gate754inter11), .b(gate754inter6), .O(gate754inter12));
  nand2 gate908(.a(gate754inter12), .b(gate754inter1), .O(N2673));
inv1 gate755( .a(N2564), .O(N2674) );

  xor2  gate1707(.a(N537), .b(N2567), .O(gate756inter0));
  nand2 gate1708(.a(gate756inter0), .b(s_118), .O(gate756inter1));
  and2  gate1709(.a(N537), .b(N2567), .O(gate756inter2));
  inv1  gate1710(.a(s_118), .O(gate756inter3));
  inv1  gate1711(.a(s_119), .O(gate756inter4));
  nand2 gate1712(.a(gate756inter4), .b(gate756inter3), .O(gate756inter5));
  nor2  gate1713(.a(gate756inter5), .b(gate756inter2), .O(gate756inter6));
  inv1  gate1714(.a(N2567), .O(gate756inter7));
  inv1  gate1715(.a(N537), .O(gate756inter8));
  nand2 gate1716(.a(gate756inter8), .b(gate756inter7), .O(gate756inter9));
  nand2 gate1717(.a(s_119), .b(gate756inter3), .O(gate756inter10));
  nor2  gate1718(.a(gate756inter10), .b(gate756inter9), .O(gate756inter11));
  nor2  gate1719(.a(gate756inter11), .b(gate756inter6), .O(gate756inter12));
  nand2 gate1720(.a(gate756inter12), .b(gate756inter1), .O(N2675));
inv1 gate757( .a(N2567), .O(N2676) );
nand2 gate758( .a(N2570), .b(N543), .O(N2682) );
inv1 gate759( .a(N2570), .O(N2683) );
nand2 gate760( .a(N2573), .b(N548), .O(N2688) );
inv1 gate761( .a(N2573), .O(N2689) );
nand2 gate762( .a(N2576), .b(N549), .O(N2690) );
inv1 gate763( .a(N2576), .O(N2691) );
and8 gate764( .a(N2627), .b(N2628), .c(N2629), .d(N2630), .e(N2631), .f(N2632), .g(N2633), .h(N2634), .O(N2710) );
nand2 gate765( .a(N343), .b(N2670), .O(N2720) );
nand2 gate766( .a(N346), .b(N2672), .O(N2721) );
nand2 gate767( .a(N349), .b(N2674), .O(N2722) );
nand2 gate768( .a(N352), .b(N2676), .O(N2723) );
nand2 gate769( .a(N2639), .b(N538), .O(N2724) );
inv1 gate770( .a(N2639), .O(N2725) );
nand2 gate771( .a(N2642), .b(N539), .O(N2726) );
inv1 gate772( .a(N2642), .O(N2727) );

  xor2  gate881(.a(N540), .b(N2645), .O(gate773inter0));
  nand2 gate882(.a(gate773inter0), .b(s_0), .O(gate773inter1));
  and2  gate883(.a(N540), .b(N2645), .O(gate773inter2));
  inv1  gate884(.a(s_0), .O(gate773inter3));
  inv1  gate885(.a(s_1), .O(gate773inter4));
  nand2 gate886(.a(gate773inter4), .b(gate773inter3), .O(gate773inter5));
  nor2  gate887(.a(gate773inter5), .b(gate773inter2), .O(gate773inter6));
  inv1  gate888(.a(N2645), .O(gate773inter7));
  inv1  gate889(.a(N540), .O(gate773inter8));
  nand2 gate890(.a(gate773inter8), .b(gate773inter7), .O(gate773inter9));
  nand2 gate891(.a(s_1), .b(gate773inter3), .O(gate773inter10));
  nor2  gate892(.a(gate773inter10), .b(gate773inter9), .O(gate773inter11));
  nor2  gate893(.a(gate773inter11), .b(gate773inter6), .O(gate773inter12));
  nand2 gate894(.a(gate773inter12), .b(gate773inter1), .O(N2728));
inv1 gate774( .a(N2645), .O(N2729) );
nand2 gate775( .a(N2648), .b(N541), .O(N2730) );
inv1 gate776( .a(N2648), .O(N2731) );
nand2 gate777( .a(N2651), .b(N542), .O(N2732) );
inv1 gate778( .a(N2651), .O(N2733) );
nand2 gate779( .a(N370), .b(N2683), .O(N2734) );

  xor2  gate1749(.a(N544), .b(N2655), .O(gate780inter0));
  nand2 gate1750(.a(gate780inter0), .b(s_124), .O(gate780inter1));
  and2  gate1751(.a(N544), .b(N2655), .O(gate780inter2));
  inv1  gate1752(.a(s_124), .O(gate780inter3));
  inv1  gate1753(.a(s_125), .O(gate780inter4));
  nand2 gate1754(.a(gate780inter4), .b(gate780inter3), .O(gate780inter5));
  nor2  gate1755(.a(gate780inter5), .b(gate780inter2), .O(gate780inter6));
  inv1  gate1756(.a(N2655), .O(gate780inter7));
  inv1  gate1757(.a(N544), .O(gate780inter8));
  nand2 gate1758(.a(gate780inter8), .b(gate780inter7), .O(gate780inter9));
  nand2 gate1759(.a(s_125), .b(gate780inter3), .O(gate780inter10));
  nor2  gate1760(.a(gate780inter10), .b(gate780inter9), .O(gate780inter11));
  nor2  gate1761(.a(gate780inter11), .b(gate780inter6), .O(gate780inter12));
  nand2 gate1762(.a(gate780inter12), .b(gate780inter1), .O(N2735));
inv1 gate781( .a(N2655), .O(N2736) );
nand2 gate782( .a(N2658), .b(N545), .O(N2737) );
inv1 gate783( .a(N2658), .O(N2738) );
nand2 gate784( .a(N2661), .b(N546), .O(N2739) );
inv1 gate785( .a(N2661), .O(N2740) );
nand2 gate786( .a(N2664), .b(N547), .O(N2741) );
inv1 gate787( .a(N2664), .O(N2742) );
nand2 gate788( .a(N385), .b(N2689), .O(N2743) );
nand2 gate789( .a(N388), .b(N2691), .O(N2744) );
nand8 gate790( .a(N2537), .b(N2540), .c(N2543), .d(N2546), .e(N2594), .f(N2597), .g(N2600), .h(N2603), .O(N2745) );
nand8 gate791( .a(N2606), .b(N2549), .c(N2611), .d(N2614), .e(N2617), .f(N2620), .g(N2552), .h(N2555), .O(N2746) );
and8 gate792( .a(N2537), .b(N2540), .c(N2543), .d(N2546), .e(N2594), .f(N2597), .g(N2600), .h(N2603), .O(N2747) );
and8 gate793( .a(N2606), .b(N2549), .c(N2611), .d(N2614), .e(N2617), .f(N2620), .g(N2552), .h(N2555), .O(N2750) );
nand2 gate794( .a(N2669), .b(N2720), .O(N2753) );
nand2 gate795( .a(N2671), .b(N2721), .O(N2754) );
nand2 gate796( .a(N2673), .b(N2722), .O(N2755) );
nand2 gate797( .a(N2675), .b(N2723), .O(N2756) );
nand2 gate798( .a(N355), .b(N2725), .O(N2757) );
nand2 gate799( .a(N358), .b(N2727), .O(N2758) );
nand2 gate800( .a(N361), .b(N2729), .O(N2759) );
nand2 gate801( .a(N364), .b(N2731), .O(N2760) );
nand2 gate802( .a(N367), .b(N2733), .O(N2761) );
nand2 gate803( .a(N2682), .b(N2734), .O(N2762) );
nand2 gate804( .a(N373), .b(N2736), .O(N2763) );

  xor2  gate1077(.a(N2738), .b(N376), .O(gate805inter0));
  nand2 gate1078(.a(gate805inter0), .b(s_28), .O(gate805inter1));
  and2  gate1079(.a(N2738), .b(N376), .O(gate805inter2));
  inv1  gate1080(.a(s_28), .O(gate805inter3));
  inv1  gate1081(.a(s_29), .O(gate805inter4));
  nand2 gate1082(.a(gate805inter4), .b(gate805inter3), .O(gate805inter5));
  nor2  gate1083(.a(gate805inter5), .b(gate805inter2), .O(gate805inter6));
  inv1  gate1084(.a(N376), .O(gate805inter7));
  inv1  gate1085(.a(N2738), .O(gate805inter8));
  nand2 gate1086(.a(gate805inter8), .b(gate805inter7), .O(gate805inter9));
  nand2 gate1087(.a(s_29), .b(gate805inter3), .O(gate805inter10));
  nor2  gate1088(.a(gate805inter10), .b(gate805inter9), .O(gate805inter11));
  nor2  gate1089(.a(gate805inter11), .b(gate805inter6), .O(gate805inter12));
  nand2 gate1090(.a(gate805inter12), .b(gate805inter1), .O(N2764));

  xor2  gate1735(.a(N2740), .b(N379), .O(gate806inter0));
  nand2 gate1736(.a(gate806inter0), .b(s_122), .O(gate806inter1));
  and2  gate1737(.a(N2740), .b(N379), .O(gate806inter2));
  inv1  gate1738(.a(s_122), .O(gate806inter3));
  inv1  gate1739(.a(s_123), .O(gate806inter4));
  nand2 gate1740(.a(gate806inter4), .b(gate806inter3), .O(gate806inter5));
  nor2  gate1741(.a(gate806inter5), .b(gate806inter2), .O(gate806inter6));
  inv1  gate1742(.a(N379), .O(gate806inter7));
  inv1  gate1743(.a(N2740), .O(gate806inter8));
  nand2 gate1744(.a(gate806inter8), .b(gate806inter7), .O(gate806inter9));
  nand2 gate1745(.a(s_123), .b(gate806inter3), .O(gate806inter10));
  nor2  gate1746(.a(gate806inter10), .b(gate806inter9), .O(gate806inter11));
  nor2  gate1747(.a(gate806inter11), .b(gate806inter6), .O(gate806inter12));
  nand2 gate1748(.a(gate806inter12), .b(gate806inter1), .O(N2765));
nand2 gate807( .a(N382), .b(N2742), .O(N2766) );
nand2 gate808( .a(N2688), .b(N2743), .O(N2767) );

  xor2  gate1021(.a(N2744), .b(N2690), .O(gate809inter0));
  nand2 gate1022(.a(gate809inter0), .b(s_20), .O(gate809inter1));
  and2  gate1023(.a(N2744), .b(N2690), .O(gate809inter2));
  inv1  gate1024(.a(s_20), .O(gate809inter3));
  inv1  gate1025(.a(s_21), .O(gate809inter4));
  nand2 gate1026(.a(gate809inter4), .b(gate809inter3), .O(gate809inter5));
  nor2  gate1027(.a(gate809inter5), .b(gate809inter2), .O(gate809inter6));
  inv1  gate1028(.a(N2690), .O(gate809inter7));
  inv1  gate1029(.a(N2744), .O(gate809inter8));
  nand2 gate1030(.a(gate809inter8), .b(gate809inter7), .O(gate809inter9));
  nand2 gate1031(.a(s_21), .b(gate809inter3), .O(gate809inter10));
  nor2  gate1032(.a(gate809inter10), .b(gate809inter9), .O(gate809inter11));
  nor2  gate1033(.a(gate809inter11), .b(gate809inter6), .O(gate809inter12));
  nand2 gate1034(.a(gate809inter12), .b(gate809inter1), .O(N2768));
and2 gate810( .a(N2745), .b(N275), .O(N2773) );
and2 gate811( .a(N2746), .b(N276), .O(N2776) );
nand2 gate812( .a(N2724), .b(N2757), .O(N2779) );
nand2 gate813( .a(N2726), .b(N2758), .O(N2780) );

  xor2  gate1665(.a(N2759), .b(N2728), .O(gate814inter0));
  nand2 gate1666(.a(gate814inter0), .b(s_112), .O(gate814inter1));
  and2  gate1667(.a(N2759), .b(N2728), .O(gate814inter2));
  inv1  gate1668(.a(s_112), .O(gate814inter3));
  inv1  gate1669(.a(s_113), .O(gate814inter4));
  nand2 gate1670(.a(gate814inter4), .b(gate814inter3), .O(gate814inter5));
  nor2  gate1671(.a(gate814inter5), .b(gate814inter2), .O(gate814inter6));
  inv1  gate1672(.a(N2728), .O(gate814inter7));
  inv1  gate1673(.a(N2759), .O(gate814inter8));
  nand2 gate1674(.a(gate814inter8), .b(gate814inter7), .O(gate814inter9));
  nand2 gate1675(.a(s_113), .b(gate814inter3), .O(gate814inter10));
  nor2  gate1676(.a(gate814inter10), .b(gate814inter9), .O(gate814inter11));
  nor2  gate1677(.a(gate814inter11), .b(gate814inter6), .O(gate814inter12));
  nand2 gate1678(.a(gate814inter12), .b(gate814inter1), .O(N2781));
nand2 gate815( .a(N2730), .b(N2760), .O(N2782) );
nand2 gate816( .a(N2732), .b(N2761), .O(N2783) );
nand2 gate817( .a(N2735), .b(N2763), .O(N2784) );
nand2 gate818( .a(N2737), .b(N2764), .O(N2785) );
nand2 gate819( .a(N2739), .b(N2765), .O(N2786) );
nand2 gate820( .a(N2741), .b(N2766), .O(N2787) );
and3 gate821( .a(N2747), .b(N2750), .c(N2710), .O(N2788) );
nand2 gate822( .a(N2747), .b(N2750), .O(N2789) );
and4 gate823( .a(N338), .b(N2279), .c(N99), .d(N2788), .O(N2800) );

  xor2  gate1245(.a(N2018), .b(N2773), .O(gate824inter0));
  nand2 gate1246(.a(gate824inter0), .b(s_52), .O(gate824inter1));
  and2  gate1247(.a(N2018), .b(N2773), .O(gate824inter2));
  inv1  gate1248(.a(s_52), .O(gate824inter3));
  inv1  gate1249(.a(s_53), .O(gate824inter4));
  nand2 gate1250(.a(gate824inter4), .b(gate824inter3), .O(gate824inter5));
  nor2  gate1251(.a(gate824inter5), .b(gate824inter2), .O(gate824inter6));
  inv1  gate1252(.a(N2773), .O(gate824inter7));
  inv1  gate1253(.a(N2018), .O(gate824inter8));
  nand2 gate1254(.a(gate824inter8), .b(gate824inter7), .O(gate824inter9));
  nand2 gate1255(.a(s_53), .b(gate824inter3), .O(gate824inter10));
  nor2  gate1256(.a(gate824inter10), .b(gate824inter9), .O(gate824inter11));
  nor2  gate1257(.a(gate824inter11), .b(gate824inter6), .O(gate824inter12));
  nand2 gate1258(.a(gate824inter12), .b(gate824inter1), .O(N2807));
inv1 gate825( .a(N2773), .O(N2808) );
nand2 gate826( .a(N2776), .b(N2019), .O(N2809) );
inv1 gate827( .a(N2776), .O(N2810) );
nor2 gate828( .a(N2384), .b(N2800), .O(N2811) );
and3 gate829( .a(N897), .b(N283), .c(N2789), .O(N2812) );
and3 gate830( .a(N76), .b(N283), .c(N2789), .O(N2815) );
and3 gate831( .a(N82), .b(N283), .c(N2789), .O(N2818) );
and3 gate832( .a(N85), .b(N283), .c(N2789), .O(N2821) );
and3 gate833( .a(N898), .b(N283), .c(N2789), .O(N2824) );
nand2 gate834( .a(N1965), .b(N2808), .O(N2827) );
nand2 gate835( .a(N1968), .b(N2810), .O(N2828) );
and3 gate836( .a(N79), .b(N283), .c(N2789), .O(N2829) );
nand2 gate837( .a(N2807), .b(N2827), .O(N2843) );
nand2 gate838( .a(N2809), .b(N2828), .O(N2846) );

  xor2  gate1637(.a(N2076), .b(N2812), .O(gate839inter0));
  nand2 gate1638(.a(gate839inter0), .b(s_108), .O(gate839inter1));
  and2  gate1639(.a(N2076), .b(N2812), .O(gate839inter2));
  inv1  gate1640(.a(s_108), .O(gate839inter3));
  inv1  gate1641(.a(s_109), .O(gate839inter4));
  nand2 gate1642(.a(gate839inter4), .b(gate839inter3), .O(gate839inter5));
  nor2  gate1643(.a(gate839inter5), .b(gate839inter2), .O(gate839inter6));
  inv1  gate1644(.a(N2812), .O(gate839inter7));
  inv1  gate1645(.a(N2076), .O(gate839inter8));
  nand2 gate1646(.a(gate839inter8), .b(gate839inter7), .O(gate839inter9));
  nand2 gate1647(.a(s_109), .b(gate839inter3), .O(gate839inter10));
  nor2  gate1648(.a(gate839inter10), .b(gate839inter9), .O(gate839inter11));
  nor2  gate1649(.a(gate839inter11), .b(gate839inter6), .O(gate839inter12));
  nand2 gate1650(.a(gate839inter12), .b(gate839inter1), .O(N2850));
nand2 gate840( .a(N2815), .b(N2077), .O(N2851) );
nand2 gate841( .a(N2818), .b(N1915), .O(N2852) );
nand2 gate842( .a(N2821), .b(N1857), .O(N2853) );
nand2 gate843( .a(N2824), .b(N1938), .O(N2854) );
inv1 gate844( .a(N2812), .O(N2857) );
inv1 gate845( .a(N2815), .O(N2858) );
inv1 gate846( .a(N2818), .O(N2859) );
inv1 gate847( .a(N2821), .O(N2860) );
inv1 gate848( .a(N2824), .O(N2861) );
inv1 gate849( .a(N2829), .O(N2862) );
nand2 gate850( .a(N2829), .b(N1985), .O(N2863) );

  xor2  gate1441(.a(N2857), .b(N2052), .O(gate851inter0));
  nand2 gate1442(.a(gate851inter0), .b(s_80), .O(gate851inter1));
  and2  gate1443(.a(N2857), .b(N2052), .O(gate851inter2));
  inv1  gate1444(.a(s_80), .O(gate851inter3));
  inv1  gate1445(.a(s_81), .O(gate851inter4));
  nand2 gate1446(.a(gate851inter4), .b(gate851inter3), .O(gate851inter5));
  nor2  gate1447(.a(gate851inter5), .b(gate851inter2), .O(gate851inter6));
  inv1  gate1448(.a(N2052), .O(gate851inter7));
  inv1  gate1449(.a(N2857), .O(gate851inter8));
  nand2 gate1450(.a(gate851inter8), .b(gate851inter7), .O(gate851inter9));
  nand2 gate1451(.a(s_81), .b(gate851inter3), .O(gate851inter10));
  nor2  gate1452(.a(gate851inter10), .b(gate851inter9), .O(gate851inter11));
  nor2  gate1453(.a(gate851inter11), .b(gate851inter6), .O(gate851inter12));
  nand2 gate1454(.a(gate851inter12), .b(gate851inter1), .O(N2866));

  xor2  gate1315(.a(N2858), .b(N2055), .O(gate852inter0));
  nand2 gate1316(.a(gate852inter0), .b(s_62), .O(gate852inter1));
  and2  gate1317(.a(N2858), .b(N2055), .O(gate852inter2));
  inv1  gate1318(.a(s_62), .O(gate852inter3));
  inv1  gate1319(.a(s_63), .O(gate852inter4));
  nand2 gate1320(.a(gate852inter4), .b(gate852inter3), .O(gate852inter5));
  nor2  gate1321(.a(gate852inter5), .b(gate852inter2), .O(gate852inter6));
  inv1  gate1322(.a(N2055), .O(gate852inter7));
  inv1  gate1323(.a(N2858), .O(gate852inter8));
  nand2 gate1324(.a(gate852inter8), .b(gate852inter7), .O(gate852inter9));
  nand2 gate1325(.a(s_63), .b(gate852inter3), .O(gate852inter10));
  nor2  gate1326(.a(gate852inter10), .b(gate852inter9), .O(gate852inter11));
  nor2  gate1327(.a(gate852inter11), .b(gate852inter6), .O(gate852inter12));
  nand2 gate1328(.a(gate852inter12), .b(gate852inter1), .O(N2867));
nand2 gate853( .a(N1866), .b(N2859), .O(N2868) );

  xor2  gate909(.a(N2860), .b(N1818), .O(gate854inter0));
  nand2 gate910(.a(gate854inter0), .b(s_4), .O(gate854inter1));
  and2  gate911(.a(N2860), .b(N1818), .O(gate854inter2));
  inv1  gate912(.a(s_4), .O(gate854inter3));
  inv1  gate913(.a(s_5), .O(gate854inter4));
  nand2 gate914(.a(gate854inter4), .b(gate854inter3), .O(gate854inter5));
  nor2  gate915(.a(gate854inter5), .b(gate854inter2), .O(gate854inter6));
  inv1  gate916(.a(N1818), .O(gate854inter7));
  inv1  gate917(.a(N2860), .O(gate854inter8));
  nand2 gate918(.a(gate854inter8), .b(gate854inter7), .O(gate854inter9));
  nand2 gate919(.a(s_5), .b(gate854inter3), .O(gate854inter10));
  nor2  gate920(.a(gate854inter10), .b(gate854inter9), .O(gate854inter11));
  nor2  gate921(.a(gate854inter11), .b(gate854inter6), .O(gate854inter12));
  nand2 gate922(.a(gate854inter12), .b(gate854inter1), .O(N2869));
nand2 gate855( .a(N1902), .b(N2861), .O(N2870) );
nand2 gate856( .a(N2843), .b(N886), .O(N2871) );
inv1 gate857( .a(N2843), .O(N2872) );
nand2 gate858( .a(N2846), .b(N887), .O(N2873) );
inv1 gate859( .a(N2846), .O(N2874) );
nand2 gate860( .a(N1933), .b(N2862), .O(N2875) );
nand2 gate861( .a(N2866), .b(N2850), .O(N2876) );

  xor2  gate1273(.a(N2851), .b(N2867), .O(gate862inter0));
  nand2 gate1274(.a(gate862inter0), .b(s_56), .O(gate862inter1));
  and2  gate1275(.a(N2851), .b(N2867), .O(gate862inter2));
  inv1  gate1276(.a(s_56), .O(gate862inter3));
  inv1  gate1277(.a(s_57), .O(gate862inter4));
  nand2 gate1278(.a(gate862inter4), .b(gate862inter3), .O(gate862inter5));
  nor2  gate1279(.a(gate862inter5), .b(gate862inter2), .O(gate862inter6));
  inv1  gate1280(.a(N2867), .O(gate862inter7));
  inv1  gate1281(.a(N2851), .O(gate862inter8));
  nand2 gate1282(.a(gate862inter8), .b(gate862inter7), .O(gate862inter9));
  nand2 gate1283(.a(s_57), .b(gate862inter3), .O(gate862inter10));
  nor2  gate1284(.a(gate862inter10), .b(gate862inter9), .O(gate862inter11));
  nor2  gate1285(.a(gate862inter11), .b(gate862inter6), .O(gate862inter12));
  nand2 gate1286(.a(gate862inter12), .b(gate862inter1), .O(N2877));
nand2 gate863( .a(N2868), .b(N2852), .O(N2878) );
nand2 gate864( .a(N2869), .b(N2853), .O(N2879) );
nand2 gate865( .a(N2870), .b(N2854), .O(N2880) );
nand2 gate866( .a(N682), .b(N2872), .O(N2881) );
nand2 gate867( .a(N685), .b(N2874), .O(N2882) );
nand2 gate868( .a(N2875), .b(N2863), .O(N2883) );
and2 gate869( .a(N2876), .b(N550), .O(N2886) );
and2 gate870( .a(N551), .b(N2877), .O(N2887) );
and2 gate871( .a(N553), .b(N2878), .O(N2888) );
and2 gate872( .a(N2879), .b(N554), .O(N2889) );
and2 gate873( .a(N555), .b(N2880), .O(N2890) );
nand2 gate874( .a(N2871), .b(N2881), .O(N2891) );
nand2 gate875( .a(N2873), .b(N2882), .O(N2892) );
nand2 gate876( .a(N2883), .b(N1461), .O(N2895) );
inv1 gate877( .a(N2883), .O(N2896) );
nand2 gate878( .a(N1383), .b(N2896), .O(N2897) );
nand2 gate879( .a(N2895), .b(N2897), .O(N2898) );
and2 gate880( .a(N2898), .b(N552), .O(N2899) );

endmodule