module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);

input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;//RE__PI;

input s_0,s_1;//RE__ALLOW(00,01,10,11);
input s_2,s_3;//RE__ALLOW(00,01,10,11);
input s_4,s_5;//RE__ALLOW(00,01,10,11);
input s_6,s_7;//RE__ALLOW(00,01,10,11);
input s_8,s_9;//RE__ALLOW(00,01,10,11);
input s_10,s_11;//RE__ALLOW(00,01,10,11);
input s_12,s_13;//RE__ALLOW(00,01,10,11);
input s_14,s_15;//RE__ALLOW(00,01,10,11);
input s_16,s_17;//RE__ALLOW(00,01,10,11);
input s_18,s_19;//RE__ALLOW(00,01,10,11);
input s_20,s_21;//RE__ALLOW(00,01,10,11);
input s_22,s_23;//RE__ALLOW(00,01,10,11);
input s_24,s_25;//RE__ALLOW(00,01,10,11);
input s_26,s_27;//RE__ALLOW(00,01,10,11);
input s_28,s_29;//RE__ALLOW(00,01,10,11);
input s_30,s_31;//RE__ALLOW(00,01,10,11);
input s_32,s_33;//RE__ALLOW(00,01,10,11);
input s_34,s_35;//RE__ALLOW(00,01,10,11);
input s_36,s_37;//RE__ALLOW(00,01,10,11);
input s_38,s_39;//RE__ALLOW(00,01,10,11);
input s_40,s_41;//RE__ALLOW(00,01,10,11);
input s_42,s_43;//RE__ALLOW(00,01,10,11);
input s_44,s_45;//RE__ALLOW(00,01,10,11);
input s_46,s_47;//RE__ALLOW(00,01,10,11);
input s_48,s_49;//RE__ALLOW(00,01,10,11);
input s_50,s_51;//RE__ALLOW(00,01,10,11);
input s_52,s_53;//RE__ALLOW(00,01,10,11);
input s_54,s_55;//RE__ALLOW(00,01,10,11);
input s_56,s_57;//RE__ALLOW(00,01,10,11);
input s_58,s_59;//RE__ALLOW(00,01,10,11);
input s_60,s_61;//RE__ALLOW(00,01,10,11);
input s_62,s_63;//RE__ALLOW(00,01,10,11);
input s_64,s_65;//RE__ALLOW(00,01,10,11);
input s_66,s_67;//RE__ALLOW(00,01,10,11);
input s_68,s_69;//RE__ALLOW(00,01,10,11);
input s_70,s_71;//RE__ALLOW(00,01,10,11);
input s_72,s_73;//RE__ALLOW(00,01,10,11);
input s_74,s_75;//RE__ALLOW(00,01,10,11);
input s_76,s_77;//RE__ALLOW(00,01,10,11);
input s_78,s_79;//RE__ALLOW(00,01,10,11);
input s_80,s_81;//RE__ALLOW(00,01,10,11);
input s_82,s_83;//RE__ALLOW(00,01,10,11);
input s_84,s_85;//RE__ALLOW(00,01,10,11);
input s_86,s_87;//RE__ALLOW(00,01,10,11);
input s_88,s_89;//RE__ALLOW(00,01,10,11);
input s_90,s_91;//RE__ALLOW(00,01,10,11);
input s_92,s_93;//RE__ALLOW(00,01,10,11);
input s_94,s_95;//RE__ALLOW(00,01,10,11);
input s_96,s_97;//RE__ALLOW(00,01,10,11);
input s_98,s_99;//RE__ALLOW(00,01,10,11);
input s_100,s_101;//RE__ALLOW(00,01,10,11);
input s_102,s_103;//RE__ALLOW(00,01,10,11);
input s_104,s_105;//RE__ALLOW(00,01,10,11);
input s_106,s_107;//RE__ALLOW(00,01,10,11);
input s_108,s_109;//RE__ALLOW(00,01,10,11);
input s_110,s_111;//RE__ALLOW(00,01,10,11);
input s_112,s_113;//RE__ALLOW(00,01,10,11);
input s_114,s_115;//RE__ALLOW(00,01,10,11);
input s_116,s_117;//RE__ALLOW(00,01,10,11);
input s_118,s_119;//RE__ALLOW(00,01,10,11);
input s_120,s_121;//RE__ALLOW(00,01,10,11);
input s_122,s_123;//RE__ALLOW(00,01,10,11);
input s_124,s_125;//RE__ALLOW(00,01,10,11);
input s_126,s_127;//RE__ALLOW(00,01,10,11);
input s_128,s_129;//RE__ALLOW(00,01,10,11);
input s_130,s_131;//RE__ALLOW(00,01,10,11);
input s_132,s_133;//RE__ALLOW(00,01,10,11);
input s_134,s_135;//RE__ALLOW(00,01,10,11);
input s_136,s_137;//RE__ALLOW(00,01,10,11);
input s_138,s_139;//RE__ALLOW(00,01,10,11);
input s_140,s_141;//RE__ALLOW(00,01,10,11);
input s_142,s_143;//RE__ALLOW(00,01,10,11);
input s_144,s_145;//RE__ALLOW(00,01,10,11);
input s_146,s_147;//RE__ALLOW(00,01,10,11);
input s_148,s_149;//RE__ALLOW(00,01,10,11);
input s_150,s_151;//RE__ALLOW(00,01,10,11);
input s_152,s_153;//RE__ALLOW(00,01,10,11);
input s_154,s_155;//RE__ALLOW(00,01,10,11);
input s_156,s_157;//RE__ALLOW(00,01,10,11);
input s_158,s_159;//RE__ALLOW(00,01,10,11);
input s_160,s_161;//RE__ALLOW(00,01,10,11);
input s_162,s_163;//RE__ALLOW(00,01,10,11);
input s_164,s_165;//RE__ALLOW(00,01,10,11);
input s_166,s_167;//RE__ALLOW(00,01,10,11);
input s_168,s_169;//RE__ALLOW(00,01,10,11);
input s_170,s_171;//RE__ALLOW(00,01,10,11);
input s_172,s_173;//RE__ALLOW(00,01,10,11);
input s_174,s_175;//RE__ALLOW(00,01,10,11);
input s_176,s_177;//RE__ALLOW(00,01,10,11);
input s_178,s_179;//RE__ALLOW(00,01,10,11);
input s_180,s_181;//RE__ALLOW(00,01,10,11);
input s_182,s_183;//RE__ALLOW(00,01,10,11);
input s_184,s_185;//RE__ALLOW(00,01,10,11);
input s_186,s_187;//RE__ALLOW(00,01,10,11);
input s_188,s_189;//RE__ALLOW(00,01,10,11);
input s_190,s_191;//RE__ALLOW(00,01,10,11);
input s_192,s_193;//RE__ALLOW(00,01,10,11);
input s_194,s_195;//RE__ALLOW(00,01,10,11);
input s_196,s_197;//RE__ALLOW(00,01,10,11);
input s_198,s_199;//RE__ALLOW(00,01,10,11);
input s_200,s_201;//RE__ALLOW(00,01,10,11);
input s_202,s_203;//RE__ALLOW(00,01,10,11);
input s_204,s_205;//RE__ALLOW(00,01,10,11);
input s_206,s_207;//RE__ALLOW(00,01,10,11);
input s_208,s_209;//RE__ALLOW(00,01,10,11);
input s_210,s_211;//RE__ALLOW(00,01,10,11);
input s_212,s_213;//RE__ALLOW(00,01,10,11);
input s_214,s_215;//RE__ALLOW(00,01,10,11);
input s_216,s_217;//RE__ALLOW(00,01,10,11);
input s_218,s_219;//RE__ALLOW(00,01,10,11);
input s_220,s_221;//RE__ALLOW(00,01,10,11);
input s_222,s_223;//RE__ALLOW(00,01,10,11);
input s_224,s_225;//RE__ALLOW(00,01,10,11);
input s_226,s_227;//RE__ALLOW(00,01,10,11);
input s_228,s_229;//RE__ALLOW(00,01,10,11);
input s_230,s_231;//RE__ALLOW(00,01,10,11);
input s_232,s_233;//RE__ALLOW(00,01,10,11);
input s_234,s_235;//RE__ALLOW(00,01,10,11);
input s_236,s_237;//RE__ALLOW(00,01,10,11);
input s_238,s_239;//RE__ALLOW(00,01,10,11);
input s_240,s_241;//RE__ALLOW(00,01,10,11);
input s_242,s_243;//RE__ALLOW(00,01,10,11);
input s_244,s_245;//RE__ALLOW(00,01,10,11);
input s_246,s_247;//RE__ALLOW(00,01,10,11);
input s_248,s_249;//RE__ALLOW(00,01,10,11);
input s_250,s_251;//RE__ALLOW(00,01,10,11);
input s_252,s_253;//RE__ALLOW(00,01,10,11);
input s_254,s_255;//RE__ALLOW(00,01,10,11);
input s_256,s_257;//RE__ALLOW(00,01,10,11);
input s_258,s_259;//RE__ALLOW(00,01,10,11);
input s_260,s_261;//RE__ALLOW(00,01,10,11);
input s_262,s_263;//RE__ALLOW(00,01,10,11);
input s_264,s_265;//RE__ALLOW(00,01,10,11);
input s_266,s_267;//RE__ALLOW(00,01,10,11);
input s_268,s_269;//RE__ALLOW(00,01,10,11);
input s_270,s_271;//RE__ALLOW(00,01,10,11);
input s_272,s_273;//RE__ALLOW(00,01,10,11);
input s_274,s_275;//RE__ALLOW(00,01,10,11);
input s_276,s_277;//RE__ALLOW(00,01,10,11);
input s_278,s_279;//RE__ALLOW(00,01,10,11);
input s_280,s_281;//RE__ALLOW(00,01,10,11);
input s_282,s_283;//RE__ALLOW(00,01,10,11);
input s_284,s_285;//RE__ALLOW(00,01,10,11);
input s_286,s_287;//RE__ALLOW(00,01,10,11);
input s_288,s_289;//RE__ALLOW(00,01,10,11);
input s_290,s_291;//RE__ALLOW(00,01,10,11);
input s_292,s_293;//RE__ALLOW(00,01,10,11);
input s_294,s_295;//RE__ALLOW(00,01,10,11);
input s_296,s_297;//RE__ALLOW(00,01,10,11);
input s_298,s_299;//RE__ALLOW(00,01,10,11);
input s_300,s_301;//RE__ALLOW(00,01,10,11);
input s_302,s_303;//RE__ALLOW(00,01,10,11);
input s_304,s_305;//RE__ALLOW(00,01,10,11);
input s_306,s_307;//RE__ALLOW(00,01,10,11);
input s_308,s_309;//RE__ALLOW(00,01,10,11);
input s_310,s_311;//RE__ALLOW(00,01,10,11);
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;

  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate84inter0, gate84inter1, gate84inter2, gate84inter3, gate84inter4, gate84inter5, gate84inter6, gate84inter7, gate84inter8, gate84inter9, gate84inter10, gate84inter11, gate84inter12, gate190inter0, gate190inter1, gate190inter2, gate190inter3, gate190inter4, gate190inter5, gate190inter6, gate190inter7, gate190inter8, gate190inter9, gate190inter10, gate190inter11, gate190inter12, gate15inter0, gate15inter1, gate15inter2, gate15inter3, gate15inter4, gate15inter5, gate15inter6, gate15inter7, gate15inter8, gate15inter9, gate15inter10, gate15inter11, gate15inter12, gate229inter0, gate229inter1, gate229inter2, gate229inter3, gate229inter4, gate229inter5, gate229inter6, gate229inter7, gate229inter8, gate229inter9, gate229inter10, gate229inter11, gate229inter12, gate452inter0, gate452inter1, gate452inter2, gate452inter3, gate452inter4, gate452inter5, gate452inter6, gate452inter7, gate452inter8, gate452inter9, gate452inter10, gate452inter11, gate452inter12, gate493inter0, gate493inter1, gate493inter2, gate493inter3, gate493inter4, gate493inter5, gate493inter6, gate493inter7, gate493inter8, gate493inter9, gate493inter10, gate493inter11, gate493inter12, gate112inter0, gate112inter1, gate112inter2, gate112inter3, gate112inter4, gate112inter5, gate112inter6, gate112inter7, gate112inter8, gate112inter9, gate112inter10, gate112inter11, gate112inter12, gate172inter0, gate172inter1, gate172inter2, gate172inter3, gate172inter4, gate172inter5, gate172inter6, gate172inter7, gate172inter8, gate172inter9, gate172inter10, gate172inter11, gate172inter12, gate415inter0, gate415inter1, gate415inter2, gate415inter3, gate415inter4, gate415inter5, gate415inter6, gate415inter7, gate415inter8, gate415inter9, gate415inter10, gate415inter11, gate415inter12, gate25inter0, gate25inter1, gate25inter2, gate25inter3, gate25inter4, gate25inter5, gate25inter6, gate25inter7, gate25inter8, gate25inter9, gate25inter10, gate25inter11, gate25inter12, gate259inter0, gate259inter1, gate259inter2, gate259inter3, gate259inter4, gate259inter5, gate259inter6, gate259inter7, gate259inter8, gate259inter9, gate259inter10, gate259inter11, gate259inter12, gate119inter0, gate119inter1, gate119inter2, gate119inter3, gate119inter4, gate119inter5, gate119inter6, gate119inter7, gate119inter8, gate119inter9, gate119inter10, gate119inter11, gate119inter12, gate466inter0, gate466inter1, gate466inter2, gate466inter3, gate466inter4, gate466inter5, gate466inter6, gate466inter7, gate466inter8, gate466inter9, gate466inter10, gate466inter11, gate466inter12, gate448inter0, gate448inter1, gate448inter2, gate448inter3, gate448inter4, gate448inter5, gate448inter6, gate448inter7, gate448inter8, gate448inter9, gate448inter10, gate448inter11, gate448inter12, gate499inter0, gate499inter1, gate499inter2, gate499inter3, gate499inter4, gate499inter5, gate499inter6, gate499inter7, gate499inter8, gate499inter9, gate499inter10, gate499inter11, gate499inter12, gate416inter0, gate416inter1, gate416inter2, gate416inter3, gate416inter4, gate416inter5, gate416inter6, gate416inter7, gate416inter8, gate416inter9, gate416inter10, gate416inter11, gate416inter12, gate49inter0, gate49inter1, gate49inter2, gate49inter3, gate49inter4, gate49inter5, gate49inter6, gate49inter7, gate49inter8, gate49inter9, gate49inter10, gate49inter11, gate49inter12, gate45inter0, gate45inter1, gate45inter2, gate45inter3, gate45inter4, gate45inter5, gate45inter6, gate45inter7, gate45inter8, gate45inter9, gate45inter10, gate45inter11, gate45inter12, gate243inter0, gate243inter1, gate243inter2, gate243inter3, gate243inter4, gate243inter5, gate243inter6, gate243inter7, gate243inter8, gate243inter9, gate243inter10, gate243inter11, gate243inter12, gate36inter0, gate36inter1, gate36inter2, gate36inter3, gate36inter4, gate36inter5, gate36inter6, gate36inter7, gate36inter8, gate36inter9, gate36inter10, gate36inter11, gate36inter12, gate220inter0, gate220inter1, gate220inter2, gate220inter3, gate220inter4, gate220inter5, gate220inter6, gate220inter7, gate220inter8, gate220inter9, gate220inter10, gate220inter11, gate220inter12, gate64inter0, gate64inter1, gate64inter2, gate64inter3, gate64inter4, gate64inter5, gate64inter6, gate64inter7, gate64inter8, gate64inter9, gate64inter10, gate64inter11, gate64inter12, gate504inter0, gate504inter1, gate504inter2, gate504inter3, gate504inter4, gate504inter5, gate504inter6, gate504inter7, gate504inter8, gate504inter9, gate504inter10, gate504inter11, gate504inter12, gate261inter0, gate261inter1, gate261inter2, gate261inter3, gate261inter4, gate261inter5, gate261inter6, gate261inter7, gate261inter8, gate261inter9, gate261inter10, gate261inter11, gate261inter12, gate295inter0, gate295inter1, gate295inter2, gate295inter3, gate295inter4, gate295inter5, gate295inter6, gate295inter7, gate295inter8, gate295inter9, gate295inter10, gate295inter11, gate295inter12, gate460inter0, gate460inter1, gate460inter2, gate460inter3, gate460inter4, gate460inter5, gate460inter6, gate460inter7, gate460inter8, gate460inter9, gate460inter10, gate460inter11, gate460inter12, gate238inter0, gate238inter1, gate238inter2, gate238inter3, gate238inter4, gate238inter5, gate238inter6, gate238inter7, gate238inter8, gate238inter9, gate238inter10, gate238inter11, gate238inter12, gate277inter0, gate277inter1, gate277inter2, gate277inter3, gate277inter4, gate277inter5, gate277inter6, gate277inter7, gate277inter8, gate277inter9, gate277inter10, gate277inter11, gate277inter12, gate126inter0, gate126inter1, gate126inter2, gate126inter3, gate126inter4, gate126inter5, gate126inter6, gate126inter7, gate126inter8, gate126inter9, gate126inter10, gate126inter11, gate126inter12, gate501inter0, gate501inter1, gate501inter2, gate501inter3, gate501inter4, gate501inter5, gate501inter6, gate501inter7, gate501inter8, gate501inter9, gate501inter10, gate501inter11, gate501inter12, gate476inter0, gate476inter1, gate476inter2, gate476inter3, gate476inter4, gate476inter5, gate476inter6, gate476inter7, gate476inter8, gate476inter9, gate476inter10, gate476inter11, gate476inter12, gate213inter0, gate213inter1, gate213inter2, gate213inter3, gate213inter4, gate213inter5, gate213inter6, gate213inter7, gate213inter8, gate213inter9, gate213inter10, gate213inter11, gate213inter12, gate188inter0, gate188inter1, gate188inter2, gate188inter3, gate188inter4, gate188inter5, gate188inter6, gate188inter7, gate188inter8, gate188inter9, gate188inter10, gate188inter11, gate188inter12, gate478inter0, gate478inter1, gate478inter2, gate478inter3, gate478inter4, gate478inter5, gate478inter6, gate478inter7, gate478inter8, gate478inter9, gate478inter10, gate478inter11, gate478inter12, gate490inter0, gate490inter1, gate490inter2, gate490inter3, gate490inter4, gate490inter5, gate490inter6, gate490inter7, gate490inter8, gate490inter9, gate490inter10, gate490inter11, gate490inter12, gate471inter0, gate471inter1, gate471inter2, gate471inter3, gate471inter4, gate471inter5, gate471inter6, gate471inter7, gate471inter8, gate471inter9, gate471inter10, gate471inter11, gate471inter12, gate450inter0, gate450inter1, gate450inter2, gate450inter3, gate450inter4, gate450inter5, gate450inter6, gate450inter7, gate450inter8, gate450inter9, gate450inter10, gate450inter11, gate450inter12, gate475inter0, gate475inter1, gate475inter2, gate475inter3, gate475inter4, gate475inter5, gate475inter6, gate475inter7, gate475inter8, gate475inter9, gate475inter10, gate475inter11, gate475inter12, gate152inter0, gate152inter1, gate152inter2, gate152inter3, gate152inter4, gate152inter5, gate152inter6, gate152inter7, gate152inter8, gate152inter9, gate152inter10, gate152inter11, gate152inter12, gate245inter0, gate245inter1, gate245inter2, gate245inter3, gate245inter4, gate245inter5, gate245inter6, gate245inter7, gate245inter8, gate245inter9, gate245inter10, gate245inter11, gate245inter12, gate403inter0, gate403inter1, gate403inter2, gate403inter3, gate403inter4, gate403inter5, gate403inter6, gate403inter7, gate403inter8, gate403inter9, gate403inter10, gate403inter11, gate403inter12, gate254inter0, gate254inter1, gate254inter2, gate254inter3, gate254inter4, gate254inter5, gate254inter6, gate254inter7, gate254inter8, gate254inter9, gate254inter10, gate254inter11, gate254inter12, gate509inter0, gate509inter1, gate509inter2, gate509inter3, gate509inter4, gate509inter5, gate509inter6, gate509inter7, gate509inter8, gate509inter9, gate509inter10, gate509inter11, gate509inter12, gate86inter0, gate86inter1, gate86inter2, gate86inter3, gate86inter4, gate86inter5, gate86inter6, gate86inter7, gate86inter8, gate86inter9, gate86inter10, gate86inter11, gate86inter12, gate437inter0, gate437inter1, gate437inter2, gate437inter3, gate437inter4, gate437inter5, gate437inter6, gate437inter7, gate437inter8, gate437inter9, gate437inter10, gate437inter11, gate437inter12, gate17inter0, gate17inter1, gate17inter2, gate17inter3, gate17inter4, gate17inter5, gate17inter6, gate17inter7, gate17inter8, gate17inter9, gate17inter10, gate17inter11, gate17inter12, gate489inter0, gate489inter1, gate489inter2, gate489inter3, gate489inter4, gate489inter5, gate489inter6, gate489inter7, gate489inter8, gate489inter9, gate489inter10, gate489inter11, gate489inter12, gate255inter0, gate255inter1, gate255inter2, gate255inter3, gate255inter4, gate255inter5, gate255inter6, gate255inter7, gate255inter8, gate255inter9, gate255inter10, gate255inter11, gate255inter12, gate407inter0, gate407inter1, gate407inter2, gate407inter3, gate407inter4, gate407inter5, gate407inter6, gate407inter7, gate407inter8, gate407inter9, gate407inter10, gate407inter11, gate407inter12, gate197inter0, gate197inter1, gate197inter2, gate197inter3, gate197inter4, gate197inter5, gate197inter6, gate197inter7, gate197inter8, gate197inter9, gate197inter10, gate197inter11, gate197inter12, gate194inter0, gate194inter1, gate194inter2, gate194inter3, gate194inter4, gate194inter5, gate194inter6, gate194inter7, gate194inter8, gate194inter9, gate194inter10, gate194inter11, gate194inter12, gate56inter0, gate56inter1, gate56inter2, gate56inter3, gate56inter4, gate56inter5, gate56inter6, gate56inter7, gate56inter8, gate56inter9, gate56inter10, gate56inter11, gate56inter12, gate420inter0, gate420inter1, gate420inter2, gate420inter3, gate420inter4, gate420inter5, gate420inter6, gate420inter7, gate420inter8, gate420inter9, gate420inter10, gate420inter11, gate420inter12, gate453inter0, gate453inter1, gate453inter2, gate453inter3, gate453inter4, gate453inter5, gate453inter6, gate453inter7, gate453inter8, gate453inter9, gate453inter10, gate453inter11, gate453inter12, gate162inter0, gate162inter1, gate162inter2, gate162inter3, gate162inter4, gate162inter5, gate162inter6, gate162inter7, gate162inter8, gate162inter9, gate162inter10, gate162inter11, gate162inter12, gate494inter0, gate494inter1, gate494inter2, gate494inter3, gate494inter4, gate494inter5, gate494inter6, gate494inter7, gate494inter8, gate494inter9, gate494inter10, gate494inter11, gate494inter12, gate201inter0, gate201inter1, gate201inter2, gate201inter3, gate201inter4, gate201inter5, gate201inter6, gate201inter7, gate201inter8, gate201inter9, gate201inter10, gate201inter11, gate201inter12, gate100inter0, gate100inter1, gate100inter2, gate100inter3, gate100inter4, gate100inter5, gate100inter6, gate100inter7, gate100inter8, gate100inter9, gate100inter10, gate100inter11, gate100inter12, gate165inter0, gate165inter1, gate165inter2, gate165inter3, gate165inter4, gate165inter5, gate165inter6, gate165inter7, gate165inter8, gate165inter9, gate165inter10, gate165inter11, gate165inter12, gate278inter0, gate278inter1, gate278inter2, gate278inter3, gate278inter4, gate278inter5, gate278inter6, gate278inter7, gate278inter8, gate278inter9, gate278inter10, gate278inter11, gate278inter12, gate429inter0, gate429inter1, gate429inter2, gate429inter3, gate429inter4, gate429inter5, gate429inter6, gate429inter7, gate429inter8, gate429inter9, gate429inter10, gate429inter11, gate429inter12, gate474inter0, gate474inter1, gate474inter2, gate474inter3, gate474inter4, gate474inter5, gate474inter6, gate474inter7, gate474inter8, gate474inter9, gate474inter10, gate474inter11, gate474inter12, gate73inter0, gate73inter1, gate73inter2, gate73inter3, gate73inter4, gate73inter5, gate73inter6, gate73inter7, gate73inter8, gate73inter9, gate73inter10, gate73inter11, gate73inter12, gate392inter0, gate392inter1, gate392inter2, gate392inter3, gate392inter4, gate392inter5, gate392inter6, gate392inter7, gate392inter8, gate392inter9, gate392inter10, gate392inter11, gate392inter12, gate426inter0, gate426inter1, gate426inter2, gate426inter3, gate426inter4, gate426inter5, gate426inter6, gate426inter7, gate426inter8, gate426inter9, gate426inter10, gate426inter11, gate426inter12, gate11inter0, gate11inter1, gate11inter2, gate11inter3, gate11inter4, gate11inter5, gate11inter6, gate11inter7, gate11inter8, gate11inter9, gate11inter10, gate11inter11, gate11inter12, gate406inter0, gate406inter1, gate406inter2, gate406inter3, gate406inter4, gate406inter5, gate406inter6, gate406inter7, gate406inter8, gate406inter9, gate406inter10, gate406inter11, gate406inter12, gate61inter0, gate61inter1, gate61inter2, gate61inter3, gate61inter4, gate61inter5, gate61inter6, gate61inter7, gate61inter8, gate61inter9, gate61inter10, gate61inter11, gate61inter12, gate198inter0, gate198inter1, gate198inter2, gate198inter3, gate198inter4, gate198inter5, gate198inter6, gate198inter7, gate198inter8, gate198inter9, gate198inter10, gate198inter11, gate198inter12, gate247inter0, gate247inter1, gate247inter2, gate247inter3, gate247inter4, gate247inter5, gate247inter6, gate247inter7, gate247inter8, gate247inter9, gate247inter10, gate247inter11, gate247inter12, gate268inter0, gate268inter1, gate268inter2, gate268inter3, gate268inter4, gate268inter5, gate268inter6, gate268inter7, gate268inter8, gate268inter9, gate268inter10, gate268inter11, gate268inter12, gate193inter0, gate193inter1, gate193inter2, gate193inter3, gate193inter4, gate193inter5, gate193inter6, gate193inter7, gate193inter8, gate193inter9, gate193inter10, gate193inter11, gate193inter12, gate68inter0, gate68inter1, gate68inter2, gate68inter3, gate68inter4, gate68inter5, gate68inter6, gate68inter7, gate68inter8, gate68inter9, gate68inter10, gate68inter11, gate68inter12, gate442inter0, gate442inter1, gate442inter2, gate442inter3, gate442inter4, gate442inter5, gate442inter6, gate442inter7, gate442inter8, gate442inter9, gate442inter10, gate442inter11, gate442inter12, gate177inter0, gate177inter1, gate177inter2, gate177inter3, gate177inter4, gate177inter5, gate177inter6, gate177inter7, gate177inter8, gate177inter9, gate177inter10, gate177inter11, gate177inter12, gate91inter0, gate91inter1, gate91inter2, gate91inter3, gate91inter4, gate91inter5, gate91inter6, gate91inter7, gate91inter8, gate91inter9, gate91inter10, gate91inter11, gate91inter12, gate513inter0, gate513inter1, gate513inter2, gate513inter3, gate513inter4, gate513inter5, gate513inter6, gate513inter7, gate513inter8, gate513inter9, gate513inter10, gate513inter11, gate513inter12, gate488inter0, gate488inter1, gate488inter2, gate488inter3, gate488inter4, gate488inter5, gate488inter6, gate488inter7, gate488inter8, gate488inter9, gate488inter10, gate488inter11, gate488inter12, gate184inter0, gate184inter1, gate184inter2, gate184inter3, gate184inter4, gate184inter5, gate184inter6, gate184inter7, gate184inter8, gate184inter9, gate184inter10, gate184inter11, gate184inter12, gate465inter0, gate465inter1, gate465inter2, gate465inter3, gate465inter4, gate465inter5, gate465inter6, gate465inter7, gate465inter8, gate465inter9, gate465inter10, gate465inter11, gate465inter12, gate274inter0, gate274inter1, gate274inter2, gate274inter3, gate274inter4, gate274inter5, gate274inter6, gate274inter7, gate274inter8, gate274inter9, gate274inter10, gate274inter11, gate274inter12, gate244inter0, gate244inter1, gate244inter2, gate244inter3, gate244inter4, gate244inter5, gate244inter6, gate244inter7, gate244inter8, gate244inter9, gate244inter10, gate244inter11, gate244inter12, gate257inter0, gate257inter1, gate257inter2, gate257inter3, gate257inter4, gate257inter5, gate257inter6, gate257inter7, gate257inter8, gate257inter9, gate257inter10, gate257inter11, gate257inter12, gate209inter0, gate209inter1, gate209inter2, gate209inter3, gate209inter4, gate209inter5, gate209inter6, gate209inter7, gate209inter8, gate209inter9, gate209inter10, gate209inter11, gate209inter12, gate13inter0, gate13inter1, gate13inter2, gate13inter3, gate13inter4, gate13inter5, gate13inter6, gate13inter7, gate13inter8, gate13inter9, gate13inter10, gate13inter11, gate13inter12, gate253inter0, gate253inter1, gate253inter2, gate253inter3, gate253inter4, gate253inter5, gate253inter6, gate253inter7, gate253inter8, gate253inter9, gate253inter10, gate253inter11, gate253inter12, gate50inter0, gate50inter1, gate50inter2, gate50inter3, gate50inter4, gate50inter5, gate50inter6, gate50inter7, gate50inter8, gate50inter9, gate50inter10, gate50inter11, gate50inter12, gate477inter0, gate477inter1, gate477inter2, gate477inter3, gate477inter4, gate477inter5, gate477inter6, gate477inter7, gate477inter8, gate477inter9, gate477inter10, gate477inter11, gate477inter12, gate225inter0, gate225inter1, gate225inter2, gate225inter3, gate225inter4, gate225inter5, gate225inter6, gate225inter7, gate225inter8, gate225inter9, gate225inter10, gate225inter11, gate225inter12, gate431inter0, gate431inter1, gate431inter2, gate431inter3, gate431inter4, gate431inter5, gate431inter6, gate431inter7, gate431inter8, gate431inter9, gate431inter10, gate431inter11, gate431inter12, gate24inter0, gate24inter1, gate24inter2, gate24inter3, gate24inter4, gate24inter5, gate24inter6, gate24inter7, gate24inter8, gate24inter9, gate24inter10, gate24inter11, gate24inter12, gate171inter0, gate171inter1, gate171inter2, gate171inter3, gate171inter4, gate171inter5, gate171inter6, gate171inter7, gate171inter8, gate171inter9, gate171inter10, gate171inter11, gate171inter12, gate92inter0, gate92inter1, gate92inter2, gate92inter3, gate92inter4, gate92inter5, gate92inter6, gate92inter7, gate92inter8, gate92inter9, gate92inter10, gate92inter11, gate92inter12, gate227inter0, gate227inter1, gate227inter2, gate227inter3, gate227inter4, gate227inter5, gate227inter6, gate227inter7, gate227inter8, gate227inter9, gate227inter10, gate227inter11, gate227inter12, gate449inter0, gate449inter1, gate449inter2, gate449inter3, gate449inter4, gate449inter5, gate449inter6, gate449inter7, gate449inter8, gate449inter9, gate449inter10, gate449inter11, gate449inter12, gate10inter0, gate10inter1, gate10inter2, gate10inter3, gate10inter4, gate10inter5, gate10inter6, gate10inter7, gate10inter8, gate10inter9, gate10inter10, gate10inter11, gate10inter12, gate502inter0, gate502inter1, gate502inter2, gate502inter3, gate502inter4, gate502inter5, gate502inter6, gate502inter7, gate502inter8, gate502inter9, gate502inter10, gate502inter11, gate502inter12, gate76inter0, gate76inter1, gate76inter2, gate76inter3, gate76inter4, gate76inter5, gate76inter6, gate76inter7, gate76inter8, gate76inter9, gate76inter10, gate76inter11, gate76inter12, gate46inter0, gate46inter1, gate46inter2, gate46inter3, gate46inter4, gate46inter5, gate46inter6, gate46inter7, gate46inter8, gate46inter9, gate46inter10, gate46inter11, gate46inter12, gate160inter0, gate160inter1, gate160inter2, gate160inter3, gate160inter4, gate160inter5, gate160inter6, gate160inter7, gate160inter8, gate160inter9, gate160inter10, gate160inter11, gate160inter12, gate109inter0, gate109inter1, gate109inter2, gate109inter3, gate109inter4, gate109inter5, gate109inter6, gate109inter7, gate109inter8, gate109inter9, gate109inter10, gate109inter11, gate109inter12, gate387inter0, gate387inter1, gate387inter2, gate387inter3, gate387inter4, gate387inter5, gate387inter6, gate387inter7, gate387inter8, gate387inter9, gate387inter10, gate387inter11, gate387inter12, gate239inter0, gate239inter1, gate239inter2, gate239inter3, gate239inter4, gate239inter5, gate239inter6, gate239inter7, gate239inter8, gate239inter9, gate239inter10, gate239inter11, gate239inter12, gate185inter0, gate185inter1, gate185inter2, gate185inter3, gate185inter4, gate185inter5, gate185inter6, gate185inter7, gate185inter8, gate185inter9, gate185inter10, gate185inter11, gate185inter12, gate296inter0, gate296inter1, gate296inter2, gate296inter3, gate296inter4, gate296inter5, gate296inter6, gate296inter7, gate296inter8, gate296inter9, gate296inter10, gate296inter11, gate296inter12, gate461inter0, gate461inter1, gate461inter2, gate461inter3, gate461inter4, gate461inter5, gate461inter6, gate461inter7, gate461inter8, gate461inter9, gate461inter10, gate461inter11, gate461inter12, gate192inter0, gate192inter1, gate192inter2, gate192inter3, gate192inter4, gate192inter5, gate192inter6, gate192inter7, gate192inter8, gate192inter9, gate192inter10, gate192inter11, gate192inter12, gate14inter0, gate14inter1, gate14inter2, gate14inter3, gate14inter4, gate14inter5, gate14inter6, gate14inter7, gate14inter8, gate14inter9, gate14inter10, gate14inter11, gate14inter12, gate151inter0, gate151inter1, gate151inter2, gate151inter3, gate151inter4, gate151inter5, gate151inter6, gate151inter7, gate151inter8, gate151inter9, gate151inter10, gate151inter11, gate151inter12, gate183inter0, gate183inter1, gate183inter2, gate183inter3, gate183inter4, gate183inter5, gate183inter6, gate183inter7, gate183inter8, gate183inter9, gate183inter10, gate183inter11, gate183inter12, gate173inter0, gate173inter1, gate173inter2, gate173inter3, gate173inter4, gate173inter5, gate173inter6, gate173inter7, gate173inter8, gate173inter9, gate173inter10, gate173inter11, gate173inter12, gate405inter0, gate405inter1, gate405inter2, gate405inter3, gate405inter4, gate405inter5, gate405inter6, gate405inter7, gate405inter8, gate405inter9, gate405inter10, gate405inter11, gate405inter12, gate432inter0, gate432inter1, gate432inter2, gate432inter3, gate432inter4, gate432inter5, gate432inter6, gate432inter7, gate432inter8, gate432inter9, gate432inter10, gate432inter11, gate432inter12, gate129inter0, gate129inter1, gate129inter2, gate129inter3, gate129inter4, gate129inter5, gate129inter6, gate129inter7, gate129inter8, gate129inter9, gate129inter10, gate129inter11, gate129inter12, gate391inter0, gate391inter1, gate391inter2, gate391inter3, gate391inter4, gate391inter5, gate391inter6, gate391inter7, gate391inter8, gate391inter9, gate391inter10, gate391inter11, gate391inter12, gate202inter0, gate202inter1, gate202inter2, gate202inter3, gate202inter4, gate202inter5, gate202inter6, gate202inter7, gate202inter8, gate202inter9, gate202inter10, gate202inter11, gate202inter12, gate270inter0, gate270inter1, gate270inter2, gate270inter3, gate270inter4, gate270inter5, gate270inter6, gate270inter7, gate270inter8, gate270inter9, gate270inter10, gate270inter11, gate270inter12, gate143inter0, gate143inter1, gate143inter2, gate143inter3, gate143inter4, gate143inter5, gate143inter6, gate143inter7, gate143inter8, gate143inter9, gate143inter10, gate143inter11, gate143inter12, gate108inter0, gate108inter1, gate108inter2, gate108inter3, gate108inter4, gate108inter5, gate108inter6, gate108inter7, gate108inter8, gate108inter9, gate108inter10, gate108inter11, gate108inter12, gate462inter0, gate462inter1, gate462inter2, gate462inter3, gate462inter4, gate462inter5, gate462inter6, gate462inter7, gate462inter8, gate462inter9, gate462inter10, gate462inter11, gate462inter12, gate237inter0, gate237inter1, gate237inter2, gate237inter3, gate237inter4, gate237inter5, gate237inter6, gate237inter7, gate237inter8, gate237inter9, gate237inter10, gate237inter11, gate237inter12, gate293inter0, gate293inter1, gate293inter2, gate293inter3, gate293inter4, gate293inter5, gate293inter6, gate293inter7, gate293inter8, gate293inter9, gate293inter10, gate293inter11, gate293inter12, gate263inter0, gate263inter1, gate263inter2, gate263inter3, gate263inter4, gate263inter5, gate263inter6, gate263inter7, gate263inter8, gate263inter9, gate263inter10, gate263inter11, gate263inter12, gate258inter0, gate258inter1, gate258inter2, gate258inter3, gate258inter4, gate258inter5, gate258inter6, gate258inter7, gate258inter8, gate258inter9, gate258inter10, gate258inter11, gate258inter12, gate414inter0, gate414inter1, gate414inter2, gate414inter3, gate414inter4, gate414inter5, gate414inter6, gate414inter7, gate414inter8, gate414inter9, gate414inter10, gate414inter11, gate414inter12, gate120inter0, gate120inter1, gate120inter2, gate120inter3, gate120inter4, gate120inter5, gate120inter6, gate120inter7, gate120inter8, gate120inter9, gate120inter10, gate120inter11, gate120inter12, gate284inter0, gate284inter1, gate284inter2, gate284inter3, gate284inter4, gate284inter5, gate284inter6, gate284inter7, gate284inter8, gate284inter9, gate284inter10, gate284inter11, gate284inter12, gate285inter0, gate285inter1, gate285inter2, gate285inter3, gate285inter4, gate285inter5, gate285inter6, gate285inter7, gate285inter8, gate285inter9, gate285inter10, gate285inter11, gate285inter12, gate215inter0, gate215inter1, gate215inter2, gate215inter3, gate215inter4, gate215inter5, gate215inter6, gate215inter7, gate215inter8, gate215inter9, gate215inter10, gate215inter11, gate215inter12, gate280inter0, gate280inter1, gate280inter2, gate280inter3, gate280inter4, gate280inter5, gate280inter6, gate280inter7, gate280inter8, gate280inter9, gate280inter10, gate280inter11, gate280inter12, gate433inter0, gate433inter1, gate433inter2, gate433inter3, gate433inter4, gate433inter5, gate433inter6, gate433inter7, gate433inter8, gate433inter9, gate433inter10, gate433inter11, gate433inter12, gate187inter0, gate187inter1, gate187inter2, gate187inter3, gate187inter4, gate187inter5, gate187inter6, gate187inter7, gate187inter8, gate187inter9, gate187inter10, gate187inter11, gate187inter12, gate458inter0, gate458inter1, gate458inter2, gate458inter3, gate458inter4, gate458inter5, gate458inter6, gate458inter7, gate458inter8, gate458inter9, gate458inter10, gate458inter11, gate458inter12, gate262inter0, gate262inter1, gate262inter2, gate262inter3, gate262inter4, gate262inter5, gate262inter6, gate262inter7, gate262inter8, gate262inter9, gate262inter10, gate262inter11, gate262inter12, gate105inter0, gate105inter1, gate105inter2, gate105inter3, gate105inter4, gate105inter5, gate105inter6, gate105inter7, gate105inter8, gate105inter9, gate105inter10, gate105inter11, gate105inter12, gate179inter0, gate179inter1, gate179inter2, gate179inter3, gate179inter4, gate179inter5, gate179inter6, gate179inter7, gate179inter8, gate179inter9, gate179inter10, gate179inter11, gate179inter12, gate246inter0, gate246inter1, gate246inter2, gate246inter3, gate246inter4, gate246inter5, gate246inter6, gate246inter7, gate246inter8, gate246inter9, gate246inter10, gate246inter11, gate246inter12, gate62inter0, gate62inter1, gate62inter2, gate62inter3, gate62inter4, gate62inter5, gate62inter6, gate62inter7, gate62inter8, gate62inter9, gate62inter10, gate62inter11, gate62inter12, gate21inter0, gate21inter1, gate21inter2, gate21inter3, gate21inter4, gate21inter5, gate21inter6, gate21inter7, gate21inter8, gate21inter9, gate21inter10, gate21inter11, gate21inter12, gate240inter0, gate240inter1, gate240inter2, gate240inter3, gate240inter4, gate240inter5, gate240inter6, gate240inter7, gate240inter8, gate240inter9, gate240inter10, gate240inter11, gate240inter12, gate485inter0, gate485inter1, gate485inter2, gate485inter3, gate485inter4, gate485inter5, gate485inter6, gate485inter7, gate485inter8, gate485inter9, gate485inter10, gate485inter11, gate485inter12, gate142inter0, gate142inter1, gate142inter2, gate142inter3, gate142inter4, gate142inter5, gate142inter6, gate142inter7, gate142inter8, gate142inter9, gate142inter10, gate142inter11, gate142inter12, gate250inter0, gate250inter1, gate250inter2, gate250inter3, gate250inter4, gate250inter5, gate250inter6, gate250inter7, gate250inter8, gate250inter9, gate250inter10, gate250inter11, gate250inter12, gate141inter0, gate141inter1, gate141inter2, gate141inter3, gate141inter4, gate141inter5, gate141inter6, gate141inter7, gate141inter8, gate141inter9, gate141inter10, gate141inter11, gate141inter12, gate398inter0, gate398inter1, gate398inter2, gate398inter3, gate398inter4, gate398inter5, gate398inter6, gate398inter7, gate398inter8, gate398inter9, gate398inter10, gate398inter11, gate398inter12, gate163inter0, gate163inter1, gate163inter2, gate163inter3, gate163inter4, gate163inter5, gate163inter6, gate163inter7, gate163inter8, gate163inter9, gate163inter10, gate163inter11, gate163inter12, gate63inter0, gate63inter1, gate63inter2, gate63inter3, gate63inter4, gate63inter5, gate63inter6, gate63inter7, gate63inter8, gate63inter9, gate63inter10, gate63inter11, gate63inter12, gate402inter0, gate402inter1, gate402inter2, gate402inter3, gate402inter4, gate402inter5, gate402inter6, gate402inter7, gate402inter8, gate402inter9, gate402inter10, gate402inter11, gate402inter12, gate482inter0, gate482inter1, gate482inter2, gate482inter3, gate482inter4, gate482inter5, gate482inter6, gate482inter7, gate482inter8, gate482inter9, gate482inter10, gate482inter11, gate482inter12, gate157inter0, gate157inter1, gate157inter2, gate157inter3, gate157inter4, gate157inter5, gate157inter6, gate157inter7, gate157inter8, gate157inter9, gate157inter10, gate157inter11, gate157inter12, gate74inter0, gate74inter1, gate74inter2, gate74inter3, gate74inter4, gate74inter5, gate74inter6, gate74inter7, gate74inter8, gate74inter9, gate74inter10, gate74inter11, gate74inter12, gate101inter0, gate101inter1, gate101inter2, gate101inter3, gate101inter4, gate101inter5, gate101inter6, gate101inter7, gate101inter8, gate101inter9, gate101inter10, gate101inter11, gate101inter12, gate71inter0, gate71inter1, gate71inter2, gate71inter3, gate71inter4, gate71inter5, gate71inter6, gate71inter7, gate71inter8, gate71inter9, gate71inter10, gate71inter11, gate71inter12, gate52inter0, gate52inter1, gate52inter2, gate52inter3, gate52inter4, gate52inter5, gate52inter6, gate52inter7, gate52inter8, gate52inter9, gate52inter10, gate52inter11, gate52inter12, gate18inter0, gate18inter1, gate18inter2, gate18inter3, gate18inter4, gate18inter5, gate18inter6, gate18inter7, gate18inter8, gate18inter9, gate18inter10, gate18inter11, gate18inter12, gate288inter0, gate288inter1, gate288inter2, gate288inter3, gate288inter4, gate288inter5, gate288inter6, gate288inter7, gate288inter8, gate288inter9, gate288inter10, gate288inter11, gate288inter12;



and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );
nand2 gate9( .a(G1), .b(G2), .O(G266) );

  xor2  gate1877(.a(G4), .b(G3), .O(gate10inter0));
  nand2 gate1878(.a(gate10inter0), .b(s_190), .O(gate10inter1));
  and2  gate1879(.a(G4), .b(G3), .O(gate10inter2));
  inv1  gate1880(.a(s_190), .O(gate10inter3));
  inv1  gate1881(.a(s_191), .O(gate10inter4));
  nand2 gate1882(.a(gate10inter4), .b(gate10inter3), .O(gate10inter5));
  nor2  gate1883(.a(gate10inter5), .b(gate10inter2), .O(gate10inter6));
  inv1  gate1884(.a(G3), .O(gate10inter7));
  inv1  gate1885(.a(G4), .O(gate10inter8));
  nand2 gate1886(.a(gate10inter8), .b(gate10inter7), .O(gate10inter9));
  nand2 gate1887(.a(s_191), .b(gate10inter3), .O(gate10inter10));
  nor2  gate1888(.a(gate10inter10), .b(gate10inter9), .O(gate10inter11));
  nor2  gate1889(.a(gate10inter11), .b(gate10inter6), .O(gate10inter12));
  nand2 gate1890(.a(gate10inter12), .b(gate10inter1), .O(G269));

  xor2  gate1457(.a(G6), .b(G5), .O(gate11inter0));
  nand2 gate1458(.a(gate11inter0), .b(s_130), .O(gate11inter1));
  and2  gate1459(.a(G6), .b(G5), .O(gate11inter2));
  inv1  gate1460(.a(s_130), .O(gate11inter3));
  inv1  gate1461(.a(s_131), .O(gate11inter4));
  nand2 gate1462(.a(gate11inter4), .b(gate11inter3), .O(gate11inter5));
  nor2  gate1463(.a(gate11inter5), .b(gate11inter2), .O(gate11inter6));
  inv1  gate1464(.a(G5), .O(gate11inter7));
  inv1  gate1465(.a(G6), .O(gate11inter8));
  nand2 gate1466(.a(gate11inter8), .b(gate11inter7), .O(gate11inter9));
  nand2 gate1467(.a(s_131), .b(gate11inter3), .O(gate11inter10));
  nor2  gate1468(.a(gate11inter10), .b(gate11inter9), .O(gate11inter11));
  nor2  gate1469(.a(gate11inter11), .b(gate11inter6), .O(gate11inter12));
  nand2 gate1470(.a(gate11inter12), .b(gate11inter1), .O(G272));
nand2 gate12( .a(G7), .b(G8), .O(G275) );

  xor2  gate1723(.a(G10), .b(G9), .O(gate13inter0));
  nand2 gate1724(.a(gate13inter0), .b(s_168), .O(gate13inter1));
  and2  gate1725(.a(G10), .b(G9), .O(gate13inter2));
  inv1  gate1726(.a(s_168), .O(gate13inter3));
  inv1  gate1727(.a(s_169), .O(gate13inter4));
  nand2 gate1728(.a(gate13inter4), .b(gate13inter3), .O(gate13inter5));
  nor2  gate1729(.a(gate13inter5), .b(gate13inter2), .O(gate13inter6));
  inv1  gate1730(.a(G9), .O(gate13inter7));
  inv1  gate1731(.a(G10), .O(gate13inter8));
  nand2 gate1732(.a(gate13inter8), .b(gate13inter7), .O(gate13inter9));
  nand2 gate1733(.a(s_169), .b(gate13inter3), .O(gate13inter10));
  nor2  gate1734(.a(gate13inter10), .b(gate13inter9), .O(gate13inter11));
  nor2  gate1735(.a(gate13inter11), .b(gate13inter6), .O(gate13inter12));
  nand2 gate1736(.a(gate13inter12), .b(gate13inter1), .O(G278));

  xor2  gate2045(.a(G12), .b(G11), .O(gate14inter0));
  nand2 gate2046(.a(gate14inter0), .b(s_214), .O(gate14inter1));
  and2  gate2047(.a(G12), .b(G11), .O(gate14inter2));
  inv1  gate2048(.a(s_214), .O(gate14inter3));
  inv1  gate2049(.a(s_215), .O(gate14inter4));
  nand2 gate2050(.a(gate14inter4), .b(gate14inter3), .O(gate14inter5));
  nor2  gate2051(.a(gate14inter5), .b(gate14inter2), .O(gate14inter6));
  inv1  gate2052(.a(G11), .O(gate14inter7));
  inv1  gate2053(.a(G12), .O(gate14inter8));
  nand2 gate2054(.a(gate14inter8), .b(gate14inter7), .O(gate14inter9));
  nand2 gate2055(.a(s_215), .b(gate14inter3), .O(gate14inter10));
  nor2  gate2056(.a(gate14inter10), .b(gate14inter9), .O(gate14inter11));
  nor2  gate2057(.a(gate14inter11), .b(gate14inter6), .O(gate14inter12));
  nand2 gate2058(.a(gate14inter12), .b(gate14inter1), .O(G281));

  xor2  gate575(.a(G14), .b(G13), .O(gate15inter0));
  nand2 gate576(.a(gate15inter0), .b(s_4), .O(gate15inter1));
  and2  gate577(.a(G14), .b(G13), .O(gate15inter2));
  inv1  gate578(.a(s_4), .O(gate15inter3));
  inv1  gate579(.a(s_5), .O(gate15inter4));
  nand2 gate580(.a(gate15inter4), .b(gate15inter3), .O(gate15inter5));
  nor2  gate581(.a(gate15inter5), .b(gate15inter2), .O(gate15inter6));
  inv1  gate582(.a(G13), .O(gate15inter7));
  inv1  gate583(.a(G14), .O(gate15inter8));
  nand2 gate584(.a(gate15inter8), .b(gate15inter7), .O(gate15inter9));
  nand2 gate585(.a(s_5), .b(gate15inter3), .O(gate15inter10));
  nor2  gate586(.a(gate15inter10), .b(gate15inter9), .O(gate15inter11));
  nor2  gate587(.a(gate15inter11), .b(gate15inter6), .O(gate15inter12));
  nand2 gate588(.a(gate15inter12), .b(gate15inter1), .O(G284));
nand2 gate16( .a(G15), .b(G16), .O(G287) );

  xor2  gate1177(.a(G18), .b(G17), .O(gate17inter0));
  nand2 gate1178(.a(gate17inter0), .b(s_90), .O(gate17inter1));
  and2  gate1179(.a(G18), .b(G17), .O(gate17inter2));
  inv1  gate1180(.a(s_90), .O(gate17inter3));
  inv1  gate1181(.a(s_91), .O(gate17inter4));
  nand2 gate1182(.a(gate17inter4), .b(gate17inter3), .O(gate17inter5));
  nor2  gate1183(.a(gate17inter5), .b(gate17inter2), .O(gate17inter6));
  inv1  gate1184(.a(G17), .O(gate17inter7));
  inv1  gate1185(.a(G18), .O(gate17inter8));
  nand2 gate1186(.a(gate17inter8), .b(gate17inter7), .O(gate17inter9));
  nand2 gate1187(.a(s_91), .b(gate17inter3), .O(gate17inter10));
  nor2  gate1188(.a(gate17inter10), .b(gate17inter9), .O(gate17inter11));
  nor2  gate1189(.a(gate17inter11), .b(gate17inter6), .O(gate17inter12));
  nand2 gate1190(.a(gate17inter12), .b(gate17inter1), .O(G290));

  xor2  gate2703(.a(G20), .b(G19), .O(gate18inter0));
  nand2 gate2704(.a(gate18inter0), .b(s_308), .O(gate18inter1));
  and2  gate2705(.a(G20), .b(G19), .O(gate18inter2));
  inv1  gate2706(.a(s_308), .O(gate18inter3));
  inv1  gate2707(.a(s_309), .O(gate18inter4));
  nand2 gate2708(.a(gate18inter4), .b(gate18inter3), .O(gate18inter5));
  nor2  gate2709(.a(gate18inter5), .b(gate18inter2), .O(gate18inter6));
  inv1  gate2710(.a(G19), .O(gate18inter7));
  inv1  gate2711(.a(G20), .O(gate18inter8));
  nand2 gate2712(.a(gate18inter8), .b(gate18inter7), .O(gate18inter9));
  nand2 gate2713(.a(s_309), .b(gate18inter3), .O(gate18inter10));
  nor2  gate2714(.a(gate18inter10), .b(gate18inter9), .O(gate18inter11));
  nor2  gate2715(.a(gate18inter11), .b(gate18inter6), .O(gate18inter12));
  nand2 gate2716(.a(gate18inter12), .b(gate18inter1), .O(G293));
nand2 gate19( .a(G21), .b(G22), .O(G296) );
nand2 gate20( .a(G23), .b(G24), .O(G299) );

  xor2  gate2479(.a(G26), .b(G25), .O(gate21inter0));
  nand2 gate2480(.a(gate21inter0), .b(s_276), .O(gate21inter1));
  and2  gate2481(.a(G26), .b(G25), .O(gate21inter2));
  inv1  gate2482(.a(s_276), .O(gate21inter3));
  inv1  gate2483(.a(s_277), .O(gate21inter4));
  nand2 gate2484(.a(gate21inter4), .b(gate21inter3), .O(gate21inter5));
  nor2  gate2485(.a(gate21inter5), .b(gate21inter2), .O(gate21inter6));
  inv1  gate2486(.a(G25), .O(gate21inter7));
  inv1  gate2487(.a(G26), .O(gate21inter8));
  nand2 gate2488(.a(gate21inter8), .b(gate21inter7), .O(gate21inter9));
  nand2 gate2489(.a(s_277), .b(gate21inter3), .O(gate21inter10));
  nor2  gate2490(.a(gate21inter10), .b(gate21inter9), .O(gate21inter11));
  nor2  gate2491(.a(gate21inter11), .b(gate21inter6), .O(gate21inter12));
  nand2 gate2492(.a(gate21inter12), .b(gate21inter1), .O(G302));
nand2 gate22( .a(G27), .b(G28), .O(G305) );
nand2 gate23( .a(G29), .b(G30), .O(G308) );

  xor2  gate1807(.a(G32), .b(G31), .O(gate24inter0));
  nand2 gate1808(.a(gate24inter0), .b(s_180), .O(gate24inter1));
  and2  gate1809(.a(G32), .b(G31), .O(gate24inter2));
  inv1  gate1810(.a(s_180), .O(gate24inter3));
  inv1  gate1811(.a(s_181), .O(gate24inter4));
  nand2 gate1812(.a(gate24inter4), .b(gate24inter3), .O(gate24inter5));
  nor2  gate1813(.a(gate24inter5), .b(gate24inter2), .O(gate24inter6));
  inv1  gate1814(.a(G31), .O(gate24inter7));
  inv1  gate1815(.a(G32), .O(gate24inter8));
  nand2 gate1816(.a(gate24inter8), .b(gate24inter7), .O(gate24inter9));
  nand2 gate1817(.a(s_181), .b(gate24inter3), .O(gate24inter10));
  nor2  gate1818(.a(gate24inter10), .b(gate24inter9), .O(gate24inter11));
  nor2  gate1819(.a(gate24inter11), .b(gate24inter6), .O(gate24inter12));
  nand2 gate1820(.a(gate24inter12), .b(gate24inter1), .O(G311));

  xor2  gate673(.a(G5), .b(G1), .O(gate25inter0));
  nand2 gate674(.a(gate25inter0), .b(s_18), .O(gate25inter1));
  and2  gate675(.a(G5), .b(G1), .O(gate25inter2));
  inv1  gate676(.a(s_18), .O(gate25inter3));
  inv1  gate677(.a(s_19), .O(gate25inter4));
  nand2 gate678(.a(gate25inter4), .b(gate25inter3), .O(gate25inter5));
  nor2  gate679(.a(gate25inter5), .b(gate25inter2), .O(gate25inter6));
  inv1  gate680(.a(G1), .O(gate25inter7));
  inv1  gate681(.a(G5), .O(gate25inter8));
  nand2 gate682(.a(gate25inter8), .b(gate25inter7), .O(gate25inter9));
  nand2 gate683(.a(s_19), .b(gate25inter3), .O(gate25inter10));
  nor2  gate684(.a(gate25inter10), .b(gate25inter9), .O(gate25inter11));
  nor2  gate685(.a(gate25inter11), .b(gate25inter6), .O(gate25inter12));
  nand2 gate686(.a(gate25inter12), .b(gate25inter1), .O(G314));
nand2 gate26( .a(G9), .b(G13), .O(G317) );
nand2 gate27( .a(G2), .b(G6), .O(G320) );
nand2 gate28( .a(G10), .b(G14), .O(G323) );
nand2 gate29( .a(G3), .b(G7), .O(G326) );
nand2 gate30( .a(G11), .b(G15), .O(G329) );
nand2 gate31( .a(G4), .b(G8), .O(G332) );
nand2 gate32( .a(G12), .b(G16), .O(G335) );
nand2 gate33( .a(G17), .b(G21), .O(G338) );
nand2 gate34( .a(G25), .b(G29), .O(G341) );
nand2 gate35( .a(G18), .b(G22), .O(G344) );

  xor2  gate813(.a(G30), .b(G26), .O(gate36inter0));
  nand2 gate814(.a(gate36inter0), .b(s_38), .O(gate36inter1));
  and2  gate815(.a(G30), .b(G26), .O(gate36inter2));
  inv1  gate816(.a(s_38), .O(gate36inter3));
  inv1  gate817(.a(s_39), .O(gate36inter4));
  nand2 gate818(.a(gate36inter4), .b(gate36inter3), .O(gate36inter5));
  nor2  gate819(.a(gate36inter5), .b(gate36inter2), .O(gate36inter6));
  inv1  gate820(.a(G26), .O(gate36inter7));
  inv1  gate821(.a(G30), .O(gate36inter8));
  nand2 gate822(.a(gate36inter8), .b(gate36inter7), .O(gate36inter9));
  nand2 gate823(.a(s_39), .b(gate36inter3), .O(gate36inter10));
  nor2  gate824(.a(gate36inter10), .b(gate36inter9), .O(gate36inter11));
  nor2  gate825(.a(gate36inter11), .b(gate36inter6), .O(gate36inter12));
  nand2 gate826(.a(gate36inter12), .b(gate36inter1), .O(G347));
nand2 gate37( .a(G19), .b(G23), .O(G350) );
nand2 gate38( .a(G27), .b(G31), .O(G353) );
nand2 gate39( .a(G20), .b(G24), .O(G356) );
nand2 gate40( .a(G28), .b(G32), .O(G359) );
nand2 gate41( .a(G1), .b(G266), .O(G362) );
nand2 gate42( .a(G2), .b(G266), .O(G363) );
nand2 gate43( .a(G3), .b(G269), .O(G364) );
nand2 gate44( .a(G4), .b(G269), .O(G365) );

  xor2  gate785(.a(G272), .b(G5), .O(gate45inter0));
  nand2 gate786(.a(gate45inter0), .b(s_34), .O(gate45inter1));
  and2  gate787(.a(G272), .b(G5), .O(gate45inter2));
  inv1  gate788(.a(s_34), .O(gate45inter3));
  inv1  gate789(.a(s_35), .O(gate45inter4));
  nand2 gate790(.a(gate45inter4), .b(gate45inter3), .O(gate45inter5));
  nor2  gate791(.a(gate45inter5), .b(gate45inter2), .O(gate45inter6));
  inv1  gate792(.a(G5), .O(gate45inter7));
  inv1  gate793(.a(G272), .O(gate45inter8));
  nand2 gate794(.a(gate45inter8), .b(gate45inter7), .O(gate45inter9));
  nand2 gate795(.a(s_35), .b(gate45inter3), .O(gate45inter10));
  nor2  gate796(.a(gate45inter10), .b(gate45inter9), .O(gate45inter11));
  nor2  gate797(.a(gate45inter11), .b(gate45inter6), .O(gate45inter12));
  nand2 gate798(.a(gate45inter12), .b(gate45inter1), .O(G366));

  xor2  gate1919(.a(G272), .b(G6), .O(gate46inter0));
  nand2 gate1920(.a(gate46inter0), .b(s_196), .O(gate46inter1));
  and2  gate1921(.a(G272), .b(G6), .O(gate46inter2));
  inv1  gate1922(.a(s_196), .O(gate46inter3));
  inv1  gate1923(.a(s_197), .O(gate46inter4));
  nand2 gate1924(.a(gate46inter4), .b(gate46inter3), .O(gate46inter5));
  nor2  gate1925(.a(gate46inter5), .b(gate46inter2), .O(gate46inter6));
  inv1  gate1926(.a(G6), .O(gate46inter7));
  inv1  gate1927(.a(G272), .O(gate46inter8));
  nand2 gate1928(.a(gate46inter8), .b(gate46inter7), .O(gate46inter9));
  nand2 gate1929(.a(s_197), .b(gate46inter3), .O(gate46inter10));
  nor2  gate1930(.a(gate46inter10), .b(gate46inter9), .O(gate46inter11));
  nor2  gate1931(.a(gate46inter11), .b(gate46inter6), .O(gate46inter12));
  nand2 gate1932(.a(gate46inter12), .b(gate46inter1), .O(G367));
nand2 gate47( .a(G7), .b(G275), .O(G368) );
nand2 gate48( .a(G8), .b(G275), .O(G369) );

  xor2  gate771(.a(G278), .b(G9), .O(gate49inter0));
  nand2 gate772(.a(gate49inter0), .b(s_32), .O(gate49inter1));
  and2  gate773(.a(G278), .b(G9), .O(gate49inter2));
  inv1  gate774(.a(s_32), .O(gate49inter3));
  inv1  gate775(.a(s_33), .O(gate49inter4));
  nand2 gate776(.a(gate49inter4), .b(gate49inter3), .O(gate49inter5));
  nor2  gate777(.a(gate49inter5), .b(gate49inter2), .O(gate49inter6));
  inv1  gate778(.a(G9), .O(gate49inter7));
  inv1  gate779(.a(G278), .O(gate49inter8));
  nand2 gate780(.a(gate49inter8), .b(gate49inter7), .O(gate49inter9));
  nand2 gate781(.a(s_33), .b(gate49inter3), .O(gate49inter10));
  nor2  gate782(.a(gate49inter10), .b(gate49inter9), .O(gate49inter11));
  nor2  gate783(.a(gate49inter11), .b(gate49inter6), .O(gate49inter12));
  nand2 gate784(.a(gate49inter12), .b(gate49inter1), .O(G370));

  xor2  gate1751(.a(G278), .b(G10), .O(gate50inter0));
  nand2 gate1752(.a(gate50inter0), .b(s_172), .O(gate50inter1));
  and2  gate1753(.a(G278), .b(G10), .O(gate50inter2));
  inv1  gate1754(.a(s_172), .O(gate50inter3));
  inv1  gate1755(.a(s_173), .O(gate50inter4));
  nand2 gate1756(.a(gate50inter4), .b(gate50inter3), .O(gate50inter5));
  nor2  gate1757(.a(gate50inter5), .b(gate50inter2), .O(gate50inter6));
  inv1  gate1758(.a(G10), .O(gate50inter7));
  inv1  gate1759(.a(G278), .O(gate50inter8));
  nand2 gate1760(.a(gate50inter8), .b(gate50inter7), .O(gate50inter9));
  nand2 gate1761(.a(s_173), .b(gate50inter3), .O(gate50inter10));
  nor2  gate1762(.a(gate50inter10), .b(gate50inter9), .O(gate50inter11));
  nor2  gate1763(.a(gate50inter11), .b(gate50inter6), .O(gate50inter12));
  nand2 gate1764(.a(gate50inter12), .b(gate50inter1), .O(G371));
nand2 gate51( .a(G11), .b(G281), .O(G372) );

  xor2  gate2689(.a(G281), .b(G12), .O(gate52inter0));
  nand2 gate2690(.a(gate52inter0), .b(s_306), .O(gate52inter1));
  and2  gate2691(.a(G281), .b(G12), .O(gate52inter2));
  inv1  gate2692(.a(s_306), .O(gate52inter3));
  inv1  gate2693(.a(s_307), .O(gate52inter4));
  nand2 gate2694(.a(gate52inter4), .b(gate52inter3), .O(gate52inter5));
  nor2  gate2695(.a(gate52inter5), .b(gate52inter2), .O(gate52inter6));
  inv1  gate2696(.a(G12), .O(gate52inter7));
  inv1  gate2697(.a(G281), .O(gate52inter8));
  nand2 gate2698(.a(gate52inter8), .b(gate52inter7), .O(gate52inter9));
  nand2 gate2699(.a(s_307), .b(gate52inter3), .O(gate52inter10));
  nor2  gate2700(.a(gate52inter10), .b(gate52inter9), .O(gate52inter11));
  nor2  gate2701(.a(gate52inter11), .b(gate52inter6), .O(gate52inter12));
  nand2 gate2702(.a(gate52inter12), .b(gate52inter1), .O(G373));
nand2 gate53( .a(G13), .b(G284), .O(G374) );
nand2 gate54( .a(G14), .b(G284), .O(G375) );
nand2 gate55( .a(G15), .b(G287), .O(G376) );

  xor2  gate1261(.a(G287), .b(G16), .O(gate56inter0));
  nand2 gate1262(.a(gate56inter0), .b(s_102), .O(gate56inter1));
  and2  gate1263(.a(G287), .b(G16), .O(gate56inter2));
  inv1  gate1264(.a(s_102), .O(gate56inter3));
  inv1  gate1265(.a(s_103), .O(gate56inter4));
  nand2 gate1266(.a(gate56inter4), .b(gate56inter3), .O(gate56inter5));
  nor2  gate1267(.a(gate56inter5), .b(gate56inter2), .O(gate56inter6));
  inv1  gate1268(.a(G16), .O(gate56inter7));
  inv1  gate1269(.a(G287), .O(gate56inter8));
  nand2 gate1270(.a(gate56inter8), .b(gate56inter7), .O(gate56inter9));
  nand2 gate1271(.a(s_103), .b(gate56inter3), .O(gate56inter10));
  nor2  gate1272(.a(gate56inter10), .b(gate56inter9), .O(gate56inter11));
  nor2  gate1273(.a(gate56inter11), .b(gate56inter6), .O(gate56inter12));
  nand2 gate1274(.a(gate56inter12), .b(gate56inter1), .O(G377));
nand2 gate57( .a(G17), .b(G290), .O(G378) );
nand2 gate58( .a(G18), .b(G290), .O(G379) );
nand2 gate59( .a(G19), .b(G293), .O(G380) );
nand2 gate60( .a(G20), .b(G293), .O(G381) );

  xor2  gate1485(.a(G296), .b(G21), .O(gate61inter0));
  nand2 gate1486(.a(gate61inter0), .b(s_134), .O(gate61inter1));
  and2  gate1487(.a(G296), .b(G21), .O(gate61inter2));
  inv1  gate1488(.a(s_134), .O(gate61inter3));
  inv1  gate1489(.a(s_135), .O(gate61inter4));
  nand2 gate1490(.a(gate61inter4), .b(gate61inter3), .O(gate61inter5));
  nor2  gate1491(.a(gate61inter5), .b(gate61inter2), .O(gate61inter6));
  inv1  gate1492(.a(G21), .O(gate61inter7));
  inv1  gate1493(.a(G296), .O(gate61inter8));
  nand2 gate1494(.a(gate61inter8), .b(gate61inter7), .O(gate61inter9));
  nand2 gate1495(.a(s_135), .b(gate61inter3), .O(gate61inter10));
  nor2  gate1496(.a(gate61inter10), .b(gate61inter9), .O(gate61inter11));
  nor2  gate1497(.a(gate61inter11), .b(gate61inter6), .O(gate61inter12));
  nand2 gate1498(.a(gate61inter12), .b(gate61inter1), .O(G382));

  xor2  gate2465(.a(G296), .b(G22), .O(gate62inter0));
  nand2 gate2466(.a(gate62inter0), .b(s_274), .O(gate62inter1));
  and2  gate2467(.a(G296), .b(G22), .O(gate62inter2));
  inv1  gate2468(.a(s_274), .O(gate62inter3));
  inv1  gate2469(.a(s_275), .O(gate62inter4));
  nand2 gate2470(.a(gate62inter4), .b(gate62inter3), .O(gate62inter5));
  nor2  gate2471(.a(gate62inter5), .b(gate62inter2), .O(gate62inter6));
  inv1  gate2472(.a(G22), .O(gate62inter7));
  inv1  gate2473(.a(G296), .O(gate62inter8));
  nand2 gate2474(.a(gate62inter8), .b(gate62inter7), .O(gate62inter9));
  nand2 gate2475(.a(s_275), .b(gate62inter3), .O(gate62inter10));
  nor2  gate2476(.a(gate62inter10), .b(gate62inter9), .O(gate62inter11));
  nor2  gate2477(.a(gate62inter11), .b(gate62inter6), .O(gate62inter12));
  nand2 gate2478(.a(gate62inter12), .b(gate62inter1), .O(G383));

  xor2  gate2591(.a(G299), .b(G23), .O(gate63inter0));
  nand2 gate2592(.a(gate63inter0), .b(s_292), .O(gate63inter1));
  and2  gate2593(.a(G299), .b(G23), .O(gate63inter2));
  inv1  gate2594(.a(s_292), .O(gate63inter3));
  inv1  gate2595(.a(s_293), .O(gate63inter4));
  nand2 gate2596(.a(gate63inter4), .b(gate63inter3), .O(gate63inter5));
  nor2  gate2597(.a(gate63inter5), .b(gate63inter2), .O(gate63inter6));
  inv1  gate2598(.a(G23), .O(gate63inter7));
  inv1  gate2599(.a(G299), .O(gate63inter8));
  nand2 gate2600(.a(gate63inter8), .b(gate63inter7), .O(gate63inter9));
  nand2 gate2601(.a(s_293), .b(gate63inter3), .O(gate63inter10));
  nor2  gate2602(.a(gate63inter10), .b(gate63inter9), .O(gate63inter11));
  nor2  gate2603(.a(gate63inter11), .b(gate63inter6), .O(gate63inter12));
  nand2 gate2604(.a(gate63inter12), .b(gate63inter1), .O(G384));

  xor2  gate841(.a(G299), .b(G24), .O(gate64inter0));
  nand2 gate842(.a(gate64inter0), .b(s_42), .O(gate64inter1));
  and2  gate843(.a(G299), .b(G24), .O(gate64inter2));
  inv1  gate844(.a(s_42), .O(gate64inter3));
  inv1  gate845(.a(s_43), .O(gate64inter4));
  nand2 gate846(.a(gate64inter4), .b(gate64inter3), .O(gate64inter5));
  nor2  gate847(.a(gate64inter5), .b(gate64inter2), .O(gate64inter6));
  inv1  gate848(.a(G24), .O(gate64inter7));
  inv1  gate849(.a(G299), .O(gate64inter8));
  nand2 gate850(.a(gate64inter8), .b(gate64inter7), .O(gate64inter9));
  nand2 gate851(.a(s_43), .b(gate64inter3), .O(gate64inter10));
  nor2  gate852(.a(gate64inter10), .b(gate64inter9), .O(gate64inter11));
  nor2  gate853(.a(gate64inter11), .b(gate64inter6), .O(gate64inter12));
  nand2 gate854(.a(gate64inter12), .b(gate64inter1), .O(G385));
nand2 gate65( .a(G25), .b(G302), .O(G386) );
nand2 gate66( .a(G26), .b(G302), .O(G387) );
nand2 gate67( .a(G27), .b(G305), .O(G388) );

  xor2  gate1555(.a(G305), .b(G28), .O(gate68inter0));
  nand2 gate1556(.a(gate68inter0), .b(s_144), .O(gate68inter1));
  and2  gate1557(.a(G305), .b(G28), .O(gate68inter2));
  inv1  gate1558(.a(s_144), .O(gate68inter3));
  inv1  gate1559(.a(s_145), .O(gate68inter4));
  nand2 gate1560(.a(gate68inter4), .b(gate68inter3), .O(gate68inter5));
  nor2  gate1561(.a(gate68inter5), .b(gate68inter2), .O(gate68inter6));
  inv1  gate1562(.a(G28), .O(gate68inter7));
  inv1  gate1563(.a(G305), .O(gate68inter8));
  nand2 gate1564(.a(gate68inter8), .b(gate68inter7), .O(gate68inter9));
  nand2 gate1565(.a(s_145), .b(gate68inter3), .O(gate68inter10));
  nor2  gate1566(.a(gate68inter10), .b(gate68inter9), .O(gate68inter11));
  nor2  gate1567(.a(gate68inter11), .b(gate68inter6), .O(gate68inter12));
  nand2 gate1568(.a(gate68inter12), .b(gate68inter1), .O(G389));
nand2 gate69( .a(G29), .b(G308), .O(G390) );
nand2 gate70( .a(G30), .b(G308), .O(G391) );

  xor2  gate2675(.a(G311), .b(G31), .O(gate71inter0));
  nand2 gate2676(.a(gate71inter0), .b(s_304), .O(gate71inter1));
  and2  gate2677(.a(G311), .b(G31), .O(gate71inter2));
  inv1  gate2678(.a(s_304), .O(gate71inter3));
  inv1  gate2679(.a(s_305), .O(gate71inter4));
  nand2 gate2680(.a(gate71inter4), .b(gate71inter3), .O(gate71inter5));
  nor2  gate2681(.a(gate71inter5), .b(gate71inter2), .O(gate71inter6));
  inv1  gate2682(.a(G31), .O(gate71inter7));
  inv1  gate2683(.a(G311), .O(gate71inter8));
  nand2 gate2684(.a(gate71inter8), .b(gate71inter7), .O(gate71inter9));
  nand2 gate2685(.a(s_305), .b(gate71inter3), .O(gate71inter10));
  nor2  gate2686(.a(gate71inter10), .b(gate71inter9), .O(gate71inter11));
  nor2  gate2687(.a(gate71inter11), .b(gate71inter6), .O(gate71inter12));
  nand2 gate2688(.a(gate71inter12), .b(gate71inter1), .O(G392));
nand2 gate72( .a(G32), .b(G311), .O(G393) );

  xor2  gate1415(.a(G314), .b(G1), .O(gate73inter0));
  nand2 gate1416(.a(gate73inter0), .b(s_124), .O(gate73inter1));
  and2  gate1417(.a(G314), .b(G1), .O(gate73inter2));
  inv1  gate1418(.a(s_124), .O(gate73inter3));
  inv1  gate1419(.a(s_125), .O(gate73inter4));
  nand2 gate1420(.a(gate73inter4), .b(gate73inter3), .O(gate73inter5));
  nor2  gate1421(.a(gate73inter5), .b(gate73inter2), .O(gate73inter6));
  inv1  gate1422(.a(G1), .O(gate73inter7));
  inv1  gate1423(.a(G314), .O(gate73inter8));
  nand2 gate1424(.a(gate73inter8), .b(gate73inter7), .O(gate73inter9));
  nand2 gate1425(.a(s_125), .b(gate73inter3), .O(gate73inter10));
  nor2  gate1426(.a(gate73inter10), .b(gate73inter9), .O(gate73inter11));
  nor2  gate1427(.a(gate73inter11), .b(gate73inter6), .O(gate73inter12));
  nand2 gate1428(.a(gate73inter12), .b(gate73inter1), .O(G394));

  xor2  gate2647(.a(G314), .b(G5), .O(gate74inter0));
  nand2 gate2648(.a(gate74inter0), .b(s_300), .O(gate74inter1));
  and2  gate2649(.a(G314), .b(G5), .O(gate74inter2));
  inv1  gate2650(.a(s_300), .O(gate74inter3));
  inv1  gate2651(.a(s_301), .O(gate74inter4));
  nand2 gate2652(.a(gate74inter4), .b(gate74inter3), .O(gate74inter5));
  nor2  gate2653(.a(gate74inter5), .b(gate74inter2), .O(gate74inter6));
  inv1  gate2654(.a(G5), .O(gate74inter7));
  inv1  gate2655(.a(G314), .O(gate74inter8));
  nand2 gate2656(.a(gate74inter8), .b(gate74inter7), .O(gate74inter9));
  nand2 gate2657(.a(s_301), .b(gate74inter3), .O(gate74inter10));
  nor2  gate2658(.a(gate74inter10), .b(gate74inter9), .O(gate74inter11));
  nor2  gate2659(.a(gate74inter11), .b(gate74inter6), .O(gate74inter12));
  nand2 gate2660(.a(gate74inter12), .b(gate74inter1), .O(G395));
nand2 gate75( .a(G9), .b(G317), .O(G396) );

  xor2  gate1905(.a(G317), .b(G13), .O(gate76inter0));
  nand2 gate1906(.a(gate76inter0), .b(s_194), .O(gate76inter1));
  and2  gate1907(.a(G317), .b(G13), .O(gate76inter2));
  inv1  gate1908(.a(s_194), .O(gate76inter3));
  inv1  gate1909(.a(s_195), .O(gate76inter4));
  nand2 gate1910(.a(gate76inter4), .b(gate76inter3), .O(gate76inter5));
  nor2  gate1911(.a(gate76inter5), .b(gate76inter2), .O(gate76inter6));
  inv1  gate1912(.a(G13), .O(gate76inter7));
  inv1  gate1913(.a(G317), .O(gate76inter8));
  nand2 gate1914(.a(gate76inter8), .b(gate76inter7), .O(gate76inter9));
  nand2 gate1915(.a(s_195), .b(gate76inter3), .O(gate76inter10));
  nor2  gate1916(.a(gate76inter10), .b(gate76inter9), .O(gate76inter11));
  nor2  gate1917(.a(gate76inter11), .b(gate76inter6), .O(gate76inter12));
  nand2 gate1918(.a(gate76inter12), .b(gate76inter1), .O(G397));
nand2 gate77( .a(G2), .b(G320), .O(G398) );
nand2 gate78( .a(G6), .b(G320), .O(G399) );
nand2 gate79( .a(G10), .b(G323), .O(G400) );
nand2 gate80( .a(G14), .b(G323), .O(G401) );
nand2 gate81( .a(G3), .b(G326), .O(G402) );
nand2 gate82( .a(G7), .b(G326), .O(G403) );
nand2 gate83( .a(G11), .b(G329), .O(G404) );

  xor2  gate547(.a(G329), .b(G15), .O(gate84inter0));
  nand2 gate548(.a(gate84inter0), .b(s_0), .O(gate84inter1));
  and2  gate549(.a(G329), .b(G15), .O(gate84inter2));
  inv1  gate550(.a(s_0), .O(gate84inter3));
  inv1  gate551(.a(s_1), .O(gate84inter4));
  nand2 gate552(.a(gate84inter4), .b(gate84inter3), .O(gate84inter5));
  nor2  gate553(.a(gate84inter5), .b(gate84inter2), .O(gate84inter6));
  inv1  gate554(.a(G15), .O(gate84inter7));
  inv1  gate555(.a(G329), .O(gate84inter8));
  nand2 gate556(.a(gate84inter8), .b(gate84inter7), .O(gate84inter9));
  nand2 gate557(.a(s_1), .b(gate84inter3), .O(gate84inter10));
  nor2  gate558(.a(gate84inter10), .b(gate84inter9), .O(gate84inter11));
  nor2  gate559(.a(gate84inter11), .b(gate84inter6), .O(gate84inter12));
  nand2 gate560(.a(gate84inter12), .b(gate84inter1), .O(G405));
nand2 gate85( .a(G4), .b(G332), .O(G406) );

  xor2  gate1149(.a(G332), .b(G8), .O(gate86inter0));
  nand2 gate1150(.a(gate86inter0), .b(s_86), .O(gate86inter1));
  and2  gate1151(.a(G332), .b(G8), .O(gate86inter2));
  inv1  gate1152(.a(s_86), .O(gate86inter3));
  inv1  gate1153(.a(s_87), .O(gate86inter4));
  nand2 gate1154(.a(gate86inter4), .b(gate86inter3), .O(gate86inter5));
  nor2  gate1155(.a(gate86inter5), .b(gate86inter2), .O(gate86inter6));
  inv1  gate1156(.a(G8), .O(gate86inter7));
  inv1  gate1157(.a(G332), .O(gate86inter8));
  nand2 gate1158(.a(gate86inter8), .b(gate86inter7), .O(gate86inter9));
  nand2 gate1159(.a(s_87), .b(gate86inter3), .O(gate86inter10));
  nor2  gate1160(.a(gate86inter10), .b(gate86inter9), .O(gate86inter11));
  nor2  gate1161(.a(gate86inter11), .b(gate86inter6), .O(gate86inter12));
  nand2 gate1162(.a(gate86inter12), .b(gate86inter1), .O(G407));
nand2 gate87( .a(G12), .b(G335), .O(G408) );
nand2 gate88( .a(G16), .b(G335), .O(G409) );
nand2 gate89( .a(G17), .b(G338), .O(G410) );
nand2 gate90( .a(G21), .b(G338), .O(G411) );

  xor2  gate1597(.a(G341), .b(G25), .O(gate91inter0));
  nand2 gate1598(.a(gate91inter0), .b(s_150), .O(gate91inter1));
  and2  gate1599(.a(G341), .b(G25), .O(gate91inter2));
  inv1  gate1600(.a(s_150), .O(gate91inter3));
  inv1  gate1601(.a(s_151), .O(gate91inter4));
  nand2 gate1602(.a(gate91inter4), .b(gate91inter3), .O(gate91inter5));
  nor2  gate1603(.a(gate91inter5), .b(gate91inter2), .O(gate91inter6));
  inv1  gate1604(.a(G25), .O(gate91inter7));
  inv1  gate1605(.a(G341), .O(gate91inter8));
  nand2 gate1606(.a(gate91inter8), .b(gate91inter7), .O(gate91inter9));
  nand2 gate1607(.a(s_151), .b(gate91inter3), .O(gate91inter10));
  nor2  gate1608(.a(gate91inter10), .b(gate91inter9), .O(gate91inter11));
  nor2  gate1609(.a(gate91inter11), .b(gate91inter6), .O(gate91inter12));
  nand2 gate1610(.a(gate91inter12), .b(gate91inter1), .O(G412));

  xor2  gate1835(.a(G341), .b(G29), .O(gate92inter0));
  nand2 gate1836(.a(gate92inter0), .b(s_184), .O(gate92inter1));
  and2  gate1837(.a(G341), .b(G29), .O(gate92inter2));
  inv1  gate1838(.a(s_184), .O(gate92inter3));
  inv1  gate1839(.a(s_185), .O(gate92inter4));
  nand2 gate1840(.a(gate92inter4), .b(gate92inter3), .O(gate92inter5));
  nor2  gate1841(.a(gate92inter5), .b(gate92inter2), .O(gate92inter6));
  inv1  gate1842(.a(G29), .O(gate92inter7));
  inv1  gate1843(.a(G341), .O(gate92inter8));
  nand2 gate1844(.a(gate92inter8), .b(gate92inter7), .O(gate92inter9));
  nand2 gate1845(.a(s_185), .b(gate92inter3), .O(gate92inter10));
  nor2  gate1846(.a(gate92inter10), .b(gate92inter9), .O(gate92inter11));
  nor2  gate1847(.a(gate92inter11), .b(gate92inter6), .O(gate92inter12));
  nand2 gate1848(.a(gate92inter12), .b(gate92inter1), .O(G413));
nand2 gate93( .a(G18), .b(G344), .O(G414) );
nand2 gate94( .a(G22), .b(G344), .O(G415) );
nand2 gate95( .a(G26), .b(G347), .O(G416) );
nand2 gate96( .a(G30), .b(G347), .O(G417) );
nand2 gate97( .a(G19), .b(G350), .O(G418) );
nand2 gate98( .a(G23), .b(G350), .O(G419) );
nand2 gate99( .a(G27), .b(G353), .O(G420) );

  xor2  gate1345(.a(G353), .b(G31), .O(gate100inter0));
  nand2 gate1346(.a(gate100inter0), .b(s_114), .O(gate100inter1));
  and2  gate1347(.a(G353), .b(G31), .O(gate100inter2));
  inv1  gate1348(.a(s_114), .O(gate100inter3));
  inv1  gate1349(.a(s_115), .O(gate100inter4));
  nand2 gate1350(.a(gate100inter4), .b(gate100inter3), .O(gate100inter5));
  nor2  gate1351(.a(gate100inter5), .b(gate100inter2), .O(gate100inter6));
  inv1  gate1352(.a(G31), .O(gate100inter7));
  inv1  gate1353(.a(G353), .O(gate100inter8));
  nand2 gate1354(.a(gate100inter8), .b(gate100inter7), .O(gate100inter9));
  nand2 gate1355(.a(s_115), .b(gate100inter3), .O(gate100inter10));
  nor2  gate1356(.a(gate100inter10), .b(gate100inter9), .O(gate100inter11));
  nor2  gate1357(.a(gate100inter11), .b(gate100inter6), .O(gate100inter12));
  nand2 gate1358(.a(gate100inter12), .b(gate100inter1), .O(G421));

  xor2  gate2661(.a(G356), .b(G20), .O(gate101inter0));
  nand2 gate2662(.a(gate101inter0), .b(s_302), .O(gate101inter1));
  and2  gate2663(.a(G356), .b(G20), .O(gate101inter2));
  inv1  gate2664(.a(s_302), .O(gate101inter3));
  inv1  gate2665(.a(s_303), .O(gate101inter4));
  nand2 gate2666(.a(gate101inter4), .b(gate101inter3), .O(gate101inter5));
  nor2  gate2667(.a(gate101inter5), .b(gate101inter2), .O(gate101inter6));
  inv1  gate2668(.a(G20), .O(gate101inter7));
  inv1  gate2669(.a(G356), .O(gate101inter8));
  nand2 gate2670(.a(gate101inter8), .b(gate101inter7), .O(gate101inter9));
  nand2 gate2671(.a(s_303), .b(gate101inter3), .O(gate101inter10));
  nor2  gate2672(.a(gate101inter10), .b(gate101inter9), .O(gate101inter11));
  nor2  gate2673(.a(gate101inter11), .b(gate101inter6), .O(gate101inter12));
  nand2 gate2674(.a(gate101inter12), .b(gate101inter1), .O(G422));
nand2 gate102( .a(G24), .b(G356), .O(G423) );
nand2 gate103( .a(G28), .b(G359), .O(G424) );
nand2 gate104( .a(G32), .b(G359), .O(G425) );

  xor2  gate2423(.a(G363), .b(G362), .O(gate105inter0));
  nand2 gate2424(.a(gate105inter0), .b(s_268), .O(gate105inter1));
  and2  gate2425(.a(G363), .b(G362), .O(gate105inter2));
  inv1  gate2426(.a(s_268), .O(gate105inter3));
  inv1  gate2427(.a(s_269), .O(gate105inter4));
  nand2 gate2428(.a(gate105inter4), .b(gate105inter3), .O(gate105inter5));
  nor2  gate2429(.a(gate105inter5), .b(gate105inter2), .O(gate105inter6));
  inv1  gate2430(.a(G362), .O(gate105inter7));
  inv1  gate2431(.a(G363), .O(gate105inter8));
  nand2 gate2432(.a(gate105inter8), .b(gate105inter7), .O(gate105inter9));
  nand2 gate2433(.a(s_269), .b(gate105inter3), .O(gate105inter10));
  nor2  gate2434(.a(gate105inter10), .b(gate105inter9), .O(gate105inter11));
  nor2  gate2435(.a(gate105inter11), .b(gate105inter6), .O(gate105inter12));
  nand2 gate2436(.a(gate105inter12), .b(gate105inter1), .O(G426));
nand2 gate106( .a(G364), .b(G365), .O(G429) );
nand2 gate107( .a(G366), .b(G367), .O(G432) );

  xor2  gate2199(.a(G369), .b(G368), .O(gate108inter0));
  nand2 gate2200(.a(gate108inter0), .b(s_236), .O(gate108inter1));
  and2  gate2201(.a(G369), .b(G368), .O(gate108inter2));
  inv1  gate2202(.a(s_236), .O(gate108inter3));
  inv1  gate2203(.a(s_237), .O(gate108inter4));
  nand2 gate2204(.a(gate108inter4), .b(gate108inter3), .O(gate108inter5));
  nor2  gate2205(.a(gate108inter5), .b(gate108inter2), .O(gate108inter6));
  inv1  gate2206(.a(G368), .O(gate108inter7));
  inv1  gate2207(.a(G369), .O(gate108inter8));
  nand2 gate2208(.a(gate108inter8), .b(gate108inter7), .O(gate108inter9));
  nand2 gate2209(.a(s_237), .b(gate108inter3), .O(gate108inter10));
  nor2  gate2210(.a(gate108inter10), .b(gate108inter9), .O(gate108inter11));
  nor2  gate2211(.a(gate108inter11), .b(gate108inter6), .O(gate108inter12));
  nand2 gate2212(.a(gate108inter12), .b(gate108inter1), .O(G435));

  xor2  gate1947(.a(G371), .b(G370), .O(gate109inter0));
  nand2 gate1948(.a(gate109inter0), .b(s_200), .O(gate109inter1));
  and2  gate1949(.a(G371), .b(G370), .O(gate109inter2));
  inv1  gate1950(.a(s_200), .O(gate109inter3));
  inv1  gate1951(.a(s_201), .O(gate109inter4));
  nand2 gate1952(.a(gate109inter4), .b(gate109inter3), .O(gate109inter5));
  nor2  gate1953(.a(gate109inter5), .b(gate109inter2), .O(gate109inter6));
  inv1  gate1954(.a(G370), .O(gate109inter7));
  inv1  gate1955(.a(G371), .O(gate109inter8));
  nand2 gate1956(.a(gate109inter8), .b(gate109inter7), .O(gate109inter9));
  nand2 gate1957(.a(s_201), .b(gate109inter3), .O(gate109inter10));
  nor2  gate1958(.a(gate109inter10), .b(gate109inter9), .O(gate109inter11));
  nor2  gate1959(.a(gate109inter11), .b(gate109inter6), .O(gate109inter12));
  nand2 gate1960(.a(gate109inter12), .b(gate109inter1), .O(G438));
nand2 gate110( .a(G372), .b(G373), .O(G441) );
nand2 gate111( .a(G374), .b(G375), .O(G444) );

  xor2  gate631(.a(G377), .b(G376), .O(gate112inter0));
  nand2 gate632(.a(gate112inter0), .b(s_12), .O(gate112inter1));
  and2  gate633(.a(G377), .b(G376), .O(gate112inter2));
  inv1  gate634(.a(s_12), .O(gate112inter3));
  inv1  gate635(.a(s_13), .O(gate112inter4));
  nand2 gate636(.a(gate112inter4), .b(gate112inter3), .O(gate112inter5));
  nor2  gate637(.a(gate112inter5), .b(gate112inter2), .O(gate112inter6));
  inv1  gate638(.a(G376), .O(gate112inter7));
  inv1  gate639(.a(G377), .O(gate112inter8));
  nand2 gate640(.a(gate112inter8), .b(gate112inter7), .O(gate112inter9));
  nand2 gate641(.a(s_13), .b(gate112inter3), .O(gate112inter10));
  nor2  gate642(.a(gate112inter10), .b(gate112inter9), .O(gate112inter11));
  nor2  gate643(.a(gate112inter11), .b(gate112inter6), .O(gate112inter12));
  nand2 gate644(.a(gate112inter12), .b(gate112inter1), .O(G447));
nand2 gate113( .a(G378), .b(G379), .O(G450) );
nand2 gate114( .a(G380), .b(G381), .O(G453) );
nand2 gate115( .a(G382), .b(G383), .O(G456) );
nand2 gate116( .a(G384), .b(G385), .O(G459) );
nand2 gate117( .a(G386), .b(G387), .O(G462) );
nand2 gate118( .a(G388), .b(G389), .O(G465) );

  xor2  gate701(.a(G391), .b(G390), .O(gate119inter0));
  nand2 gate702(.a(gate119inter0), .b(s_22), .O(gate119inter1));
  and2  gate703(.a(G391), .b(G390), .O(gate119inter2));
  inv1  gate704(.a(s_22), .O(gate119inter3));
  inv1  gate705(.a(s_23), .O(gate119inter4));
  nand2 gate706(.a(gate119inter4), .b(gate119inter3), .O(gate119inter5));
  nor2  gate707(.a(gate119inter5), .b(gate119inter2), .O(gate119inter6));
  inv1  gate708(.a(G390), .O(gate119inter7));
  inv1  gate709(.a(G391), .O(gate119inter8));
  nand2 gate710(.a(gate119inter8), .b(gate119inter7), .O(gate119inter9));
  nand2 gate711(.a(s_23), .b(gate119inter3), .O(gate119inter10));
  nor2  gate712(.a(gate119inter10), .b(gate119inter9), .O(gate119inter11));
  nor2  gate713(.a(gate119inter11), .b(gate119inter6), .O(gate119inter12));
  nand2 gate714(.a(gate119inter12), .b(gate119inter1), .O(G468));

  xor2  gate2297(.a(G393), .b(G392), .O(gate120inter0));
  nand2 gate2298(.a(gate120inter0), .b(s_250), .O(gate120inter1));
  and2  gate2299(.a(G393), .b(G392), .O(gate120inter2));
  inv1  gate2300(.a(s_250), .O(gate120inter3));
  inv1  gate2301(.a(s_251), .O(gate120inter4));
  nand2 gate2302(.a(gate120inter4), .b(gate120inter3), .O(gate120inter5));
  nor2  gate2303(.a(gate120inter5), .b(gate120inter2), .O(gate120inter6));
  inv1  gate2304(.a(G392), .O(gate120inter7));
  inv1  gate2305(.a(G393), .O(gate120inter8));
  nand2 gate2306(.a(gate120inter8), .b(gate120inter7), .O(gate120inter9));
  nand2 gate2307(.a(s_251), .b(gate120inter3), .O(gate120inter10));
  nor2  gate2308(.a(gate120inter10), .b(gate120inter9), .O(gate120inter11));
  nor2  gate2309(.a(gate120inter11), .b(gate120inter6), .O(gate120inter12));
  nand2 gate2310(.a(gate120inter12), .b(gate120inter1), .O(G471));
nand2 gate121( .a(G394), .b(G395), .O(G474) );
nand2 gate122( .a(G396), .b(G397), .O(G477) );
nand2 gate123( .a(G398), .b(G399), .O(G480) );
nand2 gate124( .a(G400), .b(G401), .O(G483) );
nand2 gate125( .a(G402), .b(G403), .O(G486) );

  xor2  gate939(.a(G405), .b(G404), .O(gate126inter0));
  nand2 gate940(.a(gate126inter0), .b(s_56), .O(gate126inter1));
  and2  gate941(.a(G405), .b(G404), .O(gate126inter2));
  inv1  gate942(.a(s_56), .O(gate126inter3));
  inv1  gate943(.a(s_57), .O(gate126inter4));
  nand2 gate944(.a(gate126inter4), .b(gate126inter3), .O(gate126inter5));
  nor2  gate945(.a(gate126inter5), .b(gate126inter2), .O(gate126inter6));
  inv1  gate946(.a(G404), .O(gate126inter7));
  inv1  gate947(.a(G405), .O(gate126inter8));
  nand2 gate948(.a(gate126inter8), .b(gate126inter7), .O(gate126inter9));
  nand2 gate949(.a(s_57), .b(gate126inter3), .O(gate126inter10));
  nor2  gate950(.a(gate126inter10), .b(gate126inter9), .O(gate126inter11));
  nor2  gate951(.a(gate126inter11), .b(gate126inter6), .O(gate126inter12));
  nand2 gate952(.a(gate126inter12), .b(gate126inter1), .O(G489));
nand2 gate127( .a(G406), .b(G407), .O(G492) );
nand2 gate128( .a(G408), .b(G409), .O(G495) );

  xor2  gate2129(.a(G411), .b(G410), .O(gate129inter0));
  nand2 gate2130(.a(gate129inter0), .b(s_226), .O(gate129inter1));
  and2  gate2131(.a(G411), .b(G410), .O(gate129inter2));
  inv1  gate2132(.a(s_226), .O(gate129inter3));
  inv1  gate2133(.a(s_227), .O(gate129inter4));
  nand2 gate2134(.a(gate129inter4), .b(gate129inter3), .O(gate129inter5));
  nor2  gate2135(.a(gate129inter5), .b(gate129inter2), .O(gate129inter6));
  inv1  gate2136(.a(G410), .O(gate129inter7));
  inv1  gate2137(.a(G411), .O(gate129inter8));
  nand2 gate2138(.a(gate129inter8), .b(gate129inter7), .O(gate129inter9));
  nand2 gate2139(.a(s_227), .b(gate129inter3), .O(gate129inter10));
  nor2  gate2140(.a(gate129inter10), .b(gate129inter9), .O(gate129inter11));
  nor2  gate2141(.a(gate129inter11), .b(gate129inter6), .O(gate129inter12));
  nand2 gate2142(.a(gate129inter12), .b(gate129inter1), .O(G498));
nand2 gate130( .a(G412), .b(G413), .O(G501) );
nand2 gate131( .a(G414), .b(G415), .O(G504) );
nand2 gate132( .a(G416), .b(G417), .O(G507) );
nand2 gate133( .a(G418), .b(G419), .O(G510) );
nand2 gate134( .a(G420), .b(G421), .O(G513) );
nand2 gate135( .a(G422), .b(G423), .O(G516) );
nand2 gate136( .a(G424), .b(G425), .O(G519) );
nand2 gate137( .a(G426), .b(G429), .O(G522) );
nand2 gate138( .a(G432), .b(G435), .O(G525) );
nand2 gate139( .a(G438), .b(G441), .O(G528) );
nand2 gate140( .a(G444), .b(G447), .O(G531) );

  xor2  gate2549(.a(G453), .b(G450), .O(gate141inter0));
  nand2 gate2550(.a(gate141inter0), .b(s_286), .O(gate141inter1));
  and2  gate2551(.a(G453), .b(G450), .O(gate141inter2));
  inv1  gate2552(.a(s_286), .O(gate141inter3));
  inv1  gate2553(.a(s_287), .O(gate141inter4));
  nand2 gate2554(.a(gate141inter4), .b(gate141inter3), .O(gate141inter5));
  nor2  gate2555(.a(gate141inter5), .b(gate141inter2), .O(gate141inter6));
  inv1  gate2556(.a(G450), .O(gate141inter7));
  inv1  gate2557(.a(G453), .O(gate141inter8));
  nand2 gate2558(.a(gate141inter8), .b(gate141inter7), .O(gate141inter9));
  nand2 gate2559(.a(s_287), .b(gate141inter3), .O(gate141inter10));
  nor2  gate2560(.a(gate141inter10), .b(gate141inter9), .O(gate141inter11));
  nor2  gate2561(.a(gate141inter11), .b(gate141inter6), .O(gate141inter12));
  nand2 gate2562(.a(gate141inter12), .b(gate141inter1), .O(G534));

  xor2  gate2521(.a(G459), .b(G456), .O(gate142inter0));
  nand2 gate2522(.a(gate142inter0), .b(s_282), .O(gate142inter1));
  and2  gate2523(.a(G459), .b(G456), .O(gate142inter2));
  inv1  gate2524(.a(s_282), .O(gate142inter3));
  inv1  gate2525(.a(s_283), .O(gate142inter4));
  nand2 gate2526(.a(gate142inter4), .b(gate142inter3), .O(gate142inter5));
  nor2  gate2527(.a(gate142inter5), .b(gate142inter2), .O(gate142inter6));
  inv1  gate2528(.a(G456), .O(gate142inter7));
  inv1  gate2529(.a(G459), .O(gate142inter8));
  nand2 gate2530(.a(gate142inter8), .b(gate142inter7), .O(gate142inter9));
  nand2 gate2531(.a(s_283), .b(gate142inter3), .O(gate142inter10));
  nor2  gate2532(.a(gate142inter10), .b(gate142inter9), .O(gate142inter11));
  nor2  gate2533(.a(gate142inter11), .b(gate142inter6), .O(gate142inter12));
  nand2 gate2534(.a(gate142inter12), .b(gate142inter1), .O(G537));

  xor2  gate2185(.a(G465), .b(G462), .O(gate143inter0));
  nand2 gate2186(.a(gate143inter0), .b(s_234), .O(gate143inter1));
  and2  gate2187(.a(G465), .b(G462), .O(gate143inter2));
  inv1  gate2188(.a(s_234), .O(gate143inter3));
  inv1  gate2189(.a(s_235), .O(gate143inter4));
  nand2 gate2190(.a(gate143inter4), .b(gate143inter3), .O(gate143inter5));
  nor2  gate2191(.a(gate143inter5), .b(gate143inter2), .O(gate143inter6));
  inv1  gate2192(.a(G462), .O(gate143inter7));
  inv1  gate2193(.a(G465), .O(gate143inter8));
  nand2 gate2194(.a(gate143inter8), .b(gate143inter7), .O(gate143inter9));
  nand2 gate2195(.a(s_235), .b(gate143inter3), .O(gate143inter10));
  nor2  gate2196(.a(gate143inter10), .b(gate143inter9), .O(gate143inter11));
  nor2  gate2197(.a(gate143inter11), .b(gate143inter6), .O(gate143inter12));
  nand2 gate2198(.a(gate143inter12), .b(gate143inter1), .O(G540));
nand2 gate144( .a(G468), .b(G471), .O(G543) );
nand2 gate145( .a(G474), .b(G477), .O(G546) );
nand2 gate146( .a(G480), .b(G483), .O(G549) );
nand2 gate147( .a(G486), .b(G489), .O(G552) );
nand2 gate148( .a(G492), .b(G495), .O(G555) );
nand2 gate149( .a(G498), .b(G501), .O(G558) );
nand2 gate150( .a(G504), .b(G507), .O(G561) );

  xor2  gate2059(.a(G513), .b(G510), .O(gate151inter0));
  nand2 gate2060(.a(gate151inter0), .b(s_216), .O(gate151inter1));
  and2  gate2061(.a(G513), .b(G510), .O(gate151inter2));
  inv1  gate2062(.a(s_216), .O(gate151inter3));
  inv1  gate2063(.a(s_217), .O(gate151inter4));
  nand2 gate2064(.a(gate151inter4), .b(gate151inter3), .O(gate151inter5));
  nor2  gate2065(.a(gate151inter5), .b(gate151inter2), .O(gate151inter6));
  inv1  gate2066(.a(G510), .O(gate151inter7));
  inv1  gate2067(.a(G513), .O(gate151inter8));
  nand2 gate2068(.a(gate151inter8), .b(gate151inter7), .O(gate151inter9));
  nand2 gate2069(.a(s_217), .b(gate151inter3), .O(gate151inter10));
  nor2  gate2070(.a(gate151inter10), .b(gate151inter9), .O(gate151inter11));
  nor2  gate2071(.a(gate151inter11), .b(gate151inter6), .O(gate151inter12));
  nand2 gate2072(.a(gate151inter12), .b(gate151inter1), .O(G564));

  xor2  gate1079(.a(G519), .b(G516), .O(gate152inter0));
  nand2 gate1080(.a(gate152inter0), .b(s_76), .O(gate152inter1));
  and2  gate1081(.a(G519), .b(G516), .O(gate152inter2));
  inv1  gate1082(.a(s_76), .O(gate152inter3));
  inv1  gate1083(.a(s_77), .O(gate152inter4));
  nand2 gate1084(.a(gate152inter4), .b(gate152inter3), .O(gate152inter5));
  nor2  gate1085(.a(gate152inter5), .b(gate152inter2), .O(gate152inter6));
  inv1  gate1086(.a(G516), .O(gate152inter7));
  inv1  gate1087(.a(G519), .O(gate152inter8));
  nand2 gate1088(.a(gate152inter8), .b(gate152inter7), .O(gate152inter9));
  nand2 gate1089(.a(s_77), .b(gate152inter3), .O(gate152inter10));
  nor2  gate1090(.a(gate152inter10), .b(gate152inter9), .O(gate152inter11));
  nor2  gate1091(.a(gate152inter11), .b(gate152inter6), .O(gate152inter12));
  nand2 gate1092(.a(gate152inter12), .b(gate152inter1), .O(G567));
nand2 gate153( .a(G426), .b(G522), .O(G570) );
nand2 gate154( .a(G429), .b(G522), .O(G571) );
nand2 gate155( .a(G432), .b(G525), .O(G572) );
nand2 gate156( .a(G435), .b(G525), .O(G573) );

  xor2  gate2633(.a(G528), .b(G438), .O(gate157inter0));
  nand2 gate2634(.a(gate157inter0), .b(s_298), .O(gate157inter1));
  and2  gate2635(.a(G528), .b(G438), .O(gate157inter2));
  inv1  gate2636(.a(s_298), .O(gate157inter3));
  inv1  gate2637(.a(s_299), .O(gate157inter4));
  nand2 gate2638(.a(gate157inter4), .b(gate157inter3), .O(gate157inter5));
  nor2  gate2639(.a(gate157inter5), .b(gate157inter2), .O(gate157inter6));
  inv1  gate2640(.a(G438), .O(gate157inter7));
  inv1  gate2641(.a(G528), .O(gate157inter8));
  nand2 gate2642(.a(gate157inter8), .b(gate157inter7), .O(gate157inter9));
  nand2 gate2643(.a(s_299), .b(gate157inter3), .O(gate157inter10));
  nor2  gate2644(.a(gate157inter10), .b(gate157inter9), .O(gate157inter11));
  nor2  gate2645(.a(gate157inter11), .b(gate157inter6), .O(gate157inter12));
  nand2 gate2646(.a(gate157inter12), .b(gate157inter1), .O(G574));
nand2 gate158( .a(G441), .b(G528), .O(G575) );
nand2 gate159( .a(G444), .b(G531), .O(G576) );

  xor2  gate1933(.a(G531), .b(G447), .O(gate160inter0));
  nand2 gate1934(.a(gate160inter0), .b(s_198), .O(gate160inter1));
  and2  gate1935(.a(G531), .b(G447), .O(gate160inter2));
  inv1  gate1936(.a(s_198), .O(gate160inter3));
  inv1  gate1937(.a(s_199), .O(gate160inter4));
  nand2 gate1938(.a(gate160inter4), .b(gate160inter3), .O(gate160inter5));
  nor2  gate1939(.a(gate160inter5), .b(gate160inter2), .O(gate160inter6));
  inv1  gate1940(.a(G447), .O(gate160inter7));
  inv1  gate1941(.a(G531), .O(gate160inter8));
  nand2 gate1942(.a(gate160inter8), .b(gate160inter7), .O(gate160inter9));
  nand2 gate1943(.a(s_199), .b(gate160inter3), .O(gate160inter10));
  nor2  gate1944(.a(gate160inter10), .b(gate160inter9), .O(gate160inter11));
  nor2  gate1945(.a(gate160inter11), .b(gate160inter6), .O(gate160inter12));
  nand2 gate1946(.a(gate160inter12), .b(gate160inter1), .O(G577));
nand2 gate161( .a(G450), .b(G534), .O(G578) );

  xor2  gate1303(.a(G534), .b(G453), .O(gate162inter0));
  nand2 gate1304(.a(gate162inter0), .b(s_108), .O(gate162inter1));
  and2  gate1305(.a(G534), .b(G453), .O(gate162inter2));
  inv1  gate1306(.a(s_108), .O(gate162inter3));
  inv1  gate1307(.a(s_109), .O(gate162inter4));
  nand2 gate1308(.a(gate162inter4), .b(gate162inter3), .O(gate162inter5));
  nor2  gate1309(.a(gate162inter5), .b(gate162inter2), .O(gate162inter6));
  inv1  gate1310(.a(G453), .O(gate162inter7));
  inv1  gate1311(.a(G534), .O(gate162inter8));
  nand2 gate1312(.a(gate162inter8), .b(gate162inter7), .O(gate162inter9));
  nand2 gate1313(.a(s_109), .b(gate162inter3), .O(gate162inter10));
  nor2  gate1314(.a(gate162inter10), .b(gate162inter9), .O(gate162inter11));
  nor2  gate1315(.a(gate162inter11), .b(gate162inter6), .O(gate162inter12));
  nand2 gate1316(.a(gate162inter12), .b(gate162inter1), .O(G579));

  xor2  gate2577(.a(G537), .b(G456), .O(gate163inter0));
  nand2 gate2578(.a(gate163inter0), .b(s_290), .O(gate163inter1));
  and2  gate2579(.a(G537), .b(G456), .O(gate163inter2));
  inv1  gate2580(.a(s_290), .O(gate163inter3));
  inv1  gate2581(.a(s_291), .O(gate163inter4));
  nand2 gate2582(.a(gate163inter4), .b(gate163inter3), .O(gate163inter5));
  nor2  gate2583(.a(gate163inter5), .b(gate163inter2), .O(gate163inter6));
  inv1  gate2584(.a(G456), .O(gate163inter7));
  inv1  gate2585(.a(G537), .O(gate163inter8));
  nand2 gate2586(.a(gate163inter8), .b(gate163inter7), .O(gate163inter9));
  nand2 gate2587(.a(s_291), .b(gate163inter3), .O(gate163inter10));
  nor2  gate2588(.a(gate163inter10), .b(gate163inter9), .O(gate163inter11));
  nor2  gate2589(.a(gate163inter11), .b(gate163inter6), .O(gate163inter12));
  nand2 gate2590(.a(gate163inter12), .b(gate163inter1), .O(G580));
nand2 gate164( .a(G459), .b(G537), .O(G581) );

  xor2  gate1359(.a(G540), .b(G462), .O(gate165inter0));
  nand2 gate1360(.a(gate165inter0), .b(s_116), .O(gate165inter1));
  and2  gate1361(.a(G540), .b(G462), .O(gate165inter2));
  inv1  gate1362(.a(s_116), .O(gate165inter3));
  inv1  gate1363(.a(s_117), .O(gate165inter4));
  nand2 gate1364(.a(gate165inter4), .b(gate165inter3), .O(gate165inter5));
  nor2  gate1365(.a(gate165inter5), .b(gate165inter2), .O(gate165inter6));
  inv1  gate1366(.a(G462), .O(gate165inter7));
  inv1  gate1367(.a(G540), .O(gate165inter8));
  nand2 gate1368(.a(gate165inter8), .b(gate165inter7), .O(gate165inter9));
  nand2 gate1369(.a(s_117), .b(gate165inter3), .O(gate165inter10));
  nor2  gate1370(.a(gate165inter10), .b(gate165inter9), .O(gate165inter11));
  nor2  gate1371(.a(gate165inter11), .b(gate165inter6), .O(gate165inter12));
  nand2 gate1372(.a(gate165inter12), .b(gate165inter1), .O(G582));
nand2 gate166( .a(G465), .b(G540), .O(G583) );
nand2 gate167( .a(G468), .b(G543), .O(G584) );
nand2 gate168( .a(G471), .b(G543), .O(G585) );
nand2 gate169( .a(G474), .b(G546), .O(G586) );
nand2 gate170( .a(G477), .b(G546), .O(G587) );

  xor2  gate1821(.a(G549), .b(G480), .O(gate171inter0));
  nand2 gate1822(.a(gate171inter0), .b(s_182), .O(gate171inter1));
  and2  gate1823(.a(G549), .b(G480), .O(gate171inter2));
  inv1  gate1824(.a(s_182), .O(gate171inter3));
  inv1  gate1825(.a(s_183), .O(gate171inter4));
  nand2 gate1826(.a(gate171inter4), .b(gate171inter3), .O(gate171inter5));
  nor2  gate1827(.a(gate171inter5), .b(gate171inter2), .O(gate171inter6));
  inv1  gate1828(.a(G480), .O(gate171inter7));
  inv1  gate1829(.a(G549), .O(gate171inter8));
  nand2 gate1830(.a(gate171inter8), .b(gate171inter7), .O(gate171inter9));
  nand2 gate1831(.a(s_183), .b(gate171inter3), .O(gate171inter10));
  nor2  gate1832(.a(gate171inter10), .b(gate171inter9), .O(gate171inter11));
  nor2  gate1833(.a(gate171inter11), .b(gate171inter6), .O(gate171inter12));
  nand2 gate1834(.a(gate171inter12), .b(gate171inter1), .O(G588));

  xor2  gate645(.a(G549), .b(G483), .O(gate172inter0));
  nand2 gate646(.a(gate172inter0), .b(s_14), .O(gate172inter1));
  and2  gate647(.a(G549), .b(G483), .O(gate172inter2));
  inv1  gate648(.a(s_14), .O(gate172inter3));
  inv1  gate649(.a(s_15), .O(gate172inter4));
  nand2 gate650(.a(gate172inter4), .b(gate172inter3), .O(gate172inter5));
  nor2  gate651(.a(gate172inter5), .b(gate172inter2), .O(gate172inter6));
  inv1  gate652(.a(G483), .O(gate172inter7));
  inv1  gate653(.a(G549), .O(gate172inter8));
  nand2 gate654(.a(gate172inter8), .b(gate172inter7), .O(gate172inter9));
  nand2 gate655(.a(s_15), .b(gate172inter3), .O(gate172inter10));
  nor2  gate656(.a(gate172inter10), .b(gate172inter9), .O(gate172inter11));
  nor2  gate657(.a(gate172inter11), .b(gate172inter6), .O(gate172inter12));
  nand2 gate658(.a(gate172inter12), .b(gate172inter1), .O(G589));

  xor2  gate2087(.a(G552), .b(G486), .O(gate173inter0));
  nand2 gate2088(.a(gate173inter0), .b(s_220), .O(gate173inter1));
  and2  gate2089(.a(G552), .b(G486), .O(gate173inter2));
  inv1  gate2090(.a(s_220), .O(gate173inter3));
  inv1  gate2091(.a(s_221), .O(gate173inter4));
  nand2 gate2092(.a(gate173inter4), .b(gate173inter3), .O(gate173inter5));
  nor2  gate2093(.a(gate173inter5), .b(gate173inter2), .O(gate173inter6));
  inv1  gate2094(.a(G486), .O(gate173inter7));
  inv1  gate2095(.a(G552), .O(gate173inter8));
  nand2 gate2096(.a(gate173inter8), .b(gate173inter7), .O(gate173inter9));
  nand2 gate2097(.a(s_221), .b(gate173inter3), .O(gate173inter10));
  nor2  gate2098(.a(gate173inter10), .b(gate173inter9), .O(gate173inter11));
  nor2  gate2099(.a(gate173inter11), .b(gate173inter6), .O(gate173inter12));
  nand2 gate2100(.a(gate173inter12), .b(gate173inter1), .O(G590));
nand2 gate174( .a(G489), .b(G552), .O(G591) );
nand2 gate175( .a(G492), .b(G555), .O(G592) );
nand2 gate176( .a(G495), .b(G555), .O(G593) );

  xor2  gate1583(.a(G558), .b(G498), .O(gate177inter0));
  nand2 gate1584(.a(gate177inter0), .b(s_148), .O(gate177inter1));
  and2  gate1585(.a(G558), .b(G498), .O(gate177inter2));
  inv1  gate1586(.a(s_148), .O(gate177inter3));
  inv1  gate1587(.a(s_149), .O(gate177inter4));
  nand2 gate1588(.a(gate177inter4), .b(gate177inter3), .O(gate177inter5));
  nor2  gate1589(.a(gate177inter5), .b(gate177inter2), .O(gate177inter6));
  inv1  gate1590(.a(G498), .O(gate177inter7));
  inv1  gate1591(.a(G558), .O(gate177inter8));
  nand2 gate1592(.a(gate177inter8), .b(gate177inter7), .O(gate177inter9));
  nand2 gate1593(.a(s_149), .b(gate177inter3), .O(gate177inter10));
  nor2  gate1594(.a(gate177inter10), .b(gate177inter9), .O(gate177inter11));
  nor2  gate1595(.a(gate177inter11), .b(gate177inter6), .O(gate177inter12));
  nand2 gate1596(.a(gate177inter12), .b(gate177inter1), .O(G594));
nand2 gate178( .a(G501), .b(G558), .O(G595) );

  xor2  gate2437(.a(G561), .b(G504), .O(gate179inter0));
  nand2 gate2438(.a(gate179inter0), .b(s_270), .O(gate179inter1));
  and2  gate2439(.a(G561), .b(G504), .O(gate179inter2));
  inv1  gate2440(.a(s_270), .O(gate179inter3));
  inv1  gate2441(.a(s_271), .O(gate179inter4));
  nand2 gate2442(.a(gate179inter4), .b(gate179inter3), .O(gate179inter5));
  nor2  gate2443(.a(gate179inter5), .b(gate179inter2), .O(gate179inter6));
  inv1  gate2444(.a(G504), .O(gate179inter7));
  inv1  gate2445(.a(G561), .O(gate179inter8));
  nand2 gate2446(.a(gate179inter8), .b(gate179inter7), .O(gate179inter9));
  nand2 gate2447(.a(s_271), .b(gate179inter3), .O(gate179inter10));
  nor2  gate2448(.a(gate179inter10), .b(gate179inter9), .O(gate179inter11));
  nor2  gate2449(.a(gate179inter11), .b(gate179inter6), .O(gate179inter12));
  nand2 gate2450(.a(gate179inter12), .b(gate179inter1), .O(G596));
nand2 gate180( .a(G507), .b(G561), .O(G597) );
nand2 gate181( .a(G510), .b(G564), .O(G598) );
nand2 gate182( .a(G513), .b(G564), .O(G599) );

  xor2  gate2073(.a(G567), .b(G516), .O(gate183inter0));
  nand2 gate2074(.a(gate183inter0), .b(s_218), .O(gate183inter1));
  and2  gate2075(.a(G567), .b(G516), .O(gate183inter2));
  inv1  gate2076(.a(s_218), .O(gate183inter3));
  inv1  gate2077(.a(s_219), .O(gate183inter4));
  nand2 gate2078(.a(gate183inter4), .b(gate183inter3), .O(gate183inter5));
  nor2  gate2079(.a(gate183inter5), .b(gate183inter2), .O(gate183inter6));
  inv1  gate2080(.a(G516), .O(gate183inter7));
  inv1  gate2081(.a(G567), .O(gate183inter8));
  nand2 gate2082(.a(gate183inter8), .b(gate183inter7), .O(gate183inter9));
  nand2 gate2083(.a(s_219), .b(gate183inter3), .O(gate183inter10));
  nor2  gate2084(.a(gate183inter10), .b(gate183inter9), .O(gate183inter11));
  nor2  gate2085(.a(gate183inter11), .b(gate183inter6), .O(gate183inter12));
  nand2 gate2086(.a(gate183inter12), .b(gate183inter1), .O(G600));

  xor2  gate1639(.a(G567), .b(G519), .O(gate184inter0));
  nand2 gate1640(.a(gate184inter0), .b(s_156), .O(gate184inter1));
  and2  gate1641(.a(G567), .b(G519), .O(gate184inter2));
  inv1  gate1642(.a(s_156), .O(gate184inter3));
  inv1  gate1643(.a(s_157), .O(gate184inter4));
  nand2 gate1644(.a(gate184inter4), .b(gate184inter3), .O(gate184inter5));
  nor2  gate1645(.a(gate184inter5), .b(gate184inter2), .O(gate184inter6));
  inv1  gate1646(.a(G519), .O(gate184inter7));
  inv1  gate1647(.a(G567), .O(gate184inter8));
  nand2 gate1648(.a(gate184inter8), .b(gate184inter7), .O(gate184inter9));
  nand2 gate1649(.a(s_157), .b(gate184inter3), .O(gate184inter10));
  nor2  gate1650(.a(gate184inter10), .b(gate184inter9), .O(gate184inter11));
  nor2  gate1651(.a(gate184inter11), .b(gate184inter6), .O(gate184inter12));
  nand2 gate1652(.a(gate184inter12), .b(gate184inter1), .O(G601));

  xor2  gate1989(.a(G571), .b(G570), .O(gate185inter0));
  nand2 gate1990(.a(gate185inter0), .b(s_206), .O(gate185inter1));
  and2  gate1991(.a(G571), .b(G570), .O(gate185inter2));
  inv1  gate1992(.a(s_206), .O(gate185inter3));
  inv1  gate1993(.a(s_207), .O(gate185inter4));
  nand2 gate1994(.a(gate185inter4), .b(gate185inter3), .O(gate185inter5));
  nor2  gate1995(.a(gate185inter5), .b(gate185inter2), .O(gate185inter6));
  inv1  gate1996(.a(G570), .O(gate185inter7));
  inv1  gate1997(.a(G571), .O(gate185inter8));
  nand2 gate1998(.a(gate185inter8), .b(gate185inter7), .O(gate185inter9));
  nand2 gate1999(.a(s_207), .b(gate185inter3), .O(gate185inter10));
  nor2  gate2000(.a(gate185inter10), .b(gate185inter9), .O(gate185inter11));
  nor2  gate2001(.a(gate185inter11), .b(gate185inter6), .O(gate185inter12));
  nand2 gate2002(.a(gate185inter12), .b(gate185inter1), .O(G602));
nand2 gate186( .a(G572), .b(G573), .O(G607) );

  xor2  gate2381(.a(G575), .b(G574), .O(gate187inter0));
  nand2 gate2382(.a(gate187inter0), .b(s_262), .O(gate187inter1));
  and2  gate2383(.a(G575), .b(G574), .O(gate187inter2));
  inv1  gate2384(.a(s_262), .O(gate187inter3));
  inv1  gate2385(.a(s_263), .O(gate187inter4));
  nand2 gate2386(.a(gate187inter4), .b(gate187inter3), .O(gate187inter5));
  nor2  gate2387(.a(gate187inter5), .b(gate187inter2), .O(gate187inter6));
  inv1  gate2388(.a(G574), .O(gate187inter7));
  inv1  gate2389(.a(G575), .O(gate187inter8));
  nand2 gate2390(.a(gate187inter8), .b(gate187inter7), .O(gate187inter9));
  nand2 gate2391(.a(s_263), .b(gate187inter3), .O(gate187inter10));
  nor2  gate2392(.a(gate187inter10), .b(gate187inter9), .O(gate187inter11));
  nor2  gate2393(.a(gate187inter11), .b(gate187inter6), .O(gate187inter12));
  nand2 gate2394(.a(gate187inter12), .b(gate187inter1), .O(G612));

  xor2  gate995(.a(G577), .b(G576), .O(gate188inter0));
  nand2 gate996(.a(gate188inter0), .b(s_64), .O(gate188inter1));
  and2  gate997(.a(G577), .b(G576), .O(gate188inter2));
  inv1  gate998(.a(s_64), .O(gate188inter3));
  inv1  gate999(.a(s_65), .O(gate188inter4));
  nand2 gate1000(.a(gate188inter4), .b(gate188inter3), .O(gate188inter5));
  nor2  gate1001(.a(gate188inter5), .b(gate188inter2), .O(gate188inter6));
  inv1  gate1002(.a(G576), .O(gate188inter7));
  inv1  gate1003(.a(G577), .O(gate188inter8));
  nand2 gate1004(.a(gate188inter8), .b(gate188inter7), .O(gate188inter9));
  nand2 gate1005(.a(s_65), .b(gate188inter3), .O(gate188inter10));
  nor2  gate1006(.a(gate188inter10), .b(gate188inter9), .O(gate188inter11));
  nor2  gate1007(.a(gate188inter11), .b(gate188inter6), .O(gate188inter12));
  nand2 gate1008(.a(gate188inter12), .b(gate188inter1), .O(G617));
nand2 gate189( .a(G578), .b(G579), .O(G622) );

  xor2  gate561(.a(G581), .b(G580), .O(gate190inter0));
  nand2 gate562(.a(gate190inter0), .b(s_2), .O(gate190inter1));
  and2  gate563(.a(G581), .b(G580), .O(gate190inter2));
  inv1  gate564(.a(s_2), .O(gate190inter3));
  inv1  gate565(.a(s_3), .O(gate190inter4));
  nand2 gate566(.a(gate190inter4), .b(gate190inter3), .O(gate190inter5));
  nor2  gate567(.a(gate190inter5), .b(gate190inter2), .O(gate190inter6));
  inv1  gate568(.a(G580), .O(gate190inter7));
  inv1  gate569(.a(G581), .O(gate190inter8));
  nand2 gate570(.a(gate190inter8), .b(gate190inter7), .O(gate190inter9));
  nand2 gate571(.a(s_3), .b(gate190inter3), .O(gate190inter10));
  nor2  gate572(.a(gate190inter10), .b(gate190inter9), .O(gate190inter11));
  nor2  gate573(.a(gate190inter11), .b(gate190inter6), .O(gate190inter12));
  nand2 gate574(.a(gate190inter12), .b(gate190inter1), .O(G627));
nand2 gate191( .a(G582), .b(G583), .O(G632) );

  xor2  gate2031(.a(G585), .b(G584), .O(gate192inter0));
  nand2 gate2032(.a(gate192inter0), .b(s_212), .O(gate192inter1));
  and2  gate2033(.a(G585), .b(G584), .O(gate192inter2));
  inv1  gate2034(.a(s_212), .O(gate192inter3));
  inv1  gate2035(.a(s_213), .O(gate192inter4));
  nand2 gate2036(.a(gate192inter4), .b(gate192inter3), .O(gate192inter5));
  nor2  gate2037(.a(gate192inter5), .b(gate192inter2), .O(gate192inter6));
  inv1  gate2038(.a(G584), .O(gate192inter7));
  inv1  gate2039(.a(G585), .O(gate192inter8));
  nand2 gate2040(.a(gate192inter8), .b(gate192inter7), .O(gate192inter9));
  nand2 gate2041(.a(s_213), .b(gate192inter3), .O(gate192inter10));
  nor2  gate2042(.a(gate192inter10), .b(gate192inter9), .O(gate192inter11));
  nor2  gate2043(.a(gate192inter11), .b(gate192inter6), .O(gate192inter12));
  nand2 gate2044(.a(gate192inter12), .b(gate192inter1), .O(G637));

  xor2  gate1541(.a(G587), .b(G586), .O(gate193inter0));
  nand2 gate1542(.a(gate193inter0), .b(s_142), .O(gate193inter1));
  and2  gate1543(.a(G587), .b(G586), .O(gate193inter2));
  inv1  gate1544(.a(s_142), .O(gate193inter3));
  inv1  gate1545(.a(s_143), .O(gate193inter4));
  nand2 gate1546(.a(gate193inter4), .b(gate193inter3), .O(gate193inter5));
  nor2  gate1547(.a(gate193inter5), .b(gate193inter2), .O(gate193inter6));
  inv1  gate1548(.a(G586), .O(gate193inter7));
  inv1  gate1549(.a(G587), .O(gate193inter8));
  nand2 gate1550(.a(gate193inter8), .b(gate193inter7), .O(gate193inter9));
  nand2 gate1551(.a(s_143), .b(gate193inter3), .O(gate193inter10));
  nor2  gate1552(.a(gate193inter10), .b(gate193inter9), .O(gate193inter11));
  nor2  gate1553(.a(gate193inter11), .b(gate193inter6), .O(gate193inter12));
  nand2 gate1554(.a(gate193inter12), .b(gate193inter1), .O(G642));

  xor2  gate1247(.a(G589), .b(G588), .O(gate194inter0));
  nand2 gate1248(.a(gate194inter0), .b(s_100), .O(gate194inter1));
  and2  gate1249(.a(G589), .b(G588), .O(gate194inter2));
  inv1  gate1250(.a(s_100), .O(gate194inter3));
  inv1  gate1251(.a(s_101), .O(gate194inter4));
  nand2 gate1252(.a(gate194inter4), .b(gate194inter3), .O(gate194inter5));
  nor2  gate1253(.a(gate194inter5), .b(gate194inter2), .O(gate194inter6));
  inv1  gate1254(.a(G588), .O(gate194inter7));
  inv1  gate1255(.a(G589), .O(gate194inter8));
  nand2 gate1256(.a(gate194inter8), .b(gate194inter7), .O(gate194inter9));
  nand2 gate1257(.a(s_101), .b(gate194inter3), .O(gate194inter10));
  nor2  gate1258(.a(gate194inter10), .b(gate194inter9), .O(gate194inter11));
  nor2  gate1259(.a(gate194inter11), .b(gate194inter6), .O(gate194inter12));
  nand2 gate1260(.a(gate194inter12), .b(gate194inter1), .O(G645));
nand2 gate195( .a(G590), .b(G591), .O(G648) );
nand2 gate196( .a(G592), .b(G593), .O(G651) );

  xor2  gate1233(.a(G595), .b(G594), .O(gate197inter0));
  nand2 gate1234(.a(gate197inter0), .b(s_98), .O(gate197inter1));
  and2  gate1235(.a(G595), .b(G594), .O(gate197inter2));
  inv1  gate1236(.a(s_98), .O(gate197inter3));
  inv1  gate1237(.a(s_99), .O(gate197inter4));
  nand2 gate1238(.a(gate197inter4), .b(gate197inter3), .O(gate197inter5));
  nor2  gate1239(.a(gate197inter5), .b(gate197inter2), .O(gate197inter6));
  inv1  gate1240(.a(G594), .O(gate197inter7));
  inv1  gate1241(.a(G595), .O(gate197inter8));
  nand2 gate1242(.a(gate197inter8), .b(gate197inter7), .O(gate197inter9));
  nand2 gate1243(.a(s_99), .b(gate197inter3), .O(gate197inter10));
  nor2  gate1244(.a(gate197inter10), .b(gate197inter9), .O(gate197inter11));
  nor2  gate1245(.a(gate197inter11), .b(gate197inter6), .O(gate197inter12));
  nand2 gate1246(.a(gate197inter12), .b(gate197inter1), .O(G654));

  xor2  gate1499(.a(G597), .b(G596), .O(gate198inter0));
  nand2 gate1500(.a(gate198inter0), .b(s_136), .O(gate198inter1));
  and2  gate1501(.a(G597), .b(G596), .O(gate198inter2));
  inv1  gate1502(.a(s_136), .O(gate198inter3));
  inv1  gate1503(.a(s_137), .O(gate198inter4));
  nand2 gate1504(.a(gate198inter4), .b(gate198inter3), .O(gate198inter5));
  nor2  gate1505(.a(gate198inter5), .b(gate198inter2), .O(gate198inter6));
  inv1  gate1506(.a(G596), .O(gate198inter7));
  inv1  gate1507(.a(G597), .O(gate198inter8));
  nand2 gate1508(.a(gate198inter8), .b(gate198inter7), .O(gate198inter9));
  nand2 gate1509(.a(s_137), .b(gate198inter3), .O(gate198inter10));
  nor2  gate1510(.a(gate198inter10), .b(gate198inter9), .O(gate198inter11));
  nor2  gate1511(.a(gate198inter11), .b(gate198inter6), .O(gate198inter12));
  nand2 gate1512(.a(gate198inter12), .b(gate198inter1), .O(G657));
nand2 gate199( .a(G598), .b(G599), .O(G660) );
nand2 gate200( .a(G600), .b(G601), .O(G663) );

  xor2  gate1331(.a(G607), .b(G602), .O(gate201inter0));
  nand2 gate1332(.a(gate201inter0), .b(s_112), .O(gate201inter1));
  and2  gate1333(.a(G607), .b(G602), .O(gate201inter2));
  inv1  gate1334(.a(s_112), .O(gate201inter3));
  inv1  gate1335(.a(s_113), .O(gate201inter4));
  nand2 gate1336(.a(gate201inter4), .b(gate201inter3), .O(gate201inter5));
  nor2  gate1337(.a(gate201inter5), .b(gate201inter2), .O(gate201inter6));
  inv1  gate1338(.a(G602), .O(gate201inter7));
  inv1  gate1339(.a(G607), .O(gate201inter8));
  nand2 gate1340(.a(gate201inter8), .b(gate201inter7), .O(gate201inter9));
  nand2 gate1341(.a(s_113), .b(gate201inter3), .O(gate201inter10));
  nor2  gate1342(.a(gate201inter10), .b(gate201inter9), .O(gate201inter11));
  nor2  gate1343(.a(gate201inter11), .b(gate201inter6), .O(gate201inter12));
  nand2 gate1344(.a(gate201inter12), .b(gate201inter1), .O(G666));

  xor2  gate2157(.a(G617), .b(G612), .O(gate202inter0));
  nand2 gate2158(.a(gate202inter0), .b(s_230), .O(gate202inter1));
  and2  gate2159(.a(G617), .b(G612), .O(gate202inter2));
  inv1  gate2160(.a(s_230), .O(gate202inter3));
  inv1  gate2161(.a(s_231), .O(gate202inter4));
  nand2 gate2162(.a(gate202inter4), .b(gate202inter3), .O(gate202inter5));
  nor2  gate2163(.a(gate202inter5), .b(gate202inter2), .O(gate202inter6));
  inv1  gate2164(.a(G612), .O(gate202inter7));
  inv1  gate2165(.a(G617), .O(gate202inter8));
  nand2 gate2166(.a(gate202inter8), .b(gate202inter7), .O(gate202inter9));
  nand2 gate2167(.a(s_231), .b(gate202inter3), .O(gate202inter10));
  nor2  gate2168(.a(gate202inter10), .b(gate202inter9), .O(gate202inter11));
  nor2  gate2169(.a(gate202inter11), .b(gate202inter6), .O(gate202inter12));
  nand2 gate2170(.a(gate202inter12), .b(gate202inter1), .O(G669));
nand2 gate203( .a(G602), .b(G612), .O(G672) );
nand2 gate204( .a(G607), .b(G617), .O(G675) );
nand2 gate205( .a(G622), .b(G627), .O(G678) );
nand2 gate206( .a(G632), .b(G637), .O(G681) );
nand2 gate207( .a(G622), .b(G632), .O(G684) );
nand2 gate208( .a(G627), .b(G637), .O(G687) );

  xor2  gate1709(.a(G666), .b(G602), .O(gate209inter0));
  nand2 gate1710(.a(gate209inter0), .b(s_166), .O(gate209inter1));
  and2  gate1711(.a(G666), .b(G602), .O(gate209inter2));
  inv1  gate1712(.a(s_166), .O(gate209inter3));
  inv1  gate1713(.a(s_167), .O(gate209inter4));
  nand2 gate1714(.a(gate209inter4), .b(gate209inter3), .O(gate209inter5));
  nor2  gate1715(.a(gate209inter5), .b(gate209inter2), .O(gate209inter6));
  inv1  gate1716(.a(G602), .O(gate209inter7));
  inv1  gate1717(.a(G666), .O(gate209inter8));
  nand2 gate1718(.a(gate209inter8), .b(gate209inter7), .O(gate209inter9));
  nand2 gate1719(.a(s_167), .b(gate209inter3), .O(gate209inter10));
  nor2  gate1720(.a(gate209inter10), .b(gate209inter9), .O(gate209inter11));
  nor2  gate1721(.a(gate209inter11), .b(gate209inter6), .O(gate209inter12));
  nand2 gate1722(.a(gate209inter12), .b(gate209inter1), .O(G690));
nand2 gate210( .a(G607), .b(G666), .O(G691) );
nand2 gate211( .a(G612), .b(G669), .O(G692) );
nand2 gate212( .a(G617), .b(G669), .O(G693) );

  xor2  gate981(.a(G672), .b(G602), .O(gate213inter0));
  nand2 gate982(.a(gate213inter0), .b(s_62), .O(gate213inter1));
  and2  gate983(.a(G672), .b(G602), .O(gate213inter2));
  inv1  gate984(.a(s_62), .O(gate213inter3));
  inv1  gate985(.a(s_63), .O(gate213inter4));
  nand2 gate986(.a(gate213inter4), .b(gate213inter3), .O(gate213inter5));
  nor2  gate987(.a(gate213inter5), .b(gate213inter2), .O(gate213inter6));
  inv1  gate988(.a(G602), .O(gate213inter7));
  inv1  gate989(.a(G672), .O(gate213inter8));
  nand2 gate990(.a(gate213inter8), .b(gate213inter7), .O(gate213inter9));
  nand2 gate991(.a(s_63), .b(gate213inter3), .O(gate213inter10));
  nor2  gate992(.a(gate213inter10), .b(gate213inter9), .O(gate213inter11));
  nor2  gate993(.a(gate213inter11), .b(gate213inter6), .O(gate213inter12));
  nand2 gate994(.a(gate213inter12), .b(gate213inter1), .O(G694));
nand2 gate214( .a(G612), .b(G672), .O(G695) );

  xor2  gate2339(.a(G675), .b(G607), .O(gate215inter0));
  nand2 gate2340(.a(gate215inter0), .b(s_256), .O(gate215inter1));
  and2  gate2341(.a(G675), .b(G607), .O(gate215inter2));
  inv1  gate2342(.a(s_256), .O(gate215inter3));
  inv1  gate2343(.a(s_257), .O(gate215inter4));
  nand2 gate2344(.a(gate215inter4), .b(gate215inter3), .O(gate215inter5));
  nor2  gate2345(.a(gate215inter5), .b(gate215inter2), .O(gate215inter6));
  inv1  gate2346(.a(G607), .O(gate215inter7));
  inv1  gate2347(.a(G675), .O(gate215inter8));
  nand2 gate2348(.a(gate215inter8), .b(gate215inter7), .O(gate215inter9));
  nand2 gate2349(.a(s_257), .b(gate215inter3), .O(gate215inter10));
  nor2  gate2350(.a(gate215inter10), .b(gate215inter9), .O(gate215inter11));
  nor2  gate2351(.a(gate215inter11), .b(gate215inter6), .O(gate215inter12));
  nand2 gate2352(.a(gate215inter12), .b(gate215inter1), .O(G696));
nand2 gate216( .a(G617), .b(G675), .O(G697) );
nand2 gate217( .a(G622), .b(G678), .O(G698) );
nand2 gate218( .a(G627), .b(G678), .O(G699) );
nand2 gate219( .a(G632), .b(G681), .O(G700) );

  xor2  gate827(.a(G681), .b(G637), .O(gate220inter0));
  nand2 gate828(.a(gate220inter0), .b(s_40), .O(gate220inter1));
  and2  gate829(.a(G681), .b(G637), .O(gate220inter2));
  inv1  gate830(.a(s_40), .O(gate220inter3));
  inv1  gate831(.a(s_41), .O(gate220inter4));
  nand2 gate832(.a(gate220inter4), .b(gate220inter3), .O(gate220inter5));
  nor2  gate833(.a(gate220inter5), .b(gate220inter2), .O(gate220inter6));
  inv1  gate834(.a(G637), .O(gate220inter7));
  inv1  gate835(.a(G681), .O(gate220inter8));
  nand2 gate836(.a(gate220inter8), .b(gate220inter7), .O(gate220inter9));
  nand2 gate837(.a(s_41), .b(gate220inter3), .O(gate220inter10));
  nor2  gate838(.a(gate220inter10), .b(gate220inter9), .O(gate220inter11));
  nor2  gate839(.a(gate220inter11), .b(gate220inter6), .O(gate220inter12));
  nand2 gate840(.a(gate220inter12), .b(gate220inter1), .O(G701));
nand2 gate221( .a(G622), .b(G684), .O(G702) );
nand2 gate222( .a(G632), .b(G684), .O(G703) );
nand2 gate223( .a(G627), .b(G687), .O(G704) );
nand2 gate224( .a(G637), .b(G687), .O(G705) );

  xor2  gate1779(.a(G691), .b(G690), .O(gate225inter0));
  nand2 gate1780(.a(gate225inter0), .b(s_176), .O(gate225inter1));
  and2  gate1781(.a(G691), .b(G690), .O(gate225inter2));
  inv1  gate1782(.a(s_176), .O(gate225inter3));
  inv1  gate1783(.a(s_177), .O(gate225inter4));
  nand2 gate1784(.a(gate225inter4), .b(gate225inter3), .O(gate225inter5));
  nor2  gate1785(.a(gate225inter5), .b(gate225inter2), .O(gate225inter6));
  inv1  gate1786(.a(G690), .O(gate225inter7));
  inv1  gate1787(.a(G691), .O(gate225inter8));
  nand2 gate1788(.a(gate225inter8), .b(gate225inter7), .O(gate225inter9));
  nand2 gate1789(.a(s_177), .b(gate225inter3), .O(gate225inter10));
  nor2  gate1790(.a(gate225inter10), .b(gate225inter9), .O(gate225inter11));
  nor2  gate1791(.a(gate225inter11), .b(gate225inter6), .O(gate225inter12));
  nand2 gate1792(.a(gate225inter12), .b(gate225inter1), .O(G706));
nand2 gate226( .a(G692), .b(G693), .O(G709) );

  xor2  gate1849(.a(G695), .b(G694), .O(gate227inter0));
  nand2 gate1850(.a(gate227inter0), .b(s_186), .O(gate227inter1));
  and2  gate1851(.a(G695), .b(G694), .O(gate227inter2));
  inv1  gate1852(.a(s_186), .O(gate227inter3));
  inv1  gate1853(.a(s_187), .O(gate227inter4));
  nand2 gate1854(.a(gate227inter4), .b(gate227inter3), .O(gate227inter5));
  nor2  gate1855(.a(gate227inter5), .b(gate227inter2), .O(gate227inter6));
  inv1  gate1856(.a(G694), .O(gate227inter7));
  inv1  gate1857(.a(G695), .O(gate227inter8));
  nand2 gate1858(.a(gate227inter8), .b(gate227inter7), .O(gate227inter9));
  nand2 gate1859(.a(s_187), .b(gate227inter3), .O(gate227inter10));
  nor2  gate1860(.a(gate227inter10), .b(gate227inter9), .O(gate227inter11));
  nor2  gate1861(.a(gate227inter11), .b(gate227inter6), .O(gate227inter12));
  nand2 gate1862(.a(gate227inter12), .b(gate227inter1), .O(G712));
nand2 gate228( .a(G696), .b(G697), .O(G715) );

  xor2  gate589(.a(G699), .b(G698), .O(gate229inter0));
  nand2 gate590(.a(gate229inter0), .b(s_6), .O(gate229inter1));
  and2  gate591(.a(G699), .b(G698), .O(gate229inter2));
  inv1  gate592(.a(s_6), .O(gate229inter3));
  inv1  gate593(.a(s_7), .O(gate229inter4));
  nand2 gate594(.a(gate229inter4), .b(gate229inter3), .O(gate229inter5));
  nor2  gate595(.a(gate229inter5), .b(gate229inter2), .O(gate229inter6));
  inv1  gate596(.a(G698), .O(gate229inter7));
  inv1  gate597(.a(G699), .O(gate229inter8));
  nand2 gate598(.a(gate229inter8), .b(gate229inter7), .O(gate229inter9));
  nand2 gate599(.a(s_7), .b(gate229inter3), .O(gate229inter10));
  nor2  gate600(.a(gate229inter10), .b(gate229inter9), .O(gate229inter11));
  nor2  gate601(.a(gate229inter11), .b(gate229inter6), .O(gate229inter12));
  nand2 gate602(.a(gate229inter12), .b(gate229inter1), .O(G718));
nand2 gate230( .a(G700), .b(G701), .O(G721) );
nand2 gate231( .a(G702), .b(G703), .O(G724) );
nand2 gate232( .a(G704), .b(G705), .O(G727) );
nand2 gate233( .a(G242), .b(G718), .O(G730) );
nand2 gate234( .a(G245), .b(G721), .O(G733) );
nand2 gate235( .a(G248), .b(G724), .O(G736) );
nand2 gate236( .a(G251), .b(G727), .O(G739) );

  xor2  gate2227(.a(G706), .b(G254), .O(gate237inter0));
  nand2 gate2228(.a(gate237inter0), .b(s_240), .O(gate237inter1));
  and2  gate2229(.a(G706), .b(G254), .O(gate237inter2));
  inv1  gate2230(.a(s_240), .O(gate237inter3));
  inv1  gate2231(.a(s_241), .O(gate237inter4));
  nand2 gate2232(.a(gate237inter4), .b(gate237inter3), .O(gate237inter5));
  nor2  gate2233(.a(gate237inter5), .b(gate237inter2), .O(gate237inter6));
  inv1  gate2234(.a(G254), .O(gate237inter7));
  inv1  gate2235(.a(G706), .O(gate237inter8));
  nand2 gate2236(.a(gate237inter8), .b(gate237inter7), .O(gate237inter9));
  nand2 gate2237(.a(s_241), .b(gate237inter3), .O(gate237inter10));
  nor2  gate2238(.a(gate237inter10), .b(gate237inter9), .O(gate237inter11));
  nor2  gate2239(.a(gate237inter11), .b(gate237inter6), .O(gate237inter12));
  nand2 gate2240(.a(gate237inter12), .b(gate237inter1), .O(G742));

  xor2  gate911(.a(G709), .b(G257), .O(gate238inter0));
  nand2 gate912(.a(gate238inter0), .b(s_52), .O(gate238inter1));
  and2  gate913(.a(G709), .b(G257), .O(gate238inter2));
  inv1  gate914(.a(s_52), .O(gate238inter3));
  inv1  gate915(.a(s_53), .O(gate238inter4));
  nand2 gate916(.a(gate238inter4), .b(gate238inter3), .O(gate238inter5));
  nor2  gate917(.a(gate238inter5), .b(gate238inter2), .O(gate238inter6));
  inv1  gate918(.a(G257), .O(gate238inter7));
  inv1  gate919(.a(G709), .O(gate238inter8));
  nand2 gate920(.a(gate238inter8), .b(gate238inter7), .O(gate238inter9));
  nand2 gate921(.a(s_53), .b(gate238inter3), .O(gate238inter10));
  nor2  gate922(.a(gate238inter10), .b(gate238inter9), .O(gate238inter11));
  nor2  gate923(.a(gate238inter11), .b(gate238inter6), .O(gate238inter12));
  nand2 gate924(.a(gate238inter12), .b(gate238inter1), .O(G745));

  xor2  gate1975(.a(G712), .b(G260), .O(gate239inter0));
  nand2 gate1976(.a(gate239inter0), .b(s_204), .O(gate239inter1));
  and2  gate1977(.a(G712), .b(G260), .O(gate239inter2));
  inv1  gate1978(.a(s_204), .O(gate239inter3));
  inv1  gate1979(.a(s_205), .O(gate239inter4));
  nand2 gate1980(.a(gate239inter4), .b(gate239inter3), .O(gate239inter5));
  nor2  gate1981(.a(gate239inter5), .b(gate239inter2), .O(gate239inter6));
  inv1  gate1982(.a(G260), .O(gate239inter7));
  inv1  gate1983(.a(G712), .O(gate239inter8));
  nand2 gate1984(.a(gate239inter8), .b(gate239inter7), .O(gate239inter9));
  nand2 gate1985(.a(s_205), .b(gate239inter3), .O(gate239inter10));
  nor2  gate1986(.a(gate239inter10), .b(gate239inter9), .O(gate239inter11));
  nor2  gate1987(.a(gate239inter11), .b(gate239inter6), .O(gate239inter12));
  nand2 gate1988(.a(gate239inter12), .b(gate239inter1), .O(G748));

  xor2  gate2493(.a(G715), .b(G263), .O(gate240inter0));
  nand2 gate2494(.a(gate240inter0), .b(s_278), .O(gate240inter1));
  and2  gate2495(.a(G715), .b(G263), .O(gate240inter2));
  inv1  gate2496(.a(s_278), .O(gate240inter3));
  inv1  gate2497(.a(s_279), .O(gate240inter4));
  nand2 gate2498(.a(gate240inter4), .b(gate240inter3), .O(gate240inter5));
  nor2  gate2499(.a(gate240inter5), .b(gate240inter2), .O(gate240inter6));
  inv1  gate2500(.a(G263), .O(gate240inter7));
  inv1  gate2501(.a(G715), .O(gate240inter8));
  nand2 gate2502(.a(gate240inter8), .b(gate240inter7), .O(gate240inter9));
  nand2 gate2503(.a(s_279), .b(gate240inter3), .O(gate240inter10));
  nor2  gate2504(.a(gate240inter10), .b(gate240inter9), .O(gate240inter11));
  nor2  gate2505(.a(gate240inter11), .b(gate240inter6), .O(gate240inter12));
  nand2 gate2506(.a(gate240inter12), .b(gate240inter1), .O(G751));
nand2 gate241( .a(G242), .b(G730), .O(G754) );
nand2 gate242( .a(G718), .b(G730), .O(G755) );

  xor2  gate799(.a(G733), .b(G245), .O(gate243inter0));
  nand2 gate800(.a(gate243inter0), .b(s_36), .O(gate243inter1));
  and2  gate801(.a(G733), .b(G245), .O(gate243inter2));
  inv1  gate802(.a(s_36), .O(gate243inter3));
  inv1  gate803(.a(s_37), .O(gate243inter4));
  nand2 gate804(.a(gate243inter4), .b(gate243inter3), .O(gate243inter5));
  nor2  gate805(.a(gate243inter5), .b(gate243inter2), .O(gate243inter6));
  inv1  gate806(.a(G245), .O(gate243inter7));
  inv1  gate807(.a(G733), .O(gate243inter8));
  nand2 gate808(.a(gate243inter8), .b(gate243inter7), .O(gate243inter9));
  nand2 gate809(.a(s_37), .b(gate243inter3), .O(gate243inter10));
  nor2  gate810(.a(gate243inter10), .b(gate243inter9), .O(gate243inter11));
  nor2  gate811(.a(gate243inter11), .b(gate243inter6), .O(gate243inter12));
  nand2 gate812(.a(gate243inter12), .b(gate243inter1), .O(G756));

  xor2  gate1681(.a(G733), .b(G721), .O(gate244inter0));
  nand2 gate1682(.a(gate244inter0), .b(s_162), .O(gate244inter1));
  and2  gate1683(.a(G733), .b(G721), .O(gate244inter2));
  inv1  gate1684(.a(s_162), .O(gate244inter3));
  inv1  gate1685(.a(s_163), .O(gate244inter4));
  nand2 gate1686(.a(gate244inter4), .b(gate244inter3), .O(gate244inter5));
  nor2  gate1687(.a(gate244inter5), .b(gate244inter2), .O(gate244inter6));
  inv1  gate1688(.a(G721), .O(gate244inter7));
  inv1  gate1689(.a(G733), .O(gate244inter8));
  nand2 gate1690(.a(gate244inter8), .b(gate244inter7), .O(gate244inter9));
  nand2 gate1691(.a(s_163), .b(gate244inter3), .O(gate244inter10));
  nor2  gate1692(.a(gate244inter10), .b(gate244inter9), .O(gate244inter11));
  nor2  gate1693(.a(gate244inter11), .b(gate244inter6), .O(gate244inter12));
  nand2 gate1694(.a(gate244inter12), .b(gate244inter1), .O(G757));

  xor2  gate1093(.a(G736), .b(G248), .O(gate245inter0));
  nand2 gate1094(.a(gate245inter0), .b(s_78), .O(gate245inter1));
  and2  gate1095(.a(G736), .b(G248), .O(gate245inter2));
  inv1  gate1096(.a(s_78), .O(gate245inter3));
  inv1  gate1097(.a(s_79), .O(gate245inter4));
  nand2 gate1098(.a(gate245inter4), .b(gate245inter3), .O(gate245inter5));
  nor2  gate1099(.a(gate245inter5), .b(gate245inter2), .O(gate245inter6));
  inv1  gate1100(.a(G248), .O(gate245inter7));
  inv1  gate1101(.a(G736), .O(gate245inter8));
  nand2 gate1102(.a(gate245inter8), .b(gate245inter7), .O(gate245inter9));
  nand2 gate1103(.a(s_79), .b(gate245inter3), .O(gate245inter10));
  nor2  gate1104(.a(gate245inter10), .b(gate245inter9), .O(gate245inter11));
  nor2  gate1105(.a(gate245inter11), .b(gate245inter6), .O(gate245inter12));
  nand2 gate1106(.a(gate245inter12), .b(gate245inter1), .O(G758));

  xor2  gate2451(.a(G736), .b(G724), .O(gate246inter0));
  nand2 gate2452(.a(gate246inter0), .b(s_272), .O(gate246inter1));
  and2  gate2453(.a(G736), .b(G724), .O(gate246inter2));
  inv1  gate2454(.a(s_272), .O(gate246inter3));
  inv1  gate2455(.a(s_273), .O(gate246inter4));
  nand2 gate2456(.a(gate246inter4), .b(gate246inter3), .O(gate246inter5));
  nor2  gate2457(.a(gate246inter5), .b(gate246inter2), .O(gate246inter6));
  inv1  gate2458(.a(G724), .O(gate246inter7));
  inv1  gate2459(.a(G736), .O(gate246inter8));
  nand2 gate2460(.a(gate246inter8), .b(gate246inter7), .O(gate246inter9));
  nand2 gate2461(.a(s_273), .b(gate246inter3), .O(gate246inter10));
  nor2  gate2462(.a(gate246inter10), .b(gate246inter9), .O(gate246inter11));
  nor2  gate2463(.a(gate246inter11), .b(gate246inter6), .O(gate246inter12));
  nand2 gate2464(.a(gate246inter12), .b(gate246inter1), .O(G759));

  xor2  gate1513(.a(G739), .b(G251), .O(gate247inter0));
  nand2 gate1514(.a(gate247inter0), .b(s_138), .O(gate247inter1));
  and2  gate1515(.a(G739), .b(G251), .O(gate247inter2));
  inv1  gate1516(.a(s_138), .O(gate247inter3));
  inv1  gate1517(.a(s_139), .O(gate247inter4));
  nand2 gate1518(.a(gate247inter4), .b(gate247inter3), .O(gate247inter5));
  nor2  gate1519(.a(gate247inter5), .b(gate247inter2), .O(gate247inter6));
  inv1  gate1520(.a(G251), .O(gate247inter7));
  inv1  gate1521(.a(G739), .O(gate247inter8));
  nand2 gate1522(.a(gate247inter8), .b(gate247inter7), .O(gate247inter9));
  nand2 gate1523(.a(s_139), .b(gate247inter3), .O(gate247inter10));
  nor2  gate1524(.a(gate247inter10), .b(gate247inter9), .O(gate247inter11));
  nor2  gate1525(.a(gate247inter11), .b(gate247inter6), .O(gate247inter12));
  nand2 gate1526(.a(gate247inter12), .b(gate247inter1), .O(G760));
nand2 gate248( .a(G727), .b(G739), .O(G761) );
nand2 gate249( .a(G254), .b(G742), .O(G762) );

  xor2  gate2535(.a(G742), .b(G706), .O(gate250inter0));
  nand2 gate2536(.a(gate250inter0), .b(s_284), .O(gate250inter1));
  and2  gate2537(.a(G742), .b(G706), .O(gate250inter2));
  inv1  gate2538(.a(s_284), .O(gate250inter3));
  inv1  gate2539(.a(s_285), .O(gate250inter4));
  nand2 gate2540(.a(gate250inter4), .b(gate250inter3), .O(gate250inter5));
  nor2  gate2541(.a(gate250inter5), .b(gate250inter2), .O(gate250inter6));
  inv1  gate2542(.a(G706), .O(gate250inter7));
  inv1  gate2543(.a(G742), .O(gate250inter8));
  nand2 gate2544(.a(gate250inter8), .b(gate250inter7), .O(gate250inter9));
  nand2 gate2545(.a(s_285), .b(gate250inter3), .O(gate250inter10));
  nor2  gate2546(.a(gate250inter10), .b(gate250inter9), .O(gate250inter11));
  nor2  gate2547(.a(gate250inter11), .b(gate250inter6), .O(gate250inter12));
  nand2 gate2548(.a(gate250inter12), .b(gate250inter1), .O(G763));
nand2 gate251( .a(G257), .b(G745), .O(G764) );
nand2 gate252( .a(G709), .b(G745), .O(G765) );

  xor2  gate1737(.a(G748), .b(G260), .O(gate253inter0));
  nand2 gate1738(.a(gate253inter0), .b(s_170), .O(gate253inter1));
  and2  gate1739(.a(G748), .b(G260), .O(gate253inter2));
  inv1  gate1740(.a(s_170), .O(gate253inter3));
  inv1  gate1741(.a(s_171), .O(gate253inter4));
  nand2 gate1742(.a(gate253inter4), .b(gate253inter3), .O(gate253inter5));
  nor2  gate1743(.a(gate253inter5), .b(gate253inter2), .O(gate253inter6));
  inv1  gate1744(.a(G260), .O(gate253inter7));
  inv1  gate1745(.a(G748), .O(gate253inter8));
  nand2 gate1746(.a(gate253inter8), .b(gate253inter7), .O(gate253inter9));
  nand2 gate1747(.a(s_171), .b(gate253inter3), .O(gate253inter10));
  nor2  gate1748(.a(gate253inter10), .b(gate253inter9), .O(gate253inter11));
  nor2  gate1749(.a(gate253inter11), .b(gate253inter6), .O(gate253inter12));
  nand2 gate1750(.a(gate253inter12), .b(gate253inter1), .O(G766));

  xor2  gate1121(.a(G748), .b(G712), .O(gate254inter0));
  nand2 gate1122(.a(gate254inter0), .b(s_82), .O(gate254inter1));
  and2  gate1123(.a(G748), .b(G712), .O(gate254inter2));
  inv1  gate1124(.a(s_82), .O(gate254inter3));
  inv1  gate1125(.a(s_83), .O(gate254inter4));
  nand2 gate1126(.a(gate254inter4), .b(gate254inter3), .O(gate254inter5));
  nor2  gate1127(.a(gate254inter5), .b(gate254inter2), .O(gate254inter6));
  inv1  gate1128(.a(G712), .O(gate254inter7));
  inv1  gate1129(.a(G748), .O(gate254inter8));
  nand2 gate1130(.a(gate254inter8), .b(gate254inter7), .O(gate254inter9));
  nand2 gate1131(.a(s_83), .b(gate254inter3), .O(gate254inter10));
  nor2  gate1132(.a(gate254inter10), .b(gate254inter9), .O(gate254inter11));
  nor2  gate1133(.a(gate254inter11), .b(gate254inter6), .O(gate254inter12));
  nand2 gate1134(.a(gate254inter12), .b(gate254inter1), .O(G767));

  xor2  gate1205(.a(G751), .b(G263), .O(gate255inter0));
  nand2 gate1206(.a(gate255inter0), .b(s_94), .O(gate255inter1));
  and2  gate1207(.a(G751), .b(G263), .O(gate255inter2));
  inv1  gate1208(.a(s_94), .O(gate255inter3));
  inv1  gate1209(.a(s_95), .O(gate255inter4));
  nand2 gate1210(.a(gate255inter4), .b(gate255inter3), .O(gate255inter5));
  nor2  gate1211(.a(gate255inter5), .b(gate255inter2), .O(gate255inter6));
  inv1  gate1212(.a(G263), .O(gate255inter7));
  inv1  gate1213(.a(G751), .O(gate255inter8));
  nand2 gate1214(.a(gate255inter8), .b(gate255inter7), .O(gate255inter9));
  nand2 gate1215(.a(s_95), .b(gate255inter3), .O(gate255inter10));
  nor2  gate1216(.a(gate255inter10), .b(gate255inter9), .O(gate255inter11));
  nor2  gate1217(.a(gate255inter11), .b(gate255inter6), .O(gate255inter12));
  nand2 gate1218(.a(gate255inter12), .b(gate255inter1), .O(G768));
nand2 gate256( .a(G715), .b(G751), .O(G769) );

  xor2  gate1695(.a(G755), .b(G754), .O(gate257inter0));
  nand2 gate1696(.a(gate257inter0), .b(s_164), .O(gate257inter1));
  and2  gate1697(.a(G755), .b(G754), .O(gate257inter2));
  inv1  gate1698(.a(s_164), .O(gate257inter3));
  inv1  gate1699(.a(s_165), .O(gate257inter4));
  nand2 gate1700(.a(gate257inter4), .b(gate257inter3), .O(gate257inter5));
  nor2  gate1701(.a(gate257inter5), .b(gate257inter2), .O(gate257inter6));
  inv1  gate1702(.a(G754), .O(gate257inter7));
  inv1  gate1703(.a(G755), .O(gate257inter8));
  nand2 gate1704(.a(gate257inter8), .b(gate257inter7), .O(gate257inter9));
  nand2 gate1705(.a(s_165), .b(gate257inter3), .O(gate257inter10));
  nor2  gate1706(.a(gate257inter10), .b(gate257inter9), .O(gate257inter11));
  nor2  gate1707(.a(gate257inter11), .b(gate257inter6), .O(gate257inter12));
  nand2 gate1708(.a(gate257inter12), .b(gate257inter1), .O(G770));

  xor2  gate2269(.a(G757), .b(G756), .O(gate258inter0));
  nand2 gate2270(.a(gate258inter0), .b(s_246), .O(gate258inter1));
  and2  gate2271(.a(G757), .b(G756), .O(gate258inter2));
  inv1  gate2272(.a(s_246), .O(gate258inter3));
  inv1  gate2273(.a(s_247), .O(gate258inter4));
  nand2 gate2274(.a(gate258inter4), .b(gate258inter3), .O(gate258inter5));
  nor2  gate2275(.a(gate258inter5), .b(gate258inter2), .O(gate258inter6));
  inv1  gate2276(.a(G756), .O(gate258inter7));
  inv1  gate2277(.a(G757), .O(gate258inter8));
  nand2 gate2278(.a(gate258inter8), .b(gate258inter7), .O(gate258inter9));
  nand2 gate2279(.a(s_247), .b(gate258inter3), .O(gate258inter10));
  nor2  gate2280(.a(gate258inter10), .b(gate258inter9), .O(gate258inter11));
  nor2  gate2281(.a(gate258inter11), .b(gate258inter6), .O(gate258inter12));
  nand2 gate2282(.a(gate258inter12), .b(gate258inter1), .O(G773));

  xor2  gate687(.a(G759), .b(G758), .O(gate259inter0));
  nand2 gate688(.a(gate259inter0), .b(s_20), .O(gate259inter1));
  and2  gate689(.a(G759), .b(G758), .O(gate259inter2));
  inv1  gate690(.a(s_20), .O(gate259inter3));
  inv1  gate691(.a(s_21), .O(gate259inter4));
  nand2 gate692(.a(gate259inter4), .b(gate259inter3), .O(gate259inter5));
  nor2  gate693(.a(gate259inter5), .b(gate259inter2), .O(gate259inter6));
  inv1  gate694(.a(G758), .O(gate259inter7));
  inv1  gate695(.a(G759), .O(gate259inter8));
  nand2 gate696(.a(gate259inter8), .b(gate259inter7), .O(gate259inter9));
  nand2 gate697(.a(s_21), .b(gate259inter3), .O(gate259inter10));
  nor2  gate698(.a(gate259inter10), .b(gate259inter9), .O(gate259inter11));
  nor2  gate699(.a(gate259inter11), .b(gate259inter6), .O(gate259inter12));
  nand2 gate700(.a(gate259inter12), .b(gate259inter1), .O(G776));
nand2 gate260( .a(G760), .b(G761), .O(G779) );

  xor2  gate869(.a(G763), .b(G762), .O(gate261inter0));
  nand2 gate870(.a(gate261inter0), .b(s_46), .O(gate261inter1));
  and2  gate871(.a(G763), .b(G762), .O(gate261inter2));
  inv1  gate872(.a(s_46), .O(gate261inter3));
  inv1  gate873(.a(s_47), .O(gate261inter4));
  nand2 gate874(.a(gate261inter4), .b(gate261inter3), .O(gate261inter5));
  nor2  gate875(.a(gate261inter5), .b(gate261inter2), .O(gate261inter6));
  inv1  gate876(.a(G762), .O(gate261inter7));
  inv1  gate877(.a(G763), .O(gate261inter8));
  nand2 gate878(.a(gate261inter8), .b(gate261inter7), .O(gate261inter9));
  nand2 gate879(.a(s_47), .b(gate261inter3), .O(gate261inter10));
  nor2  gate880(.a(gate261inter10), .b(gate261inter9), .O(gate261inter11));
  nor2  gate881(.a(gate261inter11), .b(gate261inter6), .O(gate261inter12));
  nand2 gate882(.a(gate261inter12), .b(gate261inter1), .O(G782));

  xor2  gate2409(.a(G765), .b(G764), .O(gate262inter0));
  nand2 gate2410(.a(gate262inter0), .b(s_266), .O(gate262inter1));
  and2  gate2411(.a(G765), .b(G764), .O(gate262inter2));
  inv1  gate2412(.a(s_266), .O(gate262inter3));
  inv1  gate2413(.a(s_267), .O(gate262inter4));
  nand2 gate2414(.a(gate262inter4), .b(gate262inter3), .O(gate262inter5));
  nor2  gate2415(.a(gate262inter5), .b(gate262inter2), .O(gate262inter6));
  inv1  gate2416(.a(G764), .O(gate262inter7));
  inv1  gate2417(.a(G765), .O(gate262inter8));
  nand2 gate2418(.a(gate262inter8), .b(gate262inter7), .O(gate262inter9));
  nand2 gate2419(.a(s_267), .b(gate262inter3), .O(gate262inter10));
  nor2  gate2420(.a(gate262inter10), .b(gate262inter9), .O(gate262inter11));
  nor2  gate2421(.a(gate262inter11), .b(gate262inter6), .O(gate262inter12));
  nand2 gate2422(.a(gate262inter12), .b(gate262inter1), .O(G785));

  xor2  gate2255(.a(G767), .b(G766), .O(gate263inter0));
  nand2 gate2256(.a(gate263inter0), .b(s_244), .O(gate263inter1));
  and2  gate2257(.a(G767), .b(G766), .O(gate263inter2));
  inv1  gate2258(.a(s_244), .O(gate263inter3));
  inv1  gate2259(.a(s_245), .O(gate263inter4));
  nand2 gate2260(.a(gate263inter4), .b(gate263inter3), .O(gate263inter5));
  nor2  gate2261(.a(gate263inter5), .b(gate263inter2), .O(gate263inter6));
  inv1  gate2262(.a(G766), .O(gate263inter7));
  inv1  gate2263(.a(G767), .O(gate263inter8));
  nand2 gate2264(.a(gate263inter8), .b(gate263inter7), .O(gate263inter9));
  nand2 gate2265(.a(s_245), .b(gate263inter3), .O(gate263inter10));
  nor2  gate2266(.a(gate263inter10), .b(gate263inter9), .O(gate263inter11));
  nor2  gate2267(.a(gate263inter11), .b(gate263inter6), .O(gate263inter12));
  nand2 gate2268(.a(gate263inter12), .b(gate263inter1), .O(G788));
nand2 gate264( .a(G768), .b(G769), .O(G791) );
nand2 gate265( .a(G642), .b(G770), .O(G794) );
nand2 gate266( .a(G645), .b(G773), .O(G797) );
nand2 gate267( .a(G648), .b(G776), .O(G800) );

  xor2  gate1527(.a(G779), .b(G651), .O(gate268inter0));
  nand2 gate1528(.a(gate268inter0), .b(s_140), .O(gate268inter1));
  and2  gate1529(.a(G779), .b(G651), .O(gate268inter2));
  inv1  gate1530(.a(s_140), .O(gate268inter3));
  inv1  gate1531(.a(s_141), .O(gate268inter4));
  nand2 gate1532(.a(gate268inter4), .b(gate268inter3), .O(gate268inter5));
  nor2  gate1533(.a(gate268inter5), .b(gate268inter2), .O(gate268inter6));
  inv1  gate1534(.a(G651), .O(gate268inter7));
  inv1  gate1535(.a(G779), .O(gate268inter8));
  nand2 gate1536(.a(gate268inter8), .b(gate268inter7), .O(gate268inter9));
  nand2 gate1537(.a(s_141), .b(gate268inter3), .O(gate268inter10));
  nor2  gate1538(.a(gate268inter10), .b(gate268inter9), .O(gate268inter11));
  nor2  gate1539(.a(gate268inter11), .b(gate268inter6), .O(gate268inter12));
  nand2 gate1540(.a(gate268inter12), .b(gate268inter1), .O(G803));
nand2 gate269( .a(G654), .b(G782), .O(G806) );

  xor2  gate2171(.a(G785), .b(G657), .O(gate270inter0));
  nand2 gate2172(.a(gate270inter0), .b(s_232), .O(gate270inter1));
  and2  gate2173(.a(G785), .b(G657), .O(gate270inter2));
  inv1  gate2174(.a(s_232), .O(gate270inter3));
  inv1  gate2175(.a(s_233), .O(gate270inter4));
  nand2 gate2176(.a(gate270inter4), .b(gate270inter3), .O(gate270inter5));
  nor2  gate2177(.a(gate270inter5), .b(gate270inter2), .O(gate270inter6));
  inv1  gate2178(.a(G657), .O(gate270inter7));
  inv1  gate2179(.a(G785), .O(gate270inter8));
  nand2 gate2180(.a(gate270inter8), .b(gate270inter7), .O(gate270inter9));
  nand2 gate2181(.a(s_233), .b(gate270inter3), .O(gate270inter10));
  nor2  gate2182(.a(gate270inter10), .b(gate270inter9), .O(gate270inter11));
  nor2  gate2183(.a(gate270inter11), .b(gate270inter6), .O(gate270inter12));
  nand2 gate2184(.a(gate270inter12), .b(gate270inter1), .O(G809));
nand2 gate271( .a(G660), .b(G788), .O(G812) );
nand2 gate272( .a(G663), .b(G791), .O(G815) );
nand2 gate273( .a(G642), .b(G794), .O(G818) );

  xor2  gate1667(.a(G794), .b(G770), .O(gate274inter0));
  nand2 gate1668(.a(gate274inter0), .b(s_160), .O(gate274inter1));
  and2  gate1669(.a(G794), .b(G770), .O(gate274inter2));
  inv1  gate1670(.a(s_160), .O(gate274inter3));
  inv1  gate1671(.a(s_161), .O(gate274inter4));
  nand2 gate1672(.a(gate274inter4), .b(gate274inter3), .O(gate274inter5));
  nor2  gate1673(.a(gate274inter5), .b(gate274inter2), .O(gate274inter6));
  inv1  gate1674(.a(G770), .O(gate274inter7));
  inv1  gate1675(.a(G794), .O(gate274inter8));
  nand2 gate1676(.a(gate274inter8), .b(gate274inter7), .O(gate274inter9));
  nand2 gate1677(.a(s_161), .b(gate274inter3), .O(gate274inter10));
  nor2  gate1678(.a(gate274inter10), .b(gate274inter9), .O(gate274inter11));
  nor2  gate1679(.a(gate274inter11), .b(gate274inter6), .O(gate274inter12));
  nand2 gate1680(.a(gate274inter12), .b(gate274inter1), .O(G819));
nand2 gate275( .a(G645), .b(G797), .O(G820) );
nand2 gate276( .a(G773), .b(G797), .O(G821) );

  xor2  gate925(.a(G800), .b(G648), .O(gate277inter0));
  nand2 gate926(.a(gate277inter0), .b(s_54), .O(gate277inter1));
  and2  gate927(.a(G800), .b(G648), .O(gate277inter2));
  inv1  gate928(.a(s_54), .O(gate277inter3));
  inv1  gate929(.a(s_55), .O(gate277inter4));
  nand2 gate930(.a(gate277inter4), .b(gate277inter3), .O(gate277inter5));
  nor2  gate931(.a(gate277inter5), .b(gate277inter2), .O(gate277inter6));
  inv1  gate932(.a(G648), .O(gate277inter7));
  inv1  gate933(.a(G800), .O(gate277inter8));
  nand2 gate934(.a(gate277inter8), .b(gate277inter7), .O(gate277inter9));
  nand2 gate935(.a(s_55), .b(gate277inter3), .O(gate277inter10));
  nor2  gate936(.a(gate277inter10), .b(gate277inter9), .O(gate277inter11));
  nor2  gate937(.a(gate277inter11), .b(gate277inter6), .O(gate277inter12));
  nand2 gate938(.a(gate277inter12), .b(gate277inter1), .O(G822));

  xor2  gate1373(.a(G800), .b(G776), .O(gate278inter0));
  nand2 gate1374(.a(gate278inter0), .b(s_118), .O(gate278inter1));
  and2  gate1375(.a(G800), .b(G776), .O(gate278inter2));
  inv1  gate1376(.a(s_118), .O(gate278inter3));
  inv1  gate1377(.a(s_119), .O(gate278inter4));
  nand2 gate1378(.a(gate278inter4), .b(gate278inter3), .O(gate278inter5));
  nor2  gate1379(.a(gate278inter5), .b(gate278inter2), .O(gate278inter6));
  inv1  gate1380(.a(G776), .O(gate278inter7));
  inv1  gate1381(.a(G800), .O(gate278inter8));
  nand2 gate1382(.a(gate278inter8), .b(gate278inter7), .O(gate278inter9));
  nand2 gate1383(.a(s_119), .b(gate278inter3), .O(gate278inter10));
  nor2  gate1384(.a(gate278inter10), .b(gate278inter9), .O(gate278inter11));
  nor2  gate1385(.a(gate278inter11), .b(gate278inter6), .O(gate278inter12));
  nand2 gate1386(.a(gate278inter12), .b(gate278inter1), .O(G823));
nand2 gate279( .a(G651), .b(G803), .O(G824) );

  xor2  gate2353(.a(G803), .b(G779), .O(gate280inter0));
  nand2 gate2354(.a(gate280inter0), .b(s_258), .O(gate280inter1));
  and2  gate2355(.a(G803), .b(G779), .O(gate280inter2));
  inv1  gate2356(.a(s_258), .O(gate280inter3));
  inv1  gate2357(.a(s_259), .O(gate280inter4));
  nand2 gate2358(.a(gate280inter4), .b(gate280inter3), .O(gate280inter5));
  nor2  gate2359(.a(gate280inter5), .b(gate280inter2), .O(gate280inter6));
  inv1  gate2360(.a(G779), .O(gate280inter7));
  inv1  gate2361(.a(G803), .O(gate280inter8));
  nand2 gate2362(.a(gate280inter8), .b(gate280inter7), .O(gate280inter9));
  nand2 gate2363(.a(s_259), .b(gate280inter3), .O(gate280inter10));
  nor2  gate2364(.a(gate280inter10), .b(gate280inter9), .O(gate280inter11));
  nor2  gate2365(.a(gate280inter11), .b(gate280inter6), .O(gate280inter12));
  nand2 gate2366(.a(gate280inter12), .b(gate280inter1), .O(G825));
nand2 gate281( .a(G654), .b(G806), .O(G826) );
nand2 gate282( .a(G782), .b(G806), .O(G827) );
nand2 gate283( .a(G657), .b(G809), .O(G828) );

  xor2  gate2311(.a(G809), .b(G785), .O(gate284inter0));
  nand2 gate2312(.a(gate284inter0), .b(s_252), .O(gate284inter1));
  and2  gate2313(.a(G809), .b(G785), .O(gate284inter2));
  inv1  gate2314(.a(s_252), .O(gate284inter3));
  inv1  gate2315(.a(s_253), .O(gate284inter4));
  nand2 gate2316(.a(gate284inter4), .b(gate284inter3), .O(gate284inter5));
  nor2  gate2317(.a(gate284inter5), .b(gate284inter2), .O(gate284inter6));
  inv1  gate2318(.a(G785), .O(gate284inter7));
  inv1  gate2319(.a(G809), .O(gate284inter8));
  nand2 gate2320(.a(gate284inter8), .b(gate284inter7), .O(gate284inter9));
  nand2 gate2321(.a(s_253), .b(gate284inter3), .O(gate284inter10));
  nor2  gate2322(.a(gate284inter10), .b(gate284inter9), .O(gate284inter11));
  nor2  gate2323(.a(gate284inter11), .b(gate284inter6), .O(gate284inter12));
  nand2 gate2324(.a(gate284inter12), .b(gate284inter1), .O(G829));

  xor2  gate2325(.a(G812), .b(G660), .O(gate285inter0));
  nand2 gate2326(.a(gate285inter0), .b(s_254), .O(gate285inter1));
  and2  gate2327(.a(G812), .b(G660), .O(gate285inter2));
  inv1  gate2328(.a(s_254), .O(gate285inter3));
  inv1  gate2329(.a(s_255), .O(gate285inter4));
  nand2 gate2330(.a(gate285inter4), .b(gate285inter3), .O(gate285inter5));
  nor2  gate2331(.a(gate285inter5), .b(gate285inter2), .O(gate285inter6));
  inv1  gate2332(.a(G660), .O(gate285inter7));
  inv1  gate2333(.a(G812), .O(gate285inter8));
  nand2 gate2334(.a(gate285inter8), .b(gate285inter7), .O(gate285inter9));
  nand2 gate2335(.a(s_255), .b(gate285inter3), .O(gate285inter10));
  nor2  gate2336(.a(gate285inter10), .b(gate285inter9), .O(gate285inter11));
  nor2  gate2337(.a(gate285inter11), .b(gate285inter6), .O(gate285inter12));
  nand2 gate2338(.a(gate285inter12), .b(gate285inter1), .O(G830));
nand2 gate286( .a(G788), .b(G812), .O(G831) );
nand2 gate287( .a(G663), .b(G815), .O(G832) );

  xor2  gate2717(.a(G815), .b(G791), .O(gate288inter0));
  nand2 gate2718(.a(gate288inter0), .b(s_310), .O(gate288inter1));
  and2  gate2719(.a(G815), .b(G791), .O(gate288inter2));
  inv1  gate2720(.a(s_310), .O(gate288inter3));
  inv1  gate2721(.a(s_311), .O(gate288inter4));
  nand2 gate2722(.a(gate288inter4), .b(gate288inter3), .O(gate288inter5));
  nor2  gate2723(.a(gate288inter5), .b(gate288inter2), .O(gate288inter6));
  inv1  gate2724(.a(G791), .O(gate288inter7));
  inv1  gate2725(.a(G815), .O(gate288inter8));
  nand2 gate2726(.a(gate288inter8), .b(gate288inter7), .O(gate288inter9));
  nand2 gate2727(.a(s_311), .b(gate288inter3), .O(gate288inter10));
  nor2  gate2728(.a(gate288inter10), .b(gate288inter9), .O(gate288inter11));
  nor2  gate2729(.a(gate288inter11), .b(gate288inter6), .O(gate288inter12));
  nand2 gate2730(.a(gate288inter12), .b(gate288inter1), .O(G833));
nand2 gate289( .a(G818), .b(G819), .O(G834) );
nand2 gate290( .a(G820), .b(G821), .O(G847) );
nand2 gate291( .a(G822), .b(G823), .O(G860) );
nand2 gate292( .a(G824), .b(G825), .O(G873) );

  xor2  gate2241(.a(G829), .b(G828), .O(gate293inter0));
  nand2 gate2242(.a(gate293inter0), .b(s_242), .O(gate293inter1));
  and2  gate2243(.a(G829), .b(G828), .O(gate293inter2));
  inv1  gate2244(.a(s_242), .O(gate293inter3));
  inv1  gate2245(.a(s_243), .O(gate293inter4));
  nand2 gate2246(.a(gate293inter4), .b(gate293inter3), .O(gate293inter5));
  nor2  gate2247(.a(gate293inter5), .b(gate293inter2), .O(gate293inter6));
  inv1  gate2248(.a(G828), .O(gate293inter7));
  inv1  gate2249(.a(G829), .O(gate293inter8));
  nand2 gate2250(.a(gate293inter8), .b(gate293inter7), .O(gate293inter9));
  nand2 gate2251(.a(s_243), .b(gate293inter3), .O(gate293inter10));
  nor2  gate2252(.a(gate293inter10), .b(gate293inter9), .O(gate293inter11));
  nor2  gate2253(.a(gate293inter11), .b(gate293inter6), .O(gate293inter12));
  nand2 gate2254(.a(gate293inter12), .b(gate293inter1), .O(G886));
nand2 gate294( .a(G832), .b(G833), .O(G899) );

  xor2  gate883(.a(G831), .b(G830), .O(gate295inter0));
  nand2 gate884(.a(gate295inter0), .b(s_48), .O(gate295inter1));
  and2  gate885(.a(G831), .b(G830), .O(gate295inter2));
  inv1  gate886(.a(s_48), .O(gate295inter3));
  inv1  gate887(.a(s_49), .O(gate295inter4));
  nand2 gate888(.a(gate295inter4), .b(gate295inter3), .O(gate295inter5));
  nor2  gate889(.a(gate295inter5), .b(gate295inter2), .O(gate295inter6));
  inv1  gate890(.a(G830), .O(gate295inter7));
  inv1  gate891(.a(G831), .O(gate295inter8));
  nand2 gate892(.a(gate295inter8), .b(gate295inter7), .O(gate295inter9));
  nand2 gate893(.a(s_49), .b(gate295inter3), .O(gate295inter10));
  nor2  gate894(.a(gate295inter10), .b(gate295inter9), .O(gate295inter11));
  nor2  gate895(.a(gate295inter11), .b(gate295inter6), .O(gate295inter12));
  nand2 gate896(.a(gate295inter12), .b(gate295inter1), .O(G912));

  xor2  gate2003(.a(G827), .b(G826), .O(gate296inter0));
  nand2 gate2004(.a(gate296inter0), .b(s_208), .O(gate296inter1));
  and2  gate2005(.a(G827), .b(G826), .O(gate296inter2));
  inv1  gate2006(.a(s_208), .O(gate296inter3));
  inv1  gate2007(.a(s_209), .O(gate296inter4));
  nand2 gate2008(.a(gate296inter4), .b(gate296inter3), .O(gate296inter5));
  nor2  gate2009(.a(gate296inter5), .b(gate296inter2), .O(gate296inter6));
  inv1  gate2010(.a(G826), .O(gate296inter7));
  inv1  gate2011(.a(G827), .O(gate296inter8));
  nand2 gate2012(.a(gate296inter8), .b(gate296inter7), .O(gate296inter9));
  nand2 gate2013(.a(s_209), .b(gate296inter3), .O(gate296inter10));
  nor2  gate2014(.a(gate296inter10), .b(gate296inter9), .O(gate296inter11));
  nor2  gate2015(.a(gate296inter11), .b(gate296inter6), .O(gate296inter12));
  nand2 gate2016(.a(gate296inter12), .b(gate296inter1), .O(G925));
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );

  xor2  gate1961(.a(G1036), .b(G1), .O(gate387inter0));
  nand2 gate1962(.a(gate387inter0), .b(s_202), .O(gate387inter1));
  and2  gate1963(.a(G1036), .b(G1), .O(gate387inter2));
  inv1  gate1964(.a(s_202), .O(gate387inter3));
  inv1  gate1965(.a(s_203), .O(gate387inter4));
  nand2 gate1966(.a(gate387inter4), .b(gate387inter3), .O(gate387inter5));
  nor2  gate1967(.a(gate387inter5), .b(gate387inter2), .O(gate387inter6));
  inv1  gate1968(.a(G1), .O(gate387inter7));
  inv1  gate1969(.a(G1036), .O(gate387inter8));
  nand2 gate1970(.a(gate387inter8), .b(gate387inter7), .O(gate387inter9));
  nand2 gate1971(.a(s_203), .b(gate387inter3), .O(gate387inter10));
  nor2  gate1972(.a(gate387inter10), .b(gate387inter9), .O(gate387inter11));
  nor2  gate1973(.a(gate387inter11), .b(gate387inter6), .O(gate387inter12));
  nand2 gate1974(.a(gate387inter12), .b(gate387inter1), .O(G1132));
nand2 gate388( .a(G2), .b(G1039), .O(G1135) );
nand2 gate389( .a(G3), .b(G1042), .O(G1138) );
nand2 gate390( .a(G4), .b(G1045), .O(G1141) );

  xor2  gate2143(.a(G1048), .b(G5), .O(gate391inter0));
  nand2 gate2144(.a(gate391inter0), .b(s_228), .O(gate391inter1));
  and2  gate2145(.a(G1048), .b(G5), .O(gate391inter2));
  inv1  gate2146(.a(s_228), .O(gate391inter3));
  inv1  gate2147(.a(s_229), .O(gate391inter4));
  nand2 gate2148(.a(gate391inter4), .b(gate391inter3), .O(gate391inter5));
  nor2  gate2149(.a(gate391inter5), .b(gate391inter2), .O(gate391inter6));
  inv1  gate2150(.a(G5), .O(gate391inter7));
  inv1  gate2151(.a(G1048), .O(gate391inter8));
  nand2 gate2152(.a(gate391inter8), .b(gate391inter7), .O(gate391inter9));
  nand2 gate2153(.a(s_229), .b(gate391inter3), .O(gate391inter10));
  nor2  gate2154(.a(gate391inter10), .b(gate391inter9), .O(gate391inter11));
  nor2  gate2155(.a(gate391inter11), .b(gate391inter6), .O(gate391inter12));
  nand2 gate2156(.a(gate391inter12), .b(gate391inter1), .O(G1144));

  xor2  gate1429(.a(G1051), .b(G6), .O(gate392inter0));
  nand2 gate1430(.a(gate392inter0), .b(s_126), .O(gate392inter1));
  and2  gate1431(.a(G1051), .b(G6), .O(gate392inter2));
  inv1  gate1432(.a(s_126), .O(gate392inter3));
  inv1  gate1433(.a(s_127), .O(gate392inter4));
  nand2 gate1434(.a(gate392inter4), .b(gate392inter3), .O(gate392inter5));
  nor2  gate1435(.a(gate392inter5), .b(gate392inter2), .O(gate392inter6));
  inv1  gate1436(.a(G6), .O(gate392inter7));
  inv1  gate1437(.a(G1051), .O(gate392inter8));
  nand2 gate1438(.a(gate392inter8), .b(gate392inter7), .O(gate392inter9));
  nand2 gate1439(.a(s_127), .b(gate392inter3), .O(gate392inter10));
  nor2  gate1440(.a(gate392inter10), .b(gate392inter9), .O(gate392inter11));
  nor2  gate1441(.a(gate392inter11), .b(gate392inter6), .O(gate392inter12));
  nand2 gate1442(.a(gate392inter12), .b(gate392inter1), .O(G1147));
nand2 gate393( .a(G7), .b(G1054), .O(G1150) );
nand2 gate394( .a(G8), .b(G1057), .O(G1153) );
nand2 gate395( .a(G9), .b(G1060), .O(G1156) );
nand2 gate396( .a(G10), .b(G1063), .O(G1159) );
nand2 gate397( .a(G11), .b(G1066), .O(G1162) );

  xor2  gate2563(.a(G1069), .b(G12), .O(gate398inter0));
  nand2 gate2564(.a(gate398inter0), .b(s_288), .O(gate398inter1));
  and2  gate2565(.a(G1069), .b(G12), .O(gate398inter2));
  inv1  gate2566(.a(s_288), .O(gate398inter3));
  inv1  gate2567(.a(s_289), .O(gate398inter4));
  nand2 gate2568(.a(gate398inter4), .b(gate398inter3), .O(gate398inter5));
  nor2  gate2569(.a(gate398inter5), .b(gate398inter2), .O(gate398inter6));
  inv1  gate2570(.a(G12), .O(gate398inter7));
  inv1  gate2571(.a(G1069), .O(gate398inter8));
  nand2 gate2572(.a(gate398inter8), .b(gate398inter7), .O(gate398inter9));
  nand2 gate2573(.a(s_289), .b(gate398inter3), .O(gate398inter10));
  nor2  gate2574(.a(gate398inter10), .b(gate398inter9), .O(gate398inter11));
  nor2  gate2575(.a(gate398inter11), .b(gate398inter6), .O(gate398inter12));
  nand2 gate2576(.a(gate398inter12), .b(gate398inter1), .O(G1165));
nand2 gate399( .a(G13), .b(G1072), .O(G1168) );
nand2 gate400( .a(G14), .b(G1075), .O(G1171) );
nand2 gate401( .a(G15), .b(G1078), .O(G1174) );

  xor2  gate2605(.a(G1081), .b(G16), .O(gate402inter0));
  nand2 gate2606(.a(gate402inter0), .b(s_294), .O(gate402inter1));
  and2  gate2607(.a(G1081), .b(G16), .O(gate402inter2));
  inv1  gate2608(.a(s_294), .O(gate402inter3));
  inv1  gate2609(.a(s_295), .O(gate402inter4));
  nand2 gate2610(.a(gate402inter4), .b(gate402inter3), .O(gate402inter5));
  nor2  gate2611(.a(gate402inter5), .b(gate402inter2), .O(gate402inter6));
  inv1  gate2612(.a(G16), .O(gate402inter7));
  inv1  gate2613(.a(G1081), .O(gate402inter8));
  nand2 gate2614(.a(gate402inter8), .b(gate402inter7), .O(gate402inter9));
  nand2 gate2615(.a(s_295), .b(gate402inter3), .O(gate402inter10));
  nor2  gate2616(.a(gate402inter10), .b(gate402inter9), .O(gate402inter11));
  nor2  gate2617(.a(gate402inter11), .b(gate402inter6), .O(gate402inter12));
  nand2 gate2618(.a(gate402inter12), .b(gate402inter1), .O(G1177));

  xor2  gate1107(.a(G1084), .b(G17), .O(gate403inter0));
  nand2 gate1108(.a(gate403inter0), .b(s_80), .O(gate403inter1));
  and2  gate1109(.a(G1084), .b(G17), .O(gate403inter2));
  inv1  gate1110(.a(s_80), .O(gate403inter3));
  inv1  gate1111(.a(s_81), .O(gate403inter4));
  nand2 gate1112(.a(gate403inter4), .b(gate403inter3), .O(gate403inter5));
  nor2  gate1113(.a(gate403inter5), .b(gate403inter2), .O(gate403inter6));
  inv1  gate1114(.a(G17), .O(gate403inter7));
  inv1  gate1115(.a(G1084), .O(gate403inter8));
  nand2 gate1116(.a(gate403inter8), .b(gate403inter7), .O(gate403inter9));
  nand2 gate1117(.a(s_81), .b(gate403inter3), .O(gate403inter10));
  nor2  gate1118(.a(gate403inter10), .b(gate403inter9), .O(gate403inter11));
  nor2  gate1119(.a(gate403inter11), .b(gate403inter6), .O(gate403inter12));
  nand2 gate1120(.a(gate403inter12), .b(gate403inter1), .O(G1180));
nand2 gate404( .a(G18), .b(G1087), .O(G1183) );

  xor2  gate2101(.a(G1090), .b(G19), .O(gate405inter0));
  nand2 gate2102(.a(gate405inter0), .b(s_222), .O(gate405inter1));
  and2  gate2103(.a(G1090), .b(G19), .O(gate405inter2));
  inv1  gate2104(.a(s_222), .O(gate405inter3));
  inv1  gate2105(.a(s_223), .O(gate405inter4));
  nand2 gate2106(.a(gate405inter4), .b(gate405inter3), .O(gate405inter5));
  nor2  gate2107(.a(gate405inter5), .b(gate405inter2), .O(gate405inter6));
  inv1  gate2108(.a(G19), .O(gate405inter7));
  inv1  gate2109(.a(G1090), .O(gate405inter8));
  nand2 gate2110(.a(gate405inter8), .b(gate405inter7), .O(gate405inter9));
  nand2 gate2111(.a(s_223), .b(gate405inter3), .O(gate405inter10));
  nor2  gate2112(.a(gate405inter10), .b(gate405inter9), .O(gate405inter11));
  nor2  gate2113(.a(gate405inter11), .b(gate405inter6), .O(gate405inter12));
  nand2 gate2114(.a(gate405inter12), .b(gate405inter1), .O(G1186));

  xor2  gate1471(.a(G1093), .b(G20), .O(gate406inter0));
  nand2 gate1472(.a(gate406inter0), .b(s_132), .O(gate406inter1));
  and2  gate1473(.a(G1093), .b(G20), .O(gate406inter2));
  inv1  gate1474(.a(s_132), .O(gate406inter3));
  inv1  gate1475(.a(s_133), .O(gate406inter4));
  nand2 gate1476(.a(gate406inter4), .b(gate406inter3), .O(gate406inter5));
  nor2  gate1477(.a(gate406inter5), .b(gate406inter2), .O(gate406inter6));
  inv1  gate1478(.a(G20), .O(gate406inter7));
  inv1  gate1479(.a(G1093), .O(gate406inter8));
  nand2 gate1480(.a(gate406inter8), .b(gate406inter7), .O(gate406inter9));
  nand2 gate1481(.a(s_133), .b(gate406inter3), .O(gate406inter10));
  nor2  gate1482(.a(gate406inter10), .b(gate406inter9), .O(gate406inter11));
  nor2  gate1483(.a(gate406inter11), .b(gate406inter6), .O(gate406inter12));
  nand2 gate1484(.a(gate406inter12), .b(gate406inter1), .O(G1189));

  xor2  gate1219(.a(G1096), .b(G21), .O(gate407inter0));
  nand2 gate1220(.a(gate407inter0), .b(s_96), .O(gate407inter1));
  and2  gate1221(.a(G1096), .b(G21), .O(gate407inter2));
  inv1  gate1222(.a(s_96), .O(gate407inter3));
  inv1  gate1223(.a(s_97), .O(gate407inter4));
  nand2 gate1224(.a(gate407inter4), .b(gate407inter3), .O(gate407inter5));
  nor2  gate1225(.a(gate407inter5), .b(gate407inter2), .O(gate407inter6));
  inv1  gate1226(.a(G21), .O(gate407inter7));
  inv1  gate1227(.a(G1096), .O(gate407inter8));
  nand2 gate1228(.a(gate407inter8), .b(gate407inter7), .O(gate407inter9));
  nand2 gate1229(.a(s_97), .b(gate407inter3), .O(gate407inter10));
  nor2  gate1230(.a(gate407inter10), .b(gate407inter9), .O(gate407inter11));
  nor2  gate1231(.a(gate407inter11), .b(gate407inter6), .O(gate407inter12));
  nand2 gate1232(.a(gate407inter12), .b(gate407inter1), .O(G1192));
nand2 gate408( .a(G22), .b(G1099), .O(G1195) );
nand2 gate409( .a(G23), .b(G1102), .O(G1198) );
nand2 gate410( .a(G24), .b(G1105), .O(G1201) );
nand2 gate411( .a(G25), .b(G1108), .O(G1204) );
nand2 gate412( .a(G26), .b(G1111), .O(G1207) );
nand2 gate413( .a(G27), .b(G1114), .O(G1210) );

  xor2  gate2283(.a(G1117), .b(G28), .O(gate414inter0));
  nand2 gate2284(.a(gate414inter0), .b(s_248), .O(gate414inter1));
  and2  gate2285(.a(G1117), .b(G28), .O(gate414inter2));
  inv1  gate2286(.a(s_248), .O(gate414inter3));
  inv1  gate2287(.a(s_249), .O(gate414inter4));
  nand2 gate2288(.a(gate414inter4), .b(gate414inter3), .O(gate414inter5));
  nor2  gate2289(.a(gate414inter5), .b(gate414inter2), .O(gate414inter6));
  inv1  gate2290(.a(G28), .O(gate414inter7));
  inv1  gate2291(.a(G1117), .O(gate414inter8));
  nand2 gate2292(.a(gate414inter8), .b(gate414inter7), .O(gate414inter9));
  nand2 gate2293(.a(s_249), .b(gate414inter3), .O(gate414inter10));
  nor2  gate2294(.a(gate414inter10), .b(gate414inter9), .O(gate414inter11));
  nor2  gate2295(.a(gate414inter11), .b(gate414inter6), .O(gate414inter12));
  nand2 gate2296(.a(gate414inter12), .b(gate414inter1), .O(G1213));

  xor2  gate659(.a(G1120), .b(G29), .O(gate415inter0));
  nand2 gate660(.a(gate415inter0), .b(s_16), .O(gate415inter1));
  and2  gate661(.a(G1120), .b(G29), .O(gate415inter2));
  inv1  gate662(.a(s_16), .O(gate415inter3));
  inv1  gate663(.a(s_17), .O(gate415inter4));
  nand2 gate664(.a(gate415inter4), .b(gate415inter3), .O(gate415inter5));
  nor2  gate665(.a(gate415inter5), .b(gate415inter2), .O(gate415inter6));
  inv1  gate666(.a(G29), .O(gate415inter7));
  inv1  gate667(.a(G1120), .O(gate415inter8));
  nand2 gate668(.a(gate415inter8), .b(gate415inter7), .O(gate415inter9));
  nand2 gate669(.a(s_17), .b(gate415inter3), .O(gate415inter10));
  nor2  gate670(.a(gate415inter10), .b(gate415inter9), .O(gate415inter11));
  nor2  gate671(.a(gate415inter11), .b(gate415inter6), .O(gate415inter12));
  nand2 gate672(.a(gate415inter12), .b(gate415inter1), .O(G1216));

  xor2  gate757(.a(G1123), .b(G30), .O(gate416inter0));
  nand2 gate758(.a(gate416inter0), .b(s_30), .O(gate416inter1));
  and2  gate759(.a(G1123), .b(G30), .O(gate416inter2));
  inv1  gate760(.a(s_30), .O(gate416inter3));
  inv1  gate761(.a(s_31), .O(gate416inter4));
  nand2 gate762(.a(gate416inter4), .b(gate416inter3), .O(gate416inter5));
  nor2  gate763(.a(gate416inter5), .b(gate416inter2), .O(gate416inter6));
  inv1  gate764(.a(G30), .O(gate416inter7));
  inv1  gate765(.a(G1123), .O(gate416inter8));
  nand2 gate766(.a(gate416inter8), .b(gate416inter7), .O(gate416inter9));
  nand2 gate767(.a(s_31), .b(gate416inter3), .O(gate416inter10));
  nor2  gate768(.a(gate416inter10), .b(gate416inter9), .O(gate416inter11));
  nor2  gate769(.a(gate416inter11), .b(gate416inter6), .O(gate416inter12));
  nand2 gate770(.a(gate416inter12), .b(gate416inter1), .O(G1219));
nand2 gate417( .a(G31), .b(G1126), .O(G1222) );
nand2 gate418( .a(G32), .b(G1129), .O(G1225) );
nand2 gate419( .a(G1), .b(G1132), .O(G1228) );

  xor2  gate1275(.a(G1132), .b(G1036), .O(gate420inter0));
  nand2 gate1276(.a(gate420inter0), .b(s_104), .O(gate420inter1));
  and2  gate1277(.a(G1132), .b(G1036), .O(gate420inter2));
  inv1  gate1278(.a(s_104), .O(gate420inter3));
  inv1  gate1279(.a(s_105), .O(gate420inter4));
  nand2 gate1280(.a(gate420inter4), .b(gate420inter3), .O(gate420inter5));
  nor2  gate1281(.a(gate420inter5), .b(gate420inter2), .O(gate420inter6));
  inv1  gate1282(.a(G1036), .O(gate420inter7));
  inv1  gate1283(.a(G1132), .O(gate420inter8));
  nand2 gate1284(.a(gate420inter8), .b(gate420inter7), .O(gate420inter9));
  nand2 gate1285(.a(s_105), .b(gate420inter3), .O(gate420inter10));
  nor2  gate1286(.a(gate420inter10), .b(gate420inter9), .O(gate420inter11));
  nor2  gate1287(.a(gate420inter11), .b(gate420inter6), .O(gate420inter12));
  nand2 gate1288(.a(gate420inter12), .b(gate420inter1), .O(G1229));
nand2 gate421( .a(G2), .b(G1135), .O(G1230) );
nand2 gate422( .a(G1039), .b(G1135), .O(G1231) );
nand2 gate423( .a(G3), .b(G1138), .O(G1232) );
nand2 gate424( .a(G1042), .b(G1138), .O(G1233) );
nand2 gate425( .a(G4), .b(G1141), .O(G1234) );

  xor2  gate1443(.a(G1141), .b(G1045), .O(gate426inter0));
  nand2 gate1444(.a(gate426inter0), .b(s_128), .O(gate426inter1));
  and2  gate1445(.a(G1141), .b(G1045), .O(gate426inter2));
  inv1  gate1446(.a(s_128), .O(gate426inter3));
  inv1  gate1447(.a(s_129), .O(gate426inter4));
  nand2 gate1448(.a(gate426inter4), .b(gate426inter3), .O(gate426inter5));
  nor2  gate1449(.a(gate426inter5), .b(gate426inter2), .O(gate426inter6));
  inv1  gate1450(.a(G1045), .O(gate426inter7));
  inv1  gate1451(.a(G1141), .O(gate426inter8));
  nand2 gate1452(.a(gate426inter8), .b(gate426inter7), .O(gate426inter9));
  nand2 gate1453(.a(s_129), .b(gate426inter3), .O(gate426inter10));
  nor2  gate1454(.a(gate426inter10), .b(gate426inter9), .O(gate426inter11));
  nor2  gate1455(.a(gate426inter11), .b(gate426inter6), .O(gate426inter12));
  nand2 gate1456(.a(gate426inter12), .b(gate426inter1), .O(G1235));
nand2 gate427( .a(G5), .b(G1144), .O(G1236) );
nand2 gate428( .a(G1048), .b(G1144), .O(G1237) );

  xor2  gate1387(.a(G1147), .b(G6), .O(gate429inter0));
  nand2 gate1388(.a(gate429inter0), .b(s_120), .O(gate429inter1));
  and2  gate1389(.a(G1147), .b(G6), .O(gate429inter2));
  inv1  gate1390(.a(s_120), .O(gate429inter3));
  inv1  gate1391(.a(s_121), .O(gate429inter4));
  nand2 gate1392(.a(gate429inter4), .b(gate429inter3), .O(gate429inter5));
  nor2  gate1393(.a(gate429inter5), .b(gate429inter2), .O(gate429inter6));
  inv1  gate1394(.a(G6), .O(gate429inter7));
  inv1  gate1395(.a(G1147), .O(gate429inter8));
  nand2 gate1396(.a(gate429inter8), .b(gate429inter7), .O(gate429inter9));
  nand2 gate1397(.a(s_121), .b(gate429inter3), .O(gate429inter10));
  nor2  gate1398(.a(gate429inter10), .b(gate429inter9), .O(gate429inter11));
  nor2  gate1399(.a(gate429inter11), .b(gate429inter6), .O(gate429inter12));
  nand2 gate1400(.a(gate429inter12), .b(gate429inter1), .O(G1238));
nand2 gate430( .a(G1051), .b(G1147), .O(G1239) );

  xor2  gate1793(.a(G1150), .b(G7), .O(gate431inter0));
  nand2 gate1794(.a(gate431inter0), .b(s_178), .O(gate431inter1));
  and2  gate1795(.a(G1150), .b(G7), .O(gate431inter2));
  inv1  gate1796(.a(s_178), .O(gate431inter3));
  inv1  gate1797(.a(s_179), .O(gate431inter4));
  nand2 gate1798(.a(gate431inter4), .b(gate431inter3), .O(gate431inter5));
  nor2  gate1799(.a(gate431inter5), .b(gate431inter2), .O(gate431inter6));
  inv1  gate1800(.a(G7), .O(gate431inter7));
  inv1  gate1801(.a(G1150), .O(gate431inter8));
  nand2 gate1802(.a(gate431inter8), .b(gate431inter7), .O(gate431inter9));
  nand2 gate1803(.a(s_179), .b(gate431inter3), .O(gate431inter10));
  nor2  gate1804(.a(gate431inter10), .b(gate431inter9), .O(gate431inter11));
  nor2  gate1805(.a(gate431inter11), .b(gate431inter6), .O(gate431inter12));
  nand2 gate1806(.a(gate431inter12), .b(gate431inter1), .O(G1240));

  xor2  gate2115(.a(G1150), .b(G1054), .O(gate432inter0));
  nand2 gate2116(.a(gate432inter0), .b(s_224), .O(gate432inter1));
  and2  gate2117(.a(G1150), .b(G1054), .O(gate432inter2));
  inv1  gate2118(.a(s_224), .O(gate432inter3));
  inv1  gate2119(.a(s_225), .O(gate432inter4));
  nand2 gate2120(.a(gate432inter4), .b(gate432inter3), .O(gate432inter5));
  nor2  gate2121(.a(gate432inter5), .b(gate432inter2), .O(gate432inter6));
  inv1  gate2122(.a(G1054), .O(gate432inter7));
  inv1  gate2123(.a(G1150), .O(gate432inter8));
  nand2 gate2124(.a(gate432inter8), .b(gate432inter7), .O(gate432inter9));
  nand2 gate2125(.a(s_225), .b(gate432inter3), .O(gate432inter10));
  nor2  gate2126(.a(gate432inter10), .b(gate432inter9), .O(gate432inter11));
  nor2  gate2127(.a(gate432inter11), .b(gate432inter6), .O(gate432inter12));
  nand2 gate2128(.a(gate432inter12), .b(gate432inter1), .O(G1241));

  xor2  gate2367(.a(G1153), .b(G8), .O(gate433inter0));
  nand2 gate2368(.a(gate433inter0), .b(s_260), .O(gate433inter1));
  and2  gate2369(.a(G1153), .b(G8), .O(gate433inter2));
  inv1  gate2370(.a(s_260), .O(gate433inter3));
  inv1  gate2371(.a(s_261), .O(gate433inter4));
  nand2 gate2372(.a(gate433inter4), .b(gate433inter3), .O(gate433inter5));
  nor2  gate2373(.a(gate433inter5), .b(gate433inter2), .O(gate433inter6));
  inv1  gate2374(.a(G8), .O(gate433inter7));
  inv1  gate2375(.a(G1153), .O(gate433inter8));
  nand2 gate2376(.a(gate433inter8), .b(gate433inter7), .O(gate433inter9));
  nand2 gate2377(.a(s_261), .b(gate433inter3), .O(gate433inter10));
  nor2  gate2378(.a(gate433inter10), .b(gate433inter9), .O(gate433inter11));
  nor2  gate2379(.a(gate433inter11), .b(gate433inter6), .O(gate433inter12));
  nand2 gate2380(.a(gate433inter12), .b(gate433inter1), .O(G1242));
nand2 gate434( .a(G1057), .b(G1153), .O(G1243) );
nand2 gate435( .a(G9), .b(G1156), .O(G1244) );
nand2 gate436( .a(G1060), .b(G1156), .O(G1245) );

  xor2  gate1163(.a(G1159), .b(G10), .O(gate437inter0));
  nand2 gate1164(.a(gate437inter0), .b(s_88), .O(gate437inter1));
  and2  gate1165(.a(G1159), .b(G10), .O(gate437inter2));
  inv1  gate1166(.a(s_88), .O(gate437inter3));
  inv1  gate1167(.a(s_89), .O(gate437inter4));
  nand2 gate1168(.a(gate437inter4), .b(gate437inter3), .O(gate437inter5));
  nor2  gate1169(.a(gate437inter5), .b(gate437inter2), .O(gate437inter6));
  inv1  gate1170(.a(G10), .O(gate437inter7));
  inv1  gate1171(.a(G1159), .O(gate437inter8));
  nand2 gate1172(.a(gate437inter8), .b(gate437inter7), .O(gate437inter9));
  nand2 gate1173(.a(s_89), .b(gate437inter3), .O(gate437inter10));
  nor2  gate1174(.a(gate437inter10), .b(gate437inter9), .O(gate437inter11));
  nor2  gate1175(.a(gate437inter11), .b(gate437inter6), .O(gate437inter12));
  nand2 gate1176(.a(gate437inter12), .b(gate437inter1), .O(G1246));
nand2 gate438( .a(G1063), .b(G1159), .O(G1247) );
nand2 gate439( .a(G11), .b(G1162), .O(G1248) );
nand2 gate440( .a(G1066), .b(G1162), .O(G1249) );
nand2 gate441( .a(G12), .b(G1165), .O(G1250) );

  xor2  gate1569(.a(G1165), .b(G1069), .O(gate442inter0));
  nand2 gate1570(.a(gate442inter0), .b(s_146), .O(gate442inter1));
  and2  gate1571(.a(G1165), .b(G1069), .O(gate442inter2));
  inv1  gate1572(.a(s_146), .O(gate442inter3));
  inv1  gate1573(.a(s_147), .O(gate442inter4));
  nand2 gate1574(.a(gate442inter4), .b(gate442inter3), .O(gate442inter5));
  nor2  gate1575(.a(gate442inter5), .b(gate442inter2), .O(gate442inter6));
  inv1  gate1576(.a(G1069), .O(gate442inter7));
  inv1  gate1577(.a(G1165), .O(gate442inter8));
  nand2 gate1578(.a(gate442inter8), .b(gate442inter7), .O(gate442inter9));
  nand2 gate1579(.a(s_147), .b(gate442inter3), .O(gate442inter10));
  nor2  gate1580(.a(gate442inter10), .b(gate442inter9), .O(gate442inter11));
  nor2  gate1581(.a(gate442inter11), .b(gate442inter6), .O(gate442inter12));
  nand2 gate1582(.a(gate442inter12), .b(gate442inter1), .O(G1251));
nand2 gate443( .a(G13), .b(G1168), .O(G1252) );
nand2 gate444( .a(G1072), .b(G1168), .O(G1253) );
nand2 gate445( .a(G14), .b(G1171), .O(G1254) );
nand2 gate446( .a(G1075), .b(G1171), .O(G1255) );
nand2 gate447( .a(G15), .b(G1174), .O(G1256) );

  xor2  gate729(.a(G1174), .b(G1078), .O(gate448inter0));
  nand2 gate730(.a(gate448inter0), .b(s_26), .O(gate448inter1));
  and2  gate731(.a(G1174), .b(G1078), .O(gate448inter2));
  inv1  gate732(.a(s_26), .O(gate448inter3));
  inv1  gate733(.a(s_27), .O(gate448inter4));
  nand2 gate734(.a(gate448inter4), .b(gate448inter3), .O(gate448inter5));
  nor2  gate735(.a(gate448inter5), .b(gate448inter2), .O(gate448inter6));
  inv1  gate736(.a(G1078), .O(gate448inter7));
  inv1  gate737(.a(G1174), .O(gate448inter8));
  nand2 gate738(.a(gate448inter8), .b(gate448inter7), .O(gate448inter9));
  nand2 gate739(.a(s_27), .b(gate448inter3), .O(gate448inter10));
  nor2  gate740(.a(gate448inter10), .b(gate448inter9), .O(gate448inter11));
  nor2  gate741(.a(gate448inter11), .b(gate448inter6), .O(gate448inter12));
  nand2 gate742(.a(gate448inter12), .b(gate448inter1), .O(G1257));

  xor2  gate1863(.a(G1177), .b(G16), .O(gate449inter0));
  nand2 gate1864(.a(gate449inter0), .b(s_188), .O(gate449inter1));
  and2  gate1865(.a(G1177), .b(G16), .O(gate449inter2));
  inv1  gate1866(.a(s_188), .O(gate449inter3));
  inv1  gate1867(.a(s_189), .O(gate449inter4));
  nand2 gate1868(.a(gate449inter4), .b(gate449inter3), .O(gate449inter5));
  nor2  gate1869(.a(gate449inter5), .b(gate449inter2), .O(gate449inter6));
  inv1  gate1870(.a(G16), .O(gate449inter7));
  inv1  gate1871(.a(G1177), .O(gate449inter8));
  nand2 gate1872(.a(gate449inter8), .b(gate449inter7), .O(gate449inter9));
  nand2 gate1873(.a(s_189), .b(gate449inter3), .O(gate449inter10));
  nor2  gate1874(.a(gate449inter10), .b(gate449inter9), .O(gate449inter11));
  nor2  gate1875(.a(gate449inter11), .b(gate449inter6), .O(gate449inter12));
  nand2 gate1876(.a(gate449inter12), .b(gate449inter1), .O(G1258));

  xor2  gate1051(.a(G1177), .b(G1081), .O(gate450inter0));
  nand2 gate1052(.a(gate450inter0), .b(s_72), .O(gate450inter1));
  and2  gate1053(.a(G1177), .b(G1081), .O(gate450inter2));
  inv1  gate1054(.a(s_72), .O(gate450inter3));
  inv1  gate1055(.a(s_73), .O(gate450inter4));
  nand2 gate1056(.a(gate450inter4), .b(gate450inter3), .O(gate450inter5));
  nor2  gate1057(.a(gate450inter5), .b(gate450inter2), .O(gate450inter6));
  inv1  gate1058(.a(G1081), .O(gate450inter7));
  inv1  gate1059(.a(G1177), .O(gate450inter8));
  nand2 gate1060(.a(gate450inter8), .b(gate450inter7), .O(gate450inter9));
  nand2 gate1061(.a(s_73), .b(gate450inter3), .O(gate450inter10));
  nor2  gate1062(.a(gate450inter10), .b(gate450inter9), .O(gate450inter11));
  nor2  gate1063(.a(gate450inter11), .b(gate450inter6), .O(gate450inter12));
  nand2 gate1064(.a(gate450inter12), .b(gate450inter1), .O(G1259));
nand2 gate451( .a(G17), .b(G1180), .O(G1260) );

  xor2  gate603(.a(G1180), .b(G1084), .O(gate452inter0));
  nand2 gate604(.a(gate452inter0), .b(s_8), .O(gate452inter1));
  and2  gate605(.a(G1180), .b(G1084), .O(gate452inter2));
  inv1  gate606(.a(s_8), .O(gate452inter3));
  inv1  gate607(.a(s_9), .O(gate452inter4));
  nand2 gate608(.a(gate452inter4), .b(gate452inter3), .O(gate452inter5));
  nor2  gate609(.a(gate452inter5), .b(gate452inter2), .O(gate452inter6));
  inv1  gate610(.a(G1084), .O(gate452inter7));
  inv1  gate611(.a(G1180), .O(gate452inter8));
  nand2 gate612(.a(gate452inter8), .b(gate452inter7), .O(gate452inter9));
  nand2 gate613(.a(s_9), .b(gate452inter3), .O(gate452inter10));
  nor2  gate614(.a(gate452inter10), .b(gate452inter9), .O(gate452inter11));
  nor2  gate615(.a(gate452inter11), .b(gate452inter6), .O(gate452inter12));
  nand2 gate616(.a(gate452inter12), .b(gate452inter1), .O(G1261));

  xor2  gate1289(.a(G1183), .b(G18), .O(gate453inter0));
  nand2 gate1290(.a(gate453inter0), .b(s_106), .O(gate453inter1));
  and2  gate1291(.a(G1183), .b(G18), .O(gate453inter2));
  inv1  gate1292(.a(s_106), .O(gate453inter3));
  inv1  gate1293(.a(s_107), .O(gate453inter4));
  nand2 gate1294(.a(gate453inter4), .b(gate453inter3), .O(gate453inter5));
  nor2  gate1295(.a(gate453inter5), .b(gate453inter2), .O(gate453inter6));
  inv1  gate1296(.a(G18), .O(gate453inter7));
  inv1  gate1297(.a(G1183), .O(gate453inter8));
  nand2 gate1298(.a(gate453inter8), .b(gate453inter7), .O(gate453inter9));
  nand2 gate1299(.a(s_107), .b(gate453inter3), .O(gate453inter10));
  nor2  gate1300(.a(gate453inter10), .b(gate453inter9), .O(gate453inter11));
  nor2  gate1301(.a(gate453inter11), .b(gate453inter6), .O(gate453inter12));
  nand2 gate1302(.a(gate453inter12), .b(gate453inter1), .O(G1262));
nand2 gate454( .a(G1087), .b(G1183), .O(G1263) );
nand2 gate455( .a(G19), .b(G1186), .O(G1264) );
nand2 gate456( .a(G1090), .b(G1186), .O(G1265) );
nand2 gate457( .a(G20), .b(G1189), .O(G1266) );

  xor2  gate2395(.a(G1189), .b(G1093), .O(gate458inter0));
  nand2 gate2396(.a(gate458inter0), .b(s_264), .O(gate458inter1));
  and2  gate2397(.a(G1189), .b(G1093), .O(gate458inter2));
  inv1  gate2398(.a(s_264), .O(gate458inter3));
  inv1  gate2399(.a(s_265), .O(gate458inter4));
  nand2 gate2400(.a(gate458inter4), .b(gate458inter3), .O(gate458inter5));
  nor2  gate2401(.a(gate458inter5), .b(gate458inter2), .O(gate458inter6));
  inv1  gate2402(.a(G1093), .O(gate458inter7));
  inv1  gate2403(.a(G1189), .O(gate458inter8));
  nand2 gate2404(.a(gate458inter8), .b(gate458inter7), .O(gate458inter9));
  nand2 gate2405(.a(s_265), .b(gate458inter3), .O(gate458inter10));
  nor2  gate2406(.a(gate458inter10), .b(gate458inter9), .O(gate458inter11));
  nor2  gate2407(.a(gate458inter11), .b(gate458inter6), .O(gate458inter12));
  nand2 gate2408(.a(gate458inter12), .b(gate458inter1), .O(G1267));
nand2 gate459( .a(G21), .b(G1192), .O(G1268) );

  xor2  gate897(.a(G1192), .b(G1096), .O(gate460inter0));
  nand2 gate898(.a(gate460inter0), .b(s_50), .O(gate460inter1));
  and2  gate899(.a(G1192), .b(G1096), .O(gate460inter2));
  inv1  gate900(.a(s_50), .O(gate460inter3));
  inv1  gate901(.a(s_51), .O(gate460inter4));
  nand2 gate902(.a(gate460inter4), .b(gate460inter3), .O(gate460inter5));
  nor2  gate903(.a(gate460inter5), .b(gate460inter2), .O(gate460inter6));
  inv1  gate904(.a(G1096), .O(gate460inter7));
  inv1  gate905(.a(G1192), .O(gate460inter8));
  nand2 gate906(.a(gate460inter8), .b(gate460inter7), .O(gate460inter9));
  nand2 gate907(.a(s_51), .b(gate460inter3), .O(gate460inter10));
  nor2  gate908(.a(gate460inter10), .b(gate460inter9), .O(gate460inter11));
  nor2  gate909(.a(gate460inter11), .b(gate460inter6), .O(gate460inter12));
  nand2 gate910(.a(gate460inter12), .b(gate460inter1), .O(G1269));

  xor2  gate2017(.a(G1195), .b(G22), .O(gate461inter0));
  nand2 gate2018(.a(gate461inter0), .b(s_210), .O(gate461inter1));
  and2  gate2019(.a(G1195), .b(G22), .O(gate461inter2));
  inv1  gate2020(.a(s_210), .O(gate461inter3));
  inv1  gate2021(.a(s_211), .O(gate461inter4));
  nand2 gate2022(.a(gate461inter4), .b(gate461inter3), .O(gate461inter5));
  nor2  gate2023(.a(gate461inter5), .b(gate461inter2), .O(gate461inter6));
  inv1  gate2024(.a(G22), .O(gate461inter7));
  inv1  gate2025(.a(G1195), .O(gate461inter8));
  nand2 gate2026(.a(gate461inter8), .b(gate461inter7), .O(gate461inter9));
  nand2 gate2027(.a(s_211), .b(gate461inter3), .O(gate461inter10));
  nor2  gate2028(.a(gate461inter10), .b(gate461inter9), .O(gate461inter11));
  nor2  gate2029(.a(gate461inter11), .b(gate461inter6), .O(gate461inter12));
  nand2 gate2030(.a(gate461inter12), .b(gate461inter1), .O(G1270));

  xor2  gate2213(.a(G1195), .b(G1099), .O(gate462inter0));
  nand2 gate2214(.a(gate462inter0), .b(s_238), .O(gate462inter1));
  and2  gate2215(.a(G1195), .b(G1099), .O(gate462inter2));
  inv1  gate2216(.a(s_238), .O(gate462inter3));
  inv1  gate2217(.a(s_239), .O(gate462inter4));
  nand2 gate2218(.a(gate462inter4), .b(gate462inter3), .O(gate462inter5));
  nor2  gate2219(.a(gate462inter5), .b(gate462inter2), .O(gate462inter6));
  inv1  gate2220(.a(G1099), .O(gate462inter7));
  inv1  gate2221(.a(G1195), .O(gate462inter8));
  nand2 gate2222(.a(gate462inter8), .b(gate462inter7), .O(gate462inter9));
  nand2 gate2223(.a(s_239), .b(gate462inter3), .O(gate462inter10));
  nor2  gate2224(.a(gate462inter10), .b(gate462inter9), .O(gate462inter11));
  nor2  gate2225(.a(gate462inter11), .b(gate462inter6), .O(gate462inter12));
  nand2 gate2226(.a(gate462inter12), .b(gate462inter1), .O(G1271));
nand2 gate463( .a(G23), .b(G1198), .O(G1272) );
nand2 gate464( .a(G1102), .b(G1198), .O(G1273) );

  xor2  gate1653(.a(G1201), .b(G24), .O(gate465inter0));
  nand2 gate1654(.a(gate465inter0), .b(s_158), .O(gate465inter1));
  and2  gate1655(.a(G1201), .b(G24), .O(gate465inter2));
  inv1  gate1656(.a(s_158), .O(gate465inter3));
  inv1  gate1657(.a(s_159), .O(gate465inter4));
  nand2 gate1658(.a(gate465inter4), .b(gate465inter3), .O(gate465inter5));
  nor2  gate1659(.a(gate465inter5), .b(gate465inter2), .O(gate465inter6));
  inv1  gate1660(.a(G24), .O(gate465inter7));
  inv1  gate1661(.a(G1201), .O(gate465inter8));
  nand2 gate1662(.a(gate465inter8), .b(gate465inter7), .O(gate465inter9));
  nand2 gate1663(.a(s_159), .b(gate465inter3), .O(gate465inter10));
  nor2  gate1664(.a(gate465inter10), .b(gate465inter9), .O(gate465inter11));
  nor2  gate1665(.a(gate465inter11), .b(gate465inter6), .O(gate465inter12));
  nand2 gate1666(.a(gate465inter12), .b(gate465inter1), .O(G1274));

  xor2  gate715(.a(G1201), .b(G1105), .O(gate466inter0));
  nand2 gate716(.a(gate466inter0), .b(s_24), .O(gate466inter1));
  and2  gate717(.a(G1201), .b(G1105), .O(gate466inter2));
  inv1  gate718(.a(s_24), .O(gate466inter3));
  inv1  gate719(.a(s_25), .O(gate466inter4));
  nand2 gate720(.a(gate466inter4), .b(gate466inter3), .O(gate466inter5));
  nor2  gate721(.a(gate466inter5), .b(gate466inter2), .O(gate466inter6));
  inv1  gate722(.a(G1105), .O(gate466inter7));
  inv1  gate723(.a(G1201), .O(gate466inter8));
  nand2 gate724(.a(gate466inter8), .b(gate466inter7), .O(gate466inter9));
  nand2 gate725(.a(s_25), .b(gate466inter3), .O(gate466inter10));
  nor2  gate726(.a(gate466inter10), .b(gate466inter9), .O(gate466inter11));
  nor2  gate727(.a(gate466inter11), .b(gate466inter6), .O(gate466inter12));
  nand2 gate728(.a(gate466inter12), .b(gate466inter1), .O(G1275));
nand2 gate467( .a(G25), .b(G1204), .O(G1276) );
nand2 gate468( .a(G1108), .b(G1204), .O(G1277) );
nand2 gate469( .a(G26), .b(G1207), .O(G1278) );
nand2 gate470( .a(G1111), .b(G1207), .O(G1279) );

  xor2  gate1037(.a(G1210), .b(G27), .O(gate471inter0));
  nand2 gate1038(.a(gate471inter0), .b(s_70), .O(gate471inter1));
  and2  gate1039(.a(G1210), .b(G27), .O(gate471inter2));
  inv1  gate1040(.a(s_70), .O(gate471inter3));
  inv1  gate1041(.a(s_71), .O(gate471inter4));
  nand2 gate1042(.a(gate471inter4), .b(gate471inter3), .O(gate471inter5));
  nor2  gate1043(.a(gate471inter5), .b(gate471inter2), .O(gate471inter6));
  inv1  gate1044(.a(G27), .O(gate471inter7));
  inv1  gate1045(.a(G1210), .O(gate471inter8));
  nand2 gate1046(.a(gate471inter8), .b(gate471inter7), .O(gate471inter9));
  nand2 gate1047(.a(s_71), .b(gate471inter3), .O(gate471inter10));
  nor2  gate1048(.a(gate471inter10), .b(gate471inter9), .O(gate471inter11));
  nor2  gate1049(.a(gate471inter11), .b(gate471inter6), .O(gate471inter12));
  nand2 gate1050(.a(gate471inter12), .b(gate471inter1), .O(G1280));
nand2 gate472( .a(G1114), .b(G1210), .O(G1281) );
nand2 gate473( .a(G28), .b(G1213), .O(G1282) );

  xor2  gate1401(.a(G1213), .b(G1117), .O(gate474inter0));
  nand2 gate1402(.a(gate474inter0), .b(s_122), .O(gate474inter1));
  and2  gate1403(.a(G1213), .b(G1117), .O(gate474inter2));
  inv1  gate1404(.a(s_122), .O(gate474inter3));
  inv1  gate1405(.a(s_123), .O(gate474inter4));
  nand2 gate1406(.a(gate474inter4), .b(gate474inter3), .O(gate474inter5));
  nor2  gate1407(.a(gate474inter5), .b(gate474inter2), .O(gate474inter6));
  inv1  gate1408(.a(G1117), .O(gate474inter7));
  inv1  gate1409(.a(G1213), .O(gate474inter8));
  nand2 gate1410(.a(gate474inter8), .b(gate474inter7), .O(gate474inter9));
  nand2 gate1411(.a(s_123), .b(gate474inter3), .O(gate474inter10));
  nor2  gate1412(.a(gate474inter10), .b(gate474inter9), .O(gate474inter11));
  nor2  gate1413(.a(gate474inter11), .b(gate474inter6), .O(gate474inter12));
  nand2 gate1414(.a(gate474inter12), .b(gate474inter1), .O(G1283));

  xor2  gate1065(.a(G1216), .b(G29), .O(gate475inter0));
  nand2 gate1066(.a(gate475inter0), .b(s_74), .O(gate475inter1));
  and2  gate1067(.a(G1216), .b(G29), .O(gate475inter2));
  inv1  gate1068(.a(s_74), .O(gate475inter3));
  inv1  gate1069(.a(s_75), .O(gate475inter4));
  nand2 gate1070(.a(gate475inter4), .b(gate475inter3), .O(gate475inter5));
  nor2  gate1071(.a(gate475inter5), .b(gate475inter2), .O(gate475inter6));
  inv1  gate1072(.a(G29), .O(gate475inter7));
  inv1  gate1073(.a(G1216), .O(gate475inter8));
  nand2 gate1074(.a(gate475inter8), .b(gate475inter7), .O(gate475inter9));
  nand2 gate1075(.a(s_75), .b(gate475inter3), .O(gate475inter10));
  nor2  gate1076(.a(gate475inter10), .b(gate475inter9), .O(gate475inter11));
  nor2  gate1077(.a(gate475inter11), .b(gate475inter6), .O(gate475inter12));
  nand2 gate1078(.a(gate475inter12), .b(gate475inter1), .O(G1284));

  xor2  gate967(.a(G1216), .b(G1120), .O(gate476inter0));
  nand2 gate968(.a(gate476inter0), .b(s_60), .O(gate476inter1));
  and2  gate969(.a(G1216), .b(G1120), .O(gate476inter2));
  inv1  gate970(.a(s_60), .O(gate476inter3));
  inv1  gate971(.a(s_61), .O(gate476inter4));
  nand2 gate972(.a(gate476inter4), .b(gate476inter3), .O(gate476inter5));
  nor2  gate973(.a(gate476inter5), .b(gate476inter2), .O(gate476inter6));
  inv1  gate974(.a(G1120), .O(gate476inter7));
  inv1  gate975(.a(G1216), .O(gate476inter8));
  nand2 gate976(.a(gate476inter8), .b(gate476inter7), .O(gate476inter9));
  nand2 gate977(.a(s_61), .b(gate476inter3), .O(gate476inter10));
  nor2  gate978(.a(gate476inter10), .b(gate476inter9), .O(gate476inter11));
  nor2  gate979(.a(gate476inter11), .b(gate476inter6), .O(gate476inter12));
  nand2 gate980(.a(gate476inter12), .b(gate476inter1), .O(G1285));

  xor2  gate1765(.a(G1219), .b(G30), .O(gate477inter0));
  nand2 gate1766(.a(gate477inter0), .b(s_174), .O(gate477inter1));
  and2  gate1767(.a(G1219), .b(G30), .O(gate477inter2));
  inv1  gate1768(.a(s_174), .O(gate477inter3));
  inv1  gate1769(.a(s_175), .O(gate477inter4));
  nand2 gate1770(.a(gate477inter4), .b(gate477inter3), .O(gate477inter5));
  nor2  gate1771(.a(gate477inter5), .b(gate477inter2), .O(gate477inter6));
  inv1  gate1772(.a(G30), .O(gate477inter7));
  inv1  gate1773(.a(G1219), .O(gate477inter8));
  nand2 gate1774(.a(gate477inter8), .b(gate477inter7), .O(gate477inter9));
  nand2 gate1775(.a(s_175), .b(gate477inter3), .O(gate477inter10));
  nor2  gate1776(.a(gate477inter10), .b(gate477inter9), .O(gate477inter11));
  nor2  gate1777(.a(gate477inter11), .b(gate477inter6), .O(gate477inter12));
  nand2 gate1778(.a(gate477inter12), .b(gate477inter1), .O(G1286));

  xor2  gate1009(.a(G1219), .b(G1123), .O(gate478inter0));
  nand2 gate1010(.a(gate478inter0), .b(s_66), .O(gate478inter1));
  and2  gate1011(.a(G1219), .b(G1123), .O(gate478inter2));
  inv1  gate1012(.a(s_66), .O(gate478inter3));
  inv1  gate1013(.a(s_67), .O(gate478inter4));
  nand2 gate1014(.a(gate478inter4), .b(gate478inter3), .O(gate478inter5));
  nor2  gate1015(.a(gate478inter5), .b(gate478inter2), .O(gate478inter6));
  inv1  gate1016(.a(G1123), .O(gate478inter7));
  inv1  gate1017(.a(G1219), .O(gate478inter8));
  nand2 gate1018(.a(gate478inter8), .b(gate478inter7), .O(gate478inter9));
  nand2 gate1019(.a(s_67), .b(gate478inter3), .O(gate478inter10));
  nor2  gate1020(.a(gate478inter10), .b(gate478inter9), .O(gate478inter11));
  nor2  gate1021(.a(gate478inter11), .b(gate478inter6), .O(gate478inter12));
  nand2 gate1022(.a(gate478inter12), .b(gate478inter1), .O(G1287));
nand2 gate479( .a(G31), .b(G1222), .O(G1288) );
nand2 gate480( .a(G1126), .b(G1222), .O(G1289) );
nand2 gate481( .a(G32), .b(G1225), .O(G1290) );

  xor2  gate2619(.a(G1225), .b(G1129), .O(gate482inter0));
  nand2 gate2620(.a(gate482inter0), .b(s_296), .O(gate482inter1));
  and2  gate2621(.a(G1225), .b(G1129), .O(gate482inter2));
  inv1  gate2622(.a(s_296), .O(gate482inter3));
  inv1  gate2623(.a(s_297), .O(gate482inter4));
  nand2 gate2624(.a(gate482inter4), .b(gate482inter3), .O(gate482inter5));
  nor2  gate2625(.a(gate482inter5), .b(gate482inter2), .O(gate482inter6));
  inv1  gate2626(.a(G1129), .O(gate482inter7));
  inv1  gate2627(.a(G1225), .O(gate482inter8));
  nand2 gate2628(.a(gate482inter8), .b(gate482inter7), .O(gate482inter9));
  nand2 gate2629(.a(s_297), .b(gate482inter3), .O(gate482inter10));
  nor2  gate2630(.a(gate482inter10), .b(gate482inter9), .O(gate482inter11));
  nor2  gate2631(.a(gate482inter11), .b(gate482inter6), .O(gate482inter12));
  nand2 gate2632(.a(gate482inter12), .b(gate482inter1), .O(G1291));
nand2 gate483( .a(G1228), .b(G1229), .O(G1292) );
nand2 gate484( .a(G1230), .b(G1231), .O(G1293) );

  xor2  gate2507(.a(G1233), .b(G1232), .O(gate485inter0));
  nand2 gate2508(.a(gate485inter0), .b(s_280), .O(gate485inter1));
  and2  gate2509(.a(G1233), .b(G1232), .O(gate485inter2));
  inv1  gate2510(.a(s_280), .O(gate485inter3));
  inv1  gate2511(.a(s_281), .O(gate485inter4));
  nand2 gate2512(.a(gate485inter4), .b(gate485inter3), .O(gate485inter5));
  nor2  gate2513(.a(gate485inter5), .b(gate485inter2), .O(gate485inter6));
  inv1  gate2514(.a(G1232), .O(gate485inter7));
  inv1  gate2515(.a(G1233), .O(gate485inter8));
  nand2 gate2516(.a(gate485inter8), .b(gate485inter7), .O(gate485inter9));
  nand2 gate2517(.a(s_281), .b(gate485inter3), .O(gate485inter10));
  nor2  gate2518(.a(gate485inter10), .b(gate485inter9), .O(gate485inter11));
  nor2  gate2519(.a(gate485inter11), .b(gate485inter6), .O(gate485inter12));
  nand2 gate2520(.a(gate485inter12), .b(gate485inter1), .O(G1294));
nand2 gate486( .a(G1234), .b(G1235), .O(G1295) );
nand2 gate487( .a(G1236), .b(G1237), .O(G1296) );

  xor2  gate1625(.a(G1239), .b(G1238), .O(gate488inter0));
  nand2 gate1626(.a(gate488inter0), .b(s_154), .O(gate488inter1));
  and2  gate1627(.a(G1239), .b(G1238), .O(gate488inter2));
  inv1  gate1628(.a(s_154), .O(gate488inter3));
  inv1  gate1629(.a(s_155), .O(gate488inter4));
  nand2 gate1630(.a(gate488inter4), .b(gate488inter3), .O(gate488inter5));
  nor2  gate1631(.a(gate488inter5), .b(gate488inter2), .O(gate488inter6));
  inv1  gate1632(.a(G1238), .O(gate488inter7));
  inv1  gate1633(.a(G1239), .O(gate488inter8));
  nand2 gate1634(.a(gate488inter8), .b(gate488inter7), .O(gate488inter9));
  nand2 gate1635(.a(s_155), .b(gate488inter3), .O(gate488inter10));
  nor2  gate1636(.a(gate488inter10), .b(gate488inter9), .O(gate488inter11));
  nor2  gate1637(.a(gate488inter11), .b(gate488inter6), .O(gate488inter12));
  nand2 gate1638(.a(gate488inter12), .b(gate488inter1), .O(G1297));

  xor2  gate1191(.a(G1241), .b(G1240), .O(gate489inter0));
  nand2 gate1192(.a(gate489inter0), .b(s_92), .O(gate489inter1));
  and2  gate1193(.a(G1241), .b(G1240), .O(gate489inter2));
  inv1  gate1194(.a(s_92), .O(gate489inter3));
  inv1  gate1195(.a(s_93), .O(gate489inter4));
  nand2 gate1196(.a(gate489inter4), .b(gate489inter3), .O(gate489inter5));
  nor2  gate1197(.a(gate489inter5), .b(gate489inter2), .O(gate489inter6));
  inv1  gate1198(.a(G1240), .O(gate489inter7));
  inv1  gate1199(.a(G1241), .O(gate489inter8));
  nand2 gate1200(.a(gate489inter8), .b(gate489inter7), .O(gate489inter9));
  nand2 gate1201(.a(s_93), .b(gate489inter3), .O(gate489inter10));
  nor2  gate1202(.a(gate489inter10), .b(gate489inter9), .O(gate489inter11));
  nor2  gate1203(.a(gate489inter11), .b(gate489inter6), .O(gate489inter12));
  nand2 gate1204(.a(gate489inter12), .b(gate489inter1), .O(G1298));

  xor2  gate1023(.a(G1243), .b(G1242), .O(gate490inter0));
  nand2 gate1024(.a(gate490inter0), .b(s_68), .O(gate490inter1));
  and2  gate1025(.a(G1243), .b(G1242), .O(gate490inter2));
  inv1  gate1026(.a(s_68), .O(gate490inter3));
  inv1  gate1027(.a(s_69), .O(gate490inter4));
  nand2 gate1028(.a(gate490inter4), .b(gate490inter3), .O(gate490inter5));
  nor2  gate1029(.a(gate490inter5), .b(gate490inter2), .O(gate490inter6));
  inv1  gate1030(.a(G1242), .O(gate490inter7));
  inv1  gate1031(.a(G1243), .O(gate490inter8));
  nand2 gate1032(.a(gate490inter8), .b(gate490inter7), .O(gate490inter9));
  nand2 gate1033(.a(s_69), .b(gate490inter3), .O(gate490inter10));
  nor2  gate1034(.a(gate490inter10), .b(gate490inter9), .O(gate490inter11));
  nor2  gate1035(.a(gate490inter11), .b(gate490inter6), .O(gate490inter12));
  nand2 gate1036(.a(gate490inter12), .b(gate490inter1), .O(G1299));
nand2 gate491( .a(G1244), .b(G1245), .O(G1300) );
nand2 gate492( .a(G1246), .b(G1247), .O(G1301) );

  xor2  gate617(.a(G1249), .b(G1248), .O(gate493inter0));
  nand2 gate618(.a(gate493inter0), .b(s_10), .O(gate493inter1));
  and2  gate619(.a(G1249), .b(G1248), .O(gate493inter2));
  inv1  gate620(.a(s_10), .O(gate493inter3));
  inv1  gate621(.a(s_11), .O(gate493inter4));
  nand2 gate622(.a(gate493inter4), .b(gate493inter3), .O(gate493inter5));
  nor2  gate623(.a(gate493inter5), .b(gate493inter2), .O(gate493inter6));
  inv1  gate624(.a(G1248), .O(gate493inter7));
  inv1  gate625(.a(G1249), .O(gate493inter8));
  nand2 gate626(.a(gate493inter8), .b(gate493inter7), .O(gate493inter9));
  nand2 gate627(.a(s_11), .b(gate493inter3), .O(gate493inter10));
  nor2  gate628(.a(gate493inter10), .b(gate493inter9), .O(gate493inter11));
  nor2  gate629(.a(gate493inter11), .b(gate493inter6), .O(gate493inter12));
  nand2 gate630(.a(gate493inter12), .b(gate493inter1), .O(G1302));

  xor2  gate1317(.a(G1251), .b(G1250), .O(gate494inter0));
  nand2 gate1318(.a(gate494inter0), .b(s_110), .O(gate494inter1));
  and2  gate1319(.a(G1251), .b(G1250), .O(gate494inter2));
  inv1  gate1320(.a(s_110), .O(gate494inter3));
  inv1  gate1321(.a(s_111), .O(gate494inter4));
  nand2 gate1322(.a(gate494inter4), .b(gate494inter3), .O(gate494inter5));
  nor2  gate1323(.a(gate494inter5), .b(gate494inter2), .O(gate494inter6));
  inv1  gate1324(.a(G1250), .O(gate494inter7));
  inv1  gate1325(.a(G1251), .O(gate494inter8));
  nand2 gate1326(.a(gate494inter8), .b(gate494inter7), .O(gate494inter9));
  nand2 gate1327(.a(s_111), .b(gate494inter3), .O(gate494inter10));
  nor2  gate1328(.a(gate494inter10), .b(gate494inter9), .O(gate494inter11));
  nor2  gate1329(.a(gate494inter11), .b(gate494inter6), .O(gate494inter12));
  nand2 gate1330(.a(gate494inter12), .b(gate494inter1), .O(G1303));
nand2 gate495( .a(G1252), .b(G1253), .O(G1304) );
nand2 gate496( .a(G1254), .b(G1255), .O(G1305) );
nand2 gate497( .a(G1256), .b(G1257), .O(G1306) );
nand2 gate498( .a(G1258), .b(G1259), .O(G1307) );

  xor2  gate743(.a(G1261), .b(G1260), .O(gate499inter0));
  nand2 gate744(.a(gate499inter0), .b(s_28), .O(gate499inter1));
  and2  gate745(.a(G1261), .b(G1260), .O(gate499inter2));
  inv1  gate746(.a(s_28), .O(gate499inter3));
  inv1  gate747(.a(s_29), .O(gate499inter4));
  nand2 gate748(.a(gate499inter4), .b(gate499inter3), .O(gate499inter5));
  nor2  gate749(.a(gate499inter5), .b(gate499inter2), .O(gate499inter6));
  inv1  gate750(.a(G1260), .O(gate499inter7));
  inv1  gate751(.a(G1261), .O(gate499inter8));
  nand2 gate752(.a(gate499inter8), .b(gate499inter7), .O(gate499inter9));
  nand2 gate753(.a(s_29), .b(gate499inter3), .O(gate499inter10));
  nor2  gate754(.a(gate499inter10), .b(gate499inter9), .O(gate499inter11));
  nor2  gate755(.a(gate499inter11), .b(gate499inter6), .O(gate499inter12));
  nand2 gate756(.a(gate499inter12), .b(gate499inter1), .O(G1308));
nand2 gate500( .a(G1262), .b(G1263), .O(G1309) );

  xor2  gate953(.a(G1265), .b(G1264), .O(gate501inter0));
  nand2 gate954(.a(gate501inter0), .b(s_58), .O(gate501inter1));
  and2  gate955(.a(G1265), .b(G1264), .O(gate501inter2));
  inv1  gate956(.a(s_58), .O(gate501inter3));
  inv1  gate957(.a(s_59), .O(gate501inter4));
  nand2 gate958(.a(gate501inter4), .b(gate501inter3), .O(gate501inter5));
  nor2  gate959(.a(gate501inter5), .b(gate501inter2), .O(gate501inter6));
  inv1  gate960(.a(G1264), .O(gate501inter7));
  inv1  gate961(.a(G1265), .O(gate501inter8));
  nand2 gate962(.a(gate501inter8), .b(gate501inter7), .O(gate501inter9));
  nand2 gate963(.a(s_59), .b(gate501inter3), .O(gate501inter10));
  nor2  gate964(.a(gate501inter10), .b(gate501inter9), .O(gate501inter11));
  nor2  gate965(.a(gate501inter11), .b(gate501inter6), .O(gate501inter12));
  nand2 gate966(.a(gate501inter12), .b(gate501inter1), .O(G1310));

  xor2  gate1891(.a(G1267), .b(G1266), .O(gate502inter0));
  nand2 gate1892(.a(gate502inter0), .b(s_192), .O(gate502inter1));
  and2  gate1893(.a(G1267), .b(G1266), .O(gate502inter2));
  inv1  gate1894(.a(s_192), .O(gate502inter3));
  inv1  gate1895(.a(s_193), .O(gate502inter4));
  nand2 gate1896(.a(gate502inter4), .b(gate502inter3), .O(gate502inter5));
  nor2  gate1897(.a(gate502inter5), .b(gate502inter2), .O(gate502inter6));
  inv1  gate1898(.a(G1266), .O(gate502inter7));
  inv1  gate1899(.a(G1267), .O(gate502inter8));
  nand2 gate1900(.a(gate502inter8), .b(gate502inter7), .O(gate502inter9));
  nand2 gate1901(.a(s_193), .b(gate502inter3), .O(gate502inter10));
  nor2  gate1902(.a(gate502inter10), .b(gate502inter9), .O(gate502inter11));
  nor2  gate1903(.a(gate502inter11), .b(gate502inter6), .O(gate502inter12));
  nand2 gate1904(.a(gate502inter12), .b(gate502inter1), .O(G1311));
nand2 gate503( .a(G1268), .b(G1269), .O(G1312) );

  xor2  gate855(.a(G1271), .b(G1270), .O(gate504inter0));
  nand2 gate856(.a(gate504inter0), .b(s_44), .O(gate504inter1));
  and2  gate857(.a(G1271), .b(G1270), .O(gate504inter2));
  inv1  gate858(.a(s_44), .O(gate504inter3));
  inv1  gate859(.a(s_45), .O(gate504inter4));
  nand2 gate860(.a(gate504inter4), .b(gate504inter3), .O(gate504inter5));
  nor2  gate861(.a(gate504inter5), .b(gate504inter2), .O(gate504inter6));
  inv1  gate862(.a(G1270), .O(gate504inter7));
  inv1  gate863(.a(G1271), .O(gate504inter8));
  nand2 gate864(.a(gate504inter8), .b(gate504inter7), .O(gate504inter9));
  nand2 gate865(.a(s_45), .b(gate504inter3), .O(gate504inter10));
  nor2  gate866(.a(gate504inter10), .b(gate504inter9), .O(gate504inter11));
  nor2  gate867(.a(gate504inter11), .b(gate504inter6), .O(gate504inter12));
  nand2 gate868(.a(gate504inter12), .b(gate504inter1), .O(G1313));
nand2 gate505( .a(G1272), .b(G1273), .O(G1314) );
nand2 gate506( .a(G1274), .b(G1275), .O(G1315) );
nand2 gate507( .a(G1276), .b(G1277), .O(G1316) );
nand2 gate508( .a(G1278), .b(G1279), .O(G1317) );

  xor2  gate1135(.a(G1281), .b(G1280), .O(gate509inter0));
  nand2 gate1136(.a(gate509inter0), .b(s_84), .O(gate509inter1));
  and2  gate1137(.a(G1281), .b(G1280), .O(gate509inter2));
  inv1  gate1138(.a(s_84), .O(gate509inter3));
  inv1  gate1139(.a(s_85), .O(gate509inter4));
  nand2 gate1140(.a(gate509inter4), .b(gate509inter3), .O(gate509inter5));
  nor2  gate1141(.a(gate509inter5), .b(gate509inter2), .O(gate509inter6));
  inv1  gate1142(.a(G1280), .O(gate509inter7));
  inv1  gate1143(.a(G1281), .O(gate509inter8));
  nand2 gate1144(.a(gate509inter8), .b(gate509inter7), .O(gate509inter9));
  nand2 gate1145(.a(s_85), .b(gate509inter3), .O(gate509inter10));
  nor2  gate1146(.a(gate509inter10), .b(gate509inter9), .O(gate509inter11));
  nor2  gate1147(.a(gate509inter11), .b(gate509inter6), .O(gate509inter12));
  nand2 gate1148(.a(gate509inter12), .b(gate509inter1), .O(G1318));
nand2 gate510( .a(G1282), .b(G1283), .O(G1319) );
nand2 gate511( .a(G1284), .b(G1285), .O(G1320) );
nand2 gate512( .a(G1286), .b(G1287), .O(G1321) );

  xor2  gate1611(.a(G1289), .b(G1288), .O(gate513inter0));
  nand2 gate1612(.a(gate513inter0), .b(s_152), .O(gate513inter1));
  and2  gate1613(.a(G1289), .b(G1288), .O(gate513inter2));
  inv1  gate1614(.a(s_152), .O(gate513inter3));
  inv1  gate1615(.a(s_153), .O(gate513inter4));
  nand2 gate1616(.a(gate513inter4), .b(gate513inter3), .O(gate513inter5));
  nor2  gate1617(.a(gate513inter5), .b(gate513inter2), .O(gate513inter6));
  inv1  gate1618(.a(G1288), .O(gate513inter7));
  inv1  gate1619(.a(G1289), .O(gate513inter8));
  nand2 gate1620(.a(gate513inter8), .b(gate513inter7), .O(gate513inter9));
  nand2 gate1621(.a(s_153), .b(gate513inter3), .O(gate513inter10));
  nor2  gate1622(.a(gate513inter10), .b(gate513inter9), .O(gate513inter11));
  nor2  gate1623(.a(gate513inter11), .b(gate513inter6), .O(gate513inter12));
  nand2 gate1624(.a(gate513inter12), .b(gate513inter1), .O(G1322));
nand2 gate514( .a(G1290), .b(G1291), .O(G1323) );
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule