module c3540 (N1,N13,N20,N33,N41,N45,N50,N58,N68,N77,
              N87,N97,N107,N116,N124,N125,N128,N132,N137,N143,
              N150,N159,N169,N179,N190,N200,N213,N222,N223,N226,
              N232,N238,N244,N250,N257,N264,N270,N274,N283,N294,
              N303,N311,N317,N322,N326,N329,N330,N343,N349,N350,
              N1713,N1947,N3195,N3833,N3987,N4028,N4145,N4589,N4667,N4815,
              N4944,N5002,N5045,N5047,N5078,N5102,N5120,N5121,N5192,N5231,
              N5360,N5361);

input N1,N13,N20,N33,N41,N45,N50,N58,N68,N77,
      N87,N97,N107,N116,N124,N125,N128,N132,N137,N143,
      N150,N159,N169,N179,N190,N200,N213,N222,N223,N226,
      N232,N238,N244,N250,N257,N264,N270,N274,N283,N294,
      N303,N311,N317,N322,N326,N329,N330,N343,N349,N350;//RE__PI;

input s_0,s_1;//RE__ALLOW(00,01,10,11);
input s_2,s_3;//RE__ALLOW(00,01,10,11);
input s_4,s_5;//RE__ALLOW(00,01,10,11);
input s_6,s_7;//RE__ALLOW(00,01,10,11);
input s_8,s_9;//RE__ALLOW(00,01,10,11);
input s_10,s_11;//RE__ALLOW(00,01,10,11);
input s_12,s_13;//RE__ALLOW(00,01,10,11);
input s_14,s_15;//RE__ALLOW(00,01,10,11);
input s_16,s_17;//RE__ALLOW(00,01,10,11);
input s_18,s_19;//RE__ALLOW(00,01,10,11);
input s_20,s_21;//RE__ALLOW(00,01,10,11);
input s_22,s_23;//RE__ALLOW(00,01,10,11);
input s_24,s_25;//RE__ALLOW(00,01,10,11);
input s_26,s_27;//RE__ALLOW(00,01,10,11);
input s_28,s_29;//RE__ALLOW(00,01,10,11);
input s_30,s_31;//RE__ALLOW(00,01,10,11);
input s_32,s_33;//RE__ALLOW(00,01,10,11);
input s_34,s_35;//RE__ALLOW(00,01,10,11);
input s_36,s_37;//RE__ALLOW(00,01,10,11);
input s_38,s_39;//RE__ALLOW(00,01,10,11);
input s_40,s_41;//RE__ALLOW(00,01,10,11);
input s_42,s_43;//RE__ALLOW(00,01,10,11);
input s_44,s_45;//RE__ALLOW(00,01,10,11);
input s_46,s_47;//RE__ALLOW(00,01,10,11);
input s_48,s_49;//RE__ALLOW(00,01,10,11);
input s_50,s_51;//RE__ALLOW(00,01,10,11);
input s_52,s_53;//RE__ALLOW(00,01,10,11);
input s_54,s_55;//RE__ALLOW(00,01,10,11);
input s_56,s_57;//RE__ALLOW(00,01,10,11);
input s_58,s_59;//RE__ALLOW(00,01,10,11);
input s_60,s_61;//RE__ALLOW(00,01,10,11);
input s_62,s_63;//RE__ALLOW(00,01,10,11);
input s_64,s_65;//RE__ALLOW(00,01,10,11);
input s_66,s_67;//RE__ALLOW(00,01,10,11);
input s_68,s_69;//RE__ALLOW(00,01,10,11);
input s_70,s_71;//RE__ALLOW(00,01,10,11);
input s_72,s_73;//RE__ALLOW(00,01,10,11);
input s_74,s_75;//RE__ALLOW(00,01,10,11);
input s_76,s_77;//RE__ALLOW(00,01,10,11);
input s_78,s_79;//RE__ALLOW(00,01,10,11);
input s_80,s_81;//RE__ALLOW(00,01,10,11);
input s_82,s_83;//RE__ALLOW(00,01,10,11);
input s_84,s_85;//RE__ALLOW(00,01,10,11);
input s_86,s_87;//RE__ALLOW(00,01,10,11);
input s_88,s_89;//RE__ALLOW(00,01,10,11);
input s_90,s_91;//RE__ALLOW(00,01,10,11);
input s_92,s_93;//RE__ALLOW(00,01,10,11);
input s_94,s_95;//RE__ALLOW(00,01,10,11);
input s_96,s_97;//RE__ALLOW(00,01,10,11);
input s_98,s_99;//RE__ALLOW(00,01,10,11);
input s_100,s_101;//RE__ALLOW(00,01,10,11);
input s_102,s_103;//RE__ALLOW(00,01,10,11);
input s_104,s_105;//RE__ALLOW(00,01,10,11);
input s_106,s_107;//RE__ALLOW(00,01,10,11);
input s_108,s_109;//RE__ALLOW(00,01,10,11);
input s_110,s_111;//RE__ALLOW(00,01,10,11);
input s_112,s_113;//RE__ALLOW(00,01,10,11);
input s_114,s_115;//RE__ALLOW(00,01,10,11);
input s_116,s_117;//RE__ALLOW(00,01,10,11);
input s_118,s_119;//RE__ALLOW(00,01,10,11);
input s_120,s_121;//RE__ALLOW(00,01,10,11);
input s_122,s_123;//RE__ALLOW(00,01,10,11);
input s_124,s_125;//RE__ALLOW(00,01,10,11);
input s_126,s_127;//RE__ALLOW(00,01,10,11);
input s_128,s_129;//RE__ALLOW(00,01,10,11);
input s_130,s_131;//RE__ALLOW(00,01,10,11);
input s_132,s_133;//RE__ALLOW(00,01,10,11);
input s_134,s_135;//RE__ALLOW(00,01,10,11);
input s_136,s_137;//RE__ALLOW(00,01,10,11);
input s_138,s_139;//RE__ALLOW(00,01,10,11);
input s_140,s_141;//RE__ALLOW(00,01,10,11);
input s_142,s_143;//RE__ALLOW(00,01,10,11);
input s_144,s_145;//RE__ALLOW(00,01,10,11);
input s_146,s_147;//RE__ALLOW(00,01,10,11);
input s_148,s_149;//RE__ALLOW(00,01,10,11);
input s_150,s_151;//RE__ALLOW(00,01,10,11);
input s_152,s_153;//RE__ALLOW(00,01,10,11);
input s_154,s_155;//RE__ALLOW(00,01,10,11);
input s_156,s_157;//RE__ALLOW(00,01,10,11);
input s_158,s_159;//RE__ALLOW(00,01,10,11);
input s_160,s_161;//RE__ALLOW(00,01,10,11);
input s_162,s_163;//RE__ALLOW(00,01,10,11);
input s_164,s_165;//RE__ALLOW(00,01,10,11);
input s_166,s_167;//RE__ALLOW(00,01,10,11);
input s_168,s_169;//RE__ALLOW(00,01,10,11);
input s_170,s_171;//RE__ALLOW(00,01,10,11);
input s_172,s_173;//RE__ALLOW(00,01,10,11);
input s_174,s_175;//RE__ALLOW(00,01,10,11);
input s_176,s_177;//RE__ALLOW(00,01,10,11);
input s_178,s_179;//RE__ALLOW(00,01,10,11);
input s_180,s_181;//RE__ALLOW(00,01,10,11);
input s_182,s_183;//RE__ALLOW(00,01,10,11);
input s_184,s_185;//RE__ALLOW(00,01,10,11);
input s_186,s_187;//RE__ALLOW(00,01,10,11);
input s_188,s_189;//RE__ALLOW(00,01,10,11);
input s_190,s_191;//RE__ALLOW(00,01,10,11);
input s_192,s_193;//RE__ALLOW(00,01,10,11);
input s_194,s_195;//RE__ALLOW(00,01,10,11);
input s_196,s_197;//RE__ALLOW(00,01,10,11);
input s_198,s_199;//RE__ALLOW(00,01,10,11);
input s_200,s_201;//RE__ALLOW(00,01,10,11);
input s_202,s_203;//RE__ALLOW(00,01,10,11);
input s_204,s_205;//RE__ALLOW(00,01,10,11);
input s_206,s_207;//RE__ALLOW(00,01,10,11);
input s_208,s_209;//RE__ALLOW(00,01,10,11);
input s_210,s_211;//RE__ALLOW(00,01,10,11);
input s_212,s_213;//RE__ALLOW(00,01,10,11);
input s_214,s_215;//RE__ALLOW(00,01,10,11);
input s_216,s_217;//RE__ALLOW(00,01,10,11);
input s_218,s_219;//RE__ALLOW(00,01,10,11);
input s_220,s_221;//RE__ALLOW(00,01,10,11);
input s_222,s_223;//RE__ALLOW(00,01,10,11);
input s_224,s_225;//RE__ALLOW(00,01,10,11);
input s_226,s_227;//RE__ALLOW(00,01,10,11);
input s_228,s_229;//RE__ALLOW(00,01,10,11);
input s_230,s_231;//RE__ALLOW(00,01,10,11);
input s_232,s_233;//RE__ALLOW(00,01,10,11);
input s_234,s_235;//RE__ALLOW(00,01,10,11);
input s_236,s_237;//RE__ALLOW(00,01,10,11);
input s_238,s_239;//RE__ALLOW(00,01,10,11);
input s_240,s_241;//RE__ALLOW(00,01,10,11);
input s_242,s_243;//RE__ALLOW(00,01,10,11);
input s_244,s_245;//RE__ALLOW(00,01,10,11);
input s_246,s_247;//RE__ALLOW(00,01,10,11);
input s_248,s_249;//RE__ALLOW(00,01,10,11);
input s_250,s_251;//RE__ALLOW(00,01,10,11);
input s_252,s_253;//RE__ALLOW(00,01,10,11);
input s_254,s_255;//RE__ALLOW(00,01,10,11);
input s_256,s_257;//RE__ALLOW(00,01,10,11);
input s_258,s_259;//RE__ALLOW(00,01,10,11);
input s_260,s_261;//RE__ALLOW(00,01,10,11);
input s_262,s_263;//RE__ALLOW(00,01,10,11);
input s_264,s_265;//RE__ALLOW(00,01,10,11);
input s_266,s_267;//RE__ALLOW(00,01,10,11);
input s_268,s_269;//RE__ALLOW(00,01,10,11);
input s_270,s_271;//RE__ALLOW(00,01,10,11);
input s_272,s_273;//RE__ALLOW(00,01,10,11);
input s_274,s_275;//RE__ALLOW(00,01,10,11);
input s_276,s_277;//RE__ALLOW(00,01,10,11);
input s_278,s_279;//RE__ALLOW(00,01,10,11);
input s_280,s_281;//RE__ALLOW(00,01,10,11);
input s_282,s_283;//RE__ALLOW(00,01,10,11);
input s_284,s_285;//RE__ALLOW(00,01,10,11);
input s_286,s_287;//RE__ALLOW(00,01,10,11);
input s_288,s_289;//RE__ALLOW(00,01,10,11);
input s_290,s_291;//RE__ALLOW(00,01,10,11);
input s_292,s_293;//RE__ALLOW(00,01,10,11);
input s_294,s_295;//RE__ALLOW(00,01,10,11);
input s_296,s_297;//RE__ALLOW(00,01,10,11);
input s_298,s_299;//RE__ALLOW(00,01,10,11);
input s_300,s_301;//RE__ALLOW(00,01,10,11);
input s_302,s_303;//RE__ALLOW(00,01,10,11);
input s_304,s_305;//RE__ALLOW(00,01,10,11);
input s_306,s_307;//RE__ALLOW(00,01,10,11);
input s_308,s_309;//RE__ALLOW(00,01,10,11);
input s_310,s_311;//RE__ALLOW(00,01,10,11);
input s_312,s_313;//RE__ALLOW(00,01,10,11);
input s_314,s_315;//RE__ALLOW(00,01,10,11);
input s_316,s_317;//RE__ALLOW(00,01,10,11);
input s_318,s_319;//RE__ALLOW(00,01,10,11);
input s_320,s_321;//RE__ALLOW(00,01,10,11);
input s_322,s_323;//RE__ALLOW(00,01,10,11);
input s_324,s_325;//RE__ALLOW(00,01,10,11);
input s_326,s_327;//RE__ALLOW(00,01,10,11);
input s_328,s_329;//RE__ALLOW(00,01,10,11);
input s_330,s_331;//RE__ALLOW(00,01,10,11);
input s_332,s_333;//RE__ALLOW(00,01,10,11);
input s_334,s_335;//RE__ALLOW(00,01,10,11);
input s_336,s_337;//RE__ALLOW(00,01,10,11);
input s_338,s_339;//RE__ALLOW(00,01,10,11);
input s_340,s_341;//RE__ALLOW(00,01,10,11);
input s_342,s_343;//RE__ALLOW(00,01,10,11);
input s_344,s_345;//RE__ALLOW(00,01,10,11);
input s_346,s_347;//RE__ALLOW(00,01,10,11);
input s_348,s_349;//RE__ALLOW(00,01,10,11);
input s_350,s_351;//RE__ALLOW(00,01,10,11);
input s_352,s_353;//RE__ALLOW(00,01,10,11);
input s_354,s_355;//RE__ALLOW(00,01,10,11);
input s_356,s_357;//RE__ALLOW(00,01,10,11);
input s_358,s_359;//RE__ALLOW(00,01,10,11);
input s_360,s_361;//RE__ALLOW(00,01,10,11);
input s_362,s_363;//RE__ALLOW(00,01,10,11);
input s_364,s_365;//RE__ALLOW(00,01,10,11);
input s_366,s_367;//RE__ALLOW(00,01,10,11);
input s_368,s_369;//RE__ALLOW(00,01,10,11);
input s_370,s_371;//RE__ALLOW(00,01,10,11);
input s_372,s_373;//RE__ALLOW(00,01,10,11);
input s_374,s_375;//RE__ALLOW(00,01,10,11);
input s_376,s_377;//RE__ALLOW(00,01,10,11);
input s_378,s_379;//RE__ALLOW(00,01,10,11);
input s_380,s_381;//RE__ALLOW(00,01,10,11);
input s_382,s_383;//RE__ALLOW(00,01,10,11);
input s_384,s_385;//RE__ALLOW(00,01,10,11);
input s_386,s_387;//RE__ALLOW(00,01,10,11);
input s_388,s_389;//RE__ALLOW(00,01,10,11);
input s_390,s_391;//RE__ALLOW(00,01,10,11);
output N1713,N1947,N3195,N3833,N3987,N4028,N4145,N4589,N4667,N4815,
       N4944,N5002,N5045,N5047,N5078,N5102,N5120,N5121,N5192,N5231,
       N5360,N5361;

wire N655,N665,N670,N679,N683,N686,N690,N699,N702,N706,
     N715,N724,N727,N736,N740,N749,N753,N763,N768,N769,
     N772,N779,N782,N786,N793,N794,N798,N803,N820,N821,
     N825,N829,N832,N835,N836,N839,N842,N845,N848,N851,
     N854,N858,N861,N864,N867,N870,N874,N877,N880,N883,
     N886,N889,N890,N891,N892,N895,N896,N913,N914,N915,
     N916,N917,N920,N923,N926,N929,N932,N935,N938,N941,
     N944,N947,N950,N953,N956,N959,N962,N965,N1067,N1117,
     N1179,N1196,N1197,N1202,N1219,N1250,N1251,N1252,N1253,N1254,
     N1255,N1256,N1257,N1258,N1259,N1260,N1261,N1262,N1263,N1264,
     N1267,N1268,N1271,N1272,N1273,N1276,N1279,N1298,N1302,N1306,
     N1315,N1322,N1325,N1328,N1331,N1334,N1337,N1338,N1339,N1340,
     N1343,N1344,N1345,N1346,N1347,N1348,N1349,N1350,N1351,N1352,
     N1353,N1358,N1363,N1366,N1369,N1384,N1401,N1402,N1403,N1404,
     N1405,N1406,N1407,N1408,N1409,N1426,N1427,N1452,N1459,N1460,
     N1461,N1464,N1467,N1468,N1469,N1470,N1471,N1474,N1475,N1478,
     N1481,N1484,N1487,N1490,N1493,N1496,N1499,N1502,N1505,N1507,
     N1508,N1509,N1510,N1511,N1512,N1520,N1562,N1579,N1580,N1581,
     N1582,N1583,N1584,N1585,N1586,N1587,N1588,N1589,N1590,N1591,
     N1592,N1593,N1594,N1595,N1596,N1597,N1598,N1599,N1600,N1643,
     N1644,N1645,N1646,N1647,N1648,N1649,N1650,N1667,N1670,N1673,
     N1674,N1675,N1676,N1677,N1678,N1679,N1680,N1691,N1692,N1693,
     N1694,N1714,N1715,N1718,N1721,N1722,N1725,N1726,N1727,N1728,
     N1729,N1730,N1731,N1735,N1736,N1737,N1738,N1747,N1756,N1761,
     N1764,N1765,N1766,N1767,N1768,N1769,N1770,N1787,N1788,N1789,
     N1790,N1791,N1792,N1793,N1794,N1795,N1796,N1797,N1798,N1799,
     N1800,N1801,N1802,N1803,N1806,N1809,N1812,N1815,N1818,N1821,
     N1824,N1833,N1842,N1843,N1844,N1845,N1846,N1847,N1848,N1849,
     N1850,N1851,N1852,N1853,N1854,N1855,N1856,N1857,N1858,N1859,
     N1860,N1861,N1862,N1863,N1864,N1869,N1870,N1873,N1874,N1875,
     N1878,N1879,N1880,N1883,N1884,N1885,N1888,N1889,N1890,N1893,
     N1894,N1895,N1898,N1899,N1900,N1903,N1904,N1905,N1908,N1909,
     N1912,N1913,N1917,N1922,N1926,N1930,N1933,N1936,N1939,N1940,
     N1941,N1942,N1943,N1944,N1945,N1946,N1960,N1961,N1966,N1981,
     N1982,N1983,N1986,N1987,N1988,N1989,N1990,N1991,N2022,N2023,
     N2024,N2025,N2026,N2027,N2028,N2029,N2030,N2031,N2032,N2033,
     N2034,N2035,N2036,N2037,N2038,N2043,N2052,N2057,N2068,N2073,
     N2078,N2083,N2088,N2093,N2098,N2103,N2121,N2122,N2123,N2124,
     N2125,N2126,N2127,N2128,N2133,N2134,N2135,N2136,N2137,N2138,
     N2139,N2141,N2142,N2143,N2144,N2145,N2146,N2147,N2148,N2149,
     N2150,N2151,N2152,N2153,N2154,N2155,N2156,N2157,N2158,N2175,
     N2178,N2179,N2180,N2181,N2183,N2184,N2185,N2188,N2191,N2194,
     N2197,N2200,N2203,N2206,N2209,N2210,N2211,N2212,N2221,N2230,
     N2231,N2232,N2233,N2234,N2235,N2236,N2237,N2238,N2239,N2240,
     N2241,N2242,N2243,N2244,N2245,N2270,N2277,N2282,N2287,N2294,
     N2299,N2304,N2307,N2310,N2313,N2316,N2319,N2322,N2325,N2328,
     N2331,N2334,N2341,N2342,N2347,N2348,N2349,N2350,N2351,N2352,
     N2353,N2354,N2355,N2374,N2375,N2376,N2379,N2398,N2417,N2418,
     N2419,N2420,N2421,N2422,N2425,N2426,N2427,N2430,N2431,N2432,
     N2435,N2436,N2437,N2438,N2439,N2440,N2443,N2444,N2445,N2448,
     N2449,N2450,N2467,N2468,N2469,N2470,N2471,N2474,N2475,N2476,
     N2477,N2478,N2481,N2482,N2483,N2486,N2487,N2488,N2497,N2506,
     N2515,N2524,N2533,N2542,N2551,N2560,N2569,N2578,N2587,N2596,
     N2605,N2614,N2623,N2632,N2633,N2634,N2635,N2636,N2637,N2638,
     N2639,N2640,N2641,N2642,N2643,N2644,N2645,N2646,N2647,N2648,
     N2652,N2656,N2659,N2662,N2666,N2670,N2673,N2677,N2681,N2684,
     N2688,N2692,N2697,N2702,N2706,N2710,N2715,N2719,N2723,N2728,
     N2729,N2730,N2731,N2732,N2733,N2734,N2735,N2736,N2737,N2738,
     N2739,N2740,N2741,N2742,N2743,N2744,N2745,N2746,N2748,N2749,
     N2750,N2751,N2754,N2755,N2756,N2757,N2758,N2761,N2764,N2768,
     N2769,N2898,N2899,N2900,N2901,N2962,N2966,N2967,N2970,N2973,
     N2977,N2980,N2984,N2985,N2986,N2987,N2988,N2989,N2990,N2991,
     N2992,N2993,N2994,N2995,N2996,N2997,N2998,N2999,N3000,N3001,
     N3002,N3003,N3004,N3005,N3006,N3007,N3008,N3009,N3010,N3011,
     N3012,N3013,N3014,N3015,N3016,N3017,N3018,N3019,N3020,N3021,
     N3022,N3023,N3024,N3025,N3026,N3027,N3028,N3029,N3030,N3031,
     N3032,N3033,N3034,N3035,N3036,N3037,N3038,N3039,N3040,N3041,
     N3042,N3043,N3044,N3045,N3046,N3047,N3048,N3049,N3050,N3051,
     N3052,N3053,N3054,N3055,N3056,N3057,N3058,N3059,N3060,N3061,
     N3062,N3063,N3064,N3065,N3066,N3067,N3068,N3069,N3070,N3071,
     N3072,N3073,N3074,N3075,N3076,N3077,N3078,N3079,N3080,N3081,
     N3082,N3083,N3084,N3085,N3086,N3087,N3088,N3089,N3090,N3091,
     N3092,N3093,N3094,N3095,N3096,N3097,N3098,N3099,N3100,N3101,
     N3102,N3103,N3104,N3105,N3106,N3107,N3108,N3109,N3110,N3111,
     N3112,N3115,N3118,N3119,N3122,N3125,N3128,N3131,N3134,N3135,
     N3138,N3141,N3142,N3145,N3148,N3149,N3152,N3155,N3158,N3161,
     N3164,N3165,N3168,N3171,N3172,N3175,N3178,N3181,N3184,N3187,
     N3190,N3191,N3192,N3193,N3194,N3196,N3206,N3207,N3208,N3209,
     N3210,N3211,N3212,N3213,N3214,N3215,N3216,N3217,N3218,N3219,
     N3220,N3221,N3222,N3223,N3224,N3225,N3226,N3227,N3228,N3229,
     N3230,N3231,N3232,N3233,N3234,N3235,N3236,N3237,N3238,N3239,
     N3240,N3241,N3242,N3243,N3244,N3245,N3246,N3247,N3248,N3249,
     N3250,N3251,N3252,N3253,N3254,N3255,N3256,N3257,N3258,N3259,
     N3260,N3261,N3262,N3263,N3264,N3265,N3266,N3267,N3268,N3269,
     N3270,N3271,N3272,N3273,N3274,N3275,N3276,N3277,N3278,N3279,
     N3280,N3281,N3282,N3283,N3284,N3285,N3286,N3287,N3288,N3289,
     N3290,N3291,N3292,N3293,N3294,N3295,N3296,N3297,N3298,N3299,
     N3300,N3301,N3302,N3303,N3304,N3305,N3306,N3307,N3308,N3309,
     N3310,N3311,N3312,N3313,N3314,N3315,N3316,N3317,N3318,N3319,
     N3320,N3321,N3322,N3323,N3324,N3325,N3326,N3327,N3328,N3329,
     N3330,N3331,N3332,N3333,N3334,N3383,N3384,N3387,N3388,N3389,
     N3390,N3391,N3392,N3393,N3394,N3395,N3396,N3397,N3398,N3399,
     N3400,N3401,N3402,N3403,N3404,N3405,N3406,N3407,N3410,N3413,
     N3414,N3415,N3419,N3423,N3426,N3429,N3430,N3431,N3434,N3437,
     N3438,N3439,N3442,N3445,N3446,N3447,N3451,N3455,N3458,N3461,
     N3462,N3463,N3466,N3469,N3470,N3471,N3472,N3475,N3478,N3481,
     N3484,N3487,N3490,N3493,N3496,N3499,N3502,N3505,N3508,N3511,
     N3514,N3517,N3520,N3523,N3534,N3535,N3536,N3537,N3538,N3539,
     N3540,N3541,N3542,N3543,N3544,N3545,N3546,N3547,N3548,N3549,
     N3550,N3551,N3552,N3557,N3568,N3573,N3578,N3589,N3594,N3605,
     N3626,N3627,N3628,N3629,N3630,N3631,N3632,N3633,N3634,N3635,
     N3636,N3637,N3638,N3639,N3640,N3641,N3642,N3643,N3644,N3645,
     N3648,N3651,N3652,N3653,N3654,N3657,N3658,N3661,N3662,N3663,
     N3664,N3667,N3670,N3671,N3672,N3673,N3676,N3677,N3680,N3681,
     N3682,N3685,N3686,N3687,N3688,N3689,N3690,N3693,N3694,N3695,
     N3696,N3697,N3700,N3703,N3704,N3705,N3706,N3707,N3708,N3711,
     N3712,N3713,N3714,N3715,N3716,N3717,N3718,N3719,N3720,N3721,
     N3731,N3734,N3740,N3743,N3753,N3756,N3762,N3765,N3766,N3773,
     N3774,N3775,N3776,N3777,N3778,N3779,N3780,N3786,N3789,N3800,
     N3803,N3809,N3812,N3815,N3818,N3821,N3824,N3827,N3830,N3834,
     N3835,N3838,N3845,N3850,N3855,N3858,N3861,N3865,N3868,N3884,
     N3885,N3894,N3895,N3898,N3899,N3906,N3911,N3912,N3913,N3916,
     N3917,N3920,N3921,N3924,N3925,N3926,N3930,N3931,N3932,N3935,
     N3936,N3937,N3940,N3947,N3948,N3950,N3953,N3956,N3959,N3962,
     N3965,N3968,N3971,N3974,N3977,N3980,N3983,N3992,N3996,N4013,
     N4029,N4030,N4031,N4032,N4033,N4034,N4035,N4042,N4043,N4044,
     N4045,N4046,N4047,N4048,N4049,N4050,N4051,N4052,N4053,N4054,
     N4055,N4056,N4057,N4058,N4059,N4062,N4065,N4066,N4067,N4070,
     N4073,N4074,N4075,N4076,N4077,N4078,N4079,N4080,N4085,N4086,
     N4088,N4090,N4091,N4094,N4098,N4101,N4104,N4105,N4106,N4107,
     N4108,N4109,N4110,N4111,N4112,N4113,N4114,N4115,N4116,N4119,
     N4122,N4123,N4126,N4127,N4128,N4139,N4142,N4146,N4147,N4148,
     N4149,N4150,N4151,N4152,N4153,N4154,N4161,N4167,N4174,N4182,
     N4186,N4189,N4190,N4191,N4192,N4193,N4194,N4195,N4196,N4197,
     N4200,N4203,N4209,N4213,N4218,N4223,N4238,N4239,N4241,N4242,
     N4247,N4251,N4252,N4253,N4254,N4255,N4256,N4257,N4258,N4283,
     N4284,N4287,N4291,N4295,N4296,N4299,N4303,N4304,N4305,N4310,
     N4316,N4317,N4318,N4319,N4322,N4325,N4326,N4327,N4328,N4329,
     N4330,N4331,N4335,N4338,N4341,N4344,N4347,N4350,N4353,N4356,
     N4359,N4362,N4365,N4368,N4371,N4376,N4377,N4387,N4390,N4393,
     N4398,N4413,N4416,N4421,N4427,N4430,N4435,N4442,N4443,N4446,
     N4447,N4448,N4452,N4458,N4461,N4462,N4463,N4464,N4465,N4468,
     N4472,N4475,N4479,N4484,N4486,N4487,N4491,N4493,N4496,N4497,
     N4498,N4503,N4506,N4507,N4508,N4509,N4510,N4511,N4515,N4526,
     N4527,N4528,N4529,N4530,N4531,N4534,N4537,N4540,N4545,N4549,
     N4552,N4555,N4558,N4559,N4562,N4563,N4564,N4568,N4569,N4572,
     N4573,N4576,N4581,N4584,N4587,N4588,N4593,N4596,N4597,N4599,
     N4602,N4603,N4608,N4613,N4616,N4619,N4623,N4628,N4629,N4630,
     N4635,N4636,N4640,N4641,N4642,N4643,N4644,N4647,N4650,N4656,
     N4659,N4664,N4668,N4669,N4670,N4673,N4674,N4675,N4676,N4677,
     N4678,N4679,N4687,N4688,N4691,N4694,N4697,N4700,N4704,N4705,
     N4706,N4707,N4708,N4711,N4716,N4717,N4721,N4722,N4726,N4727,
     N4730,N4733,N4740,N4743,N4747,N4748,N4749,N4750,N4753,N4754,
     N4755,N4756,N4757,N4769,N4772,N4775,N4778,N4786,N4787,N4788,
     N4789,N4794,N4797,N4800,N4805,N4808,N4812,N4816,N4817,N4818,
     N4822,N4823,N4826,N4829,N4830,N4831,N4838,N4844,N4847,N4850,
     N4854,N4859,N4860,N4868,N4870,N4872,N4873,N4876,N4880,N4885,
     N4889,N4895,N4896,N4897,N4898,N4899,N4900,N4901,N4902,N4904,
     N4905,N4906,N4907,N4913,N4916,N4920,N4921,N4924,N4925,N4926,
     N4928,N4929,N4930,N4931,N4937,N4940,N4946,N4949,N4950,N4951,
     N4952,N4953,N4954,N4957,N4964,N4965,N4968,N4969,N4970,N4973,
     N4978,N4979,N4980,N4981,N4982,N4983,N4984,N4985,N4988,N4991,
     N4996,N4999,N5007,N5010,N5013,N5018,N5021,N5026,N5029,N5030,
     N5039,N5042,N5046,N5050,N5055,N5058,N5061,N5066,N5070,N5080,
     N5085,N5094,N5095,N5097,N5103,N5108,N5109,N5110,N5111,N5114,
     N5117,N5122,N5125,N5128,N5133,N5136,N5139,N5145,N5151,N5154,
     N5159,N5160,N5163,N5166,N5173,N5174,N5177,N5182,N5183,N5184,
     N5188,N5193,N5196,N5197,N5198,N5199,N5201,N5203,N5205,N5209,
     N5212,N5215,N5217,N5219,N5220,N5221,N5222,N5223,N5224,N5225,
     N5228,N5232,N5233,N5234,N5235,N5236,N5240,N5242,N5243,N5245,
     N5246,N5250,N5253,N5254,N5257,N5258,N5261,N5266,N5269,N5277,
     N5278,N5279,N5283,N5284,N5285,N5286,N5289,N5292,N5295,N5298,
     N5303,N5306,N5309,N5312,N5313,N5322,N5323,N5324,N5327,N5332,
     N5335,N5340,N5341,N5344,N5345,N5348,N5349,N5350,N5351,N5352,
     N5353,N5354,N5355,N5356,N5357,N5358,N5359, gate235inter0, gate235inter1, gate235inter2, gate235inter3, gate235inter4, gate235inter5, gate235inter6, gate235inter7, gate235inter8, gate235inter9, gate235inter10, gate235inter11, gate235inter12, gate388inter0, gate388inter1, gate388inter2, gate388inter3, gate388inter4, gate388inter5, gate388inter6, gate388inter7, gate388inter8, gate388inter9, gate388inter10, gate388inter11, gate388inter12, gate1375inter0, gate1375inter1, gate1375inter2, gate1375inter3, gate1375inter4, gate1375inter5, gate1375inter6, gate1375inter7, gate1375inter8, gate1375inter9, gate1375inter10, gate1375inter11, gate1375inter12, gate389inter0, gate389inter1, gate389inter2, gate389inter3, gate389inter4, gate389inter5, gate389inter6, gate389inter7, gate389inter8, gate389inter9, gate389inter10, gate389inter11, gate389inter12, gate595inter0, gate595inter1, gate595inter2, gate595inter3, gate595inter4, gate595inter5, gate595inter6, gate595inter7, gate595inter8, gate595inter9, gate595inter10, gate595inter11, gate595inter12, gate233inter0, gate233inter1, gate233inter2, gate233inter3, gate233inter4, gate233inter5, gate233inter6, gate233inter7, gate233inter8, gate233inter9, gate233inter10, gate233inter11, gate233inter12, gate226inter0, gate226inter1, gate226inter2, gate226inter3, gate226inter4, gate226inter5, gate226inter6, gate226inter7, gate226inter8, gate226inter9, gate226inter10, gate226inter11, gate226inter12, gate1487inter0, gate1487inter1, gate1487inter2, gate1487inter3, gate1487inter4, gate1487inter5, gate1487inter6, gate1487inter7, gate1487inter8, gate1487inter9, gate1487inter10, gate1487inter11, gate1487inter12, gate1486inter0, gate1486inter1, gate1486inter2, gate1486inter3, gate1486inter4, gate1486inter5, gate1486inter6, gate1486inter7, gate1486inter8, gate1486inter9, gate1486inter10, gate1486inter11, gate1486inter12, gate1423inter0, gate1423inter1, gate1423inter2, gate1423inter3, gate1423inter4, gate1423inter5, gate1423inter6, gate1423inter7, gate1423inter8, gate1423inter9, gate1423inter10, gate1423inter11, gate1423inter12, gate1616inter0, gate1616inter1, gate1616inter2, gate1616inter3, gate1616inter4, gate1616inter5, gate1616inter6, gate1616inter7, gate1616inter8, gate1616inter9, gate1616inter10, gate1616inter11, gate1616inter12, gate298inter0, gate298inter1, gate298inter2, gate298inter3, gate298inter4, gate298inter5, gate298inter6, gate298inter7, gate298inter8, gate298inter9, gate298inter10, gate298inter11, gate298inter12, gate1230inter0, gate1230inter1, gate1230inter2, gate1230inter3, gate1230inter4, gate1230inter5, gate1230inter6, gate1230inter7, gate1230inter8, gate1230inter9, gate1230inter10, gate1230inter11, gate1230inter12, gate1351inter0, gate1351inter1, gate1351inter2, gate1351inter3, gate1351inter4, gate1351inter5, gate1351inter6, gate1351inter7, gate1351inter8, gate1351inter9, gate1351inter10, gate1351inter11, gate1351inter12, gate1368inter0, gate1368inter1, gate1368inter2, gate1368inter3, gate1368inter4, gate1368inter5, gate1368inter6, gate1368inter7, gate1368inter8, gate1368inter9, gate1368inter10, gate1368inter11, gate1368inter12, gate1626inter0, gate1626inter1, gate1626inter2, gate1626inter3, gate1626inter4, gate1626inter5, gate1626inter6, gate1626inter7, gate1626inter8, gate1626inter9, gate1626inter10, gate1626inter11, gate1626inter12, gate1192inter0, gate1192inter1, gate1192inter2, gate1192inter3, gate1192inter4, gate1192inter5, gate1192inter6, gate1192inter7, gate1192inter8, gate1192inter9, gate1192inter10, gate1192inter11, gate1192inter12, gate509inter0, gate509inter1, gate509inter2, gate509inter3, gate509inter4, gate509inter5, gate509inter6, gate509inter7, gate509inter8, gate509inter9, gate509inter10, gate509inter11, gate509inter12, gate591inter0, gate591inter1, gate591inter2, gate591inter3, gate591inter4, gate591inter5, gate591inter6, gate591inter7, gate591inter8, gate591inter9, gate591inter10, gate591inter11, gate591inter12, gate173inter0, gate173inter1, gate173inter2, gate173inter3, gate173inter4, gate173inter5, gate173inter6, gate173inter7, gate173inter8, gate173inter9, gate173inter10, gate173inter11, gate173inter12, gate464inter0, gate464inter1, gate464inter2, gate464inter3, gate464inter4, gate464inter5, gate464inter6, gate464inter7, gate464inter8, gate464inter9, gate464inter10, gate464inter11, gate464inter12, gate1180inter0, gate1180inter1, gate1180inter2, gate1180inter3, gate1180inter4, gate1180inter5, gate1180inter6, gate1180inter7, gate1180inter8, gate1180inter9, gate1180inter10, gate1180inter11, gate1180inter12, gate1653inter0, gate1653inter1, gate1653inter2, gate1653inter3, gate1653inter4, gate1653inter5, gate1653inter6, gate1653inter7, gate1653inter8, gate1653inter9, gate1653inter10, gate1653inter11, gate1653inter12, gate1213inter0, gate1213inter1, gate1213inter2, gate1213inter3, gate1213inter4, gate1213inter5, gate1213inter6, gate1213inter7, gate1213inter8, gate1213inter9, gate1213inter10, gate1213inter11, gate1213inter12, gate1576inter0, gate1576inter1, gate1576inter2, gate1576inter3, gate1576inter4, gate1576inter5, gate1576inter6, gate1576inter7, gate1576inter8, gate1576inter9, gate1576inter10, gate1576inter11, gate1576inter12, gate1343inter0, gate1343inter1, gate1343inter2, gate1343inter3, gate1343inter4, gate1343inter5, gate1343inter6, gate1343inter7, gate1343inter8, gate1343inter9, gate1343inter10, gate1343inter11, gate1343inter12, gate1394inter0, gate1394inter1, gate1394inter2, gate1394inter3, gate1394inter4, gate1394inter5, gate1394inter6, gate1394inter7, gate1394inter8, gate1394inter9, gate1394inter10, gate1394inter11, gate1394inter12, gate1190inter0, gate1190inter1, gate1190inter2, gate1190inter3, gate1190inter4, gate1190inter5, gate1190inter6, gate1190inter7, gate1190inter8, gate1190inter9, gate1190inter10, gate1190inter11, gate1190inter12, gate1369inter0, gate1369inter1, gate1369inter2, gate1369inter3, gate1369inter4, gate1369inter5, gate1369inter6, gate1369inter7, gate1369inter8, gate1369inter9, gate1369inter10, gate1369inter11, gate1369inter12, gate778inter0, gate778inter1, gate778inter2, gate778inter3, gate778inter4, gate778inter5, gate778inter6, gate778inter7, gate778inter8, gate778inter9, gate778inter10, gate778inter11, gate778inter12, gate391inter0, gate391inter1, gate391inter2, gate391inter3, gate391inter4, gate391inter5, gate391inter6, gate391inter7, gate391inter8, gate391inter9, gate391inter10, gate391inter11, gate391inter12, gate269inter0, gate269inter1, gate269inter2, gate269inter3, gate269inter4, gate269inter5, gate269inter6, gate269inter7, gate269inter8, gate269inter9, gate269inter10, gate269inter11, gate269inter12, gate1447inter0, gate1447inter1, gate1447inter2, gate1447inter3, gate1447inter4, gate1447inter5, gate1447inter6, gate1447inter7, gate1447inter8, gate1447inter9, gate1447inter10, gate1447inter11, gate1447inter12, gate1114inter0, gate1114inter1, gate1114inter2, gate1114inter3, gate1114inter4, gate1114inter5, gate1114inter6, gate1114inter7, gate1114inter8, gate1114inter9, gate1114inter10, gate1114inter11, gate1114inter12, gate1608inter0, gate1608inter1, gate1608inter2, gate1608inter3, gate1608inter4, gate1608inter5, gate1608inter6, gate1608inter7, gate1608inter8, gate1608inter9, gate1608inter10, gate1608inter11, gate1608inter12, gate1161inter0, gate1161inter1, gate1161inter2, gate1161inter3, gate1161inter4, gate1161inter5, gate1161inter6, gate1161inter7, gate1161inter8, gate1161inter9, gate1161inter10, gate1161inter11, gate1161inter12, gate594inter0, gate594inter1, gate594inter2, gate594inter3, gate594inter4, gate594inter5, gate594inter6, gate594inter7, gate594inter8, gate594inter9, gate594inter10, gate594inter11, gate594inter12, gate90inter0, gate90inter1, gate90inter2, gate90inter3, gate90inter4, gate90inter5, gate90inter6, gate90inter7, gate90inter8, gate90inter9, gate90inter10, gate90inter11, gate90inter12, gate1247inter0, gate1247inter1, gate1247inter2, gate1247inter3, gate1247inter4, gate1247inter5, gate1247inter6, gate1247inter7, gate1247inter8, gate1247inter9, gate1247inter10, gate1247inter11, gate1247inter12, gate1627inter0, gate1627inter1, gate1627inter2, gate1627inter3, gate1627inter4, gate1627inter5, gate1627inter6, gate1627inter7, gate1627inter8, gate1627inter9, gate1627inter10, gate1627inter11, gate1627inter12, gate1201inter0, gate1201inter1, gate1201inter2, gate1201inter3, gate1201inter4, gate1201inter5, gate1201inter6, gate1201inter7, gate1201inter8, gate1201inter9, gate1201inter10, gate1201inter11, gate1201inter12, gate1449inter0, gate1449inter1, gate1449inter2, gate1449inter3, gate1449inter4, gate1449inter5, gate1449inter6, gate1449inter7, gate1449inter8, gate1449inter9, gate1449inter10, gate1449inter11, gate1449inter12, gate1060inter0, gate1060inter1, gate1060inter2, gate1060inter3, gate1060inter4, gate1060inter5, gate1060inter6, gate1060inter7, gate1060inter8, gate1060inter9, gate1060inter10, gate1060inter11, gate1060inter12, gate175inter0, gate175inter1, gate175inter2, gate175inter3, gate175inter4, gate175inter5, gate175inter6, gate175inter7, gate175inter8, gate175inter9, gate175inter10, gate175inter11, gate175inter12, gate413inter0, gate413inter1, gate413inter2, gate413inter3, gate413inter4, gate413inter5, gate413inter6, gate413inter7, gate413inter8, gate413inter9, gate413inter10, gate413inter11, gate413inter12, gate1591inter0, gate1591inter1, gate1591inter2, gate1591inter3, gate1591inter4, gate1591inter5, gate1591inter6, gate1591inter7, gate1591inter8, gate1591inter9, gate1591inter10, gate1591inter11, gate1591inter12, gate1614inter0, gate1614inter1, gate1614inter2, gate1614inter3, gate1614inter4, gate1614inter5, gate1614inter6, gate1614inter7, gate1614inter8, gate1614inter9, gate1614inter10, gate1614inter11, gate1614inter12, gate1462inter0, gate1462inter1, gate1462inter2, gate1462inter3, gate1462inter4, gate1462inter5, gate1462inter6, gate1462inter7, gate1462inter8, gate1462inter9, gate1462inter10, gate1462inter11, gate1462inter12, gate273inter0, gate273inter1, gate273inter2, gate273inter3, gate273inter4, gate273inter5, gate273inter6, gate273inter7, gate273inter8, gate273inter9, gate273inter10, gate273inter11, gate273inter12, gate1610inter0, gate1610inter1, gate1610inter2, gate1610inter3, gate1610inter4, gate1610inter5, gate1610inter6, gate1610inter7, gate1610inter8, gate1610inter9, gate1610inter10, gate1610inter11, gate1610inter12, gate1384inter0, gate1384inter1, gate1384inter2, gate1384inter3, gate1384inter4, gate1384inter5, gate1384inter6, gate1384inter7, gate1384inter8, gate1384inter9, gate1384inter10, gate1384inter11, gate1384inter12, gate88inter0, gate88inter1, gate88inter2, gate88inter3, gate88inter4, gate88inter5, gate88inter6, gate88inter7, gate88inter8, gate88inter9, gate88inter10, gate88inter11, gate88inter12, gate980inter0, gate980inter1, gate980inter2, gate980inter3, gate980inter4, gate980inter5, gate980inter6, gate980inter7, gate980inter8, gate980inter9, gate980inter10, gate980inter11, gate980inter12, gate1221inter0, gate1221inter1, gate1221inter2, gate1221inter3, gate1221inter4, gate1221inter5, gate1221inter6, gate1221inter7, gate1221inter8, gate1221inter9, gate1221inter10, gate1221inter11, gate1221inter12, gate316inter0, gate316inter1, gate316inter2, gate316inter3, gate316inter4, gate316inter5, gate316inter6, gate316inter7, gate316inter8, gate316inter9, gate316inter10, gate316inter11, gate316inter12, gate598inter0, gate598inter1, gate598inter2, gate598inter3, gate598inter4, gate598inter5, gate598inter6, gate598inter7, gate598inter8, gate598inter9, gate598inter10, gate598inter11, gate598inter12, gate462inter0, gate462inter1, gate462inter2, gate462inter3, gate462inter4, gate462inter5, gate462inter6, gate462inter7, gate462inter8, gate462inter9, gate462inter10, gate462inter11, gate462inter12, gate423inter0, gate423inter1, gate423inter2, gate423inter3, gate423inter4, gate423inter5, gate423inter6, gate423inter7, gate423inter8, gate423inter9, gate423inter10, gate423inter11, gate423inter12, gate1607inter0, gate1607inter1, gate1607inter2, gate1607inter3, gate1607inter4, gate1607inter5, gate1607inter6, gate1607inter7, gate1607inter8, gate1607inter9, gate1607inter10, gate1607inter11, gate1607inter12, gate1639inter0, gate1639inter1, gate1639inter2, gate1639inter3, gate1639inter4, gate1639inter5, gate1639inter6, gate1639inter7, gate1639inter8, gate1639inter9, gate1639inter10, gate1639inter11, gate1639inter12, gate1484inter0, gate1484inter1, gate1484inter2, gate1484inter3, gate1484inter4, gate1484inter5, gate1484inter6, gate1484inter7, gate1484inter8, gate1484inter9, gate1484inter10, gate1484inter11, gate1484inter12, gate414inter0, gate414inter1, gate414inter2, gate414inter3, gate414inter4, gate414inter5, gate414inter6, gate414inter7, gate414inter8, gate414inter9, gate414inter10, gate414inter11, gate414inter12, gate1604inter0, gate1604inter1, gate1604inter2, gate1604inter3, gate1604inter4, gate1604inter5, gate1604inter6, gate1604inter7, gate1604inter8, gate1604inter9, gate1604inter10, gate1604inter11, gate1604inter12, gate1223inter0, gate1223inter1, gate1223inter2, gate1223inter3, gate1223inter4, gate1223inter5, gate1223inter6, gate1223inter7, gate1223inter8, gate1223inter9, gate1223inter10, gate1223inter11, gate1223inter12, gate1152inter0, gate1152inter1, gate1152inter2, gate1152inter3, gate1152inter4, gate1152inter5, gate1152inter6, gate1152inter7, gate1152inter8, gate1152inter9, gate1152inter10, gate1152inter11, gate1152inter12, gate1162inter0, gate1162inter1, gate1162inter2, gate1162inter3, gate1162inter4, gate1162inter5, gate1162inter6, gate1162inter7, gate1162inter8, gate1162inter9, gate1162inter10, gate1162inter11, gate1162inter12, gate1501inter0, gate1501inter1, gate1501inter2, gate1501inter3, gate1501inter4, gate1501inter5, gate1501inter6, gate1501inter7, gate1501inter8, gate1501inter9, gate1501inter10, gate1501inter11, gate1501inter12, gate1177inter0, gate1177inter1, gate1177inter2, gate1177inter3, gate1177inter4, gate1177inter5, gate1177inter6, gate1177inter7, gate1177inter8, gate1177inter9, gate1177inter10, gate1177inter11, gate1177inter12, gate1562inter0, gate1562inter1, gate1562inter2, gate1562inter3, gate1562inter4, gate1562inter5, gate1562inter6, gate1562inter7, gate1562inter8, gate1562inter9, gate1562inter10, gate1562inter11, gate1562inter12, gate393inter0, gate393inter1, gate393inter2, gate393inter3, gate393inter4, gate393inter5, gate393inter6, gate393inter7, gate393inter8, gate393inter9, gate393inter10, gate393inter11, gate393inter12, gate456inter0, gate456inter1, gate456inter2, gate456inter3, gate456inter4, gate456inter5, gate456inter6, gate456inter7, gate456inter8, gate456inter9, gate456inter10, gate456inter11, gate456inter12, gate331inter0, gate331inter1, gate331inter2, gate331inter3, gate331inter4, gate331inter5, gate331inter6, gate331inter7, gate331inter8, gate331inter9, gate331inter10, gate331inter11, gate331inter12, gate1448inter0, gate1448inter1, gate1448inter2, gate1448inter3, gate1448inter4, gate1448inter5, gate1448inter6, gate1448inter7, gate1448inter8, gate1448inter9, gate1448inter10, gate1448inter11, gate1448inter12, gate593inter0, gate593inter1, gate593inter2, gate593inter3, gate593inter4, gate593inter5, gate593inter6, gate593inter7, gate593inter8, gate593inter9, gate593inter10, gate593inter11, gate593inter12, gate1498inter0, gate1498inter1, gate1498inter2, gate1498inter3, gate1498inter4, gate1498inter5, gate1498inter6, gate1498inter7, gate1498inter8, gate1498inter9, gate1498inter10, gate1498inter11, gate1498inter12, gate399inter0, gate399inter1, gate399inter2, gate399inter3, gate399inter4, gate399inter5, gate399inter6, gate399inter7, gate399inter8, gate399inter9, gate399inter10, gate399inter11, gate399inter12, gate1287inter0, gate1287inter1, gate1287inter2, gate1287inter3, gate1287inter4, gate1287inter5, gate1287inter6, gate1287inter7, gate1287inter8, gate1287inter9, gate1287inter10, gate1287inter11, gate1287inter12, gate1359inter0, gate1359inter1, gate1359inter2, gate1359inter3, gate1359inter4, gate1359inter5, gate1359inter6, gate1359inter7, gate1359inter8, gate1359inter9, gate1359inter10, gate1359inter11, gate1359inter12, gate1361inter0, gate1361inter1, gate1361inter2, gate1361inter3, gate1361inter4, gate1361inter5, gate1361inter6, gate1361inter7, gate1361inter8, gate1361inter9, gate1361inter10, gate1361inter11, gate1361inter12, gate1174inter0, gate1174inter1, gate1174inter2, gate1174inter3, gate1174inter4, gate1174inter5, gate1174inter6, gate1174inter7, gate1174inter8, gate1174inter9, gate1174inter10, gate1174inter11, gate1174inter12, gate1527inter0, gate1527inter1, gate1527inter2, gate1527inter3, gate1527inter4, gate1527inter5, gate1527inter6, gate1527inter7, gate1527inter8, gate1527inter9, gate1527inter10, gate1527inter11, gate1527inter12, gate400inter0, gate400inter1, gate400inter2, gate400inter3, gate400inter4, gate400inter5, gate400inter6, gate400inter7, gate400inter8, gate400inter9, gate400inter10, gate400inter11, gate400inter12, gate1503inter0, gate1503inter1, gate1503inter2, gate1503inter3, gate1503inter4, gate1503inter5, gate1503inter6, gate1503inter7, gate1503inter8, gate1503inter9, gate1503inter10, gate1503inter11, gate1503inter12, gate1187inter0, gate1187inter1, gate1187inter2, gate1187inter3, gate1187inter4, gate1187inter5, gate1187inter6, gate1187inter7, gate1187inter8, gate1187inter9, gate1187inter10, gate1187inter11, gate1187inter12, gate1195inter0, gate1195inter1, gate1195inter2, gate1195inter3, gate1195inter4, gate1195inter5, gate1195inter6, gate1195inter7, gate1195inter8, gate1195inter9, gate1195inter10, gate1195inter11, gate1195inter12, gate390inter0, gate390inter1, gate390inter2, gate390inter3, gate390inter4, gate390inter5, gate390inter6, gate390inter7, gate390inter8, gate390inter9, gate390inter10, gate390inter11, gate390inter12, gate101inter0, gate101inter1, gate101inter2, gate101inter3, gate101inter4, gate101inter5, gate101inter6, gate101inter7, gate101inter8, gate101inter9, gate101inter10, gate101inter11, gate101inter12, gate339inter0, gate339inter1, gate339inter2, gate339inter3, gate339inter4, gate339inter5, gate339inter6, gate339inter7, gate339inter8, gate339inter9, gate339inter10, gate339inter11, gate339inter12, gate1557inter0, gate1557inter1, gate1557inter2, gate1557inter3, gate1557inter4, gate1557inter5, gate1557inter6, gate1557inter7, gate1557inter8, gate1557inter9, gate1557inter10, gate1557inter11, gate1557inter12, gate1513inter0, gate1513inter1, gate1513inter2, gate1513inter3, gate1513inter4, gate1513inter5, gate1513inter6, gate1513inter7, gate1513inter8, gate1513inter9, gate1513inter10, gate1513inter11, gate1513inter12, gate1283inter0, gate1283inter1, gate1283inter2, gate1283inter3, gate1283inter4, gate1283inter5, gate1283inter6, gate1283inter7, gate1283inter8, gate1283inter9, gate1283inter10, gate1283inter11, gate1283inter12, gate1157inter0, gate1157inter1, gate1157inter2, gate1157inter3, gate1157inter4, gate1157inter5, gate1157inter6, gate1157inter7, gate1157inter8, gate1157inter9, gate1157inter10, gate1157inter11, gate1157inter12, gate1600inter0, gate1600inter1, gate1600inter2, gate1600inter3, gate1600inter4, gate1600inter5, gate1600inter6, gate1600inter7, gate1600inter8, gate1600inter9, gate1600inter10, gate1600inter11, gate1600inter12, gate174inter0, gate174inter1, gate174inter2, gate174inter3, gate174inter4, gate174inter5, gate174inter6, gate174inter7, gate174inter8, gate174inter9, gate174inter10, gate174inter11, gate174inter12, gate1665inter0, gate1665inter1, gate1665inter2, gate1665inter3, gate1665inter4, gate1665inter5, gate1665inter6, gate1665inter7, gate1665inter8, gate1665inter9, gate1665inter10, gate1665inter11, gate1665inter12, gate328inter0, gate328inter1, gate328inter2, gate328inter3, gate328inter4, gate328inter5, gate328inter6, gate328inter7, gate328inter8, gate328inter9, gate328inter10, gate328inter11, gate328inter12, gate1094inter0, gate1094inter1, gate1094inter2, gate1094inter3, gate1094inter4, gate1094inter5, gate1094inter6, gate1094inter7, gate1094inter8, gate1094inter9, gate1094inter10, gate1094inter11, gate1094inter12, gate1411inter0, gate1411inter1, gate1411inter2, gate1411inter3, gate1411inter4, gate1411inter5, gate1411inter6, gate1411inter7, gate1411inter8, gate1411inter9, gate1411inter10, gate1411inter11, gate1411inter12, gate310inter0, gate310inter1, gate310inter2, gate310inter3, gate310inter4, gate310inter5, gate310inter6, gate310inter7, gate310inter8, gate310inter9, gate310inter10, gate310inter11, gate310inter12, gate1464inter0, gate1464inter1, gate1464inter2, gate1464inter3, gate1464inter4, gate1464inter5, gate1464inter6, gate1464inter7, gate1464inter8, gate1464inter9, gate1464inter10, gate1464inter11, gate1464inter12, gate1317inter0, gate1317inter1, gate1317inter2, gate1317inter3, gate1317inter4, gate1317inter5, gate1317inter6, gate1317inter7, gate1317inter8, gate1317inter9, gate1317inter10, gate1317inter11, gate1317inter12, gate228inter0, gate228inter1, gate228inter2, gate228inter3, gate228inter4, gate228inter5, gate228inter6, gate228inter7, gate228inter8, gate228inter9, gate228inter10, gate228inter11, gate228inter12, gate1418inter0, gate1418inter1, gate1418inter2, gate1418inter3, gate1418inter4, gate1418inter5, gate1418inter6, gate1418inter7, gate1418inter8, gate1418inter9, gate1418inter10, gate1418inter11, gate1418inter12, gate244inter0, gate244inter1, gate244inter2, gate244inter3, gate244inter4, gate244inter5, gate244inter6, gate244inter7, gate244inter8, gate244inter9, gate244inter10, gate244inter11, gate244inter12, gate1378inter0, gate1378inter1, gate1378inter2, gate1378inter3, gate1378inter4, gate1378inter5, gate1378inter6, gate1378inter7, gate1378inter8, gate1378inter9, gate1378inter10, gate1378inter11, gate1378inter12, gate1625inter0, gate1625inter1, gate1625inter2, gate1625inter3, gate1625inter4, gate1625inter5, gate1625inter6, gate1625inter7, gate1625inter8, gate1625inter9, gate1625inter10, gate1625inter11, gate1625inter12, gate1656inter0, gate1656inter1, gate1656inter2, gate1656inter3, gate1656inter4, gate1656inter5, gate1656inter6, gate1656inter7, gate1656inter8, gate1656inter9, gate1656inter10, gate1656inter11, gate1656inter12, gate1226inter0, gate1226inter1, gate1226inter2, gate1226inter3, gate1226inter4, gate1226inter5, gate1226inter6, gate1226inter7, gate1226inter8, gate1226inter9, gate1226inter10, gate1226inter11, gate1226inter12, gate1204inter0, gate1204inter1, gate1204inter2, gate1204inter3, gate1204inter4, gate1204inter5, gate1204inter6, gate1204inter7, gate1204inter8, gate1204inter9, gate1204inter10, gate1204inter11, gate1204inter12, gate1324inter0, gate1324inter1, gate1324inter2, gate1324inter3, gate1324inter4, gate1324inter5, gate1324inter6, gate1324inter7, gate1324inter8, gate1324inter9, gate1324inter10, gate1324inter11, gate1324inter12, gate463inter0, gate463inter1, gate463inter2, gate463inter3, gate463inter4, gate463inter5, gate463inter6, gate463inter7, gate463inter8, gate463inter9, gate463inter10, gate463inter11, gate463inter12, gate89inter0, gate89inter1, gate89inter2, gate89inter3, gate89inter4, gate89inter5, gate89inter6, gate89inter7, gate89inter8, gate89inter9, gate89inter10, gate89inter11, gate89inter12, gate1666inter0, gate1666inter1, gate1666inter2, gate1666inter3, gate1666inter4, gate1666inter5, gate1666inter6, gate1666inter7, gate1666inter8, gate1666inter9, gate1666inter10, gate1666inter11, gate1666inter12, gate1115inter0, gate1115inter1, gate1115inter2, gate1115inter3, gate1115inter4, gate1115inter5, gate1115inter6, gate1115inter7, gate1115inter8, gate1115inter9, gate1115inter10, gate1115inter11, gate1115inter12, gate238inter0, gate238inter1, gate238inter2, gate238inter3, gate238inter4, gate238inter5, gate238inter6, gate238inter7, gate238inter8, gate238inter9, gate238inter10, gate238inter11, gate238inter12, gate424inter0, gate424inter1, gate424inter2, gate424inter3, gate424inter4, gate424inter5, gate424inter6, gate424inter7, gate424inter8, gate424inter9, gate424inter10, gate424inter11, gate424inter12, gate94inter0, gate94inter1, gate94inter2, gate94inter3, gate94inter4, gate94inter5, gate94inter6, gate94inter7, gate94inter8, gate94inter9, gate94inter10, gate94inter11, gate94inter12, gate1222inter0, gate1222inter1, gate1222inter2, gate1222inter3, gate1222inter4, gate1222inter5, gate1222inter6, gate1222inter7, gate1222inter8, gate1222inter9, gate1222inter10, gate1222inter11, gate1222inter12, gate1435inter0, gate1435inter1, gate1435inter2, gate1435inter3, gate1435inter4, gate1435inter5, gate1435inter6, gate1435inter7, gate1435inter8, gate1435inter9, gate1435inter10, gate1435inter11, gate1435inter12, gate1472inter0, gate1472inter1, gate1472inter2, gate1472inter3, gate1472inter4, gate1472inter5, gate1472inter6, gate1472inter7, gate1472inter8, gate1472inter9, gate1472inter10, gate1472inter11, gate1472inter12, gate1158inter0, gate1158inter1, gate1158inter2, gate1158inter3, gate1158inter4, gate1158inter5, gate1158inter6, gate1158inter7, gate1158inter8, gate1158inter9, gate1158inter10, gate1158inter11, gate1158inter12, gate1233inter0, gate1233inter1, gate1233inter2, gate1233inter3, gate1233inter4, gate1233inter5, gate1233inter6, gate1233inter7, gate1233inter8, gate1233inter9, gate1233inter10, gate1233inter11, gate1233inter12, gate87inter0, gate87inter1, gate87inter2, gate87inter3, gate87inter4, gate87inter5, gate87inter6, gate87inter7, gate87inter8, gate87inter9, gate87inter10, gate87inter11, gate87inter12, gate461inter0, gate461inter1, gate461inter2, gate461inter3, gate461inter4, gate461inter5, gate461inter6, gate461inter7, gate461inter8, gate461inter9, gate461inter10, gate461inter11, gate461inter12, gate1437inter0, gate1437inter1, gate1437inter2, gate1437inter3, gate1437inter4, gate1437inter5, gate1437inter6, gate1437inter7, gate1437inter8, gate1437inter9, gate1437inter10, gate1437inter11, gate1437inter12, gate1191inter0, gate1191inter1, gate1191inter2, gate1191inter3, gate1191inter4, gate1191inter5, gate1191inter6, gate1191inter7, gate1191inter8, gate1191inter9, gate1191inter10, gate1191inter11, gate1191inter12, gate1321inter0, gate1321inter1, gate1321inter2, gate1321inter3, gate1321inter4, gate1321inter5, gate1321inter6, gate1321inter7, gate1321inter8, gate1321inter9, gate1321inter10, gate1321inter11, gate1321inter12, gate1426inter0, gate1426inter1, gate1426inter2, gate1426inter3, gate1426inter4, gate1426inter5, gate1426inter6, gate1426inter7, gate1426inter8, gate1426inter9, gate1426inter10, gate1426inter11, gate1426inter12, gate465inter0, gate465inter1, gate465inter2, gate465inter3, gate465inter4, gate465inter5, gate465inter6, gate465inter7, gate465inter8, gate465inter9, gate465inter10, gate465inter11, gate465inter12, gate221inter0, gate221inter1, gate221inter2, gate221inter3, gate221inter4, gate221inter5, gate221inter6, gate221inter7, gate221inter8, gate221inter9, gate221inter10, gate221inter11, gate221inter12, gate220inter0, gate220inter1, gate220inter2, gate220inter3, gate220inter4, gate220inter5, gate220inter6, gate220inter7, gate220inter8, gate220inter9, gate220inter10, gate220inter11, gate220inter12, gate1519inter0, gate1519inter1, gate1519inter2, gate1519inter3, gate1519inter4, gate1519inter5, gate1519inter6, gate1519inter7, gate1519inter8, gate1519inter9, gate1519inter10, gate1519inter11, gate1519inter12, gate1433inter0, gate1433inter1, gate1433inter2, gate1433inter3, gate1433inter4, gate1433inter5, gate1433inter6, gate1433inter7, gate1433inter8, gate1433inter9, gate1433inter10, gate1433inter11, gate1433inter12, gate1473inter0, gate1473inter1, gate1473inter2, gate1473inter3, gate1473inter4, gate1473inter5, gate1473inter6, gate1473inter7, gate1473inter8, gate1473inter9, gate1473inter10, gate1473inter11, gate1473inter12, gate1571inter0, gate1571inter1, gate1571inter2, gate1571inter3, gate1571inter4, gate1571inter5, gate1571inter6, gate1571inter7, gate1571inter8, gate1571inter9, gate1571inter10, gate1571inter11, gate1571inter12, gate1624inter0, gate1624inter1, gate1624inter2, gate1624inter3, gate1624inter4, gate1624inter5, gate1624inter6, gate1624inter7, gate1624inter8, gate1624inter9, gate1624inter10, gate1624inter11, gate1624inter12, gate1482inter0, gate1482inter1, gate1482inter2, gate1482inter3, gate1482inter4, gate1482inter5, gate1482inter6, gate1482inter7, gate1482inter8, gate1482inter9, gate1482inter10, gate1482inter11, gate1482inter12, gate426inter0, gate426inter1, gate426inter2, gate426inter3, gate426inter4, gate426inter5, gate426inter6, gate426inter7, gate426inter8, gate426inter9, gate426inter10, gate426inter11, gate426inter12, gate1117inter0, gate1117inter1, gate1117inter2, gate1117inter3, gate1117inter4, gate1117inter5, gate1117inter6, gate1117inter7, gate1117inter8, gate1117inter9, gate1117inter10, gate1117inter11, gate1117inter12, gate1083inter0, gate1083inter1, gate1083inter2, gate1083inter3, gate1083inter4, gate1083inter5, gate1083inter6, gate1083inter7, gate1083inter8, gate1083inter9, gate1083inter10, gate1083inter11, gate1083inter12, gate1658inter0, gate1658inter1, gate1658inter2, gate1658inter3, gate1658inter4, gate1658inter5, gate1658inter6, gate1658inter7, gate1658inter8, gate1658inter9, gate1658inter10, gate1658inter11, gate1658inter12, gate1159inter0, gate1159inter1, gate1159inter2, gate1159inter3, gate1159inter4, gate1159inter5, gate1159inter6, gate1159inter7, gate1159inter8, gate1159inter9, gate1159inter10, gate1159inter11, gate1159inter12, gate1392inter0, gate1392inter1, gate1392inter2, gate1392inter3, gate1392inter4, gate1392inter5, gate1392inter6, gate1392inter7, gate1392inter8, gate1392inter9, gate1392inter10, gate1392inter11, gate1392inter12, gate1390inter0, gate1390inter1, gate1390inter2, gate1390inter3, gate1390inter4, gate1390inter5, gate1390inter6, gate1390inter7, gate1390inter8, gate1390inter9, gate1390inter10, gate1390inter11, gate1390inter12, gate1220inter0, gate1220inter1, gate1220inter2, gate1220inter3, gate1220inter4, gate1220inter5, gate1220inter6, gate1220inter7, gate1220inter8, gate1220inter9, gate1220inter10, gate1220inter11, gate1220inter12, gate1205inter0, gate1205inter1, gate1205inter2, gate1205inter3, gate1205inter4, gate1205inter5, gate1205inter6, gate1205inter7, gate1205inter8, gate1205inter9, gate1205inter10, gate1205inter11, gate1205inter12, gate425inter0, gate425inter1, gate425inter2, gate425inter3, gate425inter4, gate425inter5, gate425inter6, gate425inter7, gate425inter8, gate425inter9, gate425inter10, gate425inter11, gate425inter12, gate1407inter0, gate1407inter1, gate1407inter2, gate1407inter3, gate1407inter4, gate1407inter5, gate1407inter6, gate1407inter7, gate1407inter8, gate1407inter9, gate1407inter10, gate1407inter11, gate1407inter12, gate1520inter0, gate1520inter1, gate1520inter2, gate1520inter3, gate1520inter4, gate1520inter5, gate1520inter6, gate1520inter7, gate1520inter8, gate1520inter9, gate1520inter10, gate1520inter11, gate1520inter12, gate1425inter0, gate1425inter1, gate1425inter2, gate1425inter3, gate1425inter4, gate1425inter5, gate1425inter6, gate1425inter7, gate1425inter8, gate1425inter9, gate1425inter10, gate1425inter11, gate1425inter12, gate1333inter0, gate1333inter1, gate1333inter2, gate1333inter3, gate1333inter4, gate1333inter5, gate1333inter6, gate1333inter7, gate1333inter8, gate1333inter9, gate1333inter10, gate1333inter11, gate1333inter12, gate1619inter0, gate1619inter1, gate1619inter2, gate1619inter3, gate1619inter4, gate1619inter5, gate1619inter6, gate1619inter7, gate1619inter8, gate1619inter9, gate1619inter10, gate1619inter11, gate1619inter12, gate1197inter0, gate1197inter1, gate1197inter2, gate1197inter3, gate1197inter4, gate1197inter5, gate1197inter6, gate1197inter7, gate1197inter8, gate1197inter9, gate1197inter10, gate1197inter11, gate1197inter12, gate1657inter0, gate1657inter1, gate1657inter2, gate1657inter3, gate1657inter4, gate1657inter5, gate1657inter6, gate1657inter7, gate1657inter8, gate1657inter9, gate1657inter10, gate1657inter11, gate1657inter12, gate1206inter0, gate1206inter1, gate1206inter2, gate1206inter3, gate1206inter4, gate1206inter5, gate1206inter6, gate1206inter7, gate1206inter8, gate1206inter9, gate1206inter10, gate1206inter11, gate1206inter12, gate1207inter0, gate1207inter1, gate1207inter2, gate1207inter3, gate1207inter4, gate1207inter5, gate1207inter6, gate1207inter7, gate1207inter8, gate1207inter9, gate1207inter10, gate1207inter11, gate1207inter12, gate1492inter0, gate1492inter1, gate1492inter2, gate1492inter3, gate1492inter4, gate1492inter5, gate1492inter6, gate1492inter7, gate1492inter8, gate1492inter9, gate1492inter10, gate1492inter11, gate1492inter12, gate1160inter0, gate1160inter1, gate1160inter2, gate1160inter3, gate1160inter4, gate1160inter5, gate1160inter6, gate1160inter7, gate1160inter8, gate1160inter9, gate1160inter10, gate1160inter11, gate1160inter12, gate342inter0, gate342inter1, gate342inter2, gate342inter3, gate342inter4, gate342inter5, gate342inter6, gate342inter7, gate342inter8, gate342inter9, gate342inter10, gate342inter11, gate342inter12, gate610inter0, gate610inter1, gate610inter2, gate610inter3, gate610inter4, gate610inter5, gate610inter6, gate610inter7, gate610inter8, gate610inter9, gate610inter10, gate610inter11, gate610inter12, gate1103inter0, gate1103inter1, gate1103inter2, gate1103inter3, gate1103inter4, gate1103inter5, gate1103inter6, gate1103inter7, gate1103inter8, gate1103inter9, gate1103inter10, gate1103inter11, gate1103inter12, gate1395inter0, gate1395inter1, gate1395inter2, gate1395inter3, gate1395inter4, gate1395inter5, gate1395inter6, gate1395inter7, gate1395inter8, gate1395inter9, gate1395inter10, gate1395inter11, gate1395inter12, gate1663inter0, gate1663inter1, gate1663inter2, gate1663inter3, gate1663inter4, gate1663inter5, gate1663inter6, gate1663inter7, gate1663inter8, gate1663inter9, gate1663inter10, gate1663inter11, gate1663inter12, gate54inter0, gate54inter1, gate54inter2, gate54inter3, gate54inter4, gate54inter5, gate54inter6, gate54inter7, gate54inter8, gate54inter9, gate54inter10, gate54inter11, gate54inter12, gate1419inter0, gate1419inter1, gate1419inter2, gate1419inter3, gate1419inter4, gate1419inter5, gate1419inter6, gate1419inter7, gate1419inter8, gate1419inter9, gate1419inter10, gate1419inter11, gate1419inter12, gate1662inter0, gate1662inter1, gate1662inter2, gate1662inter3, gate1662inter4, gate1662inter5, gate1662inter6, gate1662inter7, gate1662inter8, gate1662inter9, gate1662inter10, gate1662inter11, gate1662inter12, gate1618inter0, gate1618inter1, gate1618inter2, gate1618inter3, gate1618inter4, gate1618inter5, gate1618inter6, gate1618inter7, gate1618inter8, gate1618inter9, gate1618inter10, gate1618inter11, gate1618inter12, gate1442inter0, gate1442inter1, gate1442inter2, gate1442inter3, gate1442inter4, gate1442inter5, gate1442inter6, gate1442inter7, gate1442inter8, gate1442inter9, gate1442inter10, gate1442inter11, gate1442inter12, gate343inter0, gate343inter1, gate343inter2, gate343inter3, gate343inter4, gate343inter5, gate343inter6, gate343inter7, gate343inter8, gate343inter9, gate343inter10, gate343inter11, gate343inter12, gate419inter0, gate419inter1, gate419inter2, gate419inter3, gate419inter4, gate419inter5, gate419inter6, gate419inter7, gate419inter8, gate419inter9, gate419inter10, gate419inter11, gate419inter12, gate1594inter0, gate1594inter1, gate1594inter2, gate1594inter3, gate1594inter4, gate1594inter5, gate1594inter6, gate1594inter7, gate1594inter8, gate1594inter9, gate1594inter10, gate1594inter11, gate1594inter12, gate1033inter0, gate1033inter1, gate1033inter2, gate1033inter3, gate1033inter4, gate1033inter5, gate1033inter6, gate1033inter7, gate1033inter8, gate1033inter9, gate1033inter10, gate1033inter11, gate1033inter12, gate219inter0, gate219inter1, gate219inter2, gate219inter3, gate219inter4, gate219inter5, gate219inter6, gate219inter7, gate219inter8, gate219inter9, gate219inter10, gate219inter11, gate219inter12, gate1059inter0, gate1059inter1, gate1059inter2, gate1059inter3, gate1059inter4, gate1059inter5, gate1059inter6, gate1059inter7, gate1059inter8, gate1059inter9, gate1059inter10, gate1059inter11, gate1059inter12, gate1491inter0, gate1491inter1, gate1491inter2, gate1491inter3, gate1491inter4, gate1491inter5, gate1491inter6, gate1491inter7, gate1491inter8, gate1491inter9, gate1491inter10, gate1491inter11, gate1491inter12, gate1605inter0, gate1605inter1, gate1605inter2, gate1605inter3, gate1605inter4, gate1605inter5, gate1605inter6, gate1605inter7, gate1605inter8, gate1605inter9, gate1605inter10, gate1605inter11, gate1605inter12, gate1643inter0, gate1643inter1, gate1643inter2, gate1643inter3, gate1643inter4, gate1643inter5, gate1643inter6, gate1643inter7, gate1643inter8, gate1643inter9, gate1643inter10, gate1643inter11, gate1643inter12, gate230inter0, gate230inter1, gate230inter2, gate230inter3, gate230inter4, gate230inter5, gate230inter6, gate230inter7, gate230inter8, gate230inter9, gate230inter10, gate230inter11, gate230inter12, gate93inter0, gate93inter1, gate93inter2, gate93inter3, gate93inter4, gate93inter5, gate93inter6, gate93inter7, gate93inter8, gate93inter9, gate93inter10, gate93inter11, gate93inter12, gate1509inter0, gate1509inter1, gate1509inter2, gate1509inter3, gate1509inter4, gate1509inter5, gate1509inter6, gate1509inter7, gate1509inter8, gate1509inter9, gate1509inter10, gate1509inter11, gate1509inter12, gate1620inter0, gate1620inter1, gate1620inter2, gate1620inter3, gate1620inter4, gate1620inter5, gate1620inter6, gate1620inter7, gate1620inter8, gate1620inter9, gate1620inter10, gate1620inter11, gate1620inter12, gate1461inter0, gate1461inter1, gate1461inter2, gate1461inter3, gate1461inter4, gate1461inter5, gate1461inter6, gate1461inter7, gate1461inter8, gate1461inter9, gate1461inter10, gate1461inter11, gate1461inter12, gate1210inter0, gate1210inter1, gate1210inter2, gate1210inter3, gate1210inter4, gate1210inter5, gate1210inter6, gate1210inter7, gate1210inter8, gate1210inter9, gate1210inter10, gate1210inter11, gate1210inter12, gate92inter0, gate92inter1, gate92inter2, gate92inter3, gate92inter4, gate92inter5, gate92inter6, gate92inter7, gate92inter8, gate92inter9, gate92inter10, gate92inter11, gate92inter12, gate132inter0, gate132inter1, gate132inter2, gate132inter3, gate132inter4, gate132inter5, gate132inter6, gate132inter7, gate132inter8, gate132inter9, gate132inter10, gate132inter11, gate132inter12, gate1409inter0, gate1409inter1, gate1409inter2, gate1409inter3, gate1409inter4, gate1409inter5, gate1409inter6, gate1409inter7, gate1409inter8, gate1409inter9, gate1409inter10, gate1409inter11, gate1409inter12, gate1240inter0, gate1240inter1, gate1240inter2, gate1240inter3, gate1240inter4, gate1240inter5, gate1240inter6, gate1240inter7, gate1240inter8, gate1240inter9, gate1240inter10, gate1240inter11, gate1240inter12, gate1029inter0, gate1029inter1, gate1029inter2, gate1029inter3, gate1029inter4, gate1029inter5, gate1029inter6, gate1029inter7, gate1029inter8, gate1029inter9, gate1029inter10, gate1029inter11, gate1029inter12, gate1499inter0, gate1499inter1, gate1499inter2, gate1499inter3, gate1499inter4, gate1499inter5, gate1499inter6, gate1499inter7, gate1499inter8, gate1499inter9, gate1499inter10, gate1499inter11, gate1499inter12, gate340inter0, gate340inter1, gate340inter2, gate340inter3, gate340inter4, gate340inter5, gate340inter6, gate340inter7, gate340inter8, gate340inter9, gate340inter10, gate340inter11, gate340inter12, gate301inter0, gate301inter1, gate301inter2, gate301inter3, gate301inter4, gate301inter5, gate301inter6, gate301inter7, gate301inter8, gate301inter9, gate301inter10, gate301inter11, gate301inter12, gate169inter0, gate169inter1, gate169inter2, gate169inter3, gate169inter4, gate169inter5, gate169inter6, gate169inter7, gate169inter8, gate169inter9, gate169inter10, gate169inter11, gate169inter12, gate1564inter0, gate1564inter1, gate1564inter2, gate1564inter3, gate1564inter4, gate1564inter5, gate1564inter6, gate1564inter7, gate1564inter8, gate1564inter9, gate1564inter10, gate1564inter11, gate1564inter12, gate592inter0, gate592inter1, gate592inter2, gate592inter3, gate592inter4, gate592inter5, gate592inter6, gate592inter7, gate592inter8, gate592inter9, gate592inter10, gate592inter11, gate592inter12, gate1202inter0, gate1202inter1, gate1202inter2, gate1202inter3, gate1202inter4, gate1202inter5, gate1202inter6, gate1202inter7, gate1202inter8, gate1202inter9, gate1202inter10, gate1202inter11, gate1202inter12, gate1104inter0, gate1104inter1, gate1104inter2, gate1104inter3, gate1104inter4, gate1104inter5, gate1104inter6, gate1104inter7, gate1104inter8, gate1104inter9, gate1104inter10, gate1104inter11, gate1104inter12;



buf1 gate1( .a(N50), .O(N655) );
inv1 gate2( .a(N50), .O(N665) );
buf1 gate3( .a(N58), .O(N670) );
inv1 gate4( .a(N58), .O(N679) );
buf1 gate5( .a(N68), .O(N683) );
inv1 gate6( .a(N68), .O(N686) );
buf1 gate7( .a(N68), .O(N690) );
buf1 gate8( .a(N77), .O(N699) );
inv1 gate9( .a(N77), .O(N702) );
buf1 gate10( .a(N77), .O(N706) );
buf1 gate11( .a(N87), .O(N715) );
inv1 gate12( .a(N87), .O(N724) );
buf1 gate13( .a(N97), .O(N727) );
inv1 gate14( .a(N97), .O(N736) );
buf1 gate15( .a(N107), .O(N740) );
inv1 gate16( .a(N107), .O(N749) );
buf1 gate17( .a(N116), .O(N753) );
inv1 gate18( .a(N116), .O(N763) );
or2 gate19( .a(N257), .b(N264), .O(N768) );
inv1 gate20( .a(N1), .O(N769) );
buf1 gate21( .a(N1), .O(N772) );
inv1 gate22( .a(N1), .O(N779) );
buf1 gate23( .a(N13), .O(N782) );
inv1 gate24( .a(N13), .O(N786) );
and2 gate25( .a(N13), .b(N20), .O(N793) );
inv1 gate26( .a(N20), .O(N794) );
buf1 gate27( .a(N20), .O(N798) );
inv1 gate28( .a(N20), .O(N803) );
inv1 gate29( .a(N33), .O(N820) );
buf1 gate30( .a(N33), .O(N821) );
inv1 gate31( .a(N33), .O(N825) );
and2 gate32( .a(N33), .b(N41), .O(N829) );
inv1 gate33( .a(N41), .O(N832) );
or2 gate34( .a(N41), .b(N45), .O(N835) );
buf1 gate35( .a(N45), .O(N836) );
inv1 gate36( .a(N45), .O(N839) );
inv1 gate37( .a(N50), .O(N842) );
buf1 gate38( .a(N58), .O(N845) );
inv1 gate39( .a(N58), .O(N848) );
buf1 gate40( .a(N68), .O(N851) );
inv1 gate41( .a(N68), .O(N854) );
buf1 gate42( .a(N87), .O(N858) );
inv1 gate43( .a(N87), .O(N861) );
buf1 gate44( .a(N97), .O(N864) );
inv1 gate45( .a(N97), .O(N867) );
inv1 gate46( .a(N107), .O(N870) );
buf1 gate47( .a(N1), .O(N874) );
buf1 gate48( .a(N68), .O(N877) );
buf1 gate49( .a(N107), .O(N880) );
inv1 gate50( .a(N20), .O(N883) );
buf1 gate51( .a(N190), .O(N886) );
inv1 gate52( .a(N200), .O(N889) );
and2 gate53( .a(N20), .b(N200), .O(N890) );

  xor2  gate3952(.a(N200), .b(N20), .O(gate54inter0));
  nand2 gate3953(.a(gate54inter0), .b(s_326), .O(gate54inter1));
  and2  gate3954(.a(N200), .b(N20), .O(gate54inter2));
  inv1  gate3955(.a(s_326), .O(gate54inter3));
  inv1  gate3956(.a(s_327), .O(gate54inter4));
  nand2 gate3957(.a(gate54inter4), .b(gate54inter3), .O(gate54inter5));
  nor2  gate3958(.a(gate54inter5), .b(gate54inter2), .O(gate54inter6));
  inv1  gate3959(.a(N20), .O(gate54inter7));
  inv1  gate3960(.a(N200), .O(gate54inter8));
  nand2 gate3961(.a(gate54inter8), .b(gate54inter7), .O(gate54inter9));
  nand2 gate3962(.a(s_327), .b(gate54inter3), .O(gate54inter10));
  nor2  gate3963(.a(gate54inter10), .b(gate54inter9), .O(gate54inter11));
  nor2  gate3964(.a(gate54inter11), .b(gate54inter6), .O(gate54inter12));
  nand2 gate3965(.a(gate54inter12), .b(gate54inter1), .O(N891));
and2 gate55( .a(N20), .b(N179), .O(N892) );
inv1 gate56( .a(N20), .O(N895) );
or2 gate57( .a(N349), .b(N33), .O(N896) );
nand2 gate58( .a(N1), .b(N13), .O(N913) );
nand3 gate59( .a(N1), .b(N20), .c(N33), .O(N914) );
inv1 gate60( .a(N20), .O(N915) );
inv1 gate61( .a(N33), .O(N916) );
buf1 gate62( .a(N179), .O(N917) );
inv1 gate63( .a(N213), .O(N920) );
buf1 gate64( .a(N343), .O(N923) );
buf1 gate65( .a(N226), .O(N926) );
buf1 gate66( .a(N232), .O(N929) );
buf1 gate67( .a(N238), .O(N932) );
buf1 gate68( .a(N244), .O(N935) );
buf1 gate69( .a(N250), .O(N938) );
buf1 gate70( .a(N257), .O(N941) );
buf1 gate71( .a(N264), .O(N944) );
buf1 gate72( .a(N270), .O(N947) );
buf1 gate73( .a(N50), .O(N950) );
buf1 gate74( .a(N58), .O(N953) );
buf1 gate75( .a(N58), .O(N956) );
buf1 gate76( .a(N97), .O(N959) );
buf1 gate77( .a(N97), .O(N962) );
buf1 gate78( .a(N330), .O(N965) );
and2 gate79( .a(N250), .b(N768), .O(N1067) );
or2 gate80( .a(N820), .b(N20), .O(N1117) );
or2 gate81( .a(N895), .b(N169), .O(N1179) );
inv1 gate82( .a(N793), .O(N1196) );
or2 gate83( .a(N915), .b(N1), .O(N1197) );
and2 gate84( .a(N913), .b(N914), .O(N1202) );
or2 gate85( .a(N916), .b(N1), .O(N1219) );
and3 gate86( .a(N842), .b(N848), .c(N854), .O(N1250) );

  xor2  gate3378(.a(N655), .b(N226), .O(gate87inter0));
  nand2 gate3379(.a(gate87inter0), .b(s_244), .O(gate87inter1));
  and2  gate3380(.a(N655), .b(N226), .O(gate87inter2));
  inv1  gate3381(.a(s_244), .O(gate87inter3));
  inv1  gate3382(.a(s_245), .O(gate87inter4));
  nand2 gate3383(.a(gate87inter4), .b(gate87inter3), .O(gate87inter5));
  nor2  gate3384(.a(gate87inter5), .b(gate87inter2), .O(gate87inter6));
  inv1  gate3385(.a(N226), .O(gate87inter7));
  inv1  gate3386(.a(N655), .O(gate87inter8));
  nand2 gate3387(.a(gate87inter8), .b(gate87inter7), .O(gate87inter9));
  nand2 gate3388(.a(s_245), .b(gate87inter3), .O(gate87inter10));
  nor2  gate3389(.a(gate87inter10), .b(gate87inter9), .O(gate87inter11));
  nor2  gate3390(.a(gate87inter11), .b(gate87inter6), .O(gate87inter12));
  nand2 gate3391(.a(gate87inter12), .b(gate87inter1), .O(N1251));

  xor2  gate2384(.a(N670), .b(N232), .O(gate88inter0));
  nand2 gate2385(.a(gate88inter0), .b(s_102), .O(gate88inter1));
  and2  gate2386(.a(N670), .b(N232), .O(gate88inter2));
  inv1  gate2387(.a(s_102), .O(gate88inter3));
  inv1  gate2388(.a(s_103), .O(gate88inter4));
  nand2 gate2389(.a(gate88inter4), .b(gate88inter3), .O(gate88inter5));
  nor2  gate2390(.a(gate88inter5), .b(gate88inter2), .O(gate88inter6));
  inv1  gate2391(.a(N232), .O(gate88inter7));
  inv1  gate2392(.a(N670), .O(gate88inter8));
  nand2 gate2393(.a(gate88inter8), .b(gate88inter7), .O(gate88inter9));
  nand2 gate2394(.a(s_103), .b(gate88inter3), .O(gate88inter10));
  nor2  gate2395(.a(gate88inter10), .b(gate88inter9), .O(gate88inter11));
  nor2  gate2396(.a(gate88inter11), .b(gate88inter6), .O(gate88inter12));
  nand2 gate2397(.a(gate88inter12), .b(gate88inter1), .O(N1252));

  xor2  gate3224(.a(N690), .b(N238), .O(gate89inter0));
  nand2 gate3225(.a(gate89inter0), .b(s_222), .O(gate89inter1));
  and2  gate3226(.a(N690), .b(N238), .O(gate89inter2));
  inv1  gate3227(.a(s_222), .O(gate89inter3));
  inv1  gate3228(.a(s_223), .O(gate89inter4));
  nand2 gate3229(.a(gate89inter4), .b(gate89inter3), .O(gate89inter5));
  nor2  gate3230(.a(gate89inter5), .b(gate89inter2), .O(gate89inter6));
  inv1  gate3231(.a(N238), .O(gate89inter7));
  inv1  gate3232(.a(N690), .O(gate89inter8));
  nand2 gate3233(.a(gate89inter8), .b(gate89inter7), .O(gate89inter9));
  nand2 gate3234(.a(s_223), .b(gate89inter3), .O(gate89inter10));
  nor2  gate3235(.a(gate89inter10), .b(gate89inter9), .O(gate89inter11));
  nor2  gate3236(.a(gate89inter11), .b(gate89inter6), .O(gate89inter12));
  nand2 gate3237(.a(gate89inter12), .b(gate89inter1), .O(N1253));

  xor2  gate2188(.a(N706), .b(N244), .O(gate90inter0));
  nand2 gate2189(.a(gate90inter0), .b(s_74), .O(gate90inter1));
  and2  gate2190(.a(N706), .b(N244), .O(gate90inter2));
  inv1  gate2191(.a(s_74), .O(gate90inter3));
  inv1  gate2192(.a(s_75), .O(gate90inter4));
  nand2 gate2193(.a(gate90inter4), .b(gate90inter3), .O(gate90inter5));
  nor2  gate2194(.a(gate90inter5), .b(gate90inter2), .O(gate90inter6));
  inv1  gate2195(.a(N244), .O(gate90inter7));
  inv1  gate2196(.a(N706), .O(gate90inter8));
  nand2 gate2197(.a(gate90inter8), .b(gate90inter7), .O(gate90inter9));
  nand2 gate2198(.a(s_75), .b(gate90inter3), .O(gate90inter10));
  nor2  gate2199(.a(gate90inter10), .b(gate90inter9), .O(gate90inter11));
  nor2  gate2200(.a(gate90inter11), .b(gate90inter6), .O(gate90inter12));
  nand2 gate2201(.a(gate90inter12), .b(gate90inter1), .O(N1254));
nand2 gate91( .a(N250), .b(N715), .O(N1255) );

  xor2  gate4232(.a(N727), .b(N257), .O(gate92inter0));
  nand2 gate4233(.a(gate92inter0), .b(s_366), .O(gate92inter1));
  and2  gate4234(.a(N727), .b(N257), .O(gate92inter2));
  inv1  gate4235(.a(s_366), .O(gate92inter3));
  inv1  gate4236(.a(s_367), .O(gate92inter4));
  nand2 gate4237(.a(gate92inter4), .b(gate92inter3), .O(gate92inter5));
  nor2  gate4238(.a(gate92inter5), .b(gate92inter2), .O(gate92inter6));
  inv1  gate4239(.a(N257), .O(gate92inter7));
  inv1  gate4240(.a(N727), .O(gate92inter8));
  nand2 gate4241(.a(gate92inter8), .b(gate92inter7), .O(gate92inter9));
  nand2 gate4242(.a(s_367), .b(gate92inter3), .O(gate92inter10));
  nor2  gate4243(.a(gate92inter10), .b(gate92inter9), .O(gate92inter11));
  nor2  gate4244(.a(gate92inter11), .b(gate92inter6), .O(gate92inter12));
  nand2 gate4245(.a(gate92inter12), .b(gate92inter1), .O(N1256));

  xor2  gate4162(.a(N740), .b(N264), .O(gate93inter0));
  nand2 gate4163(.a(gate93inter0), .b(s_356), .O(gate93inter1));
  and2  gate4164(.a(N740), .b(N264), .O(gate93inter2));
  inv1  gate4165(.a(s_356), .O(gate93inter3));
  inv1  gate4166(.a(s_357), .O(gate93inter4));
  nand2 gate4167(.a(gate93inter4), .b(gate93inter3), .O(gate93inter5));
  nor2  gate4168(.a(gate93inter5), .b(gate93inter2), .O(gate93inter6));
  inv1  gate4169(.a(N264), .O(gate93inter7));
  inv1  gate4170(.a(N740), .O(gate93inter8));
  nand2 gate4171(.a(gate93inter8), .b(gate93inter7), .O(gate93inter9));
  nand2 gate4172(.a(s_357), .b(gate93inter3), .O(gate93inter10));
  nor2  gate4173(.a(gate93inter10), .b(gate93inter9), .O(gate93inter11));
  nor2  gate4174(.a(gate93inter11), .b(gate93inter6), .O(gate93inter12));
  nand2 gate4175(.a(gate93inter12), .b(gate93inter1), .O(N1257));

  xor2  gate3294(.a(N753), .b(N270), .O(gate94inter0));
  nand2 gate3295(.a(gate94inter0), .b(s_232), .O(gate94inter1));
  and2  gate3296(.a(N753), .b(N270), .O(gate94inter2));
  inv1  gate3297(.a(s_232), .O(gate94inter3));
  inv1  gate3298(.a(s_233), .O(gate94inter4));
  nand2 gate3299(.a(gate94inter4), .b(gate94inter3), .O(gate94inter5));
  nor2  gate3300(.a(gate94inter5), .b(gate94inter2), .O(gate94inter6));
  inv1  gate3301(.a(N270), .O(gate94inter7));
  inv1  gate3302(.a(N753), .O(gate94inter8));
  nand2 gate3303(.a(gate94inter8), .b(gate94inter7), .O(gate94inter9));
  nand2 gate3304(.a(s_233), .b(gate94inter3), .O(gate94inter10));
  nor2  gate3305(.a(gate94inter10), .b(gate94inter9), .O(gate94inter11));
  nor2  gate3306(.a(gate94inter11), .b(gate94inter6), .O(gate94inter12));
  nand2 gate3307(.a(gate94inter12), .b(gate94inter1), .O(N1258));
inv1 gate95( .a(N926), .O(N1259) );
inv1 gate96( .a(N929), .O(N1260) );
inv1 gate97( .a(N932), .O(N1261) );
inv1 gate98( .a(N935), .O(N1262) );
nand2 gate99( .a(N679), .b(N686), .O(N1263) );
nand2 gate100( .a(N736), .b(N749), .O(N1264) );

  xor2  gate2874(.a(N699), .b(N683), .O(gate101inter0));
  nand2 gate2875(.a(gate101inter0), .b(s_172), .O(gate101inter1));
  and2  gate2876(.a(N699), .b(N683), .O(gate101inter2));
  inv1  gate2877(.a(s_172), .O(gate101inter3));
  inv1  gate2878(.a(s_173), .O(gate101inter4));
  nand2 gate2879(.a(gate101inter4), .b(gate101inter3), .O(gate101inter5));
  nor2  gate2880(.a(gate101inter5), .b(gate101inter2), .O(gate101inter6));
  inv1  gate2881(.a(N683), .O(gate101inter7));
  inv1  gate2882(.a(N699), .O(gate101inter8));
  nand2 gate2883(.a(gate101inter8), .b(gate101inter7), .O(gate101inter9));
  nand2 gate2884(.a(s_173), .b(gate101inter3), .O(gate101inter10));
  nor2  gate2885(.a(gate101inter10), .b(gate101inter9), .O(gate101inter11));
  nor2  gate2886(.a(gate101inter11), .b(gate101inter6), .O(gate101inter12));
  nand2 gate2887(.a(gate101inter12), .b(gate101inter1), .O(N1267));
buf1 gate102( .a(N665), .O(N1268) );
inv1 gate103( .a(N953), .O(N1271) );
inv1 gate104( .a(N959), .O(N1272) );
buf1 gate105( .a(N839), .O(N1273) );
buf1 gate106( .a(N839), .O(N1276) );
buf1 gate107( .a(N782), .O(N1279) );
buf1 gate108( .a(N825), .O(N1298) );
buf1 gate109( .a(N832), .O(N1302) );
and2 gate110( .a(N779), .b(N835), .O(N1306) );
and3 gate111( .a(N779), .b(N836), .c(N832), .O(N1315) );
and2 gate112( .a(N769), .b(N836), .O(N1322) );
and3 gate113( .a(N772), .b(N786), .c(N798), .O(N1325) );
nand3 gate114( .a(N772), .b(N786), .c(N798), .O(N1328) );
nand2 gate115( .a(N772), .b(N786), .O(N1331) );
buf1 gate116( .a(N874), .O(N1334) );
nand3 gate117( .a(N782), .b(N794), .c(N45), .O(N1337) );
nand3 gate118( .a(N842), .b(N848), .c(N854), .O(N1338) );
inv1 gate119( .a(N956), .O(N1339) );
and3 gate120( .a(N861), .b(N867), .c(N870), .O(N1340) );
nand3 gate121( .a(N861), .b(N867), .c(N870), .O(N1343) );
inv1 gate122( .a(N962), .O(N1344) );
inv1 gate123( .a(N803), .O(N1345) );
inv1 gate124( .a(N803), .O(N1346) );
inv1 gate125( .a(N803), .O(N1347) );
inv1 gate126( .a(N803), .O(N1348) );
inv1 gate127( .a(N803), .O(N1349) );
inv1 gate128( .a(N803), .O(N1350) );
inv1 gate129( .a(N803), .O(N1351) );
inv1 gate130( .a(N803), .O(N1352) );
or2 gate131( .a(N883), .b(N886), .O(N1353) );

  xor2  gate4246(.a(N886), .b(N883), .O(gate132inter0));
  nand2 gate4247(.a(gate132inter0), .b(s_368), .O(gate132inter1));
  and2  gate4248(.a(N886), .b(N883), .O(gate132inter2));
  inv1  gate4249(.a(s_368), .O(gate132inter3));
  inv1  gate4250(.a(s_369), .O(gate132inter4));
  nand2 gate4251(.a(gate132inter4), .b(gate132inter3), .O(gate132inter5));
  nor2  gate4252(.a(gate132inter5), .b(gate132inter2), .O(gate132inter6));
  inv1  gate4253(.a(N883), .O(gate132inter7));
  inv1  gate4254(.a(N886), .O(gate132inter8));
  nand2 gate4255(.a(gate132inter8), .b(gate132inter7), .O(gate132inter9));
  nand2 gate4256(.a(s_369), .b(gate132inter3), .O(gate132inter10));
  nor2  gate4257(.a(gate132inter10), .b(gate132inter9), .O(gate132inter11));
  nor2  gate4258(.a(gate132inter11), .b(gate132inter6), .O(gate132inter12));
  nand2 gate4259(.a(gate132inter12), .b(gate132inter1), .O(N1358));
buf1 gate133( .a(N892), .O(N1363) );
inv1 gate134( .a(N892), .O(N1366) );
buf1 gate135( .a(N821), .O(N1369) );
buf1 gate136( .a(N825), .O(N1384) );
inv1 gate137( .a(N896), .O(N1401) );
inv1 gate138( .a(N896), .O(N1402) );
inv1 gate139( .a(N896), .O(N1403) );
inv1 gate140( .a(N896), .O(N1404) );
inv1 gate141( .a(N896), .O(N1405) );
inv1 gate142( .a(N896), .O(N1406) );
inv1 gate143( .a(N896), .O(N1407) );
inv1 gate144( .a(N896), .O(N1408) );
or2 gate145( .a(N1), .b(N1196), .O(N1409) );
inv1 gate146( .a(N829), .O(N1426) );
inv1 gate147( .a(N829), .O(N1427) );
and3 gate148( .a(N769), .b(N782), .c(N794), .O(N1452) );
inv1 gate149( .a(N917), .O(N1459) );
inv1 gate150( .a(N965), .O(N1460) );
or2 gate151( .a(N920), .b(N923), .O(N1461) );
nor2 gate152( .a(N920), .b(N923), .O(N1464) );
inv1 gate153( .a(N938), .O(N1467) );
inv1 gate154( .a(N941), .O(N1468) );
inv1 gate155( .a(N944), .O(N1469) );
inv1 gate156( .a(N947), .O(N1470) );
buf1 gate157( .a(N679), .O(N1471) );
inv1 gate158( .a(N950), .O(N1474) );
buf1 gate159( .a(N686), .O(N1475) );
buf1 gate160( .a(N702), .O(N1478) );
buf1 gate161( .a(N724), .O(N1481) );
buf1 gate162( .a(N736), .O(N1484) );
buf1 gate163( .a(N749), .O(N1487) );
buf1 gate164( .a(N763), .O(N1490) );
buf1 gate165( .a(N877), .O(N1493) );
buf1 gate166( .a(N877), .O(N1496) );
buf1 gate167( .a(N880), .O(N1499) );
buf1 gate168( .a(N880), .O(N1502) );

  xor2  gate4344(.a(N1250), .b(N702), .O(gate169inter0));
  nand2 gate4345(.a(gate169inter0), .b(s_382), .O(gate169inter1));
  and2  gate4346(.a(N1250), .b(N702), .O(gate169inter2));
  inv1  gate4347(.a(s_382), .O(gate169inter3));
  inv1  gate4348(.a(s_383), .O(gate169inter4));
  nand2 gate4349(.a(gate169inter4), .b(gate169inter3), .O(gate169inter5));
  nor2  gate4350(.a(gate169inter5), .b(gate169inter2), .O(gate169inter6));
  inv1  gate4351(.a(N702), .O(gate169inter7));
  inv1  gate4352(.a(N1250), .O(gate169inter8));
  nand2 gate4353(.a(gate169inter8), .b(gate169inter7), .O(gate169inter9));
  nand2 gate4354(.a(s_383), .b(gate169inter3), .O(gate169inter10));
  nor2  gate4355(.a(gate169inter10), .b(gate169inter9), .O(gate169inter11));
  nor2  gate4356(.a(gate169inter11), .b(gate169inter6), .O(gate169inter12));
  nand2 gate4357(.a(gate169inter12), .b(gate169inter1), .O(N1505));
and4 gate170( .a(N1251), .b(N1252), .c(N1253), .d(N1254), .O(N1507) );
and4 gate171( .a(N1255), .b(N1256), .c(N1257), .d(N1258), .O(N1508) );
nand2 gate172( .a(N929), .b(N1259), .O(N1509) );

  xor2  gate1936(.a(N1260), .b(N926), .O(gate173inter0));
  nand2 gate1937(.a(gate173inter0), .b(s_38), .O(gate173inter1));
  and2  gate1938(.a(N1260), .b(N926), .O(gate173inter2));
  inv1  gate1939(.a(s_38), .O(gate173inter3));
  inv1  gate1940(.a(s_39), .O(gate173inter4));
  nand2 gate1941(.a(gate173inter4), .b(gate173inter3), .O(gate173inter5));
  nor2  gate1942(.a(gate173inter5), .b(gate173inter2), .O(gate173inter6));
  inv1  gate1943(.a(N926), .O(gate173inter7));
  inv1  gate1944(.a(N1260), .O(gate173inter8));
  nand2 gate1945(.a(gate173inter8), .b(gate173inter7), .O(gate173inter9));
  nand2 gate1946(.a(s_39), .b(gate173inter3), .O(gate173inter10));
  nor2  gate1947(.a(gate173inter10), .b(gate173inter9), .O(gate173inter11));
  nor2  gate1948(.a(gate173inter11), .b(gate173inter6), .O(gate173inter12));
  nand2 gate1949(.a(gate173inter12), .b(gate173inter1), .O(N1510));

  xor2  gate2972(.a(N1261), .b(N935), .O(gate174inter0));
  nand2 gate2973(.a(gate174inter0), .b(s_186), .O(gate174inter1));
  and2  gate2974(.a(N1261), .b(N935), .O(gate174inter2));
  inv1  gate2975(.a(s_186), .O(gate174inter3));
  inv1  gate2976(.a(s_187), .O(gate174inter4));
  nand2 gate2977(.a(gate174inter4), .b(gate174inter3), .O(gate174inter5));
  nor2  gate2978(.a(gate174inter5), .b(gate174inter2), .O(gate174inter6));
  inv1  gate2979(.a(N935), .O(gate174inter7));
  inv1  gate2980(.a(N1261), .O(gate174inter8));
  nand2 gate2981(.a(gate174inter8), .b(gate174inter7), .O(gate174inter9));
  nand2 gate2982(.a(s_187), .b(gate174inter3), .O(gate174inter10));
  nor2  gate2983(.a(gate174inter10), .b(gate174inter9), .O(gate174inter11));
  nor2  gate2984(.a(gate174inter11), .b(gate174inter6), .O(gate174inter12));
  nand2 gate2985(.a(gate174inter12), .b(gate174inter1), .O(N1511));

  xor2  gate2272(.a(N1262), .b(N932), .O(gate175inter0));
  nand2 gate2273(.a(gate175inter0), .b(s_86), .O(gate175inter1));
  and2  gate2274(.a(N1262), .b(N932), .O(gate175inter2));
  inv1  gate2275(.a(s_86), .O(gate175inter3));
  inv1  gate2276(.a(s_87), .O(gate175inter4));
  nand2 gate2277(.a(gate175inter4), .b(gate175inter3), .O(gate175inter5));
  nor2  gate2278(.a(gate175inter5), .b(gate175inter2), .O(gate175inter6));
  inv1  gate2279(.a(N932), .O(gate175inter7));
  inv1  gate2280(.a(N1262), .O(gate175inter8));
  nand2 gate2281(.a(gate175inter8), .b(gate175inter7), .O(gate175inter9));
  nand2 gate2282(.a(s_87), .b(gate175inter3), .O(gate175inter10));
  nor2  gate2283(.a(gate175inter10), .b(gate175inter9), .O(gate175inter11));
  nor2  gate2284(.a(gate175inter11), .b(gate175inter6), .O(gate175inter12));
  nand2 gate2285(.a(gate175inter12), .b(gate175inter1), .O(N1512));
and2 gate176( .a(N655), .b(N1263), .O(N1520) );
and2 gate177( .a(N874), .b(N1337), .O(N1562) );
inv1 gate178( .a(N1117), .O(N1579) );
and2 gate179( .a(N803), .b(N1117), .O(N1580) );
and2 gate180( .a(N1338), .b(N1345), .O(N1581) );
inv1 gate181( .a(N1117), .O(N1582) );
and2 gate182( .a(N803), .b(N1117), .O(N1583) );
inv1 gate183( .a(N1117), .O(N1584) );
and2 gate184( .a(N803), .b(N1117), .O(N1585) );
and2 gate185( .a(N854), .b(N1347), .O(N1586) );
inv1 gate186( .a(N1117), .O(N1587) );
and2 gate187( .a(N803), .b(N1117), .O(N1588) );
and2 gate188( .a(N77), .b(N1348), .O(N1589) );
inv1 gate189( .a(N1117), .O(N1590) );
and2 gate190( .a(N803), .b(N1117), .O(N1591) );
and2 gate191( .a(N1343), .b(N1349), .O(N1592) );
inv1 gate192( .a(N1117), .O(N1593) );
and2 gate193( .a(N803), .b(N1117), .O(N1594) );
inv1 gate194( .a(N1117), .O(N1595) );
and2 gate195( .a(N803), .b(N1117), .O(N1596) );
and2 gate196( .a(N870), .b(N1351), .O(N1597) );
inv1 gate197( .a(N1117), .O(N1598) );
and2 gate198( .a(N803), .b(N1117), .O(N1599) );
and2 gate199( .a(N116), .b(N1352), .O(N1600) );
and2 gate200( .a(N222), .b(N1401), .O(N1643) );
and2 gate201( .a(N223), .b(N1402), .O(N1644) );
and2 gate202( .a(N226), .b(N1403), .O(N1645) );
and2 gate203( .a(N232), .b(N1404), .O(N1646) );
and2 gate204( .a(N238), .b(N1405), .O(N1647) );
and2 gate205( .a(N244), .b(N1406), .O(N1648) );
and2 gate206( .a(N250), .b(N1407), .O(N1649) );
and2 gate207( .a(N257), .b(N1408), .O(N1650) );
and3 gate208( .a(N1), .b(N13), .c(N1426), .O(N1667) );
and3 gate209( .a(N1), .b(N13), .c(N1427), .O(N1670) );
inv1 gate210( .a(N1202), .O(N1673) );
inv1 gate211( .a(N1202), .O(N1674) );
inv1 gate212( .a(N1202), .O(N1675) );
inv1 gate213( .a(N1202), .O(N1676) );
inv1 gate214( .a(N1202), .O(N1677) );
inv1 gate215( .a(N1202), .O(N1678) );
inv1 gate216( .a(N1202), .O(N1679) );
inv1 gate217( .a(N1202), .O(N1680) );
nand2 gate218( .a(N941), .b(N1467), .O(N1691) );

  xor2  gate4078(.a(N1468), .b(N938), .O(gate219inter0));
  nand2 gate4079(.a(gate219inter0), .b(s_344), .O(gate219inter1));
  and2  gate4080(.a(N1468), .b(N938), .O(gate219inter2));
  inv1  gate4081(.a(s_344), .O(gate219inter3));
  inv1  gate4082(.a(s_345), .O(gate219inter4));
  nand2 gate4083(.a(gate219inter4), .b(gate219inter3), .O(gate219inter5));
  nor2  gate4084(.a(gate219inter5), .b(gate219inter2), .O(gate219inter6));
  inv1  gate4085(.a(N938), .O(gate219inter7));
  inv1  gate4086(.a(N1468), .O(gate219inter8));
  nand2 gate4087(.a(gate219inter8), .b(gate219inter7), .O(gate219inter9));
  nand2 gate4088(.a(s_345), .b(gate219inter3), .O(gate219inter10));
  nor2  gate4089(.a(gate219inter10), .b(gate219inter9), .O(gate219inter11));
  nor2  gate4090(.a(gate219inter11), .b(gate219inter6), .O(gate219inter12));
  nand2 gate4091(.a(gate219inter12), .b(gate219inter1), .O(N1692));

  xor2  gate3490(.a(N1469), .b(N947), .O(gate220inter0));
  nand2 gate3491(.a(gate220inter0), .b(s_260), .O(gate220inter1));
  and2  gate3492(.a(N1469), .b(N947), .O(gate220inter2));
  inv1  gate3493(.a(s_260), .O(gate220inter3));
  inv1  gate3494(.a(s_261), .O(gate220inter4));
  nand2 gate3495(.a(gate220inter4), .b(gate220inter3), .O(gate220inter5));
  nor2  gate3496(.a(gate220inter5), .b(gate220inter2), .O(gate220inter6));
  inv1  gate3497(.a(N947), .O(gate220inter7));
  inv1  gate3498(.a(N1469), .O(gate220inter8));
  nand2 gate3499(.a(gate220inter8), .b(gate220inter7), .O(gate220inter9));
  nand2 gate3500(.a(s_261), .b(gate220inter3), .O(gate220inter10));
  nor2  gate3501(.a(gate220inter10), .b(gate220inter9), .O(gate220inter11));
  nor2  gate3502(.a(gate220inter11), .b(gate220inter6), .O(gate220inter12));
  nand2 gate3503(.a(gate220inter12), .b(gate220inter1), .O(N1693));

  xor2  gate3476(.a(N1470), .b(N944), .O(gate221inter0));
  nand2 gate3477(.a(gate221inter0), .b(s_258), .O(gate221inter1));
  and2  gate3478(.a(N1470), .b(N944), .O(gate221inter2));
  inv1  gate3479(.a(s_258), .O(gate221inter3));
  inv1  gate3480(.a(s_259), .O(gate221inter4));
  nand2 gate3481(.a(gate221inter4), .b(gate221inter3), .O(gate221inter5));
  nor2  gate3482(.a(gate221inter5), .b(gate221inter2), .O(gate221inter6));
  inv1  gate3483(.a(N944), .O(gate221inter7));
  inv1  gate3484(.a(N1470), .O(gate221inter8));
  nand2 gate3485(.a(gate221inter8), .b(gate221inter7), .O(gate221inter9));
  nand2 gate3486(.a(s_259), .b(gate221inter3), .O(gate221inter10));
  nor2  gate3487(.a(gate221inter10), .b(gate221inter9), .O(gate221inter11));
  nor2  gate3488(.a(gate221inter11), .b(gate221inter6), .O(gate221inter12));
  nand2 gate3489(.a(gate221inter12), .b(gate221inter1), .O(N1694));
inv1 gate222( .a(N1505), .O(N1713) );
and2 gate223( .a(N87), .b(N1264), .O(N1714) );
nand2 gate224( .a(N1509), .b(N1510), .O(N1715) );
nand2 gate225( .a(N1511), .b(N1512), .O(N1718) );

  xor2  gate1754(.a(N1508), .b(N1507), .O(gate226inter0));
  nand2 gate1755(.a(gate226inter0), .b(s_12), .O(gate226inter1));
  and2  gate1756(.a(N1508), .b(N1507), .O(gate226inter2));
  inv1  gate1757(.a(s_12), .O(gate226inter3));
  inv1  gate1758(.a(s_13), .O(gate226inter4));
  nand2 gate1759(.a(gate226inter4), .b(gate226inter3), .O(gate226inter5));
  nor2  gate1760(.a(gate226inter5), .b(gate226inter2), .O(gate226inter6));
  inv1  gate1761(.a(N1507), .O(gate226inter7));
  inv1  gate1762(.a(N1508), .O(gate226inter8));
  nand2 gate1763(.a(gate226inter8), .b(gate226inter7), .O(gate226inter9));
  nand2 gate1764(.a(s_13), .b(gate226inter3), .O(gate226inter10));
  nor2  gate1765(.a(gate226inter10), .b(gate226inter9), .O(gate226inter11));
  nor2  gate1766(.a(gate226inter11), .b(gate226inter6), .O(gate226inter12));
  nand2 gate1767(.a(gate226inter12), .b(gate226inter1), .O(N1721));
and2 gate227( .a(N763), .b(N1340), .O(N1722) );

  xor2  gate3084(.a(N1340), .b(N763), .O(gate228inter0));
  nand2 gate3085(.a(gate228inter0), .b(s_202), .O(gate228inter1));
  and2  gate3086(.a(N1340), .b(N763), .O(gate228inter2));
  inv1  gate3087(.a(s_202), .O(gate228inter3));
  inv1  gate3088(.a(s_203), .O(gate228inter4));
  nand2 gate3089(.a(gate228inter4), .b(gate228inter3), .O(gate228inter5));
  nor2  gate3090(.a(gate228inter5), .b(gate228inter2), .O(gate228inter6));
  inv1  gate3091(.a(N763), .O(gate228inter7));
  inv1  gate3092(.a(N1340), .O(gate228inter8));
  nand2 gate3093(.a(gate228inter8), .b(gate228inter7), .O(gate228inter9));
  nand2 gate3094(.a(s_203), .b(gate228inter3), .O(gate228inter10));
  nor2  gate3095(.a(gate228inter10), .b(gate228inter9), .O(gate228inter11));
  nor2  gate3096(.a(gate228inter11), .b(gate228inter6), .O(gate228inter12));
  nand2 gate3097(.a(gate228inter12), .b(gate228inter1), .O(N1725));
inv1 gate229( .a(N1268), .O(N1726) );

  xor2  gate4148(.a(N1271), .b(N1493), .O(gate230inter0));
  nand2 gate4149(.a(gate230inter0), .b(s_354), .O(gate230inter1));
  and2  gate4150(.a(N1271), .b(N1493), .O(gate230inter2));
  inv1  gate4151(.a(s_354), .O(gate230inter3));
  inv1  gate4152(.a(s_355), .O(gate230inter4));
  nand2 gate4153(.a(gate230inter4), .b(gate230inter3), .O(gate230inter5));
  nor2  gate4154(.a(gate230inter5), .b(gate230inter2), .O(gate230inter6));
  inv1  gate4155(.a(N1493), .O(gate230inter7));
  inv1  gate4156(.a(N1271), .O(gate230inter8));
  nand2 gate4157(.a(gate230inter8), .b(gate230inter7), .O(gate230inter9));
  nand2 gate4158(.a(s_355), .b(gate230inter3), .O(gate230inter10));
  nor2  gate4159(.a(gate230inter10), .b(gate230inter9), .O(gate230inter11));
  nor2  gate4160(.a(gate230inter11), .b(gate230inter6), .O(gate230inter12));
  nand2 gate4161(.a(gate230inter12), .b(gate230inter1), .O(N1727));
inv1 gate231( .a(N1493), .O(N1728) );
and2 gate232( .a(N683), .b(N1268), .O(N1729) );

  xor2  gate1740(.a(N1272), .b(N1499), .O(gate233inter0));
  nand2 gate1741(.a(gate233inter0), .b(s_10), .O(gate233inter1));
  and2  gate1742(.a(N1272), .b(N1499), .O(gate233inter2));
  inv1  gate1743(.a(s_10), .O(gate233inter3));
  inv1  gate1744(.a(s_11), .O(gate233inter4));
  nand2 gate1745(.a(gate233inter4), .b(gate233inter3), .O(gate233inter5));
  nor2  gate1746(.a(gate233inter5), .b(gate233inter2), .O(gate233inter6));
  inv1  gate1747(.a(N1499), .O(gate233inter7));
  inv1  gate1748(.a(N1272), .O(gate233inter8));
  nand2 gate1749(.a(gate233inter8), .b(gate233inter7), .O(gate233inter9));
  nand2 gate1750(.a(s_11), .b(gate233inter3), .O(gate233inter10));
  nor2  gate1751(.a(gate233inter10), .b(gate233inter9), .O(gate233inter11));
  nor2  gate1752(.a(gate233inter11), .b(gate233inter6), .O(gate233inter12));
  nand2 gate1753(.a(gate233inter12), .b(gate233inter1), .O(N1730));
inv1 gate234( .a(N1499), .O(N1731) );

  xor2  gate1670(.a(N1264), .b(N87), .O(gate235inter0));
  nand2 gate1671(.a(gate235inter0), .b(s_0), .O(gate235inter1));
  and2  gate1672(.a(N1264), .b(N87), .O(gate235inter2));
  inv1  gate1673(.a(s_0), .O(gate235inter3));
  inv1  gate1674(.a(s_1), .O(gate235inter4));
  nand2 gate1675(.a(gate235inter4), .b(gate235inter3), .O(gate235inter5));
  nor2  gate1676(.a(gate235inter5), .b(gate235inter2), .O(gate235inter6));
  inv1  gate1677(.a(N87), .O(gate235inter7));
  inv1  gate1678(.a(N1264), .O(gate235inter8));
  nand2 gate1679(.a(gate235inter8), .b(gate235inter7), .O(gate235inter9));
  nand2 gate1680(.a(s_1), .b(gate235inter3), .O(gate235inter10));
  nor2  gate1681(.a(gate235inter10), .b(gate235inter9), .O(gate235inter11));
  nor2  gate1682(.a(gate235inter11), .b(gate235inter6), .O(gate235inter12));
  nand2 gate1683(.a(gate235inter12), .b(gate235inter1), .O(N1735));
inv1 gate236( .a(N1273), .O(N1736) );
inv1 gate237( .a(N1276), .O(N1737) );

  xor2  gate3266(.a(N821), .b(N1325), .O(gate238inter0));
  nand2 gate3267(.a(gate238inter0), .b(s_228), .O(gate238inter1));
  and2  gate3268(.a(N821), .b(N1325), .O(gate238inter2));
  inv1  gate3269(.a(s_228), .O(gate238inter3));
  inv1  gate3270(.a(s_229), .O(gate238inter4));
  nand2 gate3271(.a(gate238inter4), .b(gate238inter3), .O(gate238inter5));
  nor2  gate3272(.a(gate238inter5), .b(gate238inter2), .O(gate238inter6));
  inv1  gate3273(.a(N1325), .O(gate238inter7));
  inv1  gate3274(.a(N821), .O(gate238inter8));
  nand2 gate3275(.a(gate238inter8), .b(gate238inter7), .O(gate238inter9));
  nand2 gate3276(.a(s_229), .b(gate238inter3), .O(gate238inter10));
  nor2  gate3277(.a(gate238inter10), .b(gate238inter9), .O(gate238inter11));
  nor2  gate3278(.a(gate238inter11), .b(gate238inter6), .O(gate238inter12));
  nand2 gate3279(.a(gate238inter12), .b(gate238inter1), .O(N1738));
nand2 gate239( .a(N1325), .b(N825), .O(N1747) );
nand3 gate240( .a(N772), .b(N1279), .c(N798), .O(N1756) );
nand4 gate241( .a(N772), .b(N786), .c(N798), .d(N1302), .O(N1761) );
nand2 gate242( .a(N1496), .b(N1339), .O(N1764) );
inv1 gate243( .a(N1496), .O(N1765) );

  xor2  gate3112(.a(N1344), .b(N1502), .O(gate244inter0));
  nand2 gate3113(.a(gate244inter0), .b(s_206), .O(gate244inter1));
  and2  gate3114(.a(N1344), .b(N1502), .O(gate244inter2));
  inv1  gate3115(.a(s_206), .O(gate244inter3));
  inv1  gate3116(.a(s_207), .O(gate244inter4));
  nand2 gate3117(.a(gate244inter4), .b(gate244inter3), .O(gate244inter5));
  nor2  gate3118(.a(gate244inter5), .b(gate244inter2), .O(gate244inter6));
  inv1  gate3119(.a(N1502), .O(gate244inter7));
  inv1  gate3120(.a(N1344), .O(gate244inter8));
  nand2 gate3121(.a(gate244inter8), .b(gate244inter7), .O(gate244inter9));
  nand2 gate3122(.a(s_207), .b(gate244inter3), .O(gate244inter10));
  nor2  gate3123(.a(gate244inter10), .b(gate244inter9), .O(gate244inter11));
  nor2  gate3124(.a(gate244inter11), .b(gate244inter6), .O(gate244inter12));
  nand2 gate3125(.a(gate244inter12), .b(gate244inter1), .O(N1766));
inv1 gate245( .a(N1502), .O(N1767) );
inv1 gate246( .a(N1328), .O(N1768) );
inv1 gate247( .a(N1334), .O(N1769) );
inv1 gate248( .a(N1331), .O(N1770) );
and2 gate249( .a(N845), .b(N1579), .O(N1787) );
and2 gate250( .a(N150), .b(N1580), .O(N1788) );
and2 gate251( .a(N851), .b(N1582), .O(N1789) );
and2 gate252( .a(N159), .b(N1583), .O(N1790) );
and2 gate253( .a(N77), .b(N1584), .O(N1791) );
and2 gate254( .a(N50), .b(N1585), .O(N1792) );
and2 gate255( .a(N858), .b(N1587), .O(N1793) );
and2 gate256( .a(N845), .b(N1588), .O(N1794) );
and2 gate257( .a(N864), .b(N1590), .O(N1795) );
and2 gate258( .a(N851), .b(N1591), .O(N1796) );
and2 gate259( .a(N107), .b(N1593), .O(N1797) );
and2 gate260( .a(N77), .b(N1594), .O(N1798) );
and2 gate261( .a(N116), .b(N1595), .O(N1799) );
and2 gate262( .a(N858), .b(N1596), .O(N1800) );
and2 gate263( .a(N283), .b(N1598), .O(N1801) );
and2 gate264( .a(N864), .b(N1599), .O(N1802) );
and2 gate265( .a(N200), .b(N1363), .O(N1803) );
and2 gate266( .a(N889), .b(N1363), .O(N1806) );
and2 gate267( .a(N890), .b(N1366), .O(N1809) );
and2 gate268( .a(N891), .b(N1366), .O(N1812) );

  xor2  gate2104(.a(N1302), .b(N1298), .O(gate269inter0));
  nand2 gate2105(.a(gate269inter0), .b(s_62), .O(gate269inter1));
  and2  gate2106(.a(N1302), .b(N1298), .O(gate269inter2));
  inv1  gate2107(.a(s_62), .O(gate269inter3));
  inv1  gate2108(.a(s_63), .O(gate269inter4));
  nand2 gate2109(.a(gate269inter4), .b(gate269inter3), .O(gate269inter5));
  nor2  gate2110(.a(gate269inter5), .b(gate269inter2), .O(gate269inter6));
  inv1  gate2111(.a(N1298), .O(gate269inter7));
  inv1  gate2112(.a(N1302), .O(gate269inter8));
  nand2 gate2113(.a(gate269inter8), .b(gate269inter7), .O(gate269inter9));
  nand2 gate2114(.a(s_63), .b(gate269inter3), .O(gate269inter10));
  nor2  gate2115(.a(gate269inter10), .b(gate269inter9), .O(gate269inter11));
  nor2  gate2116(.a(gate269inter11), .b(gate269inter6), .O(gate269inter12));
  nand2 gate2117(.a(gate269inter12), .b(gate269inter1), .O(N1815));
nand2 gate270( .a(N821), .b(N1302), .O(N1818) );
nand3 gate271( .a(N772), .b(N1279), .c(N1179), .O(N1821) );
nand3 gate272( .a(N786), .b(N794), .c(N1298), .O(N1824) );

  xor2  gate2342(.a(N1298), .b(N786), .O(gate273inter0));
  nand2 gate2343(.a(gate273inter0), .b(s_96), .O(gate273inter1));
  and2  gate2344(.a(N1298), .b(N786), .O(gate273inter2));
  inv1  gate2345(.a(s_96), .O(gate273inter3));
  inv1  gate2346(.a(s_97), .O(gate273inter4));
  nand2 gate2347(.a(gate273inter4), .b(gate273inter3), .O(gate273inter5));
  nor2  gate2348(.a(gate273inter5), .b(gate273inter2), .O(gate273inter6));
  inv1  gate2349(.a(N786), .O(gate273inter7));
  inv1  gate2350(.a(N1298), .O(gate273inter8));
  nand2 gate2351(.a(gate273inter8), .b(gate273inter7), .O(gate273inter9));
  nand2 gate2352(.a(s_97), .b(gate273inter3), .O(gate273inter10));
  nor2  gate2353(.a(gate273inter10), .b(gate273inter9), .O(gate273inter11));
  nor2  gate2354(.a(gate273inter11), .b(gate273inter6), .O(gate273inter12));
  nand2 gate2355(.a(gate273inter12), .b(gate273inter1), .O(N1833));
inv1 gate274( .a(N1369), .O(N1842) );
inv1 gate275( .a(N1369), .O(N1843) );
inv1 gate276( .a(N1369), .O(N1844) );
inv1 gate277( .a(N1369), .O(N1845) );
inv1 gate278( .a(N1369), .O(N1846) );
inv1 gate279( .a(N1369), .O(N1847) );
inv1 gate280( .a(N1369), .O(N1848) );
inv1 gate281( .a(N1384), .O(N1849) );
and2 gate282( .a(N1384), .b(N896), .O(N1850) );
inv1 gate283( .a(N1384), .O(N1851) );
and2 gate284( .a(N1384), .b(N896), .O(N1852) );
inv1 gate285( .a(N1384), .O(N1853) );
and2 gate286( .a(N1384), .b(N896), .O(N1854) );
inv1 gate287( .a(N1384), .O(N1855) );
and2 gate288( .a(N1384), .b(N896), .O(N1856) );
inv1 gate289( .a(N1384), .O(N1857) );
and2 gate290( .a(N1384), .b(N896), .O(N1858) );
inv1 gate291( .a(N1384), .O(N1859) );
and2 gate292( .a(N1384), .b(N896), .O(N1860) );
inv1 gate293( .a(N1384), .O(N1861) );
and2 gate294( .a(N1384), .b(N896), .O(N1862) );
inv1 gate295( .a(N1384), .O(N1863) );
and2 gate296( .a(N1384), .b(N896), .O(N1864) );
and2 gate297( .a(N1202), .b(N1409), .O(N1869) );

  xor2  gate1824(.a(N1409), .b(N50), .O(gate298inter0));
  nand2 gate1825(.a(gate298inter0), .b(s_22), .O(gate298inter1));
  and2  gate1826(.a(N1409), .b(N50), .O(gate298inter2));
  inv1  gate1827(.a(s_22), .O(gate298inter3));
  inv1  gate1828(.a(s_23), .O(gate298inter4));
  nand2 gate1829(.a(gate298inter4), .b(gate298inter3), .O(gate298inter5));
  nor2  gate1830(.a(gate298inter5), .b(gate298inter2), .O(gate298inter6));
  inv1  gate1831(.a(N50), .O(gate298inter7));
  inv1  gate1832(.a(N1409), .O(gate298inter8));
  nand2 gate1833(.a(gate298inter8), .b(gate298inter7), .O(gate298inter9));
  nand2 gate1834(.a(s_23), .b(gate298inter3), .O(gate298inter10));
  nor2  gate1835(.a(gate298inter10), .b(gate298inter9), .O(gate298inter11));
  nor2  gate1836(.a(gate298inter11), .b(gate298inter6), .O(gate298inter12));
  nand2 gate1837(.a(gate298inter12), .b(gate298inter1), .O(N1870));
inv1 gate299( .a(N1306), .O(N1873) );
and2 gate300( .a(N1202), .b(N1409), .O(N1874) );

  xor2  gate4330(.a(N1409), .b(N58), .O(gate301inter0));
  nand2 gate4331(.a(gate301inter0), .b(s_380), .O(gate301inter1));
  and2  gate4332(.a(N1409), .b(N58), .O(gate301inter2));
  inv1  gate4333(.a(s_380), .O(gate301inter3));
  inv1  gate4334(.a(s_381), .O(gate301inter4));
  nand2 gate4335(.a(gate301inter4), .b(gate301inter3), .O(gate301inter5));
  nor2  gate4336(.a(gate301inter5), .b(gate301inter2), .O(gate301inter6));
  inv1  gate4337(.a(N58), .O(gate301inter7));
  inv1  gate4338(.a(N1409), .O(gate301inter8));
  nand2 gate4339(.a(gate301inter8), .b(gate301inter7), .O(gate301inter9));
  nand2 gate4340(.a(s_381), .b(gate301inter3), .O(gate301inter10));
  nor2  gate4341(.a(gate301inter10), .b(gate301inter9), .O(gate301inter11));
  nor2  gate4342(.a(gate301inter11), .b(gate301inter6), .O(gate301inter12));
  nand2 gate4343(.a(gate301inter12), .b(gate301inter1), .O(N1875));
inv1 gate302( .a(N1306), .O(N1878) );
and2 gate303( .a(N1202), .b(N1409), .O(N1879) );
nor2 gate304( .a(N68), .b(N1409), .O(N1880) );
inv1 gate305( .a(N1306), .O(N1883) );
and2 gate306( .a(N1202), .b(N1409), .O(N1884) );
nor2 gate307( .a(N77), .b(N1409), .O(N1885) );
inv1 gate308( .a(N1306), .O(N1888) );
and2 gate309( .a(N1202), .b(N1409), .O(N1889) );

  xor2  gate3042(.a(N1409), .b(N87), .O(gate310inter0));
  nand2 gate3043(.a(gate310inter0), .b(s_196), .O(gate310inter1));
  and2  gate3044(.a(N1409), .b(N87), .O(gate310inter2));
  inv1  gate3045(.a(s_196), .O(gate310inter3));
  inv1  gate3046(.a(s_197), .O(gate310inter4));
  nand2 gate3047(.a(gate310inter4), .b(gate310inter3), .O(gate310inter5));
  nor2  gate3048(.a(gate310inter5), .b(gate310inter2), .O(gate310inter6));
  inv1  gate3049(.a(N87), .O(gate310inter7));
  inv1  gate3050(.a(N1409), .O(gate310inter8));
  nand2 gate3051(.a(gate310inter8), .b(gate310inter7), .O(gate310inter9));
  nand2 gate3052(.a(s_197), .b(gate310inter3), .O(gate310inter10));
  nor2  gate3053(.a(gate310inter10), .b(gate310inter9), .O(gate310inter11));
  nor2  gate3054(.a(gate310inter11), .b(gate310inter6), .O(gate310inter12));
  nand2 gate3055(.a(gate310inter12), .b(gate310inter1), .O(N1890));
inv1 gate311( .a(N1322), .O(N1893) );
and2 gate312( .a(N1202), .b(N1409), .O(N1894) );
nor2 gate313( .a(N97), .b(N1409), .O(N1895) );
inv1 gate314( .a(N1315), .O(N1898) );
and2 gate315( .a(N1202), .b(N1409), .O(N1899) );

  xor2  gate2426(.a(N1409), .b(N107), .O(gate316inter0));
  nand2 gate2427(.a(gate316inter0), .b(s_108), .O(gate316inter1));
  and2  gate2428(.a(N1409), .b(N107), .O(gate316inter2));
  inv1  gate2429(.a(s_108), .O(gate316inter3));
  inv1  gate2430(.a(s_109), .O(gate316inter4));
  nand2 gate2431(.a(gate316inter4), .b(gate316inter3), .O(gate316inter5));
  nor2  gate2432(.a(gate316inter5), .b(gate316inter2), .O(gate316inter6));
  inv1  gate2433(.a(N107), .O(gate316inter7));
  inv1  gate2434(.a(N1409), .O(gate316inter8));
  nand2 gate2435(.a(gate316inter8), .b(gate316inter7), .O(gate316inter9));
  nand2 gate2436(.a(s_109), .b(gate316inter3), .O(gate316inter10));
  nor2  gate2437(.a(gate316inter10), .b(gate316inter9), .O(gate316inter11));
  nor2  gate2438(.a(gate316inter11), .b(gate316inter6), .O(gate316inter12));
  nand2 gate2439(.a(gate316inter12), .b(gate316inter1), .O(N1900));
inv1 gate317( .a(N1315), .O(N1903) );
and2 gate318( .a(N1202), .b(N1409), .O(N1904) );
nor2 gate319( .a(N116), .b(N1409), .O(N1905) );
inv1 gate320( .a(N1315), .O(N1908) );
and2 gate321( .a(N1452), .b(N213), .O(N1909) );
nand2 gate322( .a(N1452), .b(N213), .O(N1912) );
and3 gate323( .a(N1452), .b(N213), .c(N343), .O(N1913) );
nand3 gate324( .a(N1452), .b(N213), .c(N343), .O(N1917) );
and3 gate325( .a(N1452), .b(N213), .c(N343), .O(N1922) );
nand3 gate326( .a(N1452), .b(N213), .c(N343), .O(N1926) );
buf1 gate327( .a(N1464), .O(N1930) );

  xor2  gate3000(.a(N1692), .b(N1691), .O(gate328inter0));
  nand2 gate3001(.a(gate328inter0), .b(s_190), .O(gate328inter1));
  and2  gate3002(.a(N1692), .b(N1691), .O(gate328inter2));
  inv1  gate3003(.a(s_190), .O(gate328inter3));
  inv1  gate3004(.a(s_191), .O(gate328inter4));
  nand2 gate3005(.a(gate328inter4), .b(gate328inter3), .O(gate328inter5));
  nor2  gate3006(.a(gate328inter5), .b(gate328inter2), .O(gate328inter6));
  inv1  gate3007(.a(N1691), .O(gate328inter7));
  inv1  gate3008(.a(N1692), .O(gate328inter8));
  nand2 gate3009(.a(gate328inter8), .b(gate328inter7), .O(gate328inter9));
  nand2 gate3010(.a(s_191), .b(gate328inter3), .O(gate328inter10));
  nor2  gate3011(.a(gate328inter10), .b(gate328inter9), .O(gate328inter11));
  nor2  gate3012(.a(gate328inter11), .b(gate328inter6), .O(gate328inter12));
  nand2 gate3013(.a(gate328inter12), .b(gate328inter1), .O(N1933));
nand2 gate329( .a(N1693), .b(N1694), .O(N1936) );
inv1 gate330( .a(N1471), .O(N1939) );

  xor2  gate2664(.a(N1474), .b(N1471), .O(gate331inter0));
  nand2 gate2665(.a(gate331inter0), .b(s_142), .O(gate331inter1));
  and2  gate2666(.a(N1474), .b(N1471), .O(gate331inter2));
  inv1  gate2667(.a(s_142), .O(gate331inter3));
  inv1  gate2668(.a(s_143), .O(gate331inter4));
  nand2 gate2669(.a(gate331inter4), .b(gate331inter3), .O(gate331inter5));
  nor2  gate2670(.a(gate331inter5), .b(gate331inter2), .O(gate331inter6));
  inv1  gate2671(.a(N1471), .O(gate331inter7));
  inv1  gate2672(.a(N1474), .O(gate331inter8));
  nand2 gate2673(.a(gate331inter8), .b(gate331inter7), .O(gate331inter9));
  nand2 gate2674(.a(s_143), .b(gate331inter3), .O(gate331inter10));
  nor2  gate2675(.a(gate331inter10), .b(gate331inter9), .O(gate331inter11));
  nor2  gate2676(.a(gate331inter11), .b(gate331inter6), .O(gate331inter12));
  nand2 gate2677(.a(gate331inter12), .b(gate331inter1), .O(N1940));
inv1 gate332( .a(N1475), .O(N1941) );
inv1 gate333( .a(N1478), .O(N1942) );
inv1 gate334( .a(N1481), .O(N1943) );
inv1 gate335( .a(N1484), .O(N1944) );
inv1 gate336( .a(N1487), .O(N1945) );
inv1 gate337( .a(N1490), .O(N1946) );
inv1 gate338( .a(N1714), .O(N1947) );

  xor2  gate2888(.a(N1728), .b(N953), .O(gate339inter0));
  nand2 gate2889(.a(gate339inter0), .b(s_174), .O(gate339inter1));
  and2  gate2890(.a(N1728), .b(N953), .O(gate339inter2));
  inv1  gate2891(.a(s_174), .O(gate339inter3));
  inv1  gate2892(.a(s_175), .O(gate339inter4));
  nand2 gate2893(.a(gate339inter4), .b(gate339inter3), .O(gate339inter5));
  nor2  gate2894(.a(gate339inter5), .b(gate339inter2), .O(gate339inter6));
  inv1  gate2895(.a(N953), .O(gate339inter7));
  inv1  gate2896(.a(N1728), .O(gate339inter8));
  nand2 gate2897(.a(gate339inter8), .b(gate339inter7), .O(gate339inter9));
  nand2 gate2898(.a(s_175), .b(gate339inter3), .O(gate339inter10));
  nor2  gate2899(.a(gate339inter10), .b(gate339inter9), .O(gate339inter11));
  nor2  gate2900(.a(gate339inter11), .b(gate339inter6), .O(gate339inter12));
  nand2 gate2901(.a(gate339inter12), .b(gate339inter1), .O(N1960));

  xor2  gate4316(.a(N1731), .b(N959), .O(gate340inter0));
  nand2 gate4317(.a(gate340inter0), .b(s_378), .O(gate340inter1));
  and2  gate4318(.a(N1731), .b(N959), .O(gate340inter2));
  inv1  gate4319(.a(s_378), .O(gate340inter3));
  inv1  gate4320(.a(s_379), .O(gate340inter4));
  nand2 gate4321(.a(gate340inter4), .b(gate340inter3), .O(gate340inter5));
  nor2  gate4322(.a(gate340inter5), .b(gate340inter2), .O(gate340inter6));
  inv1  gate4323(.a(N959), .O(gate340inter7));
  inv1  gate4324(.a(N1731), .O(gate340inter8));
  nand2 gate4325(.a(gate340inter8), .b(gate340inter7), .O(gate340inter9));
  nand2 gate4326(.a(s_379), .b(gate340inter3), .O(gate340inter10));
  nor2  gate4327(.a(gate340inter10), .b(gate340inter9), .O(gate340inter11));
  nor2  gate4328(.a(gate340inter11), .b(gate340inter6), .O(gate340inter12));
  nand2 gate4329(.a(gate340inter12), .b(gate340inter1), .O(N1961));
and2 gate341( .a(N1520), .b(N1276), .O(N1966) );

  xor2  gate3882(.a(N1765), .b(N956), .O(gate342inter0));
  nand2 gate3883(.a(gate342inter0), .b(s_316), .O(gate342inter1));
  and2  gate3884(.a(N1765), .b(N956), .O(gate342inter2));
  inv1  gate3885(.a(s_316), .O(gate342inter3));
  inv1  gate3886(.a(s_317), .O(gate342inter4));
  nand2 gate3887(.a(gate342inter4), .b(gate342inter3), .O(gate342inter5));
  nor2  gate3888(.a(gate342inter5), .b(gate342inter2), .O(gate342inter6));
  inv1  gate3889(.a(N956), .O(gate342inter7));
  inv1  gate3890(.a(N1765), .O(gate342inter8));
  nand2 gate3891(.a(gate342inter8), .b(gate342inter7), .O(gate342inter9));
  nand2 gate3892(.a(s_317), .b(gate342inter3), .O(gate342inter10));
  nor2  gate3893(.a(gate342inter10), .b(gate342inter9), .O(gate342inter11));
  nor2  gate3894(.a(gate342inter11), .b(gate342inter6), .O(gate342inter12));
  nand2 gate3895(.a(gate342inter12), .b(gate342inter1), .O(N1981));

  xor2  gate4022(.a(N1767), .b(N962), .O(gate343inter0));
  nand2 gate4023(.a(gate343inter0), .b(s_336), .O(gate343inter1));
  and2  gate4024(.a(N1767), .b(N962), .O(gate343inter2));
  inv1  gate4025(.a(s_336), .O(gate343inter3));
  inv1  gate4026(.a(s_337), .O(gate343inter4));
  nand2 gate4027(.a(gate343inter4), .b(gate343inter3), .O(gate343inter5));
  nor2  gate4028(.a(gate343inter5), .b(gate343inter2), .O(gate343inter6));
  inv1  gate4029(.a(N962), .O(gate343inter7));
  inv1  gate4030(.a(N1767), .O(gate343inter8));
  nand2 gate4031(.a(gate343inter8), .b(gate343inter7), .O(gate343inter9));
  nand2 gate4032(.a(s_337), .b(gate343inter3), .O(gate343inter10));
  nor2  gate4033(.a(gate343inter10), .b(gate343inter9), .O(gate343inter11));
  nor2  gate4034(.a(gate343inter11), .b(gate343inter6), .O(gate343inter12));
  nand2 gate4035(.a(gate343inter12), .b(gate343inter1), .O(N1982));
and2 gate344( .a(N1067), .b(N1768), .O(N1983) );
or3 gate345( .a(N1581), .b(N1787), .c(N1788), .O(N1986) );
or3 gate346( .a(N1586), .b(N1791), .c(N1792), .O(N1987) );
or3 gate347( .a(N1589), .b(N1793), .c(N1794), .O(N1988) );
or3 gate348( .a(N1592), .b(N1795), .c(N1796), .O(N1989) );
or3 gate349( .a(N1597), .b(N1799), .c(N1800), .O(N1990) );
or3 gate350( .a(N1600), .b(N1801), .c(N1802), .O(N1991) );
and2 gate351( .a(N77), .b(N1849), .O(N2022) );
and2 gate352( .a(N223), .b(N1850), .O(N2023) );
and2 gate353( .a(N87), .b(N1851), .O(N2024) );
and2 gate354( .a(N226), .b(N1852), .O(N2025) );
and2 gate355( .a(N97), .b(N1853), .O(N2026) );
and2 gate356( .a(N232), .b(N1854), .O(N2027) );
and2 gate357( .a(N107), .b(N1855), .O(N2028) );
and2 gate358( .a(N238), .b(N1856), .O(N2029) );
and2 gate359( .a(N116), .b(N1857), .O(N2030) );
and2 gate360( .a(N244), .b(N1858), .O(N2031) );
and2 gate361( .a(N283), .b(N1859), .O(N2032) );
and2 gate362( .a(N250), .b(N1860), .O(N2033) );
and2 gate363( .a(N294), .b(N1861), .O(N2034) );
and2 gate364( .a(N257), .b(N1862), .O(N2035) );
and2 gate365( .a(N303), .b(N1863), .O(N2036) );
and2 gate366( .a(N264), .b(N1864), .O(N2037) );
buf1 gate367( .a(N1667), .O(N2038) );
inv1 gate368( .a(N1667), .O(N2043) );
buf1 gate369( .a(N1670), .O(N2052) );
inv1 gate370( .a(N1670), .O(N2057) );
and3 gate371( .a(N50), .b(N1197), .c(N1869), .O(N2068) );
and3 gate372( .a(N58), .b(N1197), .c(N1874), .O(N2073) );
and3 gate373( .a(N68), .b(N1197), .c(N1879), .O(N2078) );
and3 gate374( .a(N77), .b(N1197), .c(N1884), .O(N2083) );
and3 gate375( .a(N87), .b(N1219), .c(N1889), .O(N2088) );
and3 gate376( .a(N97), .b(N1219), .c(N1894), .O(N2093) );
and3 gate377( .a(N107), .b(N1219), .c(N1899), .O(N2098) );
and3 gate378( .a(N116), .b(N1219), .c(N1904), .O(N2103) );
inv1 gate379( .a(N1562), .O(N2121) );
inv1 gate380( .a(N1562), .O(N2122) );
inv1 gate381( .a(N1562), .O(N2123) );
inv1 gate382( .a(N1562), .O(N2124) );
inv1 gate383( .a(N1562), .O(N2125) );
inv1 gate384( .a(N1562), .O(N2126) );
inv1 gate385( .a(N1562), .O(N2127) );
inv1 gate386( .a(N1562), .O(N2128) );
nand2 gate387( .a(N950), .b(N1939), .O(N2133) );

  xor2  gate1684(.a(N1941), .b(N1478), .O(gate388inter0));
  nand2 gate1685(.a(gate388inter0), .b(s_2), .O(gate388inter1));
  and2  gate1686(.a(N1941), .b(N1478), .O(gate388inter2));
  inv1  gate1687(.a(s_2), .O(gate388inter3));
  inv1  gate1688(.a(s_3), .O(gate388inter4));
  nand2 gate1689(.a(gate388inter4), .b(gate388inter3), .O(gate388inter5));
  nor2  gate1690(.a(gate388inter5), .b(gate388inter2), .O(gate388inter6));
  inv1  gate1691(.a(N1478), .O(gate388inter7));
  inv1  gate1692(.a(N1941), .O(gate388inter8));
  nand2 gate1693(.a(gate388inter8), .b(gate388inter7), .O(gate388inter9));
  nand2 gate1694(.a(s_3), .b(gate388inter3), .O(gate388inter10));
  nor2  gate1695(.a(gate388inter10), .b(gate388inter9), .O(gate388inter11));
  nor2  gate1696(.a(gate388inter11), .b(gate388inter6), .O(gate388inter12));
  nand2 gate1697(.a(gate388inter12), .b(gate388inter1), .O(N2134));

  xor2  gate1712(.a(N1942), .b(N1475), .O(gate389inter0));
  nand2 gate1713(.a(gate389inter0), .b(s_6), .O(gate389inter1));
  and2  gate1714(.a(N1942), .b(N1475), .O(gate389inter2));
  inv1  gate1715(.a(s_6), .O(gate389inter3));
  inv1  gate1716(.a(s_7), .O(gate389inter4));
  nand2 gate1717(.a(gate389inter4), .b(gate389inter3), .O(gate389inter5));
  nor2  gate1718(.a(gate389inter5), .b(gate389inter2), .O(gate389inter6));
  inv1  gate1719(.a(N1475), .O(gate389inter7));
  inv1  gate1720(.a(N1942), .O(gate389inter8));
  nand2 gate1721(.a(gate389inter8), .b(gate389inter7), .O(gate389inter9));
  nand2 gate1722(.a(s_7), .b(gate389inter3), .O(gate389inter10));
  nor2  gate1723(.a(gate389inter10), .b(gate389inter9), .O(gate389inter11));
  nor2  gate1724(.a(gate389inter11), .b(gate389inter6), .O(gate389inter12));
  nand2 gate1725(.a(gate389inter12), .b(gate389inter1), .O(N2135));

  xor2  gate2860(.a(N1943), .b(N1484), .O(gate390inter0));
  nand2 gate2861(.a(gate390inter0), .b(s_170), .O(gate390inter1));
  and2  gate2862(.a(N1943), .b(N1484), .O(gate390inter2));
  inv1  gate2863(.a(s_170), .O(gate390inter3));
  inv1  gate2864(.a(s_171), .O(gate390inter4));
  nand2 gate2865(.a(gate390inter4), .b(gate390inter3), .O(gate390inter5));
  nor2  gate2866(.a(gate390inter5), .b(gate390inter2), .O(gate390inter6));
  inv1  gate2867(.a(N1484), .O(gate390inter7));
  inv1  gate2868(.a(N1943), .O(gate390inter8));
  nand2 gate2869(.a(gate390inter8), .b(gate390inter7), .O(gate390inter9));
  nand2 gate2870(.a(s_171), .b(gate390inter3), .O(gate390inter10));
  nor2  gate2871(.a(gate390inter10), .b(gate390inter9), .O(gate390inter11));
  nor2  gate2872(.a(gate390inter11), .b(gate390inter6), .O(gate390inter12));
  nand2 gate2873(.a(gate390inter12), .b(gate390inter1), .O(N2136));

  xor2  gate2090(.a(N1944), .b(N1481), .O(gate391inter0));
  nand2 gate2091(.a(gate391inter0), .b(s_60), .O(gate391inter1));
  and2  gate2092(.a(N1944), .b(N1481), .O(gate391inter2));
  inv1  gate2093(.a(s_60), .O(gate391inter3));
  inv1  gate2094(.a(s_61), .O(gate391inter4));
  nand2 gate2095(.a(gate391inter4), .b(gate391inter3), .O(gate391inter5));
  nor2  gate2096(.a(gate391inter5), .b(gate391inter2), .O(gate391inter6));
  inv1  gate2097(.a(N1481), .O(gate391inter7));
  inv1  gate2098(.a(N1944), .O(gate391inter8));
  nand2 gate2099(.a(gate391inter8), .b(gate391inter7), .O(gate391inter9));
  nand2 gate2100(.a(s_61), .b(gate391inter3), .O(gate391inter10));
  nor2  gate2101(.a(gate391inter10), .b(gate391inter9), .O(gate391inter11));
  nor2  gate2102(.a(gate391inter11), .b(gate391inter6), .O(gate391inter12));
  nand2 gate2103(.a(gate391inter12), .b(gate391inter1), .O(N2137));
nand2 gate392( .a(N1490), .b(N1945), .O(N2138) );

  xor2  gate2636(.a(N1946), .b(N1487), .O(gate393inter0));
  nand2 gate2637(.a(gate393inter0), .b(s_138), .O(gate393inter1));
  and2  gate2638(.a(N1946), .b(N1487), .O(gate393inter2));
  inv1  gate2639(.a(s_138), .O(gate393inter3));
  inv1  gate2640(.a(s_139), .O(gate393inter4));
  nand2 gate2641(.a(gate393inter4), .b(gate393inter3), .O(gate393inter5));
  nor2  gate2642(.a(gate393inter5), .b(gate393inter2), .O(gate393inter6));
  inv1  gate2643(.a(N1487), .O(gate393inter7));
  inv1  gate2644(.a(N1946), .O(gate393inter8));
  nand2 gate2645(.a(gate393inter8), .b(gate393inter7), .O(gate393inter9));
  nand2 gate2646(.a(s_139), .b(gate393inter3), .O(gate393inter10));
  nor2  gate2647(.a(gate393inter10), .b(gate393inter9), .O(gate393inter11));
  nor2  gate2648(.a(gate393inter11), .b(gate393inter6), .O(gate393inter12));
  nand2 gate2649(.a(gate393inter12), .b(gate393inter1), .O(N2139));
inv1 gate394( .a(N1933), .O(N2141) );
inv1 gate395( .a(N1936), .O(N2142) );
inv1 gate396( .a(N1738), .O(N2143) );
and2 gate397( .a(N1738), .b(N1747), .O(N2144) );
inv1 gate398( .a(N1747), .O(N2145) );

  xor2  gate2720(.a(N1960), .b(N1727), .O(gate399inter0));
  nand2 gate2721(.a(gate399inter0), .b(s_150), .O(gate399inter1));
  and2  gate2722(.a(N1960), .b(N1727), .O(gate399inter2));
  inv1  gate2723(.a(s_150), .O(gate399inter3));
  inv1  gate2724(.a(s_151), .O(gate399inter4));
  nand2 gate2725(.a(gate399inter4), .b(gate399inter3), .O(gate399inter5));
  nor2  gate2726(.a(gate399inter5), .b(gate399inter2), .O(gate399inter6));
  inv1  gate2727(.a(N1727), .O(gate399inter7));
  inv1  gate2728(.a(N1960), .O(gate399inter8));
  nand2 gate2729(.a(gate399inter8), .b(gate399inter7), .O(gate399inter9));
  nand2 gate2730(.a(s_151), .b(gate399inter3), .O(gate399inter10));
  nor2  gate2731(.a(gate399inter10), .b(gate399inter9), .O(gate399inter11));
  nor2  gate2732(.a(gate399inter11), .b(gate399inter6), .O(gate399inter12));
  nand2 gate2733(.a(gate399inter12), .b(gate399inter1), .O(N2146));

  xor2  gate2804(.a(N1961), .b(N1730), .O(gate400inter0));
  nand2 gate2805(.a(gate400inter0), .b(s_162), .O(gate400inter1));
  and2  gate2806(.a(N1961), .b(N1730), .O(gate400inter2));
  inv1  gate2807(.a(s_162), .O(gate400inter3));
  inv1  gate2808(.a(s_163), .O(gate400inter4));
  nand2 gate2809(.a(gate400inter4), .b(gate400inter3), .O(gate400inter5));
  nor2  gate2810(.a(gate400inter5), .b(gate400inter2), .O(gate400inter6));
  inv1  gate2811(.a(N1730), .O(gate400inter7));
  inv1  gate2812(.a(N1961), .O(gate400inter8));
  nand2 gate2813(.a(gate400inter8), .b(gate400inter7), .O(gate400inter9));
  nand2 gate2814(.a(s_163), .b(gate400inter3), .O(gate400inter10));
  nor2  gate2815(.a(gate400inter10), .b(gate400inter9), .O(gate400inter11));
  nor2  gate2816(.a(gate400inter11), .b(gate400inter6), .O(gate400inter12));
  nand2 gate2817(.a(gate400inter12), .b(gate400inter1), .O(N2147));
and4 gate401( .a(N1722), .b(N1267), .c(N665), .d(N58), .O(N2148) );
inv1 gate402( .a(N1738), .O(N2149) );
and2 gate403( .a(N1738), .b(N1747), .O(N2150) );
inv1 gate404( .a(N1747), .O(N2151) );
inv1 gate405( .a(N1738), .O(N2152) );
inv1 gate406( .a(N1747), .O(N2153) );
and2 gate407( .a(N1738), .b(N1747), .O(N2154) );
inv1 gate408( .a(N1738), .O(N2155) );
inv1 gate409( .a(N1747), .O(N2156) );
and2 gate410( .a(N1738), .b(N1747), .O(N2157) );
buf1 gate411( .a(N1761), .O(N2158) );
buf1 gate412( .a(N1761), .O(N2175) );

  xor2  gate2286(.a(N1981), .b(N1764), .O(gate413inter0));
  nand2 gate2287(.a(gate413inter0), .b(s_88), .O(gate413inter1));
  and2  gate2288(.a(N1981), .b(N1764), .O(gate413inter2));
  inv1  gate2289(.a(s_88), .O(gate413inter3));
  inv1  gate2290(.a(s_89), .O(gate413inter4));
  nand2 gate2291(.a(gate413inter4), .b(gate413inter3), .O(gate413inter5));
  nor2  gate2292(.a(gate413inter5), .b(gate413inter2), .O(gate413inter6));
  inv1  gate2293(.a(N1764), .O(gate413inter7));
  inv1  gate2294(.a(N1981), .O(gate413inter8));
  nand2 gate2295(.a(gate413inter8), .b(gate413inter7), .O(gate413inter9));
  nand2 gate2296(.a(s_89), .b(gate413inter3), .O(gate413inter10));
  nor2  gate2297(.a(gate413inter10), .b(gate413inter9), .O(gate413inter11));
  nor2  gate2298(.a(gate413inter11), .b(gate413inter6), .O(gate413inter12));
  nand2 gate2299(.a(gate413inter12), .b(gate413inter1), .O(N2178));

  xor2  gate2524(.a(N1982), .b(N1766), .O(gate414inter0));
  nand2 gate2525(.a(gate414inter0), .b(s_122), .O(gate414inter1));
  and2  gate2526(.a(N1982), .b(N1766), .O(gate414inter2));
  inv1  gate2527(.a(s_122), .O(gate414inter3));
  inv1  gate2528(.a(s_123), .O(gate414inter4));
  nand2 gate2529(.a(gate414inter4), .b(gate414inter3), .O(gate414inter5));
  nor2  gate2530(.a(gate414inter5), .b(gate414inter2), .O(gate414inter6));
  inv1  gate2531(.a(N1766), .O(gate414inter7));
  inv1  gate2532(.a(N1982), .O(gate414inter8));
  nand2 gate2533(.a(gate414inter8), .b(gate414inter7), .O(gate414inter9));
  nand2 gate2534(.a(s_123), .b(gate414inter3), .O(gate414inter10));
  nor2  gate2535(.a(gate414inter10), .b(gate414inter9), .O(gate414inter11));
  nor2  gate2536(.a(gate414inter11), .b(gate414inter6), .O(gate414inter12));
  nand2 gate2537(.a(gate414inter12), .b(gate414inter1), .O(N2179));
inv1 gate415( .a(N1756), .O(N2180) );
and2 gate416( .a(N1756), .b(N1328), .O(N2181) );
inv1 gate417( .a(N1756), .O(N2183) );
and2 gate418( .a(N1331), .b(N1756), .O(N2184) );

  xor2  gate4036(.a(N1812), .b(N1358), .O(gate419inter0));
  nand2 gate4037(.a(gate419inter0), .b(s_338), .O(gate419inter1));
  and2  gate4038(.a(N1812), .b(N1358), .O(gate419inter2));
  inv1  gate4039(.a(s_338), .O(gate419inter3));
  inv1  gate4040(.a(s_339), .O(gate419inter4));
  nand2 gate4041(.a(gate419inter4), .b(gate419inter3), .O(gate419inter5));
  nor2  gate4042(.a(gate419inter5), .b(gate419inter2), .O(gate419inter6));
  inv1  gate4043(.a(N1358), .O(gate419inter7));
  inv1  gate4044(.a(N1812), .O(gate419inter8));
  nand2 gate4045(.a(gate419inter8), .b(gate419inter7), .O(gate419inter9));
  nand2 gate4046(.a(s_339), .b(gate419inter3), .O(gate419inter10));
  nor2  gate4047(.a(gate419inter10), .b(gate419inter9), .O(gate419inter11));
  nor2  gate4048(.a(gate419inter11), .b(gate419inter6), .O(gate419inter12));
  nand2 gate4049(.a(gate419inter12), .b(gate419inter1), .O(N2185));
nand2 gate420( .a(N1358), .b(N1809), .O(N2188) );
nand2 gate421( .a(N1353), .b(N1812), .O(N2191) );
nand2 gate422( .a(N1353), .b(N1809), .O(N2194) );

  xor2  gate2468(.a(N1806), .b(N1358), .O(gate423inter0));
  nand2 gate2469(.a(gate423inter0), .b(s_114), .O(gate423inter1));
  and2  gate2470(.a(N1806), .b(N1358), .O(gate423inter2));
  inv1  gate2471(.a(s_114), .O(gate423inter3));
  inv1  gate2472(.a(s_115), .O(gate423inter4));
  nand2 gate2473(.a(gate423inter4), .b(gate423inter3), .O(gate423inter5));
  nor2  gate2474(.a(gate423inter5), .b(gate423inter2), .O(gate423inter6));
  inv1  gate2475(.a(N1358), .O(gate423inter7));
  inv1  gate2476(.a(N1806), .O(gate423inter8));
  nand2 gate2477(.a(gate423inter8), .b(gate423inter7), .O(gate423inter9));
  nand2 gate2478(.a(s_115), .b(gate423inter3), .O(gate423inter10));
  nor2  gate2479(.a(gate423inter10), .b(gate423inter9), .O(gate423inter11));
  nor2  gate2480(.a(gate423inter11), .b(gate423inter6), .O(gate423inter12));
  nand2 gate2481(.a(gate423inter12), .b(gate423inter1), .O(N2197));

  xor2  gate3280(.a(N1803), .b(N1358), .O(gate424inter0));
  nand2 gate3281(.a(gate424inter0), .b(s_230), .O(gate424inter1));
  and2  gate3282(.a(N1803), .b(N1358), .O(gate424inter2));
  inv1  gate3283(.a(s_230), .O(gate424inter3));
  inv1  gate3284(.a(s_231), .O(gate424inter4));
  nand2 gate3285(.a(gate424inter4), .b(gate424inter3), .O(gate424inter5));
  nor2  gate3286(.a(gate424inter5), .b(gate424inter2), .O(gate424inter6));
  inv1  gate3287(.a(N1358), .O(gate424inter7));
  inv1  gate3288(.a(N1803), .O(gate424inter8));
  nand2 gate3289(.a(gate424inter8), .b(gate424inter7), .O(gate424inter9));
  nand2 gate3290(.a(s_231), .b(gate424inter3), .O(gate424inter10));
  nor2  gate3291(.a(gate424inter10), .b(gate424inter9), .O(gate424inter11));
  nor2  gate3292(.a(gate424inter11), .b(gate424inter6), .O(gate424inter12));
  nand2 gate3293(.a(gate424inter12), .b(gate424inter1), .O(N2200));

  xor2  gate3714(.a(N1806), .b(N1353), .O(gate425inter0));
  nand2 gate3715(.a(gate425inter0), .b(s_292), .O(gate425inter1));
  and2  gate3716(.a(N1806), .b(N1353), .O(gate425inter2));
  inv1  gate3717(.a(s_292), .O(gate425inter3));
  inv1  gate3718(.a(s_293), .O(gate425inter4));
  nand2 gate3719(.a(gate425inter4), .b(gate425inter3), .O(gate425inter5));
  nor2  gate3720(.a(gate425inter5), .b(gate425inter2), .O(gate425inter6));
  inv1  gate3721(.a(N1353), .O(gate425inter7));
  inv1  gate3722(.a(N1806), .O(gate425inter8));
  nand2 gate3723(.a(gate425inter8), .b(gate425inter7), .O(gate425inter9));
  nand2 gate3724(.a(s_293), .b(gate425inter3), .O(gate425inter10));
  nor2  gate3725(.a(gate425inter10), .b(gate425inter9), .O(gate425inter11));
  nor2  gate3726(.a(gate425inter11), .b(gate425inter6), .O(gate425inter12));
  nand2 gate3727(.a(gate425inter12), .b(gate425inter1), .O(N2203));

  xor2  gate3588(.a(N1803), .b(N1353), .O(gate426inter0));
  nand2 gate3589(.a(gate426inter0), .b(s_274), .O(gate426inter1));
  and2  gate3590(.a(N1803), .b(N1353), .O(gate426inter2));
  inv1  gate3591(.a(s_274), .O(gate426inter3));
  inv1  gate3592(.a(s_275), .O(gate426inter4));
  nand2 gate3593(.a(gate426inter4), .b(gate426inter3), .O(gate426inter5));
  nor2  gate3594(.a(gate426inter5), .b(gate426inter2), .O(gate426inter6));
  inv1  gate3595(.a(N1353), .O(gate426inter7));
  inv1  gate3596(.a(N1803), .O(gate426inter8));
  nand2 gate3597(.a(gate426inter8), .b(gate426inter7), .O(gate426inter9));
  nand2 gate3598(.a(s_275), .b(gate426inter3), .O(gate426inter10));
  nor2  gate3599(.a(gate426inter10), .b(gate426inter9), .O(gate426inter11));
  nor2  gate3600(.a(gate426inter11), .b(gate426inter6), .O(gate426inter12));
  nand2 gate3601(.a(gate426inter12), .b(gate426inter1), .O(N2206));
inv1 gate427( .a(N1815), .O(N2209) );
inv1 gate428( .a(N1818), .O(N2210) );
and2 gate429( .a(N1815), .b(N1818), .O(N2211) );
buf1 gate430( .a(N1821), .O(N2212) );
buf1 gate431( .a(N1821), .O(N2221) );
inv1 gate432( .a(N1833), .O(N2230) );
inv1 gate433( .a(N1833), .O(N2231) );
inv1 gate434( .a(N1833), .O(N2232) );
inv1 gate435( .a(N1833), .O(N2233) );
inv1 gate436( .a(N1824), .O(N2234) );
inv1 gate437( .a(N1824), .O(N2235) );
inv1 gate438( .a(N1824), .O(N2236) );
inv1 gate439( .a(N1824), .O(N2237) );
or3 gate440( .a(N2022), .b(N1643), .c(N2023), .O(N2238) );
or3 gate441( .a(N2024), .b(N1644), .c(N2025), .O(N2239) );
or3 gate442( .a(N2026), .b(N1645), .c(N2027), .O(N2240) );
or3 gate443( .a(N2028), .b(N1646), .c(N2029), .O(N2241) );
or3 gate444( .a(N2030), .b(N1647), .c(N2031), .O(N2242) );
or3 gate445( .a(N2032), .b(N1648), .c(N2033), .O(N2243) );
or3 gate446( .a(N2034), .b(N1649), .c(N2035), .O(N2244) );
or3 gate447( .a(N2036), .b(N1650), .c(N2037), .O(N2245) );
and2 gate448( .a(N1986), .b(N1673), .O(N2270) );
and2 gate449( .a(N1987), .b(N1675), .O(N2277) );
and2 gate450( .a(N1988), .b(N1676), .O(N2282) );
and2 gate451( .a(N1989), .b(N1677), .O(N2287) );
and2 gate452( .a(N1990), .b(N1679), .O(N2294) );
and2 gate453( .a(N1991), .b(N1680), .O(N2299) );
buf1 gate454( .a(N1917), .O(N2304) );
and2 gate455( .a(N1930), .b(N350), .O(N2307) );

  xor2  gate2650(.a(N350), .b(N1930), .O(gate456inter0));
  nand2 gate2651(.a(gate456inter0), .b(s_140), .O(gate456inter1));
  and2  gate2652(.a(N350), .b(N1930), .O(gate456inter2));
  inv1  gate2653(.a(s_140), .O(gate456inter3));
  inv1  gate2654(.a(s_141), .O(gate456inter4));
  nand2 gate2655(.a(gate456inter4), .b(gate456inter3), .O(gate456inter5));
  nor2  gate2656(.a(gate456inter5), .b(gate456inter2), .O(gate456inter6));
  inv1  gate2657(.a(N1930), .O(gate456inter7));
  inv1  gate2658(.a(N350), .O(gate456inter8));
  nand2 gate2659(.a(gate456inter8), .b(gate456inter7), .O(gate456inter9));
  nand2 gate2660(.a(s_141), .b(gate456inter3), .O(gate456inter10));
  nor2  gate2661(.a(gate456inter10), .b(gate456inter9), .O(gate456inter11));
  nor2  gate2662(.a(gate456inter11), .b(gate456inter6), .O(gate456inter12));
  nand2 gate2663(.a(gate456inter12), .b(gate456inter1), .O(N2310));
buf1 gate457( .a(N1715), .O(N2313) );
buf1 gate458( .a(N1718), .O(N2316) );
buf1 gate459( .a(N1715), .O(N2319) );
buf1 gate460( .a(N1718), .O(N2322) );

  xor2  gate3392(.a(N2133), .b(N1940), .O(gate461inter0));
  nand2 gate3393(.a(gate461inter0), .b(s_246), .O(gate461inter1));
  and2  gate3394(.a(N2133), .b(N1940), .O(gate461inter2));
  inv1  gate3395(.a(s_246), .O(gate461inter3));
  inv1  gate3396(.a(s_247), .O(gate461inter4));
  nand2 gate3397(.a(gate461inter4), .b(gate461inter3), .O(gate461inter5));
  nor2  gate3398(.a(gate461inter5), .b(gate461inter2), .O(gate461inter6));
  inv1  gate3399(.a(N1940), .O(gate461inter7));
  inv1  gate3400(.a(N2133), .O(gate461inter8));
  nand2 gate3401(.a(gate461inter8), .b(gate461inter7), .O(gate461inter9));
  nand2 gate3402(.a(s_247), .b(gate461inter3), .O(gate461inter10));
  nor2  gate3403(.a(gate461inter10), .b(gate461inter9), .O(gate461inter11));
  nor2  gate3404(.a(gate461inter11), .b(gate461inter6), .O(gate461inter12));
  nand2 gate3405(.a(gate461inter12), .b(gate461inter1), .O(N2325));

  xor2  gate2454(.a(N2135), .b(N2134), .O(gate462inter0));
  nand2 gate2455(.a(gate462inter0), .b(s_112), .O(gate462inter1));
  and2  gate2456(.a(N2135), .b(N2134), .O(gate462inter2));
  inv1  gate2457(.a(s_112), .O(gate462inter3));
  inv1  gate2458(.a(s_113), .O(gate462inter4));
  nand2 gate2459(.a(gate462inter4), .b(gate462inter3), .O(gate462inter5));
  nor2  gate2460(.a(gate462inter5), .b(gate462inter2), .O(gate462inter6));
  inv1  gate2461(.a(N2134), .O(gate462inter7));
  inv1  gate2462(.a(N2135), .O(gate462inter8));
  nand2 gate2463(.a(gate462inter8), .b(gate462inter7), .O(gate462inter9));
  nand2 gate2464(.a(s_113), .b(gate462inter3), .O(gate462inter10));
  nor2  gate2465(.a(gate462inter10), .b(gate462inter9), .O(gate462inter11));
  nor2  gate2466(.a(gate462inter11), .b(gate462inter6), .O(gate462inter12));
  nand2 gate2467(.a(gate462inter12), .b(gate462inter1), .O(N2328));

  xor2  gate3210(.a(N2137), .b(N2136), .O(gate463inter0));
  nand2 gate3211(.a(gate463inter0), .b(s_220), .O(gate463inter1));
  and2  gate3212(.a(N2137), .b(N2136), .O(gate463inter2));
  inv1  gate3213(.a(s_220), .O(gate463inter3));
  inv1  gate3214(.a(s_221), .O(gate463inter4));
  nand2 gate3215(.a(gate463inter4), .b(gate463inter3), .O(gate463inter5));
  nor2  gate3216(.a(gate463inter5), .b(gate463inter2), .O(gate463inter6));
  inv1  gate3217(.a(N2136), .O(gate463inter7));
  inv1  gate3218(.a(N2137), .O(gate463inter8));
  nand2 gate3219(.a(gate463inter8), .b(gate463inter7), .O(gate463inter9));
  nand2 gate3220(.a(s_221), .b(gate463inter3), .O(gate463inter10));
  nor2  gate3221(.a(gate463inter10), .b(gate463inter9), .O(gate463inter11));
  nor2  gate3222(.a(gate463inter11), .b(gate463inter6), .O(gate463inter12));
  nand2 gate3223(.a(gate463inter12), .b(gate463inter1), .O(N2331));

  xor2  gate1950(.a(N2139), .b(N2138), .O(gate464inter0));
  nand2 gate1951(.a(gate464inter0), .b(s_40), .O(gate464inter1));
  and2  gate1952(.a(N2139), .b(N2138), .O(gate464inter2));
  inv1  gate1953(.a(s_40), .O(gate464inter3));
  inv1  gate1954(.a(s_41), .O(gate464inter4));
  nand2 gate1955(.a(gate464inter4), .b(gate464inter3), .O(gate464inter5));
  nor2  gate1956(.a(gate464inter5), .b(gate464inter2), .O(gate464inter6));
  inv1  gate1957(.a(N2138), .O(gate464inter7));
  inv1  gate1958(.a(N2139), .O(gate464inter8));
  nand2 gate1959(.a(gate464inter8), .b(gate464inter7), .O(gate464inter9));
  nand2 gate1960(.a(s_41), .b(gate464inter3), .O(gate464inter10));
  nor2  gate1961(.a(gate464inter10), .b(gate464inter9), .O(gate464inter11));
  nor2  gate1962(.a(gate464inter11), .b(gate464inter6), .O(gate464inter12));
  nand2 gate1963(.a(gate464inter12), .b(gate464inter1), .O(N2334));

  xor2  gate3462(.a(N2141), .b(N1936), .O(gate465inter0));
  nand2 gate3463(.a(gate465inter0), .b(s_256), .O(gate465inter1));
  and2  gate3464(.a(N2141), .b(N1936), .O(gate465inter2));
  inv1  gate3465(.a(s_256), .O(gate465inter3));
  inv1  gate3466(.a(s_257), .O(gate465inter4));
  nand2 gate3467(.a(gate465inter4), .b(gate465inter3), .O(gate465inter5));
  nor2  gate3468(.a(gate465inter5), .b(gate465inter2), .O(gate465inter6));
  inv1  gate3469(.a(N1936), .O(gate465inter7));
  inv1  gate3470(.a(N2141), .O(gate465inter8));
  nand2 gate3471(.a(gate465inter8), .b(gate465inter7), .O(gate465inter9));
  nand2 gate3472(.a(s_257), .b(gate465inter3), .O(gate465inter10));
  nor2  gate3473(.a(gate465inter10), .b(gate465inter9), .O(gate465inter11));
  nor2  gate3474(.a(gate465inter11), .b(gate465inter6), .O(gate465inter12));
  nand2 gate3475(.a(gate465inter12), .b(gate465inter1), .O(N2341));
nand2 gate466( .a(N1933), .b(N2142), .O(N2342) );
and2 gate467( .a(N724), .b(N2144), .O(N2347) );
and3 gate468( .a(N2146), .b(N699), .c(N1726), .O(N2348) );
and2 gate469( .a(N753), .b(N2147), .O(N2349) );
and2 gate470( .a(N2148), .b(N1273), .O(N2350) );
and2 gate471( .a(N736), .b(N2150), .O(N2351) );
and2 gate472( .a(N1735), .b(N2153), .O(N2352) );
and2 gate473( .a(N763), .b(N2154), .O(N2353) );
and2 gate474( .a(N1725), .b(N2156), .O(N2354) );
and2 gate475( .a(N749), .b(N2157), .O(N2355) );
inv1 gate476( .a(N2178), .O(N2374) );
inv1 gate477( .a(N2179), .O(N2375) );
and2 gate478( .a(N1520), .b(N2180), .O(N2376) );
and2 gate479( .a(N1721), .b(N2181), .O(N2379) );
and2 gate480( .a(N665), .b(N2211), .O(N2398) );
and3 gate481( .a(N2057), .b(N226), .c(N1873), .O(N2417) );
and3 gate482( .a(N2057), .b(N274), .c(N1306), .O(N2418) );
and2 gate483( .a(N2052), .b(N2238), .O(N2419) );
and3 gate484( .a(N2057), .b(N232), .c(N1878), .O(N2420) );
and3 gate485( .a(N2057), .b(N274), .c(N1306), .O(N2421) );
and2 gate486( .a(N2052), .b(N2239), .O(N2422) );
and3 gate487( .a(N2057), .b(N238), .c(N1883), .O(N2425) );
and3 gate488( .a(N2057), .b(N274), .c(N1306), .O(N2426) );
and2 gate489( .a(N2052), .b(N2240), .O(N2427) );
and3 gate490( .a(N2057), .b(N244), .c(N1888), .O(N2430) );
and3 gate491( .a(N2057), .b(N274), .c(N1306), .O(N2431) );
and2 gate492( .a(N2052), .b(N2241), .O(N2432) );
and3 gate493( .a(N2043), .b(N250), .c(N1893), .O(N2435) );
and3 gate494( .a(N2043), .b(N274), .c(N1322), .O(N2436) );
and2 gate495( .a(N2038), .b(N2242), .O(N2437) );
and3 gate496( .a(N2043), .b(N257), .c(N1898), .O(N2438) );
and3 gate497( .a(N2043), .b(N274), .c(N1315), .O(N2439) );
and2 gate498( .a(N2038), .b(N2243), .O(N2440) );
and3 gate499( .a(N2043), .b(N264), .c(N1903), .O(N2443) );
and3 gate500( .a(N2043), .b(N274), .c(N1315), .O(N2444) );
and2 gate501( .a(N2038), .b(N2244), .O(N2445) );
and3 gate502( .a(N2043), .b(N270), .c(N1908), .O(N2448) );
and3 gate503( .a(N2043), .b(N274), .c(N1315), .O(N2449) );
and2 gate504( .a(N2038), .b(N2245), .O(N2450) );
inv1 gate505( .a(N2313), .O(N2467) );
inv1 gate506( .a(N2316), .O(N2468) );
inv1 gate507( .a(N2319), .O(N2469) );
inv1 gate508( .a(N2322), .O(N2470) );

  xor2  gate1908(.a(N2342), .b(N2341), .O(gate509inter0));
  nand2 gate1909(.a(gate509inter0), .b(s_34), .O(gate509inter1));
  and2  gate1910(.a(N2342), .b(N2341), .O(gate509inter2));
  inv1  gate1911(.a(s_34), .O(gate509inter3));
  inv1  gate1912(.a(s_35), .O(gate509inter4));
  nand2 gate1913(.a(gate509inter4), .b(gate509inter3), .O(gate509inter5));
  nor2  gate1914(.a(gate509inter5), .b(gate509inter2), .O(gate509inter6));
  inv1  gate1915(.a(N2341), .O(gate509inter7));
  inv1  gate1916(.a(N2342), .O(gate509inter8));
  nand2 gate1917(.a(gate509inter8), .b(gate509inter7), .O(gate509inter9));
  nand2 gate1918(.a(s_35), .b(gate509inter3), .O(gate509inter10));
  nor2  gate1919(.a(gate509inter10), .b(gate509inter9), .O(gate509inter11));
  nor2  gate1920(.a(gate509inter11), .b(gate509inter6), .O(gate509inter12));
  nand2 gate1921(.a(gate509inter12), .b(gate509inter1), .O(N2471));
inv1 gate510( .a(N2325), .O(N2474) );
inv1 gate511( .a(N2328), .O(N2475) );
inv1 gate512( .a(N2331), .O(N2476) );
inv1 gate513( .a(N2334), .O(N2477) );
or2 gate514( .a(N2348), .b(N1729), .O(N2478) );
inv1 gate515( .a(N2175), .O(N2481) );
and2 gate516( .a(N2175), .b(N1334), .O(N2482) );
and2 gate517( .a(N2349), .b(N2183), .O(N2483) );
and2 gate518( .a(N2374), .b(N1346), .O(N2486) );
and2 gate519( .a(N2375), .b(N1350), .O(N2487) );
buf1 gate520( .a(N2185), .O(N2488) );
buf1 gate521( .a(N2188), .O(N2497) );
buf1 gate522( .a(N2191), .O(N2506) );
buf1 gate523( .a(N2194), .O(N2515) );
buf1 gate524( .a(N2197), .O(N2524) );
buf1 gate525( .a(N2200), .O(N2533) );
buf1 gate526( .a(N2203), .O(N2542) );
buf1 gate527( .a(N2206), .O(N2551) );
buf1 gate528( .a(N2185), .O(N2560) );
buf1 gate529( .a(N2188), .O(N2569) );
buf1 gate530( .a(N2191), .O(N2578) );
buf1 gate531( .a(N2194), .O(N2587) );
buf1 gate532( .a(N2197), .O(N2596) );
buf1 gate533( .a(N2200), .O(N2605) );
buf1 gate534( .a(N2203), .O(N2614) );
buf1 gate535( .a(N2206), .O(N2623) );
inv1 gate536( .a(N2212), .O(N2632) );
and2 gate537( .a(N2212), .b(N1833), .O(N2633) );
inv1 gate538( .a(N2212), .O(N2634) );
and2 gate539( .a(N2212), .b(N1833), .O(N2635) );
inv1 gate540( .a(N2212), .O(N2636) );
and2 gate541( .a(N2212), .b(N1833), .O(N2637) );
inv1 gate542( .a(N2212), .O(N2638) );
and2 gate543( .a(N2212), .b(N1833), .O(N2639) );
inv1 gate544( .a(N2221), .O(N2640) );
and2 gate545( .a(N2221), .b(N1824), .O(N2641) );
inv1 gate546( .a(N2221), .O(N2642) );
and2 gate547( .a(N2221), .b(N1824), .O(N2643) );
inv1 gate548( .a(N2221), .O(N2644) );
and2 gate549( .a(N2221), .b(N1824), .O(N2645) );
inv1 gate550( .a(N2221), .O(N2646) );
and2 gate551( .a(N2221), .b(N1824), .O(N2647) );
or3 gate552( .a(N2270), .b(N1870), .c(N2068), .O(N2648) );
nor3 gate553( .a(N2270), .b(N1870), .c(N2068), .O(N2652) );
or3 gate554( .a(N2417), .b(N2418), .c(N2419), .O(N2656) );
or3 gate555( .a(N2420), .b(N2421), .c(N2422), .O(N2659) );
or3 gate556( .a(N2277), .b(N1880), .c(N2078), .O(N2662) );
nor3 gate557( .a(N2277), .b(N1880), .c(N2078), .O(N2666) );
or3 gate558( .a(N2425), .b(N2426), .c(N2427), .O(N2670) );
or3 gate559( .a(N2282), .b(N1885), .c(N2083), .O(N2673) );
nor3 gate560( .a(N2282), .b(N1885), .c(N2083), .O(N2677) );
or3 gate561( .a(N2430), .b(N2431), .c(N2432), .O(N2681) );
or3 gate562( .a(N2287), .b(N1890), .c(N2088), .O(N2684) );
nor3 gate563( .a(N2287), .b(N1890), .c(N2088), .O(N2688) );
or3 gate564( .a(N2435), .b(N2436), .c(N2437), .O(N2692) );
or3 gate565( .a(N2438), .b(N2439), .c(N2440), .O(N2697) );
or3 gate566( .a(N2294), .b(N1900), .c(N2098), .O(N2702) );
nor3 gate567( .a(N2294), .b(N1900), .c(N2098), .O(N2706) );
or3 gate568( .a(N2443), .b(N2444), .c(N2445), .O(N2710) );
or3 gate569( .a(N2299), .b(N1905), .c(N2103), .O(N2715) );
nor3 gate570( .a(N2299), .b(N1905), .c(N2103), .O(N2719) );
or3 gate571( .a(N2448), .b(N2449), .c(N2450), .O(N2723) );
inv1 gate572( .a(N2304), .O(N2728) );
inv1 gate573( .a(N2158), .O(N2729) );
and2 gate574( .a(N1562), .b(N2158), .O(N2730) );
inv1 gate575( .a(N2158), .O(N2731) );
and2 gate576( .a(N1562), .b(N2158), .O(N2732) );
inv1 gate577( .a(N2158), .O(N2733) );
and2 gate578( .a(N1562), .b(N2158), .O(N2734) );
inv1 gate579( .a(N2158), .O(N2735) );
and2 gate580( .a(N1562), .b(N2158), .O(N2736) );
inv1 gate581( .a(N2158), .O(N2737) );
and2 gate582( .a(N1562), .b(N2158), .O(N2738) );
inv1 gate583( .a(N2158), .O(N2739) );
and2 gate584( .a(N1562), .b(N2158), .O(N2740) );
inv1 gate585( .a(N2158), .O(N2741) );
and2 gate586( .a(N1562), .b(N2158), .O(N2742) );
inv1 gate587( .a(N2158), .O(N2743) );
and2 gate588( .a(N1562), .b(N2158), .O(N2744) );
or3 gate589( .a(N2376), .b(N1983), .c(N2379), .O(N2745) );
nor3 gate590( .a(N2376), .b(N1983), .c(N2379), .O(N2746) );

  xor2  gate1922(.a(N2467), .b(N2316), .O(gate591inter0));
  nand2 gate1923(.a(gate591inter0), .b(s_36), .O(gate591inter1));
  and2  gate1924(.a(N2467), .b(N2316), .O(gate591inter2));
  inv1  gate1925(.a(s_36), .O(gate591inter3));
  inv1  gate1926(.a(s_37), .O(gate591inter4));
  nand2 gate1927(.a(gate591inter4), .b(gate591inter3), .O(gate591inter5));
  nor2  gate1928(.a(gate591inter5), .b(gate591inter2), .O(gate591inter6));
  inv1  gate1929(.a(N2316), .O(gate591inter7));
  inv1  gate1930(.a(N2467), .O(gate591inter8));
  nand2 gate1931(.a(gate591inter8), .b(gate591inter7), .O(gate591inter9));
  nand2 gate1932(.a(s_37), .b(gate591inter3), .O(gate591inter10));
  nor2  gate1933(.a(gate591inter10), .b(gate591inter9), .O(gate591inter11));
  nor2  gate1934(.a(gate591inter11), .b(gate591inter6), .O(gate591inter12));
  nand2 gate1935(.a(gate591inter12), .b(gate591inter1), .O(N2748));

  xor2  gate4372(.a(N2468), .b(N2313), .O(gate592inter0));
  nand2 gate4373(.a(gate592inter0), .b(s_386), .O(gate592inter1));
  and2  gate4374(.a(N2468), .b(N2313), .O(gate592inter2));
  inv1  gate4375(.a(s_386), .O(gate592inter3));
  inv1  gate4376(.a(s_387), .O(gate592inter4));
  nand2 gate4377(.a(gate592inter4), .b(gate592inter3), .O(gate592inter5));
  nor2  gate4378(.a(gate592inter5), .b(gate592inter2), .O(gate592inter6));
  inv1  gate4379(.a(N2313), .O(gate592inter7));
  inv1  gate4380(.a(N2468), .O(gate592inter8));
  nand2 gate4381(.a(gate592inter8), .b(gate592inter7), .O(gate592inter9));
  nand2 gate4382(.a(s_387), .b(gate592inter3), .O(gate592inter10));
  nor2  gate4383(.a(gate592inter10), .b(gate592inter9), .O(gate592inter11));
  nor2  gate4384(.a(gate592inter11), .b(gate592inter6), .O(gate592inter12));
  nand2 gate4385(.a(gate592inter12), .b(gate592inter1), .O(N2749));

  xor2  gate2692(.a(N2469), .b(N2322), .O(gate593inter0));
  nand2 gate2693(.a(gate593inter0), .b(s_146), .O(gate593inter1));
  and2  gate2694(.a(N2469), .b(N2322), .O(gate593inter2));
  inv1  gate2695(.a(s_146), .O(gate593inter3));
  inv1  gate2696(.a(s_147), .O(gate593inter4));
  nand2 gate2697(.a(gate593inter4), .b(gate593inter3), .O(gate593inter5));
  nor2  gate2698(.a(gate593inter5), .b(gate593inter2), .O(gate593inter6));
  inv1  gate2699(.a(N2322), .O(gate593inter7));
  inv1  gate2700(.a(N2469), .O(gate593inter8));
  nand2 gate2701(.a(gate593inter8), .b(gate593inter7), .O(gate593inter9));
  nand2 gate2702(.a(s_147), .b(gate593inter3), .O(gate593inter10));
  nor2  gate2703(.a(gate593inter10), .b(gate593inter9), .O(gate593inter11));
  nor2  gate2704(.a(gate593inter11), .b(gate593inter6), .O(gate593inter12));
  nand2 gate2705(.a(gate593inter12), .b(gate593inter1), .O(N2750));

  xor2  gate2174(.a(N2470), .b(N2319), .O(gate594inter0));
  nand2 gate2175(.a(gate594inter0), .b(s_72), .O(gate594inter1));
  and2  gate2176(.a(N2470), .b(N2319), .O(gate594inter2));
  inv1  gate2177(.a(s_72), .O(gate594inter3));
  inv1  gate2178(.a(s_73), .O(gate594inter4));
  nand2 gate2179(.a(gate594inter4), .b(gate594inter3), .O(gate594inter5));
  nor2  gate2180(.a(gate594inter5), .b(gate594inter2), .O(gate594inter6));
  inv1  gate2181(.a(N2319), .O(gate594inter7));
  inv1  gate2182(.a(N2470), .O(gate594inter8));
  nand2 gate2183(.a(gate594inter8), .b(gate594inter7), .O(gate594inter9));
  nand2 gate2184(.a(s_73), .b(gate594inter3), .O(gate594inter10));
  nor2  gate2185(.a(gate594inter10), .b(gate594inter9), .O(gate594inter11));
  nor2  gate2186(.a(gate594inter11), .b(gate594inter6), .O(gate594inter12));
  nand2 gate2187(.a(gate594inter12), .b(gate594inter1), .O(N2751));

  xor2  gate1726(.a(N2474), .b(N2328), .O(gate595inter0));
  nand2 gate1727(.a(gate595inter0), .b(s_8), .O(gate595inter1));
  and2  gate1728(.a(N2474), .b(N2328), .O(gate595inter2));
  inv1  gate1729(.a(s_8), .O(gate595inter3));
  inv1  gate1730(.a(s_9), .O(gate595inter4));
  nand2 gate1731(.a(gate595inter4), .b(gate595inter3), .O(gate595inter5));
  nor2  gate1732(.a(gate595inter5), .b(gate595inter2), .O(gate595inter6));
  inv1  gate1733(.a(N2328), .O(gate595inter7));
  inv1  gate1734(.a(N2474), .O(gate595inter8));
  nand2 gate1735(.a(gate595inter8), .b(gate595inter7), .O(gate595inter9));
  nand2 gate1736(.a(s_9), .b(gate595inter3), .O(gate595inter10));
  nor2  gate1737(.a(gate595inter10), .b(gate595inter9), .O(gate595inter11));
  nor2  gate1738(.a(gate595inter11), .b(gate595inter6), .O(gate595inter12));
  nand2 gate1739(.a(gate595inter12), .b(gate595inter1), .O(N2754));
nand2 gate596( .a(N2325), .b(N2475), .O(N2755) );
nand2 gate597( .a(N2334), .b(N2476), .O(N2756) );

  xor2  gate2440(.a(N2477), .b(N2331), .O(gate598inter0));
  nand2 gate2441(.a(gate598inter0), .b(s_110), .O(gate598inter1));
  and2  gate2442(.a(N2477), .b(N2331), .O(gate598inter2));
  inv1  gate2443(.a(s_110), .O(gate598inter3));
  inv1  gate2444(.a(s_111), .O(gate598inter4));
  nand2 gate2445(.a(gate598inter4), .b(gate598inter3), .O(gate598inter5));
  nor2  gate2446(.a(gate598inter5), .b(gate598inter2), .O(gate598inter6));
  inv1  gate2447(.a(N2331), .O(gate598inter7));
  inv1  gate2448(.a(N2477), .O(gate598inter8));
  nand2 gate2449(.a(gate598inter8), .b(gate598inter7), .O(gate598inter9));
  nand2 gate2450(.a(s_111), .b(gate598inter3), .O(gate598inter10));
  nor2  gate2451(.a(gate598inter10), .b(gate598inter9), .O(gate598inter11));
  nor2  gate2452(.a(gate598inter11), .b(gate598inter6), .O(gate598inter12));
  nand2 gate2453(.a(gate598inter12), .b(gate598inter1), .O(N2757));
and2 gate599( .a(N1520), .b(N2481), .O(N2758) );
and2 gate600( .a(N1722), .b(N2482), .O(N2761) );
and2 gate601( .a(N2478), .b(N1770), .O(N2764) );
or3 gate602( .a(N2486), .b(N1789), .c(N1790), .O(N2768) );
or3 gate603( .a(N2487), .b(N1797), .c(N1798), .O(N2769) );
and2 gate604( .a(N665), .b(N2633), .O(N2898) );
and2 gate605( .a(N679), .b(N2635), .O(N2899) );
and2 gate606( .a(N686), .b(N2637), .O(N2900) );
and2 gate607( .a(N702), .b(N2639), .O(N2901) );
inv1 gate608( .a(N2746), .O(N2962) );
nand2 gate609( .a(N2748), .b(N2749), .O(N2966) );

  xor2  gate3896(.a(N2751), .b(N2750), .O(gate610inter0));
  nand2 gate3897(.a(gate610inter0), .b(s_318), .O(gate610inter1));
  and2  gate3898(.a(N2751), .b(N2750), .O(gate610inter2));
  inv1  gate3899(.a(s_318), .O(gate610inter3));
  inv1  gate3900(.a(s_319), .O(gate610inter4));
  nand2 gate3901(.a(gate610inter4), .b(gate610inter3), .O(gate610inter5));
  nor2  gate3902(.a(gate610inter5), .b(gate610inter2), .O(gate610inter6));
  inv1  gate3903(.a(N2750), .O(gate610inter7));
  inv1  gate3904(.a(N2751), .O(gate610inter8));
  nand2 gate3905(.a(gate610inter8), .b(gate610inter7), .O(gate610inter9));
  nand2 gate3906(.a(s_319), .b(gate610inter3), .O(gate610inter10));
  nor2  gate3907(.a(gate610inter10), .b(gate610inter9), .O(gate610inter11));
  nor2  gate3908(.a(gate610inter11), .b(gate610inter6), .O(gate610inter12));
  nand2 gate3909(.a(gate610inter12), .b(gate610inter1), .O(N2967));
buf1 gate611( .a(N2471), .O(N2970) );
nand2 gate612( .a(N2754), .b(N2755), .O(N2973) );
nand2 gate613( .a(N2756), .b(N2757), .O(N2977) );
and2 gate614( .a(N2471), .b(N2143), .O(N2980) );
inv1 gate615( .a(N2488), .O(N2984) );
inv1 gate616( .a(N2497), .O(N2985) );
inv1 gate617( .a(N2506), .O(N2986) );
inv1 gate618( .a(N2515), .O(N2987) );
inv1 gate619( .a(N2524), .O(N2988) );
inv1 gate620( .a(N2533), .O(N2989) );
inv1 gate621( .a(N2542), .O(N2990) );
inv1 gate622( .a(N2551), .O(N2991) );
inv1 gate623( .a(N2488), .O(N2992) );
inv1 gate624( .a(N2497), .O(N2993) );
inv1 gate625( .a(N2506), .O(N2994) );
inv1 gate626( .a(N2515), .O(N2995) );
inv1 gate627( .a(N2524), .O(N2996) );
inv1 gate628( .a(N2533), .O(N2997) );
inv1 gate629( .a(N2542), .O(N2998) );
inv1 gate630( .a(N2551), .O(N2999) );
inv1 gate631( .a(N2488), .O(N3000) );
inv1 gate632( .a(N2497), .O(N3001) );
inv1 gate633( .a(N2506), .O(N3002) );
inv1 gate634( .a(N2515), .O(N3003) );
inv1 gate635( .a(N2524), .O(N3004) );
inv1 gate636( .a(N2533), .O(N3005) );
inv1 gate637( .a(N2542), .O(N3006) );
inv1 gate638( .a(N2551), .O(N3007) );
inv1 gate639( .a(N2488), .O(N3008) );
inv1 gate640( .a(N2497), .O(N3009) );
inv1 gate641( .a(N2506), .O(N3010) );
inv1 gate642( .a(N2515), .O(N3011) );
inv1 gate643( .a(N2524), .O(N3012) );
inv1 gate644( .a(N2533), .O(N3013) );
inv1 gate645( .a(N2542), .O(N3014) );
inv1 gate646( .a(N2551), .O(N3015) );
inv1 gate647( .a(N2488), .O(N3016) );
inv1 gate648( .a(N2497), .O(N3017) );
inv1 gate649( .a(N2506), .O(N3018) );
inv1 gate650( .a(N2515), .O(N3019) );
inv1 gate651( .a(N2524), .O(N3020) );
inv1 gate652( .a(N2533), .O(N3021) );
inv1 gate653( .a(N2542), .O(N3022) );
inv1 gate654( .a(N2551), .O(N3023) );
inv1 gate655( .a(N2488), .O(N3024) );
inv1 gate656( .a(N2497), .O(N3025) );
inv1 gate657( .a(N2506), .O(N3026) );
inv1 gate658( .a(N2515), .O(N3027) );
inv1 gate659( .a(N2524), .O(N3028) );
inv1 gate660( .a(N2533), .O(N3029) );
inv1 gate661( .a(N2542), .O(N3030) );
inv1 gate662( .a(N2551), .O(N3031) );
inv1 gate663( .a(N2488), .O(N3032) );
inv1 gate664( .a(N2497), .O(N3033) );
inv1 gate665( .a(N2506), .O(N3034) );
inv1 gate666( .a(N2515), .O(N3035) );
inv1 gate667( .a(N2524), .O(N3036) );
inv1 gate668( .a(N2533), .O(N3037) );
inv1 gate669( .a(N2542), .O(N3038) );
inv1 gate670( .a(N2551), .O(N3039) );
inv1 gate671( .a(N2488), .O(N3040) );
inv1 gate672( .a(N2497), .O(N3041) );
inv1 gate673( .a(N2506), .O(N3042) );
inv1 gate674( .a(N2515), .O(N3043) );
inv1 gate675( .a(N2524), .O(N3044) );
inv1 gate676( .a(N2533), .O(N3045) );
inv1 gate677( .a(N2542), .O(N3046) );
inv1 gate678( .a(N2551), .O(N3047) );
inv1 gate679( .a(N2560), .O(N3048) );
inv1 gate680( .a(N2569), .O(N3049) );
inv1 gate681( .a(N2578), .O(N3050) );
inv1 gate682( .a(N2587), .O(N3051) );
inv1 gate683( .a(N2596), .O(N3052) );
inv1 gate684( .a(N2605), .O(N3053) );
inv1 gate685( .a(N2614), .O(N3054) );
inv1 gate686( .a(N2623), .O(N3055) );
inv1 gate687( .a(N2560), .O(N3056) );
inv1 gate688( .a(N2569), .O(N3057) );
inv1 gate689( .a(N2578), .O(N3058) );
inv1 gate690( .a(N2587), .O(N3059) );
inv1 gate691( .a(N2596), .O(N3060) );
inv1 gate692( .a(N2605), .O(N3061) );
inv1 gate693( .a(N2614), .O(N3062) );
inv1 gate694( .a(N2623), .O(N3063) );
inv1 gate695( .a(N2560), .O(N3064) );
inv1 gate696( .a(N2569), .O(N3065) );
inv1 gate697( .a(N2578), .O(N3066) );
inv1 gate698( .a(N2587), .O(N3067) );
inv1 gate699( .a(N2596), .O(N3068) );
inv1 gate700( .a(N2605), .O(N3069) );
inv1 gate701( .a(N2614), .O(N3070) );
inv1 gate702( .a(N2623), .O(N3071) );
inv1 gate703( .a(N2560), .O(N3072) );
inv1 gate704( .a(N2569), .O(N3073) );
inv1 gate705( .a(N2578), .O(N3074) );
inv1 gate706( .a(N2587), .O(N3075) );
inv1 gate707( .a(N2596), .O(N3076) );
inv1 gate708( .a(N2605), .O(N3077) );
inv1 gate709( .a(N2614), .O(N3078) );
inv1 gate710( .a(N2623), .O(N3079) );
inv1 gate711( .a(N2560), .O(N3080) );
inv1 gate712( .a(N2569), .O(N3081) );
inv1 gate713( .a(N2578), .O(N3082) );
inv1 gate714( .a(N2587), .O(N3083) );
inv1 gate715( .a(N2596), .O(N3084) );
inv1 gate716( .a(N2605), .O(N3085) );
inv1 gate717( .a(N2614), .O(N3086) );
inv1 gate718( .a(N2623), .O(N3087) );
inv1 gate719( .a(N2560), .O(N3088) );
inv1 gate720( .a(N2569), .O(N3089) );
inv1 gate721( .a(N2578), .O(N3090) );
inv1 gate722( .a(N2587), .O(N3091) );
inv1 gate723( .a(N2596), .O(N3092) );
inv1 gate724( .a(N2605), .O(N3093) );
inv1 gate725( .a(N2614), .O(N3094) );
inv1 gate726( .a(N2623), .O(N3095) );
inv1 gate727( .a(N2560), .O(N3096) );
inv1 gate728( .a(N2569), .O(N3097) );
inv1 gate729( .a(N2578), .O(N3098) );
inv1 gate730( .a(N2587), .O(N3099) );
inv1 gate731( .a(N2596), .O(N3100) );
inv1 gate732( .a(N2605), .O(N3101) );
inv1 gate733( .a(N2614), .O(N3102) );
inv1 gate734( .a(N2623), .O(N3103) );
inv1 gate735( .a(N2560), .O(N3104) );
inv1 gate736( .a(N2569), .O(N3105) );
inv1 gate737( .a(N2578), .O(N3106) );
inv1 gate738( .a(N2587), .O(N3107) );
inv1 gate739( .a(N2596), .O(N3108) );
inv1 gate740( .a(N2605), .O(N3109) );
inv1 gate741( .a(N2614), .O(N3110) );
inv1 gate742( .a(N2623), .O(N3111) );
buf1 gate743( .a(N2656), .O(N3112) );
inv1 gate744( .a(N2656), .O(N3115) );
inv1 gate745( .a(N2652), .O(N3118) );
and2 gate746( .a(N2768), .b(N1674), .O(N3119) );
buf1 gate747( .a(N2659), .O(N3122) );
inv1 gate748( .a(N2659), .O(N3125) );
buf1 gate749( .a(N2670), .O(N3128) );
inv1 gate750( .a(N2670), .O(N3131) );
inv1 gate751( .a(N2666), .O(N3134) );
buf1 gate752( .a(N2681), .O(N3135) );
inv1 gate753( .a(N2681), .O(N3138) );
inv1 gate754( .a(N2677), .O(N3141) );
buf1 gate755( .a(N2692), .O(N3142) );
inv1 gate756( .a(N2692), .O(N3145) );
inv1 gate757( .a(N2688), .O(N3148) );
and2 gate758( .a(N2769), .b(N1678), .O(N3149) );
buf1 gate759( .a(N2697), .O(N3152) );
inv1 gate760( .a(N2697), .O(N3155) );
buf1 gate761( .a(N2710), .O(N3158) );
inv1 gate762( .a(N2710), .O(N3161) );
inv1 gate763( .a(N2706), .O(N3164) );
buf1 gate764( .a(N2723), .O(N3165) );
inv1 gate765( .a(N2723), .O(N3168) );
inv1 gate766( .a(N2719), .O(N3171) );
and2 gate767( .a(N1909), .b(N2648), .O(N3172) );
and2 gate768( .a(N1913), .b(N2662), .O(N3175) );
and2 gate769( .a(N1913), .b(N2673), .O(N3178) );
and2 gate770( .a(N1913), .b(N2684), .O(N3181) );
and2 gate771( .a(N1922), .b(N2702), .O(N3184) );
and2 gate772( .a(N1922), .b(N2715), .O(N3187) );
inv1 gate773( .a(N2692), .O(N3190) );
inv1 gate774( .a(N2697), .O(N3191) );
inv1 gate775( .a(N2710), .O(N3192) );
inv1 gate776( .a(N2723), .O(N3193) );
and5 gate777( .a(N2692), .b(N2697), .c(N2710), .d(N2723), .e(N1459), .O(N3194) );

  xor2  gate2076(.a(N2962), .b(N2745), .O(gate778inter0));
  nand2 gate2077(.a(gate778inter0), .b(s_58), .O(gate778inter1));
  and2  gate2078(.a(N2962), .b(N2745), .O(gate778inter2));
  inv1  gate2079(.a(s_58), .O(gate778inter3));
  inv1  gate2080(.a(s_59), .O(gate778inter4));
  nand2 gate2081(.a(gate778inter4), .b(gate778inter3), .O(gate778inter5));
  nor2  gate2082(.a(gate778inter5), .b(gate778inter2), .O(gate778inter6));
  inv1  gate2083(.a(N2745), .O(gate778inter7));
  inv1  gate2084(.a(N2962), .O(gate778inter8));
  nand2 gate2085(.a(gate778inter8), .b(gate778inter7), .O(gate778inter9));
  nand2 gate2086(.a(s_59), .b(gate778inter3), .O(gate778inter10));
  nor2  gate2087(.a(gate778inter10), .b(gate778inter9), .O(gate778inter11));
  nor2  gate2088(.a(gate778inter11), .b(gate778inter6), .O(gate778inter12));
  nand2 gate2089(.a(gate778inter12), .b(gate778inter1), .O(N3195));
inv1 gate779( .a(N2966), .O(N3196) );
or3 gate780( .a(N2980), .b(N2145), .c(N2347), .O(N3206) );
and2 gate781( .a(N124), .b(N2984), .O(N3207) );
and2 gate782( .a(N159), .b(N2985), .O(N3208) );
and2 gate783( .a(N150), .b(N2986), .O(N3209) );
and2 gate784( .a(N143), .b(N2987), .O(N3210) );
and2 gate785( .a(N137), .b(N2988), .O(N3211) );
and2 gate786( .a(N132), .b(N2989), .O(N3212) );
and2 gate787( .a(N128), .b(N2990), .O(N3213) );
and2 gate788( .a(N125), .b(N2991), .O(N3214) );
and2 gate789( .a(N125), .b(N2992), .O(N3215) );
and2 gate790( .a(N655), .b(N2993), .O(N3216) );
and2 gate791( .a(N159), .b(N2994), .O(N3217) );
and2 gate792( .a(N150), .b(N2995), .O(N3218) );
and2 gate793( .a(N143), .b(N2996), .O(N3219) );
and2 gate794( .a(N137), .b(N2997), .O(N3220) );
and2 gate795( .a(N132), .b(N2998), .O(N3221) );
and2 gate796( .a(N128), .b(N2999), .O(N3222) );
and2 gate797( .a(N128), .b(N3000), .O(N3223) );
and2 gate798( .a(N670), .b(N3001), .O(N3224) );
and2 gate799( .a(N655), .b(N3002), .O(N3225) );
and2 gate800( .a(N159), .b(N3003), .O(N3226) );
and2 gate801( .a(N150), .b(N3004), .O(N3227) );
and2 gate802( .a(N143), .b(N3005), .O(N3228) );
and2 gate803( .a(N137), .b(N3006), .O(N3229) );
and2 gate804( .a(N132), .b(N3007), .O(N3230) );
and2 gate805( .a(N132), .b(N3008), .O(N3231) );
and2 gate806( .a(N690), .b(N3009), .O(N3232) );
and2 gate807( .a(N670), .b(N3010), .O(N3233) );
and2 gate808( .a(N655), .b(N3011), .O(N3234) );
and2 gate809( .a(N159), .b(N3012), .O(N3235) );
and2 gate810( .a(N150), .b(N3013), .O(N3236) );
and2 gate811( .a(N143), .b(N3014), .O(N3237) );
and2 gate812( .a(N137), .b(N3015), .O(N3238) );
and2 gate813( .a(N137), .b(N3016), .O(N3239) );
and2 gate814( .a(N706), .b(N3017), .O(N3240) );
and2 gate815( .a(N690), .b(N3018), .O(N3241) );
and2 gate816( .a(N670), .b(N3019), .O(N3242) );
and2 gate817( .a(N655), .b(N3020), .O(N3243) );
and2 gate818( .a(N159), .b(N3021), .O(N3244) );
and2 gate819( .a(N150), .b(N3022), .O(N3245) );
and2 gate820( .a(N143), .b(N3023), .O(N3246) );
and2 gate821( .a(N143), .b(N3024), .O(N3247) );
and2 gate822( .a(N715), .b(N3025), .O(N3248) );
and2 gate823( .a(N706), .b(N3026), .O(N3249) );
and2 gate824( .a(N690), .b(N3027), .O(N3250) );
and2 gate825( .a(N670), .b(N3028), .O(N3251) );
and2 gate826( .a(N655), .b(N3029), .O(N3252) );
and2 gate827( .a(N159), .b(N3030), .O(N3253) );
and2 gate828( .a(N150), .b(N3031), .O(N3254) );
and2 gate829( .a(N150), .b(N3032), .O(N3255) );
and2 gate830( .a(N727), .b(N3033), .O(N3256) );
and2 gate831( .a(N715), .b(N3034), .O(N3257) );
and2 gate832( .a(N706), .b(N3035), .O(N3258) );
and2 gate833( .a(N690), .b(N3036), .O(N3259) );
and2 gate834( .a(N670), .b(N3037), .O(N3260) );
and2 gate835( .a(N655), .b(N3038), .O(N3261) );
and2 gate836( .a(N159), .b(N3039), .O(N3262) );
and2 gate837( .a(N159), .b(N3040), .O(N3263) );
and2 gate838( .a(N740), .b(N3041), .O(N3264) );
and2 gate839( .a(N727), .b(N3042), .O(N3265) );
and2 gate840( .a(N715), .b(N3043), .O(N3266) );
and2 gate841( .a(N706), .b(N3044), .O(N3267) );
and2 gate842( .a(N690), .b(N3045), .O(N3268) );
and2 gate843( .a(N670), .b(N3046), .O(N3269) );
and2 gate844( .a(N655), .b(N3047), .O(N3270) );
and2 gate845( .a(N283), .b(N3048), .O(N3271) );
and2 gate846( .a(N670), .b(N3049), .O(N3272) );
and2 gate847( .a(N690), .b(N3050), .O(N3273) );
and2 gate848( .a(N706), .b(N3051), .O(N3274) );
and2 gate849( .a(N715), .b(N3052), .O(N3275) );
and2 gate850( .a(N727), .b(N3053), .O(N3276) );
and2 gate851( .a(N740), .b(N3054), .O(N3277) );
and2 gate852( .a(N753), .b(N3055), .O(N3278) );
and2 gate853( .a(N294), .b(N3056), .O(N3279) );
and2 gate854( .a(N690), .b(N3057), .O(N3280) );
and2 gate855( .a(N706), .b(N3058), .O(N3281) );
and2 gate856( .a(N715), .b(N3059), .O(N3282) );
and2 gate857( .a(N727), .b(N3060), .O(N3283) );
and2 gate858( .a(N740), .b(N3061), .O(N3284) );
and2 gate859( .a(N753), .b(N3062), .O(N3285) );
and2 gate860( .a(N283), .b(N3063), .O(N3286) );
and2 gate861( .a(N303), .b(N3064), .O(N3287) );
and2 gate862( .a(N706), .b(N3065), .O(N3288) );
and2 gate863( .a(N715), .b(N3066), .O(N3289) );
and2 gate864( .a(N727), .b(N3067), .O(N3290) );
and2 gate865( .a(N740), .b(N3068), .O(N3291) );
and2 gate866( .a(N753), .b(N3069), .O(N3292) );
and2 gate867( .a(N283), .b(N3070), .O(N3293) );
and2 gate868( .a(N294), .b(N3071), .O(N3294) );
and2 gate869( .a(N311), .b(N3072), .O(N3295) );
and2 gate870( .a(N715), .b(N3073), .O(N3296) );
and2 gate871( .a(N727), .b(N3074), .O(N3297) );
and2 gate872( .a(N740), .b(N3075), .O(N3298) );
and2 gate873( .a(N753), .b(N3076), .O(N3299) );
and2 gate874( .a(N283), .b(N3077), .O(N3300) );
and2 gate875( .a(N294), .b(N3078), .O(N3301) );
and2 gate876( .a(N303), .b(N3079), .O(N3302) );
and2 gate877( .a(N317), .b(N3080), .O(N3303) );
and2 gate878( .a(N727), .b(N3081), .O(N3304) );
and2 gate879( .a(N740), .b(N3082), .O(N3305) );
and2 gate880( .a(N753), .b(N3083), .O(N3306) );
and2 gate881( .a(N283), .b(N3084), .O(N3307) );
and2 gate882( .a(N294), .b(N3085), .O(N3308) );
and2 gate883( .a(N303), .b(N3086), .O(N3309) );
and2 gate884( .a(N311), .b(N3087), .O(N3310) );
and2 gate885( .a(N322), .b(N3088), .O(N3311) );
and2 gate886( .a(N740), .b(N3089), .O(N3312) );
and2 gate887( .a(N753), .b(N3090), .O(N3313) );
and2 gate888( .a(N283), .b(N3091), .O(N3314) );
and2 gate889( .a(N294), .b(N3092), .O(N3315) );
and2 gate890( .a(N303), .b(N3093), .O(N3316) );
and2 gate891( .a(N311), .b(N3094), .O(N3317) );
and2 gate892( .a(N317), .b(N3095), .O(N3318) );
and2 gate893( .a(N326), .b(N3096), .O(N3319) );
and2 gate894( .a(N753), .b(N3097), .O(N3320) );
and2 gate895( .a(N283), .b(N3098), .O(N3321) );
and2 gate896( .a(N294), .b(N3099), .O(N3322) );
and2 gate897( .a(N303), .b(N3100), .O(N3323) );
and2 gate898( .a(N311), .b(N3101), .O(N3324) );
and2 gate899( .a(N317), .b(N3102), .O(N3325) );
and2 gate900( .a(N322), .b(N3103), .O(N3326) );
and2 gate901( .a(N329), .b(N3104), .O(N3327) );
and2 gate902( .a(N283), .b(N3105), .O(N3328) );
and2 gate903( .a(N294), .b(N3106), .O(N3329) );
and2 gate904( .a(N303), .b(N3107), .O(N3330) );
and2 gate905( .a(N311), .b(N3108), .O(N3331) );
and2 gate906( .a(N317), .b(N3109), .O(N3332) );
and2 gate907( .a(N322), .b(N3110), .O(N3333) );
and2 gate908( .a(N326), .b(N3111), .O(N3334) );
and5 gate909( .a(N3190), .b(N3191), .c(N3192), .d(N3193), .e(N917), .O(N3383) );
buf1 gate910( .a(N2977), .O(N3384) );
and2 gate911( .a(N3196), .b(N1736), .O(N3387) );
and2 gate912( .a(N2977), .b(N2149), .O(N3388) );
and2 gate913( .a(N2973), .b(N1737), .O(N3389) );
nor8 gate914( .a(N3207), .b(N3208), .c(N3209), .d(N3210), .e(N3211), .f(N3212), .g(N3213), .h(N3214), .O(N3390) );
nor8 gate915( .a(N3215), .b(N3216), .c(N3217), .d(N3218), .e(N3219), .f(N3220), .g(N3221), .h(N3222), .O(N3391) );
nor8 gate916( .a(N3223), .b(N3224), .c(N3225), .d(N3226), .e(N3227), .f(N3228), .g(N3229), .h(N3230), .O(N3392) );
nor8 gate917( .a(N3231), .b(N3232), .c(N3233), .d(N3234), .e(N3235), .f(N3236), .g(N3237), .h(N3238), .O(N3393) );
nor8 gate918( .a(N3239), .b(N3240), .c(N3241), .d(N3242), .e(N3243), .f(N3244), .g(N3245), .h(N3246), .O(N3394) );
nor8 gate919( .a(N3247), .b(N3248), .c(N3249), .d(N3250), .e(N3251), .f(N3252), .g(N3253), .h(N3254), .O(N3395) );
nor8 gate920( .a(N3255), .b(N3256), .c(N3257), .d(N3258), .e(N3259), .f(N3260), .g(N3261), .h(N3262), .O(N3396) );
nor8 gate921( .a(N3263), .b(N3264), .c(N3265), .d(N3266), .e(N3267), .f(N3268), .g(N3269), .h(N3270), .O(N3397) );
nor8 gate922( .a(N3271), .b(N3272), .c(N3273), .d(N3274), .e(N3275), .f(N3276), .g(N3277), .h(N3278), .O(N3398) );
nor8 gate923( .a(N3279), .b(N3280), .c(N3281), .d(N3282), .e(N3283), .f(N3284), .g(N3285), .h(N3286), .O(N3399) );
nor8 gate924( .a(N3287), .b(N3288), .c(N3289), .d(N3290), .e(N3291), .f(N3292), .g(N3293), .h(N3294), .O(N3400) );
nor8 gate925( .a(N3295), .b(N3296), .c(N3297), .d(N3298), .e(N3299), .f(N3300), .g(N3301), .h(N3302), .O(N3401) );
nor8 gate926( .a(N3303), .b(N3304), .c(N3305), .d(N3306), .e(N3307), .f(N3308), .g(N3309), .h(N3310), .O(N3402) );
nor8 gate927( .a(N3311), .b(N3312), .c(N3313), .d(N3314), .e(N3315), .f(N3316), .g(N3317), .h(N3318), .O(N3403) );
nor8 gate928( .a(N3319), .b(N3320), .c(N3321), .d(N3322), .e(N3323), .f(N3324), .g(N3325), .h(N3326), .O(N3404) );
nor8 gate929( .a(N3327), .b(N3328), .c(N3329), .d(N3330), .e(N3331), .f(N3332), .g(N3333), .h(N3334), .O(N3405) );
and2 gate930( .a(N3206), .b(N2641), .O(N3406) );
and3 gate931( .a(N169), .b(N2648), .c(N3112), .O(N3407) );
and3 gate932( .a(N179), .b(N2648), .c(N3115), .O(N3410) );
and3 gate933( .a(N190), .b(N2652), .c(N3115), .O(N3413) );
and3 gate934( .a(N200), .b(N2652), .c(N3112), .O(N3414) );
or3 gate935( .a(N3119), .b(N1875), .c(N2073), .O(N3415) );
nor3 gate936( .a(N3119), .b(N1875), .c(N2073), .O(N3419) );
and3 gate937( .a(N169), .b(N2662), .c(N3128), .O(N3423) );
and3 gate938( .a(N179), .b(N2662), .c(N3131), .O(N3426) );
and3 gate939( .a(N190), .b(N2666), .c(N3131), .O(N3429) );
and3 gate940( .a(N200), .b(N2666), .c(N3128), .O(N3430) );
and3 gate941( .a(N169), .b(N2673), .c(N3135), .O(N3431) );
and3 gate942( .a(N179), .b(N2673), .c(N3138), .O(N3434) );
and3 gate943( .a(N190), .b(N2677), .c(N3138), .O(N3437) );
and3 gate944( .a(N200), .b(N2677), .c(N3135), .O(N3438) );
and3 gate945( .a(N169), .b(N2684), .c(N3142), .O(N3439) );
and3 gate946( .a(N179), .b(N2684), .c(N3145), .O(N3442) );
and3 gate947( .a(N190), .b(N2688), .c(N3145), .O(N3445) );
and3 gate948( .a(N200), .b(N2688), .c(N3142), .O(N3446) );
or3 gate949( .a(N3149), .b(N1895), .c(N2093), .O(N3447) );
nor3 gate950( .a(N3149), .b(N1895), .c(N2093), .O(N3451) );
and3 gate951( .a(N169), .b(N2702), .c(N3158), .O(N3455) );
and3 gate952( .a(N179), .b(N2702), .c(N3161), .O(N3458) );
and3 gate953( .a(N190), .b(N2706), .c(N3161), .O(N3461) );
and3 gate954( .a(N200), .b(N2706), .c(N3158), .O(N3462) );
and3 gate955( .a(N169), .b(N2715), .c(N3165), .O(N3463) );
and3 gate956( .a(N179), .b(N2715), .c(N3168), .O(N3466) );
and3 gate957( .a(N190), .b(N2719), .c(N3168), .O(N3469) );
and3 gate958( .a(N200), .b(N2719), .c(N3165), .O(N3470) );
or2 gate959( .a(N3194), .b(N3383), .O(N3471) );
buf1 gate960( .a(N2967), .O(N3472) );
buf1 gate961( .a(N2970), .O(N3475) );
buf1 gate962( .a(N2967), .O(N3478) );
buf1 gate963( .a(N2970), .O(N3481) );
buf1 gate964( .a(N2973), .O(N3484) );
buf1 gate965( .a(N2973), .O(N3487) );
buf1 gate966( .a(N3172), .O(N3490) );
buf1 gate967( .a(N3172), .O(N3493) );
buf1 gate968( .a(N3175), .O(N3496) );
buf1 gate969( .a(N3175), .O(N3499) );
buf1 gate970( .a(N3178), .O(N3502) );
buf1 gate971( .a(N3178), .O(N3505) );
buf1 gate972( .a(N3181), .O(N3508) );
buf1 gate973( .a(N3181), .O(N3511) );
buf1 gate974( .a(N3184), .O(N3514) );
buf1 gate975( .a(N3184), .O(N3517) );
buf1 gate976( .a(N3187), .O(N3520) );
buf1 gate977( .a(N3187), .O(N3523) );
nor2 gate978( .a(N3387), .b(N2350), .O(N3534) );
or3 gate979( .a(N3388), .b(N2151), .c(N2351), .O(N3535) );

  xor2  gate2398(.a(N1966), .b(N3389), .O(gate980inter0));
  nand2 gate2399(.a(gate980inter0), .b(s_104), .O(gate980inter1));
  and2  gate2400(.a(N1966), .b(N3389), .O(gate980inter2));
  inv1  gate2401(.a(s_104), .O(gate980inter3));
  inv1  gate2402(.a(s_105), .O(gate980inter4));
  nand2 gate2403(.a(gate980inter4), .b(gate980inter3), .O(gate980inter5));
  nor2  gate2404(.a(gate980inter5), .b(gate980inter2), .O(gate980inter6));
  inv1  gate2405(.a(N3389), .O(gate980inter7));
  inv1  gate2406(.a(N1966), .O(gate980inter8));
  nand2 gate2407(.a(gate980inter8), .b(gate980inter7), .O(gate980inter9));
  nand2 gate2408(.a(s_105), .b(gate980inter3), .O(gate980inter10));
  nor2  gate2409(.a(gate980inter10), .b(gate980inter9), .O(gate980inter11));
  nor2  gate2410(.a(gate980inter11), .b(gate980inter6), .O(gate980inter12));
  nand2 gate2411(.a(gate980inter12), .b(gate980inter1), .O(N3536));
and2 gate981( .a(N3390), .b(N2209), .O(N3537) );
and2 gate982( .a(N3398), .b(N2210), .O(N3538) );
and2 gate983( .a(N3391), .b(N1842), .O(N3539) );
and2 gate984( .a(N3399), .b(N1369), .O(N3540) );
and2 gate985( .a(N3392), .b(N1843), .O(N3541) );
and2 gate986( .a(N3400), .b(N1369), .O(N3542) );
and2 gate987( .a(N3393), .b(N1844), .O(N3543) );
and2 gate988( .a(N3401), .b(N1369), .O(N3544) );
and2 gate989( .a(N3394), .b(N1845), .O(N3545) );
and2 gate990( .a(N3402), .b(N1369), .O(N3546) );
and2 gate991( .a(N3395), .b(N1846), .O(N3547) );
and2 gate992( .a(N3403), .b(N1369), .O(N3548) );
and2 gate993( .a(N3396), .b(N1847), .O(N3549) );
and2 gate994( .a(N3404), .b(N1369), .O(N3550) );
and2 gate995( .a(N3397), .b(N1848), .O(N3551) );
and2 gate996( .a(N3405), .b(N1369), .O(N3552) );
or3 gate997( .a(N3413), .b(N3414), .c(N3118), .O(N3557) );
or3 gate998( .a(N3429), .b(N3430), .c(N3134), .O(N3568) );
or3 gate999( .a(N3437), .b(N3438), .c(N3141), .O(N3573) );
or3 gate1000( .a(N3445), .b(N3446), .c(N3148), .O(N3578) );
or3 gate1001( .a(N3461), .b(N3462), .c(N3164), .O(N3589) );
or3 gate1002( .a(N3469), .b(N3470), .c(N3171), .O(N3594) );
and2 gate1003( .a(N3471), .b(N2728), .O(N3605) );
inv1 gate1004( .a(N3478), .O(N3626) );
inv1 gate1005( .a(N3481), .O(N3627) );
inv1 gate1006( .a(N3487), .O(N3628) );
inv1 gate1007( .a(N3484), .O(N3629) );
inv1 gate1008( .a(N3472), .O(N3630) );
inv1 gate1009( .a(N3475), .O(N3631) );
and2 gate1010( .a(N3536), .b(N2152), .O(N3632) );
and2 gate1011( .a(N3534), .b(N2155), .O(N3633) );
or3 gate1012( .a(N3537), .b(N3538), .c(N2398), .O(N3634) );
or2 gate1013( .a(N3539), .b(N3540), .O(N3635) );
or2 gate1014( .a(N3541), .b(N3542), .O(N3636) );
or2 gate1015( .a(N3543), .b(N3544), .O(N3637) );
or2 gate1016( .a(N3545), .b(N3546), .O(N3638) );
or2 gate1017( .a(N3547), .b(N3548), .O(N3639) );
or2 gate1018( .a(N3549), .b(N3550), .O(N3640) );
or2 gate1019( .a(N3551), .b(N3552), .O(N3641) );
and2 gate1020( .a(N3535), .b(N2643), .O(N3642) );
or2 gate1021( .a(N3407), .b(N3410), .O(N3643) );
nor2 gate1022( .a(N3407), .b(N3410), .O(N3644) );
and3 gate1023( .a(N169), .b(N3415), .c(N3122), .O(N3645) );
and3 gate1024( .a(N179), .b(N3415), .c(N3125), .O(N3648) );
and3 gate1025( .a(N190), .b(N3419), .c(N3125), .O(N3651) );
and3 gate1026( .a(N200), .b(N3419), .c(N3122), .O(N3652) );
inv1 gate1027( .a(N3419), .O(N3653) );
or2 gate1028( .a(N3423), .b(N3426), .O(N3654) );

  xor2  gate4288(.a(N3426), .b(N3423), .O(gate1029inter0));
  nand2 gate4289(.a(gate1029inter0), .b(s_374), .O(gate1029inter1));
  and2  gate4290(.a(N3426), .b(N3423), .O(gate1029inter2));
  inv1  gate4291(.a(s_374), .O(gate1029inter3));
  inv1  gate4292(.a(s_375), .O(gate1029inter4));
  nand2 gate4293(.a(gate1029inter4), .b(gate1029inter3), .O(gate1029inter5));
  nor2  gate4294(.a(gate1029inter5), .b(gate1029inter2), .O(gate1029inter6));
  inv1  gate4295(.a(N3423), .O(gate1029inter7));
  inv1  gate4296(.a(N3426), .O(gate1029inter8));
  nand2 gate4297(.a(gate1029inter8), .b(gate1029inter7), .O(gate1029inter9));
  nand2 gate4298(.a(s_375), .b(gate1029inter3), .O(gate1029inter10));
  nor2  gate4299(.a(gate1029inter10), .b(gate1029inter9), .O(gate1029inter11));
  nor2  gate4300(.a(gate1029inter11), .b(gate1029inter6), .O(gate1029inter12));
  nand2 gate4301(.a(gate1029inter12), .b(gate1029inter1), .O(N3657));
or2 gate1030( .a(N3431), .b(N3434), .O(N3658) );
nor2 gate1031( .a(N3431), .b(N3434), .O(N3661) );
or2 gate1032( .a(N3439), .b(N3442), .O(N3662) );

  xor2  gate4064(.a(N3442), .b(N3439), .O(gate1033inter0));
  nand2 gate4065(.a(gate1033inter0), .b(s_342), .O(gate1033inter1));
  and2  gate4066(.a(N3442), .b(N3439), .O(gate1033inter2));
  inv1  gate4067(.a(s_342), .O(gate1033inter3));
  inv1  gate4068(.a(s_343), .O(gate1033inter4));
  nand2 gate4069(.a(gate1033inter4), .b(gate1033inter3), .O(gate1033inter5));
  nor2  gate4070(.a(gate1033inter5), .b(gate1033inter2), .O(gate1033inter6));
  inv1  gate4071(.a(N3439), .O(gate1033inter7));
  inv1  gate4072(.a(N3442), .O(gate1033inter8));
  nand2 gate4073(.a(gate1033inter8), .b(gate1033inter7), .O(gate1033inter9));
  nand2 gate4074(.a(s_343), .b(gate1033inter3), .O(gate1033inter10));
  nor2  gate4075(.a(gate1033inter10), .b(gate1033inter9), .O(gate1033inter11));
  nor2  gate4076(.a(gate1033inter11), .b(gate1033inter6), .O(gate1033inter12));
  nand2 gate4077(.a(gate1033inter12), .b(gate1033inter1), .O(N3663));
and3 gate1034( .a(N169), .b(N3447), .c(N3152), .O(N3664) );
and3 gate1035( .a(N179), .b(N3447), .c(N3155), .O(N3667) );
and3 gate1036( .a(N190), .b(N3451), .c(N3155), .O(N3670) );
and3 gate1037( .a(N200), .b(N3451), .c(N3152), .O(N3671) );
inv1 gate1038( .a(N3451), .O(N3672) );
or2 gate1039( .a(N3455), .b(N3458), .O(N3673) );
nor2 gate1040( .a(N3455), .b(N3458), .O(N3676) );
or2 gate1041( .a(N3463), .b(N3466), .O(N3677) );
nor2 gate1042( .a(N3463), .b(N3466), .O(N3680) );
inv1 gate1043( .a(N3493), .O(N3681) );
and2 gate1044( .a(N1909), .b(N3415), .O(N3682) );
inv1 gate1045( .a(N3496), .O(N3685) );
inv1 gate1046( .a(N3499), .O(N3686) );
inv1 gate1047( .a(N3502), .O(N3687) );
inv1 gate1048( .a(N3505), .O(N3688) );
inv1 gate1049( .a(N3511), .O(N3689) );
and2 gate1050( .a(N1922), .b(N3447), .O(N3690) );
inv1 gate1051( .a(N3517), .O(N3693) );
inv1 gate1052( .a(N3520), .O(N3694) );
inv1 gate1053( .a(N3523), .O(N3695) );
inv1 gate1054( .a(N3514), .O(N3696) );
buf1 gate1055( .a(N3384), .O(N3697) );
buf1 gate1056( .a(N3384), .O(N3700) );
inv1 gate1057( .a(N3490), .O(N3703) );
inv1 gate1058( .a(N3508), .O(N3704) );

  xor2  gate4092(.a(N3630), .b(N3475), .O(gate1059inter0));
  nand2 gate4093(.a(gate1059inter0), .b(s_346), .O(gate1059inter1));
  and2  gate4094(.a(N3630), .b(N3475), .O(gate1059inter2));
  inv1  gate4095(.a(s_346), .O(gate1059inter3));
  inv1  gate4096(.a(s_347), .O(gate1059inter4));
  nand2 gate4097(.a(gate1059inter4), .b(gate1059inter3), .O(gate1059inter5));
  nor2  gate4098(.a(gate1059inter5), .b(gate1059inter2), .O(gate1059inter6));
  inv1  gate4099(.a(N3475), .O(gate1059inter7));
  inv1  gate4100(.a(N3630), .O(gate1059inter8));
  nand2 gate4101(.a(gate1059inter8), .b(gate1059inter7), .O(gate1059inter9));
  nand2 gate4102(.a(s_347), .b(gate1059inter3), .O(gate1059inter10));
  nor2  gate4103(.a(gate1059inter10), .b(gate1059inter9), .O(gate1059inter11));
  nor2  gate4104(.a(gate1059inter11), .b(gate1059inter6), .O(gate1059inter12));
  nand2 gate4105(.a(gate1059inter12), .b(gate1059inter1), .O(N3705));

  xor2  gate2258(.a(N3631), .b(N3472), .O(gate1060inter0));
  nand2 gate2259(.a(gate1060inter0), .b(s_84), .O(gate1060inter1));
  and2  gate2260(.a(N3631), .b(N3472), .O(gate1060inter2));
  inv1  gate2261(.a(s_84), .O(gate1060inter3));
  inv1  gate2262(.a(s_85), .O(gate1060inter4));
  nand2 gate2263(.a(gate1060inter4), .b(gate1060inter3), .O(gate1060inter5));
  nor2  gate2264(.a(gate1060inter5), .b(gate1060inter2), .O(gate1060inter6));
  inv1  gate2265(.a(N3472), .O(gate1060inter7));
  inv1  gate2266(.a(N3631), .O(gate1060inter8));
  nand2 gate2267(.a(gate1060inter8), .b(gate1060inter7), .O(gate1060inter9));
  nand2 gate2268(.a(s_85), .b(gate1060inter3), .O(gate1060inter10));
  nor2  gate2269(.a(gate1060inter10), .b(gate1060inter9), .O(gate1060inter11));
  nor2  gate2270(.a(gate1060inter11), .b(gate1060inter6), .O(gate1060inter12));
  nand2 gate2271(.a(gate1060inter12), .b(gate1060inter1), .O(N3706));
nand2 gate1061( .a(N3481), .b(N3626), .O(N3707) );
nand2 gate1062( .a(N3478), .b(N3627), .O(N3708) );
or3 gate1063( .a(N3632), .b(N2352), .c(N2353), .O(N3711) );
or3 gate1064( .a(N3633), .b(N2354), .c(N2355), .O(N3712) );
and2 gate1065( .a(N3634), .b(N2632), .O(N3713) );
and2 gate1066( .a(N3635), .b(N2634), .O(N3714) );
and2 gate1067( .a(N3636), .b(N2636), .O(N3715) );
and2 gate1068( .a(N3637), .b(N2638), .O(N3716) );
and2 gate1069( .a(N3638), .b(N2640), .O(N3717) );
and2 gate1070( .a(N3639), .b(N2642), .O(N3718) );
and2 gate1071( .a(N3640), .b(N2644), .O(N3719) );
and2 gate1072( .a(N3641), .b(N2646), .O(N3720) );
and2 gate1073( .a(N3644), .b(N3557), .O(N3721) );
or3 gate1074( .a(N3651), .b(N3652), .c(N3653), .O(N3731) );
and2 gate1075( .a(N3657), .b(N3568), .O(N3734) );
and2 gate1076( .a(N3661), .b(N3573), .O(N3740) );
and2 gate1077( .a(N3663), .b(N3578), .O(N3743) );
or3 gate1078( .a(N3670), .b(N3671), .c(N3672), .O(N3753) );
and2 gate1079( .a(N3676), .b(N3589), .O(N3756) );
and2 gate1080( .a(N3680), .b(N3594), .O(N3762) );
inv1 gate1081( .a(N3643), .O(N3765) );
inv1 gate1082( .a(N3662), .O(N3766) );

  xor2  gate3616(.a(N3706), .b(N3705), .O(gate1083inter0));
  nand2 gate3617(.a(gate1083inter0), .b(s_278), .O(gate1083inter1));
  and2  gate3618(.a(N3706), .b(N3705), .O(gate1083inter2));
  inv1  gate3619(.a(s_278), .O(gate1083inter3));
  inv1  gate3620(.a(s_279), .O(gate1083inter4));
  nand2 gate3621(.a(gate1083inter4), .b(gate1083inter3), .O(gate1083inter5));
  nor2  gate3622(.a(gate1083inter5), .b(gate1083inter2), .O(gate1083inter6));
  inv1  gate3623(.a(N3705), .O(gate1083inter7));
  inv1  gate3624(.a(N3706), .O(gate1083inter8));
  nand2 gate3625(.a(gate1083inter8), .b(gate1083inter7), .O(gate1083inter9));
  nand2 gate3626(.a(s_279), .b(gate1083inter3), .O(gate1083inter10));
  nor2  gate3627(.a(gate1083inter10), .b(gate1083inter9), .O(gate1083inter11));
  nor2  gate3628(.a(gate1083inter11), .b(gate1083inter6), .O(gate1083inter12));
  nand2 gate3629(.a(gate1083inter12), .b(gate1083inter1), .O(N3773));
nand2 gate1084( .a(N3707), .b(N3708), .O(N3774) );
nand2 gate1085( .a(N3700), .b(N3628), .O(N3775) );
inv1 gate1086( .a(N3700), .O(N3776) );
nand2 gate1087( .a(N3697), .b(N3629), .O(N3777) );
inv1 gate1088( .a(N3697), .O(N3778) );
and2 gate1089( .a(N3712), .b(N2645), .O(N3779) );
and2 gate1090( .a(N3711), .b(N2647), .O(N3780) );
or2 gate1091( .a(N3645), .b(N3648), .O(N3786) );
nor2 gate1092( .a(N3645), .b(N3648), .O(N3789) );
or2 gate1093( .a(N3664), .b(N3667), .O(N3800) );

  xor2  gate3014(.a(N3667), .b(N3664), .O(gate1094inter0));
  nand2 gate3015(.a(gate1094inter0), .b(s_192), .O(gate1094inter1));
  and2  gate3016(.a(N3667), .b(N3664), .O(gate1094inter2));
  inv1  gate3017(.a(s_192), .O(gate1094inter3));
  inv1  gate3018(.a(s_193), .O(gate1094inter4));
  nand2 gate3019(.a(gate1094inter4), .b(gate1094inter3), .O(gate1094inter5));
  nor2  gate3020(.a(gate1094inter5), .b(gate1094inter2), .O(gate1094inter6));
  inv1  gate3021(.a(N3664), .O(gate1094inter7));
  inv1  gate3022(.a(N3667), .O(gate1094inter8));
  nand2 gate3023(.a(gate1094inter8), .b(gate1094inter7), .O(gate1094inter9));
  nand2 gate3024(.a(s_193), .b(gate1094inter3), .O(gate1094inter10));
  nor2  gate3025(.a(gate1094inter10), .b(gate1094inter9), .O(gate1094inter11));
  nor2  gate3026(.a(gate1094inter11), .b(gate1094inter6), .O(gate1094inter12));
  nand2 gate3027(.a(gate1094inter12), .b(gate1094inter1), .O(N3803));
and2 gate1095( .a(N3654), .b(N1917), .O(N3809) );
and2 gate1096( .a(N3658), .b(N1917), .O(N3812) );
and2 gate1097( .a(N3673), .b(N1926), .O(N3815) );
and2 gate1098( .a(N3677), .b(N1926), .O(N3818) );
buf1 gate1099( .a(N3682), .O(N3821) );
buf1 gate1100( .a(N3682), .O(N3824) );
buf1 gate1101( .a(N3690), .O(N3827) );
buf1 gate1102( .a(N3690), .O(N3830) );

  xor2  gate3910(.a(N3774), .b(N3773), .O(gate1103inter0));
  nand2 gate3911(.a(gate1103inter0), .b(s_320), .O(gate1103inter1));
  and2  gate3912(.a(N3774), .b(N3773), .O(gate1103inter2));
  inv1  gate3913(.a(s_320), .O(gate1103inter3));
  inv1  gate3914(.a(s_321), .O(gate1103inter4));
  nand2 gate3915(.a(gate1103inter4), .b(gate1103inter3), .O(gate1103inter5));
  nor2  gate3916(.a(gate1103inter5), .b(gate1103inter2), .O(gate1103inter6));
  inv1  gate3917(.a(N3773), .O(gate1103inter7));
  inv1  gate3918(.a(N3774), .O(gate1103inter8));
  nand2 gate3919(.a(gate1103inter8), .b(gate1103inter7), .O(gate1103inter9));
  nand2 gate3920(.a(s_321), .b(gate1103inter3), .O(gate1103inter10));
  nor2  gate3921(.a(gate1103inter10), .b(gate1103inter9), .O(gate1103inter11));
  nor2  gate3922(.a(gate1103inter11), .b(gate1103inter6), .O(gate1103inter12));
  nand2 gate3923(.a(gate1103inter12), .b(gate1103inter1), .O(N3833));

  xor2  gate4400(.a(N3776), .b(N3487), .O(gate1104inter0));
  nand2 gate4401(.a(gate1104inter0), .b(s_390), .O(gate1104inter1));
  and2  gate4402(.a(N3776), .b(N3487), .O(gate1104inter2));
  inv1  gate4403(.a(s_390), .O(gate1104inter3));
  inv1  gate4404(.a(s_391), .O(gate1104inter4));
  nand2 gate4405(.a(gate1104inter4), .b(gate1104inter3), .O(gate1104inter5));
  nor2  gate4406(.a(gate1104inter5), .b(gate1104inter2), .O(gate1104inter6));
  inv1  gate4407(.a(N3487), .O(gate1104inter7));
  inv1  gate4408(.a(N3776), .O(gate1104inter8));
  nand2 gate4409(.a(gate1104inter8), .b(gate1104inter7), .O(gate1104inter9));
  nand2 gate4410(.a(s_391), .b(gate1104inter3), .O(gate1104inter10));
  nor2  gate4411(.a(gate1104inter10), .b(gate1104inter9), .O(gate1104inter11));
  nor2  gate4412(.a(gate1104inter11), .b(gate1104inter6), .O(gate1104inter12));
  nand2 gate4413(.a(gate1104inter12), .b(gate1104inter1), .O(N3834));
nand2 gate1105( .a(N3484), .b(N3778), .O(N3835) );
and2 gate1106( .a(N3789), .b(N3731), .O(N3838) );
and2 gate1107( .a(N3803), .b(N3753), .O(N3845) );
buf1 gate1108( .a(N3721), .O(N3850) );
buf1 gate1109( .a(N3734), .O(N3855) );
buf1 gate1110( .a(N3740), .O(N3858) );
buf1 gate1111( .a(N3743), .O(N3861) );
buf1 gate1112( .a(N3756), .O(N3865) );
buf1 gate1113( .a(N3762), .O(N3868) );

  xor2  gate2132(.a(N3834), .b(N3775), .O(gate1114inter0));
  nand2 gate2133(.a(gate1114inter0), .b(s_66), .O(gate1114inter1));
  and2  gate2134(.a(N3834), .b(N3775), .O(gate1114inter2));
  inv1  gate2135(.a(s_66), .O(gate1114inter3));
  inv1  gate2136(.a(s_67), .O(gate1114inter4));
  nand2 gate2137(.a(gate1114inter4), .b(gate1114inter3), .O(gate1114inter5));
  nor2  gate2138(.a(gate1114inter5), .b(gate1114inter2), .O(gate1114inter6));
  inv1  gate2139(.a(N3775), .O(gate1114inter7));
  inv1  gate2140(.a(N3834), .O(gate1114inter8));
  nand2 gate2141(.a(gate1114inter8), .b(gate1114inter7), .O(gate1114inter9));
  nand2 gate2142(.a(s_67), .b(gate1114inter3), .O(gate1114inter10));
  nor2  gate2143(.a(gate1114inter10), .b(gate1114inter9), .O(gate1114inter11));
  nor2  gate2144(.a(gate1114inter11), .b(gate1114inter6), .O(gate1114inter12));
  nand2 gate2145(.a(gate1114inter12), .b(gate1114inter1), .O(N3884));

  xor2  gate3252(.a(N3835), .b(N3777), .O(gate1115inter0));
  nand2 gate3253(.a(gate1115inter0), .b(s_226), .O(gate1115inter1));
  and2  gate3254(.a(N3835), .b(N3777), .O(gate1115inter2));
  inv1  gate3255(.a(s_226), .O(gate1115inter3));
  inv1  gate3256(.a(s_227), .O(gate1115inter4));
  nand2 gate3257(.a(gate1115inter4), .b(gate1115inter3), .O(gate1115inter5));
  nor2  gate3258(.a(gate1115inter5), .b(gate1115inter2), .O(gate1115inter6));
  inv1  gate3259(.a(N3777), .O(gate1115inter7));
  inv1  gate3260(.a(N3835), .O(gate1115inter8));
  nand2 gate3261(.a(gate1115inter8), .b(gate1115inter7), .O(gate1115inter9));
  nand2 gate3262(.a(s_227), .b(gate1115inter3), .O(gate1115inter10));
  nor2  gate3263(.a(gate1115inter10), .b(gate1115inter9), .O(gate1115inter11));
  nor2  gate3264(.a(gate1115inter11), .b(gate1115inter6), .O(gate1115inter12));
  nand2 gate3265(.a(gate1115inter12), .b(gate1115inter1), .O(N3885));
nand2 gate1116( .a(N3721), .b(N3786), .O(N3894) );

  xor2  gate3602(.a(N3800), .b(N3743), .O(gate1117inter0));
  nand2 gate3603(.a(gate1117inter0), .b(s_276), .O(gate1117inter1));
  and2  gate3604(.a(N3800), .b(N3743), .O(gate1117inter2));
  inv1  gate3605(.a(s_276), .O(gate1117inter3));
  inv1  gate3606(.a(s_277), .O(gate1117inter4));
  nand2 gate3607(.a(gate1117inter4), .b(gate1117inter3), .O(gate1117inter5));
  nor2  gate3608(.a(gate1117inter5), .b(gate1117inter2), .O(gate1117inter6));
  inv1  gate3609(.a(N3743), .O(gate1117inter7));
  inv1  gate3610(.a(N3800), .O(gate1117inter8));
  nand2 gate3611(.a(gate1117inter8), .b(gate1117inter7), .O(gate1117inter9));
  nand2 gate3612(.a(s_277), .b(gate1117inter3), .O(gate1117inter10));
  nor2  gate3613(.a(gate1117inter10), .b(gate1117inter9), .O(gate1117inter11));
  nor2  gate3614(.a(gate1117inter11), .b(gate1117inter6), .O(gate1117inter12));
  nand2 gate3615(.a(gate1117inter12), .b(gate1117inter1), .O(N3895));
inv1 gate1118( .a(N3821), .O(N3898) );
inv1 gate1119( .a(N3824), .O(N3899) );
inv1 gate1120( .a(N3830), .O(N3906) );
inv1 gate1121( .a(N3827), .O(N3911) );
and2 gate1122( .a(N3786), .b(N1912), .O(N3912) );
buf1 gate1123( .a(N3812), .O(N3913) );
and2 gate1124( .a(N3800), .b(N1917), .O(N3916) );
buf1 gate1125( .a(N3818), .O(N3917) );
inv1 gate1126( .a(N3809), .O(N3920) );
buf1 gate1127( .a(N3818), .O(N3921) );
inv1 gate1128( .a(N3884), .O(N3924) );
inv1 gate1129( .a(N3885), .O(N3925) );
and4 gate1130( .a(N3721), .b(N3838), .c(N3734), .d(N3740), .O(N3926) );
nand3 gate1131( .a(N3721), .b(N3838), .c(N3654), .O(N3930) );
nand4 gate1132( .a(N3658), .b(N3838), .c(N3734), .d(N3721), .O(N3931) );
and4 gate1133( .a(N3743), .b(N3845), .c(N3756), .d(N3762), .O(N3932) );
nand3 gate1134( .a(N3743), .b(N3845), .c(N3673), .O(N3935) );
nand4 gate1135( .a(N3677), .b(N3845), .c(N3756), .d(N3743), .O(N3936) );
buf1 gate1136( .a(N3838), .O(N3937) );
buf1 gate1137( .a(N3845), .O(N3940) );
inv1 gate1138( .a(N3912), .O(N3947) );
inv1 gate1139( .a(N3916), .O(N3948) );
buf1 gate1140( .a(N3850), .O(N3950) );
buf1 gate1141( .a(N3850), .O(N3953) );
buf1 gate1142( .a(N3855), .O(N3956) );
buf1 gate1143( .a(N3855), .O(N3959) );
buf1 gate1144( .a(N3858), .O(N3962) );
buf1 gate1145( .a(N3858), .O(N3965) );
buf1 gate1146( .a(N3861), .O(N3968) );
buf1 gate1147( .a(N3861), .O(N3971) );
buf1 gate1148( .a(N3865), .O(N3974) );
buf1 gate1149( .a(N3865), .O(N3977) );
buf1 gate1150( .a(N3868), .O(N3980) );
buf1 gate1151( .a(N3868), .O(N3983) );

  xor2  gate2566(.a(N3925), .b(N3924), .O(gate1152inter0));
  nand2 gate2567(.a(gate1152inter0), .b(s_128), .O(gate1152inter1));
  and2  gate2568(.a(N3925), .b(N3924), .O(gate1152inter2));
  inv1  gate2569(.a(s_128), .O(gate1152inter3));
  inv1  gate2570(.a(s_129), .O(gate1152inter4));
  nand2 gate2571(.a(gate1152inter4), .b(gate1152inter3), .O(gate1152inter5));
  nor2  gate2572(.a(gate1152inter5), .b(gate1152inter2), .O(gate1152inter6));
  inv1  gate2573(.a(N3924), .O(gate1152inter7));
  inv1  gate2574(.a(N3925), .O(gate1152inter8));
  nand2 gate2575(.a(gate1152inter8), .b(gate1152inter7), .O(gate1152inter9));
  nand2 gate2576(.a(s_129), .b(gate1152inter3), .O(gate1152inter10));
  nor2  gate2577(.a(gate1152inter10), .b(gate1152inter9), .O(gate1152inter11));
  nor2  gate2578(.a(gate1152inter11), .b(gate1152inter6), .O(gate1152inter12));
  nand2 gate2579(.a(gate1152inter12), .b(gate1152inter1), .O(N3987));
nand4 gate1153( .a(N3765), .b(N3894), .c(N3930), .d(N3931), .O(N3992) );
nand4 gate1154( .a(N3766), .b(N3895), .c(N3935), .d(N3936), .O(N3996) );
inv1 gate1155( .a(N3921), .O(N4013) );
and2 gate1156( .a(N3932), .b(N3926), .O(N4028) );

  xor2  gate2944(.a(N3681), .b(N3953), .O(gate1157inter0));
  nand2 gate2945(.a(gate1157inter0), .b(s_182), .O(gate1157inter1));
  and2  gate2946(.a(N3681), .b(N3953), .O(gate1157inter2));
  inv1  gate2947(.a(s_182), .O(gate1157inter3));
  inv1  gate2948(.a(s_183), .O(gate1157inter4));
  nand2 gate2949(.a(gate1157inter4), .b(gate1157inter3), .O(gate1157inter5));
  nor2  gate2950(.a(gate1157inter5), .b(gate1157inter2), .O(gate1157inter6));
  inv1  gate2951(.a(N3953), .O(gate1157inter7));
  inv1  gate2952(.a(N3681), .O(gate1157inter8));
  nand2 gate2953(.a(gate1157inter8), .b(gate1157inter7), .O(gate1157inter9));
  nand2 gate2954(.a(s_183), .b(gate1157inter3), .O(gate1157inter10));
  nor2  gate2955(.a(gate1157inter10), .b(gate1157inter9), .O(gate1157inter11));
  nor2  gate2956(.a(gate1157inter11), .b(gate1157inter6), .O(gate1157inter12));
  nand2 gate2957(.a(gate1157inter12), .b(gate1157inter1), .O(N4029));

  xor2  gate3350(.a(N3686), .b(N3959), .O(gate1158inter0));
  nand2 gate3351(.a(gate1158inter0), .b(s_240), .O(gate1158inter1));
  and2  gate3352(.a(N3686), .b(N3959), .O(gate1158inter2));
  inv1  gate3353(.a(s_240), .O(gate1158inter3));
  inv1  gate3354(.a(s_241), .O(gate1158inter4));
  nand2 gate3355(.a(gate1158inter4), .b(gate1158inter3), .O(gate1158inter5));
  nor2  gate3356(.a(gate1158inter5), .b(gate1158inter2), .O(gate1158inter6));
  inv1  gate3357(.a(N3959), .O(gate1158inter7));
  inv1  gate3358(.a(N3686), .O(gate1158inter8));
  nand2 gate3359(.a(gate1158inter8), .b(gate1158inter7), .O(gate1158inter9));
  nand2 gate3360(.a(s_241), .b(gate1158inter3), .O(gate1158inter10));
  nor2  gate3361(.a(gate1158inter10), .b(gate1158inter9), .O(gate1158inter11));
  nor2  gate3362(.a(gate1158inter11), .b(gate1158inter6), .O(gate1158inter12));
  nand2 gate3363(.a(gate1158inter12), .b(gate1158inter1), .O(N4030));

  xor2  gate3644(.a(N3688), .b(N3965), .O(gate1159inter0));
  nand2 gate3645(.a(gate1159inter0), .b(s_282), .O(gate1159inter1));
  and2  gate3646(.a(N3688), .b(N3965), .O(gate1159inter2));
  inv1  gate3647(.a(s_282), .O(gate1159inter3));
  inv1  gate3648(.a(s_283), .O(gate1159inter4));
  nand2 gate3649(.a(gate1159inter4), .b(gate1159inter3), .O(gate1159inter5));
  nor2  gate3650(.a(gate1159inter5), .b(gate1159inter2), .O(gate1159inter6));
  inv1  gate3651(.a(N3965), .O(gate1159inter7));
  inv1  gate3652(.a(N3688), .O(gate1159inter8));
  nand2 gate3653(.a(gate1159inter8), .b(gate1159inter7), .O(gate1159inter9));
  nand2 gate3654(.a(s_283), .b(gate1159inter3), .O(gate1159inter10));
  nor2  gate3655(.a(gate1159inter10), .b(gate1159inter9), .O(gate1159inter11));
  nor2  gate3656(.a(gate1159inter11), .b(gate1159inter6), .O(gate1159inter12));
  nand2 gate3657(.a(gate1159inter12), .b(gate1159inter1), .O(N4031));

  xor2  gate3868(.a(N3689), .b(N3971), .O(gate1160inter0));
  nand2 gate3869(.a(gate1160inter0), .b(s_314), .O(gate1160inter1));
  and2  gate3870(.a(N3689), .b(N3971), .O(gate1160inter2));
  inv1  gate3871(.a(s_314), .O(gate1160inter3));
  inv1  gate3872(.a(s_315), .O(gate1160inter4));
  nand2 gate3873(.a(gate1160inter4), .b(gate1160inter3), .O(gate1160inter5));
  nor2  gate3874(.a(gate1160inter5), .b(gate1160inter2), .O(gate1160inter6));
  inv1  gate3875(.a(N3971), .O(gate1160inter7));
  inv1  gate3876(.a(N3689), .O(gate1160inter8));
  nand2 gate3877(.a(gate1160inter8), .b(gate1160inter7), .O(gate1160inter9));
  nand2 gate3878(.a(s_315), .b(gate1160inter3), .O(gate1160inter10));
  nor2  gate3879(.a(gate1160inter10), .b(gate1160inter9), .O(gate1160inter11));
  nor2  gate3880(.a(gate1160inter11), .b(gate1160inter6), .O(gate1160inter12));
  nand2 gate3881(.a(gate1160inter12), .b(gate1160inter1), .O(N4032));

  xor2  gate2160(.a(N3693), .b(N3977), .O(gate1161inter0));
  nand2 gate2161(.a(gate1161inter0), .b(s_70), .O(gate1161inter1));
  and2  gate2162(.a(N3693), .b(N3977), .O(gate1161inter2));
  inv1  gate2163(.a(s_70), .O(gate1161inter3));
  inv1  gate2164(.a(s_71), .O(gate1161inter4));
  nand2 gate2165(.a(gate1161inter4), .b(gate1161inter3), .O(gate1161inter5));
  nor2  gate2166(.a(gate1161inter5), .b(gate1161inter2), .O(gate1161inter6));
  inv1  gate2167(.a(N3977), .O(gate1161inter7));
  inv1  gate2168(.a(N3693), .O(gate1161inter8));
  nand2 gate2169(.a(gate1161inter8), .b(gate1161inter7), .O(gate1161inter9));
  nand2 gate2170(.a(s_71), .b(gate1161inter3), .O(gate1161inter10));
  nor2  gate2171(.a(gate1161inter10), .b(gate1161inter9), .O(gate1161inter11));
  nor2  gate2172(.a(gate1161inter11), .b(gate1161inter6), .O(gate1161inter12));
  nand2 gate2173(.a(gate1161inter12), .b(gate1161inter1), .O(N4033));

  xor2  gate2580(.a(N3695), .b(N3983), .O(gate1162inter0));
  nand2 gate2581(.a(gate1162inter0), .b(s_130), .O(gate1162inter1));
  and2  gate2582(.a(N3695), .b(N3983), .O(gate1162inter2));
  inv1  gate2583(.a(s_130), .O(gate1162inter3));
  inv1  gate2584(.a(s_131), .O(gate1162inter4));
  nand2 gate2585(.a(gate1162inter4), .b(gate1162inter3), .O(gate1162inter5));
  nor2  gate2586(.a(gate1162inter5), .b(gate1162inter2), .O(gate1162inter6));
  inv1  gate2587(.a(N3983), .O(gate1162inter7));
  inv1  gate2588(.a(N3695), .O(gate1162inter8));
  nand2 gate2589(.a(gate1162inter8), .b(gate1162inter7), .O(gate1162inter9));
  nand2 gate2590(.a(s_131), .b(gate1162inter3), .O(gate1162inter10));
  nor2  gate2591(.a(gate1162inter10), .b(gate1162inter9), .O(gate1162inter11));
  nor2  gate2592(.a(gate1162inter11), .b(gate1162inter6), .O(gate1162inter12));
  nand2 gate2593(.a(gate1162inter12), .b(gate1162inter1), .O(N4034));
buf1 gate1163( .a(N3926), .O(N4035) );
inv1 gate1164( .a(N3953), .O(N4042) );
inv1 gate1165( .a(N3956), .O(N4043) );
nand2 gate1166( .a(N3956), .b(N3685), .O(N4044) );
inv1 gate1167( .a(N3959), .O(N4045) );
inv1 gate1168( .a(N3962), .O(N4046) );
nand2 gate1169( .a(N3962), .b(N3687), .O(N4047) );
inv1 gate1170( .a(N3965), .O(N4048) );
inv1 gate1171( .a(N3971), .O(N4049) );
inv1 gate1172( .a(N3977), .O(N4050) );
inv1 gate1173( .a(N3980), .O(N4051) );

  xor2  gate2776(.a(N3694), .b(N3980), .O(gate1174inter0));
  nand2 gate2777(.a(gate1174inter0), .b(s_158), .O(gate1174inter1));
  and2  gate2778(.a(N3694), .b(N3980), .O(gate1174inter2));
  inv1  gate2779(.a(s_158), .O(gate1174inter3));
  inv1  gate2780(.a(s_159), .O(gate1174inter4));
  nand2 gate2781(.a(gate1174inter4), .b(gate1174inter3), .O(gate1174inter5));
  nor2  gate2782(.a(gate1174inter5), .b(gate1174inter2), .O(gate1174inter6));
  inv1  gate2783(.a(N3980), .O(gate1174inter7));
  inv1  gate2784(.a(N3694), .O(gate1174inter8));
  nand2 gate2785(.a(gate1174inter8), .b(gate1174inter7), .O(gate1174inter9));
  nand2 gate2786(.a(s_159), .b(gate1174inter3), .O(gate1174inter10));
  nor2  gate2787(.a(gate1174inter10), .b(gate1174inter9), .O(gate1174inter11));
  nor2  gate2788(.a(gate1174inter11), .b(gate1174inter6), .O(gate1174inter12));
  nand2 gate2789(.a(gate1174inter12), .b(gate1174inter1), .O(N4052));
inv1 gate1175( .a(N3983), .O(N4053) );
inv1 gate1176( .a(N3974), .O(N4054) );

  xor2  gate2608(.a(N3696), .b(N3974), .O(gate1177inter0));
  nand2 gate2609(.a(gate1177inter0), .b(s_134), .O(gate1177inter1));
  and2  gate2610(.a(N3696), .b(N3974), .O(gate1177inter2));
  inv1  gate2611(.a(s_134), .O(gate1177inter3));
  inv1  gate2612(.a(s_135), .O(gate1177inter4));
  nand2 gate2613(.a(gate1177inter4), .b(gate1177inter3), .O(gate1177inter5));
  nor2  gate2614(.a(gate1177inter5), .b(gate1177inter2), .O(gate1177inter6));
  inv1  gate2615(.a(N3974), .O(gate1177inter7));
  inv1  gate2616(.a(N3696), .O(gate1177inter8));
  nand2 gate2617(.a(gate1177inter8), .b(gate1177inter7), .O(gate1177inter9));
  nand2 gate2618(.a(s_135), .b(gate1177inter3), .O(gate1177inter10));
  nor2  gate2619(.a(gate1177inter10), .b(gate1177inter9), .O(gate1177inter11));
  nor2  gate2620(.a(gate1177inter11), .b(gate1177inter6), .O(gate1177inter12));
  nand2 gate2621(.a(gate1177inter12), .b(gate1177inter1), .O(N4055));
and2 gate1178( .a(N3932), .b(N2304), .O(N4056) );
inv1 gate1179( .a(N3950), .O(N4057) );

  xor2  gate1964(.a(N3703), .b(N3950), .O(gate1180inter0));
  nand2 gate1965(.a(gate1180inter0), .b(s_42), .O(gate1180inter1));
  and2  gate1966(.a(N3703), .b(N3950), .O(gate1180inter2));
  inv1  gate1967(.a(s_42), .O(gate1180inter3));
  inv1  gate1968(.a(s_43), .O(gate1180inter4));
  nand2 gate1969(.a(gate1180inter4), .b(gate1180inter3), .O(gate1180inter5));
  nor2  gate1970(.a(gate1180inter5), .b(gate1180inter2), .O(gate1180inter6));
  inv1  gate1971(.a(N3950), .O(gate1180inter7));
  inv1  gate1972(.a(N3703), .O(gate1180inter8));
  nand2 gate1973(.a(gate1180inter8), .b(gate1180inter7), .O(gate1180inter9));
  nand2 gate1974(.a(s_43), .b(gate1180inter3), .O(gate1180inter10));
  nor2  gate1975(.a(gate1180inter10), .b(gate1180inter9), .O(gate1180inter11));
  nor2  gate1976(.a(gate1180inter11), .b(gate1180inter6), .O(gate1180inter12));
  nand2 gate1977(.a(gate1180inter12), .b(gate1180inter1), .O(N4058));
buf1 gate1181( .a(N3937), .O(N4059) );
buf1 gate1182( .a(N3937), .O(N4062) );
inv1 gate1183( .a(N3968), .O(N4065) );
nand2 gate1184( .a(N3968), .b(N3704), .O(N4066) );
buf1 gate1185( .a(N3940), .O(N4067) );
buf1 gate1186( .a(N3940), .O(N4070) );

  xor2  gate2832(.a(N3996), .b(N3926), .O(gate1187inter0));
  nand2 gate2833(.a(gate1187inter0), .b(s_166), .O(gate1187inter1));
  and2  gate2834(.a(N3996), .b(N3926), .O(gate1187inter2));
  inv1  gate2835(.a(s_166), .O(gate1187inter3));
  inv1  gate2836(.a(s_167), .O(gate1187inter4));
  nand2 gate2837(.a(gate1187inter4), .b(gate1187inter3), .O(gate1187inter5));
  nor2  gate2838(.a(gate1187inter5), .b(gate1187inter2), .O(gate1187inter6));
  inv1  gate2839(.a(N3926), .O(gate1187inter7));
  inv1  gate2840(.a(N3996), .O(gate1187inter8));
  nand2 gate2841(.a(gate1187inter8), .b(gate1187inter7), .O(gate1187inter9));
  nand2 gate2842(.a(s_167), .b(gate1187inter3), .O(gate1187inter10));
  nor2  gate2843(.a(gate1187inter10), .b(gate1187inter9), .O(gate1187inter11));
  nor2  gate2844(.a(gate1187inter11), .b(gate1187inter6), .O(gate1187inter12));
  nand2 gate2845(.a(gate1187inter12), .b(gate1187inter1), .O(N4073));
inv1 gate1188( .a(N3992), .O(N4074) );
nand2 gate1189( .a(N3493), .b(N4042), .O(N4075) );

  xor2  gate2048(.a(N4045), .b(N3499), .O(gate1190inter0));
  nand2 gate2049(.a(gate1190inter0), .b(s_54), .O(gate1190inter1));
  and2  gate2050(.a(N4045), .b(N3499), .O(gate1190inter2));
  inv1  gate2051(.a(s_54), .O(gate1190inter3));
  inv1  gate2052(.a(s_55), .O(gate1190inter4));
  nand2 gate2053(.a(gate1190inter4), .b(gate1190inter3), .O(gate1190inter5));
  nor2  gate2054(.a(gate1190inter5), .b(gate1190inter2), .O(gate1190inter6));
  inv1  gate2055(.a(N3499), .O(gate1190inter7));
  inv1  gate2056(.a(N4045), .O(gate1190inter8));
  nand2 gate2057(.a(gate1190inter8), .b(gate1190inter7), .O(gate1190inter9));
  nand2 gate2058(.a(s_55), .b(gate1190inter3), .O(gate1190inter10));
  nor2  gate2059(.a(gate1190inter10), .b(gate1190inter9), .O(gate1190inter11));
  nor2  gate2060(.a(gate1190inter11), .b(gate1190inter6), .O(gate1190inter12));
  nand2 gate2061(.a(gate1190inter12), .b(gate1190inter1), .O(N4076));

  xor2  gate3420(.a(N4048), .b(N3505), .O(gate1191inter0));
  nand2 gate3421(.a(gate1191inter0), .b(s_250), .O(gate1191inter1));
  and2  gate3422(.a(N4048), .b(N3505), .O(gate1191inter2));
  inv1  gate3423(.a(s_250), .O(gate1191inter3));
  inv1  gate3424(.a(s_251), .O(gate1191inter4));
  nand2 gate3425(.a(gate1191inter4), .b(gate1191inter3), .O(gate1191inter5));
  nor2  gate3426(.a(gate1191inter5), .b(gate1191inter2), .O(gate1191inter6));
  inv1  gate3427(.a(N3505), .O(gate1191inter7));
  inv1  gate3428(.a(N4048), .O(gate1191inter8));
  nand2 gate3429(.a(gate1191inter8), .b(gate1191inter7), .O(gate1191inter9));
  nand2 gate3430(.a(s_251), .b(gate1191inter3), .O(gate1191inter10));
  nor2  gate3431(.a(gate1191inter10), .b(gate1191inter9), .O(gate1191inter11));
  nor2  gate3432(.a(gate1191inter11), .b(gate1191inter6), .O(gate1191inter12));
  nand2 gate3433(.a(gate1191inter12), .b(gate1191inter1), .O(N4077));

  xor2  gate1894(.a(N4049), .b(N3511), .O(gate1192inter0));
  nand2 gate1895(.a(gate1192inter0), .b(s_32), .O(gate1192inter1));
  and2  gate1896(.a(N4049), .b(N3511), .O(gate1192inter2));
  inv1  gate1897(.a(s_32), .O(gate1192inter3));
  inv1  gate1898(.a(s_33), .O(gate1192inter4));
  nand2 gate1899(.a(gate1192inter4), .b(gate1192inter3), .O(gate1192inter5));
  nor2  gate1900(.a(gate1192inter5), .b(gate1192inter2), .O(gate1192inter6));
  inv1  gate1901(.a(N3511), .O(gate1192inter7));
  inv1  gate1902(.a(N4049), .O(gate1192inter8));
  nand2 gate1903(.a(gate1192inter8), .b(gate1192inter7), .O(gate1192inter9));
  nand2 gate1904(.a(s_33), .b(gate1192inter3), .O(gate1192inter10));
  nor2  gate1905(.a(gate1192inter10), .b(gate1192inter9), .O(gate1192inter11));
  nor2  gate1906(.a(gate1192inter11), .b(gate1192inter6), .O(gate1192inter12));
  nand2 gate1907(.a(gate1192inter12), .b(gate1192inter1), .O(N4078));
nand2 gate1193( .a(N3517), .b(N4050), .O(N4079) );
nand2 gate1194( .a(N3523), .b(N4053), .O(N4080) );

  xor2  gate2846(.a(N4043), .b(N3496), .O(gate1195inter0));
  nand2 gate2847(.a(gate1195inter0), .b(s_168), .O(gate1195inter1));
  and2  gate2848(.a(N4043), .b(N3496), .O(gate1195inter2));
  inv1  gate2849(.a(s_168), .O(gate1195inter3));
  inv1  gate2850(.a(s_169), .O(gate1195inter4));
  nand2 gate2851(.a(gate1195inter4), .b(gate1195inter3), .O(gate1195inter5));
  nor2  gate2852(.a(gate1195inter5), .b(gate1195inter2), .O(gate1195inter6));
  inv1  gate2853(.a(N3496), .O(gate1195inter7));
  inv1  gate2854(.a(N4043), .O(gate1195inter8));
  nand2 gate2855(.a(gate1195inter8), .b(gate1195inter7), .O(gate1195inter9));
  nand2 gate2856(.a(s_169), .b(gate1195inter3), .O(gate1195inter10));
  nor2  gate2857(.a(gate1195inter10), .b(gate1195inter9), .O(gate1195inter11));
  nor2  gate2858(.a(gate1195inter11), .b(gate1195inter6), .O(gate1195inter12));
  nand2 gate2859(.a(gate1195inter12), .b(gate1195inter1), .O(N4085));
nand2 gate1196( .a(N3502), .b(N4046), .O(N4086) );

  xor2  gate3798(.a(N4051), .b(N3520), .O(gate1197inter0));
  nand2 gate3799(.a(gate1197inter0), .b(s_304), .O(gate1197inter1));
  and2  gate3800(.a(N4051), .b(N3520), .O(gate1197inter2));
  inv1  gate3801(.a(s_304), .O(gate1197inter3));
  inv1  gate3802(.a(s_305), .O(gate1197inter4));
  nand2 gate3803(.a(gate1197inter4), .b(gate1197inter3), .O(gate1197inter5));
  nor2  gate3804(.a(gate1197inter5), .b(gate1197inter2), .O(gate1197inter6));
  inv1  gate3805(.a(N3520), .O(gate1197inter7));
  inv1  gate3806(.a(N4051), .O(gate1197inter8));
  nand2 gate3807(.a(gate1197inter8), .b(gate1197inter7), .O(gate1197inter9));
  nand2 gate3808(.a(s_305), .b(gate1197inter3), .O(gate1197inter10));
  nor2  gate3809(.a(gate1197inter10), .b(gate1197inter9), .O(gate1197inter11));
  nor2  gate3810(.a(gate1197inter11), .b(gate1197inter6), .O(gate1197inter12));
  nand2 gate3811(.a(gate1197inter12), .b(gate1197inter1), .O(N4088));
nand2 gate1198( .a(N3514), .b(N4054), .O(N4090) );
and2 gate1199( .a(N3996), .b(N1926), .O(N4091) );
or2 gate1200( .a(N3605), .b(N4056), .O(N4094) );

  xor2  gate2230(.a(N4057), .b(N3490), .O(gate1201inter0));
  nand2 gate2231(.a(gate1201inter0), .b(s_80), .O(gate1201inter1));
  and2  gate2232(.a(N4057), .b(N3490), .O(gate1201inter2));
  inv1  gate2233(.a(s_80), .O(gate1201inter3));
  inv1  gate2234(.a(s_81), .O(gate1201inter4));
  nand2 gate2235(.a(gate1201inter4), .b(gate1201inter3), .O(gate1201inter5));
  nor2  gate2236(.a(gate1201inter5), .b(gate1201inter2), .O(gate1201inter6));
  inv1  gate2237(.a(N3490), .O(gate1201inter7));
  inv1  gate2238(.a(N4057), .O(gate1201inter8));
  nand2 gate2239(.a(gate1201inter8), .b(gate1201inter7), .O(gate1201inter9));
  nand2 gate2240(.a(s_81), .b(gate1201inter3), .O(gate1201inter10));
  nor2  gate2241(.a(gate1201inter10), .b(gate1201inter9), .O(gate1201inter11));
  nor2  gate2242(.a(gate1201inter11), .b(gate1201inter6), .O(gate1201inter12));
  nand2 gate2243(.a(gate1201inter12), .b(gate1201inter1), .O(N4098));

  xor2  gate4386(.a(N4065), .b(N3508), .O(gate1202inter0));
  nand2 gate4387(.a(gate1202inter0), .b(s_388), .O(gate1202inter1));
  and2  gate4388(.a(N4065), .b(N3508), .O(gate1202inter2));
  inv1  gate4389(.a(s_388), .O(gate1202inter3));
  inv1  gate4390(.a(s_389), .O(gate1202inter4));
  nand2 gate4391(.a(gate1202inter4), .b(gate1202inter3), .O(gate1202inter5));
  nor2  gate4392(.a(gate1202inter5), .b(gate1202inter2), .O(gate1202inter6));
  inv1  gate4393(.a(N3508), .O(gate1202inter7));
  inv1  gate4394(.a(N4065), .O(gate1202inter8));
  nand2 gate4395(.a(gate1202inter8), .b(gate1202inter7), .O(gate1202inter9));
  nand2 gate4396(.a(s_389), .b(gate1202inter3), .O(gate1202inter10));
  nor2  gate4397(.a(gate1202inter10), .b(gate1202inter9), .O(gate1202inter11));
  nor2  gate4398(.a(gate1202inter11), .b(gate1202inter6), .O(gate1202inter12));
  nand2 gate4399(.a(gate1202inter12), .b(gate1202inter1), .O(N4101));
and2 gate1203( .a(N4073), .b(N4074), .O(N4104) );

  xor2  gate3182(.a(N4029), .b(N4075), .O(gate1204inter0));
  nand2 gate3183(.a(gate1204inter0), .b(s_216), .O(gate1204inter1));
  and2  gate3184(.a(N4029), .b(N4075), .O(gate1204inter2));
  inv1  gate3185(.a(s_216), .O(gate1204inter3));
  inv1  gate3186(.a(s_217), .O(gate1204inter4));
  nand2 gate3187(.a(gate1204inter4), .b(gate1204inter3), .O(gate1204inter5));
  nor2  gate3188(.a(gate1204inter5), .b(gate1204inter2), .O(gate1204inter6));
  inv1  gate3189(.a(N4075), .O(gate1204inter7));
  inv1  gate3190(.a(N4029), .O(gate1204inter8));
  nand2 gate3191(.a(gate1204inter8), .b(gate1204inter7), .O(gate1204inter9));
  nand2 gate3192(.a(s_217), .b(gate1204inter3), .O(gate1204inter10));
  nor2  gate3193(.a(gate1204inter10), .b(gate1204inter9), .O(gate1204inter11));
  nor2  gate3194(.a(gate1204inter11), .b(gate1204inter6), .O(gate1204inter12));
  nand2 gate3195(.a(gate1204inter12), .b(gate1204inter1), .O(N4105));

  xor2  gate3700(.a(N3899), .b(N4062), .O(gate1205inter0));
  nand2 gate3701(.a(gate1205inter0), .b(s_290), .O(gate1205inter1));
  and2  gate3702(.a(N3899), .b(N4062), .O(gate1205inter2));
  inv1  gate3703(.a(s_290), .O(gate1205inter3));
  inv1  gate3704(.a(s_291), .O(gate1205inter4));
  nand2 gate3705(.a(gate1205inter4), .b(gate1205inter3), .O(gate1205inter5));
  nor2  gate3706(.a(gate1205inter5), .b(gate1205inter2), .O(gate1205inter6));
  inv1  gate3707(.a(N4062), .O(gate1205inter7));
  inv1  gate3708(.a(N3899), .O(gate1205inter8));
  nand2 gate3709(.a(gate1205inter8), .b(gate1205inter7), .O(gate1205inter9));
  nand2 gate3710(.a(s_291), .b(gate1205inter3), .O(gate1205inter10));
  nor2  gate3711(.a(gate1205inter10), .b(gate1205inter9), .O(gate1205inter11));
  nor2  gate3712(.a(gate1205inter11), .b(gate1205inter6), .O(gate1205inter12));
  nand2 gate3713(.a(gate1205inter12), .b(gate1205inter1), .O(N4106));

  xor2  gate3826(.a(N4030), .b(N4076), .O(gate1206inter0));
  nand2 gate3827(.a(gate1206inter0), .b(s_308), .O(gate1206inter1));
  and2  gate3828(.a(N4030), .b(N4076), .O(gate1206inter2));
  inv1  gate3829(.a(s_308), .O(gate1206inter3));
  inv1  gate3830(.a(s_309), .O(gate1206inter4));
  nand2 gate3831(.a(gate1206inter4), .b(gate1206inter3), .O(gate1206inter5));
  nor2  gate3832(.a(gate1206inter5), .b(gate1206inter2), .O(gate1206inter6));
  inv1  gate3833(.a(N4076), .O(gate1206inter7));
  inv1  gate3834(.a(N4030), .O(gate1206inter8));
  nand2 gate3835(.a(gate1206inter8), .b(gate1206inter7), .O(gate1206inter9));
  nand2 gate3836(.a(s_309), .b(gate1206inter3), .O(gate1206inter10));
  nor2  gate3837(.a(gate1206inter10), .b(gate1206inter9), .O(gate1206inter11));
  nor2  gate3838(.a(gate1206inter11), .b(gate1206inter6), .O(gate1206inter12));
  nand2 gate3839(.a(gate1206inter12), .b(gate1206inter1), .O(N4107));

  xor2  gate3840(.a(N4031), .b(N4077), .O(gate1207inter0));
  nand2 gate3841(.a(gate1207inter0), .b(s_310), .O(gate1207inter1));
  and2  gate3842(.a(N4031), .b(N4077), .O(gate1207inter2));
  inv1  gate3843(.a(s_310), .O(gate1207inter3));
  inv1  gate3844(.a(s_311), .O(gate1207inter4));
  nand2 gate3845(.a(gate1207inter4), .b(gate1207inter3), .O(gate1207inter5));
  nor2  gate3846(.a(gate1207inter5), .b(gate1207inter2), .O(gate1207inter6));
  inv1  gate3847(.a(N4077), .O(gate1207inter7));
  inv1  gate3848(.a(N4031), .O(gate1207inter8));
  nand2 gate3849(.a(gate1207inter8), .b(gate1207inter7), .O(gate1207inter9));
  nand2 gate3850(.a(s_311), .b(gate1207inter3), .O(gate1207inter10));
  nor2  gate3851(.a(gate1207inter10), .b(gate1207inter9), .O(gate1207inter11));
  nor2  gate3852(.a(gate1207inter11), .b(gate1207inter6), .O(gate1207inter12));
  nand2 gate3853(.a(gate1207inter12), .b(gate1207inter1), .O(N4108));
nand2 gate1208( .a(N4078), .b(N4032), .O(N4109) );
nand2 gate1209( .a(N4070), .b(N3906), .O(N4110) );

  xor2  gate4218(.a(N4033), .b(N4079), .O(gate1210inter0));
  nand2 gate4219(.a(gate1210inter0), .b(s_364), .O(gate1210inter1));
  and2  gate4220(.a(N4033), .b(N4079), .O(gate1210inter2));
  inv1  gate4221(.a(s_364), .O(gate1210inter3));
  inv1  gate4222(.a(s_365), .O(gate1210inter4));
  nand2 gate4223(.a(gate1210inter4), .b(gate1210inter3), .O(gate1210inter5));
  nor2  gate4224(.a(gate1210inter5), .b(gate1210inter2), .O(gate1210inter6));
  inv1  gate4225(.a(N4079), .O(gate1210inter7));
  inv1  gate4226(.a(N4033), .O(gate1210inter8));
  nand2 gate4227(.a(gate1210inter8), .b(gate1210inter7), .O(gate1210inter9));
  nand2 gate4228(.a(s_365), .b(gate1210inter3), .O(gate1210inter10));
  nor2  gate4229(.a(gate1210inter10), .b(gate1210inter9), .O(gate1210inter11));
  nor2  gate4230(.a(gate1210inter11), .b(gate1210inter6), .O(gate1210inter12));
  nand2 gate4231(.a(gate1210inter12), .b(gate1210inter1), .O(N4111));
nand2 gate1211( .a(N4080), .b(N4034), .O(N4112) );
inv1 gate1212( .a(N4059), .O(N4113) );

  xor2  gate1992(.a(N3898), .b(N4059), .O(gate1213inter0));
  nand2 gate1993(.a(gate1213inter0), .b(s_46), .O(gate1213inter1));
  and2  gate1994(.a(N3898), .b(N4059), .O(gate1213inter2));
  inv1  gate1995(.a(s_46), .O(gate1213inter3));
  inv1  gate1996(.a(s_47), .O(gate1213inter4));
  nand2 gate1997(.a(gate1213inter4), .b(gate1213inter3), .O(gate1213inter5));
  nor2  gate1998(.a(gate1213inter5), .b(gate1213inter2), .O(gate1213inter6));
  inv1  gate1999(.a(N4059), .O(gate1213inter7));
  inv1  gate2000(.a(N3898), .O(gate1213inter8));
  nand2 gate2001(.a(gate1213inter8), .b(gate1213inter7), .O(gate1213inter9));
  nand2 gate2002(.a(s_47), .b(gate1213inter3), .O(gate1213inter10));
  nor2  gate2003(.a(gate1213inter10), .b(gate1213inter9), .O(gate1213inter11));
  nor2  gate2004(.a(gate1213inter11), .b(gate1213inter6), .O(gate1213inter12));
  nand2 gate2005(.a(gate1213inter12), .b(gate1213inter1), .O(N4114));
inv1 gate1214( .a(N4062), .O(N4115) );
nand2 gate1215( .a(N4085), .b(N4044), .O(N4116) );
nand2 gate1216( .a(N4086), .b(N4047), .O(N4119) );
inv1 gate1217( .a(N4070), .O(N4122) );
nand2 gate1218( .a(N4088), .b(N4052), .O(N4123) );
inv1 gate1219( .a(N4067), .O(N4126) );

  xor2  gate3686(.a(N3911), .b(N4067), .O(gate1220inter0));
  nand2 gate3687(.a(gate1220inter0), .b(s_288), .O(gate1220inter1));
  and2  gate3688(.a(N3911), .b(N4067), .O(gate1220inter2));
  inv1  gate3689(.a(s_288), .O(gate1220inter3));
  inv1  gate3690(.a(s_289), .O(gate1220inter4));
  nand2 gate3691(.a(gate1220inter4), .b(gate1220inter3), .O(gate1220inter5));
  nor2  gate3692(.a(gate1220inter5), .b(gate1220inter2), .O(gate1220inter6));
  inv1  gate3693(.a(N4067), .O(gate1220inter7));
  inv1  gate3694(.a(N3911), .O(gate1220inter8));
  nand2 gate3695(.a(gate1220inter8), .b(gate1220inter7), .O(gate1220inter9));
  nand2 gate3696(.a(s_289), .b(gate1220inter3), .O(gate1220inter10));
  nor2  gate3697(.a(gate1220inter10), .b(gate1220inter9), .O(gate1220inter11));
  nor2  gate3698(.a(gate1220inter11), .b(gate1220inter6), .O(gate1220inter12));
  nand2 gate3699(.a(gate1220inter12), .b(gate1220inter1), .O(N4127));

  xor2  gate2412(.a(N4055), .b(N4090), .O(gate1221inter0));
  nand2 gate2413(.a(gate1221inter0), .b(s_106), .O(gate1221inter1));
  and2  gate2414(.a(N4055), .b(N4090), .O(gate1221inter2));
  inv1  gate2415(.a(s_106), .O(gate1221inter3));
  inv1  gate2416(.a(s_107), .O(gate1221inter4));
  nand2 gate2417(.a(gate1221inter4), .b(gate1221inter3), .O(gate1221inter5));
  nor2  gate2418(.a(gate1221inter5), .b(gate1221inter2), .O(gate1221inter6));
  inv1  gate2419(.a(N4090), .O(gate1221inter7));
  inv1  gate2420(.a(N4055), .O(gate1221inter8));
  nand2 gate2421(.a(gate1221inter8), .b(gate1221inter7), .O(gate1221inter9));
  nand2 gate2422(.a(s_107), .b(gate1221inter3), .O(gate1221inter10));
  nor2  gate2423(.a(gate1221inter10), .b(gate1221inter9), .O(gate1221inter11));
  nor2  gate2424(.a(gate1221inter11), .b(gate1221inter6), .O(gate1221inter12));
  nand2 gate2425(.a(gate1221inter12), .b(gate1221inter1), .O(N4128));

  xor2  gate3308(.a(N4058), .b(N4098), .O(gate1222inter0));
  nand2 gate3309(.a(gate1222inter0), .b(s_234), .O(gate1222inter1));
  and2  gate3310(.a(N4058), .b(N4098), .O(gate1222inter2));
  inv1  gate3311(.a(s_234), .O(gate1222inter3));
  inv1  gate3312(.a(s_235), .O(gate1222inter4));
  nand2 gate3313(.a(gate1222inter4), .b(gate1222inter3), .O(gate1222inter5));
  nor2  gate3314(.a(gate1222inter5), .b(gate1222inter2), .O(gate1222inter6));
  inv1  gate3315(.a(N4098), .O(gate1222inter7));
  inv1  gate3316(.a(N4058), .O(gate1222inter8));
  nand2 gate3317(.a(gate1222inter8), .b(gate1222inter7), .O(gate1222inter9));
  nand2 gate3318(.a(s_235), .b(gate1222inter3), .O(gate1222inter10));
  nor2  gate3319(.a(gate1222inter10), .b(gate1222inter9), .O(gate1222inter11));
  nor2  gate3320(.a(gate1222inter11), .b(gate1222inter6), .O(gate1222inter12));
  nand2 gate3321(.a(gate1222inter12), .b(gate1222inter1), .O(N4139));

  xor2  gate2552(.a(N4066), .b(N4101), .O(gate1223inter0));
  nand2 gate2553(.a(gate1223inter0), .b(s_126), .O(gate1223inter1));
  and2  gate2554(.a(N4066), .b(N4101), .O(gate1223inter2));
  inv1  gate2555(.a(s_126), .O(gate1223inter3));
  inv1  gate2556(.a(s_127), .O(gate1223inter4));
  nand2 gate2557(.a(gate1223inter4), .b(gate1223inter3), .O(gate1223inter5));
  nor2  gate2558(.a(gate1223inter5), .b(gate1223inter2), .O(gate1223inter6));
  inv1  gate2559(.a(N4101), .O(gate1223inter7));
  inv1  gate2560(.a(N4066), .O(gate1223inter8));
  nand2 gate2561(.a(gate1223inter8), .b(gate1223inter7), .O(gate1223inter9));
  nand2 gate2562(.a(s_127), .b(gate1223inter3), .O(gate1223inter10));
  nor2  gate2563(.a(gate1223inter10), .b(gate1223inter9), .O(gate1223inter11));
  nor2  gate2564(.a(gate1223inter11), .b(gate1223inter6), .O(gate1223inter12));
  nand2 gate2565(.a(gate1223inter12), .b(gate1223inter1), .O(N4142));
inv1 gate1224( .a(N4104), .O(N4145) );
inv1 gate1225( .a(N4105), .O(N4146) );

  xor2  gate3168(.a(N4115), .b(N3824), .O(gate1226inter0));
  nand2 gate3169(.a(gate1226inter0), .b(s_214), .O(gate1226inter1));
  and2  gate3170(.a(N4115), .b(N3824), .O(gate1226inter2));
  inv1  gate3171(.a(s_214), .O(gate1226inter3));
  inv1  gate3172(.a(s_215), .O(gate1226inter4));
  nand2 gate3173(.a(gate1226inter4), .b(gate1226inter3), .O(gate1226inter5));
  nor2  gate3174(.a(gate1226inter5), .b(gate1226inter2), .O(gate1226inter6));
  inv1  gate3175(.a(N3824), .O(gate1226inter7));
  inv1  gate3176(.a(N4115), .O(gate1226inter8));
  nand2 gate3177(.a(gate1226inter8), .b(gate1226inter7), .O(gate1226inter9));
  nand2 gate3178(.a(s_215), .b(gate1226inter3), .O(gate1226inter10));
  nor2  gate3179(.a(gate1226inter10), .b(gate1226inter9), .O(gate1226inter11));
  nor2  gate3180(.a(gate1226inter11), .b(gate1226inter6), .O(gate1226inter12));
  nand2 gate3181(.a(gate1226inter12), .b(gate1226inter1), .O(N4147));
inv1 gate1227( .a(N4107), .O(N4148) );
inv1 gate1228( .a(N4108), .O(N4149) );
inv1 gate1229( .a(N4109), .O(N4150) );

  xor2  gate1838(.a(N4122), .b(N3830), .O(gate1230inter0));
  nand2 gate1839(.a(gate1230inter0), .b(s_24), .O(gate1230inter1));
  and2  gate1840(.a(N4122), .b(N3830), .O(gate1230inter2));
  inv1  gate1841(.a(s_24), .O(gate1230inter3));
  inv1  gate1842(.a(s_25), .O(gate1230inter4));
  nand2 gate1843(.a(gate1230inter4), .b(gate1230inter3), .O(gate1230inter5));
  nor2  gate1844(.a(gate1230inter5), .b(gate1230inter2), .O(gate1230inter6));
  inv1  gate1845(.a(N3830), .O(gate1230inter7));
  inv1  gate1846(.a(N4122), .O(gate1230inter8));
  nand2 gate1847(.a(gate1230inter8), .b(gate1230inter7), .O(gate1230inter9));
  nand2 gate1848(.a(s_25), .b(gate1230inter3), .O(gate1230inter10));
  nor2  gate1849(.a(gate1230inter10), .b(gate1230inter9), .O(gate1230inter11));
  nor2  gate1850(.a(gate1230inter11), .b(gate1230inter6), .O(gate1230inter12));
  nand2 gate1851(.a(gate1230inter12), .b(gate1230inter1), .O(N4151));
inv1 gate1231( .a(N4111), .O(N4152) );
inv1 gate1232( .a(N4112), .O(N4153) );

  xor2  gate3364(.a(N4113), .b(N3821), .O(gate1233inter0));
  nand2 gate3365(.a(gate1233inter0), .b(s_242), .O(gate1233inter1));
  and2  gate3366(.a(N4113), .b(N3821), .O(gate1233inter2));
  inv1  gate3367(.a(s_242), .O(gate1233inter3));
  inv1  gate3368(.a(s_243), .O(gate1233inter4));
  nand2 gate3369(.a(gate1233inter4), .b(gate1233inter3), .O(gate1233inter5));
  nor2  gate3370(.a(gate1233inter5), .b(gate1233inter2), .O(gate1233inter6));
  inv1  gate3371(.a(N3821), .O(gate1233inter7));
  inv1  gate3372(.a(N4113), .O(gate1233inter8));
  nand2 gate3373(.a(gate1233inter8), .b(gate1233inter7), .O(gate1233inter9));
  nand2 gate3374(.a(s_243), .b(gate1233inter3), .O(gate1233inter10));
  nor2  gate3375(.a(gate1233inter10), .b(gate1233inter9), .O(gate1233inter11));
  nor2  gate3376(.a(gate1233inter11), .b(gate1233inter6), .O(gate1233inter12));
  nand2 gate3377(.a(gate1233inter12), .b(gate1233inter1), .O(N4154));
nand2 gate1234( .a(N3827), .b(N4126), .O(N4161) );
buf1 gate1235( .a(N4091), .O(N4167) );
buf1 gate1236( .a(N4094), .O(N4174) );
buf1 gate1237( .a(N4091), .O(N4182) );
and2 gate1238( .a(N330), .b(N4094), .O(N4186) );
and2 gate1239( .a(N4146), .b(N2230), .O(N4189) );

  xor2  gate4274(.a(N4106), .b(N4147), .O(gate1240inter0));
  nand2 gate4275(.a(gate1240inter0), .b(s_372), .O(gate1240inter1));
  and2  gate4276(.a(N4106), .b(N4147), .O(gate1240inter2));
  inv1  gate4277(.a(s_372), .O(gate1240inter3));
  inv1  gate4278(.a(s_373), .O(gate1240inter4));
  nand2 gate4279(.a(gate1240inter4), .b(gate1240inter3), .O(gate1240inter5));
  nor2  gate4280(.a(gate1240inter5), .b(gate1240inter2), .O(gate1240inter6));
  inv1  gate4281(.a(N4147), .O(gate1240inter7));
  inv1  gate4282(.a(N4106), .O(gate1240inter8));
  nand2 gate4283(.a(gate1240inter8), .b(gate1240inter7), .O(gate1240inter9));
  nand2 gate4284(.a(s_373), .b(gate1240inter3), .O(gate1240inter10));
  nor2  gate4285(.a(gate1240inter10), .b(gate1240inter9), .O(gate1240inter11));
  nor2  gate4286(.a(gate1240inter11), .b(gate1240inter6), .O(gate1240inter12));
  nand2 gate4287(.a(gate1240inter12), .b(gate1240inter1), .O(N4190));
and2 gate1241( .a(N4148), .b(N2232), .O(N4191) );
and2 gate1242( .a(N4149), .b(N2233), .O(N4192) );
and2 gate1243( .a(N4150), .b(N2234), .O(N4193) );
nand2 gate1244( .a(N4151), .b(N4110), .O(N4194) );
and2 gate1245( .a(N4152), .b(N2236), .O(N4195) );
and2 gate1246( .a(N4153), .b(N2237), .O(N4196) );

  xor2  gate2202(.a(N4114), .b(N4154), .O(gate1247inter0));
  nand2 gate2203(.a(gate1247inter0), .b(s_76), .O(gate1247inter1));
  and2  gate2204(.a(N4114), .b(N4154), .O(gate1247inter2));
  inv1  gate2205(.a(s_76), .O(gate1247inter3));
  inv1  gate2206(.a(s_77), .O(gate1247inter4));
  nand2 gate2207(.a(gate1247inter4), .b(gate1247inter3), .O(gate1247inter5));
  nor2  gate2208(.a(gate1247inter5), .b(gate1247inter2), .O(gate1247inter6));
  inv1  gate2209(.a(N4154), .O(gate1247inter7));
  inv1  gate2210(.a(N4114), .O(gate1247inter8));
  nand2 gate2211(.a(gate1247inter8), .b(gate1247inter7), .O(gate1247inter9));
  nand2 gate2212(.a(s_77), .b(gate1247inter3), .O(gate1247inter10));
  nor2  gate2213(.a(gate1247inter10), .b(gate1247inter9), .O(gate1247inter11));
  nor2  gate2214(.a(gate1247inter11), .b(gate1247inter6), .O(gate1247inter12));
  nand2 gate2215(.a(gate1247inter12), .b(gate1247inter1), .O(N4197));
buf1 gate1248( .a(N4116), .O(N4200) );
buf1 gate1249( .a(N4116), .O(N4203) );
buf1 gate1250( .a(N4119), .O(N4209) );
buf1 gate1251( .a(N4119), .O(N4213) );
nand2 gate1252( .a(N4161), .b(N4127), .O(N4218) );
buf1 gate1253( .a(N4123), .O(N4223) );
and2 gate1254( .a(N4128), .b(N3917), .O(N4238) );
inv1 gate1255( .a(N4139), .O(N4239) );
inv1 gate1256( .a(N4142), .O(N4241) );
and2 gate1257( .a(N330), .b(N4123), .O(N4242) );
buf1 gate1258( .a(N4128), .O(N4247) );
nor3 gate1259( .a(N3713), .b(N4189), .c(N2898), .O(N4251) );
inv1 gate1260( .a(N4190), .O(N4252) );
nor3 gate1261( .a(N3715), .b(N4191), .c(N2900), .O(N4253) );
nor3 gate1262( .a(N3716), .b(N4192), .c(N2901), .O(N4254) );
nor3 gate1263( .a(N3717), .b(N4193), .c(N3406), .O(N4255) );
inv1 gate1264( .a(N4194), .O(N4256) );
nor3 gate1265( .a(N3719), .b(N4195), .c(N3779), .O(N4257) );
nor3 gate1266( .a(N3720), .b(N4196), .c(N3780), .O(N4258) );
and2 gate1267( .a(N4167), .b(N4035), .O(N4283) );
and2 gate1268( .a(N4174), .b(N4035), .O(N4284) );
or2 gate1269( .a(N3815), .b(N4238), .O(N4287) );
inv1 gate1270( .a(N4186), .O(N4291) );
inv1 gate1271( .a(N4167), .O(N4295) );
buf1 gate1272( .a(N4167), .O(N4296) );
inv1 gate1273( .a(N4182), .O(N4299) );
and2 gate1274( .a(N4252), .b(N2231), .O(N4303) );
and2 gate1275( .a(N4256), .b(N2235), .O(N4304) );
buf1 gate1276( .a(N4197), .O(N4305) );
or2 gate1277( .a(N3992), .b(N4283), .O(N4310) );
and3 gate1278( .a(N4174), .b(N4213), .c(N4203), .O(N4316) );
and2 gate1279( .a(N4174), .b(N4209), .O(N4317) );
and3 gate1280( .a(N4223), .b(N4128), .c(N4218), .O(N4318) );
and2 gate1281( .a(N4223), .b(N4128), .O(N4319) );
and2 gate1282( .a(N4167), .b(N4209), .O(N4322) );

  xor2  gate2930(.a(N3913), .b(N4203), .O(gate1283inter0));
  nand2 gate2931(.a(gate1283inter0), .b(s_180), .O(gate1283inter1));
  and2  gate2932(.a(N3913), .b(N4203), .O(gate1283inter2));
  inv1  gate2933(.a(s_180), .O(gate1283inter3));
  inv1  gate2934(.a(s_181), .O(gate1283inter4));
  nand2 gate2935(.a(gate1283inter4), .b(gate1283inter3), .O(gate1283inter5));
  nor2  gate2936(.a(gate1283inter5), .b(gate1283inter2), .O(gate1283inter6));
  inv1  gate2937(.a(N4203), .O(gate1283inter7));
  inv1  gate2938(.a(N3913), .O(gate1283inter8));
  nand2 gate2939(.a(gate1283inter8), .b(gate1283inter7), .O(gate1283inter9));
  nand2 gate2940(.a(s_181), .b(gate1283inter3), .O(gate1283inter10));
  nor2  gate2941(.a(gate1283inter10), .b(gate1283inter9), .O(gate1283inter11));
  nor2  gate2942(.a(gate1283inter11), .b(gate1283inter6), .O(gate1283inter12));
  nand2 gate2943(.a(gate1283inter12), .b(gate1283inter1), .O(N4325));
nand3 gate1284( .a(N4203), .b(N4213), .c(N4167), .O(N4326) );
nand2 gate1285( .a(N4218), .b(N3815), .O(N4327) );
nand3 gate1286( .a(N4218), .b(N4128), .c(N3917), .O(N4328) );

  xor2  gate2734(.a(N4013), .b(N4247), .O(gate1287inter0));
  nand2 gate2735(.a(gate1287inter0), .b(s_152), .O(gate1287inter1));
  and2  gate2736(.a(N4013), .b(N4247), .O(gate1287inter2));
  inv1  gate2737(.a(s_152), .O(gate1287inter3));
  inv1  gate2738(.a(s_153), .O(gate1287inter4));
  nand2 gate2739(.a(gate1287inter4), .b(gate1287inter3), .O(gate1287inter5));
  nor2  gate2740(.a(gate1287inter5), .b(gate1287inter2), .O(gate1287inter6));
  inv1  gate2741(.a(N4247), .O(gate1287inter7));
  inv1  gate2742(.a(N4013), .O(gate1287inter8));
  nand2 gate2743(.a(gate1287inter8), .b(gate1287inter7), .O(gate1287inter9));
  nand2 gate2744(.a(s_153), .b(gate1287inter3), .O(gate1287inter10));
  nor2  gate2745(.a(gate1287inter10), .b(gate1287inter9), .O(gate1287inter11));
  nor2  gate2746(.a(gate1287inter11), .b(gate1287inter6), .O(gate1287inter12));
  nand2 gate2747(.a(gate1287inter12), .b(gate1287inter1), .O(N4329));
inv1 gate1288( .a(N4247), .O(N4330) );
and3 gate1289( .a(N330), .b(N4094), .c(N4295), .O(N4331) );
and2 gate1290( .a(N4251), .b(N2730), .O(N4335) );
and2 gate1291( .a(N4253), .b(N2734), .O(N4338) );
and2 gate1292( .a(N4254), .b(N2736), .O(N4341) );
and2 gate1293( .a(N4255), .b(N2738), .O(N4344) );
and2 gate1294( .a(N4257), .b(N2742), .O(N4347) );
and2 gate1295( .a(N4258), .b(N2744), .O(N4350) );
buf1 gate1296( .a(N4197), .O(N4353) );
buf1 gate1297( .a(N4203), .O(N4356) );
buf1 gate1298( .a(N4209), .O(N4359) );
buf1 gate1299( .a(N4218), .O(N4362) );
buf1 gate1300( .a(N4242), .O(N4365) );
buf1 gate1301( .a(N4242), .O(N4368) );
and2 gate1302( .a(N4223), .b(N4223), .O(N4371) );
nor3 gate1303( .a(N3714), .b(N4303), .c(N2899), .O(N4376) );
nor3 gate1304( .a(N3718), .b(N4304), .c(N3642), .O(N4377) );
and2 gate1305( .a(N330), .b(N4317), .O(N4387) );
and2 gate1306( .a(N330), .b(N4318), .O(N4390) );
nand2 gate1307( .a(N3921), .b(N4330), .O(N4393) );
buf1 gate1308( .a(N4287), .O(N4398) );
buf1 gate1309( .a(N4284), .O(N4413) );
nand3 gate1310( .a(N3920), .b(N4325), .c(N4326), .O(N4416) );
or2 gate1311( .a(N3812), .b(N4322), .O(N4421) );
nand3 gate1312( .a(N3948), .b(N4327), .c(N4328), .O(N4427) );
buf1 gate1313( .a(N4287), .O(N4430) );
and2 gate1314( .a(N330), .b(N4316), .O(N4435) );
or2 gate1315( .a(N4331), .b(N4296), .O(N4442) );
and4 gate1316( .a(N4174), .b(N4305), .c(N4203), .d(N4213), .O(N4443) );

  xor2  gate3070(.a(N3809), .b(N4305), .O(gate1317inter0));
  nand2 gate3071(.a(gate1317inter0), .b(s_200), .O(gate1317inter1));
  and2  gate3072(.a(N3809), .b(N4305), .O(gate1317inter2));
  inv1  gate3073(.a(s_200), .O(gate1317inter3));
  inv1  gate3074(.a(s_201), .O(gate1317inter4));
  nand2 gate3075(.a(gate1317inter4), .b(gate1317inter3), .O(gate1317inter5));
  nor2  gate3076(.a(gate1317inter5), .b(gate1317inter2), .O(gate1317inter6));
  inv1  gate3077(.a(N4305), .O(gate1317inter7));
  inv1  gate3078(.a(N3809), .O(gate1317inter8));
  nand2 gate3079(.a(gate1317inter8), .b(gate1317inter7), .O(gate1317inter9));
  nand2 gate3080(.a(s_201), .b(gate1317inter3), .O(gate1317inter10));
  nor2  gate3081(.a(gate1317inter10), .b(gate1317inter9), .O(gate1317inter11));
  nor2  gate3082(.a(gate1317inter11), .b(gate1317inter6), .O(gate1317inter12));
  nand2 gate3083(.a(gate1317inter12), .b(gate1317inter1), .O(N4446));
nand3 gate1318( .a(N4305), .b(N4200), .c(N3913), .O(N4447) );
nand4 gate1319( .a(N4305), .b(N4200), .c(N4213), .d(N4167), .O(N4448) );
inv1 gate1320( .a(N4356), .O(N4452) );

  xor2  gate3434(.a(N4393), .b(N4329), .O(gate1321inter0));
  nand2 gate3435(.a(gate1321inter0), .b(s_252), .O(gate1321inter1));
  and2  gate3436(.a(N4393), .b(N4329), .O(gate1321inter2));
  inv1  gate3437(.a(s_252), .O(gate1321inter3));
  inv1  gate3438(.a(s_253), .O(gate1321inter4));
  nand2 gate3439(.a(gate1321inter4), .b(gate1321inter3), .O(gate1321inter5));
  nor2  gate3440(.a(gate1321inter5), .b(gate1321inter2), .O(gate1321inter6));
  inv1  gate3441(.a(N4329), .O(gate1321inter7));
  inv1  gate3442(.a(N4393), .O(gate1321inter8));
  nand2 gate3443(.a(gate1321inter8), .b(gate1321inter7), .O(gate1321inter9));
  nand2 gate3444(.a(s_253), .b(gate1321inter3), .O(gate1321inter10));
  nor2  gate3445(.a(gate1321inter10), .b(gate1321inter9), .O(gate1321inter11));
  nor2  gate3446(.a(gate1321inter11), .b(gate1321inter6), .O(gate1321inter12));
  nand2 gate3447(.a(gate1321inter12), .b(gate1321inter1), .O(N4458));
inv1 gate1322( .a(N4365), .O(N4461) );
inv1 gate1323( .a(N4368), .O(N4462) );

  xor2  gate3196(.a(N1460), .b(N4371), .O(gate1324inter0));
  nand2 gate3197(.a(gate1324inter0), .b(s_218), .O(gate1324inter1));
  and2  gate3198(.a(N1460), .b(N4371), .O(gate1324inter2));
  inv1  gate3199(.a(s_218), .O(gate1324inter3));
  inv1  gate3200(.a(s_219), .O(gate1324inter4));
  nand2 gate3201(.a(gate1324inter4), .b(gate1324inter3), .O(gate1324inter5));
  nor2  gate3202(.a(gate1324inter5), .b(gate1324inter2), .O(gate1324inter6));
  inv1  gate3203(.a(N4371), .O(gate1324inter7));
  inv1  gate3204(.a(N1460), .O(gate1324inter8));
  nand2 gate3205(.a(gate1324inter8), .b(gate1324inter7), .O(gate1324inter9));
  nand2 gate3206(.a(s_219), .b(gate1324inter3), .O(gate1324inter10));
  nor2  gate3207(.a(gate1324inter10), .b(gate1324inter9), .O(gate1324inter11));
  nor2  gate3208(.a(gate1324inter11), .b(gate1324inter6), .O(gate1324inter12));
  nand2 gate3209(.a(gate1324inter12), .b(gate1324inter1), .O(N4463));
inv1 gate1325( .a(N4371), .O(N4464) );
buf1 gate1326( .a(N4310), .O(N4465) );
nor2 gate1327( .a(N4331), .b(N4296), .O(N4468) );
and2 gate1328( .a(N4376), .b(N2732), .O(N4472) );
and2 gate1329( .a(N4377), .b(N2740), .O(N4475) );
buf1 gate1330( .a(N4310), .O(N4479) );
inv1 gate1331( .a(N4353), .O(N4484) );
inv1 gate1332( .a(N4359), .O(N4486) );

  xor2  gate3770(.a(N4299), .b(N4359), .O(gate1333inter0));
  nand2 gate3771(.a(gate1333inter0), .b(s_300), .O(gate1333inter1));
  and2  gate3772(.a(N4299), .b(N4359), .O(gate1333inter2));
  inv1  gate3773(.a(s_300), .O(gate1333inter3));
  inv1  gate3774(.a(s_301), .O(gate1333inter4));
  nand2 gate3775(.a(gate1333inter4), .b(gate1333inter3), .O(gate1333inter5));
  nor2  gate3776(.a(gate1333inter5), .b(gate1333inter2), .O(gate1333inter6));
  inv1  gate3777(.a(N4359), .O(gate1333inter7));
  inv1  gate3778(.a(N4299), .O(gate1333inter8));
  nand2 gate3779(.a(gate1333inter8), .b(gate1333inter7), .O(gate1333inter9));
  nand2 gate3780(.a(s_301), .b(gate1333inter3), .O(gate1333inter10));
  nor2  gate3781(.a(gate1333inter10), .b(gate1333inter9), .O(gate1333inter11));
  nor2  gate3782(.a(gate1333inter11), .b(gate1333inter6), .O(gate1333inter12));
  nand2 gate3783(.a(gate1333inter12), .b(gate1333inter1), .O(N4487));
inv1 gate1334( .a(N4362), .O(N4491) );
and2 gate1335( .a(N330), .b(N4319), .O(N4493) );
inv1 gate1336( .a(N4398), .O(N4496) );
and2 gate1337( .a(N4287), .b(N4398), .O(N4497) );
and2 gate1338( .a(N4442), .b(N1769), .O(N4498) );
nand4 gate1339( .a(N3947), .b(N4446), .c(N4447), .d(N4448), .O(N4503) );
inv1 gate1340( .a(N4413), .O(N4506) );
inv1 gate1341( .a(N4435), .O(N4507) );
inv1 gate1342( .a(N4421), .O(N4508) );

  xor2  gate2020(.a(N4452), .b(N4421), .O(gate1343inter0));
  nand2 gate2021(.a(gate1343inter0), .b(s_50), .O(gate1343inter1));
  and2  gate2022(.a(N4452), .b(N4421), .O(gate1343inter2));
  inv1  gate2023(.a(s_50), .O(gate1343inter3));
  inv1  gate2024(.a(s_51), .O(gate1343inter4));
  nand2 gate2025(.a(gate1343inter4), .b(gate1343inter3), .O(gate1343inter5));
  nor2  gate2026(.a(gate1343inter5), .b(gate1343inter2), .O(gate1343inter6));
  inv1  gate2027(.a(N4421), .O(gate1343inter7));
  inv1  gate2028(.a(N4452), .O(gate1343inter8));
  nand2 gate2029(.a(gate1343inter8), .b(gate1343inter7), .O(gate1343inter9));
  nand2 gate2030(.a(s_51), .b(gate1343inter3), .O(gate1343inter10));
  nor2  gate2031(.a(gate1343inter10), .b(gate1343inter9), .O(gate1343inter11));
  nor2  gate2032(.a(gate1343inter11), .b(gate1343inter6), .O(gate1343inter12));
  nand2 gate2033(.a(gate1343inter12), .b(gate1343inter1), .O(N4509));
inv1 gate1344( .a(N4427), .O(N4510) );
nand2 gate1345( .a(N4427), .b(N4241), .O(N4511) );
nand2 gate1346( .a(N965), .b(N4464), .O(N4515) );
inv1 gate1347( .a(N4416), .O(N4526) );
nand2 gate1348( .a(N4416), .b(N4484), .O(N4527) );
nand2 gate1349( .a(N4182), .b(N4486), .O(N4528) );
inv1 gate1350( .a(N4430), .O(N4529) );

  xor2  gate1852(.a(N4491), .b(N4430), .O(gate1351inter0));
  nand2 gate1853(.a(gate1351inter0), .b(s_26), .O(gate1351inter1));
  and2  gate1854(.a(N4491), .b(N4430), .O(gate1351inter2));
  inv1  gate1855(.a(s_26), .O(gate1351inter3));
  inv1  gate1856(.a(s_27), .O(gate1351inter4));
  nand2 gate1857(.a(gate1351inter4), .b(gate1351inter3), .O(gate1351inter5));
  nor2  gate1858(.a(gate1351inter5), .b(gate1351inter2), .O(gate1351inter6));
  inv1  gate1859(.a(N4430), .O(gate1351inter7));
  inv1  gate1860(.a(N4491), .O(gate1351inter8));
  nand2 gate1861(.a(gate1351inter8), .b(gate1351inter7), .O(gate1351inter9));
  nand2 gate1862(.a(s_27), .b(gate1351inter3), .O(gate1351inter10));
  nor2  gate1863(.a(gate1351inter10), .b(gate1351inter9), .O(gate1351inter11));
  nor2  gate1864(.a(gate1351inter11), .b(gate1351inter6), .O(gate1351inter12));
  nand2 gate1865(.a(gate1351inter12), .b(gate1351inter1), .O(N4530));
buf1 gate1352( .a(N4387), .O(N4531) );
buf1 gate1353( .a(N4387), .O(N4534) );
buf1 gate1354( .a(N4390), .O(N4537) );
buf1 gate1355( .a(N4390), .O(N4540) );
and3 gate1356( .a(N330), .b(N4319), .c(N4496), .O(N4545) );
and2 gate1357( .a(N330), .b(N4443), .O(N4549) );
nand2 gate1358( .a(N4356), .b(N4508), .O(N4552) );

  xor2  gate2748(.a(N4510), .b(N4142), .O(gate1359inter0));
  nand2 gate2749(.a(gate1359inter0), .b(s_154), .O(gate1359inter1));
  and2  gate2750(.a(N4510), .b(N4142), .O(gate1359inter2));
  inv1  gate2751(.a(s_154), .O(gate1359inter3));
  inv1  gate2752(.a(s_155), .O(gate1359inter4));
  nand2 gate2753(.a(gate1359inter4), .b(gate1359inter3), .O(gate1359inter5));
  nor2  gate2754(.a(gate1359inter5), .b(gate1359inter2), .O(gate1359inter6));
  inv1  gate2755(.a(N4142), .O(gate1359inter7));
  inv1  gate2756(.a(N4510), .O(gate1359inter8));
  nand2 gate2757(.a(gate1359inter8), .b(gate1359inter7), .O(gate1359inter9));
  nand2 gate2758(.a(s_155), .b(gate1359inter3), .O(gate1359inter10));
  nor2  gate2759(.a(gate1359inter10), .b(gate1359inter9), .O(gate1359inter11));
  nor2  gate2760(.a(gate1359inter11), .b(gate1359inter6), .O(gate1359inter12));
  nand2 gate2761(.a(gate1359inter12), .b(gate1359inter1), .O(N4555));
inv1 gate1360( .a(N4493), .O(N4558) );

  xor2  gate2762(.a(N4515), .b(N4463), .O(gate1361inter0));
  nand2 gate2763(.a(gate1361inter0), .b(s_156), .O(gate1361inter1));
  and2  gate2764(.a(N4515), .b(N4463), .O(gate1361inter2));
  inv1  gate2765(.a(s_156), .O(gate1361inter3));
  inv1  gate2766(.a(s_157), .O(gate1361inter4));
  nand2 gate2767(.a(gate1361inter4), .b(gate1361inter3), .O(gate1361inter5));
  nor2  gate2768(.a(gate1361inter5), .b(gate1361inter2), .O(gate1361inter6));
  inv1  gate2769(.a(N4463), .O(gate1361inter7));
  inv1  gate2770(.a(N4515), .O(gate1361inter8));
  nand2 gate2771(.a(gate1361inter8), .b(gate1361inter7), .O(gate1361inter9));
  nand2 gate2772(.a(s_157), .b(gate1361inter3), .O(gate1361inter10));
  nor2  gate2773(.a(gate1361inter10), .b(gate1361inter9), .O(gate1361inter11));
  nor2  gate2774(.a(gate1361inter11), .b(gate1361inter6), .O(gate1361inter12));
  nand2 gate2775(.a(gate1361inter12), .b(gate1361inter1), .O(N4559));
inv1 gate1362( .a(N4465), .O(N4562) );
and2 gate1363( .a(N4310), .b(N4465), .O(N4563) );
buf1 gate1364( .a(N4468), .O(N4564) );
inv1 gate1365( .a(N4479), .O(N4568) );
buf1 gate1366( .a(N4443), .O(N4569) );
nand2 gate1367( .a(N4353), .b(N4526), .O(N4572) );

  xor2  gate1866(.a(N4529), .b(N4362), .O(gate1368inter0));
  nand2 gate1867(.a(gate1368inter0), .b(s_28), .O(gate1368inter1));
  and2  gate1868(.a(N4529), .b(N4362), .O(gate1368inter2));
  inv1  gate1869(.a(s_28), .O(gate1368inter3));
  inv1  gate1870(.a(s_29), .O(gate1368inter4));
  nand2 gate1871(.a(gate1368inter4), .b(gate1368inter3), .O(gate1368inter5));
  nor2  gate1872(.a(gate1368inter5), .b(gate1368inter2), .O(gate1368inter6));
  inv1  gate1873(.a(N4362), .O(gate1368inter7));
  inv1  gate1874(.a(N4529), .O(gate1368inter8));
  nand2 gate1875(.a(gate1368inter8), .b(gate1368inter7), .O(gate1368inter9));
  nand2 gate1876(.a(s_29), .b(gate1368inter3), .O(gate1368inter10));
  nor2  gate1877(.a(gate1368inter10), .b(gate1368inter9), .O(gate1368inter11));
  nor2  gate1878(.a(gate1368inter11), .b(gate1368inter6), .O(gate1368inter12));
  nand2 gate1879(.a(gate1368inter12), .b(gate1368inter1), .O(N4573));

  xor2  gate2062(.a(N4528), .b(N4487), .O(gate1369inter0));
  nand2 gate2063(.a(gate1369inter0), .b(s_56), .O(gate1369inter1));
  and2  gate2064(.a(N4528), .b(N4487), .O(gate1369inter2));
  inv1  gate2065(.a(s_56), .O(gate1369inter3));
  inv1  gate2066(.a(s_57), .O(gate1369inter4));
  nand2 gate2067(.a(gate1369inter4), .b(gate1369inter3), .O(gate1369inter5));
  nor2  gate2068(.a(gate1369inter5), .b(gate1369inter2), .O(gate1369inter6));
  inv1  gate2069(.a(N4487), .O(gate1369inter7));
  inv1  gate2070(.a(N4528), .O(gate1369inter8));
  nand2 gate2071(.a(gate1369inter8), .b(gate1369inter7), .O(gate1369inter9));
  nand2 gate2072(.a(s_57), .b(gate1369inter3), .O(gate1369inter10));
  nor2  gate2073(.a(gate1369inter10), .b(gate1369inter9), .O(gate1369inter11));
  nor2  gate2074(.a(gate1369inter11), .b(gate1369inter6), .O(gate1369inter12));
  nand2 gate2075(.a(gate1369inter12), .b(gate1369inter1), .O(N4576));
buf1 gate1370( .a(N4458), .O(N4581) );
buf1 gate1371( .a(N4458), .O(N4584) );
or3 gate1372( .a(N2758), .b(N4498), .c(N2761), .O(N4587) );
nor3 gate1373( .a(N2758), .b(N4498), .c(N2761), .O(N4588) );
or2 gate1374( .a(N4545), .b(N4497), .O(N4589) );

  xor2  gate1698(.a(N4509), .b(N4552), .O(gate1375inter0));
  nand2 gate1699(.a(gate1375inter0), .b(s_4), .O(gate1375inter1));
  and2  gate1700(.a(N4509), .b(N4552), .O(gate1375inter2));
  inv1  gate1701(.a(s_4), .O(gate1375inter3));
  inv1  gate1702(.a(s_5), .O(gate1375inter4));
  nand2 gate1703(.a(gate1375inter4), .b(gate1375inter3), .O(gate1375inter5));
  nor2  gate1704(.a(gate1375inter5), .b(gate1375inter2), .O(gate1375inter6));
  inv1  gate1705(.a(N4552), .O(gate1375inter7));
  inv1  gate1706(.a(N4509), .O(gate1375inter8));
  nand2 gate1707(.a(gate1375inter8), .b(gate1375inter7), .O(gate1375inter9));
  nand2 gate1708(.a(s_5), .b(gate1375inter3), .O(gate1375inter10));
  nor2  gate1709(.a(gate1375inter10), .b(gate1375inter9), .O(gate1375inter11));
  nor2  gate1710(.a(gate1375inter11), .b(gate1375inter6), .O(gate1375inter12));
  nand2 gate1711(.a(gate1375inter12), .b(gate1375inter1), .O(N4593));
inv1 gate1376( .a(N4531), .O(N4596) );
inv1 gate1377( .a(N4534), .O(N4597) );

  xor2  gate3126(.a(N4511), .b(N4555), .O(gate1378inter0));
  nand2 gate3127(.a(gate1378inter0), .b(s_208), .O(gate1378inter1));
  and2  gate3128(.a(N4511), .b(N4555), .O(gate1378inter2));
  inv1  gate3129(.a(s_208), .O(gate1378inter3));
  inv1  gate3130(.a(s_209), .O(gate1378inter4));
  nand2 gate3131(.a(gate1378inter4), .b(gate1378inter3), .O(gate1378inter5));
  nor2  gate3132(.a(gate1378inter5), .b(gate1378inter2), .O(gate1378inter6));
  inv1  gate3133(.a(N4555), .O(gate1378inter7));
  inv1  gate3134(.a(N4511), .O(gate1378inter8));
  nand2 gate3135(.a(gate1378inter8), .b(gate1378inter7), .O(gate1378inter9));
  nand2 gate3136(.a(s_209), .b(gate1378inter3), .O(gate1378inter10));
  nor2  gate3137(.a(gate1378inter10), .b(gate1378inter9), .O(gate1378inter11));
  nor2  gate3138(.a(gate1378inter11), .b(gate1378inter6), .O(gate1378inter12));
  nand2 gate3139(.a(gate1378inter12), .b(gate1378inter1), .O(N4599));
inv1 gate1379( .a(N4537), .O(N4602) );
inv1 gate1380( .a(N4540), .O(N4603) );
and3 gate1381( .a(N330), .b(N4284), .c(N4562), .O(N4608) );
buf1 gate1382( .a(N4503), .O(N4613) );
buf1 gate1383( .a(N4503), .O(N4616) );

  xor2  gate2370(.a(N4527), .b(N4572), .O(gate1384inter0));
  nand2 gate2371(.a(gate1384inter0), .b(s_100), .O(gate1384inter1));
  and2  gate2372(.a(N4527), .b(N4572), .O(gate1384inter2));
  inv1  gate2373(.a(s_100), .O(gate1384inter3));
  inv1  gate2374(.a(s_101), .O(gate1384inter4));
  nand2 gate2375(.a(gate1384inter4), .b(gate1384inter3), .O(gate1384inter5));
  nor2  gate2376(.a(gate1384inter5), .b(gate1384inter2), .O(gate1384inter6));
  inv1  gate2377(.a(N4572), .O(gate1384inter7));
  inv1  gate2378(.a(N4527), .O(gate1384inter8));
  nand2 gate2379(.a(gate1384inter8), .b(gate1384inter7), .O(gate1384inter9));
  nand2 gate2380(.a(s_101), .b(gate1384inter3), .O(gate1384inter10));
  nor2  gate2381(.a(gate1384inter10), .b(gate1384inter9), .O(gate1384inter11));
  nor2  gate2382(.a(gate1384inter11), .b(gate1384inter6), .O(gate1384inter12));
  nand2 gate2383(.a(gate1384inter12), .b(gate1384inter1), .O(N4619));
nand2 gate1385( .a(N4573), .b(N4530), .O(N4623) );
inv1 gate1386( .a(N4588), .O(N4628) );
nand2 gate1387( .a(N4569), .b(N4506), .O(N4629) );
inv1 gate1388( .a(N4569), .O(N4630) );
inv1 gate1389( .a(N4576), .O(N4635) );

  xor2  gate3672(.a(N4291), .b(N4576), .O(gate1390inter0));
  nand2 gate3673(.a(gate1390inter0), .b(s_286), .O(gate1390inter1));
  and2  gate3674(.a(N4291), .b(N4576), .O(gate1390inter2));
  inv1  gate3675(.a(s_286), .O(gate1390inter3));
  inv1  gate3676(.a(s_287), .O(gate1390inter4));
  nand2 gate3677(.a(gate1390inter4), .b(gate1390inter3), .O(gate1390inter5));
  nor2  gate3678(.a(gate1390inter5), .b(gate1390inter2), .O(gate1390inter6));
  inv1  gate3679(.a(N4576), .O(gate1390inter7));
  inv1  gate3680(.a(N4291), .O(gate1390inter8));
  nand2 gate3681(.a(gate1390inter8), .b(gate1390inter7), .O(gate1390inter9));
  nand2 gate3682(.a(s_287), .b(gate1390inter3), .O(gate1390inter10));
  nor2  gate3683(.a(gate1390inter10), .b(gate1390inter9), .O(gate1390inter11));
  nor2  gate3684(.a(gate1390inter11), .b(gate1390inter6), .O(gate1390inter12));
  nand2 gate3685(.a(gate1390inter12), .b(gate1390inter1), .O(N4636));
inv1 gate1391( .a(N4581), .O(N4640) );

  xor2  gate3658(.a(N4461), .b(N4581), .O(gate1392inter0));
  nand2 gate3659(.a(gate1392inter0), .b(s_284), .O(gate1392inter1));
  and2  gate3660(.a(N4461), .b(N4581), .O(gate1392inter2));
  inv1  gate3661(.a(s_284), .O(gate1392inter3));
  inv1  gate3662(.a(s_285), .O(gate1392inter4));
  nand2 gate3663(.a(gate1392inter4), .b(gate1392inter3), .O(gate1392inter5));
  nor2  gate3664(.a(gate1392inter5), .b(gate1392inter2), .O(gate1392inter6));
  inv1  gate3665(.a(N4581), .O(gate1392inter7));
  inv1  gate3666(.a(N4461), .O(gate1392inter8));
  nand2 gate3667(.a(gate1392inter8), .b(gate1392inter7), .O(gate1392inter9));
  nand2 gate3668(.a(s_285), .b(gate1392inter3), .O(gate1392inter10));
  nor2  gate3669(.a(gate1392inter10), .b(gate1392inter9), .O(gate1392inter11));
  nor2  gate3670(.a(gate1392inter11), .b(gate1392inter6), .O(gate1392inter12));
  nand2 gate3671(.a(gate1392inter12), .b(gate1392inter1), .O(N4641));
inv1 gate1393( .a(N4584), .O(N4642) );

  xor2  gate2034(.a(N4462), .b(N4584), .O(gate1394inter0));
  nand2 gate2035(.a(gate1394inter0), .b(s_52), .O(gate1394inter1));
  and2  gate2036(.a(N4462), .b(N4584), .O(gate1394inter2));
  inv1  gate2037(.a(s_52), .O(gate1394inter3));
  inv1  gate2038(.a(s_53), .O(gate1394inter4));
  nand2 gate2039(.a(gate1394inter4), .b(gate1394inter3), .O(gate1394inter5));
  nor2  gate2040(.a(gate1394inter5), .b(gate1394inter2), .O(gate1394inter6));
  inv1  gate2041(.a(N4584), .O(gate1394inter7));
  inv1  gate2042(.a(N4462), .O(gate1394inter8));
  nand2 gate2043(.a(gate1394inter8), .b(gate1394inter7), .O(gate1394inter9));
  nand2 gate2044(.a(s_53), .b(gate1394inter3), .O(gate1394inter10));
  nor2  gate2045(.a(gate1394inter10), .b(gate1394inter9), .O(gate1394inter11));
  nor2  gate2046(.a(gate1394inter11), .b(gate1394inter6), .O(gate1394inter12));
  nand2 gate2047(.a(gate1394inter12), .b(gate1394inter1), .O(N4643));

  xor2  gate3924(.a(N4563), .b(N4608), .O(gate1395inter0));
  nand2 gate3925(.a(gate1395inter0), .b(s_322), .O(gate1395inter1));
  and2  gate3926(.a(N4563), .b(N4608), .O(gate1395inter2));
  inv1  gate3927(.a(s_322), .O(gate1395inter3));
  inv1  gate3928(.a(s_323), .O(gate1395inter4));
  nand2 gate3929(.a(gate1395inter4), .b(gate1395inter3), .O(gate1395inter5));
  nor2  gate3930(.a(gate1395inter5), .b(gate1395inter2), .O(gate1395inter6));
  inv1  gate3931(.a(N4608), .O(gate1395inter7));
  inv1  gate3932(.a(N4563), .O(gate1395inter8));
  nand2 gate3933(.a(gate1395inter8), .b(gate1395inter7), .O(gate1395inter9));
  nand2 gate3934(.a(s_323), .b(gate1395inter3), .O(gate1395inter10));
  nor2  gate3935(.a(gate1395inter10), .b(gate1395inter9), .O(gate1395inter11));
  nor2  gate3936(.a(gate1395inter11), .b(gate1395inter6), .O(gate1395inter12));
  nand2 gate3937(.a(gate1395inter12), .b(gate1395inter1), .O(N4644));
and2 gate1396( .a(N4559), .b(N2128), .O(N4647) );
and2 gate1397( .a(N4559), .b(N2743), .O(N4650) );
buf1 gate1398( .a(N4549), .O(N4656) );
buf1 gate1399( .a(N4549), .O(N4659) );
buf1 gate1400( .a(N4564), .O(N4664) );
and2 gate1401( .a(N4587), .b(N4628), .O(N4667) );
nand2 gate1402( .a(N4413), .b(N4630), .O(N4668) );
inv1 gate1403( .a(N4616), .O(N4669) );
nand2 gate1404( .a(N4616), .b(N4239), .O(N4670) );
inv1 gate1405( .a(N4619), .O(N4673) );
nand2 gate1406( .a(N4619), .b(N4507), .O(N4674) );

  xor2  gate3728(.a(N4635), .b(N4186), .O(gate1407inter0));
  nand2 gate3729(.a(gate1407inter0), .b(s_294), .O(gate1407inter1));
  and2  gate3730(.a(N4635), .b(N4186), .O(gate1407inter2));
  inv1  gate3731(.a(s_294), .O(gate1407inter3));
  inv1  gate3732(.a(s_295), .O(gate1407inter4));
  nand2 gate3733(.a(gate1407inter4), .b(gate1407inter3), .O(gate1407inter5));
  nor2  gate3734(.a(gate1407inter5), .b(gate1407inter2), .O(gate1407inter6));
  inv1  gate3735(.a(N4186), .O(gate1407inter7));
  inv1  gate3736(.a(N4635), .O(gate1407inter8));
  nand2 gate3737(.a(gate1407inter8), .b(gate1407inter7), .O(gate1407inter9));
  nand2 gate3738(.a(s_295), .b(gate1407inter3), .O(gate1407inter10));
  nor2  gate3739(.a(gate1407inter10), .b(gate1407inter9), .O(gate1407inter11));
  nor2  gate3740(.a(gate1407inter11), .b(gate1407inter6), .O(gate1407inter12));
  nand2 gate3741(.a(gate1407inter12), .b(gate1407inter1), .O(N4675));
inv1 gate1408( .a(N4623), .O(N4676) );

  xor2  gate4260(.a(N4558), .b(N4623), .O(gate1409inter0));
  nand2 gate4261(.a(gate1409inter0), .b(s_370), .O(gate1409inter1));
  and2  gate4262(.a(N4558), .b(N4623), .O(gate1409inter2));
  inv1  gate4263(.a(s_370), .O(gate1409inter3));
  inv1  gate4264(.a(s_371), .O(gate1409inter4));
  nand2 gate4265(.a(gate1409inter4), .b(gate1409inter3), .O(gate1409inter5));
  nor2  gate4266(.a(gate1409inter5), .b(gate1409inter2), .O(gate1409inter6));
  inv1  gate4267(.a(N4623), .O(gate1409inter7));
  inv1  gate4268(.a(N4558), .O(gate1409inter8));
  nand2 gate4269(.a(gate1409inter8), .b(gate1409inter7), .O(gate1409inter9));
  nand2 gate4270(.a(s_371), .b(gate1409inter3), .O(gate1409inter10));
  nor2  gate4271(.a(gate1409inter10), .b(gate1409inter9), .O(gate1409inter11));
  nor2  gate4272(.a(gate1409inter11), .b(gate1409inter6), .O(gate1409inter12));
  nand2 gate4273(.a(gate1409inter12), .b(gate1409inter1), .O(N4677));
nand2 gate1410( .a(N4365), .b(N4640), .O(N4678) );

  xor2  gate3028(.a(N4642), .b(N4368), .O(gate1411inter0));
  nand2 gate3029(.a(gate1411inter0), .b(s_194), .O(gate1411inter1));
  and2  gate3030(.a(N4642), .b(N4368), .O(gate1411inter2));
  inv1  gate3031(.a(s_194), .O(gate1411inter3));
  inv1  gate3032(.a(s_195), .O(gate1411inter4));
  nand2 gate3033(.a(gate1411inter4), .b(gate1411inter3), .O(gate1411inter5));
  nor2  gate3034(.a(gate1411inter5), .b(gate1411inter2), .O(gate1411inter6));
  inv1  gate3035(.a(N4368), .O(gate1411inter7));
  inv1  gate3036(.a(N4642), .O(gate1411inter8));
  nand2 gate3037(.a(gate1411inter8), .b(gate1411inter7), .O(gate1411inter9));
  nand2 gate3038(.a(s_195), .b(gate1411inter3), .O(gate1411inter10));
  nor2  gate3039(.a(gate1411inter10), .b(gate1411inter9), .O(gate1411inter11));
  nor2  gate3040(.a(gate1411inter11), .b(gate1411inter6), .O(gate1411inter12));
  nand2 gate3041(.a(gate1411inter12), .b(gate1411inter1), .O(N4679));
inv1 gate1412( .a(N4613), .O(N4687) );
nand2 gate1413( .a(N4613), .b(N4568), .O(N4688) );
buf1 gate1414( .a(N4593), .O(N4691) );
buf1 gate1415( .a(N4593), .O(N4694) );
buf1 gate1416( .a(N4599), .O(N4697) );
buf1 gate1417( .a(N4599), .O(N4700) );

  xor2  gate3098(.a(N4668), .b(N4629), .O(gate1418inter0));
  nand2 gate3099(.a(gate1418inter0), .b(s_204), .O(gate1418inter1));
  and2  gate3100(.a(N4668), .b(N4629), .O(gate1418inter2));
  inv1  gate3101(.a(s_204), .O(gate1418inter3));
  inv1  gate3102(.a(s_205), .O(gate1418inter4));
  nand2 gate3103(.a(gate1418inter4), .b(gate1418inter3), .O(gate1418inter5));
  nor2  gate3104(.a(gate1418inter5), .b(gate1418inter2), .O(gate1418inter6));
  inv1  gate3105(.a(N4629), .O(gate1418inter7));
  inv1  gate3106(.a(N4668), .O(gate1418inter8));
  nand2 gate3107(.a(gate1418inter8), .b(gate1418inter7), .O(gate1418inter9));
  nand2 gate3108(.a(s_205), .b(gate1418inter3), .O(gate1418inter10));
  nor2  gate3109(.a(gate1418inter10), .b(gate1418inter9), .O(gate1418inter11));
  nor2  gate3110(.a(gate1418inter11), .b(gate1418inter6), .O(gate1418inter12));
  nand2 gate3111(.a(gate1418inter12), .b(gate1418inter1), .O(N4704));

  xor2  gate3966(.a(N4669), .b(N4139), .O(gate1419inter0));
  nand2 gate3967(.a(gate1419inter0), .b(s_328), .O(gate1419inter1));
  and2  gate3968(.a(N4669), .b(N4139), .O(gate1419inter2));
  inv1  gate3969(.a(s_328), .O(gate1419inter3));
  inv1  gate3970(.a(s_329), .O(gate1419inter4));
  nand2 gate3971(.a(gate1419inter4), .b(gate1419inter3), .O(gate1419inter5));
  nor2  gate3972(.a(gate1419inter5), .b(gate1419inter2), .O(gate1419inter6));
  inv1  gate3973(.a(N4139), .O(gate1419inter7));
  inv1  gate3974(.a(N4669), .O(gate1419inter8));
  nand2 gate3975(.a(gate1419inter8), .b(gate1419inter7), .O(gate1419inter9));
  nand2 gate3976(.a(s_329), .b(gate1419inter3), .O(gate1419inter10));
  nor2  gate3977(.a(gate1419inter10), .b(gate1419inter9), .O(gate1419inter11));
  nor2  gate3978(.a(gate1419inter11), .b(gate1419inter6), .O(gate1419inter12));
  nand2 gate3979(.a(gate1419inter12), .b(gate1419inter1), .O(N4705));
inv1 gate1420( .a(N4656), .O(N4706) );
inv1 gate1421( .a(N4659), .O(N4707) );
nand2 gate1422( .a(N4435), .b(N4673), .O(N4708) );

  xor2  gate1796(.a(N4636), .b(N4675), .O(gate1423inter0));
  nand2 gate1797(.a(gate1423inter0), .b(s_18), .O(gate1423inter1));
  and2  gate1798(.a(N4636), .b(N4675), .O(gate1423inter2));
  inv1  gate1799(.a(s_18), .O(gate1423inter3));
  inv1  gate1800(.a(s_19), .O(gate1423inter4));
  nand2 gate1801(.a(gate1423inter4), .b(gate1423inter3), .O(gate1423inter5));
  nor2  gate1802(.a(gate1423inter5), .b(gate1423inter2), .O(gate1423inter6));
  inv1  gate1803(.a(N4675), .O(gate1423inter7));
  inv1  gate1804(.a(N4636), .O(gate1423inter8));
  nand2 gate1805(.a(gate1423inter8), .b(gate1423inter7), .O(gate1423inter9));
  nand2 gate1806(.a(s_19), .b(gate1423inter3), .O(gate1423inter10));
  nor2  gate1807(.a(gate1423inter10), .b(gate1423inter9), .O(gate1423inter11));
  nor2  gate1808(.a(gate1423inter11), .b(gate1423inter6), .O(gate1423inter12));
  nand2 gate1809(.a(gate1423inter12), .b(gate1423inter1), .O(N4711));
nand2 gate1424( .a(N4493), .b(N4676), .O(N4716) );

  xor2  gate3756(.a(N4641), .b(N4678), .O(gate1425inter0));
  nand2 gate3757(.a(gate1425inter0), .b(s_298), .O(gate1425inter1));
  and2  gate3758(.a(N4641), .b(N4678), .O(gate1425inter2));
  inv1  gate3759(.a(s_298), .O(gate1425inter3));
  inv1  gate3760(.a(s_299), .O(gate1425inter4));
  nand2 gate3761(.a(gate1425inter4), .b(gate1425inter3), .O(gate1425inter5));
  nor2  gate3762(.a(gate1425inter5), .b(gate1425inter2), .O(gate1425inter6));
  inv1  gate3763(.a(N4678), .O(gate1425inter7));
  inv1  gate3764(.a(N4641), .O(gate1425inter8));
  nand2 gate3765(.a(gate1425inter8), .b(gate1425inter7), .O(gate1425inter9));
  nand2 gate3766(.a(s_299), .b(gate1425inter3), .O(gate1425inter10));
  nor2  gate3767(.a(gate1425inter10), .b(gate1425inter9), .O(gate1425inter11));
  nor2  gate3768(.a(gate1425inter11), .b(gate1425inter6), .O(gate1425inter12));
  nand2 gate3769(.a(gate1425inter12), .b(gate1425inter1), .O(N4717));

  xor2  gate3448(.a(N4643), .b(N4679), .O(gate1426inter0));
  nand2 gate3449(.a(gate1426inter0), .b(s_254), .O(gate1426inter1));
  and2  gate3450(.a(N4643), .b(N4679), .O(gate1426inter2));
  inv1  gate3451(.a(s_254), .O(gate1426inter3));
  inv1  gate3452(.a(s_255), .O(gate1426inter4));
  nand2 gate3453(.a(gate1426inter4), .b(gate1426inter3), .O(gate1426inter5));
  nor2  gate3454(.a(gate1426inter5), .b(gate1426inter2), .O(gate1426inter6));
  inv1  gate3455(.a(N4679), .O(gate1426inter7));
  inv1  gate3456(.a(N4643), .O(gate1426inter8));
  nand2 gate3457(.a(gate1426inter8), .b(gate1426inter7), .O(gate1426inter9));
  nand2 gate3458(.a(s_255), .b(gate1426inter3), .O(gate1426inter10));
  nor2  gate3459(.a(gate1426inter10), .b(gate1426inter9), .O(gate1426inter11));
  nor2  gate3460(.a(gate1426inter11), .b(gate1426inter6), .O(gate1426inter12));
  nand2 gate3461(.a(gate1426inter12), .b(gate1426inter1), .O(N4721));
buf1 gate1427( .a(N4644), .O(N4722) );
inv1 gate1428( .a(N4664), .O(N4726) );
or3 gate1429( .a(N4647), .b(N4650), .c(N4350), .O(N4727) );
nor3 gate1430( .a(N4647), .b(N4650), .c(N4350), .O(N4730) );
nand2 gate1431( .a(N4479), .b(N4687), .O(N4733) );
nand2 gate1432( .a(N4705), .b(N4670), .O(N4740) );

  xor2  gate3518(.a(N4674), .b(N4708), .O(gate1433inter0));
  nand2 gate3519(.a(gate1433inter0), .b(s_264), .O(gate1433inter1));
  and2  gate3520(.a(N4674), .b(N4708), .O(gate1433inter2));
  inv1  gate3521(.a(s_264), .O(gate1433inter3));
  inv1  gate3522(.a(s_265), .O(gate1433inter4));
  nand2 gate3523(.a(gate1433inter4), .b(gate1433inter3), .O(gate1433inter5));
  nor2  gate3524(.a(gate1433inter5), .b(gate1433inter2), .O(gate1433inter6));
  inv1  gate3525(.a(N4708), .O(gate1433inter7));
  inv1  gate3526(.a(N4674), .O(gate1433inter8));
  nand2 gate3527(.a(gate1433inter8), .b(gate1433inter7), .O(gate1433inter9));
  nand2 gate3528(.a(s_265), .b(gate1433inter3), .O(gate1433inter10));
  nor2  gate3529(.a(gate1433inter10), .b(gate1433inter9), .O(gate1433inter11));
  nor2  gate3530(.a(gate1433inter11), .b(gate1433inter6), .O(gate1433inter12));
  nand2 gate3531(.a(gate1433inter12), .b(gate1433inter1), .O(N4743));
inv1 gate1434( .a(N4691), .O(N4747) );

  xor2  gate3322(.a(N4596), .b(N4691), .O(gate1435inter0));
  nand2 gate3323(.a(gate1435inter0), .b(s_236), .O(gate1435inter1));
  and2  gate3324(.a(N4596), .b(N4691), .O(gate1435inter2));
  inv1  gate3325(.a(s_236), .O(gate1435inter3));
  inv1  gate3326(.a(s_237), .O(gate1435inter4));
  nand2 gate3327(.a(gate1435inter4), .b(gate1435inter3), .O(gate1435inter5));
  nor2  gate3328(.a(gate1435inter5), .b(gate1435inter2), .O(gate1435inter6));
  inv1  gate3329(.a(N4691), .O(gate1435inter7));
  inv1  gate3330(.a(N4596), .O(gate1435inter8));
  nand2 gate3331(.a(gate1435inter8), .b(gate1435inter7), .O(gate1435inter9));
  nand2 gate3332(.a(s_237), .b(gate1435inter3), .O(gate1435inter10));
  nor2  gate3333(.a(gate1435inter10), .b(gate1435inter9), .O(gate1435inter11));
  nor2  gate3334(.a(gate1435inter11), .b(gate1435inter6), .O(gate1435inter12));
  nand2 gate3335(.a(gate1435inter12), .b(gate1435inter1), .O(N4748));
inv1 gate1436( .a(N4694), .O(N4749) );

  xor2  gate3406(.a(N4597), .b(N4694), .O(gate1437inter0));
  nand2 gate3407(.a(gate1437inter0), .b(s_248), .O(gate1437inter1));
  and2  gate3408(.a(N4597), .b(N4694), .O(gate1437inter2));
  inv1  gate3409(.a(s_248), .O(gate1437inter3));
  inv1  gate3410(.a(s_249), .O(gate1437inter4));
  nand2 gate3411(.a(gate1437inter4), .b(gate1437inter3), .O(gate1437inter5));
  nor2  gate3412(.a(gate1437inter5), .b(gate1437inter2), .O(gate1437inter6));
  inv1  gate3413(.a(N4694), .O(gate1437inter7));
  inv1  gate3414(.a(N4597), .O(gate1437inter8));
  nand2 gate3415(.a(gate1437inter8), .b(gate1437inter7), .O(gate1437inter9));
  nand2 gate3416(.a(s_249), .b(gate1437inter3), .O(gate1437inter10));
  nor2  gate3417(.a(gate1437inter10), .b(gate1437inter9), .O(gate1437inter11));
  nor2  gate3418(.a(gate1437inter11), .b(gate1437inter6), .O(gate1437inter12));
  nand2 gate3419(.a(gate1437inter12), .b(gate1437inter1), .O(N4750));
inv1 gate1438( .a(N4697), .O(N4753) );
nand2 gate1439( .a(N4697), .b(N4602), .O(N4754) );
inv1 gate1440( .a(N4700), .O(N4755) );
nand2 gate1441( .a(N4700), .b(N4603), .O(N4756) );

  xor2  gate4008(.a(N4677), .b(N4716), .O(gate1442inter0));
  nand2 gate4009(.a(gate1442inter0), .b(s_334), .O(gate1442inter1));
  and2  gate4010(.a(N4677), .b(N4716), .O(gate1442inter2));
  inv1  gate4011(.a(s_334), .O(gate1442inter3));
  inv1  gate4012(.a(s_335), .O(gate1442inter4));
  nand2 gate4013(.a(gate1442inter4), .b(gate1442inter3), .O(gate1442inter5));
  nor2  gate4014(.a(gate1442inter5), .b(gate1442inter2), .O(gate1442inter6));
  inv1  gate4015(.a(N4716), .O(gate1442inter7));
  inv1  gate4016(.a(N4677), .O(gate1442inter8));
  nand2 gate4017(.a(gate1442inter8), .b(gate1442inter7), .O(gate1442inter9));
  nand2 gate4018(.a(s_335), .b(gate1442inter3), .O(gate1442inter10));
  nor2  gate4019(.a(gate1442inter10), .b(gate1442inter9), .O(gate1442inter11));
  nor2  gate4020(.a(gate1442inter11), .b(gate1442inter6), .O(gate1442inter12));
  nand2 gate4021(.a(gate1442inter12), .b(gate1442inter1), .O(N4757));
nand2 gate1443( .a(N4733), .b(N4688), .O(N4769) );
and2 gate1444( .a(N330), .b(N4704), .O(N4772) );
inv1 gate1445( .a(N4721), .O(N4775) );
inv1 gate1446( .a(N4730), .O(N4778) );

  xor2  gate2118(.a(N4747), .b(N4531), .O(gate1447inter0));
  nand2 gate2119(.a(gate1447inter0), .b(s_64), .O(gate1447inter1));
  and2  gate2120(.a(N4747), .b(N4531), .O(gate1447inter2));
  inv1  gate2121(.a(s_64), .O(gate1447inter3));
  inv1  gate2122(.a(s_65), .O(gate1447inter4));
  nand2 gate2123(.a(gate1447inter4), .b(gate1447inter3), .O(gate1447inter5));
  nor2  gate2124(.a(gate1447inter5), .b(gate1447inter2), .O(gate1447inter6));
  inv1  gate2125(.a(N4531), .O(gate1447inter7));
  inv1  gate2126(.a(N4747), .O(gate1447inter8));
  nand2 gate2127(.a(gate1447inter8), .b(gate1447inter7), .O(gate1447inter9));
  nand2 gate2128(.a(s_65), .b(gate1447inter3), .O(gate1447inter10));
  nor2  gate2129(.a(gate1447inter10), .b(gate1447inter9), .O(gate1447inter11));
  nor2  gate2130(.a(gate1447inter11), .b(gate1447inter6), .O(gate1447inter12));
  nand2 gate2131(.a(gate1447inter12), .b(gate1447inter1), .O(N4786));

  xor2  gate2678(.a(N4749), .b(N4534), .O(gate1448inter0));
  nand2 gate2679(.a(gate1448inter0), .b(s_144), .O(gate1448inter1));
  and2  gate2680(.a(N4749), .b(N4534), .O(gate1448inter2));
  inv1  gate2681(.a(s_144), .O(gate1448inter3));
  inv1  gate2682(.a(s_145), .O(gate1448inter4));
  nand2 gate2683(.a(gate1448inter4), .b(gate1448inter3), .O(gate1448inter5));
  nor2  gate2684(.a(gate1448inter5), .b(gate1448inter2), .O(gate1448inter6));
  inv1  gate2685(.a(N4534), .O(gate1448inter7));
  inv1  gate2686(.a(N4749), .O(gate1448inter8));
  nand2 gate2687(.a(gate1448inter8), .b(gate1448inter7), .O(gate1448inter9));
  nand2 gate2688(.a(s_145), .b(gate1448inter3), .O(gate1448inter10));
  nor2  gate2689(.a(gate1448inter10), .b(gate1448inter9), .O(gate1448inter11));
  nor2  gate2690(.a(gate1448inter11), .b(gate1448inter6), .O(gate1448inter12));
  nand2 gate2691(.a(gate1448inter12), .b(gate1448inter1), .O(N4787));

  xor2  gate2244(.a(N4753), .b(N4537), .O(gate1449inter0));
  nand2 gate2245(.a(gate1449inter0), .b(s_82), .O(gate1449inter1));
  and2  gate2246(.a(N4753), .b(N4537), .O(gate1449inter2));
  inv1  gate2247(.a(s_82), .O(gate1449inter3));
  inv1  gate2248(.a(s_83), .O(gate1449inter4));
  nand2 gate2249(.a(gate1449inter4), .b(gate1449inter3), .O(gate1449inter5));
  nor2  gate2250(.a(gate1449inter5), .b(gate1449inter2), .O(gate1449inter6));
  inv1  gate2251(.a(N4537), .O(gate1449inter7));
  inv1  gate2252(.a(N4753), .O(gate1449inter8));
  nand2 gate2253(.a(gate1449inter8), .b(gate1449inter7), .O(gate1449inter9));
  nand2 gate2254(.a(s_83), .b(gate1449inter3), .O(gate1449inter10));
  nor2  gate2255(.a(gate1449inter10), .b(gate1449inter9), .O(gate1449inter11));
  nor2  gate2256(.a(gate1449inter11), .b(gate1449inter6), .O(gate1449inter12));
  nand2 gate2257(.a(gate1449inter12), .b(gate1449inter1), .O(N4788));
nand2 gate1450( .a(N4540), .b(N4755), .O(N4789) );
and2 gate1451( .a(N4711), .b(N2124), .O(N4794) );
and2 gate1452( .a(N4711), .b(N2735), .O(N4797) );
and2 gate1453( .a(N4717), .b(N2127), .O(N4800) );
buf1 gate1454( .a(N4722), .O(N4805) );
and2 gate1455( .a(N4717), .b(N4468), .O(N4808) );
buf1 gate1456( .a(N4727), .O(N4812) );
and2 gate1457( .a(N4727), .b(N4778), .O(N4815) );
inv1 gate1458( .a(N4769), .O(N4816) );
inv1 gate1459( .a(N4772), .O(N4817) );
nand2 gate1460( .a(N4786), .b(N4748), .O(N4818) );

  xor2  gate4204(.a(N4750), .b(N4787), .O(gate1461inter0));
  nand2 gate4205(.a(gate1461inter0), .b(s_362), .O(gate1461inter1));
  and2  gate4206(.a(N4750), .b(N4787), .O(gate1461inter2));
  inv1  gate4207(.a(s_362), .O(gate1461inter3));
  inv1  gate4208(.a(s_363), .O(gate1461inter4));
  nand2 gate4209(.a(gate1461inter4), .b(gate1461inter3), .O(gate1461inter5));
  nor2  gate4210(.a(gate1461inter5), .b(gate1461inter2), .O(gate1461inter6));
  inv1  gate4211(.a(N4787), .O(gate1461inter7));
  inv1  gate4212(.a(N4750), .O(gate1461inter8));
  nand2 gate4213(.a(gate1461inter8), .b(gate1461inter7), .O(gate1461inter9));
  nand2 gate4214(.a(s_363), .b(gate1461inter3), .O(gate1461inter10));
  nor2  gate4215(.a(gate1461inter10), .b(gate1461inter9), .O(gate1461inter11));
  nor2  gate4216(.a(gate1461inter11), .b(gate1461inter6), .O(gate1461inter12));
  nand2 gate4217(.a(gate1461inter12), .b(gate1461inter1), .O(N4822));

  xor2  gate2328(.a(N4754), .b(N4788), .O(gate1462inter0));
  nand2 gate2329(.a(gate1462inter0), .b(s_94), .O(gate1462inter1));
  and2  gate2330(.a(N4754), .b(N4788), .O(gate1462inter2));
  inv1  gate2331(.a(s_94), .O(gate1462inter3));
  inv1  gate2332(.a(s_95), .O(gate1462inter4));
  nand2 gate2333(.a(gate1462inter4), .b(gate1462inter3), .O(gate1462inter5));
  nor2  gate2334(.a(gate1462inter5), .b(gate1462inter2), .O(gate1462inter6));
  inv1  gate2335(.a(N4788), .O(gate1462inter7));
  inv1  gate2336(.a(N4754), .O(gate1462inter8));
  nand2 gate2337(.a(gate1462inter8), .b(gate1462inter7), .O(gate1462inter9));
  nand2 gate2338(.a(s_95), .b(gate1462inter3), .O(gate1462inter10));
  nor2  gate2339(.a(gate1462inter10), .b(gate1462inter9), .O(gate1462inter11));
  nor2  gate2340(.a(gate1462inter11), .b(gate1462inter6), .O(gate1462inter12));
  nand2 gate2341(.a(gate1462inter12), .b(gate1462inter1), .O(N4823));
nand2 gate1463( .a(N4789), .b(N4756), .O(N4826) );

  xor2  gate3056(.a(N4726), .b(N4775), .O(gate1464inter0));
  nand2 gate3057(.a(gate1464inter0), .b(s_198), .O(gate1464inter1));
  and2  gate3058(.a(N4726), .b(N4775), .O(gate1464inter2));
  inv1  gate3059(.a(s_198), .O(gate1464inter3));
  inv1  gate3060(.a(s_199), .O(gate1464inter4));
  nand2 gate3061(.a(gate1464inter4), .b(gate1464inter3), .O(gate1464inter5));
  nor2  gate3062(.a(gate1464inter5), .b(gate1464inter2), .O(gate1464inter6));
  inv1  gate3063(.a(N4775), .O(gate1464inter7));
  inv1  gate3064(.a(N4726), .O(gate1464inter8));
  nand2 gate3065(.a(gate1464inter8), .b(gate1464inter7), .O(gate1464inter9));
  nand2 gate3066(.a(s_199), .b(gate1464inter3), .O(gate1464inter10));
  nor2  gate3067(.a(gate1464inter10), .b(gate1464inter9), .O(gate1464inter11));
  nor2  gate3068(.a(gate1464inter11), .b(gate1464inter6), .O(gate1464inter12));
  nand2 gate3069(.a(gate1464inter12), .b(gate1464inter1), .O(N4829));
inv1 gate1465( .a(N4775), .O(N4830) );
and2 gate1466( .a(N4743), .b(N2122), .O(N4831) );
and2 gate1467( .a(N4757), .b(N2126), .O(N4838) );
buf1 gate1468( .a(N4740), .O(N4844) );
buf1 gate1469( .a(N4740), .O(N4847) );
buf1 gate1470( .a(N4743), .O(N4850) );
buf1 gate1471( .a(N4757), .O(N4854) );

  xor2  gate3336(.a(N4816), .b(N4772), .O(gate1472inter0));
  nand2 gate3337(.a(gate1472inter0), .b(s_238), .O(gate1472inter1));
  and2  gate3338(.a(N4816), .b(N4772), .O(gate1472inter2));
  inv1  gate3339(.a(s_238), .O(gate1472inter3));
  inv1  gate3340(.a(s_239), .O(gate1472inter4));
  nand2 gate3341(.a(gate1472inter4), .b(gate1472inter3), .O(gate1472inter5));
  nor2  gate3342(.a(gate1472inter5), .b(gate1472inter2), .O(gate1472inter6));
  inv1  gate3343(.a(N4772), .O(gate1472inter7));
  inv1  gate3344(.a(N4816), .O(gate1472inter8));
  nand2 gate3345(.a(gate1472inter8), .b(gate1472inter7), .O(gate1472inter9));
  nand2 gate3346(.a(s_239), .b(gate1472inter3), .O(gate1472inter10));
  nor2  gate3347(.a(gate1472inter10), .b(gate1472inter9), .O(gate1472inter11));
  nor2  gate3348(.a(gate1472inter11), .b(gate1472inter6), .O(gate1472inter12));
  nand2 gate3349(.a(gate1472inter12), .b(gate1472inter1), .O(N4859));

  xor2  gate3532(.a(N4817), .b(N4769), .O(gate1473inter0));
  nand2 gate3533(.a(gate1473inter0), .b(s_266), .O(gate1473inter1));
  and2  gate3534(.a(N4817), .b(N4769), .O(gate1473inter2));
  inv1  gate3535(.a(s_266), .O(gate1473inter3));
  inv1  gate3536(.a(s_267), .O(gate1473inter4));
  nand2 gate3537(.a(gate1473inter4), .b(gate1473inter3), .O(gate1473inter5));
  nor2  gate3538(.a(gate1473inter5), .b(gate1473inter2), .O(gate1473inter6));
  inv1  gate3539(.a(N4769), .O(gate1473inter7));
  inv1  gate3540(.a(N4817), .O(gate1473inter8));
  nand2 gate3541(.a(gate1473inter8), .b(gate1473inter7), .O(gate1473inter9));
  nand2 gate3542(.a(s_267), .b(gate1473inter3), .O(gate1473inter10));
  nor2  gate3543(.a(gate1473inter10), .b(gate1473inter9), .O(gate1473inter11));
  nor2  gate3544(.a(gate1473inter11), .b(gate1473inter6), .O(gate1473inter12));
  nand2 gate3545(.a(gate1473inter12), .b(gate1473inter1), .O(N4860));
inv1 gate1474( .a(N4826), .O(N4868) );
inv1 gate1475( .a(N4805), .O(N4870) );
inv1 gate1476( .a(N4808), .O(N4872) );
nand2 gate1477( .a(N4664), .b(N4830), .O(N4873) );
or3 gate1478( .a(N4794), .b(N4797), .c(N4341), .O(N4876) );
nor3 gate1479( .a(N4794), .b(N4797), .c(N4341), .O(N4880) );
inv1 gate1480( .a(N4812), .O(N4885) );
inv1 gate1481( .a(N4822), .O(N4889) );

  xor2  gate3574(.a(N4860), .b(N4859), .O(gate1482inter0));
  nand2 gate3575(.a(gate1482inter0), .b(s_272), .O(gate1482inter1));
  and2  gate3576(.a(N4860), .b(N4859), .O(gate1482inter2));
  inv1  gate3577(.a(s_272), .O(gate1482inter3));
  inv1  gate3578(.a(s_273), .O(gate1482inter4));
  nand2 gate3579(.a(gate1482inter4), .b(gate1482inter3), .O(gate1482inter5));
  nor2  gate3580(.a(gate1482inter5), .b(gate1482inter2), .O(gate1482inter6));
  inv1  gate3581(.a(N4859), .O(gate1482inter7));
  inv1  gate3582(.a(N4860), .O(gate1482inter8));
  nand2 gate3583(.a(gate1482inter8), .b(gate1482inter7), .O(gate1482inter9));
  nand2 gate3584(.a(s_273), .b(gate1482inter3), .O(gate1482inter10));
  nor2  gate3585(.a(gate1482inter10), .b(gate1482inter9), .O(gate1482inter11));
  nor2  gate3586(.a(gate1482inter11), .b(gate1482inter6), .O(gate1482inter12));
  nand2 gate3587(.a(gate1482inter12), .b(gate1482inter1), .O(N4895));
inv1 gate1483( .a(N4844), .O(N4896) );

  xor2  gate2510(.a(N4706), .b(N4844), .O(gate1484inter0));
  nand2 gate2511(.a(gate1484inter0), .b(s_120), .O(gate1484inter1));
  and2  gate2512(.a(N4706), .b(N4844), .O(gate1484inter2));
  inv1  gate2513(.a(s_120), .O(gate1484inter3));
  inv1  gate2514(.a(s_121), .O(gate1484inter4));
  nand2 gate2515(.a(gate1484inter4), .b(gate1484inter3), .O(gate1484inter5));
  nor2  gate2516(.a(gate1484inter5), .b(gate1484inter2), .O(gate1484inter6));
  inv1  gate2517(.a(N4844), .O(gate1484inter7));
  inv1  gate2518(.a(N4706), .O(gate1484inter8));
  nand2 gate2519(.a(gate1484inter8), .b(gate1484inter7), .O(gate1484inter9));
  nand2 gate2520(.a(s_121), .b(gate1484inter3), .O(gate1484inter10));
  nor2  gate2521(.a(gate1484inter10), .b(gate1484inter9), .O(gate1484inter11));
  nor2  gate2522(.a(gate1484inter11), .b(gate1484inter6), .O(gate1484inter12));
  nand2 gate2523(.a(gate1484inter12), .b(gate1484inter1), .O(N4897));
inv1 gate1485( .a(N4847), .O(N4898) );

  xor2  gate1782(.a(N4707), .b(N4847), .O(gate1486inter0));
  nand2 gate1783(.a(gate1486inter0), .b(s_16), .O(gate1486inter1));
  and2  gate1784(.a(N4707), .b(N4847), .O(gate1486inter2));
  inv1  gate1785(.a(s_16), .O(gate1486inter3));
  inv1  gate1786(.a(s_17), .O(gate1486inter4));
  nand2 gate1787(.a(gate1486inter4), .b(gate1486inter3), .O(gate1486inter5));
  nor2  gate1788(.a(gate1486inter5), .b(gate1486inter2), .O(gate1486inter6));
  inv1  gate1789(.a(N4847), .O(gate1486inter7));
  inv1  gate1790(.a(N4707), .O(gate1486inter8));
  nand2 gate1791(.a(gate1486inter8), .b(gate1486inter7), .O(gate1486inter9));
  nand2 gate1792(.a(s_17), .b(gate1486inter3), .O(gate1486inter10));
  nor2  gate1793(.a(gate1486inter10), .b(gate1486inter9), .O(gate1486inter11));
  nor2  gate1794(.a(gate1486inter11), .b(gate1486inter6), .O(gate1486inter12));
  nand2 gate1795(.a(gate1486inter12), .b(gate1486inter1), .O(N4899));

  xor2  gate1768(.a(N4564), .b(N4868), .O(gate1487inter0));
  nand2 gate1769(.a(gate1487inter0), .b(s_14), .O(gate1487inter1));
  and2  gate1770(.a(N4564), .b(N4868), .O(gate1487inter2));
  inv1  gate1771(.a(s_14), .O(gate1487inter3));
  inv1  gate1772(.a(s_15), .O(gate1487inter4));
  nand2 gate1773(.a(gate1487inter4), .b(gate1487inter3), .O(gate1487inter5));
  nor2  gate1774(.a(gate1487inter5), .b(gate1487inter2), .O(gate1487inter6));
  inv1  gate1775(.a(N4868), .O(gate1487inter7));
  inv1  gate1776(.a(N4564), .O(gate1487inter8));
  nand2 gate1777(.a(gate1487inter8), .b(gate1487inter7), .O(gate1487inter9));
  nand2 gate1778(.a(s_15), .b(gate1487inter3), .O(gate1487inter10));
  nor2  gate1779(.a(gate1487inter10), .b(gate1487inter9), .O(gate1487inter11));
  nor2  gate1780(.a(gate1487inter11), .b(gate1487inter6), .O(gate1487inter12));
  nand2 gate1781(.a(gate1487inter12), .b(gate1487inter1), .O(N4900));
and4 gate1488( .a(N4717), .b(N4757), .c(N4823), .d(N4564), .O(N4901) );
inv1 gate1489( .a(N4850), .O(N4902) );
inv1 gate1490( .a(N4854), .O(N4904) );

  xor2  gate4106(.a(N4872), .b(N4854), .O(gate1491inter0));
  nand2 gate4107(.a(gate1491inter0), .b(s_348), .O(gate1491inter1));
  and2  gate4108(.a(N4872), .b(N4854), .O(gate1491inter2));
  inv1  gate4109(.a(s_348), .O(gate1491inter3));
  inv1  gate4110(.a(s_349), .O(gate1491inter4));
  nand2 gate4111(.a(gate1491inter4), .b(gate1491inter3), .O(gate1491inter5));
  nor2  gate4112(.a(gate1491inter5), .b(gate1491inter2), .O(gate1491inter6));
  inv1  gate4113(.a(N4854), .O(gate1491inter7));
  inv1  gate4114(.a(N4872), .O(gate1491inter8));
  nand2 gate4115(.a(gate1491inter8), .b(gate1491inter7), .O(gate1491inter9));
  nand2 gate4116(.a(s_349), .b(gate1491inter3), .O(gate1491inter10));
  nor2  gate4117(.a(gate1491inter10), .b(gate1491inter9), .O(gate1491inter11));
  nor2  gate4118(.a(gate1491inter11), .b(gate1491inter6), .O(gate1491inter12));
  nand2 gate4119(.a(gate1491inter12), .b(gate1491inter1), .O(N4905));

  xor2  gate3854(.a(N4829), .b(N4873), .O(gate1492inter0));
  nand2 gate3855(.a(gate1492inter0), .b(s_312), .O(gate1492inter1));
  and2  gate3856(.a(N4829), .b(N4873), .O(gate1492inter2));
  inv1  gate3857(.a(s_312), .O(gate1492inter3));
  inv1  gate3858(.a(s_313), .O(gate1492inter4));
  nand2 gate3859(.a(gate1492inter4), .b(gate1492inter3), .O(gate1492inter5));
  nor2  gate3860(.a(gate1492inter5), .b(gate1492inter2), .O(gate1492inter6));
  inv1  gate3861(.a(N4873), .O(gate1492inter7));
  inv1  gate3862(.a(N4829), .O(gate1492inter8));
  nand2 gate3863(.a(gate1492inter8), .b(gate1492inter7), .O(gate1492inter9));
  nand2 gate3864(.a(s_313), .b(gate1492inter3), .O(gate1492inter10));
  nor2  gate3865(.a(gate1492inter10), .b(gate1492inter9), .O(gate1492inter11));
  nor2  gate3866(.a(gate1492inter11), .b(gate1492inter6), .O(gate1492inter12));
  nand2 gate3867(.a(gate1492inter12), .b(gate1492inter1), .O(N4906));
and2 gate1493( .a(N4818), .b(N2123), .O(N4907) );
and2 gate1494( .a(N4823), .b(N2125), .O(N4913) );
and2 gate1495( .a(N4818), .b(N4644), .O(N4916) );
inv1 gate1496( .a(N4880), .O(N4920) );
and2 gate1497( .a(N4895), .b(N2184), .O(N4921) );

  xor2  gate2706(.a(N4896), .b(N4656), .O(gate1498inter0));
  nand2 gate2707(.a(gate1498inter0), .b(s_148), .O(gate1498inter1));
  and2  gate2708(.a(N4896), .b(N4656), .O(gate1498inter2));
  inv1  gate2709(.a(s_148), .O(gate1498inter3));
  inv1  gate2710(.a(s_149), .O(gate1498inter4));
  nand2 gate2711(.a(gate1498inter4), .b(gate1498inter3), .O(gate1498inter5));
  nor2  gate2712(.a(gate1498inter5), .b(gate1498inter2), .O(gate1498inter6));
  inv1  gate2713(.a(N4656), .O(gate1498inter7));
  inv1  gate2714(.a(N4896), .O(gate1498inter8));
  nand2 gate2715(.a(gate1498inter8), .b(gate1498inter7), .O(gate1498inter9));
  nand2 gate2716(.a(s_149), .b(gate1498inter3), .O(gate1498inter10));
  nor2  gate2717(.a(gate1498inter10), .b(gate1498inter9), .O(gate1498inter11));
  nor2  gate2718(.a(gate1498inter11), .b(gate1498inter6), .O(gate1498inter12));
  nand2 gate2719(.a(gate1498inter12), .b(gate1498inter1), .O(N4924));

  xor2  gate4302(.a(N4898), .b(N4659), .O(gate1499inter0));
  nand2 gate4303(.a(gate1499inter0), .b(s_376), .O(gate1499inter1));
  and2  gate4304(.a(N4898), .b(N4659), .O(gate1499inter2));
  inv1  gate4305(.a(s_376), .O(gate1499inter3));
  inv1  gate4306(.a(s_377), .O(gate1499inter4));
  nand2 gate4307(.a(gate1499inter4), .b(gate1499inter3), .O(gate1499inter5));
  nor2  gate4308(.a(gate1499inter5), .b(gate1499inter2), .O(gate1499inter6));
  inv1  gate4309(.a(N4659), .O(gate1499inter7));
  inv1  gate4310(.a(N4898), .O(gate1499inter8));
  nand2 gate4311(.a(gate1499inter8), .b(gate1499inter7), .O(gate1499inter9));
  nand2 gate4312(.a(s_377), .b(gate1499inter3), .O(gate1499inter10));
  nor2  gate4313(.a(gate1499inter10), .b(gate1499inter9), .O(gate1499inter11));
  nor2  gate4314(.a(gate1499inter11), .b(gate1499inter6), .O(gate1499inter12));
  nand2 gate4315(.a(gate1499inter12), .b(gate1499inter1), .O(N4925));
or2 gate1500( .a(N4900), .b(N4901), .O(N4926) );

  xor2  gate2594(.a(N4870), .b(N4889), .O(gate1501inter0));
  nand2 gate2595(.a(gate1501inter0), .b(s_132), .O(gate1501inter1));
  and2  gate2596(.a(N4870), .b(N4889), .O(gate1501inter2));
  inv1  gate2597(.a(s_132), .O(gate1501inter3));
  inv1  gate2598(.a(s_133), .O(gate1501inter4));
  nand2 gate2599(.a(gate1501inter4), .b(gate1501inter3), .O(gate1501inter5));
  nor2  gate2600(.a(gate1501inter5), .b(gate1501inter2), .O(gate1501inter6));
  inv1  gate2601(.a(N4889), .O(gate1501inter7));
  inv1  gate2602(.a(N4870), .O(gate1501inter8));
  nand2 gate2603(.a(gate1501inter8), .b(gate1501inter7), .O(gate1501inter9));
  nand2 gate2604(.a(s_133), .b(gate1501inter3), .O(gate1501inter10));
  nor2  gate2605(.a(gate1501inter10), .b(gate1501inter9), .O(gate1501inter11));
  nor2  gate2606(.a(gate1501inter11), .b(gate1501inter6), .O(gate1501inter12));
  nand2 gate2607(.a(gate1501inter12), .b(gate1501inter1), .O(N4928));
inv1 gate1502( .a(N4889), .O(N4929) );

  xor2  gate2818(.a(N4904), .b(N4808), .O(gate1503inter0));
  nand2 gate2819(.a(gate1503inter0), .b(s_164), .O(gate1503inter1));
  and2  gate2820(.a(N4904), .b(N4808), .O(gate1503inter2));
  inv1  gate2821(.a(s_164), .O(gate1503inter3));
  inv1  gate2822(.a(s_165), .O(gate1503inter4));
  nand2 gate2823(.a(gate1503inter4), .b(gate1503inter3), .O(gate1503inter5));
  nor2  gate2824(.a(gate1503inter5), .b(gate1503inter2), .O(gate1503inter6));
  inv1  gate2825(.a(N4808), .O(gate1503inter7));
  inv1  gate2826(.a(N4904), .O(gate1503inter8));
  nand2 gate2827(.a(gate1503inter8), .b(gate1503inter7), .O(gate1503inter9));
  nand2 gate2828(.a(s_165), .b(gate1503inter3), .O(gate1503inter10));
  nor2  gate2829(.a(gate1503inter10), .b(gate1503inter9), .O(gate1503inter11));
  nor2  gate2830(.a(gate1503inter11), .b(gate1503inter6), .O(gate1503inter12));
  nand2 gate2831(.a(gate1503inter12), .b(gate1503inter1), .O(N4930));
inv1 gate1504( .a(N4906), .O(N4931) );
buf1 gate1505( .a(N4876), .O(N4937) );
buf1 gate1506( .a(N4876), .O(N4940) );
and2 gate1507( .a(N4876), .b(N4920), .O(N4944) );
nand2 gate1508( .a(N4924), .b(N4897), .O(N4946) );

  xor2  gate4176(.a(N4899), .b(N4925), .O(gate1509inter0));
  nand2 gate4177(.a(gate1509inter0), .b(s_358), .O(gate1509inter1));
  and2  gate4178(.a(N4899), .b(N4925), .O(gate1509inter2));
  inv1  gate4179(.a(s_358), .O(gate1509inter3));
  inv1  gate4180(.a(s_359), .O(gate1509inter4));
  nand2 gate4181(.a(gate1509inter4), .b(gate1509inter3), .O(gate1509inter5));
  nor2  gate4182(.a(gate1509inter5), .b(gate1509inter2), .O(gate1509inter6));
  inv1  gate4183(.a(N4925), .O(gate1509inter7));
  inv1  gate4184(.a(N4899), .O(gate1509inter8));
  nand2 gate4185(.a(gate1509inter8), .b(gate1509inter7), .O(gate1509inter9));
  nand2 gate4186(.a(s_359), .b(gate1509inter3), .O(gate1509inter10));
  nor2  gate4187(.a(gate1509inter10), .b(gate1509inter9), .O(gate1509inter11));
  nor2  gate4188(.a(gate1509inter11), .b(gate1509inter6), .O(gate1509inter12));
  nand2 gate4189(.a(gate1509inter12), .b(gate1509inter1), .O(N4949));
nand2 gate1510( .a(N4916), .b(N4902), .O(N4950) );
inv1 gate1511( .a(N4916), .O(N4951) );
nand2 gate1512( .a(N4805), .b(N4929), .O(N4952) );

  xor2  gate2916(.a(N4905), .b(N4930), .O(gate1513inter0));
  nand2 gate2917(.a(gate1513inter0), .b(s_178), .O(gate1513inter1));
  and2  gate2918(.a(N4905), .b(N4930), .O(gate1513inter2));
  inv1  gate2919(.a(s_178), .O(gate1513inter3));
  inv1  gate2920(.a(s_179), .O(gate1513inter4));
  nand2 gate2921(.a(gate1513inter4), .b(gate1513inter3), .O(gate1513inter5));
  nor2  gate2922(.a(gate1513inter5), .b(gate1513inter2), .O(gate1513inter6));
  inv1  gate2923(.a(N4930), .O(gate1513inter7));
  inv1  gate2924(.a(N4905), .O(gate1513inter8));
  nand2 gate2925(.a(gate1513inter8), .b(gate1513inter7), .O(gate1513inter9));
  nand2 gate2926(.a(s_179), .b(gate1513inter3), .O(gate1513inter10));
  nor2  gate2927(.a(gate1513inter10), .b(gate1513inter9), .O(gate1513inter11));
  nor2  gate2928(.a(gate1513inter11), .b(gate1513inter6), .O(gate1513inter12));
  nand2 gate2929(.a(gate1513inter12), .b(gate1513inter1), .O(N4953));
and2 gate1514( .a(N4926), .b(N2737), .O(N4954) );
and2 gate1515( .a(N4931), .b(N2741), .O(N4957) );
or3 gate1516( .a(N2764), .b(N2483), .c(N4921), .O(N4964) );
nor3 gate1517( .a(N2764), .b(N2483), .c(N4921), .O(N4965) );
inv1 gate1518( .a(N4949), .O(N4968) );

  xor2  gate3504(.a(N4951), .b(N4850), .O(gate1519inter0));
  nand2 gate3505(.a(gate1519inter0), .b(s_262), .O(gate1519inter1));
  and2  gate3506(.a(N4951), .b(N4850), .O(gate1519inter2));
  inv1  gate3507(.a(s_262), .O(gate1519inter3));
  inv1  gate3508(.a(s_263), .O(gate1519inter4));
  nand2 gate3509(.a(gate1519inter4), .b(gate1519inter3), .O(gate1519inter5));
  nor2  gate3510(.a(gate1519inter5), .b(gate1519inter2), .O(gate1519inter6));
  inv1  gate3511(.a(N4850), .O(gate1519inter7));
  inv1  gate3512(.a(N4951), .O(gate1519inter8));
  nand2 gate3513(.a(gate1519inter8), .b(gate1519inter7), .O(gate1519inter9));
  nand2 gate3514(.a(s_263), .b(gate1519inter3), .O(gate1519inter10));
  nor2  gate3515(.a(gate1519inter10), .b(gate1519inter9), .O(gate1519inter11));
  nor2  gate3516(.a(gate1519inter11), .b(gate1519inter6), .O(gate1519inter12));
  nand2 gate3517(.a(gate1519inter12), .b(gate1519inter1), .O(N4969));

  xor2  gate3742(.a(N4928), .b(N4952), .O(gate1520inter0));
  nand2 gate3743(.a(gate1520inter0), .b(s_296), .O(gate1520inter1));
  and2  gate3744(.a(N4928), .b(N4952), .O(gate1520inter2));
  inv1  gate3745(.a(s_296), .O(gate1520inter3));
  inv1  gate3746(.a(s_297), .O(gate1520inter4));
  nand2 gate3747(.a(gate1520inter4), .b(gate1520inter3), .O(gate1520inter5));
  nor2  gate3748(.a(gate1520inter5), .b(gate1520inter2), .O(gate1520inter6));
  inv1  gate3749(.a(N4952), .O(gate1520inter7));
  inv1  gate3750(.a(N4928), .O(gate1520inter8));
  nand2 gate3751(.a(gate1520inter8), .b(gate1520inter7), .O(gate1520inter9));
  nand2 gate3752(.a(s_297), .b(gate1520inter3), .O(gate1520inter10));
  nor2  gate3753(.a(gate1520inter10), .b(gate1520inter9), .O(gate1520inter11));
  nor2  gate3754(.a(gate1520inter11), .b(gate1520inter6), .O(gate1520inter12));
  nand2 gate3755(.a(gate1520inter12), .b(gate1520inter1), .O(N4970));
and2 gate1521( .a(N4953), .b(N2739), .O(N4973) );
inv1 gate1522( .a(N4937), .O(N4978) );
inv1 gate1523( .a(N4940), .O(N4979) );
inv1 gate1524( .a(N4965), .O(N4980) );
nor2 gate1525( .a(N4968), .b(N4722), .O(N4981) );
and4 gate1526( .a(N4818), .b(N4743), .c(N4946), .d(N4722), .O(N4982) );

  xor2  gate2790(.a(N4969), .b(N4950), .O(gate1527inter0));
  nand2 gate2791(.a(gate1527inter0), .b(s_160), .O(gate1527inter1));
  and2  gate2792(.a(N4969), .b(N4950), .O(gate1527inter2));
  inv1  gate2793(.a(s_160), .O(gate1527inter3));
  inv1  gate2794(.a(s_161), .O(gate1527inter4));
  nand2 gate2795(.a(gate1527inter4), .b(gate1527inter3), .O(gate1527inter5));
  nor2  gate2796(.a(gate1527inter5), .b(gate1527inter2), .O(gate1527inter6));
  inv1  gate2797(.a(N4950), .O(gate1527inter7));
  inv1  gate2798(.a(N4969), .O(gate1527inter8));
  nand2 gate2799(.a(gate1527inter8), .b(gate1527inter7), .O(gate1527inter9));
  nand2 gate2800(.a(s_161), .b(gate1527inter3), .O(gate1527inter10));
  nor2  gate2801(.a(gate1527inter10), .b(gate1527inter9), .O(gate1527inter11));
  nor2  gate2802(.a(gate1527inter11), .b(gate1527inter6), .O(gate1527inter12));
  nand2 gate2803(.a(gate1527inter12), .b(gate1527inter1), .O(N4983));
inv1 gate1528( .a(N4970), .O(N4984) );
and2 gate1529( .a(N4946), .b(N2121), .O(N4985) );
or3 gate1530( .a(N4913), .b(N4954), .c(N4344), .O(N4988) );
nor3 gate1531( .a(N4913), .b(N4954), .c(N4344), .O(N4991) );
or3 gate1532( .a(N4800), .b(N4957), .c(N4347), .O(N4996) );
nor3 gate1533( .a(N4800), .b(N4957), .c(N4347), .O(N4999) );
and2 gate1534( .a(N4964), .b(N4980), .O(N5002) );
or2 gate1535( .a(N4981), .b(N4982), .O(N5007) );
and2 gate1536( .a(N4983), .b(N2731), .O(N5010) );
and2 gate1537( .a(N4984), .b(N2733), .O(N5013) );
or3 gate1538( .a(N4838), .b(N4973), .c(N4475), .O(N5018) );
nor3 gate1539( .a(N4838), .b(N4973), .c(N4475), .O(N5021) );
inv1 gate1540( .a(N4991), .O(N5026) );
inv1 gate1541( .a(N4999), .O(N5029) );
and2 gate1542( .a(N5007), .b(N2729), .O(N5030) );
buf1 gate1543( .a(N4996), .O(N5039) );
buf1 gate1544( .a(N4988), .O(N5042) );
and2 gate1545( .a(N4988), .b(N5026), .O(N5045) );
inv1 gate1546( .a(N5021), .O(N5046) );
and2 gate1547( .a(N4996), .b(N5029), .O(N5047) );
or3 gate1548( .a(N4831), .b(N5010), .c(N4472), .O(N5050) );
nor3 gate1549( .a(N4831), .b(N5010), .c(N4472), .O(N5055) );
or3 gate1550( .a(N4907), .b(N5013), .c(N4338), .O(N5058) );
nor3 gate1551( .a(N4907), .b(N5013), .c(N4338), .O(N5061) );
and4 gate1552( .a(N4730), .b(N4999), .c(N5021), .d(N4991), .O(N5066) );
buf1 gate1553( .a(N5018), .O(N5070) );
and2 gate1554( .a(N5018), .b(N5046), .O(N5078) );
or3 gate1555( .a(N4985), .b(N5030), .c(N4335), .O(N5080) );
nor3 gate1556( .a(N4985), .b(N5030), .c(N4335), .O(N5085) );

  xor2  gate2902(.a(N4885), .b(N5039), .O(gate1557inter0));
  nand2 gate2903(.a(gate1557inter0), .b(s_176), .O(gate1557inter1));
  and2  gate2904(.a(N4885), .b(N5039), .O(gate1557inter2));
  inv1  gate2905(.a(s_176), .O(gate1557inter3));
  inv1  gate2906(.a(s_177), .O(gate1557inter4));
  nand2 gate2907(.a(gate1557inter4), .b(gate1557inter3), .O(gate1557inter5));
  nor2  gate2908(.a(gate1557inter5), .b(gate1557inter2), .O(gate1557inter6));
  inv1  gate2909(.a(N5039), .O(gate1557inter7));
  inv1  gate2910(.a(N4885), .O(gate1557inter8));
  nand2 gate2911(.a(gate1557inter8), .b(gate1557inter7), .O(gate1557inter9));
  nand2 gate2912(.a(s_177), .b(gate1557inter3), .O(gate1557inter10));
  nor2  gate2913(.a(gate1557inter10), .b(gate1557inter9), .O(gate1557inter11));
  nor2  gate2914(.a(gate1557inter11), .b(gate1557inter6), .O(gate1557inter12));
  nand2 gate2915(.a(gate1557inter12), .b(gate1557inter1), .O(N5094));
inv1 gate1558( .a(N5039), .O(N5095) );
inv1 gate1559( .a(N5042), .O(N5097) );
and2 gate1560( .a(N5050), .b(N5050), .O(N5102) );
inv1 gate1561( .a(N5061), .O(N5103) );

  xor2  gate2622(.a(N5095), .b(N4812), .O(gate1562inter0));
  nand2 gate2623(.a(gate1562inter0), .b(s_136), .O(gate1562inter1));
  and2  gate2624(.a(N5095), .b(N4812), .O(gate1562inter2));
  inv1  gate2625(.a(s_136), .O(gate1562inter3));
  inv1  gate2626(.a(s_137), .O(gate1562inter4));
  nand2 gate2627(.a(gate1562inter4), .b(gate1562inter3), .O(gate1562inter5));
  nor2  gate2628(.a(gate1562inter5), .b(gate1562inter2), .O(gate1562inter6));
  inv1  gate2629(.a(N4812), .O(gate1562inter7));
  inv1  gate2630(.a(N5095), .O(gate1562inter8));
  nand2 gate2631(.a(gate1562inter8), .b(gate1562inter7), .O(gate1562inter9));
  nand2 gate2632(.a(s_137), .b(gate1562inter3), .O(gate1562inter10));
  nor2  gate2633(.a(gate1562inter10), .b(gate1562inter9), .O(gate1562inter11));
  nor2  gate2634(.a(gate1562inter11), .b(gate1562inter6), .O(gate1562inter12));
  nand2 gate2635(.a(gate1562inter12), .b(gate1562inter1), .O(N5108));
inv1 gate1563( .a(N5070), .O(N5109) );

  xor2  gate4358(.a(N5097), .b(N5070), .O(gate1564inter0));
  nand2 gate4359(.a(gate1564inter0), .b(s_384), .O(gate1564inter1));
  and2  gate4360(.a(N5097), .b(N5070), .O(gate1564inter2));
  inv1  gate4361(.a(s_384), .O(gate1564inter3));
  inv1  gate4362(.a(s_385), .O(gate1564inter4));
  nand2 gate4363(.a(gate1564inter4), .b(gate1564inter3), .O(gate1564inter5));
  nor2  gate4364(.a(gate1564inter5), .b(gate1564inter2), .O(gate1564inter6));
  inv1  gate4365(.a(N5070), .O(gate1564inter7));
  inv1  gate4366(.a(N5097), .O(gate1564inter8));
  nand2 gate4367(.a(gate1564inter8), .b(gate1564inter7), .O(gate1564inter9));
  nand2 gate4368(.a(s_385), .b(gate1564inter3), .O(gate1564inter10));
  nor2  gate4369(.a(gate1564inter10), .b(gate1564inter9), .O(gate1564inter11));
  nor2  gate4370(.a(gate1564inter11), .b(gate1564inter6), .O(gate1564inter12));
  nand2 gate4371(.a(gate1564inter12), .b(gate1564inter1), .O(N5110));
buf1 gate1565( .a(N5058), .O(N5111) );
and2 gate1566( .a(N5050), .b(N1461), .O(N5114) );
buf1 gate1567( .a(N5050), .O(N5117) );
and2 gate1568( .a(N5080), .b(N5080), .O(N5120) );
and2 gate1569( .a(N5058), .b(N5103), .O(N5121) );
nand2 gate1570( .a(N5094), .b(N5108), .O(N5122) );

  xor2  gate3546(.a(N5109), .b(N5042), .O(gate1571inter0));
  nand2 gate3547(.a(gate1571inter0), .b(s_268), .O(gate1571inter1));
  and2  gate3548(.a(N5109), .b(N5042), .O(gate1571inter2));
  inv1  gate3549(.a(s_268), .O(gate1571inter3));
  inv1  gate3550(.a(s_269), .O(gate1571inter4));
  nand2 gate3551(.a(gate1571inter4), .b(gate1571inter3), .O(gate1571inter5));
  nor2  gate3552(.a(gate1571inter5), .b(gate1571inter2), .O(gate1571inter6));
  inv1  gate3553(.a(N5042), .O(gate1571inter7));
  inv1  gate3554(.a(N5109), .O(gate1571inter8));
  nand2 gate3555(.a(gate1571inter8), .b(gate1571inter7), .O(gate1571inter9));
  nand2 gate3556(.a(s_269), .b(gate1571inter3), .O(gate1571inter10));
  nor2  gate3557(.a(gate1571inter10), .b(gate1571inter9), .O(gate1571inter11));
  nor2  gate3558(.a(gate1571inter11), .b(gate1571inter6), .O(gate1571inter12));
  nand2 gate3559(.a(gate1571inter12), .b(gate1571inter1), .O(N5125));
and2 gate1572( .a(N1461), .b(N5080), .O(N5128) );
and4 gate1573( .a(N4880), .b(N5061), .c(N5055), .d(N5085), .O(N5133) );
and3 gate1574( .a(N5055), .b(N5085), .c(N1464), .O(N5136) );
buf1 gate1575( .a(N5080), .O(N5139) );

  xor2  gate2006(.a(N5110), .b(N5125), .O(gate1576inter0));
  nand2 gate2007(.a(gate1576inter0), .b(s_48), .O(gate1576inter1));
  and2  gate2008(.a(N5110), .b(N5125), .O(gate1576inter2));
  inv1  gate2009(.a(s_48), .O(gate1576inter3));
  inv1  gate2010(.a(s_49), .O(gate1576inter4));
  nand2 gate2011(.a(gate1576inter4), .b(gate1576inter3), .O(gate1576inter5));
  nor2  gate2012(.a(gate1576inter5), .b(gate1576inter2), .O(gate1576inter6));
  inv1  gate2013(.a(N5125), .O(gate1576inter7));
  inv1  gate2014(.a(N5110), .O(gate1576inter8));
  nand2 gate2015(.a(gate1576inter8), .b(gate1576inter7), .O(gate1576inter9));
  nand2 gate2016(.a(s_49), .b(gate1576inter3), .O(gate1576inter10));
  nor2  gate2017(.a(gate1576inter10), .b(gate1576inter9), .O(gate1576inter11));
  nor2  gate2018(.a(gate1576inter11), .b(gate1576inter6), .O(gate1576inter12));
  nand2 gate2019(.a(gate1576inter12), .b(gate1576inter1), .O(N5145));
buf1 gate1577( .a(N5111), .O(N5151) );
buf1 gate1578( .a(N5111), .O(N5154) );
inv1 gate1579( .a(N5117), .O(N5159) );
buf1 gate1580( .a(N5114), .O(N5160) );
buf1 gate1581( .a(N5114), .O(N5163) );
and2 gate1582( .a(N5066), .b(N5133), .O(N5166) );
and2 gate1583( .a(N5066), .b(N5133), .O(N5173) );
buf1 gate1584( .a(N5122), .O(N5174) );
buf1 gate1585( .a(N5122), .O(N5177) );
inv1 gate1586( .a(N5139), .O(N5182) );
nand2 gate1587( .a(N5139), .b(N5159), .O(N5183) );
buf1 gate1588( .a(N5128), .O(N5184) );
buf1 gate1589( .a(N5128), .O(N5188) );
inv1 gate1590( .a(N5166), .O(N5192) );

  xor2  gate2300(.a(N5173), .b(N5136), .O(gate1591inter0));
  nand2 gate2301(.a(gate1591inter0), .b(s_90), .O(gate1591inter1));
  and2  gate2302(.a(N5173), .b(N5136), .O(gate1591inter2));
  inv1  gate2303(.a(s_90), .O(gate1591inter3));
  inv1  gate2304(.a(s_91), .O(gate1591inter4));
  nand2 gate2305(.a(gate1591inter4), .b(gate1591inter3), .O(gate1591inter5));
  nor2  gate2306(.a(gate1591inter5), .b(gate1591inter2), .O(gate1591inter6));
  inv1  gate2307(.a(N5136), .O(gate1591inter7));
  inv1  gate2308(.a(N5173), .O(gate1591inter8));
  nand2 gate2309(.a(gate1591inter8), .b(gate1591inter7), .O(gate1591inter9));
  nand2 gate2310(.a(s_91), .b(gate1591inter3), .O(gate1591inter10));
  nor2  gate2311(.a(gate1591inter10), .b(gate1591inter9), .O(gate1591inter11));
  nor2  gate2312(.a(gate1591inter11), .b(gate1591inter6), .O(gate1591inter12));
  nand2 gate2313(.a(gate1591inter12), .b(gate1591inter1), .O(N5193));
nand2 gate1592( .a(N5151), .b(N4978), .O(N5196) );
inv1 gate1593( .a(N5151), .O(N5197) );

  xor2  gate4050(.a(N4979), .b(N5154), .O(gate1594inter0));
  nand2 gate4051(.a(gate1594inter0), .b(s_340), .O(gate1594inter1));
  and2  gate4052(.a(N4979), .b(N5154), .O(gate1594inter2));
  inv1  gate4053(.a(s_340), .O(gate1594inter3));
  inv1  gate4054(.a(s_341), .O(gate1594inter4));
  nand2 gate4055(.a(gate1594inter4), .b(gate1594inter3), .O(gate1594inter5));
  nor2  gate4056(.a(gate1594inter5), .b(gate1594inter2), .O(gate1594inter6));
  inv1  gate4057(.a(N5154), .O(gate1594inter7));
  inv1  gate4058(.a(N4979), .O(gate1594inter8));
  nand2 gate4059(.a(gate1594inter8), .b(gate1594inter7), .O(gate1594inter9));
  nand2 gate4060(.a(s_341), .b(gate1594inter3), .O(gate1594inter10));
  nor2  gate4061(.a(gate1594inter10), .b(gate1594inter9), .O(gate1594inter11));
  nor2  gate4062(.a(gate1594inter11), .b(gate1594inter6), .O(gate1594inter12));
  nand2 gate4063(.a(gate1594inter12), .b(gate1594inter1), .O(N5198));
inv1 gate1595( .a(N5154), .O(N5199) );
inv1 gate1596( .a(N5160), .O(N5201) );
inv1 gate1597( .a(N5163), .O(N5203) );
buf1 gate1598( .a(N5145), .O(N5205) );
buf1 gate1599( .a(N5145), .O(N5209) );

  xor2  gate2958(.a(N5182), .b(N5117), .O(gate1600inter0));
  nand2 gate2959(.a(gate1600inter0), .b(s_184), .O(gate1600inter1));
  and2  gate2960(.a(N5182), .b(N5117), .O(gate1600inter2));
  inv1  gate2961(.a(s_184), .O(gate1600inter3));
  inv1  gate2962(.a(s_185), .O(gate1600inter4));
  nand2 gate2963(.a(gate1600inter4), .b(gate1600inter3), .O(gate1600inter5));
  nor2  gate2964(.a(gate1600inter5), .b(gate1600inter2), .O(gate1600inter6));
  inv1  gate2965(.a(N5117), .O(gate1600inter7));
  inv1  gate2966(.a(N5182), .O(gate1600inter8));
  nand2 gate2967(.a(gate1600inter8), .b(gate1600inter7), .O(gate1600inter9));
  nand2 gate2968(.a(s_185), .b(gate1600inter3), .O(gate1600inter10));
  nor2  gate2969(.a(gate1600inter10), .b(gate1600inter9), .O(gate1600inter11));
  nor2  gate2970(.a(gate1600inter11), .b(gate1600inter6), .O(gate1600inter12));
  nand2 gate2971(.a(gate1600inter12), .b(gate1600inter1), .O(N5212));
and2 gate1601( .a(N213), .b(N5193), .O(N5215) );
inv1 gate1602( .a(N5174), .O(N5217) );
inv1 gate1603( .a(N5177), .O(N5219) );

  xor2  gate2538(.a(N5197), .b(N4937), .O(gate1604inter0));
  nand2 gate2539(.a(gate1604inter0), .b(s_124), .O(gate1604inter1));
  and2  gate2540(.a(N5197), .b(N4937), .O(gate1604inter2));
  inv1  gate2541(.a(s_124), .O(gate1604inter3));
  inv1  gate2542(.a(s_125), .O(gate1604inter4));
  nand2 gate2543(.a(gate1604inter4), .b(gate1604inter3), .O(gate1604inter5));
  nor2  gate2544(.a(gate1604inter5), .b(gate1604inter2), .O(gate1604inter6));
  inv1  gate2545(.a(N4937), .O(gate1604inter7));
  inv1  gate2546(.a(N5197), .O(gate1604inter8));
  nand2 gate2547(.a(gate1604inter8), .b(gate1604inter7), .O(gate1604inter9));
  nand2 gate2548(.a(s_125), .b(gate1604inter3), .O(gate1604inter10));
  nor2  gate2549(.a(gate1604inter10), .b(gate1604inter9), .O(gate1604inter11));
  nor2  gate2550(.a(gate1604inter11), .b(gate1604inter6), .O(gate1604inter12));
  nand2 gate2551(.a(gate1604inter12), .b(gate1604inter1), .O(N5220));

  xor2  gate4120(.a(N5199), .b(N4940), .O(gate1605inter0));
  nand2 gate4121(.a(gate1605inter0), .b(s_350), .O(gate1605inter1));
  and2  gate4122(.a(N5199), .b(N4940), .O(gate1605inter2));
  inv1  gate4123(.a(s_350), .O(gate1605inter3));
  inv1  gate4124(.a(s_351), .O(gate1605inter4));
  nand2 gate4125(.a(gate1605inter4), .b(gate1605inter3), .O(gate1605inter5));
  nor2  gate4126(.a(gate1605inter5), .b(gate1605inter2), .O(gate1605inter6));
  inv1  gate4127(.a(N4940), .O(gate1605inter7));
  inv1  gate4128(.a(N5199), .O(gate1605inter8));
  nand2 gate4129(.a(gate1605inter8), .b(gate1605inter7), .O(gate1605inter9));
  nand2 gate4130(.a(s_351), .b(gate1605inter3), .O(gate1605inter10));
  nor2  gate4131(.a(gate1605inter10), .b(gate1605inter9), .O(gate1605inter11));
  nor2  gate4132(.a(gate1605inter11), .b(gate1605inter6), .O(gate1605inter12));
  nand2 gate4133(.a(gate1605inter12), .b(gate1605inter1), .O(N5221));
inv1 gate1606( .a(N5184), .O(N5222) );

  xor2  gate2482(.a(N5201), .b(N5184), .O(gate1607inter0));
  nand2 gate2483(.a(gate1607inter0), .b(s_116), .O(gate1607inter1));
  and2  gate2484(.a(N5201), .b(N5184), .O(gate1607inter2));
  inv1  gate2485(.a(s_116), .O(gate1607inter3));
  inv1  gate2486(.a(s_117), .O(gate1607inter4));
  nand2 gate2487(.a(gate1607inter4), .b(gate1607inter3), .O(gate1607inter5));
  nor2  gate2488(.a(gate1607inter5), .b(gate1607inter2), .O(gate1607inter6));
  inv1  gate2489(.a(N5184), .O(gate1607inter7));
  inv1  gate2490(.a(N5201), .O(gate1607inter8));
  nand2 gate2491(.a(gate1607inter8), .b(gate1607inter7), .O(gate1607inter9));
  nand2 gate2492(.a(s_117), .b(gate1607inter3), .O(gate1607inter10));
  nor2  gate2493(.a(gate1607inter10), .b(gate1607inter9), .O(gate1607inter11));
  nor2  gate2494(.a(gate1607inter11), .b(gate1607inter6), .O(gate1607inter12));
  nand2 gate2495(.a(gate1607inter12), .b(gate1607inter1), .O(N5223));

  xor2  gate2146(.a(N5203), .b(N5188), .O(gate1608inter0));
  nand2 gate2147(.a(gate1608inter0), .b(s_68), .O(gate1608inter1));
  and2  gate2148(.a(N5203), .b(N5188), .O(gate1608inter2));
  inv1  gate2149(.a(s_68), .O(gate1608inter3));
  inv1  gate2150(.a(s_69), .O(gate1608inter4));
  nand2 gate2151(.a(gate1608inter4), .b(gate1608inter3), .O(gate1608inter5));
  nor2  gate2152(.a(gate1608inter5), .b(gate1608inter2), .O(gate1608inter6));
  inv1  gate2153(.a(N5188), .O(gate1608inter7));
  inv1  gate2154(.a(N5203), .O(gate1608inter8));
  nand2 gate2155(.a(gate1608inter8), .b(gate1608inter7), .O(gate1608inter9));
  nand2 gate2156(.a(s_69), .b(gate1608inter3), .O(gate1608inter10));
  nor2  gate2157(.a(gate1608inter10), .b(gate1608inter9), .O(gate1608inter11));
  nor2  gate2158(.a(gate1608inter11), .b(gate1608inter6), .O(gate1608inter12));
  nand2 gate2159(.a(gate1608inter12), .b(gate1608inter1), .O(N5224));
inv1 gate1609( .a(N5188), .O(N5225) );

  xor2  gate2356(.a(N5212), .b(N5183), .O(gate1610inter0));
  nand2 gate2357(.a(gate1610inter0), .b(s_98), .O(gate1610inter1));
  and2  gate2358(.a(N5212), .b(N5183), .O(gate1610inter2));
  inv1  gate2359(.a(s_98), .O(gate1610inter3));
  inv1  gate2360(.a(s_99), .O(gate1610inter4));
  nand2 gate2361(.a(gate1610inter4), .b(gate1610inter3), .O(gate1610inter5));
  nor2  gate2362(.a(gate1610inter5), .b(gate1610inter2), .O(gate1610inter6));
  inv1  gate2363(.a(N5183), .O(gate1610inter7));
  inv1  gate2364(.a(N5212), .O(gate1610inter8));
  nand2 gate2365(.a(gate1610inter8), .b(gate1610inter7), .O(gate1610inter9));
  nand2 gate2366(.a(s_99), .b(gate1610inter3), .O(gate1610inter10));
  nor2  gate2367(.a(gate1610inter10), .b(gate1610inter9), .O(gate1610inter11));
  nor2  gate2368(.a(gate1610inter11), .b(gate1610inter6), .O(gate1610inter12));
  nand2 gate2369(.a(gate1610inter12), .b(gate1610inter1), .O(N5228));
inv1 gate1611( .a(N5215), .O(N5231) );
nand2 gate1612( .a(N5205), .b(N5217), .O(N5232) );
inv1 gate1613( .a(N5205), .O(N5233) );

  xor2  gate2314(.a(N5219), .b(N5209), .O(gate1614inter0));
  nand2 gate2315(.a(gate1614inter0), .b(s_92), .O(gate1614inter1));
  and2  gate2316(.a(N5219), .b(N5209), .O(gate1614inter2));
  inv1  gate2317(.a(s_92), .O(gate1614inter3));
  inv1  gate2318(.a(s_93), .O(gate1614inter4));
  nand2 gate2319(.a(gate1614inter4), .b(gate1614inter3), .O(gate1614inter5));
  nor2  gate2320(.a(gate1614inter5), .b(gate1614inter2), .O(gate1614inter6));
  inv1  gate2321(.a(N5209), .O(gate1614inter7));
  inv1  gate2322(.a(N5219), .O(gate1614inter8));
  nand2 gate2323(.a(gate1614inter8), .b(gate1614inter7), .O(gate1614inter9));
  nand2 gate2324(.a(s_93), .b(gate1614inter3), .O(gate1614inter10));
  nor2  gate2325(.a(gate1614inter10), .b(gate1614inter9), .O(gate1614inter11));
  nor2  gate2326(.a(gate1614inter11), .b(gate1614inter6), .O(gate1614inter12));
  nand2 gate2327(.a(gate1614inter12), .b(gate1614inter1), .O(N5234));
inv1 gate1615( .a(N5209), .O(N5235) );

  xor2  gate1810(.a(N5220), .b(N5196), .O(gate1616inter0));
  nand2 gate1811(.a(gate1616inter0), .b(s_20), .O(gate1616inter1));
  and2  gate1812(.a(N5220), .b(N5196), .O(gate1616inter2));
  inv1  gate1813(.a(s_20), .O(gate1616inter3));
  inv1  gate1814(.a(s_21), .O(gate1616inter4));
  nand2 gate1815(.a(gate1616inter4), .b(gate1616inter3), .O(gate1616inter5));
  nor2  gate1816(.a(gate1616inter5), .b(gate1616inter2), .O(gate1616inter6));
  inv1  gate1817(.a(N5196), .O(gate1616inter7));
  inv1  gate1818(.a(N5220), .O(gate1616inter8));
  nand2 gate1819(.a(gate1616inter8), .b(gate1616inter7), .O(gate1616inter9));
  nand2 gate1820(.a(s_21), .b(gate1616inter3), .O(gate1616inter10));
  nor2  gate1821(.a(gate1616inter10), .b(gate1616inter9), .O(gate1616inter11));
  nor2  gate1822(.a(gate1616inter11), .b(gate1616inter6), .O(gate1616inter12));
  nand2 gate1823(.a(gate1616inter12), .b(gate1616inter1), .O(N5236));
nand2 gate1617( .a(N5198), .b(N5221), .O(N5240) );

  xor2  gate3994(.a(N5222), .b(N5160), .O(gate1618inter0));
  nand2 gate3995(.a(gate1618inter0), .b(s_332), .O(gate1618inter1));
  and2  gate3996(.a(N5222), .b(N5160), .O(gate1618inter2));
  inv1  gate3997(.a(s_332), .O(gate1618inter3));
  inv1  gate3998(.a(s_333), .O(gate1618inter4));
  nand2 gate3999(.a(gate1618inter4), .b(gate1618inter3), .O(gate1618inter5));
  nor2  gate4000(.a(gate1618inter5), .b(gate1618inter2), .O(gate1618inter6));
  inv1  gate4001(.a(N5160), .O(gate1618inter7));
  inv1  gate4002(.a(N5222), .O(gate1618inter8));
  nand2 gate4003(.a(gate1618inter8), .b(gate1618inter7), .O(gate1618inter9));
  nand2 gate4004(.a(s_333), .b(gate1618inter3), .O(gate1618inter10));
  nor2  gate4005(.a(gate1618inter10), .b(gate1618inter9), .O(gate1618inter11));
  nor2  gate4006(.a(gate1618inter11), .b(gate1618inter6), .O(gate1618inter12));
  nand2 gate4007(.a(gate1618inter12), .b(gate1618inter1), .O(N5242));

  xor2  gate3784(.a(N5225), .b(N5163), .O(gate1619inter0));
  nand2 gate3785(.a(gate1619inter0), .b(s_302), .O(gate1619inter1));
  and2  gate3786(.a(N5225), .b(N5163), .O(gate1619inter2));
  inv1  gate3787(.a(s_302), .O(gate1619inter3));
  inv1  gate3788(.a(s_303), .O(gate1619inter4));
  nand2 gate3789(.a(gate1619inter4), .b(gate1619inter3), .O(gate1619inter5));
  nor2  gate3790(.a(gate1619inter5), .b(gate1619inter2), .O(gate1619inter6));
  inv1  gate3791(.a(N5163), .O(gate1619inter7));
  inv1  gate3792(.a(N5225), .O(gate1619inter8));
  nand2 gate3793(.a(gate1619inter8), .b(gate1619inter7), .O(gate1619inter9));
  nand2 gate3794(.a(s_303), .b(gate1619inter3), .O(gate1619inter10));
  nor2  gate3795(.a(gate1619inter10), .b(gate1619inter9), .O(gate1619inter11));
  nor2  gate3796(.a(gate1619inter11), .b(gate1619inter6), .O(gate1619inter12));
  nand2 gate3797(.a(gate1619inter12), .b(gate1619inter1), .O(N5243));

  xor2  gate4190(.a(N5233), .b(N5174), .O(gate1620inter0));
  nand2 gate4191(.a(gate1620inter0), .b(s_360), .O(gate1620inter1));
  and2  gate4192(.a(N5233), .b(N5174), .O(gate1620inter2));
  inv1  gate4193(.a(s_360), .O(gate1620inter3));
  inv1  gate4194(.a(s_361), .O(gate1620inter4));
  nand2 gate4195(.a(gate1620inter4), .b(gate1620inter3), .O(gate1620inter5));
  nor2  gate4196(.a(gate1620inter5), .b(gate1620inter2), .O(gate1620inter6));
  inv1  gate4197(.a(N5174), .O(gate1620inter7));
  inv1  gate4198(.a(N5233), .O(gate1620inter8));
  nand2 gate4199(.a(gate1620inter8), .b(gate1620inter7), .O(gate1620inter9));
  nand2 gate4200(.a(s_361), .b(gate1620inter3), .O(gate1620inter10));
  nor2  gate4201(.a(gate1620inter10), .b(gate1620inter9), .O(gate1620inter11));
  nor2  gate4202(.a(gate1620inter11), .b(gate1620inter6), .O(gate1620inter12));
  nand2 gate4203(.a(gate1620inter12), .b(gate1620inter1), .O(N5245));
nand2 gate1621( .a(N5177), .b(N5235), .O(N5246) );
inv1 gate1622( .a(N5240), .O(N5250) );
inv1 gate1623( .a(N5228), .O(N5253) );

  xor2  gate3560(.a(N5223), .b(N5242), .O(gate1624inter0));
  nand2 gate3561(.a(gate1624inter0), .b(s_270), .O(gate1624inter1));
  and2  gate3562(.a(N5223), .b(N5242), .O(gate1624inter2));
  inv1  gate3563(.a(s_270), .O(gate1624inter3));
  inv1  gate3564(.a(s_271), .O(gate1624inter4));
  nand2 gate3565(.a(gate1624inter4), .b(gate1624inter3), .O(gate1624inter5));
  nor2  gate3566(.a(gate1624inter5), .b(gate1624inter2), .O(gate1624inter6));
  inv1  gate3567(.a(N5242), .O(gate1624inter7));
  inv1  gate3568(.a(N5223), .O(gate1624inter8));
  nand2 gate3569(.a(gate1624inter8), .b(gate1624inter7), .O(gate1624inter9));
  nand2 gate3570(.a(s_271), .b(gate1624inter3), .O(gate1624inter10));
  nor2  gate3571(.a(gate1624inter10), .b(gate1624inter9), .O(gate1624inter11));
  nor2  gate3572(.a(gate1624inter11), .b(gate1624inter6), .O(gate1624inter12));
  nand2 gate3573(.a(gate1624inter12), .b(gate1624inter1), .O(N5254));

  xor2  gate3140(.a(N5224), .b(N5243), .O(gate1625inter0));
  nand2 gate3141(.a(gate1625inter0), .b(s_210), .O(gate1625inter1));
  and2  gate3142(.a(N5224), .b(N5243), .O(gate1625inter2));
  inv1  gate3143(.a(s_210), .O(gate1625inter3));
  inv1  gate3144(.a(s_211), .O(gate1625inter4));
  nand2 gate3145(.a(gate1625inter4), .b(gate1625inter3), .O(gate1625inter5));
  nor2  gate3146(.a(gate1625inter5), .b(gate1625inter2), .O(gate1625inter6));
  inv1  gate3147(.a(N5243), .O(gate1625inter7));
  inv1  gate3148(.a(N5224), .O(gate1625inter8));
  nand2 gate3149(.a(gate1625inter8), .b(gate1625inter7), .O(gate1625inter9));
  nand2 gate3150(.a(s_211), .b(gate1625inter3), .O(gate1625inter10));
  nor2  gate3151(.a(gate1625inter10), .b(gate1625inter9), .O(gate1625inter11));
  nor2  gate3152(.a(gate1625inter11), .b(gate1625inter6), .O(gate1625inter12));
  nand2 gate3153(.a(gate1625inter12), .b(gate1625inter1), .O(N5257));

  xor2  gate1880(.a(N5245), .b(N5232), .O(gate1626inter0));
  nand2 gate1881(.a(gate1626inter0), .b(s_30), .O(gate1626inter1));
  and2  gate1882(.a(N5245), .b(N5232), .O(gate1626inter2));
  inv1  gate1883(.a(s_30), .O(gate1626inter3));
  inv1  gate1884(.a(s_31), .O(gate1626inter4));
  nand2 gate1885(.a(gate1626inter4), .b(gate1626inter3), .O(gate1626inter5));
  nor2  gate1886(.a(gate1626inter5), .b(gate1626inter2), .O(gate1626inter6));
  inv1  gate1887(.a(N5232), .O(gate1626inter7));
  inv1  gate1888(.a(N5245), .O(gate1626inter8));
  nand2 gate1889(.a(gate1626inter8), .b(gate1626inter7), .O(gate1626inter9));
  nand2 gate1890(.a(s_31), .b(gate1626inter3), .O(gate1626inter10));
  nor2  gate1891(.a(gate1626inter10), .b(gate1626inter9), .O(gate1626inter11));
  nor2  gate1892(.a(gate1626inter11), .b(gate1626inter6), .O(gate1626inter12));
  nand2 gate1893(.a(gate1626inter12), .b(gate1626inter1), .O(N5258));

  xor2  gate2216(.a(N5246), .b(N5234), .O(gate1627inter0));
  nand2 gate2217(.a(gate1627inter0), .b(s_78), .O(gate1627inter1));
  and2  gate2218(.a(N5246), .b(N5234), .O(gate1627inter2));
  inv1  gate2219(.a(s_78), .O(gate1627inter3));
  inv1  gate2220(.a(s_79), .O(gate1627inter4));
  nand2 gate2221(.a(gate1627inter4), .b(gate1627inter3), .O(gate1627inter5));
  nor2  gate2222(.a(gate1627inter5), .b(gate1627inter2), .O(gate1627inter6));
  inv1  gate2223(.a(N5234), .O(gate1627inter7));
  inv1  gate2224(.a(N5246), .O(gate1627inter8));
  nand2 gate2225(.a(gate1627inter8), .b(gate1627inter7), .O(gate1627inter9));
  nand2 gate2226(.a(s_79), .b(gate1627inter3), .O(gate1627inter10));
  nor2  gate2227(.a(gate1627inter10), .b(gate1627inter9), .O(gate1627inter11));
  nor2  gate2228(.a(gate1627inter11), .b(gate1627inter6), .O(gate1627inter12));
  nand2 gate2229(.a(gate1627inter12), .b(gate1627inter1), .O(N5261));
inv1 gate1628( .a(N5257), .O(N5266) );
buf1 gate1629( .a(N5236), .O(N5269) );
and3 gate1630( .a(N5236), .b(N5254), .c(N2307), .O(N5277) );
and3 gate1631( .a(N5250), .b(N5254), .c(N2310), .O(N5278) );
inv1 gate1632( .a(N5261), .O(N5279) );
inv1 gate1633( .a(N5269), .O(N5283) );
nand2 gate1634( .a(N5269), .b(N5253), .O(N5284) );
and3 gate1635( .a(N5236), .b(N5266), .c(N2310), .O(N5285) );
and3 gate1636( .a(N5250), .b(N5266), .c(N2307), .O(N5286) );
buf1 gate1637( .a(N5258), .O(N5289) );
buf1 gate1638( .a(N5258), .O(N5292) );

  xor2  gate2496(.a(N5283), .b(N5228), .O(gate1639inter0));
  nand2 gate2497(.a(gate1639inter0), .b(s_118), .O(gate1639inter1));
  and2  gate2498(.a(N5283), .b(N5228), .O(gate1639inter2));
  inv1  gate2499(.a(s_118), .O(gate1639inter3));
  inv1  gate2500(.a(s_119), .O(gate1639inter4));
  nand2 gate2501(.a(gate1639inter4), .b(gate1639inter3), .O(gate1639inter5));
  nor2  gate2502(.a(gate1639inter5), .b(gate1639inter2), .O(gate1639inter6));
  inv1  gate2503(.a(N5228), .O(gate1639inter7));
  inv1  gate2504(.a(N5283), .O(gate1639inter8));
  nand2 gate2505(.a(gate1639inter8), .b(gate1639inter7), .O(gate1639inter9));
  nand2 gate2506(.a(s_119), .b(gate1639inter3), .O(gate1639inter10));
  nor2  gate2507(.a(gate1639inter10), .b(gate1639inter9), .O(gate1639inter11));
  nor2  gate2508(.a(gate1639inter11), .b(gate1639inter6), .O(gate1639inter12));
  nand2 gate2509(.a(gate1639inter12), .b(gate1639inter1), .O(N5295));
or4 gate1640( .a(N5277), .b(N5285), .c(N5278), .d(N5286), .O(N5298) );
buf1 gate1641( .a(N5279), .O(N5303) );
buf1 gate1642( .a(N5279), .O(N5306) );

  xor2  gate4134(.a(N5284), .b(N5295), .O(gate1643inter0));
  nand2 gate4135(.a(gate1643inter0), .b(s_352), .O(gate1643inter1));
  and2  gate4136(.a(N5284), .b(N5295), .O(gate1643inter2));
  inv1  gate4137(.a(s_352), .O(gate1643inter3));
  inv1  gate4138(.a(s_353), .O(gate1643inter4));
  nand2 gate4139(.a(gate1643inter4), .b(gate1643inter3), .O(gate1643inter5));
  nor2  gate4140(.a(gate1643inter5), .b(gate1643inter2), .O(gate1643inter6));
  inv1  gate4141(.a(N5295), .O(gate1643inter7));
  inv1  gate4142(.a(N5284), .O(gate1643inter8));
  nand2 gate4143(.a(gate1643inter8), .b(gate1643inter7), .O(gate1643inter9));
  nand2 gate4144(.a(s_353), .b(gate1643inter3), .O(gate1643inter10));
  nor2  gate4145(.a(gate1643inter10), .b(gate1643inter9), .O(gate1643inter11));
  nor2  gate4146(.a(gate1643inter11), .b(gate1643inter6), .O(gate1643inter12));
  nand2 gate4147(.a(gate1643inter12), .b(gate1643inter1), .O(N5309));
inv1 gate1644( .a(N5292), .O(N5312) );
inv1 gate1645( .a(N5289), .O(N5313) );
inv1 gate1646( .a(N5306), .O(N5322) );
inv1 gate1647( .a(N5303), .O(N5323) );
buf1 gate1648( .a(N5298), .O(N5324) );
buf1 gate1649( .a(N5298), .O(N5327) );
buf1 gate1650( .a(N5309), .O(N5332) );
buf1 gate1651( .a(N5309), .O(N5335) );
nand2 gate1652( .a(N5324), .b(N5323), .O(N5340) );

  xor2  gate1978(.a(N5322), .b(N5327), .O(gate1653inter0));
  nand2 gate1979(.a(gate1653inter0), .b(s_44), .O(gate1653inter1));
  and2  gate1980(.a(N5322), .b(N5327), .O(gate1653inter2));
  inv1  gate1981(.a(s_44), .O(gate1653inter3));
  inv1  gate1982(.a(s_45), .O(gate1653inter4));
  nand2 gate1983(.a(gate1653inter4), .b(gate1653inter3), .O(gate1653inter5));
  nor2  gate1984(.a(gate1653inter5), .b(gate1653inter2), .O(gate1653inter6));
  inv1  gate1985(.a(N5327), .O(gate1653inter7));
  inv1  gate1986(.a(N5322), .O(gate1653inter8));
  nand2 gate1987(.a(gate1653inter8), .b(gate1653inter7), .O(gate1653inter9));
  nand2 gate1988(.a(s_45), .b(gate1653inter3), .O(gate1653inter10));
  nor2  gate1989(.a(gate1653inter10), .b(gate1653inter9), .O(gate1653inter11));
  nor2  gate1990(.a(gate1653inter11), .b(gate1653inter6), .O(gate1653inter12));
  nand2 gate1991(.a(gate1653inter12), .b(gate1653inter1), .O(N5341));
inv1 gate1654( .a(N5327), .O(N5344) );
inv1 gate1655( .a(N5324), .O(N5345) );

  xor2  gate3154(.a(N5313), .b(N5332), .O(gate1656inter0));
  nand2 gate3155(.a(gate1656inter0), .b(s_212), .O(gate1656inter1));
  and2  gate3156(.a(N5313), .b(N5332), .O(gate1656inter2));
  inv1  gate3157(.a(s_212), .O(gate1656inter3));
  inv1  gate3158(.a(s_213), .O(gate1656inter4));
  nand2 gate3159(.a(gate1656inter4), .b(gate1656inter3), .O(gate1656inter5));
  nor2  gate3160(.a(gate1656inter5), .b(gate1656inter2), .O(gate1656inter6));
  inv1  gate3161(.a(N5332), .O(gate1656inter7));
  inv1  gate3162(.a(N5313), .O(gate1656inter8));
  nand2 gate3163(.a(gate1656inter8), .b(gate1656inter7), .O(gate1656inter9));
  nand2 gate3164(.a(s_213), .b(gate1656inter3), .O(gate1656inter10));
  nor2  gate3165(.a(gate1656inter10), .b(gate1656inter9), .O(gate1656inter11));
  nor2  gate3166(.a(gate1656inter11), .b(gate1656inter6), .O(gate1656inter12));
  nand2 gate3167(.a(gate1656inter12), .b(gate1656inter1), .O(N5348));

  xor2  gate3812(.a(N5312), .b(N5335), .O(gate1657inter0));
  nand2 gate3813(.a(gate1657inter0), .b(s_306), .O(gate1657inter1));
  and2  gate3814(.a(N5312), .b(N5335), .O(gate1657inter2));
  inv1  gate3815(.a(s_306), .O(gate1657inter3));
  inv1  gate3816(.a(s_307), .O(gate1657inter4));
  nand2 gate3817(.a(gate1657inter4), .b(gate1657inter3), .O(gate1657inter5));
  nor2  gate3818(.a(gate1657inter5), .b(gate1657inter2), .O(gate1657inter6));
  inv1  gate3819(.a(N5335), .O(gate1657inter7));
  inv1  gate3820(.a(N5312), .O(gate1657inter8));
  nand2 gate3821(.a(gate1657inter8), .b(gate1657inter7), .O(gate1657inter9));
  nand2 gate3822(.a(s_307), .b(gate1657inter3), .O(gate1657inter10));
  nor2  gate3823(.a(gate1657inter10), .b(gate1657inter9), .O(gate1657inter11));
  nor2  gate3824(.a(gate1657inter11), .b(gate1657inter6), .O(gate1657inter12));
  nand2 gate3825(.a(gate1657inter12), .b(gate1657inter1), .O(N5349));

  xor2  gate3630(.a(N5345), .b(N5303), .O(gate1658inter0));
  nand2 gate3631(.a(gate1658inter0), .b(s_280), .O(gate1658inter1));
  and2  gate3632(.a(N5345), .b(N5303), .O(gate1658inter2));
  inv1  gate3633(.a(s_280), .O(gate1658inter3));
  inv1  gate3634(.a(s_281), .O(gate1658inter4));
  nand2 gate3635(.a(gate1658inter4), .b(gate1658inter3), .O(gate1658inter5));
  nor2  gate3636(.a(gate1658inter5), .b(gate1658inter2), .O(gate1658inter6));
  inv1  gate3637(.a(N5303), .O(gate1658inter7));
  inv1  gate3638(.a(N5345), .O(gate1658inter8));
  nand2 gate3639(.a(gate1658inter8), .b(gate1658inter7), .O(gate1658inter9));
  nand2 gate3640(.a(s_281), .b(gate1658inter3), .O(gate1658inter10));
  nor2  gate3641(.a(gate1658inter10), .b(gate1658inter9), .O(gate1658inter11));
  nor2  gate3642(.a(gate1658inter11), .b(gate1658inter6), .O(gate1658inter12));
  nand2 gate3643(.a(gate1658inter12), .b(gate1658inter1), .O(N5350));
nand2 gate1659( .a(N5306), .b(N5344), .O(N5351) );
inv1 gate1660( .a(N5335), .O(N5352) );
inv1 gate1661( .a(N5332), .O(N5353) );

  xor2  gate3980(.a(N5353), .b(N5289), .O(gate1662inter0));
  nand2 gate3981(.a(gate1662inter0), .b(s_330), .O(gate1662inter1));
  and2  gate3982(.a(N5353), .b(N5289), .O(gate1662inter2));
  inv1  gate3983(.a(s_330), .O(gate1662inter3));
  inv1  gate3984(.a(s_331), .O(gate1662inter4));
  nand2 gate3985(.a(gate1662inter4), .b(gate1662inter3), .O(gate1662inter5));
  nor2  gate3986(.a(gate1662inter5), .b(gate1662inter2), .O(gate1662inter6));
  inv1  gate3987(.a(N5289), .O(gate1662inter7));
  inv1  gate3988(.a(N5353), .O(gate1662inter8));
  nand2 gate3989(.a(gate1662inter8), .b(gate1662inter7), .O(gate1662inter9));
  nand2 gate3990(.a(s_331), .b(gate1662inter3), .O(gate1662inter10));
  nor2  gate3991(.a(gate1662inter10), .b(gate1662inter9), .O(gate1662inter11));
  nor2  gate3992(.a(gate1662inter11), .b(gate1662inter6), .O(gate1662inter12));
  nand2 gate3993(.a(gate1662inter12), .b(gate1662inter1), .O(N5354));

  xor2  gate3938(.a(N5352), .b(N5292), .O(gate1663inter0));
  nand2 gate3939(.a(gate1663inter0), .b(s_324), .O(gate1663inter1));
  and2  gate3940(.a(N5352), .b(N5292), .O(gate1663inter2));
  inv1  gate3941(.a(s_324), .O(gate1663inter3));
  inv1  gate3942(.a(s_325), .O(gate1663inter4));
  nand2 gate3943(.a(gate1663inter4), .b(gate1663inter3), .O(gate1663inter5));
  nor2  gate3944(.a(gate1663inter5), .b(gate1663inter2), .O(gate1663inter6));
  inv1  gate3945(.a(N5292), .O(gate1663inter7));
  inv1  gate3946(.a(N5352), .O(gate1663inter8));
  nand2 gate3947(.a(gate1663inter8), .b(gate1663inter7), .O(gate1663inter9));
  nand2 gate3948(.a(s_325), .b(gate1663inter3), .O(gate1663inter10));
  nor2  gate3949(.a(gate1663inter10), .b(gate1663inter9), .O(gate1663inter11));
  nor2  gate3950(.a(gate1663inter11), .b(gate1663inter6), .O(gate1663inter12));
  nand2 gate3951(.a(gate1663inter12), .b(gate1663inter1), .O(N5355));
nand2 gate1664( .a(N5350), .b(N5340), .O(N5356) );

  xor2  gate2986(.a(N5341), .b(N5351), .O(gate1665inter0));
  nand2 gate2987(.a(gate1665inter0), .b(s_188), .O(gate1665inter1));
  and2  gate2988(.a(N5341), .b(N5351), .O(gate1665inter2));
  inv1  gate2989(.a(s_188), .O(gate1665inter3));
  inv1  gate2990(.a(s_189), .O(gate1665inter4));
  nand2 gate2991(.a(gate1665inter4), .b(gate1665inter3), .O(gate1665inter5));
  nor2  gate2992(.a(gate1665inter5), .b(gate1665inter2), .O(gate1665inter6));
  inv1  gate2993(.a(N5351), .O(gate1665inter7));
  inv1  gate2994(.a(N5341), .O(gate1665inter8));
  nand2 gate2995(.a(gate1665inter8), .b(gate1665inter7), .O(gate1665inter9));
  nand2 gate2996(.a(s_189), .b(gate1665inter3), .O(gate1665inter10));
  nor2  gate2997(.a(gate1665inter10), .b(gate1665inter9), .O(gate1665inter11));
  nor2  gate2998(.a(gate1665inter11), .b(gate1665inter6), .O(gate1665inter12));
  nand2 gate2999(.a(gate1665inter12), .b(gate1665inter1), .O(N5357));

  xor2  gate3238(.a(N5354), .b(N5348), .O(gate1666inter0));
  nand2 gate3239(.a(gate1666inter0), .b(s_224), .O(gate1666inter1));
  and2  gate3240(.a(N5354), .b(N5348), .O(gate1666inter2));
  inv1  gate3241(.a(s_224), .O(gate1666inter3));
  inv1  gate3242(.a(s_225), .O(gate1666inter4));
  nand2 gate3243(.a(gate1666inter4), .b(gate1666inter3), .O(gate1666inter5));
  nor2  gate3244(.a(gate1666inter5), .b(gate1666inter2), .O(gate1666inter6));
  inv1  gate3245(.a(N5348), .O(gate1666inter7));
  inv1  gate3246(.a(N5354), .O(gate1666inter8));
  nand2 gate3247(.a(gate1666inter8), .b(gate1666inter7), .O(gate1666inter9));
  nand2 gate3248(.a(s_225), .b(gate1666inter3), .O(gate1666inter10));
  nor2  gate3249(.a(gate1666inter10), .b(gate1666inter9), .O(gate1666inter11));
  nor2  gate3250(.a(gate1666inter11), .b(gate1666inter6), .O(gate1666inter12));
  nand2 gate3251(.a(gate1666inter12), .b(gate1666inter1), .O(N5358));
nand2 gate1667( .a(N5349), .b(N5355), .O(N5359) );
and2 gate1668( .a(N5356), .b(N5357), .O(N5360) );
nand2 gate1669( .a(N5358), .b(N5359), .O(N5361) );

endmodule