module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);

input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;//RE__PI;

input s_0,s_1;//RE__ALLOW(00,01,10,11);
input s_2,s_3;//RE__ALLOW(00,01,10,11);
input s_4,s_5;//RE__ALLOW(00,01,10,11);
input s_6,s_7;//RE__ALLOW(00,01,10,11);
input s_8,s_9;//RE__ALLOW(00,01,10,11);
input s_10,s_11;//RE__ALLOW(00,01,10,11);
input s_12,s_13;//RE__ALLOW(00,01,10,11);
input s_14,s_15;//RE__ALLOW(00,01,10,11);
input s_16,s_17;//RE__ALLOW(00,01,10,11);
input s_18,s_19;//RE__ALLOW(00,01,10,11);
input s_20,s_21;//RE__ALLOW(00,01,10,11);
input s_22,s_23;//RE__ALLOW(00,01,10,11);
input s_24,s_25;//RE__ALLOW(00,01,10,11);
input s_26,s_27;//RE__ALLOW(00,01,10,11);
input s_28,s_29;//RE__ALLOW(00,01,10,11);
input s_30,s_31;//RE__ALLOW(00,01,10,11);
input s_32,s_33;//RE__ALLOW(00,01,10,11);
input s_34,s_35;//RE__ALLOW(00,01,10,11);
input s_36,s_37;//RE__ALLOW(00,01,10,11);
input s_38,s_39;//RE__ALLOW(00,01,10,11);
input s_40,s_41;//RE__ALLOW(00,01,10,11);
input s_42,s_43;//RE__ALLOW(00,01,10,11);
input s_44,s_45;//RE__ALLOW(00,01,10,11);
input s_46,s_47;//RE__ALLOW(00,01,10,11);
input s_48,s_49;//RE__ALLOW(00,01,10,11);
input s_50,s_51;//RE__ALLOW(00,01,10,11);
input s_52,s_53;//RE__ALLOW(00,01,10,11);
input s_54,s_55;//RE__ALLOW(00,01,10,11);
input s_56,s_57;//RE__ALLOW(00,01,10,11);
input s_58,s_59;//RE__ALLOW(00,01,10,11);
input s_60,s_61;//RE__ALLOW(00,01,10,11);
input s_62,s_63;//RE__ALLOW(00,01,10,11);
input s_64,s_65;//RE__ALLOW(00,01,10,11);
input s_66,s_67;//RE__ALLOW(00,01,10,11);
input s_68,s_69;//RE__ALLOW(00,01,10,11);
input s_70,s_71;//RE__ALLOW(00,01,10,11);
input s_72,s_73;//RE__ALLOW(00,01,10,11);
input s_74,s_75;//RE__ALLOW(00,01,10,11);
input s_76,s_77;//RE__ALLOW(00,01,10,11);
input s_78,s_79;//RE__ALLOW(00,01,10,11);
input s_80,s_81;//RE__ALLOW(00,01,10,11);
input s_82,s_83;//RE__ALLOW(00,01,10,11);
input s_84,s_85;//RE__ALLOW(00,01,10,11);
input s_86,s_87;//RE__ALLOW(00,01,10,11);
input s_88,s_89;//RE__ALLOW(00,01,10,11);
input s_90,s_91;//RE__ALLOW(00,01,10,11);
input s_92,s_93;//RE__ALLOW(00,01,10,11);
input s_94,s_95;//RE__ALLOW(00,01,10,11);
input s_96,s_97;//RE__ALLOW(00,01,10,11);
input s_98,s_99;//RE__ALLOW(00,01,10,11);
input s_100,s_101;//RE__ALLOW(00,01,10,11);
input s_102,s_103;//RE__ALLOW(00,01,10,11);
input s_104,s_105;//RE__ALLOW(00,01,10,11);
input s_106,s_107;//RE__ALLOW(00,01,10,11);
input s_108,s_109;//RE__ALLOW(00,01,10,11);
input s_110,s_111;//RE__ALLOW(00,01,10,11);
input s_112,s_113;//RE__ALLOW(00,01,10,11);
input s_114,s_115;//RE__ALLOW(00,01,10,11);
input s_116,s_117;//RE__ALLOW(00,01,10,11);
input s_118,s_119;//RE__ALLOW(00,01,10,11);
input s_120,s_121;//RE__ALLOW(00,01,10,11);
input s_122,s_123;//RE__ALLOW(00,01,10,11);
input s_124,s_125;//RE__ALLOW(00,01,10,11);
input s_126,s_127;//RE__ALLOW(00,01,10,11);
input s_128,s_129;//RE__ALLOW(00,01,10,11);
input s_130,s_131;//RE__ALLOW(00,01,10,11);
input s_132,s_133;//RE__ALLOW(00,01,10,11);
input s_134,s_135;//RE__ALLOW(00,01,10,11);
input s_136,s_137;//RE__ALLOW(00,01,10,11);
input s_138,s_139;//RE__ALLOW(00,01,10,11);
input s_140,s_141;//RE__ALLOW(00,01,10,11);
input s_142,s_143;//RE__ALLOW(00,01,10,11);
input s_144,s_145;//RE__ALLOW(00,01,10,11);
input s_146,s_147;//RE__ALLOW(00,01,10,11);
input s_148,s_149;//RE__ALLOW(00,01,10,11);
input s_150,s_151;//RE__ALLOW(00,01,10,11);
input s_152,s_153;//RE__ALLOW(00,01,10,11);
input s_154,s_155;//RE__ALLOW(00,01,10,11);
input s_156,s_157;//RE__ALLOW(00,01,10,11);
input s_158,s_159;//RE__ALLOW(00,01,10,11);
input s_160,s_161;//RE__ALLOW(00,01,10,11);
input s_162,s_163;//RE__ALLOW(00,01,10,11);
input s_164,s_165;//RE__ALLOW(00,01,10,11);
input s_166,s_167;//RE__ALLOW(00,01,10,11);
input s_168,s_169;//RE__ALLOW(00,01,10,11);
input s_170,s_171;//RE__ALLOW(00,01,10,11);
input s_172,s_173;//RE__ALLOW(00,01,10,11);
input s_174,s_175;//RE__ALLOW(00,01,10,11);
input s_176,s_177;//RE__ALLOW(00,01,10,11);
input s_178,s_179;//RE__ALLOW(00,01,10,11);
input s_180,s_181;//RE__ALLOW(00,01,10,11);
input s_182,s_183;//RE__ALLOW(00,01,10,11);
input s_184,s_185;//RE__ALLOW(00,01,10,11);
input s_186,s_187;//RE__ALLOW(00,01,10,11);
input s_188,s_189;//RE__ALLOW(00,01,10,11);
input s_190,s_191;//RE__ALLOW(00,01,10,11);
input s_192,s_193;//RE__ALLOW(00,01,10,11);
input s_194,s_195;//RE__ALLOW(00,01,10,11);
input s_196,s_197;//RE__ALLOW(00,01,10,11);
input s_198,s_199;//RE__ALLOW(00,01,10,11);
input s_200,s_201;//RE__ALLOW(00,01,10,11);
input s_202,s_203;//RE__ALLOW(00,01,10,11);
input s_204,s_205;//RE__ALLOW(00,01,10,11);
input s_206,s_207;//RE__ALLOW(00,01,10,11);
input s_208,s_209;//RE__ALLOW(00,01,10,11);
input s_210,s_211;//RE__ALLOW(00,01,10,11);
input s_212,s_213;//RE__ALLOW(00,01,10,11);
input s_214,s_215;//RE__ALLOW(00,01,10,11);
input s_216,s_217;//RE__ALLOW(00,01,10,11);
input s_218,s_219;//RE__ALLOW(00,01,10,11);
input s_220,s_221;//RE__ALLOW(00,01,10,11);
input s_222,s_223;//RE__ALLOW(00,01,10,11);
input s_224,s_225;//RE__ALLOW(00,01,10,11);
input s_226,s_227;//RE__ALLOW(00,01,10,11);
input s_228,s_229;//RE__ALLOW(00,01,10,11);
input s_230,s_231;//RE__ALLOW(00,01,10,11);
input s_232,s_233;//RE__ALLOW(00,01,10,11);
input s_234,s_235;//RE__ALLOW(00,01,10,11);
input s_236,s_237;//RE__ALLOW(00,01,10,11);
input s_238,s_239;//RE__ALLOW(00,01,10,11);
input s_240,s_241;//RE__ALLOW(00,01,10,11);
input s_242,s_243;//RE__ALLOW(00,01,10,11);
input s_244,s_245;//RE__ALLOW(00,01,10,11);
input s_246,s_247;//RE__ALLOW(00,01,10,11);
input s_248,s_249;//RE__ALLOW(00,01,10,11);
input s_250,s_251;//RE__ALLOW(00,01,10,11);
input s_252,s_253;//RE__ALLOW(00,01,10,11);
input s_254,s_255;//RE__ALLOW(00,01,10,11);
input s_256,s_257;//RE__ALLOW(00,01,10,11);
input s_258,s_259;//RE__ALLOW(00,01,10,11);
input s_260,s_261;//RE__ALLOW(00,01,10,11);
input s_262,s_263;//RE__ALLOW(00,01,10,11);
input s_264,s_265;//RE__ALLOW(00,01,10,11);
input s_266,s_267;//RE__ALLOW(00,01,10,11);
input s_268,s_269;//RE__ALLOW(00,01,10,11);
input s_270,s_271;//RE__ALLOW(00,01,10,11);
input s_272,s_273;//RE__ALLOW(00,01,10,11);
input s_274,s_275;//RE__ALLOW(00,01,10,11);
input s_276,s_277;//RE__ALLOW(00,01,10,11);
input s_278,s_279;//RE__ALLOW(00,01,10,11);
input s_280,s_281;//RE__ALLOW(00,01,10,11);
input s_282,s_283;//RE__ALLOW(00,01,10,11);
input s_284,s_285;//RE__ALLOW(00,01,10,11);
input s_286,s_287;//RE__ALLOW(00,01,10,11);
input s_288,s_289;//RE__ALLOW(00,01,10,11);
input s_290,s_291;//RE__ALLOW(00,01,10,11);
input s_292,s_293;//RE__ALLOW(00,01,10,11);
input s_294,s_295;//RE__ALLOW(00,01,10,11);
input s_296,s_297;//RE__ALLOW(00,01,10,11);
input s_298,s_299;//RE__ALLOW(00,01,10,11);
input s_300,s_301;//RE__ALLOW(00,01,10,11);
input s_302,s_303;//RE__ALLOW(00,01,10,11);
input s_304,s_305;//RE__ALLOW(00,01,10,11);
input s_306,s_307;//RE__ALLOW(00,01,10,11);
input s_308,s_309;//RE__ALLOW(00,01,10,11);
input s_310,s_311;//RE__ALLOW(00,01,10,11);
input s_312,s_313;//RE__ALLOW(00,01,10,11);
input s_314,s_315;//RE__ALLOW(00,01,10,11);
input s_316,s_317;//RE__ALLOW(00,01,10,11);
input s_318,s_319;//RE__ALLOW(00,01,10,11);
input s_320,s_321;//RE__ALLOW(00,01,10,11);
input s_322,s_323;//RE__ALLOW(00,01,10,11);
input s_324,s_325;//RE__ALLOW(00,01,10,11);
input s_326,s_327;//RE__ALLOW(00,01,10,11);
input s_328,s_329;//RE__ALLOW(00,01,10,11);
input s_330,s_331;//RE__ALLOW(00,01,10,11);
input s_332,s_333;//RE__ALLOW(00,01,10,11);
input s_334,s_335;//RE__ALLOW(00,01,10,11);
input s_336,s_337;//RE__ALLOW(00,01,10,11);
input s_338,s_339;//RE__ALLOW(00,01,10,11);
input s_340,s_341;//RE__ALLOW(00,01,10,11);
input s_342,s_343;//RE__ALLOW(00,01,10,11);
input s_344,s_345;//RE__ALLOW(00,01,10,11);
input s_346,s_347;//RE__ALLOW(00,01,10,11);
input s_348,s_349;//RE__ALLOW(00,01,10,11);
input s_350,s_351;//RE__ALLOW(00,01,10,11);
input s_352,s_353;//RE__ALLOW(00,01,10,11);
input s_354,s_355;//RE__ALLOW(00,01,10,11);
input s_356,s_357;//RE__ALLOW(00,01,10,11);
input s_358,s_359;//RE__ALLOW(00,01,10,11);
input s_360,s_361;//RE__ALLOW(00,01,10,11);
input s_362,s_363;//RE__ALLOW(00,01,10,11);
input s_364,s_365;//RE__ALLOW(00,01,10,11);
input s_366,s_367;//RE__ALLOW(00,01,10,11);
input s_368,s_369;//RE__ALLOW(00,01,10,11);
input s_370,s_371;//RE__ALLOW(00,01,10,11);
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;

  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate211inter0, gate211inter1, gate211inter2, gate211inter3, gate211inter4, gate211inter5, gate211inter6, gate211inter7, gate211inter8, gate211inter9, gate211inter10, gate211inter11, gate211inter12, gate100inter0, gate100inter1, gate100inter2, gate100inter3, gate100inter4, gate100inter5, gate100inter6, gate100inter7, gate100inter8, gate100inter9, gate100inter10, gate100inter11, gate100inter12, gate86inter0, gate86inter1, gate86inter2, gate86inter3, gate86inter4, gate86inter5, gate86inter6, gate86inter7, gate86inter8, gate86inter9, gate86inter10, gate86inter11, gate86inter12, gate435inter0, gate435inter1, gate435inter2, gate435inter3, gate435inter4, gate435inter5, gate435inter6, gate435inter7, gate435inter8, gate435inter9, gate435inter10, gate435inter11, gate435inter12, gate405inter0, gate405inter1, gate405inter2, gate405inter3, gate405inter4, gate405inter5, gate405inter6, gate405inter7, gate405inter8, gate405inter9, gate405inter10, gate405inter11, gate405inter12, gate489inter0, gate489inter1, gate489inter2, gate489inter3, gate489inter4, gate489inter5, gate489inter6, gate489inter7, gate489inter8, gate489inter9, gate489inter10, gate489inter11, gate489inter12, gate165inter0, gate165inter1, gate165inter2, gate165inter3, gate165inter4, gate165inter5, gate165inter6, gate165inter7, gate165inter8, gate165inter9, gate165inter10, gate165inter11, gate165inter12, gate286inter0, gate286inter1, gate286inter2, gate286inter3, gate286inter4, gate286inter5, gate286inter6, gate286inter7, gate286inter8, gate286inter9, gate286inter10, gate286inter11, gate286inter12, gate112inter0, gate112inter1, gate112inter2, gate112inter3, gate112inter4, gate112inter5, gate112inter6, gate112inter7, gate112inter8, gate112inter9, gate112inter10, gate112inter11, gate112inter12, gate79inter0, gate79inter1, gate79inter2, gate79inter3, gate79inter4, gate79inter5, gate79inter6, gate79inter7, gate79inter8, gate79inter9, gate79inter10, gate79inter11, gate79inter12, gate284inter0, gate284inter1, gate284inter2, gate284inter3, gate284inter4, gate284inter5, gate284inter6, gate284inter7, gate284inter8, gate284inter9, gate284inter10, gate284inter11, gate284inter12, gate38inter0, gate38inter1, gate38inter2, gate38inter3, gate38inter4, gate38inter5, gate38inter6, gate38inter7, gate38inter8, gate38inter9, gate38inter10, gate38inter11, gate38inter12, gate406inter0, gate406inter1, gate406inter2, gate406inter3, gate406inter4, gate406inter5, gate406inter6, gate406inter7, gate406inter8, gate406inter9, gate406inter10, gate406inter11, gate406inter12, gate294inter0, gate294inter1, gate294inter2, gate294inter3, gate294inter4, gate294inter5, gate294inter6, gate294inter7, gate294inter8, gate294inter9, gate294inter10, gate294inter11, gate294inter12, gate136inter0, gate136inter1, gate136inter2, gate136inter3, gate136inter4, gate136inter5, gate136inter6, gate136inter7, gate136inter8, gate136inter9, gate136inter10, gate136inter11, gate136inter12, gate30inter0, gate30inter1, gate30inter2, gate30inter3, gate30inter4, gate30inter5, gate30inter6, gate30inter7, gate30inter8, gate30inter9, gate30inter10, gate30inter11, gate30inter12, gate222inter0, gate222inter1, gate222inter2, gate222inter3, gate222inter4, gate222inter5, gate222inter6, gate222inter7, gate222inter8, gate222inter9, gate222inter10, gate222inter11, gate222inter12, gate271inter0, gate271inter1, gate271inter2, gate271inter3, gate271inter4, gate271inter5, gate271inter6, gate271inter7, gate271inter8, gate271inter9, gate271inter10, gate271inter11, gate271inter12, gate119inter0, gate119inter1, gate119inter2, gate119inter3, gate119inter4, gate119inter5, gate119inter6, gate119inter7, gate119inter8, gate119inter9, gate119inter10, gate119inter11, gate119inter12, gate400inter0, gate400inter1, gate400inter2, gate400inter3, gate400inter4, gate400inter5, gate400inter6, gate400inter7, gate400inter8, gate400inter9, gate400inter10, gate400inter11, gate400inter12, gate508inter0, gate508inter1, gate508inter2, gate508inter3, gate508inter4, gate508inter5, gate508inter6, gate508inter7, gate508inter8, gate508inter9, gate508inter10, gate508inter11, gate508inter12, gate502inter0, gate502inter1, gate502inter2, gate502inter3, gate502inter4, gate502inter5, gate502inter6, gate502inter7, gate502inter8, gate502inter9, gate502inter10, gate502inter11, gate502inter12, gate266inter0, gate266inter1, gate266inter2, gate266inter3, gate266inter4, gate266inter5, gate266inter6, gate266inter7, gate266inter8, gate266inter9, gate266inter10, gate266inter11, gate266inter12, gate482inter0, gate482inter1, gate482inter2, gate482inter3, gate482inter4, gate482inter5, gate482inter6, gate482inter7, gate482inter8, gate482inter9, gate482inter10, gate482inter11, gate482inter12, gate110inter0, gate110inter1, gate110inter2, gate110inter3, gate110inter4, gate110inter5, gate110inter6, gate110inter7, gate110inter8, gate110inter9, gate110inter10, gate110inter11, gate110inter12, gate13inter0, gate13inter1, gate13inter2, gate13inter3, gate13inter4, gate13inter5, gate13inter6, gate13inter7, gate13inter8, gate13inter9, gate13inter10, gate13inter11, gate13inter12, gate418inter0, gate418inter1, gate418inter2, gate418inter3, gate418inter4, gate418inter5, gate418inter6, gate418inter7, gate418inter8, gate418inter9, gate418inter10, gate418inter11, gate418inter12, gate433inter0, gate433inter1, gate433inter2, gate433inter3, gate433inter4, gate433inter5, gate433inter6, gate433inter7, gate433inter8, gate433inter9, gate433inter10, gate433inter11, gate433inter12, gate134inter0, gate134inter1, gate134inter2, gate134inter3, gate134inter4, gate134inter5, gate134inter6, gate134inter7, gate134inter8, gate134inter9, gate134inter10, gate134inter11, gate134inter12, gate421inter0, gate421inter1, gate421inter2, gate421inter3, gate421inter4, gate421inter5, gate421inter6, gate421inter7, gate421inter8, gate421inter9, gate421inter10, gate421inter11, gate421inter12, gate214inter0, gate214inter1, gate214inter2, gate214inter3, gate214inter4, gate214inter5, gate214inter6, gate214inter7, gate214inter8, gate214inter9, gate214inter10, gate214inter11, gate214inter12, gate68inter0, gate68inter1, gate68inter2, gate68inter3, gate68inter4, gate68inter5, gate68inter6, gate68inter7, gate68inter8, gate68inter9, gate68inter10, gate68inter11, gate68inter12, gate111inter0, gate111inter1, gate111inter2, gate111inter3, gate111inter4, gate111inter5, gate111inter6, gate111inter7, gate111inter8, gate111inter9, gate111inter10, gate111inter11, gate111inter12, gate94inter0, gate94inter1, gate94inter2, gate94inter3, gate94inter4, gate94inter5, gate94inter6, gate94inter7, gate94inter8, gate94inter9, gate94inter10, gate94inter11, gate94inter12, gate231inter0, gate231inter1, gate231inter2, gate231inter3, gate231inter4, gate231inter5, gate231inter6, gate231inter7, gate231inter8, gate231inter9, gate231inter10, gate231inter11, gate231inter12, gate448inter0, gate448inter1, gate448inter2, gate448inter3, gate448inter4, gate448inter5, gate448inter6, gate448inter7, gate448inter8, gate448inter9, gate448inter10, gate448inter11, gate448inter12, gate487inter0, gate487inter1, gate487inter2, gate487inter3, gate487inter4, gate487inter5, gate487inter6, gate487inter7, gate487inter8, gate487inter9, gate487inter10, gate487inter11, gate487inter12, gate166inter0, gate166inter1, gate166inter2, gate166inter3, gate166inter4, gate166inter5, gate166inter6, gate166inter7, gate166inter8, gate166inter9, gate166inter10, gate166inter11, gate166inter12, gate187inter0, gate187inter1, gate187inter2, gate187inter3, gate187inter4, gate187inter5, gate187inter6, gate187inter7, gate187inter8, gate187inter9, gate187inter10, gate187inter11, gate187inter12, gate51inter0, gate51inter1, gate51inter2, gate51inter3, gate51inter4, gate51inter5, gate51inter6, gate51inter7, gate51inter8, gate51inter9, gate51inter10, gate51inter11, gate51inter12, gate124inter0, gate124inter1, gate124inter2, gate124inter3, gate124inter4, gate124inter5, gate124inter6, gate124inter7, gate124inter8, gate124inter9, gate124inter10, gate124inter11, gate124inter12, gate164inter0, gate164inter1, gate164inter2, gate164inter3, gate164inter4, gate164inter5, gate164inter6, gate164inter7, gate164inter8, gate164inter9, gate164inter10, gate164inter11, gate164inter12, gate99inter0, gate99inter1, gate99inter2, gate99inter3, gate99inter4, gate99inter5, gate99inter6, gate99inter7, gate99inter8, gate99inter9, gate99inter10, gate99inter11, gate99inter12, gate185inter0, gate185inter1, gate185inter2, gate185inter3, gate185inter4, gate185inter5, gate185inter6, gate185inter7, gate185inter8, gate185inter9, gate185inter10, gate185inter11, gate185inter12, gate457inter0, gate457inter1, gate457inter2, gate457inter3, gate457inter4, gate457inter5, gate457inter6, gate457inter7, gate457inter8, gate457inter9, gate457inter10, gate457inter11, gate457inter12, gate275inter0, gate275inter1, gate275inter2, gate275inter3, gate275inter4, gate275inter5, gate275inter6, gate275inter7, gate275inter8, gate275inter9, gate275inter10, gate275inter11, gate275inter12, gate103inter0, gate103inter1, gate103inter2, gate103inter3, gate103inter4, gate103inter5, gate103inter6, gate103inter7, gate103inter8, gate103inter9, gate103inter10, gate103inter11, gate103inter12, gate198inter0, gate198inter1, gate198inter2, gate198inter3, gate198inter4, gate198inter5, gate198inter6, gate198inter7, gate198inter8, gate198inter9, gate198inter10, gate198inter11, gate198inter12, gate408inter0, gate408inter1, gate408inter2, gate408inter3, gate408inter4, gate408inter5, gate408inter6, gate408inter7, gate408inter8, gate408inter9, gate408inter10, gate408inter11, gate408inter12, gate9inter0, gate9inter1, gate9inter2, gate9inter3, gate9inter4, gate9inter5, gate9inter6, gate9inter7, gate9inter8, gate9inter9, gate9inter10, gate9inter11, gate9inter12, gate42inter0, gate42inter1, gate42inter2, gate42inter3, gate42inter4, gate42inter5, gate42inter6, gate42inter7, gate42inter8, gate42inter9, gate42inter10, gate42inter11, gate42inter12, gate92inter0, gate92inter1, gate92inter2, gate92inter3, gate92inter4, gate92inter5, gate92inter6, gate92inter7, gate92inter8, gate92inter9, gate92inter10, gate92inter11, gate92inter12, gate97inter0, gate97inter1, gate97inter2, gate97inter3, gate97inter4, gate97inter5, gate97inter6, gate97inter7, gate97inter8, gate97inter9, gate97inter10, gate97inter11, gate97inter12, gate235inter0, gate235inter1, gate235inter2, gate235inter3, gate235inter4, gate235inter5, gate235inter6, gate235inter7, gate235inter8, gate235inter9, gate235inter10, gate235inter11, gate235inter12, gate497inter0, gate497inter1, gate497inter2, gate497inter3, gate497inter4, gate497inter5, gate497inter6, gate497inter7, gate497inter8, gate497inter9, gate497inter10, gate497inter11, gate497inter12, gate459inter0, gate459inter1, gate459inter2, gate459inter3, gate459inter4, gate459inter5, gate459inter6, gate459inter7, gate459inter8, gate459inter9, gate459inter10, gate459inter11, gate459inter12, gate105inter0, gate105inter1, gate105inter2, gate105inter3, gate105inter4, gate105inter5, gate105inter6, gate105inter7, gate105inter8, gate105inter9, gate105inter10, gate105inter11, gate105inter12, gate414inter0, gate414inter1, gate414inter2, gate414inter3, gate414inter4, gate414inter5, gate414inter6, gate414inter7, gate414inter8, gate414inter9, gate414inter10, gate414inter11, gate414inter12, gate27inter0, gate27inter1, gate27inter2, gate27inter3, gate27inter4, gate27inter5, gate27inter6, gate27inter7, gate27inter8, gate27inter9, gate27inter10, gate27inter11, gate27inter12, gate84inter0, gate84inter1, gate84inter2, gate84inter3, gate84inter4, gate84inter5, gate84inter6, gate84inter7, gate84inter8, gate84inter9, gate84inter10, gate84inter11, gate84inter12, gate394inter0, gate394inter1, gate394inter2, gate394inter3, gate394inter4, gate394inter5, gate394inter6, gate394inter7, gate394inter8, gate394inter9, gate394inter10, gate394inter11, gate394inter12, gate36inter0, gate36inter1, gate36inter2, gate36inter3, gate36inter4, gate36inter5, gate36inter6, gate36inter7, gate36inter8, gate36inter9, gate36inter10, gate36inter11, gate36inter12, gate44inter0, gate44inter1, gate44inter2, gate44inter3, gate44inter4, gate44inter5, gate44inter6, gate44inter7, gate44inter8, gate44inter9, gate44inter10, gate44inter11, gate44inter12, gate283inter0, gate283inter1, gate283inter2, gate283inter3, gate283inter4, gate283inter5, gate283inter6, gate283inter7, gate283inter8, gate283inter9, gate283inter10, gate283inter11, gate283inter12, gate441inter0, gate441inter1, gate441inter2, gate441inter3, gate441inter4, gate441inter5, gate441inter6, gate441inter7, gate441inter8, gate441inter9, gate441inter10, gate441inter11, gate441inter12, gate428inter0, gate428inter1, gate428inter2, gate428inter3, gate428inter4, gate428inter5, gate428inter6, gate428inter7, gate428inter8, gate428inter9, gate428inter10, gate428inter11, gate428inter12, gate210inter0, gate210inter1, gate210inter2, gate210inter3, gate210inter4, gate210inter5, gate210inter6, gate210inter7, gate210inter8, gate210inter9, gate210inter10, gate210inter11, gate210inter12, gate415inter0, gate415inter1, gate415inter2, gate415inter3, gate415inter4, gate415inter5, gate415inter6, gate415inter7, gate415inter8, gate415inter9, gate415inter10, gate415inter11, gate415inter12, gate288inter0, gate288inter1, gate288inter2, gate288inter3, gate288inter4, gate288inter5, gate288inter6, gate288inter7, gate288inter8, gate288inter9, gate288inter10, gate288inter11, gate288inter12, gate144inter0, gate144inter1, gate144inter2, gate144inter3, gate144inter4, gate144inter5, gate144inter6, gate144inter7, gate144inter8, gate144inter9, gate144inter10, gate144inter11, gate144inter12, gate416inter0, gate416inter1, gate416inter2, gate416inter3, gate416inter4, gate416inter5, gate416inter6, gate416inter7, gate416inter8, gate416inter9, gate416inter10, gate416inter11, gate416inter12, gate131inter0, gate131inter1, gate131inter2, gate131inter3, gate131inter4, gate131inter5, gate131inter6, gate131inter7, gate131inter8, gate131inter9, gate131inter10, gate131inter11, gate131inter12, gate48inter0, gate48inter1, gate48inter2, gate48inter3, gate48inter4, gate48inter5, gate48inter6, gate48inter7, gate48inter8, gate48inter9, gate48inter10, gate48inter11, gate48inter12, gate46inter0, gate46inter1, gate46inter2, gate46inter3, gate46inter4, gate46inter5, gate46inter6, gate46inter7, gate46inter8, gate46inter9, gate46inter10, gate46inter11, gate46inter12, gate200inter0, gate200inter1, gate200inter2, gate200inter3, gate200inter4, gate200inter5, gate200inter6, gate200inter7, gate200inter8, gate200inter9, gate200inter10, gate200inter11, gate200inter12, gate137inter0, gate137inter1, gate137inter2, gate137inter3, gate137inter4, gate137inter5, gate137inter6, gate137inter7, gate137inter8, gate137inter9, gate137inter10, gate137inter11, gate137inter12, gate504inter0, gate504inter1, gate504inter2, gate504inter3, gate504inter4, gate504inter5, gate504inter6, gate504inter7, gate504inter8, gate504inter9, gate504inter10, gate504inter11, gate504inter12, gate201inter0, gate201inter1, gate201inter2, gate201inter3, gate201inter4, gate201inter5, gate201inter6, gate201inter7, gate201inter8, gate201inter9, gate201inter10, gate201inter11, gate201inter12, gate499inter0, gate499inter1, gate499inter2, gate499inter3, gate499inter4, gate499inter5, gate499inter6, gate499inter7, gate499inter8, gate499inter9, gate499inter10, gate499inter11, gate499inter12, gate63inter0, gate63inter1, gate63inter2, gate63inter3, gate63inter4, gate63inter5, gate63inter6, gate63inter7, gate63inter8, gate63inter9, gate63inter10, gate63inter11, gate63inter12, gate184inter0, gate184inter1, gate184inter2, gate184inter3, gate184inter4, gate184inter5, gate184inter6, gate184inter7, gate184inter8, gate184inter9, gate184inter10, gate184inter11, gate184inter12, gate228inter0, gate228inter1, gate228inter2, gate228inter3, gate228inter4, gate228inter5, gate228inter6, gate228inter7, gate228inter8, gate228inter9, gate228inter10, gate228inter11, gate228inter12, gate477inter0, gate477inter1, gate477inter2, gate477inter3, gate477inter4, gate477inter5, gate477inter6, gate477inter7, gate477inter8, gate477inter9, gate477inter10, gate477inter11, gate477inter12, gate221inter0, gate221inter1, gate221inter2, gate221inter3, gate221inter4, gate221inter5, gate221inter6, gate221inter7, gate221inter8, gate221inter9, gate221inter10, gate221inter11, gate221inter12, gate130inter0, gate130inter1, gate130inter2, gate130inter3, gate130inter4, gate130inter5, gate130inter6, gate130inter7, gate130inter8, gate130inter9, gate130inter10, gate130inter11, gate130inter12, gate280inter0, gate280inter1, gate280inter2, gate280inter3, gate280inter4, gate280inter5, gate280inter6, gate280inter7, gate280inter8, gate280inter9, gate280inter10, gate280inter11, gate280inter12, gate429inter0, gate429inter1, gate429inter2, gate429inter3, gate429inter4, gate429inter5, gate429inter6, gate429inter7, gate429inter8, gate429inter9, gate429inter10, gate429inter11, gate429inter12, gate253inter0, gate253inter1, gate253inter2, gate253inter3, gate253inter4, gate253inter5, gate253inter6, gate253inter7, gate253inter8, gate253inter9, gate253inter10, gate253inter11, gate253inter12, gate495inter0, gate495inter1, gate495inter2, gate495inter3, gate495inter4, gate495inter5, gate495inter6, gate495inter7, gate495inter8, gate495inter9, gate495inter10, gate495inter11, gate495inter12, gate26inter0, gate26inter1, gate26inter2, gate26inter3, gate26inter4, gate26inter5, gate26inter6, gate26inter7, gate26inter8, gate26inter9, gate26inter10, gate26inter11, gate26inter12, gate256inter0, gate256inter1, gate256inter2, gate256inter3, gate256inter4, gate256inter5, gate256inter6, gate256inter7, gate256inter8, gate256inter9, gate256inter10, gate256inter11, gate256inter12, gate81inter0, gate81inter1, gate81inter2, gate81inter3, gate81inter4, gate81inter5, gate81inter6, gate81inter7, gate81inter8, gate81inter9, gate81inter10, gate81inter11, gate81inter12, gate402inter0, gate402inter1, gate402inter2, gate402inter3, gate402inter4, gate402inter5, gate402inter6, gate402inter7, gate402inter8, gate402inter9, gate402inter10, gate402inter11, gate402inter12, gate106inter0, gate106inter1, gate106inter2, gate106inter3, gate106inter4, gate106inter5, gate106inter6, gate106inter7, gate106inter8, gate106inter9, gate106inter10, gate106inter11, gate106inter12, gate163inter0, gate163inter1, gate163inter2, gate163inter3, gate163inter4, gate163inter5, gate163inter6, gate163inter7, gate163inter8, gate163inter9, gate163inter10, gate163inter11, gate163inter12, gate181inter0, gate181inter1, gate181inter2, gate181inter3, gate181inter4, gate181inter5, gate181inter6, gate181inter7, gate181inter8, gate181inter9, gate181inter10, gate181inter11, gate181inter12, gate436inter0, gate436inter1, gate436inter2, gate436inter3, gate436inter4, gate436inter5, gate436inter6, gate436inter7, gate436inter8, gate436inter9, gate436inter10, gate436inter11, gate436inter12, gate391inter0, gate391inter1, gate391inter2, gate391inter3, gate391inter4, gate391inter5, gate391inter6, gate391inter7, gate391inter8, gate391inter9, gate391inter10, gate391inter11, gate391inter12, gate195inter0, gate195inter1, gate195inter2, gate195inter3, gate195inter4, gate195inter5, gate195inter6, gate195inter7, gate195inter8, gate195inter9, gate195inter10, gate195inter11, gate195inter12, gate456inter0, gate456inter1, gate456inter2, gate456inter3, gate456inter4, gate456inter5, gate456inter6, gate456inter7, gate456inter8, gate456inter9, gate456inter10, gate456inter11, gate456inter12, gate35inter0, gate35inter1, gate35inter2, gate35inter3, gate35inter4, gate35inter5, gate35inter6, gate35inter7, gate35inter8, gate35inter9, gate35inter10, gate35inter11, gate35inter12, gate237inter0, gate237inter1, gate237inter2, gate237inter3, gate237inter4, gate237inter5, gate237inter6, gate237inter7, gate237inter8, gate237inter9, gate237inter10, gate237inter11, gate237inter12, gate173inter0, gate173inter1, gate173inter2, gate173inter3, gate173inter4, gate173inter5, gate173inter6, gate173inter7, gate173inter8, gate173inter9, gate173inter10, gate173inter11, gate173inter12, gate32inter0, gate32inter1, gate32inter2, gate32inter3, gate32inter4, gate32inter5, gate32inter6, gate32inter7, gate32inter8, gate32inter9, gate32inter10, gate32inter11, gate32inter12, gate147inter0, gate147inter1, gate147inter2, gate147inter3, gate147inter4, gate147inter5, gate147inter6, gate147inter7, gate147inter8, gate147inter9, gate147inter10, gate147inter11, gate147inter12, gate258inter0, gate258inter1, gate258inter2, gate258inter3, gate258inter4, gate258inter5, gate258inter6, gate258inter7, gate258inter8, gate258inter9, gate258inter10, gate258inter11, gate258inter12, gate156inter0, gate156inter1, gate156inter2, gate156inter3, gate156inter4, gate156inter5, gate156inter6, gate156inter7, gate156inter8, gate156inter9, gate156inter10, gate156inter11, gate156inter12, gate212inter0, gate212inter1, gate212inter2, gate212inter3, gate212inter4, gate212inter5, gate212inter6, gate212inter7, gate212inter8, gate212inter9, gate212inter10, gate212inter11, gate212inter12, gate460inter0, gate460inter1, gate460inter2, gate460inter3, gate460inter4, gate460inter5, gate460inter6, gate460inter7, gate460inter8, gate460inter9, gate460inter10, gate460inter11, gate460inter12, gate56inter0, gate56inter1, gate56inter2, gate56inter3, gate56inter4, gate56inter5, gate56inter6, gate56inter7, gate56inter8, gate56inter9, gate56inter10, gate56inter11, gate56inter12, gate76inter0, gate76inter1, gate76inter2, gate76inter3, gate76inter4, gate76inter5, gate76inter6, gate76inter7, gate76inter8, gate76inter9, gate76inter10, gate76inter11, gate76inter12, gate215inter0, gate215inter1, gate215inter2, gate215inter3, gate215inter4, gate215inter5, gate215inter6, gate215inter7, gate215inter8, gate215inter9, gate215inter10, gate215inter11, gate215inter12, gate138inter0, gate138inter1, gate138inter2, gate138inter3, gate138inter4, gate138inter5, gate138inter6, gate138inter7, gate138inter8, gate138inter9, gate138inter10, gate138inter11, gate138inter12, gate19inter0, gate19inter1, gate19inter2, gate19inter3, gate19inter4, gate19inter5, gate19inter6, gate19inter7, gate19inter8, gate19inter9, gate19inter10, gate19inter11, gate19inter12, gate511inter0, gate511inter1, gate511inter2, gate511inter3, gate511inter4, gate511inter5, gate511inter6, gate511inter7, gate511inter8, gate511inter9, gate511inter10, gate511inter11, gate511inter12, gate483inter0, gate483inter1, gate483inter2, gate483inter3, gate483inter4, gate483inter5, gate483inter6, gate483inter7, gate483inter8, gate483inter9, gate483inter10, gate483inter11, gate483inter12, gate188inter0, gate188inter1, gate188inter2, gate188inter3, gate188inter4, gate188inter5, gate188inter6, gate188inter7, gate188inter8, gate188inter9, gate188inter10, gate188inter11, gate188inter12, gate470inter0, gate470inter1, gate470inter2, gate470inter3, gate470inter4, gate470inter5, gate470inter6, gate470inter7, gate470inter8, gate470inter9, gate470inter10, gate470inter11, gate470inter12, gate10inter0, gate10inter1, gate10inter2, gate10inter3, gate10inter4, gate10inter5, gate10inter6, gate10inter7, gate10inter8, gate10inter9, gate10inter10, gate10inter11, gate10inter12, gate290inter0, gate290inter1, gate290inter2, gate290inter3, gate290inter4, gate290inter5, gate290inter6, gate290inter7, gate290inter8, gate290inter9, gate290inter10, gate290inter11, gate290inter12, gate479inter0, gate479inter1, gate479inter2, gate479inter3, gate479inter4, gate479inter5, gate479inter6, gate479inter7, gate479inter8, gate479inter9, gate479inter10, gate479inter11, gate479inter12, gate189inter0, gate189inter1, gate189inter2, gate189inter3, gate189inter4, gate189inter5, gate189inter6, gate189inter7, gate189inter8, gate189inter9, gate189inter10, gate189inter11, gate189inter12, gate128inter0, gate128inter1, gate128inter2, gate128inter3, gate128inter4, gate128inter5, gate128inter6, gate128inter7, gate128inter8, gate128inter9, gate128inter10, gate128inter11, gate128inter12, gate155inter0, gate155inter1, gate155inter2, gate155inter3, gate155inter4, gate155inter5, gate155inter6, gate155inter7, gate155inter8, gate155inter9, gate155inter10, gate155inter11, gate155inter12, gate407inter0, gate407inter1, gate407inter2, gate407inter3, gate407inter4, gate407inter5, gate407inter6, gate407inter7, gate407inter8, gate407inter9, gate407inter10, gate407inter11, gate407inter12, gate403inter0, gate403inter1, gate403inter2, gate403inter3, gate403inter4, gate403inter5, gate403inter6, gate403inter7, gate403inter8, gate403inter9, gate403inter10, gate403inter11, gate403inter12, gate170inter0, gate170inter1, gate170inter2, gate170inter3, gate170inter4, gate170inter5, gate170inter6, gate170inter7, gate170inter8, gate170inter9, gate170inter10, gate170inter11, gate170inter12, gate430inter0, gate430inter1, gate430inter2, gate430inter3, gate430inter4, gate430inter5, gate430inter6, gate430inter7, gate430inter8, gate430inter9, gate430inter10, gate430inter11, gate430inter12, gate229inter0, gate229inter1, gate229inter2, gate229inter3, gate229inter4, gate229inter5, gate229inter6, gate229inter7, gate229inter8, gate229inter9, gate229inter10, gate229inter11, gate229inter12, gate116inter0, gate116inter1, gate116inter2, gate116inter3, gate116inter4, gate116inter5, gate116inter6, gate116inter7, gate116inter8, gate116inter9, gate116inter10, gate116inter11, gate116inter12, gate149inter0, gate149inter1, gate149inter2, gate149inter3, gate149inter4, gate149inter5, gate149inter6, gate149inter7, gate149inter8, gate149inter9, gate149inter10, gate149inter11, gate149inter12, gate91inter0, gate91inter1, gate91inter2, gate91inter3, gate91inter4, gate91inter5, gate91inter6, gate91inter7, gate91inter8, gate91inter9, gate91inter10, gate91inter11, gate91inter12, gate70inter0, gate70inter1, gate70inter2, gate70inter3, gate70inter4, gate70inter5, gate70inter6, gate70inter7, gate70inter8, gate70inter9, gate70inter10, gate70inter11, gate70inter12, gate14inter0, gate14inter1, gate14inter2, gate14inter3, gate14inter4, gate14inter5, gate14inter6, gate14inter7, gate14inter8, gate14inter9, gate14inter10, gate14inter11, gate14inter12, gate85inter0, gate85inter1, gate85inter2, gate85inter3, gate85inter4, gate85inter5, gate85inter6, gate85inter7, gate85inter8, gate85inter9, gate85inter10, gate85inter11, gate85inter12, gate118inter0, gate118inter1, gate118inter2, gate118inter3, gate118inter4, gate118inter5, gate118inter6, gate118inter7, gate118inter8, gate118inter9, gate118inter10, gate118inter11, gate118inter12, gate208inter0, gate208inter1, gate208inter2, gate208inter3, gate208inter4, gate208inter5, gate208inter6, gate208inter7, gate208inter8, gate208inter9, gate208inter10, gate208inter11, gate208inter12, gate153inter0, gate153inter1, gate153inter2, gate153inter3, gate153inter4, gate153inter5, gate153inter6, gate153inter7, gate153inter8, gate153inter9, gate153inter10, gate153inter11, gate153inter12, gate439inter0, gate439inter1, gate439inter2, gate439inter3, gate439inter4, gate439inter5, gate439inter6, gate439inter7, gate439inter8, gate439inter9, gate439inter10, gate439inter11, gate439inter12, gate404inter0, gate404inter1, gate404inter2, gate404inter3, gate404inter4, gate404inter5, gate404inter6, gate404inter7, gate404inter8, gate404inter9, gate404inter10, gate404inter11, gate404inter12, gate254inter0, gate254inter1, gate254inter2, gate254inter3, gate254inter4, gate254inter5, gate254inter6, gate254inter7, gate254inter8, gate254inter9, gate254inter10, gate254inter11, gate254inter12, gate467inter0, gate467inter1, gate467inter2, gate467inter3, gate467inter4, gate467inter5, gate467inter6, gate467inter7, gate467inter8, gate467inter9, gate467inter10, gate467inter11, gate467inter12, gate104inter0, gate104inter1, gate104inter2, gate104inter3, gate104inter4, gate104inter5, gate104inter6, gate104inter7, gate104inter8, gate104inter9, gate104inter10, gate104inter11, gate104inter12, gate126inter0, gate126inter1, gate126inter2, gate126inter3, gate126inter4, gate126inter5, gate126inter6, gate126inter7, gate126inter8, gate126inter9, gate126inter10, gate126inter11, gate126inter12, gate31inter0, gate31inter1, gate31inter2, gate31inter3, gate31inter4, gate31inter5, gate31inter6, gate31inter7, gate31inter8, gate31inter9, gate31inter10, gate31inter11, gate31inter12, gate98inter0, gate98inter1, gate98inter2, gate98inter3, gate98inter4, gate98inter5, gate98inter6, gate98inter7, gate98inter8, gate98inter9, gate98inter10, gate98inter11, gate98inter12, gate218inter0, gate218inter1, gate218inter2, gate218inter3, gate218inter4, gate218inter5, gate218inter6, gate218inter7, gate218inter8, gate218inter9, gate218inter10, gate218inter11, gate218inter12, gate207inter0, gate207inter1, gate207inter2, gate207inter3, gate207inter4, gate207inter5, gate207inter6, gate207inter7, gate207inter8, gate207inter9, gate207inter10, gate207inter11, gate207inter12, gate485inter0, gate485inter1, gate485inter2, gate485inter3, gate485inter4, gate485inter5, gate485inter6, gate485inter7, gate485inter8, gate485inter9, gate485inter10, gate485inter11, gate485inter12, gate16inter0, gate16inter1, gate16inter2, gate16inter3, gate16inter4, gate16inter5, gate16inter6, gate16inter7, gate16inter8, gate16inter9, gate16inter10, gate16inter11, gate16inter12, gate50inter0, gate50inter1, gate50inter2, gate50inter3, gate50inter4, gate50inter5, gate50inter6, gate50inter7, gate50inter8, gate50inter9, gate50inter10, gate50inter11, gate50inter12, gate480inter0, gate480inter1, gate480inter2, gate480inter3, gate480inter4, gate480inter5, gate480inter6, gate480inter7, gate480inter8, gate480inter9, gate480inter10, gate480inter11, gate480inter12, gate78inter0, gate78inter1, gate78inter2, gate78inter3, gate78inter4, gate78inter5, gate78inter6, gate78inter7, gate78inter8, gate78inter9, gate78inter10, gate78inter11, gate78inter12, gate510inter0, gate510inter1, gate510inter2, gate510inter3, gate510inter4, gate510inter5, gate510inter6, gate510inter7, gate510inter8, gate510inter9, gate510inter10, gate510inter11, gate510inter12, gate82inter0, gate82inter1, gate82inter2, gate82inter3, gate82inter4, gate82inter5, gate82inter6, gate82inter7, gate82inter8, gate82inter9, gate82inter10, gate82inter11, gate82inter12, gate220inter0, gate220inter1, gate220inter2, gate220inter3, gate220inter4, gate220inter5, gate220inter6, gate220inter7, gate220inter8, gate220inter9, gate220inter10, gate220inter11, gate220inter12, gate176inter0, gate176inter1, gate176inter2, gate176inter3, gate176inter4, gate176inter5, gate176inter6, gate176inter7, gate176inter8, gate176inter9, gate176inter10, gate176inter11, gate176inter12, gate39inter0, gate39inter1, gate39inter2, gate39inter3, gate39inter4, gate39inter5, gate39inter6, gate39inter7, gate39inter8, gate39inter9, gate39inter10, gate39inter11, gate39inter12, gate473inter0, gate473inter1, gate473inter2, gate473inter3, gate473inter4, gate473inter5, gate473inter6, gate473inter7, gate473inter8, gate473inter9, gate473inter10, gate473inter11, gate473inter12, gate241inter0, gate241inter1, gate241inter2, gate241inter3, gate241inter4, gate241inter5, gate241inter6, gate241inter7, gate241inter8, gate241inter9, gate241inter10, gate241inter11, gate241inter12, gate247inter0, gate247inter1, gate247inter2, gate247inter3, gate247inter4, gate247inter5, gate247inter6, gate247inter7, gate247inter8, gate247inter9, gate247inter10, gate247inter11, gate247inter12, gate224inter0, gate224inter1, gate224inter2, gate224inter3, gate224inter4, gate224inter5, gate224inter6, gate224inter7, gate224inter8, gate224inter9, gate224inter10, gate224inter11, gate224inter12, gate196inter0, gate196inter1, gate196inter2, gate196inter3, gate196inter4, gate196inter5, gate196inter6, gate196inter7, gate196inter8, gate196inter9, gate196inter10, gate196inter11, gate196inter12, gate180inter0, gate180inter1, gate180inter2, gate180inter3, gate180inter4, gate180inter5, gate180inter6, gate180inter7, gate180inter8, gate180inter9, gate180inter10, gate180inter11, gate180inter12, gate238inter0, gate238inter1, gate238inter2, gate238inter3, gate238inter4, gate238inter5, gate238inter6, gate238inter7, gate238inter8, gate238inter9, gate238inter10, gate238inter11, gate238inter12, gate17inter0, gate17inter1, gate17inter2, gate17inter3, gate17inter4, gate17inter5, gate17inter6, gate17inter7, gate17inter8, gate17inter9, gate17inter10, gate17inter11, gate17inter12, gate469inter0, gate469inter1, gate469inter2, gate469inter3, gate469inter4, gate469inter5, gate469inter6, gate469inter7, gate469inter8, gate469inter9, gate469inter10, gate469inter11, gate469inter12, gate267inter0, gate267inter1, gate267inter2, gate267inter3, gate267inter4, gate267inter5, gate267inter6, gate267inter7, gate267inter8, gate267inter9, gate267inter10, gate267inter11, gate267inter12, gate513inter0, gate513inter1, gate513inter2, gate513inter3, gate513inter4, gate513inter5, gate513inter6, gate513inter7, gate513inter8, gate513inter9, gate513inter10, gate513inter11, gate513inter12, gate453inter0, gate453inter1, gate453inter2, gate453inter3, gate453inter4, gate453inter5, gate453inter6, gate453inter7, gate453inter8, gate453inter9, gate453inter10, gate453inter11, gate453inter12, gate243inter0, gate243inter1, gate243inter2, gate243inter3, gate243inter4, gate243inter5, gate243inter6, gate243inter7, gate243inter8, gate243inter9, gate243inter10, gate243inter11, gate243inter12, gate233inter0, gate233inter1, gate233inter2, gate233inter3, gate233inter4, gate233inter5, gate233inter6, gate233inter7, gate233inter8, gate233inter9, gate233inter10, gate233inter11, gate233inter12, gate264inter0, gate264inter1, gate264inter2, gate264inter3, gate264inter4, gate264inter5, gate264inter6, gate264inter7, gate264inter8, gate264inter9, gate264inter10, gate264inter11, gate264inter12, gate419inter0, gate419inter1, gate419inter2, gate419inter3, gate419inter4, gate419inter5, gate419inter6, gate419inter7, gate419inter8, gate419inter9, gate419inter10, gate419inter11, gate419inter12, gate249inter0, gate249inter1, gate249inter2, gate249inter3, gate249inter4, gate249inter5, gate249inter6, gate249inter7, gate249inter8, gate249inter9, gate249inter10, gate249inter11, gate249inter12, gate102inter0, gate102inter1, gate102inter2, gate102inter3, gate102inter4, gate102inter5, gate102inter6, gate102inter7, gate102inter8, gate102inter9, gate102inter10, gate102inter11, gate102inter12, gate67inter0, gate67inter1, gate67inter2, gate67inter3, gate67inter4, gate67inter5, gate67inter6, gate67inter7, gate67inter8, gate67inter9, gate67inter10, gate67inter11, gate67inter12, gate129inter0, gate129inter1, gate129inter2, gate129inter3, gate129inter4, gate129inter5, gate129inter6, gate129inter7, gate129inter8, gate129inter9, gate129inter10, gate129inter11, gate129inter12, gate115inter0, gate115inter1, gate115inter2, gate115inter3, gate115inter4, gate115inter5, gate115inter6, gate115inter7, gate115inter8, gate115inter9, gate115inter10, gate115inter11, gate115inter12, gate397inter0, gate397inter1, gate397inter2, gate397inter3, gate397inter4, gate397inter5, gate397inter6, gate397inter7, gate397inter8, gate397inter9, gate397inter10, gate397inter11, gate397inter12, gate505inter0, gate505inter1, gate505inter2, gate505inter3, gate505inter4, gate505inter5, gate505inter6, gate505inter7, gate505inter8, gate505inter9, gate505inter10, gate505inter11, gate505inter12, gate89inter0, gate89inter1, gate89inter2, gate89inter3, gate89inter4, gate89inter5, gate89inter6, gate89inter7, gate89inter8, gate89inter9, gate89inter10, gate89inter11, gate89inter12, gate447inter0, gate447inter1, gate447inter2, gate447inter3, gate447inter4, gate447inter5, gate447inter6, gate447inter7, gate447inter8, gate447inter9, gate447inter10, gate447inter11, gate447inter12, gate449inter0, gate449inter1, gate449inter2, gate449inter3, gate449inter4, gate449inter5, gate449inter6, gate449inter7, gate449inter8, gate449inter9, gate449inter10, gate449inter11, gate449inter12, gate514inter0, gate514inter1, gate514inter2, gate514inter3, gate514inter4, gate514inter5, gate514inter6, gate514inter7, gate514inter8, gate514inter9, gate514inter10, gate514inter11, gate514inter12, gate395inter0, gate395inter1, gate395inter2, gate395inter3, gate395inter4, gate395inter5, gate395inter6, gate395inter7, gate395inter8, gate395inter9, gate395inter10, gate395inter11, gate395inter12;



and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );

  xor2  gate1233(.a(G2), .b(G1), .O(gate9inter0));
  nand2 gate1234(.a(gate9inter0), .b(s_98), .O(gate9inter1));
  and2  gate1235(.a(G2), .b(G1), .O(gate9inter2));
  inv1  gate1236(.a(s_98), .O(gate9inter3));
  inv1  gate1237(.a(s_99), .O(gate9inter4));
  nand2 gate1238(.a(gate9inter4), .b(gate9inter3), .O(gate9inter5));
  nor2  gate1239(.a(gate9inter5), .b(gate9inter2), .O(gate9inter6));
  inv1  gate1240(.a(G1), .O(gate9inter7));
  inv1  gate1241(.a(G2), .O(gate9inter8));
  nand2 gate1242(.a(gate9inter8), .b(gate9inter7), .O(gate9inter9));
  nand2 gate1243(.a(s_99), .b(gate9inter3), .O(gate9inter10));
  nor2  gate1244(.a(gate9inter10), .b(gate9inter9), .O(gate9inter11));
  nor2  gate1245(.a(gate9inter11), .b(gate9inter6), .O(gate9inter12));
  nand2 gate1246(.a(gate9inter12), .b(gate9inter1), .O(G266));

  xor2  gate2199(.a(G4), .b(G3), .O(gate10inter0));
  nand2 gate2200(.a(gate10inter0), .b(s_236), .O(gate10inter1));
  and2  gate2201(.a(G4), .b(G3), .O(gate10inter2));
  inv1  gate2202(.a(s_236), .O(gate10inter3));
  inv1  gate2203(.a(s_237), .O(gate10inter4));
  nand2 gate2204(.a(gate10inter4), .b(gate10inter3), .O(gate10inter5));
  nor2  gate2205(.a(gate10inter5), .b(gate10inter2), .O(gate10inter6));
  inv1  gate2206(.a(G3), .O(gate10inter7));
  inv1  gate2207(.a(G4), .O(gate10inter8));
  nand2 gate2208(.a(gate10inter8), .b(gate10inter7), .O(gate10inter9));
  nand2 gate2209(.a(s_237), .b(gate10inter3), .O(gate10inter10));
  nor2  gate2210(.a(gate10inter10), .b(gate10inter9), .O(gate10inter11));
  nor2  gate2211(.a(gate10inter11), .b(gate10inter6), .O(gate10inter12));
  nand2 gate2212(.a(gate10inter12), .b(gate10inter1), .O(G269));
nand2 gate11( .a(G5), .b(G6), .O(G272) );
nand2 gate12( .a(G7), .b(G8), .O(G275) );

  xor2  gate897(.a(G10), .b(G9), .O(gate13inter0));
  nand2 gate898(.a(gate13inter0), .b(s_50), .O(gate13inter1));
  and2  gate899(.a(G10), .b(G9), .O(gate13inter2));
  inv1  gate900(.a(s_50), .O(gate13inter3));
  inv1  gate901(.a(s_51), .O(gate13inter4));
  nand2 gate902(.a(gate13inter4), .b(gate13inter3), .O(gate13inter5));
  nor2  gate903(.a(gate13inter5), .b(gate13inter2), .O(gate13inter6));
  inv1  gate904(.a(G9), .O(gate13inter7));
  inv1  gate905(.a(G10), .O(gate13inter8));
  nand2 gate906(.a(gate13inter8), .b(gate13inter7), .O(gate13inter9));
  nand2 gate907(.a(s_51), .b(gate13inter3), .O(gate13inter10));
  nor2  gate908(.a(gate13inter10), .b(gate13inter9), .O(gate13inter11));
  nor2  gate909(.a(gate13inter11), .b(gate13inter6), .O(gate13inter12));
  nand2 gate910(.a(gate13inter12), .b(gate13inter1), .O(G278));

  xor2  gate2409(.a(G12), .b(G11), .O(gate14inter0));
  nand2 gate2410(.a(gate14inter0), .b(s_266), .O(gate14inter1));
  and2  gate2411(.a(G12), .b(G11), .O(gate14inter2));
  inv1  gate2412(.a(s_266), .O(gate14inter3));
  inv1  gate2413(.a(s_267), .O(gate14inter4));
  nand2 gate2414(.a(gate14inter4), .b(gate14inter3), .O(gate14inter5));
  nor2  gate2415(.a(gate14inter5), .b(gate14inter2), .O(gate14inter6));
  inv1  gate2416(.a(G11), .O(gate14inter7));
  inv1  gate2417(.a(G12), .O(gate14inter8));
  nand2 gate2418(.a(gate14inter8), .b(gate14inter7), .O(gate14inter9));
  nand2 gate2419(.a(s_267), .b(gate14inter3), .O(gate14inter10));
  nor2  gate2420(.a(gate14inter10), .b(gate14inter9), .O(gate14inter11));
  nor2  gate2421(.a(gate14inter11), .b(gate14inter6), .O(gate14inter12));
  nand2 gate2422(.a(gate14inter12), .b(gate14inter1), .O(G281));
nand2 gate15( .a(G13), .b(G14), .O(G284) );

  xor2  gate2633(.a(G16), .b(G15), .O(gate16inter0));
  nand2 gate2634(.a(gate16inter0), .b(s_298), .O(gate16inter1));
  and2  gate2635(.a(G16), .b(G15), .O(gate16inter2));
  inv1  gate2636(.a(s_298), .O(gate16inter3));
  inv1  gate2637(.a(s_299), .O(gate16inter4));
  nand2 gate2638(.a(gate16inter4), .b(gate16inter3), .O(gate16inter5));
  nor2  gate2639(.a(gate16inter5), .b(gate16inter2), .O(gate16inter6));
  inv1  gate2640(.a(G15), .O(gate16inter7));
  inv1  gate2641(.a(G16), .O(gate16inter8));
  nand2 gate2642(.a(gate16inter8), .b(gate16inter7), .O(gate16inter9));
  nand2 gate2643(.a(s_299), .b(gate16inter3), .O(gate16inter10));
  nor2  gate2644(.a(gate16inter10), .b(gate16inter9), .O(gate16inter11));
  nor2  gate2645(.a(gate16inter11), .b(gate16inter6), .O(gate16inter12));
  nand2 gate2646(.a(gate16inter12), .b(gate16inter1), .O(G287));

  xor2  gate2857(.a(G18), .b(G17), .O(gate17inter0));
  nand2 gate2858(.a(gate17inter0), .b(s_330), .O(gate17inter1));
  and2  gate2859(.a(G18), .b(G17), .O(gate17inter2));
  inv1  gate2860(.a(s_330), .O(gate17inter3));
  inv1  gate2861(.a(s_331), .O(gate17inter4));
  nand2 gate2862(.a(gate17inter4), .b(gate17inter3), .O(gate17inter5));
  nor2  gate2863(.a(gate17inter5), .b(gate17inter2), .O(gate17inter6));
  inv1  gate2864(.a(G17), .O(gate17inter7));
  inv1  gate2865(.a(G18), .O(gate17inter8));
  nand2 gate2866(.a(gate17inter8), .b(gate17inter7), .O(gate17inter9));
  nand2 gate2867(.a(s_331), .b(gate17inter3), .O(gate17inter10));
  nor2  gate2868(.a(gate17inter10), .b(gate17inter9), .O(gate17inter11));
  nor2  gate2869(.a(gate17inter11), .b(gate17inter6), .O(gate17inter12));
  nand2 gate2870(.a(gate17inter12), .b(gate17inter1), .O(G290));
nand2 gate18( .a(G19), .b(G20), .O(G293) );

  xor2  gate2129(.a(G22), .b(G21), .O(gate19inter0));
  nand2 gate2130(.a(gate19inter0), .b(s_226), .O(gate19inter1));
  and2  gate2131(.a(G22), .b(G21), .O(gate19inter2));
  inv1  gate2132(.a(s_226), .O(gate19inter3));
  inv1  gate2133(.a(s_227), .O(gate19inter4));
  nand2 gate2134(.a(gate19inter4), .b(gate19inter3), .O(gate19inter5));
  nor2  gate2135(.a(gate19inter5), .b(gate19inter2), .O(gate19inter6));
  inv1  gate2136(.a(G21), .O(gate19inter7));
  inv1  gate2137(.a(G22), .O(gate19inter8));
  nand2 gate2138(.a(gate19inter8), .b(gate19inter7), .O(gate19inter9));
  nand2 gate2139(.a(s_227), .b(gate19inter3), .O(gate19inter10));
  nor2  gate2140(.a(gate19inter10), .b(gate19inter9), .O(gate19inter11));
  nor2  gate2141(.a(gate19inter11), .b(gate19inter6), .O(gate19inter12));
  nand2 gate2142(.a(gate19inter12), .b(gate19inter1), .O(G296));
nand2 gate20( .a(G23), .b(G24), .O(G299) );
nand2 gate21( .a(G25), .b(G26), .O(G302) );
nand2 gate22( .a(G27), .b(G28), .O(G305) );
nand2 gate23( .a(G29), .b(G30), .O(G308) );
nand2 gate24( .a(G31), .b(G32), .O(G311) );
nand2 gate25( .a(G1), .b(G5), .O(G314) );

  xor2  gate1793(.a(G13), .b(G9), .O(gate26inter0));
  nand2 gate1794(.a(gate26inter0), .b(s_178), .O(gate26inter1));
  and2  gate1795(.a(G13), .b(G9), .O(gate26inter2));
  inv1  gate1796(.a(s_178), .O(gate26inter3));
  inv1  gate1797(.a(s_179), .O(gate26inter4));
  nand2 gate1798(.a(gate26inter4), .b(gate26inter3), .O(gate26inter5));
  nor2  gate1799(.a(gate26inter5), .b(gate26inter2), .O(gate26inter6));
  inv1  gate1800(.a(G9), .O(gate26inter7));
  inv1  gate1801(.a(G13), .O(gate26inter8));
  nand2 gate1802(.a(gate26inter8), .b(gate26inter7), .O(gate26inter9));
  nand2 gate1803(.a(s_179), .b(gate26inter3), .O(gate26inter10));
  nor2  gate1804(.a(gate26inter10), .b(gate26inter9), .O(gate26inter11));
  nor2  gate1805(.a(gate26inter11), .b(gate26inter6), .O(gate26inter12));
  nand2 gate1806(.a(gate26inter12), .b(gate26inter1), .O(G317));

  xor2  gate1359(.a(G6), .b(G2), .O(gate27inter0));
  nand2 gate1360(.a(gate27inter0), .b(s_116), .O(gate27inter1));
  and2  gate1361(.a(G6), .b(G2), .O(gate27inter2));
  inv1  gate1362(.a(s_116), .O(gate27inter3));
  inv1  gate1363(.a(s_117), .O(gate27inter4));
  nand2 gate1364(.a(gate27inter4), .b(gate27inter3), .O(gate27inter5));
  nor2  gate1365(.a(gate27inter5), .b(gate27inter2), .O(gate27inter6));
  inv1  gate1366(.a(G2), .O(gate27inter7));
  inv1  gate1367(.a(G6), .O(gate27inter8));
  nand2 gate1368(.a(gate27inter8), .b(gate27inter7), .O(gate27inter9));
  nand2 gate1369(.a(s_117), .b(gate27inter3), .O(gate27inter10));
  nor2  gate1370(.a(gate27inter10), .b(gate27inter9), .O(gate27inter11));
  nor2  gate1371(.a(gate27inter11), .b(gate27inter6), .O(gate27inter12));
  nand2 gate1372(.a(gate27inter12), .b(gate27inter1), .O(G320));
nand2 gate28( .a(G10), .b(G14), .O(G323) );
nand2 gate29( .a(G3), .b(G7), .O(G326) );

  xor2  gate757(.a(G15), .b(G11), .O(gate30inter0));
  nand2 gate758(.a(gate30inter0), .b(s_30), .O(gate30inter1));
  and2  gate759(.a(G15), .b(G11), .O(gate30inter2));
  inv1  gate760(.a(s_30), .O(gate30inter3));
  inv1  gate761(.a(s_31), .O(gate30inter4));
  nand2 gate762(.a(gate30inter4), .b(gate30inter3), .O(gate30inter5));
  nor2  gate763(.a(gate30inter5), .b(gate30inter2), .O(gate30inter6));
  inv1  gate764(.a(G11), .O(gate30inter7));
  inv1  gate765(.a(G15), .O(gate30inter8));
  nand2 gate766(.a(gate30inter8), .b(gate30inter7), .O(gate30inter9));
  nand2 gate767(.a(s_31), .b(gate30inter3), .O(gate30inter10));
  nor2  gate768(.a(gate30inter10), .b(gate30inter9), .O(gate30inter11));
  nor2  gate769(.a(gate30inter11), .b(gate30inter6), .O(gate30inter12));
  nand2 gate770(.a(gate30inter12), .b(gate30inter1), .O(G329));

  xor2  gate2563(.a(G8), .b(G4), .O(gate31inter0));
  nand2 gate2564(.a(gate31inter0), .b(s_288), .O(gate31inter1));
  and2  gate2565(.a(G8), .b(G4), .O(gate31inter2));
  inv1  gate2566(.a(s_288), .O(gate31inter3));
  inv1  gate2567(.a(s_289), .O(gate31inter4));
  nand2 gate2568(.a(gate31inter4), .b(gate31inter3), .O(gate31inter5));
  nor2  gate2569(.a(gate31inter5), .b(gate31inter2), .O(gate31inter6));
  inv1  gate2570(.a(G4), .O(gate31inter7));
  inv1  gate2571(.a(G8), .O(gate31inter8));
  nand2 gate2572(.a(gate31inter8), .b(gate31inter7), .O(gate31inter9));
  nand2 gate2573(.a(s_289), .b(gate31inter3), .O(gate31inter10));
  nor2  gate2574(.a(gate31inter10), .b(gate31inter9), .O(gate31inter11));
  nor2  gate2575(.a(gate31inter11), .b(gate31inter6), .O(gate31inter12));
  nand2 gate2576(.a(gate31inter12), .b(gate31inter1), .O(G332));

  xor2  gate1989(.a(G16), .b(G12), .O(gate32inter0));
  nand2 gate1990(.a(gate32inter0), .b(s_206), .O(gate32inter1));
  and2  gate1991(.a(G16), .b(G12), .O(gate32inter2));
  inv1  gate1992(.a(s_206), .O(gate32inter3));
  inv1  gate1993(.a(s_207), .O(gate32inter4));
  nand2 gate1994(.a(gate32inter4), .b(gate32inter3), .O(gate32inter5));
  nor2  gate1995(.a(gate32inter5), .b(gate32inter2), .O(gate32inter6));
  inv1  gate1996(.a(G12), .O(gate32inter7));
  inv1  gate1997(.a(G16), .O(gate32inter8));
  nand2 gate1998(.a(gate32inter8), .b(gate32inter7), .O(gate32inter9));
  nand2 gate1999(.a(s_207), .b(gate32inter3), .O(gate32inter10));
  nor2  gate2000(.a(gate32inter10), .b(gate32inter9), .O(gate32inter11));
  nor2  gate2001(.a(gate32inter11), .b(gate32inter6), .O(gate32inter12));
  nand2 gate2002(.a(gate32inter12), .b(gate32inter1), .O(G335));
nand2 gate33( .a(G17), .b(G21), .O(G338) );
nand2 gate34( .a(G25), .b(G29), .O(G341) );

  xor2  gate1947(.a(G22), .b(G18), .O(gate35inter0));
  nand2 gate1948(.a(gate35inter0), .b(s_200), .O(gate35inter1));
  and2  gate1949(.a(G22), .b(G18), .O(gate35inter2));
  inv1  gate1950(.a(s_200), .O(gate35inter3));
  inv1  gate1951(.a(s_201), .O(gate35inter4));
  nand2 gate1952(.a(gate35inter4), .b(gate35inter3), .O(gate35inter5));
  nor2  gate1953(.a(gate35inter5), .b(gate35inter2), .O(gate35inter6));
  inv1  gate1954(.a(G18), .O(gate35inter7));
  inv1  gate1955(.a(G22), .O(gate35inter8));
  nand2 gate1956(.a(gate35inter8), .b(gate35inter7), .O(gate35inter9));
  nand2 gate1957(.a(s_201), .b(gate35inter3), .O(gate35inter10));
  nor2  gate1958(.a(gate35inter10), .b(gate35inter9), .O(gate35inter11));
  nor2  gate1959(.a(gate35inter11), .b(gate35inter6), .O(gate35inter12));
  nand2 gate1960(.a(gate35inter12), .b(gate35inter1), .O(G344));

  xor2  gate1401(.a(G30), .b(G26), .O(gate36inter0));
  nand2 gate1402(.a(gate36inter0), .b(s_122), .O(gate36inter1));
  and2  gate1403(.a(G30), .b(G26), .O(gate36inter2));
  inv1  gate1404(.a(s_122), .O(gate36inter3));
  inv1  gate1405(.a(s_123), .O(gate36inter4));
  nand2 gate1406(.a(gate36inter4), .b(gate36inter3), .O(gate36inter5));
  nor2  gate1407(.a(gate36inter5), .b(gate36inter2), .O(gate36inter6));
  inv1  gate1408(.a(G26), .O(gate36inter7));
  inv1  gate1409(.a(G30), .O(gate36inter8));
  nand2 gate1410(.a(gate36inter8), .b(gate36inter7), .O(gate36inter9));
  nand2 gate1411(.a(s_123), .b(gate36inter3), .O(gate36inter10));
  nor2  gate1412(.a(gate36inter10), .b(gate36inter9), .O(gate36inter11));
  nor2  gate1413(.a(gate36inter11), .b(gate36inter6), .O(gate36inter12));
  nand2 gate1414(.a(gate36inter12), .b(gate36inter1), .O(G347));
nand2 gate37( .a(G19), .b(G23), .O(G350) );

  xor2  gate701(.a(G31), .b(G27), .O(gate38inter0));
  nand2 gate702(.a(gate38inter0), .b(s_22), .O(gate38inter1));
  and2  gate703(.a(G31), .b(G27), .O(gate38inter2));
  inv1  gate704(.a(s_22), .O(gate38inter3));
  inv1  gate705(.a(s_23), .O(gate38inter4));
  nand2 gate706(.a(gate38inter4), .b(gate38inter3), .O(gate38inter5));
  nor2  gate707(.a(gate38inter5), .b(gate38inter2), .O(gate38inter6));
  inv1  gate708(.a(G27), .O(gate38inter7));
  inv1  gate709(.a(G31), .O(gate38inter8));
  nand2 gate710(.a(gate38inter8), .b(gate38inter7), .O(gate38inter9));
  nand2 gate711(.a(s_23), .b(gate38inter3), .O(gate38inter10));
  nor2  gate712(.a(gate38inter10), .b(gate38inter9), .O(gate38inter11));
  nor2  gate713(.a(gate38inter11), .b(gate38inter6), .O(gate38inter12));
  nand2 gate714(.a(gate38inter12), .b(gate38inter1), .O(G353));

  xor2  gate2745(.a(G24), .b(G20), .O(gate39inter0));
  nand2 gate2746(.a(gate39inter0), .b(s_314), .O(gate39inter1));
  and2  gate2747(.a(G24), .b(G20), .O(gate39inter2));
  inv1  gate2748(.a(s_314), .O(gate39inter3));
  inv1  gate2749(.a(s_315), .O(gate39inter4));
  nand2 gate2750(.a(gate39inter4), .b(gate39inter3), .O(gate39inter5));
  nor2  gate2751(.a(gate39inter5), .b(gate39inter2), .O(gate39inter6));
  inv1  gate2752(.a(G20), .O(gate39inter7));
  inv1  gate2753(.a(G24), .O(gate39inter8));
  nand2 gate2754(.a(gate39inter8), .b(gate39inter7), .O(gate39inter9));
  nand2 gate2755(.a(s_315), .b(gate39inter3), .O(gate39inter10));
  nor2  gate2756(.a(gate39inter10), .b(gate39inter9), .O(gate39inter11));
  nor2  gate2757(.a(gate39inter11), .b(gate39inter6), .O(gate39inter12));
  nand2 gate2758(.a(gate39inter12), .b(gate39inter1), .O(G356));
nand2 gate40( .a(G28), .b(G32), .O(G359) );
nand2 gate41( .a(G1), .b(G266), .O(G362) );

  xor2  gate1247(.a(G266), .b(G2), .O(gate42inter0));
  nand2 gate1248(.a(gate42inter0), .b(s_100), .O(gate42inter1));
  and2  gate1249(.a(G266), .b(G2), .O(gate42inter2));
  inv1  gate1250(.a(s_100), .O(gate42inter3));
  inv1  gate1251(.a(s_101), .O(gate42inter4));
  nand2 gate1252(.a(gate42inter4), .b(gate42inter3), .O(gate42inter5));
  nor2  gate1253(.a(gate42inter5), .b(gate42inter2), .O(gate42inter6));
  inv1  gate1254(.a(G2), .O(gate42inter7));
  inv1  gate1255(.a(G266), .O(gate42inter8));
  nand2 gate1256(.a(gate42inter8), .b(gate42inter7), .O(gate42inter9));
  nand2 gate1257(.a(s_101), .b(gate42inter3), .O(gate42inter10));
  nor2  gate1258(.a(gate42inter10), .b(gate42inter9), .O(gate42inter11));
  nor2  gate1259(.a(gate42inter11), .b(gate42inter6), .O(gate42inter12));
  nand2 gate1260(.a(gate42inter12), .b(gate42inter1), .O(G363));
nand2 gate43( .a(G3), .b(G269), .O(G364) );

  xor2  gate1415(.a(G269), .b(G4), .O(gate44inter0));
  nand2 gate1416(.a(gate44inter0), .b(s_124), .O(gate44inter1));
  and2  gate1417(.a(G269), .b(G4), .O(gate44inter2));
  inv1  gate1418(.a(s_124), .O(gate44inter3));
  inv1  gate1419(.a(s_125), .O(gate44inter4));
  nand2 gate1420(.a(gate44inter4), .b(gate44inter3), .O(gate44inter5));
  nor2  gate1421(.a(gate44inter5), .b(gate44inter2), .O(gate44inter6));
  inv1  gate1422(.a(G4), .O(gate44inter7));
  inv1  gate1423(.a(G269), .O(gate44inter8));
  nand2 gate1424(.a(gate44inter8), .b(gate44inter7), .O(gate44inter9));
  nand2 gate1425(.a(s_125), .b(gate44inter3), .O(gate44inter10));
  nor2  gate1426(.a(gate44inter10), .b(gate44inter9), .O(gate44inter11));
  nor2  gate1427(.a(gate44inter11), .b(gate44inter6), .O(gate44inter12));
  nand2 gate1428(.a(gate44inter12), .b(gate44inter1), .O(G365));
nand2 gate45( .a(G5), .b(G272), .O(G366) );

  xor2  gate1569(.a(G272), .b(G6), .O(gate46inter0));
  nand2 gate1570(.a(gate46inter0), .b(s_146), .O(gate46inter1));
  and2  gate1571(.a(G272), .b(G6), .O(gate46inter2));
  inv1  gate1572(.a(s_146), .O(gate46inter3));
  inv1  gate1573(.a(s_147), .O(gate46inter4));
  nand2 gate1574(.a(gate46inter4), .b(gate46inter3), .O(gate46inter5));
  nor2  gate1575(.a(gate46inter5), .b(gate46inter2), .O(gate46inter6));
  inv1  gate1576(.a(G6), .O(gate46inter7));
  inv1  gate1577(.a(G272), .O(gate46inter8));
  nand2 gate1578(.a(gate46inter8), .b(gate46inter7), .O(gate46inter9));
  nand2 gate1579(.a(s_147), .b(gate46inter3), .O(gate46inter10));
  nor2  gate1580(.a(gate46inter10), .b(gate46inter9), .O(gate46inter11));
  nor2  gate1581(.a(gate46inter11), .b(gate46inter6), .O(gate46inter12));
  nand2 gate1582(.a(gate46inter12), .b(gate46inter1), .O(G367));
nand2 gate47( .a(G7), .b(G275), .O(G368) );

  xor2  gate1555(.a(G275), .b(G8), .O(gate48inter0));
  nand2 gate1556(.a(gate48inter0), .b(s_144), .O(gate48inter1));
  and2  gate1557(.a(G275), .b(G8), .O(gate48inter2));
  inv1  gate1558(.a(s_144), .O(gate48inter3));
  inv1  gate1559(.a(s_145), .O(gate48inter4));
  nand2 gate1560(.a(gate48inter4), .b(gate48inter3), .O(gate48inter5));
  nor2  gate1561(.a(gate48inter5), .b(gate48inter2), .O(gate48inter6));
  inv1  gate1562(.a(G8), .O(gate48inter7));
  inv1  gate1563(.a(G275), .O(gate48inter8));
  nand2 gate1564(.a(gate48inter8), .b(gate48inter7), .O(gate48inter9));
  nand2 gate1565(.a(s_145), .b(gate48inter3), .O(gate48inter10));
  nor2  gate1566(.a(gate48inter10), .b(gate48inter9), .O(gate48inter11));
  nor2  gate1567(.a(gate48inter11), .b(gate48inter6), .O(gate48inter12));
  nand2 gate1568(.a(gate48inter12), .b(gate48inter1), .O(G369));
nand2 gate49( .a(G9), .b(G278), .O(G370) );

  xor2  gate2647(.a(G278), .b(G10), .O(gate50inter0));
  nand2 gate2648(.a(gate50inter0), .b(s_300), .O(gate50inter1));
  and2  gate2649(.a(G278), .b(G10), .O(gate50inter2));
  inv1  gate2650(.a(s_300), .O(gate50inter3));
  inv1  gate2651(.a(s_301), .O(gate50inter4));
  nand2 gate2652(.a(gate50inter4), .b(gate50inter3), .O(gate50inter5));
  nor2  gate2653(.a(gate50inter5), .b(gate50inter2), .O(gate50inter6));
  inv1  gate2654(.a(G10), .O(gate50inter7));
  inv1  gate2655(.a(G278), .O(gate50inter8));
  nand2 gate2656(.a(gate50inter8), .b(gate50inter7), .O(gate50inter9));
  nand2 gate2657(.a(s_301), .b(gate50inter3), .O(gate50inter10));
  nor2  gate2658(.a(gate50inter10), .b(gate50inter9), .O(gate50inter11));
  nor2  gate2659(.a(gate50inter11), .b(gate50inter6), .O(gate50inter12));
  nand2 gate2660(.a(gate50inter12), .b(gate50inter1), .O(G371));

  xor2  gate1093(.a(G281), .b(G11), .O(gate51inter0));
  nand2 gate1094(.a(gate51inter0), .b(s_78), .O(gate51inter1));
  and2  gate1095(.a(G281), .b(G11), .O(gate51inter2));
  inv1  gate1096(.a(s_78), .O(gate51inter3));
  inv1  gate1097(.a(s_79), .O(gate51inter4));
  nand2 gate1098(.a(gate51inter4), .b(gate51inter3), .O(gate51inter5));
  nor2  gate1099(.a(gate51inter5), .b(gate51inter2), .O(gate51inter6));
  inv1  gate1100(.a(G11), .O(gate51inter7));
  inv1  gate1101(.a(G281), .O(gate51inter8));
  nand2 gate1102(.a(gate51inter8), .b(gate51inter7), .O(gate51inter9));
  nand2 gate1103(.a(s_79), .b(gate51inter3), .O(gate51inter10));
  nor2  gate1104(.a(gate51inter10), .b(gate51inter9), .O(gate51inter11));
  nor2  gate1105(.a(gate51inter11), .b(gate51inter6), .O(gate51inter12));
  nand2 gate1106(.a(gate51inter12), .b(gate51inter1), .O(G372));
nand2 gate52( .a(G12), .b(G281), .O(G373) );
nand2 gate53( .a(G13), .b(G284), .O(G374) );
nand2 gate54( .a(G14), .b(G284), .O(G375) );
nand2 gate55( .a(G15), .b(G287), .O(G376) );

  xor2  gate2073(.a(G287), .b(G16), .O(gate56inter0));
  nand2 gate2074(.a(gate56inter0), .b(s_218), .O(gate56inter1));
  and2  gate2075(.a(G287), .b(G16), .O(gate56inter2));
  inv1  gate2076(.a(s_218), .O(gate56inter3));
  inv1  gate2077(.a(s_219), .O(gate56inter4));
  nand2 gate2078(.a(gate56inter4), .b(gate56inter3), .O(gate56inter5));
  nor2  gate2079(.a(gate56inter5), .b(gate56inter2), .O(gate56inter6));
  inv1  gate2080(.a(G16), .O(gate56inter7));
  inv1  gate2081(.a(G287), .O(gate56inter8));
  nand2 gate2082(.a(gate56inter8), .b(gate56inter7), .O(gate56inter9));
  nand2 gate2083(.a(s_219), .b(gate56inter3), .O(gate56inter10));
  nor2  gate2084(.a(gate56inter10), .b(gate56inter9), .O(gate56inter11));
  nor2  gate2085(.a(gate56inter11), .b(gate56inter6), .O(gate56inter12));
  nand2 gate2086(.a(gate56inter12), .b(gate56inter1), .O(G377));
nand2 gate57( .a(G17), .b(G290), .O(G378) );
nand2 gate58( .a(G18), .b(G290), .O(G379) );
nand2 gate59( .a(G19), .b(G293), .O(G380) );
nand2 gate60( .a(G20), .b(G293), .O(G381) );
nand2 gate61( .a(G21), .b(G296), .O(G382) );
nand2 gate62( .a(G22), .b(G296), .O(G383) );

  xor2  gate1653(.a(G299), .b(G23), .O(gate63inter0));
  nand2 gate1654(.a(gate63inter0), .b(s_158), .O(gate63inter1));
  and2  gate1655(.a(G299), .b(G23), .O(gate63inter2));
  inv1  gate1656(.a(s_158), .O(gate63inter3));
  inv1  gate1657(.a(s_159), .O(gate63inter4));
  nand2 gate1658(.a(gate63inter4), .b(gate63inter3), .O(gate63inter5));
  nor2  gate1659(.a(gate63inter5), .b(gate63inter2), .O(gate63inter6));
  inv1  gate1660(.a(G23), .O(gate63inter7));
  inv1  gate1661(.a(G299), .O(gate63inter8));
  nand2 gate1662(.a(gate63inter8), .b(gate63inter7), .O(gate63inter9));
  nand2 gate1663(.a(s_159), .b(gate63inter3), .O(gate63inter10));
  nor2  gate1664(.a(gate63inter10), .b(gate63inter9), .O(gate63inter11));
  nor2  gate1665(.a(gate63inter11), .b(gate63inter6), .O(gate63inter12));
  nand2 gate1666(.a(gate63inter12), .b(gate63inter1), .O(G384));
nand2 gate64( .a(G24), .b(G299), .O(G385) );
nand2 gate65( .a(G25), .b(G302), .O(G386) );
nand2 gate66( .a(G26), .b(G302), .O(G387) );

  xor2  gate3011(.a(G305), .b(G27), .O(gate67inter0));
  nand2 gate3012(.a(gate67inter0), .b(s_352), .O(gate67inter1));
  and2  gate3013(.a(G305), .b(G27), .O(gate67inter2));
  inv1  gate3014(.a(s_352), .O(gate67inter3));
  inv1  gate3015(.a(s_353), .O(gate67inter4));
  nand2 gate3016(.a(gate67inter4), .b(gate67inter3), .O(gate67inter5));
  nor2  gate3017(.a(gate67inter5), .b(gate67inter2), .O(gate67inter6));
  inv1  gate3018(.a(G27), .O(gate67inter7));
  inv1  gate3019(.a(G305), .O(gate67inter8));
  nand2 gate3020(.a(gate67inter8), .b(gate67inter7), .O(gate67inter9));
  nand2 gate3021(.a(s_353), .b(gate67inter3), .O(gate67inter10));
  nor2  gate3022(.a(gate67inter10), .b(gate67inter9), .O(gate67inter11));
  nor2  gate3023(.a(gate67inter11), .b(gate67inter6), .O(gate67inter12));
  nand2 gate3024(.a(gate67inter12), .b(gate67inter1), .O(G388));

  xor2  gate981(.a(G305), .b(G28), .O(gate68inter0));
  nand2 gate982(.a(gate68inter0), .b(s_62), .O(gate68inter1));
  and2  gate983(.a(G305), .b(G28), .O(gate68inter2));
  inv1  gate984(.a(s_62), .O(gate68inter3));
  inv1  gate985(.a(s_63), .O(gate68inter4));
  nand2 gate986(.a(gate68inter4), .b(gate68inter3), .O(gate68inter5));
  nor2  gate987(.a(gate68inter5), .b(gate68inter2), .O(gate68inter6));
  inv1  gate988(.a(G28), .O(gate68inter7));
  inv1  gate989(.a(G305), .O(gate68inter8));
  nand2 gate990(.a(gate68inter8), .b(gate68inter7), .O(gate68inter9));
  nand2 gate991(.a(s_63), .b(gate68inter3), .O(gate68inter10));
  nor2  gate992(.a(gate68inter10), .b(gate68inter9), .O(gate68inter11));
  nor2  gate993(.a(gate68inter11), .b(gate68inter6), .O(gate68inter12));
  nand2 gate994(.a(gate68inter12), .b(gate68inter1), .O(G389));
nand2 gate69( .a(G29), .b(G308), .O(G390) );

  xor2  gate2395(.a(G308), .b(G30), .O(gate70inter0));
  nand2 gate2396(.a(gate70inter0), .b(s_264), .O(gate70inter1));
  and2  gate2397(.a(G308), .b(G30), .O(gate70inter2));
  inv1  gate2398(.a(s_264), .O(gate70inter3));
  inv1  gate2399(.a(s_265), .O(gate70inter4));
  nand2 gate2400(.a(gate70inter4), .b(gate70inter3), .O(gate70inter5));
  nor2  gate2401(.a(gate70inter5), .b(gate70inter2), .O(gate70inter6));
  inv1  gate2402(.a(G30), .O(gate70inter7));
  inv1  gate2403(.a(G308), .O(gate70inter8));
  nand2 gate2404(.a(gate70inter8), .b(gate70inter7), .O(gate70inter9));
  nand2 gate2405(.a(s_265), .b(gate70inter3), .O(gate70inter10));
  nor2  gate2406(.a(gate70inter10), .b(gate70inter9), .O(gate70inter11));
  nor2  gate2407(.a(gate70inter11), .b(gate70inter6), .O(gate70inter12));
  nand2 gate2408(.a(gate70inter12), .b(gate70inter1), .O(G391));
nand2 gate71( .a(G31), .b(G311), .O(G392) );
nand2 gate72( .a(G32), .b(G311), .O(G393) );
nand2 gate73( .a(G1), .b(G314), .O(G394) );
nand2 gate74( .a(G5), .b(G314), .O(G395) );
nand2 gate75( .a(G9), .b(G317), .O(G396) );

  xor2  gate2087(.a(G317), .b(G13), .O(gate76inter0));
  nand2 gate2088(.a(gate76inter0), .b(s_220), .O(gate76inter1));
  and2  gate2089(.a(G317), .b(G13), .O(gate76inter2));
  inv1  gate2090(.a(s_220), .O(gate76inter3));
  inv1  gate2091(.a(s_221), .O(gate76inter4));
  nand2 gate2092(.a(gate76inter4), .b(gate76inter3), .O(gate76inter5));
  nor2  gate2093(.a(gate76inter5), .b(gate76inter2), .O(gate76inter6));
  inv1  gate2094(.a(G13), .O(gate76inter7));
  inv1  gate2095(.a(G317), .O(gate76inter8));
  nand2 gate2096(.a(gate76inter8), .b(gate76inter7), .O(gate76inter9));
  nand2 gate2097(.a(s_221), .b(gate76inter3), .O(gate76inter10));
  nor2  gate2098(.a(gate76inter10), .b(gate76inter9), .O(gate76inter11));
  nor2  gate2099(.a(gate76inter11), .b(gate76inter6), .O(gate76inter12));
  nand2 gate2100(.a(gate76inter12), .b(gate76inter1), .O(G397));
nand2 gate77( .a(G2), .b(G320), .O(G398) );

  xor2  gate2675(.a(G320), .b(G6), .O(gate78inter0));
  nand2 gate2676(.a(gate78inter0), .b(s_304), .O(gate78inter1));
  and2  gate2677(.a(G320), .b(G6), .O(gate78inter2));
  inv1  gate2678(.a(s_304), .O(gate78inter3));
  inv1  gate2679(.a(s_305), .O(gate78inter4));
  nand2 gate2680(.a(gate78inter4), .b(gate78inter3), .O(gate78inter5));
  nor2  gate2681(.a(gate78inter5), .b(gate78inter2), .O(gate78inter6));
  inv1  gate2682(.a(G6), .O(gate78inter7));
  inv1  gate2683(.a(G320), .O(gate78inter8));
  nand2 gate2684(.a(gate78inter8), .b(gate78inter7), .O(gate78inter9));
  nand2 gate2685(.a(s_305), .b(gate78inter3), .O(gate78inter10));
  nor2  gate2686(.a(gate78inter10), .b(gate78inter9), .O(gate78inter11));
  nor2  gate2687(.a(gate78inter11), .b(gate78inter6), .O(gate78inter12));
  nand2 gate2688(.a(gate78inter12), .b(gate78inter1), .O(G399));

  xor2  gate673(.a(G323), .b(G10), .O(gate79inter0));
  nand2 gate674(.a(gate79inter0), .b(s_18), .O(gate79inter1));
  and2  gate675(.a(G323), .b(G10), .O(gate79inter2));
  inv1  gate676(.a(s_18), .O(gate79inter3));
  inv1  gate677(.a(s_19), .O(gate79inter4));
  nand2 gate678(.a(gate79inter4), .b(gate79inter3), .O(gate79inter5));
  nor2  gate679(.a(gate79inter5), .b(gate79inter2), .O(gate79inter6));
  inv1  gate680(.a(G10), .O(gate79inter7));
  inv1  gate681(.a(G323), .O(gate79inter8));
  nand2 gate682(.a(gate79inter8), .b(gate79inter7), .O(gate79inter9));
  nand2 gate683(.a(s_19), .b(gate79inter3), .O(gate79inter10));
  nor2  gate684(.a(gate79inter10), .b(gate79inter9), .O(gate79inter11));
  nor2  gate685(.a(gate79inter11), .b(gate79inter6), .O(gate79inter12));
  nand2 gate686(.a(gate79inter12), .b(gate79inter1), .O(G400));
nand2 gate80( .a(G14), .b(G323), .O(G401) );

  xor2  gate1821(.a(G326), .b(G3), .O(gate81inter0));
  nand2 gate1822(.a(gate81inter0), .b(s_182), .O(gate81inter1));
  and2  gate1823(.a(G326), .b(G3), .O(gate81inter2));
  inv1  gate1824(.a(s_182), .O(gate81inter3));
  inv1  gate1825(.a(s_183), .O(gate81inter4));
  nand2 gate1826(.a(gate81inter4), .b(gate81inter3), .O(gate81inter5));
  nor2  gate1827(.a(gate81inter5), .b(gate81inter2), .O(gate81inter6));
  inv1  gate1828(.a(G3), .O(gate81inter7));
  inv1  gate1829(.a(G326), .O(gate81inter8));
  nand2 gate1830(.a(gate81inter8), .b(gate81inter7), .O(gate81inter9));
  nand2 gate1831(.a(s_183), .b(gate81inter3), .O(gate81inter10));
  nor2  gate1832(.a(gate81inter10), .b(gate81inter9), .O(gate81inter11));
  nor2  gate1833(.a(gate81inter11), .b(gate81inter6), .O(gate81inter12));
  nand2 gate1834(.a(gate81inter12), .b(gate81inter1), .O(G402));

  xor2  gate2703(.a(G326), .b(G7), .O(gate82inter0));
  nand2 gate2704(.a(gate82inter0), .b(s_308), .O(gate82inter1));
  and2  gate2705(.a(G326), .b(G7), .O(gate82inter2));
  inv1  gate2706(.a(s_308), .O(gate82inter3));
  inv1  gate2707(.a(s_309), .O(gate82inter4));
  nand2 gate2708(.a(gate82inter4), .b(gate82inter3), .O(gate82inter5));
  nor2  gate2709(.a(gate82inter5), .b(gate82inter2), .O(gate82inter6));
  inv1  gate2710(.a(G7), .O(gate82inter7));
  inv1  gate2711(.a(G326), .O(gate82inter8));
  nand2 gate2712(.a(gate82inter8), .b(gate82inter7), .O(gate82inter9));
  nand2 gate2713(.a(s_309), .b(gate82inter3), .O(gate82inter10));
  nor2  gate2714(.a(gate82inter10), .b(gate82inter9), .O(gate82inter11));
  nor2  gate2715(.a(gate82inter11), .b(gate82inter6), .O(gate82inter12));
  nand2 gate2716(.a(gate82inter12), .b(gate82inter1), .O(G403));
nand2 gate83( .a(G11), .b(G329), .O(G404) );

  xor2  gate1373(.a(G329), .b(G15), .O(gate84inter0));
  nand2 gate1374(.a(gate84inter0), .b(s_118), .O(gate84inter1));
  and2  gate1375(.a(G329), .b(G15), .O(gate84inter2));
  inv1  gate1376(.a(s_118), .O(gate84inter3));
  inv1  gate1377(.a(s_119), .O(gate84inter4));
  nand2 gate1378(.a(gate84inter4), .b(gate84inter3), .O(gate84inter5));
  nor2  gate1379(.a(gate84inter5), .b(gate84inter2), .O(gate84inter6));
  inv1  gate1380(.a(G15), .O(gate84inter7));
  inv1  gate1381(.a(G329), .O(gate84inter8));
  nand2 gate1382(.a(gate84inter8), .b(gate84inter7), .O(gate84inter9));
  nand2 gate1383(.a(s_119), .b(gate84inter3), .O(gate84inter10));
  nor2  gate1384(.a(gate84inter10), .b(gate84inter9), .O(gate84inter11));
  nor2  gate1385(.a(gate84inter11), .b(gate84inter6), .O(gate84inter12));
  nand2 gate1386(.a(gate84inter12), .b(gate84inter1), .O(G405));

  xor2  gate2423(.a(G332), .b(G4), .O(gate85inter0));
  nand2 gate2424(.a(gate85inter0), .b(s_268), .O(gate85inter1));
  and2  gate2425(.a(G332), .b(G4), .O(gate85inter2));
  inv1  gate2426(.a(s_268), .O(gate85inter3));
  inv1  gate2427(.a(s_269), .O(gate85inter4));
  nand2 gate2428(.a(gate85inter4), .b(gate85inter3), .O(gate85inter5));
  nor2  gate2429(.a(gate85inter5), .b(gate85inter2), .O(gate85inter6));
  inv1  gate2430(.a(G4), .O(gate85inter7));
  inv1  gate2431(.a(G332), .O(gate85inter8));
  nand2 gate2432(.a(gate85inter8), .b(gate85inter7), .O(gate85inter9));
  nand2 gate2433(.a(s_269), .b(gate85inter3), .O(gate85inter10));
  nor2  gate2434(.a(gate85inter10), .b(gate85inter9), .O(gate85inter11));
  nor2  gate2435(.a(gate85inter11), .b(gate85inter6), .O(gate85inter12));
  nand2 gate2436(.a(gate85inter12), .b(gate85inter1), .O(G406));

  xor2  gate575(.a(G332), .b(G8), .O(gate86inter0));
  nand2 gate576(.a(gate86inter0), .b(s_4), .O(gate86inter1));
  and2  gate577(.a(G332), .b(G8), .O(gate86inter2));
  inv1  gate578(.a(s_4), .O(gate86inter3));
  inv1  gate579(.a(s_5), .O(gate86inter4));
  nand2 gate580(.a(gate86inter4), .b(gate86inter3), .O(gate86inter5));
  nor2  gate581(.a(gate86inter5), .b(gate86inter2), .O(gate86inter6));
  inv1  gate582(.a(G8), .O(gate86inter7));
  inv1  gate583(.a(G332), .O(gate86inter8));
  nand2 gate584(.a(gate86inter8), .b(gate86inter7), .O(gate86inter9));
  nand2 gate585(.a(s_5), .b(gate86inter3), .O(gate86inter10));
  nor2  gate586(.a(gate86inter10), .b(gate86inter9), .O(gate86inter11));
  nor2  gate587(.a(gate86inter11), .b(gate86inter6), .O(gate86inter12));
  nand2 gate588(.a(gate86inter12), .b(gate86inter1), .O(G407));
nand2 gate87( .a(G12), .b(G335), .O(G408) );
nand2 gate88( .a(G16), .b(G335), .O(G409) );

  xor2  gate3081(.a(G338), .b(G17), .O(gate89inter0));
  nand2 gate3082(.a(gate89inter0), .b(s_362), .O(gate89inter1));
  and2  gate3083(.a(G338), .b(G17), .O(gate89inter2));
  inv1  gate3084(.a(s_362), .O(gate89inter3));
  inv1  gate3085(.a(s_363), .O(gate89inter4));
  nand2 gate3086(.a(gate89inter4), .b(gate89inter3), .O(gate89inter5));
  nor2  gate3087(.a(gate89inter5), .b(gate89inter2), .O(gate89inter6));
  inv1  gate3088(.a(G17), .O(gate89inter7));
  inv1  gate3089(.a(G338), .O(gate89inter8));
  nand2 gate3090(.a(gate89inter8), .b(gate89inter7), .O(gate89inter9));
  nand2 gate3091(.a(s_363), .b(gate89inter3), .O(gate89inter10));
  nor2  gate3092(.a(gate89inter10), .b(gate89inter9), .O(gate89inter11));
  nor2  gate3093(.a(gate89inter11), .b(gate89inter6), .O(gate89inter12));
  nand2 gate3094(.a(gate89inter12), .b(gate89inter1), .O(G410));
nand2 gate90( .a(G21), .b(G338), .O(G411) );

  xor2  gate2381(.a(G341), .b(G25), .O(gate91inter0));
  nand2 gate2382(.a(gate91inter0), .b(s_262), .O(gate91inter1));
  and2  gate2383(.a(G341), .b(G25), .O(gate91inter2));
  inv1  gate2384(.a(s_262), .O(gate91inter3));
  inv1  gate2385(.a(s_263), .O(gate91inter4));
  nand2 gate2386(.a(gate91inter4), .b(gate91inter3), .O(gate91inter5));
  nor2  gate2387(.a(gate91inter5), .b(gate91inter2), .O(gate91inter6));
  inv1  gate2388(.a(G25), .O(gate91inter7));
  inv1  gate2389(.a(G341), .O(gate91inter8));
  nand2 gate2390(.a(gate91inter8), .b(gate91inter7), .O(gate91inter9));
  nand2 gate2391(.a(s_263), .b(gate91inter3), .O(gate91inter10));
  nor2  gate2392(.a(gate91inter10), .b(gate91inter9), .O(gate91inter11));
  nor2  gate2393(.a(gate91inter11), .b(gate91inter6), .O(gate91inter12));
  nand2 gate2394(.a(gate91inter12), .b(gate91inter1), .O(G412));

  xor2  gate1261(.a(G341), .b(G29), .O(gate92inter0));
  nand2 gate1262(.a(gate92inter0), .b(s_102), .O(gate92inter1));
  and2  gate1263(.a(G341), .b(G29), .O(gate92inter2));
  inv1  gate1264(.a(s_102), .O(gate92inter3));
  inv1  gate1265(.a(s_103), .O(gate92inter4));
  nand2 gate1266(.a(gate92inter4), .b(gate92inter3), .O(gate92inter5));
  nor2  gate1267(.a(gate92inter5), .b(gate92inter2), .O(gate92inter6));
  inv1  gate1268(.a(G29), .O(gate92inter7));
  inv1  gate1269(.a(G341), .O(gate92inter8));
  nand2 gate1270(.a(gate92inter8), .b(gate92inter7), .O(gate92inter9));
  nand2 gate1271(.a(s_103), .b(gate92inter3), .O(gate92inter10));
  nor2  gate1272(.a(gate92inter10), .b(gate92inter9), .O(gate92inter11));
  nor2  gate1273(.a(gate92inter11), .b(gate92inter6), .O(gate92inter12));
  nand2 gate1274(.a(gate92inter12), .b(gate92inter1), .O(G413));
nand2 gate93( .a(G18), .b(G344), .O(G414) );

  xor2  gate1009(.a(G344), .b(G22), .O(gate94inter0));
  nand2 gate1010(.a(gate94inter0), .b(s_66), .O(gate94inter1));
  and2  gate1011(.a(G344), .b(G22), .O(gate94inter2));
  inv1  gate1012(.a(s_66), .O(gate94inter3));
  inv1  gate1013(.a(s_67), .O(gate94inter4));
  nand2 gate1014(.a(gate94inter4), .b(gate94inter3), .O(gate94inter5));
  nor2  gate1015(.a(gate94inter5), .b(gate94inter2), .O(gate94inter6));
  inv1  gate1016(.a(G22), .O(gate94inter7));
  inv1  gate1017(.a(G344), .O(gate94inter8));
  nand2 gate1018(.a(gate94inter8), .b(gate94inter7), .O(gate94inter9));
  nand2 gate1019(.a(s_67), .b(gate94inter3), .O(gate94inter10));
  nor2  gate1020(.a(gate94inter10), .b(gate94inter9), .O(gate94inter11));
  nor2  gate1021(.a(gate94inter11), .b(gate94inter6), .O(gate94inter12));
  nand2 gate1022(.a(gate94inter12), .b(gate94inter1), .O(G415));
nand2 gate95( .a(G26), .b(G347), .O(G416) );
nand2 gate96( .a(G30), .b(G347), .O(G417) );

  xor2  gate1275(.a(G350), .b(G19), .O(gate97inter0));
  nand2 gate1276(.a(gate97inter0), .b(s_104), .O(gate97inter1));
  and2  gate1277(.a(G350), .b(G19), .O(gate97inter2));
  inv1  gate1278(.a(s_104), .O(gate97inter3));
  inv1  gate1279(.a(s_105), .O(gate97inter4));
  nand2 gate1280(.a(gate97inter4), .b(gate97inter3), .O(gate97inter5));
  nor2  gate1281(.a(gate97inter5), .b(gate97inter2), .O(gate97inter6));
  inv1  gate1282(.a(G19), .O(gate97inter7));
  inv1  gate1283(.a(G350), .O(gate97inter8));
  nand2 gate1284(.a(gate97inter8), .b(gate97inter7), .O(gate97inter9));
  nand2 gate1285(.a(s_105), .b(gate97inter3), .O(gate97inter10));
  nor2  gate1286(.a(gate97inter10), .b(gate97inter9), .O(gate97inter11));
  nor2  gate1287(.a(gate97inter11), .b(gate97inter6), .O(gate97inter12));
  nand2 gate1288(.a(gate97inter12), .b(gate97inter1), .O(G418));

  xor2  gate2577(.a(G350), .b(G23), .O(gate98inter0));
  nand2 gate2578(.a(gate98inter0), .b(s_290), .O(gate98inter1));
  and2  gate2579(.a(G350), .b(G23), .O(gate98inter2));
  inv1  gate2580(.a(s_290), .O(gate98inter3));
  inv1  gate2581(.a(s_291), .O(gate98inter4));
  nand2 gate2582(.a(gate98inter4), .b(gate98inter3), .O(gate98inter5));
  nor2  gate2583(.a(gate98inter5), .b(gate98inter2), .O(gate98inter6));
  inv1  gate2584(.a(G23), .O(gate98inter7));
  inv1  gate2585(.a(G350), .O(gate98inter8));
  nand2 gate2586(.a(gate98inter8), .b(gate98inter7), .O(gate98inter9));
  nand2 gate2587(.a(s_291), .b(gate98inter3), .O(gate98inter10));
  nor2  gate2588(.a(gate98inter10), .b(gate98inter9), .O(gate98inter11));
  nor2  gate2589(.a(gate98inter11), .b(gate98inter6), .O(gate98inter12));
  nand2 gate2590(.a(gate98inter12), .b(gate98inter1), .O(G419));

  xor2  gate1135(.a(G353), .b(G27), .O(gate99inter0));
  nand2 gate1136(.a(gate99inter0), .b(s_84), .O(gate99inter1));
  and2  gate1137(.a(G353), .b(G27), .O(gate99inter2));
  inv1  gate1138(.a(s_84), .O(gate99inter3));
  inv1  gate1139(.a(s_85), .O(gate99inter4));
  nand2 gate1140(.a(gate99inter4), .b(gate99inter3), .O(gate99inter5));
  nor2  gate1141(.a(gate99inter5), .b(gate99inter2), .O(gate99inter6));
  inv1  gate1142(.a(G27), .O(gate99inter7));
  inv1  gate1143(.a(G353), .O(gate99inter8));
  nand2 gate1144(.a(gate99inter8), .b(gate99inter7), .O(gate99inter9));
  nand2 gate1145(.a(s_85), .b(gate99inter3), .O(gate99inter10));
  nor2  gate1146(.a(gate99inter10), .b(gate99inter9), .O(gate99inter11));
  nor2  gate1147(.a(gate99inter11), .b(gate99inter6), .O(gate99inter12));
  nand2 gate1148(.a(gate99inter12), .b(gate99inter1), .O(G420));

  xor2  gate561(.a(G353), .b(G31), .O(gate100inter0));
  nand2 gate562(.a(gate100inter0), .b(s_2), .O(gate100inter1));
  and2  gate563(.a(G353), .b(G31), .O(gate100inter2));
  inv1  gate564(.a(s_2), .O(gate100inter3));
  inv1  gate565(.a(s_3), .O(gate100inter4));
  nand2 gate566(.a(gate100inter4), .b(gate100inter3), .O(gate100inter5));
  nor2  gate567(.a(gate100inter5), .b(gate100inter2), .O(gate100inter6));
  inv1  gate568(.a(G31), .O(gate100inter7));
  inv1  gate569(.a(G353), .O(gate100inter8));
  nand2 gate570(.a(gate100inter8), .b(gate100inter7), .O(gate100inter9));
  nand2 gate571(.a(s_3), .b(gate100inter3), .O(gate100inter10));
  nor2  gate572(.a(gate100inter10), .b(gate100inter9), .O(gate100inter11));
  nor2  gate573(.a(gate100inter11), .b(gate100inter6), .O(gate100inter12));
  nand2 gate574(.a(gate100inter12), .b(gate100inter1), .O(G421));
nand2 gate101( .a(G20), .b(G356), .O(G422) );

  xor2  gate2997(.a(G356), .b(G24), .O(gate102inter0));
  nand2 gate2998(.a(gate102inter0), .b(s_350), .O(gate102inter1));
  and2  gate2999(.a(G356), .b(G24), .O(gate102inter2));
  inv1  gate3000(.a(s_350), .O(gate102inter3));
  inv1  gate3001(.a(s_351), .O(gate102inter4));
  nand2 gate3002(.a(gate102inter4), .b(gate102inter3), .O(gate102inter5));
  nor2  gate3003(.a(gate102inter5), .b(gate102inter2), .O(gate102inter6));
  inv1  gate3004(.a(G24), .O(gate102inter7));
  inv1  gate3005(.a(G356), .O(gate102inter8));
  nand2 gate3006(.a(gate102inter8), .b(gate102inter7), .O(gate102inter9));
  nand2 gate3007(.a(s_351), .b(gate102inter3), .O(gate102inter10));
  nor2  gate3008(.a(gate102inter10), .b(gate102inter9), .O(gate102inter11));
  nor2  gate3009(.a(gate102inter11), .b(gate102inter6), .O(gate102inter12));
  nand2 gate3010(.a(gate102inter12), .b(gate102inter1), .O(G423));

  xor2  gate1191(.a(G359), .b(G28), .O(gate103inter0));
  nand2 gate1192(.a(gate103inter0), .b(s_92), .O(gate103inter1));
  and2  gate1193(.a(G359), .b(G28), .O(gate103inter2));
  inv1  gate1194(.a(s_92), .O(gate103inter3));
  inv1  gate1195(.a(s_93), .O(gate103inter4));
  nand2 gate1196(.a(gate103inter4), .b(gate103inter3), .O(gate103inter5));
  nor2  gate1197(.a(gate103inter5), .b(gate103inter2), .O(gate103inter6));
  inv1  gate1198(.a(G28), .O(gate103inter7));
  inv1  gate1199(.a(G359), .O(gate103inter8));
  nand2 gate1200(.a(gate103inter8), .b(gate103inter7), .O(gate103inter9));
  nand2 gate1201(.a(s_93), .b(gate103inter3), .O(gate103inter10));
  nor2  gate1202(.a(gate103inter10), .b(gate103inter9), .O(gate103inter11));
  nor2  gate1203(.a(gate103inter11), .b(gate103inter6), .O(gate103inter12));
  nand2 gate1204(.a(gate103inter12), .b(gate103inter1), .O(G424));

  xor2  gate2535(.a(G359), .b(G32), .O(gate104inter0));
  nand2 gate2536(.a(gate104inter0), .b(s_284), .O(gate104inter1));
  and2  gate2537(.a(G359), .b(G32), .O(gate104inter2));
  inv1  gate2538(.a(s_284), .O(gate104inter3));
  inv1  gate2539(.a(s_285), .O(gate104inter4));
  nand2 gate2540(.a(gate104inter4), .b(gate104inter3), .O(gate104inter5));
  nor2  gate2541(.a(gate104inter5), .b(gate104inter2), .O(gate104inter6));
  inv1  gate2542(.a(G32), .O(gate104inter7));
  inv1  gate2543(.a(G359), .O(gate104inter8));
  nand2 gate2544(.a(gate104inter8), .b(gate104inter7), .O(gate104inter9));
  nand2 gate2545(.a(s_285), .b(gate104inter3), .O(gate104inter10));
  nor2  gate2546(.a(gate104inter10), .b(gate104inter9), .O(gate104inter11));
  nor2  gate2547(.a(gate104inter11), .b(gate104inter6), .O(gate104inter12));
  nand2 gate2548(.a(gate104inter12), .b(gate104inter1), .O(G425));

  xor2  gate1331(.a(G363), .b(G362), .O(gate105inter0));
  nand2 gate1332(.a(gate105inter0), .b(s_112), .O(gate105inter1));
  and2  gate1333(.a(G363), .b(G362), .O(gate105inter2));
  inv1  gate1334(.a(s_112), .O(gate105inter3));
  inv1  gate1335(.a(s_113), .O(gate105inter4));
  nand2 gate1336(.a(gate105inter4), .b(gate105inter3), .O(gate105inter5));
  nor2  gate1337(.a(gate105inter5), .b(gate105inter2), .O(gate105inter6));
  inv1  gate1338(.a(G362), .O(gate105inter7));
  inv1  gate1339(.a(G363), .O(gate105inter8));
  nand2 gate1340(.a(gate105inter8), .b(gate105inter7), .O(gate105inter9));
  nand2 gate1341(.a(s_113), .b(gate105inter3), .O(gate105inter10));
  nor2  gate1342(.a(gate105inter10), .b(gate105inter9), .O(gate105inter11));
  nor2  gate1343(.a(gate105inter11), .b(gate105inter6), .O(gate105inter12));
  nand2 gate1344(.a(gate105inter12), .b(gate105inter1), .O(G426));

  xor2  gate1849(.a(G365), .b(G364), .O(gate106inter0));
  nand2 gate1850(.a(gate106inter0), .b(s_186), .O(gate106inter1));
  and2  gate1851(.a(G365), .b(G364), .O(gate106inter2));
  inv1  gate1852(.a(s_186), .O(gate106inter3));
  inv1  gate1853(.a(s_187), .O(gate106inter4));
  nand2 gate1854(.a(gate106inter4), .b(gate106inter3), .O(gate106inter5));
  nor2  gate1855(.a(gate106inter5), .b(gate106inter2), .O(gate106inter6));
  inv1  gate1856(.a(G364), .O(gate106inter7));
  inv1  gate1857(.a(G365), .O(gate106inter8));
  nand2 gate1858(.a(gate106inter8), .b(gate106inter7), .O(gate106inter9));
  nand2 gate1859(.a(s_187), .b(gate106inter3), .O(gate106inter10));
  nor2  gate1860(.a(gate106inter10), .b(gate106inter9), .O(gate106inter11));
  nor2  gate1861(.a(gate106inter11), .b(gate106inter6), .O(gate106inter12));
  nand2 gate1862(.a(gate106inter12), .b(gate106inter1), .O(G429));
nand2 gate107( .a(G366), .b(G367), .O(G432) );
nand2 gate108( .a(G368), .b(G369), .O(G435) );
nand2 gate109( .a(G370), .b(G371), .O(G438) );

  xor2  gate883(.a(G373), .b(G372), .O(gate110inter0));
  nand2 gate884(.a(gate110inter0), .b(s_48), .O(gate110inter1));
  and2  gate885(.a(G373), .b(G372), .O(gate110inter2));
  inv1  gate886(.a(s_48), .O(gate110inter3));
  inv1  gate887(.a(s_49), .O(gate110inter4));
  nand2 gate888(.a(gate110inter4), .b(gate110inter3), .O(gate110inter5));
  nor2  gate889(.a(gate110inter5), .b(gate110inter2), .O(gate110inter6));
  inv1  gate890(.a(G372), .O(gate110inter7));
  inv1  gate891(.a(G373), .O(gate110inter8));
  nand2 gate892(.a(gate110inter8), .b(gate110inter7), .O(gate110inter9));
  nand2 gate893(.a(s_49), .b(gate110inter3), .O(gate110inter10));
  nor2  gate894(.a(gate110inter10), .b(gate110inter9), .O(gate110inter11));
  nor2  gate895(.a(gate110inter11), .b(gate110inter6), .O(gate110inter12));
  nand2 gate896(.a(gate110inter12), .b(gate110inter1), .O(G441));

  xor2  gate995(.a(G375), .b(G374), .O(gate111inter0));
  nand2 gate996(.a(gate111inter0), .b(s_64), .O(gate111inter1));
  and2  gate997(.a(G375), .b(G374), .O(gate111inter2));
  inv1  gate998(.a(s_64), .O(gate111inter3));
  inv1  gate999(.a(s_65), .O(gate111inter4));
  nand2 gate1000(.a(gate111inter4), .b(gate111inter3), .O(gate111inter5));
  nor2  gate1001(.a(gate111inter5), .b(gate111inter2), .O(gate111inter6));
  inv1  gate1002(.a(G374), .O(gate111inter7));
  inv1  gate1003(.a(G375), .O(gate111inter8));
  nand2 gate1004(.a(gate111inter8), .b(gate111inter7), .O(gate111inter9));
  nand2 gate1005(.a(s_65), .b(gate111inter3), .O(gate111inter10));
  nor2  gate1006(.a(gate111inter10), .b(gate111inter9), .O(gate111inter11));
  nor2  gate1007(.a(gate111inter11), .b(gate111inter6), .O(gate111inter12));
  nand2 gate1008(.a(gate111inter12), .b(gate111inter1), .O(G444));

  xor2  gate659(.a(G377), .b(G376), .O(gate112inter0));
  nand2 gate660(.a(gate112inter0), .b(s_16), .O(gate112inter1));
  and2  gate661(.a(G377), .b(G376), .O(gate112inter2));
  inv1  gate662(.a(s_16), .O(gate112inter3));
  inv1  gate663(.a(s_17), .O(gate112inter4));
  nand2 gate664(.a(gate112inter4), .b(gate112inter3), .O(gate112inter5));
  nor2  gate665(.a(gate112inter5), .b(gate112inter2), .O(gate112inter6));
  inv1  gate666(.a(G376), .O(gate112inter7));
  inv1  gate667(.a(G377), .O(gate112inter8));
  nand2 gate668(.a(gate112inter8), .b(gate112inter7), .O(gate112inter9));
  nand2 gate669(.a(s_17), .b(gate112inter3), .O(gate112inter10));
  nor2  gate670(.a(gate112inter10), .b(gate112inter9), .O(gate112inter11));
  nor2  gate671(.a(gate112inter11), .b(gate112inter6), .O(gate112inter12));
  nand2 gate672(.a(gate112inter12), .b(gate112inter1), .O(G447));
nand2 gate113( .a(G378), .b(G379), .O(G450) );
nand2 gate114( .a(G380), .b(G381), .O(G453) );

  xor2  gate3039(.a(G383), .b(G382), .O(gate115inter0));
  nand2 gate3040(.a(gate115inter0), .b(s_356), .O(gate115inter1));
  and2  gate3041(.a(G383), .b(G382), .O(gate115inter2));
  inv1  gate3042(.a(s_356), .O(gate115inter3));
  inv1  gate3043(.a(s_357), .O(gate115inter4));
  nand2 gate3044(.a(gate115inter4), .b(gate115inter3), .O(gate115inter5));
  nor2  gate3045(.a(gate115inter5), .b(gate115inter2), .O(gate115inter6));
  inv1  gate3046(.a(G382), .O(gate115inter7));
  inv1  gate3047(.a(G383), .O(gate115inter8));
  nand2 gate3048(.a(gate115inter8), .b(gate115inter7), .O(gate115inter9));
  nand2 gate3049(.a(s_357), .b(gate115inter3), .O(gate115inter10));
  nor2  gate3050(.a(gate115inter10), .b(gate115inter9), .O(gate115inter11));
  nor2  gate3051(.a(gate115inter11), .b(gate115inter6), .O(gate115inter12));
  nand2 gate3052(.a(gate115inter12), .b(gate115inter1), .O(G456));

  xor2  gate2353(.a(G385), .b(G384), .O(gate116inter0));
  nand2 gate2354(.a(gate116inter0), .b(s_258), .O(gate116inter1));
  and2  gate2355(.a(G385), .b(G384), .O(gate116inter2));
  inv1  gate2356(.a(s_258), .O(gate116inter3));
  inv1  gate2357(.a(s_259), .O(gate116inter4));
  nand2 gate2358(.a(gate116inter4), .b(gate116inter3), .O(gate116inter5));
  nor2  gate2359(.a(gate116inter5), .b(gate116inter2), .O(gate116inter6));
  inv1  gate2360(.a(G384), .O(gate116inter7));
  inv1  gate2361(.a(G385), .O(gate116inter8));
  nand2 gate2362(.a(gate116inter8), .b(gate116inter7), .O(gate116inter9));
  nand2 gate2363(.a(s_259), .b(gate116inter3), .O(gate116inter10));
  nor2  gate2364(.a(gate116inter10), .b(gate116inter9), .O(gate116inter11));
  nor2  gate2365(.a(gate116inter11), .b(gate116inter6), .O(gate116inter12));
  nand2 gate2366(.a(gate116inter12), .b(gate116inter1), .O(G459));
nand2 gate117( .a(G386), .b(G387), .O(G462) );

  xor2  gate2437(.a(G389), .b(G388), .O(gate118inter0));
  nand2 gate2438(.a(gate118inter0), .b(s_270), .O(gate118inter1));
  and2  gate2439(.a(G389), .b(G388), .O(gate118inter2));
  inv1  gate2440(.a(s_270), .O(gate118inter3));
  inv1  gate2441(.a(s_271), .O(gate118inter4));
  nand2 gate2442(.a(gate118inter4), .b(gate118inter3), .O(gate118inter5));
  nor2  gate2443(.a(gate118inter5), .b(gate118inter2), .O(gate118inter6));
  inv1  gate2444(.a(G388), .O(gate118inter7));
  inv1  gate2445(.a(G389), .O(gate118inter8));
  nand2 gate2446(.a(gate118inter8), .b(gate118inter7), .O(gate118inter9));
  nand2 gate2447(.a(s_271), .b(gate118inter3), .O(gate118inter10));
  nor2  gate2448(.a(gate118inter10), .b(gate118inter9), .O(gate118inter11));
  nor2  gate2449(.a(gate118inter11), .b(gate118inter6), .O(gate118inter12));
  nand2 gate2450(.a(gate118inter12), .b(gate118inter1), .O(G465));

  xor2  gate799(.a(G391), .b(G390), .O(gate119inter0));
  nand2 gate800(.a(gate119inter0), .b(s_36), .O(gate119inter1));
  and2  gate801(.a(G391), .b(G390), .O(gate119inter2));
  inv1  gate802(.a(s_36), .O(gate119inter3));
  inv1  gate803(.a(s_37), .O(gate119inter4));
  nand2 gate804(.a(gate119inter4), .b(gate119inter3), .O(gate119inter5));
  nor2  gate805(.a(gate119inter5), .b(gate119inter2), .O(gate119inter6));
  inv1  gate806(.a(G390), .O(gate119inter7));
  inv1  gate807(.a(G391), .O(gate119inter8));
  nand2 gate808(.a(gate119inter8), .b(gate119inter7), .O(gate119inter9));
  nand2 gate809(.a(s_37), .b(gate119inter3), .O(gate119inter10));
  nor2  gate810(.a(gate119inter10), .b(gate119inter9), .O(gate119inter11));
  nor2  gate811(.a(gate119inter11), .b(gate119inter6), .O(gate119inter12));
  nand2 gate812(.a(gate119inter12), .b(gate119inter1), .O(G468));
nand2 gate120( .a(G392), .b(G393), .O(G471) );
nand2 gate121( .a(G394), .b(G395), .O(G474) );
nand2 gate122( .a(G396), .b(G397), .O(G477) );
nand2 gate123( .a(G398), .b(G399), .O(G480) );

  xor2  gate1107(.a(G401), .b(G400), .O(gate124inter0));
  nand2 gate1108(.a(gate124inter0), .b(s_80), .O(gate124inter1));
  and2  gate1109(.a(G401), .b(G400), .O(gate124inter2));
  inv1  gate1110(.a(s_80), .O(gate124inter3));
  inv1  gate1111(.a(s_81), .O(gate124inter4));
  nand2 gate1112(.a(gate124inter4), .b(gate124inter3), .O(gate124inter5));
  nor2  gate1113(.a(gate124inter5), .b(gate124inter2), .O(gate124inter6));
  inv1  gate1114(.a(G400), .O(gate124inter7));
  inv1  gate1115(.a(G401), .O(gate124inter8));
  nand2 gate1116(.a(gate124inter8), .b(gate124inter7), .O(gate124inter9));
  nand2 gate1117(.a(s_81), .b(gate124inter3), .O(gate124inter10));
  nor2  gate1118(.a(gate124inter10), .b(gate124inter9), .O(gate124inter11));
  nor2  gate1119(.a(gate124inter11), .b(gate124inter6), .O(gate124inter12));
  nand2 gate1120(.a(gate124inter12), .b(gate124inter1), .O(G483));
nand2 gate125( .a(G402), .b(G403), .O(G486) );

  xor2  gate2549(.a(G405), .b(G404), .O(gate126inter0));
  nand2 gate2550(.a(gate126inter0), .b(s_286), .O(gate126inter1));
  and2  gate2551(.a(G405), .b(G404), .O(gate126inter2));
  inv1  gate2552(.a(s_286), .O(gate126inter3));
  inv1  gate2553(.a(s_287), .O(gate126inter4));
  nand2 gate2554(.a(gate126inter4), .b(gate126inter3), .O(gate126inter5));
  nor2  gate2555(.a(gate126inter5), .b(gate126inter2), .O(gate126inter6));
  inv1  gate2556(.a(G404), .O(gate126inter7));
  inv1  gate2557(.a(G405), .O(gate126inter8));
  nand2 gate2558(.a(gate126inter8), .b(gate126inter7), .O(gate126inter9));
  nand2 gate2559(.a(s_287), .b(gate126inter3), .O(gate126inter10));
  nor2  gate2560(.a(gate126inter10), .b(gate126inter9), .O(gate126inter11));
  nor2  gate2561(.a(gate126inter11), .b(gate126inter6), .O(gate126inter12));
  nand2 gate2562(.a(gate126inter12), .b(gate126inter1), .O(G489));
nand2 gate127( .a(G406), .b(G407), .O(G492) );

  xor2  gate2255(.a(G409), .b(G408), .O(gate128inter0));
  nand2 gate2256(.a(gate128inter0), .b(s_244), .O(gate128inter1));
  and2  gate2257(.a(G409), .b(G408), .O(gate128inter2));
  inv1  gate2258(.a(s_244), .O(gate128inter3));
  inv1  gate2259(.a(s_245), .O(gate128inter4));
  nand2 gate2260(.a(gate128inter4), .b(gate128inter3), .O(gate128inter5));
  nor2  gate2261(.a(gate128inter5), .b(gate128inter2), .O(gate128inter6));
  inv1  gate2262(.a(G408), .O(gate128inter7));
  inv1  gate2263(.a(G409), .O(gate128inter8));
  nand2 gate2264(.a(gate128inter8), .b(gate128inter7), .O(gate128inter9));
  nand2 gate2265(.a(s_245), .b(gate128inter3), .O(gate128inter10));
  nor2  gate2266(.a(gate128inter10), .b(gate128inter9), .O(gate128inter11));
  nor2  gate2267(.a(gate128inter11), .b(gate128inter6), .O(gate128inter12));
  nand2 gate2268(.a(gate128inter12), .b(gate128inter1), .O(G495));

  xor2  gate3025(.a(G411), .b(G410), .O(gate129inter0));
  nand2 gate3026(.a(gate129inter0), .b(s_354), .O(gate129inter1));
  and2  gate3027(.a(G411), .b(G410), .O(gate129inter2));
  inv1  gate3028(.a(s_354), .O(gate129inter3));
  inv1  gate3029(.a(s_355), .O(gate129inter4));
  nand2 gate3030(.a(gate129inter4), .b(gate129inter3), .O(gate129inter5));
  nor2  gate3031(.a(gate129inter5), .b(gate129inter2), .O(gate129inter6));
  inv1  gate3032(.a(G410), .O(gate129inter7));
  inv1  gate3033(.a(G411), .O(gate129inter8));
  nand2 gate3034(.a(gate129inter8), .b(gate129inter7), .O(gate129inter9));
  nand2 gate3035(.a(s_355), .b(gate129inter3), .O(gate129inter10));
  nor2  gate3036(.a(gate129inter10), .b(gate129inter9), .O(gate129inter11));
  nor2  gate3037(.a(gate129inter11), .b(gate129inter6), .O(gate129inter12));
  nand2 gate3038(.a(gate129inter12), .b(gate129inter1), .O(G498));

  xor2  gate1723(.a(G413), .b(G412), .O(gate130inter0));
  nand2 gate1724(.a(gate130inter0), .b(s_168), .O(gate130inter1));
  and2  gate1725(.a(G413), .b(G412), .O(gate130inter2));
  inv1  gate1726(.a(s_168), .O(gate130inter3));
  inv1  gate1727(.a(s_169), .O(gate130inter4));
  nand2 gate1728(.a(gate130inter4), .b(gate130inter3), .O(gate130inter5));
  nor2  gate1729(.a(gate130inter5), .b(gate130inter2), .O(gate130inter6));
  inv1  gate1730(.a(G412), .O(gate130inter7));
  inv1  gate1731(.a(G413), .O(gate130inter8));
  nand2 gate1732(.a(gate130inter8), .b(gate130inter7), .O(gate130inter9));
  nand2 gate1733(.a(s_169), .b(gate130inter3), .O(gate130inter10));
  nor2  gate1734(.a(gate130inter10), .b(gate130inter9), .O(gate130inter11));
  nor2  gate1735(.a(gate130inter11), .b(gate130inter6), .O(gate130inter12));
  nand2 gate1736(.a(gate130inter12), .b(gate130inter1), .O(G501));

  xor2  gate1541(.a(G415), .b(G414), .O(gate131inter0));
  nand2 gate1542(.a(gate131inter0), .b(s_142), .O(gate131inter1));
  and2  gate1543(.a(G415), .b(G414), .O(gate131inter2));
  inv1  gate1544(.a(s_142), .O(gate131inter3));
  inv1  gate1545(.a(s_143), .O(gate131inter4));
  nand2 gate1546(.a(gate131inter4), .b(gate131inter3), .O(gate131inter5));
  nor2  gate1547(.a(gate131inter5), .b(gate131inter2), .O(gate131inter6));
  inv1  gate1548(.a(G414), .O(gate131inter7));
  inv1  gate1549(.a(G415), .O(gate131inter8));
  nand2 gate1550(.a(gate131inter8), .b(gate131inter7), .O(gate131inter9));
  nand2 gate1551(.a(s_143), .b(gate131inter3), .O(gate131inter10));
  nor2  gate1552(.a(gate131inter10), .b(gate131inter9), .O(gate131inter11));
  nor2  gate1553(.a(gate131inter11), .b(gate131inter6), .O(gate131inter12));
  nand2 gate1554(.a(gate131inter12), .b(gate131inter1), .O(G504));
nand2 gate132( .a(G416), .b(G417), .O(G507) );
nand2 gate133( .a(G418), .b(G419), .O(G510) );

  xor2  gate939(.a(G421), .b(G420), .O(gate134inter0));
  nand2 gate940(.a(gate134inter0), .b(s_56), .O(gate134inter1));
  and2  gate941(.a(G421), .b(G420), .O(gate134inter2));
  inv1  gate942(.a(s_56), .O(gate134inter3));
  inv1  gate943(.a(s_57), .O(gate134inter4));
  nand2 gate944(.a(gate134inter4), .b(gate134inter3), .O(gate134inter5));
  nor2  gate945(.a(gate134inter5), .b(gate134inter2), .O(gate134inter6));
  inv1  gate946(.a(G420), .O(gate134inter7));
  inv1  gate947(.a(G421), .O(gate134inter8));
  nand2 gate948(.a(gate134inter8), .b(gate134inter7), .O(gate134inter9));
  nand2 gate949(.a(s_57), .b(gate134inter3), .O(gate134inter10));
  nor2  gate950(.a(gate134inter10), .b(gate134inter9), .O(gate134inter11));
  nor2  gate951(.a(gate134inter11), .b(gate134inter6), .O(gate134inter12));
  nand2 gate952(.a(gate134inter12), .b(gate134inter1), .O(G513));
nand2 gate135( .a(G422), .b(G423), .O(G516) );

  xor2  gate743(.a(G425), .b(G424), .O(gate136inter0));
  nand2 gate744(.a(gate136inter0), .b(s_28), .O(gate136inter1));
  and2  gate745(.a(G425), .b(G424), .O(gate136inter2));
  inv1  gate746(.a(s_28), .O(gate136inter3));
  inv1  gate747(.a(s_29), .O(gate136inter4));
  nand2 gate748(.a(gate136inter4), .b(gate136inter3), .O(gate136inter5));
  nor2  gate749(.a(gate136inter5), .b(gate136inter2), .O(gate136inter6));
  inv1  gate750(.a(G424), .O(gate136inter7));
  inv1  gate751(.a(G425), .O(gate136inter8));
  nand2 gate752(.a(gate136inter8), .b(gate136inter7), .O(gate136inter9));
  nand2 gate753(.a(s_29), .b(gate136inter3), .O(gate136inter10));
  nor2  gate754(.a(gate136inter10), .b(gate136inter9), .O(gate136inter11));
  nor2  gate755(.a(gate136inter11), .b(gate136inter6), .O(gate136inter12));
  nand2 gate756(.a(gate136inter12), .b(gate136inter1), .O(G519));

  xor2  gate1597(.a(G429), .b(G426), .O(gate137inter0));
  nand2 gate1598(.a(gate137inter0), .b(s_150), .O(gate137inter1));
  and2  gate1599(.a(G429), .b(G426), .O(gate137inter2));
  inv1  gate1600(.a(s_150), .O(gate137inter3));
  inv1  gate1601(.a(s_151), .O(gate137inter4));
  nand2 gate1602(.a(gate137inter4), .b(gate137inter3), .O(gate137inter5));
  nor2  gate1603(.a(gate137inter5), .b(gate137inter2), .O(gate137inter6));
  inv1  gate1604(.a(G426), .O(gate137inter7));
  inv1  gate1605(.a(G429), .O(gate137inter8));
  nand2 gate1606(.a(gate137inter8), .b(gate137inter7), .O(gate137inter9));
  nand2 gate1607(.a(s_151), .b(gate137inter3), .O(gate137inter10));
  nor2  gate1608(.a(gate137inter10), .b(gate137inter9), .O(gate137inter11));
  nor2  gate1609(.a(gate137inter11), .b(gate137inter6), .O(gate137inter12));
  nand2 gate1610(.a(gate137inter12), .b(gate137inter1), .O(G522));

  xor2  gate2115(.a(G435), .b(G432), .O(gate138inter0));
  nand2 gate2116(.a(gate138inter0), .b(s_224), .O(gate138inter1));
  and2  gate2117(.a(G435), .b(G432), .O(gate138inter2));
  inv1  gate2118(.a(s_224), .O(gate138inter3));
  inv1  gate2119(.a(s_225), .O(gate138inter4));
  nand2 gate2120(.a(gate138inter4), .b(gate138inter3), .O(gate138inter5));
  nor2  gate2121(.a(gate138inter5), .b(gate138inter2), .O(gate138inter6));
  inv1  gate2122(.a(G432), .O(gate138inter7));
  inv1  gate2123(.a(G435), .O(gate138inter8));
  nand2 gate2124(.a(gate138inter8), .b(gate138inter7), .O(gate138inter9));
  nand2 gate2125(.a(s_225), .b(gate138inter3), .O(gate138inter10));
  nor2  gate2126(.a(gate138inter10), .b(gate138inter9), .O(gate138inter11));
  nor2  gate2127(.a(gate138inter11), .b(gate138inter6), .O(gate138inter12));
  nand2 gate2128(.a(gate138inter12), .b(gate138inter1), .O(G525));
nand2 gate139( .a(G438), .b(G441), .O(G528) );
nand2 gate140( .a(G444), .b(G447), .O(G531) );
nand2 gate141( .a(G450), .b(G453), .O(G534) );
nand2 gate142( .a(G456), .b(G459), .O(G537) );
nand2 gate143( .a(G462), .b(G465), .O(G540) );

  xor2  gate1513(.a(G471), .b(G468), .O(gate144inter0));
  nand2 gate1514(.a(gate144inter0), .b(s_138), .O(gate144inter1));
  and2  gate1515(.a(G471), .b(G468), .O(gate144inter2));
  inv1  gate1516(.a(s_138), .O(gate144inter3));
  inv1  gate1517(.a(s_139), .O(gate144inter4));
  nand2 gate1518(.a(gate144inter4), .b(gate144inter3), .O(gate144inter5));
  nor2  gate1519(.a(gate144inter5), .b(gate144inter2), .O(gate144inter6));
  inv1  gate1520(.a(G468), .O(gate144inter7));
  inv1  gate1521(.a(G471), .O(gate144inter8));
  nand2 gate1522(.a(gate144inter8), .b(gate144inter7), .O(gate144inter9));
  nand2 gate1523(.a(s_139), .b(gate144inter3), .O(gate144inter10));
  nor2  gate1524(.a(gate144inter10), .b(gate144inter9), .O(gate144inter11));
  nor2  gate1525(.a(gate144inter11), .b(gate144inter6), .O(gate144inter12));
  nand2 gate1526(.a(gate144inter12), .b(gate144inter1), .O(G543));
nand2 gate145( .a(G474), .b(G477), .O(G546) );
nand2 gate146( .a(G480), .b(G483), .O(G549) );

  xor2  gate2003(.a(G489), .b(G486), .O(gate147inter0));
  nand2 gate2004(.a(gate147inter0), .b(s_208), .O(gate147inter1));
  and2  gate2005(.a(G489), .b(G486), .O(gate147inter2));
  inv1  gate2006(.a(s_208), .O(gate147inter3));
  inv1  gate2007(.a(s_209), .O(gate147inter4));
  nand2 gate2008(.a(gate147inter4), .b(gate147inter3), .O(gate147inter5));
  nor2  gate2009(.a(gate147inter5), .b(gate147inter2), .O(gate147inter6));
  inv1  gate2010(.a(G486), .O(gate147inter7));
  inv1  gate2011(.a(G489), .O(gate147inter8));
  nand2 gate2012(.a(gate147inter8), .b(gate147inter7), .O(gate147inter9));
  nand2 gate2013(.a(s_209), .b(gate147inter3), .O(gate147inter10));
  nor2  gate2014(.a(gate147inter10), .b(gate147inter9), .O(gate147inter11));
  nor2  gate2015(.a(gate147inter11), .b(gate147inter6), .O(gate147inter12));
  nand2 gate2016(.a(gate147inter12), .b(gate147inter1), .O(G552));
nand2 gate148( .a(G492), .b(G495), .O(G555) );

  xor2  gate2367(.a(G501), .b(G498), .O(gate149inter0));
  nand2 gate2368(.a(gate149inter0), .b(s_260), .O(gate149inter1));
  and2  gate2369(.a(G501), .b(G498), .O(gate149inter2));
  inv1  gate2370(.a(s_260), .O(gate149inter3));
  inv1  gate2371(.a(s_261), .O(gate149inter4));
  nand2 gate2372(.a(gate149inter4), .b(gate149inter3), .O(gate149inter5));
  nor2  gate2373(.a(gate149inter5), .b(gate149inter2), .O(gate149inter6));
  inv1  gate2374(.a(G498), .O(gate149inter7));
  inv1  gate2375(.a(G501), .O(gate149inter8));
  nand2 gate2376(.a(gate149inter8), .b(gate149inter7), .O(gate149inter9));
  nand2 gate2377(.a(s_261), .b(gate149inter3), .O(gate149inter10));
  nor2  gate2378(.a(gate149inter10), .b(gate149inter9), .O(gate149inter11));
  nor2  gate2379(.a(gate149inter11), .b(gate149inter6), .O(gate149inter12));
  nand2 gate2380(.a(gate149inter12), .b(gate149inter1), .O(G558));
nand2 gate150( .a(G504), .b(G507), .O(G561) );
nand2 gate151( .a(G510), .b(G513), .O(G564) );
nand2 gate152( .a(G516), .b(G519), .O(G567) );

  xor2  gate2465(.a(G522), .b(G426), .O(gate153inter0));
  nand2 gate2466(.a(gate153inter0), .b(s_274), .O(gate153inter1));
  and2  gate2467(.a(G522), .b(G426), .O(gate153inter2));
  inv1  gate2468(.a(s_274), .O(gate153inter3));
  inv1  gate2469(.a(s_275), .O(gate153inter4));
  nand2 gate2470(.a(gate153inter4), .b(gate153inter3), .O(gate153inter5));
  nor2  gate2471(.a(gate153inter5), .b(gate153inter2), .O(gate153inter6));
  inv1  gate2472(.a(G426), .O(gate153inter7));
  inv1  gate2473(.a(G522), .O(gate153inter8));
  nand2 gate2474(.a(gate153inter8), .b(gate153inter7), .O(gate153inter9));
  nand2 gate2475(.a(s_275), .b(gate153inter3), .O(gate153inter10));
  nor2  gate2476(.a(gate153inter10), .b(gate153inter9), .O(gate153inter11));
  nor2  gate2477(.a(gate153inter11), .b(gate153inter6), .O(gate153inter12));
  nand2 gate2478(.a(gate153inter12), .b(gate153inter1), .O(G570));
nand2 gate154( .a(G429), .b(G522), .O(G571) );

  xor2  gate2269(.a(G525), .b(G432), .O(gate155inter0));
  nand2 gate2270(.a(gate155inter0), .b(s_246), .O(gate155inter1));
  and2  gate2271(.a(G525), .b(G432), .O(gate155inter2));
  inv1  gate2272(.a(s_246), .O(gate155inter3));
  inv1  gate2273(.a(s_247), .O(gate155inter4));
  nand2 gate2274(.a(gate155inter4), .b(gate155inter3), .O(gate155inter5));
  nor2  gate2275(.a(gate155inter5), .b(gate155inter2), .O(gate155inter6));
  inv1  gate2276(.a(G432), .O(gate155inter7));
  inv1  gate2277(.a(G525), .O(gate155inter8));
  nand2 gate2278(.a(gate155inter8), .b(gate155inter7), .O(gate155inter9));
  nand2 gate2279(.a(s_247), .b(gate155inter3), .O(gate155inter10));
  nor2  gate2280(.a(gate155inter10), .b(gate155inter9), .O(gate155inter11));
  nor2  gate2281(.a(gate155inter11), .b(gate155inter6), .O(gate155inter12));
  nand2 gate2282(.a(gate155inter12), .b(gate155inter1), .O(G572));

  xor2  gate2031(.a(G525), .b(G435), .O(gate156inter0));
  nand2 gate2032(.a(gate156inter0), .b(s_212), .O(gate156inter1));
  and2  gate2033(.a(G525), .b(G435), .O(gate156inter2));
  inv1  gate2034(.a(s_212), .O(gate156inter3));
  inv1  gate2035(.a(s_213), .O(gate156inter4));
  nand2 gate2036(.a(gate156inter4), .b(gate156inter3), .O(gate156inter5));
  nor2  gate2037(.a(gate156inter5), .b(gate156inter2), .O(gate156inter6));
  inv1  gate2038(.a(G435), .O(gate156inter7));
  inv1  gate2039(.a(G525), .O(gate156inter8));
  nand2 gate2040(.a(gate156inter8), .b(gate156inter7), .O(gate156inter9));
  nand2 gate2041(.a(s_213), .b(gate156inter3), .O(gate156inter10));
  nor2  gate2042(.a(gate156inter10), .b(gate156inter9), .O(gate156inter11));
  nor2  gate2043(.a(gate156inter11), .b(gate156inter6), .O(gate156inter12));
  nand2 gate2044(.a(gate156inter12), .b(gate156inter1), .O(G573));
nand2 gate157( .a(G438), .b(G528), .O(G574) );
nand2 gate158( .a(G441), .b(G528), .O(G575) );
nand2 gate159( .a(G444), .b(G531), .O(G576) );
nand2 gate160( .a(G447), .b(G531), .O(G577) );
nand2 gate161( .a(G450), .b(G534), .O(G578) );
nand2 gate162( .a(G453), .b(G534), .O(G579) );

  xor2  gate1863(.a(G537), .b(G456), .O(gate163inter0));
  nand2 gate1864(.a(gate163inter0), .b(s_188), .O(gate163inter1));
  and2  gate1865(.a(G537), .b(G456), .O(gate163inter2));
  inv1  gate1866(.a(s_188), .O(gate163inter3));
  inv1  gate1867(.a(s_189), .O(gate163inter4));
  nand2 gate1868(.a(gate163inter4), .b(gate163inter3), .O(gate163inter5));
  nor2  gate1869(.a(gate163inter5), .b(gate163inter2), .O(gate163inter6));
  inv1  gate1870(.a(G456), .O(gate163inter7));
  inv1  gate1871(.a(G537), .O(gate163inter8));
  nand2 gate1872(.a(gate163inter8), .b(gate163inter7), .O(gate163inter9));
  nand2 gate1873(.a(s_189), .b(gate163inter3), .O(gate163inter10));
  nor2  gate1874(.a(gate163inter10), .b(gate163inter9), .O(gate163inter11));
  nor2  gate1875(.a(gate163inter11), .b(gate163inter6), .O(gate163inter12));
  nand2 gate1876(.a(gate163inter12), .b(gate163inter1), .O(G580));

  xor2  gate1121(.a(G537), .b(G459), .O(gate164inter0));
  nand2 gate1122(.a(gate164inter0), .b(s_82), .O(gate164inter1));
  and2  gate1123(.a(G537), .b(G459), .O(gate164inter2));
  inv1  gate1124(.a(s_82), .O(gate164inter3));
  inv1  gate1125(.a(s_83), .O(gate164inter4));
  nand2 gate1126(.a(gate164inter4), .b(gate164inter3), .O(gate164inter5));
  nor2  gate1127(.a(gate164inter5), .b(gate164inter2), .O(gate164inter6));
  inv1  gate1128(.a(G459), .O(gate164inter7));
  inv1  gate1129(.a(G537), .O(gate164inter8));
  nand2 gate1130(.a(gate164inter8), .b(gate164inter7), .O(gate164inter9));
  nand2 gate1131(.a(s_83), .b(gate164inter3), .O(gate164inter10));
  nor2  gate1132(.a(gate164inter10), .b(gate164inter9), .O(gate164inter11));
  nor2  gate1133(.a(gate164inter11), .b(gate164inter6), .O(gate164inter12));
  nand2 gate1134(.a(gate164inter12), .b(gate164inter1), .O(G581));

  xor2  gate631(.a(G540), .b(G462), .O(gate165inter0));
  nand2 gate632(.a(gate165inter0), .b(s_12), .O(gate165inter1));
  and2  gate633(.a(G540), .b(G462), .O(gate165inter2));
  inv1  gate634(.a(s_12), .O(gate165inter3));
  inv1  gate635(.a(s_13), .O(gate165inter4));
  nand2 gate636(.a(gate165inter4), .b(gate165inter3), .O(gate165inter5));
  nor2  gate637(.a(gate165inter5), .b(gate165inter2), .O(gate165inter6));
  inv1  gate638(.a(G462), .O(gate165inter7));
  inv1  gate639(.a(G540), .O(gate165inter8));
  nand2 gate640(.a(gate165inter8), .b(gate165inter7), .O(gate165inter9));
  nand2 gate641(.a(s_13), .b(gate165inter3), .O(gate165inter10));
  nor2  gate642(.a(gate165inter10), .b(gate165inter9), .O(gate165inter11));
  nor2  gate643(.a(gate165inter11), .b(gate165inter6), .O(gate165inter12));
  nand2 gate644(.a(gate165inter12), .b(gate165inter1), .O(G582));

  xor2  gate1065(.a(G540), .b(G465), .O(gate166inter0));
  nand2 gate1066(.a(gate166inter0), .b(s_74), .O(gate166inter1));
  and2  gate1067(.a(G540), .b(G465), .O(gate166inter2));
  inv1  gate1068(.a(s_74), .O(gate166inter3));
  inv1  gate1069(.a(s_75), .O(gate166inter4));
  nand2 gate1070(.a(gate166inter4), .b(gate166inter3), .O(gate166inter5));
  nor2  gate1071(.a(gate166inter5), .b(gate166inter2), .O(gate166inter6));
  inv1  gate1072(.a(G465), .O(gate166inter7));
  inv1  gate1073(.a(G540), .O(gate166inter8));
  nand2 gate1074(.a(gate166inter8), .b(gate166inter7), .O(gate166inter9));
  nand2 gate1075(.a(s_75), .b(gate166inter3), .O(gate166inter10));
  nor2  gate1076(.a(gate166inter10), .b(gate166inter9), .O(gate166inter11));
  nor2  gate1077(.a(gate166inter11), .b(gate166inter6), .O(gate166inter12));
  nand2 gate1078(.a(gate166inter12), .b(gate166inter1), .O(G583));
nand2 gate167( .a(G468), .b(G543), .O(G584) );
nand2 gate168( .a(G471), .b(G543), .O(G585) );
nand2 gate169( .a(G474), .b(G546), .O(G586) );

  xor2  gate2311(.a(G546), .b(G477), .O(gate170inter0));
  nand2 gate2312(.a(gate170inter0), .b(s_252), .O(gate170inter1));
  and2  gate2313(.a(G546), .b(G477), .O(gate170inter2));
  inv1  gate2314(.a(s_252), .O(gate170inter3));
  inv1  gate2315(.a(s_253), .O(gate170inter4));
  nand2 gate2316(.a(gate170inter4), .b(gate170inter3), .O(gate170inter5));
  nor2  gate2317(.a(gate170inter5), .b(gate170inter2), .O(gate170inter6));
  inv1  gate2318(.a(G477), .O(gate170inter7));
  inv1  gate2319(.a(G546), .O(gate170inter8));
  nand2 gate2320(.a(gate170inter8), .b(gate170inter7), .O(gate170inter9));
  nand2 gate2321(.a(s_253), .b(gate170inter3), .O(gate170inter10));
  nor2  gate2322(.a(gate170inter10), .b(gate170inter9), .O(gate170inter11));
  nor2  gate2323(.a(gate170inter11), .b(gate170inter6), .O(gate170inter12));
  nand2 gate2324(.a(gate170inter12), .b(gate170inter1), .O(G587));
nand2 gate171( .a(G480), .b(G549), .O(G588) );
nand2 gate172( .a(G483), .b(G549), .O(G589) );

  xor2  gate1975(.a(G552), .b(G486), .O(gate173inter0));
  nand2 gate1976(.a(gate173inter0), .b(s_204), .O(gate173inter1));
  and2  gate1977(.a(G552), .b(G486), .O(gate173inter2));
  inv1  gate1978(.a(s_204), .O(gate173inter3));
  inv1  gate1979(.a(s_205), .O(gate173inter4));
  nand2 gate1980(.a(gate173inter4), .b(gate173inter3), .O(gate173inter5));
  nor2  gate1981(.a(gate173inter5), .b(gate173inter2), .O(gate173inter6));
  inv1  gate1982(.a(G486), .O(gate173inter7));
  inv1  gate1983(.a(G552), .O(gate173inter8));
  nand2 gate1984(.a(gate173inter8), .b(gate173inter7), .O(gate173inter9));
  nand2 gate1985(.a(s_205), .b(gate173inter3), .O(gate173inter10));
  nor2  gate1986(.a(gate173inter10), .b(gate173inter9), .O(gate173inter11));
  nor2  gate1987(.a(gate173inter11), .b(gate173inter6), .O(gate173inter12));
  nand2 gate1988(.a(gate173inter12), .b(gate173inter1), .O(G590));
nand2 gate174( .a(G489), .b(G552), .O(G591) );
nand2 gate175( .a(G492), .b(G555), .O(G592) );

  xor2  gate2731(.a(G555), .b(G495), .O(gate176inter0));
  nand2 gate2732(.a(gate176inter0), .b(s_312), .O(gate176inter1));
  and2  gate2733(.a(G555), .b(G495), .O(gate176inter2));
  inv1  gate2734(.a(s_312), .O(gate176inter3));
  inv1  gate2735(.a(s_313), .O(gate176inter4));
  nand2 gate2736(.a(gate176inter4), .b(gate176inter3), .O(gate176inter5));
  nor2  gate2737(.a(gate176inter5), .b(gate176inter2), .O(gate176inter6));
  inv1  gate2738(.a(G495), .O(gate176inter7));
  inv1  gate2739(.a(G555), .O(gate176inter8));
  nand2 gate2740(.a(gate176inter8), .b(gate176inter7), .O(gate176inter9));
  nand2 gate2741(.a(s_313), .b(gate176inter3), .O(gate176inter10));
  nor2  gate2742(.a(gate176inter10), .b(gate176inter9), .O(gate176inter11));
  nor2  gate2743(.a(gate176inter11), .b(gate176inter6), .O(gate176inter12));
  nand2 gate2744(.a(gate176inter12), .b(gate176inter1), .O(G593));
nand2 gate177( .a(G498), .b(G558), .O(G594) );
nand2 gate178( .a(G501), .b(G558), .O(G595) );
nand2 gate179( .a(G504), .b(G561), .O(G596) );

  xor2  gate2829(.a(G561), .b(G507), .O(gate180inter0));
  nand2 gate2830(.a(gate180inter0), .b(s_326), .O(gate180inter1));
  and2  gate2831(.a(G561), .b(G507), .O(gate180inter2));
  inv1  gate2832(.a(s_326), .O(gate180inter3));
  inv1  gate2833(.a(s_327), .O(gate180inter4));
  nand2 gate2834(.a(gate180inter4), .b(gate180inter3), .O(gate180inter5));
  nor2  gate2835(.a(gate180inter5), .b(gate180inter2), .O(gate180inter6));
  inv1  gate2836(.a(G507), .O(gate180inter7));
  inv1  gate2837(.a(G561), .O(gate180inter8));
  nand2 gate2838(.a(gate180inter8), .b(gate180inter7), .O(gate180inter9));
  nand2 gate2839(.a(s_327), .b(gate180inter3), .O(gate180inter10));
  nor2  gate2840(.a(gate180inter10), .b(gate180inter9), .O(gate180inter11));
  nor2  gate2841(.a(gate180inter11), .b(gate180inter6), .O(gate180inter12));
  nand2 gate2842(.a(gate180inter12), .b(gate180inter1), .O(G597));

  xor2  gate1877(.a(G564), .b(G510), .O(gate181inter0));
  nand2 gate1878(.a(gate181inter0), .b(s_190), .O(gate181inter1));
  and2  gate1879(.a(G564), .b(G510), .O(gate181inter2));
  inv1  gate1880(.a(s_190), .O(gate181inter3));
  inv1  gate1881(.a(s_191), .O(gate181inter4));
  nand2 gate1882(.a(gate181inter4), .b(gate181inter3), .O(gate181inter5));
  nor2  gate1883(.a(gate181inter5), .b(gate181inter2), .O(gate181inter6));
  inv1  gate1884(.a(G510), .O(gate181inter7));
  inv1  gate1885(.a(G564), .O(gate181inter8));
  nand2 gate1886(.a(gate181inter8), .b(gate181inter7), .O(gate181inter9));
  nand2 gate1887(.a(s_191), .b(gate181inter3), .O(gate181inter10));
  nor2  gate1888(.a(gate181inter10), .b(gate181inter9), .O(gate181inter11));
  nor2  gate1889(.a(gate181inter11), .b(gate181inter6), .O(gate181inter12));
  nand2 gate1890(.a(gate181inter12), .b(gate181inter1), .O(G598));
nand2 gate182( .a(G513), .b(G564), .O(G599) );
nand2 gate183( .a(G516), .b(G567), .O(G600) );

  xor2  gate1667(.a(G567), .b(G519), .O(gate184inter0));
  nand2 gate1668(.a(gate184inter0), .b(s_160), .O(gate184inter1));
  and2  gate1669(.a(G567), .b(G519), .O(gate184inter2));
  inv1  gate1670(.a(s_160), .O(gate184inter3));
  inv1  gate1671(.a(s_161), .O(gate184inter4));
  nand2 gate1672(.a(gate184inter4), .b(gate184inter3), .O(gate184inter5));
  nor2  gate1673(.a(gate184inter5), .b(gate184inter2), .O(gate184inter6));
  inv1  gate1674(.a(G519), .O(gate184inter7));
  inv1  gate1675(.a(G567), .O(gate184inter8));
  nand2 gate1676(.a(gate184inter8), .b(gate184inter7), .O(gate184inter9));
  nand2 gate1677(.a(s_161), .b(gate184inter3), .O(gate184inter10));
  nor2  gate1678(.a(gate184inter10), .b(gate184inter9), .O(gate184inter11));
  nor2  gate1679(.a(gate184inter11), .b(gate184inter6), .O(gate184inter12));
  nand2 gate1680(.a(gate184inter12), .b(gate184inter1), .O(G601));

  xor2  gate1149(.a(G571), .b(G570), .O(gate185inter0));
  nand2 gate1150(.a(gate185inter0), .b(s_86), .O(gate185inter1));
  and2  gate1151(.a(G571), .b(G570), .O(gate185inter2));
  inv1  gate1152(.a(s_86), .O(gate185inter3));
  inv1  gate1153(.a(s_87), .O(gate185inter4));
  nand2 gate1154(.a(gate185inter4), .b(gate185inter3), .O(gate185inter5));
  nor2  gate1155(.a(gate185inter5), .b(gate185inter2), .O(gate185inter6));
  inv1  gate1156(.a(G570), .O(gate185inter7));
  inv1  gate1157(.a(G571), .O(gate185inter8));
  nand2 gate1158(.a(gate185inter8), .b(gate185inter7), .O(gate185inter9));
  nand2 gate1159(.a(s_87), .b(gate185inter3), .O(gate185inter10));
  nor2  gate1160(.a(gate185inter10), .b(gate185inter9), .O(gate185inter11));
  nor2  gate1161(.a(gate185inter11), .b(gate185inter6), .O(gate185inter12));
  nand2 gate1162(.a(gate185inter12), .b(gate185inter1), .O(G602));
nand2 gate186( .a(G572), .b(G573), .O(G607) );

  xor2  gate1079(.a(G575), .b(G574), .O(gate187inter0));
  nand2 gate1080(.a(gate187inter0), .b(s_76), .O(gate187inter1));
  and2  gate1081(.a(G575), .b(G574), .O(gate187inter2));
  inv1  gate1082(.a(s_76), .O(gate187inter3));
  inv1  gate1083(.a(s_77), .O(gate187inter4));
  nand2 gate1084(.a(gate187inter4), .b(gate187inter3), .O(gate187inter5));
  nor2  gate1085(.a(gate187inter5), .b(gate187inter2), .O(gate187inter6));
  inv1  gate1086(.a(G574), .O(gate187inter7));
  inv1  gate1087(.a(G575), .O(gate187inter8));
  nand2 gate1088(.a(gate187inter8), .b(gate187inter7), .O(gate187inter9));
  nand2 gate1089(.a(s_77), .b(gate187inter3), .O(gate187inter10));
  nor2  gate1090(.a(gate187inter10), .b(gate187inter9), .O(gate187inter11));
  nor2  gate1091(.a(gate187inter11), .b(gate187inter6), .O(gate187inter12));
  nand2 gate1092(.a(gate187inter12), .b(gate187inter1), .O(G612));

  xor2  gate2171(.a(G577), .b(G576), .O(gate188inter0));
  nand2 gate2172(.a(gate188inter0), .b(s_232), .O(gate188inter1));
  and2  gate2173(.a(G577), .b(G576), .O(gate188inter2));
  inv1  gate2174(.a(s_232), .O(gate188inter3));
  inv1  gate2175(.a(s_233), .O(gate188inter4));
  nand2 gate2176(.a(gate188inter4), .b(gate188inter3), .O(gate188inter5));
  nor2  gate2177(.a(gate188inter5), .b(gate188inter2), .O(gate188inter6));
  inv1  gate2178(.a(G576), .O(gate188inter7));
  inv1  gate2179(.a(G577), .O(gate188inter8));
  nand2 gate2180(.a(gate188inter8), .b(gate188inter7), .O(gate188inter9));
  nand2 gate2181(.a(s_233), .b(gate188inter3), .O(gate188inter10));
  nor2  gate2182(.a(gate188inter10), .b(gate188inter9), .O(gate188inter11));
  nor2  gate2183(.a(gate188inter11), .b(gate188inter6), .O(gate188inter12));
  nand2 gate2184(.a(gate188inter12), .b(gate188inter1), .O(G617));

  xor2  gate2241(.a(G579), .b(G578), .O(gate189inter0));
  nand2 gate2242(.a(gate189inter0), .b(s_242), .O(gate189inter1));
  and2  gate2243(.a(G579), .b(G578), .O(gate189inter2));
  inv1  gate2244(.a(s_242), .O(gate189inter3));
  inv1  gate2245(.a(s_243), .O(gate189inter4));
  nand2 gate2246(.a(gate189inter4), .b(gate189inter3), .O(gate189inter5));
  nor2  gate2247(.a(gate189inter5), .b(gate189inter2), .O(gate189inter6));
  inv1  gate2248(.a(G578), .O(gate189inter7));
  inv1  gate2249(.a(G579), .O(gate189inter8));
  nand2 gate2250(.a(gate189inter8), .b(gate189inter7), .O(gate189inter9));
  nand2 gate2251(.a(s_243), .b(gate189inter3), .O(gate189inter10));
  nor2  gate2252(.a(gate189inter10), .b(gate189inter9), .O(gate189inter11));
  nor2  gate2253(.a(gate189inter11), .b(gate189inter6), .O(gate189inter12));
  nand2 gate2254(.a(gate189inter12), .b(gate189inter1), .O(G622));
nand2 gate190( .a(G580), .b(G581), .O(G627) );
nand2 gate191( .a(G582), .b(G583), .O(G632) );
nand2 gate192( .a(G584), .b(G585), .O(G637) );
nand2 gate193( .a(G586), .b(G587), .O(G642) );
nand2 gate194( .a(G588), .b(G589), .O(G645) );

  xor2  gate1919(.a(G591), .b(G590), .O(gate195inter0));
  nand2 gate1920(.a(gate195inter0), .b(s_196), .O(gate195inter1));
  and2  gate1921(.a(G591), .b(G590), .O(gate195inter2));
  inv1  gate1922(.a(s_196), .O(gate195inter3));
  inv1  gate1923(.a(s_197), .O(gate195inter4));
  nand2 gate1924(.a(gate195inter4), .b(gate195inter3), .O(gate195inter5));
  nor2  gate1925(.a(gate195inter5), .b(gate195inter2), .O(gate195inter6));
  inv1  gate1926(.a(G590), .O(gate195inter7));
  inv1  gate1927(.a(G591), .O(gate195inter8));
  nand2 gate1928(.a(gate195inter8), .b(gate195inter7), .O(gate195inter9));
  nand2 gate1929(.a(s_197), .b(gate195inter3), .O(gate195inter10));
  nor2  gate1930(.a(gate195inter10), .b(gate195inter9), .O(gate195inter11));
  nor2  gate1931(.a(gate195inter11), .b(gate195inter6), .O(gate195inter12));
  nand2 gate1932(.a(gate195inter12), .b(gate195inter1), .O(G648));

  xor2  gate2815(.a(G593), .b(G592), .O(gate196inter0));
  nand2 gate2816(.a(gate196inter0), .b(s_324), .O(gate196inter1));
  and2  gate2817(.a(G593), .b(G592), .O(gate196inter2));
  inv1  gate2818(.a(s_324), .O(gate196inter3));
  inv1  gate2819(.a(s_325), .O(gate196inter4));
  nand2 gate2820(.a(gate196inter4), .b(gate196inter3), .O(gate196inter5));
  nor2  gate2821(.a(gate196inter5), .b(gate196inter2), .O(gate196inter6));
  inv1  gate2822(.a(G592), .O(gate196inter7));
  inv1  gate2823(.a(G593), .O(gate196inter8));
  nand2 gate2824(.a(gate196inter8), .b(gate196inter7), .O(gate196inter9));
  nand2 gate2825(.a(s_325), .b(gate196inter3), .O(gate196inter10));
  nor2  gate2826(.a(gate196inter10), .b(gate196inter9), .O(gate196inter11));
  nor2  gate2827(.a(gate196inter11), .b(gate196inter6), .O(gate196inter12));
  nand2 gate2828(.a(gate196inter12), .b(gate196inter1), .O(G651));
nand2 gate197( .a(G594), .b(G595), .O(G654) );

  xor2  gate1205(.a(G597), .b(G596), .O(gate198inter0));
  nand2 gate1206(.a(gate198inter0), .b(s_94), .O(gate198inter1));
  and2  gate1207(.a(G597), .b(G596), .O(gate198inter2));
  inv1  gate1208(.a(s_94), .O(gate198inter3));
  inv1  gate1209(.a(s_95), .O(gate198inter4));
  nand2 gate1210(.a(gate198inter4), .b(gate198inter3), .O(gate198inter5));
  nor2  gate1211(.a(gate198inter5), .b(gate198inter2), .O(gate198inter6));
  inv1  gate1212(.a(G596), .O(gate198inter7));
  inv1  gate1213(.a(G597), .O(gate198inter8));
  nand2 gate1214(.a(gate198inter8), .b(gate198inter7), .O(gate198inter9));
  nand2 gate1215(.a(s_95), .b(gate198inter3), .O(gate198inter10));
  nor2  gate1216(.a(gate198inter10), .b(gate198inter9), .O(gate198inter11));
  nor2  gate1217(.a(gate198inter11), .b(gate198inter6), .O(gate198inter12));
  nand2 gate1218(.a(gate198inter12), .b(gate198inter1), .O(G657));
nand2 gate199( .a(G598), .b(G599), .O(G660) );

  xor2  gate1583(.a(G601), .b(G600), .O(gate200inter0));
  nand2 gate1584(.a(gate200inter0), .b(s_148), .O(gate200inter1));
  and2  gate1585(.a(G601), .b(G600), .O(gate200inter2));
  inv1  gate1586(.a(s_148), .O(gate200inter3));
  inv1  gate1587(.a(s_149), .O(gate200inter4));
  nand2 gate1588(.a(gate200inter4), .b(gate200inter3), .O(gate200inter5));
  nor2  gate1589(.a(gate200inter5), .b(gate200inter2), .O(gate200inter6));
  inv1  gate1590(.a(G600), .O(gate200inter7));
  inv1  gate1591(.a(G601), .O(gate200inter8));
  nand2 gate1592(.a(gate200inter8), .b(gate200inter7), .O(gate200inter9));
  nand2 gate1593(.a(s_149), .b(gate200inter3), .O(gate200inter10));
  nor2  gate1594(.a(gate200inter10), .b(gate200inter9), .O(gate200inter11));
  nor2  gate1595(.a(gate200inter11), .b(gate200inter6), .O(gate200inter12));
  nand2 gate1596(.a(gate200inter12), .b(gate200inter1), .O(G663));

  xor2  gate1625(.a(G607), .b(G602), .O(gate201inter0));
  nand2 gate1626(.a(gate201inter0), .b(s_154), .O(gate201inter1));
  and2  gate1627(.a(G607), .b(G602), .O(gate201inter2));
  inv1  gate1628(.a(s_154), .O(gate201inter3));
  inv1  gate1629(.a(s_155), .O(gate201inter4));
  nand2 gate1630(.a(gate201inter4), .b(gate201inter3), .O(gate201inter5));
  nor2  gate1631(.a(gate201inter5), .b(gate201inter2), .O(gate201inter6));
  inv1  gate1632(.a(G602), .O(gate201inter7));
  inv1  gate1633(.a(G607), .O(gate201inter8));
  nand2 gate1634(.a(gate201inter8), .b(gate201inter7), .O(gate201inter9));
  nand2 gate1635(.a(s_155), .b(gate201inter3), .O(gate201inter10));
  nor2  gate1636(.a(gate201inter10), .b(gate201inter9), .O(gate201inter11));
  nor2  gate1637(.a(gate201inter11), .b(gate201inter6), .O(gate201inter12));
  nand2 gate1638(.a(gate201inter12), .b(gate201inter1), .O(G666));
nand2 gate202( .a(G612), .b(G617), .O(G669) );
nand2 gate203( .a(G602), .b(G612), .O(G672) );
nand2 gate204( .a(G607), .b(G617), .O(G675) );
nand2 gate205( .a(G622), .b(G627), .O(G678) );
nand2 gate206( .a(G632), .b(G637), .O(G681) );

  xor2  gate2605(.a(G632), .b(G622), .O(gate207inter0));
  nand2 gate2606(.a(gate207inter0), .b(s_294), .O(gate207inter1));
  and2  gate2607(.a(G632), .b(G622), .O(gate207inter2));
  inv1  gate2608(.a(s_294), .O(gate207inter3));
  inv1  gate2609(.a(s_295), .O(gate207inter4));
  nand2 gate2610(.a(gate207inter4), .b(gate207inter3), .O(gate207inter5));
  nor2  gate2611(.a(gate207inter5), .b(gate207inter2), .O(gate207inter6));
  inv1  gate2612(.a(G622), .O(gate207inter7));
  inv1  gate2613(.a(G632), .O(gate207inter8));
  nand2 gate2614(.a(gate207inter8), .b(gate207inter7), .O(gate207inter9));
  nand2 gate2615(.a(s_295), .b(gate207inter3), .O(gate207inter10));
  nor2  gate2616(.a(gate207inter10), .b(gate207inter9), .O(gate207inter11));
  nor2  gate2617(.a(gate207inter11), .b(gate207inter6), .O(gate207inter12));
  nand2 gate2618(.a(gate207inter12), .b(gate207inter1), .O(G684));

  xor2  gate2451(.a(G637), .b(G627), .O(gate208inter0));
  nand2 gate2452(.a(gate208inter0), .b(s_272), .O(gate208inter1));
  and2  gate2453(.a(G637), .b(G627), .O(gate208inter2));
  inv1  gate2454(.a(s_272), .O(gate208inter3));
  inv1  gate2455(.a(s_273), .O(gate208inter4));
  nand2 gate2456(.a(gate208inter4), .b(gate208inter3), .O(gate208inter5));
  nor2  gate2457(.a(gate208inter5), .b(gate208inter2), .O(gate208inter6));
  inv1  gate2458(.a(G627), .O(gate208inter7));
  inv1  gate2459(.a(G637), .O(gate208inter8));
  nand2 gate2460(.a(gate208inter8), .b(gate208inter7), .O(gate208inter9));
  nand2 gate2461(.a(s_273), .b(gate208inter3), .O(gate208inter10));
  nor2  gate2462(.a(gate208inter10), .b(gate208inter9), .O(gate208inter11));
  nor2  gate2463(.a(gate208inter11), .b(gate208inter6), .O(gate208inter12));
  nand2 gate2464(.a(gate208inter12), .b(gate208inter1), .O(G687));
nand2 gate209( .a(G602), .b(G666), .O(G690) );

  xor2  gate1471(.a(G666), .b(G607), .O(gate210inter0));
  nand2 gate1472(.a(gate210inter0), .b(s_132), .O(gate210inter1));
  and2  gate1473(.a(G666), .b(G607), .O(gate210inter2));
  inv1  gate1474(.a(s_132), .O(gate210inter3));
  inv1  gate1475(.a(s_133), .O(gate210inter4));
  nand2 gate1476(.a(gate210inter4), .b(gate210inter3), .O(gate210inter5));
  nor2  gate1477(.a(gate210inter5), .b(gate210inter2), .O(gate210inter6));
  inv1  gate1478(.a(G607), .O(gate210inter7));
  inv1  gate1479(.a(G666), .O(gate210inter8));
  nand2 gate1480(.a(gate210inter8), .b(gate210inter7), .O(gate210inter9));
  nand2 gate1481(.a(s_133), .b(gate210inter3), .O(gate210inter10));
  nor2  gate1482(.a(gate210inter10), .b(gate210inter9), .O(gate210inter11));
  nor2  gate1483(.a(gate210inter11), .b(gate210inter6), .O(gate210inter12));
  nand2 gate1484(.a(gate210inter12), .b(gate210inter1), .O(G691));

  xor2  gate547(.a(G669), .b(G612), .O(gate211inter0));
  nand2 gate548(.a(gate211inter0), .b(s_0), .O(gate211inter1));
  and2  gate549(.a(G669), .b(G612), .O(gate211inter2));
  inv1  gate550(.a(s_0), .O(gate211inter3));
  inv1  gate551(.a(s_1), .O(gate211inter4));
  nand2 gate552(.a(gate211inter4), .b(gate211inter3), .O(gate211inter5));
  nor2  gate553(.a(gate211inter5), .b(gate211inter2), .O(gate211inter6));
  inv1  gate554(.a(G612), .O(gate211inter7));
  inv1  gate555(.a(G669), .O(gate211inter8));
  nand2 gate556(.a(gate211inter8), .b(gate211inter7), .O(gate211inter9));
  nand2 gate557(.a(s_1), .b(gate211inter3), .O(gate211inter10));
  nor2  gate558(.a(gate211inter10), .b(gate211inter9), .O(gate211inter11));
  nor2  gate559(.a(gate211inter11), .b(gate211inter6), .O(gate211inter12));
  nand2 gate560(.a(gate211inter12), .b(gate211inter1), .O(G692));

  xor2  gate2045(.a(G669), .b(G617), .O(gate212inter0));
  nand2 gate2046(.a(gate212inter0), .b(s_214), .O(gate212inter1));
  and2  gate2047(.a(G669), .b(G617), .O(gate212inter2));
  inv1  gate2048(.a(s_214), .O(gate212inter3));
  inv1  gate2049(.a(s_215), .O(gate212inter4));
  nand2 gate2050(.a(gate212inter4), .b(gate212inter3), .O(gate212inter5));
  nor2  gate2051(.a(gate212inter5), .b(gate212inter2), .O(gate212inter6));
  inv1  gate2052(.a(G617), .O(gate212inter7));
  inv1  gate2053(.a(G669), .O(gate212inter8));
  nand2 gate2054(.a(gate212inter8), .b(gate212inter7), .O(gate212inter9));
  nand2 gate2055(.a(s_215), .b(gate212inter3), .O(gate212inter10));
  nor2  gate2056(.a(gate212inter10), .b(gate212inter9), .O(gate212inter11));
  nor2  gate2057(.a(gate212inter11), .b(gate212inter6), .O(gate212inter12));
  nand2 gate2058(.a(gate212inter12), .b(gate212inter1), .O(G693));
nand2 gate213( .a(G602), .b(G672), .O(G694) );

  xor2  gate967(.a(G672), .b(G612), .O(gate214inter0));
  nand2 gate968(.a(gate214inter0), .b(s_60), .O(gate214inter1));
  and2  gate969(.a(G672), .b(G612), .O(gate214inter2));
  inv1  gate970(.a(s_60), .O(gate214inter3));
  inv1  gate971(.a(s_61), .O(gate214inter4));
  nand2 gate972(.a(gate214inter4), .b(gate214inter3), .O(gate214inter5));
  nor2  gate973(.a(gate214inter5), .b(gate214inter2), .O(gate214inter6));
  inv1  gate974(.a(G612), .O(gate214inter7));
  inv1  gate975(.a(G672), .O(gate214inter8));
  nand2 gate976(.a(gate214inter8), .b(gate214inter7), .O(gate214inter9));
  nand2 gate977(.a(s_61), .b(gate214inter3), .O(gate214inter10));
  nor2  gate978(.a(gate214inter10), .b(gate214inter9), .O(gate214inter11));
  nor2  gate979(.a(gate214inter11), .b(gate214inter6), .O(gate214inter12));
  nand2 gate980(.a(gate214inter12), .b(gate214inter1), .O(G695));

  xor2  gate2101(.a(G675), .b(G607), .O(gate215inter0));
  nand2 gate2102(.a(gate215inter0), .b(s_222), .O(gate215inter1));
  and2  gate2103(.a(G675), .b(G607), .O(gate215inter2));
  inv1  gate2104(.a(s_222), .O(gate215inter3));
  inv1  gate2105(.a(s_223), .O(gate215inter4));
  nand2 gate2106(.a(gate215inter4), .b(gate215inter3), .O(gate215inter5));
  nor2  gate2107(.a(gate215inter5), .b(gate215inter2), .O(gate215inter6));
  inv1  gate2108(.a(G607), .O(gate215inter7));
  inv1  gate2109(.a(G675), .O(gate215inter8));
  nand2 gate2110(.a(gate215inter8), .b(gate215inter7), .O(gate215inter9));
  nand2 gate2111(.a(s_223), .b(gate215inter3), .O(gate215inter10));
  nor2  gate2112(.a(gate215inter10), .b(gate215inter9), .O(gate215inter11));
  nor2  gate2113(.a(gate215inter11), .b(gate215inter6), .O(gate215inter12));
  nand2 gate2114(.a(gate215inter12), .b(gate215inter1), .O(G696));
nand2 gate216( .a(G617), .b(G675), .O(G697) );
nand2 gate217( .a(G622), .b(G678), .O(G698) );

  xor2  gate2591(.a(G678), .b(G627), .O(gate218inter0));
  nand2 gate2592(.a(gate218inter0), .b(s_292), .O(gate218inter1));
  and2  gate2593(.a(G678), .b(G627), .O(gate218inter2));
  inv1  gate2594(.a(s_292), .O(gate218inter3));
  inv1  gate2595(.a(s_293), .O(gate218inter4));
  nand2 gate2596(.a(gate218inter4), .b(gate218inter3), .O(gate218inter5));
  nor2  gate2597(.a(gate218inter5), .b(gate218inter2), .O(gate218inter6));
  inv1  gate2598(.a(G627), .O(gate218inter7));
  inv1  gate2599(.a(G678), .O(gate218inter8));
  nand2 gate2600(.a(gate218inter8), .b(gate218inter7), .O(gate218inter9));
  nand2 gate2601(.a(s_293), .b(gate218inter3), .O(gate218inter10));
  nor2  gate2602(.a(gate218inter10), .b(gate218inter9), .O(gate218inter11));
  nor2  gate2603(.a(gate218inter11), .b(gate218inter6), .O(gate218inter12));
  nand2 gate2604(.a(gate218inter12), .b(gate218inter1), .O(G699));
nand2 gate219( .a(G632), .b(G681), .O(G700) );

  xor2  gate2717(.a(G681), .b(G637), .O(gate220inter0));
  nand2 gate2718(.a(gate220inter0), .b(s_310), .O(gate220inter1));
  and2  gate2719(.a(G681), .b(G637), .O(gate220inter2));
  inv1  gate2720(.a(s_310), .O(gate220inter3));
  inv1  gate2721(.a(s_311), .O(gate220inter4));
  nand2 gate2722(.a(gate220inter4), .b(gate220inter3), .O(gate220inter5));
  nor2  gate2723(.a(gate220inter5), .b(gate220inter2), .O(gate220inter6));
  inv1  gate2724(.a(G637), .O(gate220inter7));
  inv1  gate2725(.a(G681), .O(gate220inter8));
  nand2 gate2726(.a(gate220inter8), .b(gate220inter7), .O(gate220inter9));
  nand2 gate2727(.a(s_311), .b(gate220inter3), .O(gate220inter10));
  nor2  gate2728(.a(gate220inter10), .b(gate220inter9), .O(gate220inter11));
  nor2  gate2729(.a(gate220inter11), .b(gate220inter6), .O(gate220inter12));
  nand2 gate2730(.a(gate220inter12), .b(gate220inter1), .O(G701));

  xor2  gate1709(.a(G684), .b(G622), .O(gate221inter0));
  nand2 gate1710(.a(gate221inter0), .b(s_166), .O(gate221inter1));
  and2  gate1711(.a(G684), .b(G622), .O(gate221inter2));
  inv1  gate1712(.a(s_166), .O(gate221inter3));
  inv1  gate1713(.a(s_167), .O(gate221inter4));
  nand2 gate1714(.a(gate221inter4), .b(gate221inter3), .O(gate221inter5));
  nor2  gate1715(.a(gate221inter5), .b(gate221inter2), .O(gate221inter6));
  inv1  gate1716(.a(G622), .O(gate221inter7));
  inv1  gate1717(.a(G684), .O(gate221inter8));
  nand2 gate1718(.a(gate221inter8), .b(gate221inter7), .O(gate221inter9));
  nand2 gate1719(.a(s_167), .b(gate221inter3), .O(gate221inter10));
  nor2  gate1720(.a(gate221inter10), .b(gate221inter9), .O(gate221inter11));
  nor2  gate1721(.a(gate221inter11), .b(gate221inter6), .O(gate221inter12));
  nand2 gate1722(.a(gate221inter12), .b(gate221inter1), .O(G702));

  xor2  gate771(.a(G684), .b(G632), .O(gate222inter0));
  nand2 gate772(.a(gate222inter0), .b(s_32), .O(gate222inter1));
  and2  gate773(.a(G684), .b(G632), .O(gate222inter2));
  inv1  gate774(.a(s_32), .O(gate222inter3));
  inv1  gate775(.a(s_33), .O(gate222inter4));
  nand2 gate776(.a(gate222inter4), .b(gate222inter3), .O(gate222inter5));
  nor2  gate777(.a(gate222inter5), .b(gate222inter2), .O(gate222inter6));
  inv1  gate778(.a(G632), .O(gate222inter7));
  inv1  gate779(.a(G684), .O(gate222inter8));
  nand2 gate780(.a(gate222inter8), .b(gate222inter7), .O(gate222inter9));
  nand2 gate781(.a(s_33), .b(gate222inter3), .O(gate222inter10));
  nor2  gate782(.a(gate222inter10), .b(gate222inter9), .O(gate222inter11));
  nor2  gate783(.a(gate222inter11), .b(gate222inter6), .O(gate222inter12));
  nand2 gate784(.a(gate222inter12), .b(gate222inter1), .O(G703));
nand2 gate223( .a(G627), .b(G687), .O(G704) );

  xor2  gate2801(.a(G687), .b(G637), .O(gate224inter0));
  nand2 gate2802(.a(gate224inter0), .b(s_322), .O(gate224inter1));
  and2  gate2803(.a(G687), .b(G637), .O(gate224inter2));
  inv1  gate2804(.a(s_322), .O(gate224inter3));
  inv1  gate2805(.a(s_323), .O(gate224inter4));
  nand2 gate2806(.a(gate224inter4), .b(gate224inter3), .O(gate224inter5));
  nor2  gate2807(.a(gate224inter5), .b(gate224inter2), .O(gate224inter6));
  inv1  gate2808(.a(G637), .O(gate224inter7));
  inv1  gate2809(.a(G687), .O(gate224inter8));
  nand2 gate2810(.a(gate224inter8), .b(gate224inter7), .O(gate224inter9));
  nand2 gate2811(.a(s_323), .b(gate224inter3), .O(gate224inter10));
  nor2  gate2812(.a(gate224inter10), .b(gate224inter9), .O(gate224inter11));
  nor2  gate2813(.a(gate224inter11), .b(gate224inter6), .O(gate224inter12));
  nand2 gate2814(.a(gate224inter12), .b(gate224inter1), .O(G705));
nand2 gate225( .a(G690), .b(G691), .O(G706) );
nand2 gate226( .a(G692), .b(G693), .O(G709) );
nand2 gate227( .a(G694), .b(G695), .O(G712) );

  xor2  gate1681(.a(G697), .b(G696), .O(gate228inter0));
  nand2 gate1682(.a(gate228inter0), .b(s_162), .O(gate228inter1));
  and2  gate1683(.a(G697), .b(G696), .O(gate228inter2));
  inv1  gate1684(.a(s_162), .O(gate228inter3));
  inv1  gate1685(.a(s_163), .O(gate228inter4));
  nand2 gate1686(.a(gate228inter4), .b(gate228inter3), .O(gate228inter5));
  nor2  gate1687(.a(gate228inter5), .b(gate228inter2), .O(gate228inter6));
  inv1  gate1688(.a(G696), .O(gate228inter7));
  inv1  gate1689(.a(G697), .O(gate228inter8));
  nand2 gate1690(.a(gate228inter8), .b(gate228inter7), .O(gate228inter9));
  nand2 gate1691(.a(s_163), .b(gate228inter3), .O(gate228inter10));
  nor2  gate1692(.a(gate228inter10), .b(gate228inter9), .O(gate228inter11));
  nor2  gate1693(.a(gate228inter11), .b(gate228inter6), .O(gate228inter12));
  nand2 gate1694(.a(gate228inter12), .b(gate228inter1), .O(G715));

  xor2  gate2339(.a(G699), .b(G698), .O(gate229inter0));
  nand2 gate2340(.a(gate229inter0), .b(s_256), .O(gate229inter1));
  and2  gate2341(.a(G699), .b(G698), .O(gate229inter2));
  inv1  gate2342(.a(s_256), .O(gate229inter3));
  inv1  gate2343(.a(s_257), .O(gate229inter4));
  nand2 gate2344(.a(gate229inter4), .b(gate229inter3), .O(gate229inter5));
  nor2  gate2345(.a(gate229inter5), .b(gate229inter2), .O(gate229inter6));
  inv1  gate2346(.a(G698), .O(gate229inter7));
  inv1  gate2347(.a(G699), .O(gate229inter8));
  nand2 gate2348(.a(gate229inter8), .b(gate229inter7), .O(gate229inter9));
  nand2 gate2349(.a(s_257), .b(gate229inter3), .O(gate229inter10));
  nor2  gate2350(.a(gate229inter10), .b(gate229inter9), .O(gate229inter11));
  nor2  gate2351(.a(gate229inter11), .b(gate229inter6), .O(gate229inter12));
  nand2 gate2352(.a(gate229inter12), .b(gate229inter1), .O(G718));
nand2 gate230( .a(G700), .b(G701), .O(G721) );

  xor2  gate1023(.a(G703), .b(G702), .O(gate231inter0));
  nand2 gate1024(.a(gate231inter0), .b(s_68), .O(gate231inter1));
  and2  gate1025(.a(G703), .b(G702), .O(gate231inter2));
  inv1  gate1026(.a(s_68), .O(gate231inter3));
  inv1  gate1027(.a(s_69), .O(gate231inter4));
  nand2 gate1028(.a(gate231inter4), .b(gate231inter3), .O(gate231inter5));
  nor2  gate1029(.a(gate231inter5), .b(gate231inter2), .O(gate231inter6));
  inv1  gate1030(.a(G702), .O(gate231inter7));
  inv1  gate1031(.a(G703), .O(gate231inter8));
  nand2 gate1032(.a(gate231inter8), .b(gate231inter7), .O(gate231inter9));
  nand2 gate1033(.a(s_69), .b(gate231inter3), .O(gate231inter10));
  nor2  gate1034(.a(gate231inter10), .b(gate231inter9), .O(gate231inter11));
  nor2  gate1035(.a(gate231inter11), .b(gate231inter6), .O(gate231inter12));
  nand2 gate1036(.a(gate231inter12), .b(gate231inter1), .O(G724));
nand2 gate232( .a(G704), .b(G705), .O(G727) );

  xor2  gate2941(.a(G718), .b(G242), .O(gate233inter0));
  nand2 gate2942(.a(gate233inter0), .b(s_342), .O(gate233inter1));
  and2  gate2943(.a(G718), .b(G242), .O(gate233inter2));
  inv1  gate2944(.a(s_342), .O(gate233inter3));
  inv1  gate2945(.a(s_343), .O(gate233inter4));
  nand2 gate2946(.a(gate233inter4), .b(gate233inter3), .O(gate233inter5));
  nor2  gate2947(.a(gate233inter5), .b(gate233inter2), .O(gate233inter6));
  inv1  gate2948(.a(G242), .O(gate233inter7));
  inv1  gate2949(.a(G718), .O(gate233inter8));
  nand2 gate2950(.a(gate233inter8), .b(gate233inter7), .O(gate233inter9));
  nand2 gate2951(.a(s_343), .b(gate233inter3), .O(gate233inter10));
  nor2  gate2952(.a(gate233inter10), .b(gate233inter9), .O(gate233inter11));
  nor2  gate2953(.a(gate233inter11), .b(gate233inter6), .O(gate233inter12));
  nand2 gate2954(.a(gate233inter12), .b(gate233inter1), .O(G730));
nand2 gate234( .a(G245), .b(G721), .O(G733) );

  xor2  gate1289(.a(G724), .b(G248), .O(gate235inter0));
  nand2 gate1290(.a(gate235inter0), .b(s_106), .O(gate235inter1));
  and2  gate1291(.a(G724), .b(G248), .O(gate235inter2));
  inv1  gate1292(.a(s_106), .O(gate235inter3));
  inv1  gate1293(.a(s_107), .O(gate235inter4));
  nand2 gate1294(.a(gate235inter4), .b(gate235inter3), .O(gate235inter5));
  nor2  gate1295(.a(gate235inter5), .b(gate235inter2), .O(gate235inter6));
  inv1  gate1296(.a(G248), .O(gate235inter7));
  inv1  gate1297(.a(G724), .O(gate235inter8));
  nand2 gate1298(.a(gate235inter8), .b(gate235inter7), .O(gate235inter9));
  nand2 gate1299(.a(s_107), .b(gate235inter3), .O(gate235inter10));
  nor2  gate1300(.a(gate235inter10), .b(gate235inter9), .O(gate235inter11));
  nor2  gate1301(.a(gate235inter11), .b(gate235inter6), .O(gate235inter12));
  nand2 gate1302(.a(gate235inter12), .b(gate235inter1), .O(G736));
nand2 gate236( .a(G251), .b(G727), .O(G739) );

  xor2  gate1961(.a(G706), .b(G254), .O(gate237inter0));
  nand2 gate1962(.a(gate237inter0), .b(s_202), .O(gate237inter1));
  and2  gate1963(.a(G706), .b(G254), .O(gate237inter2));
  inv1  gate1964(.a(s_202), .O(gate237inter3));
  inv1  gate1965(.a(s_203), .O(gate237inter4));
  nand2 gate1966(.a(gate237inter4), .b(gate237inter3), .O(gate237inter5));
  nor2  gate1967(.a(gate237inter5), .b(gate237inter2), .O(gate237inter6));
  inv1  gate1968(.a(G254), .O(gate237inter7));
  inv1  gate1969(.a(G706), .O(gate237inter8));
  nand2 gate1970(.a(gate237inter8), .b(gate237inter7), .O(gate237inter9));
  nand2 gate1971(.a(s_203), .b(gate237inter3), .O(gate237inter10));
  nor2  gate1972(.a(gate237inter10), .b(gate237inter9), .O(gate237inter11));
  nor2  gate1973(.a(gate237inter11), .b(gate237inter6), .O(gate237inter12));
  nand2 gate1974(.a(gate237inter12), .b(gate237inter1), .O(G742));

  xor2  gate2843(.a(G709), .b(G257), .O(gate238inter0));
  nand2 gate2844(.a(gate238inter0), .b(s_328), .O(gate238inter1));
  and2  gate2845(.a(G709), .b(G257), .O(gate238inter2));
  inv1  gate2846(.a(s_328), .O(gate238inter3));
  inv1  gate2847(.a(s_329), .O(gate238inter4));
  nand2 gate2848(.a(gate238inter4), .b(gate238inter3), .O(gate238inter5));
  nor2  gate2849(.a(gate238inter5), .b(gate238inter2), .O(gate238inter6));
  inv1  gate2850(.a(G257), .O(gate238inter7));
  inv1  gate2851(.a(G709), .O(gate238inter8));
  nand2 gate2852(.a(gate238inter8), .b(gate238inter7), .O(gate238inter9));
  nand2 gate2853(.a(s_329), .b(gate238inter3), .O(gate238inter10));
  nor2  gate2854(.a(gate238inter10), .b(gate238inter9), .O(gate238inter11));
  nor2  gate2855(.a(gate238inter11), .b(gate238inter6), .O(gate238inter12));
  nand2 gate2856(.a(gate238inter12), .b(gate238inter1), .O(G745));
nand2 gate239( .a(G260), .b(G712), .O(G748) );
nand2 gate240( .a(G263), .b(G715), .O(G751) );

  xor2  gate2773(.a(G730), .b(G242), .O(gate241inter0));
  nand2 gate2774(.a(gate241inter0), .b(s_318), .O(gate241inter1));
  and2  gate2775(.a(G730), .b(G242), .O(gate241inter2));
  inv1  gate2776(.a(s_318), .O(gate241inter3));
  inv1  gate2777(.a(s_319), .O(gate241inter4));
  nand2 gate2778(.a(gate241inter4), .b(gate241inter3), .O(gate241inter5));
  nor2  gate2779(.a(gate241inter5), .b(gate241inter2), .O(gate241inter6));
  inv1  gate2780(.a(G242), .O(gate241inter7));
  inv1  gate2781(.a(G730), .O(gate241inter8));
  nand2 gate2782(.a(gate241inter8), .b(gate241inter7), .O(gate241inter9));
  nand2 gate2783(.a(s_319), .b(gate241inter3), .O(gate241inter10));
  nor2  gate2784(.a(gate241inter10), .b(gate241inter9), .O(gate241inter11));
  nor2  gate2785(.a(gate241inter11), .b(gate241inter6), .O(gate241inter12));
  nand2 gate2786(.a(gate241inter12), .b(gate241inter1), .O(G754));
nand2 gate242( .a(G718), .b(G730), .O(G755) );

  xor2  gate2927(.a(G733), .b(G245), .O(gate243inter0));
  nand2 gate2928(.a(gate243inter0), .b(s_340), .O(gate243inter1));
  and2  gate2929(.a(G733), .b(G245), .O(gate243inter2));
  inv1  gate2930(.a(s_340), .O(gate243inter3));
  inv1  gate2931(.a(s_341), .O(gate243inter4));
  nand2 gate2932(.a(gate243inter4), .b(gate243inter3), .O(gate243inter5));
  nor2  gate2933(.a(gate243inter5), .b(gate243inter2), .O(gate243inter6));
  inv1  gate2934(.a(G245), .O(gate243inter7));
  inv1  gate2935(.a(G733), .O(gate243inter8));
  nand2 gate2936(.a(gate243inter8), .b(gate243inter7), .O(gate243inter9));
  nand2 gate2937(.a(s_341), .b(gate243inter3), .O(gate243inter10));
  nor2  gate2938(.a(gate243inter10), .b(gate243inter9), .O(gate243inter11));
  nor2  gate2939(.a(gate243inter11), .b(gate243inter6), .O(gate243inter12));
  nand2 gate2940(.a(gate243inter12), .b(gate243inter1), .O(G756));
nand2 gate244( .a(G721), .b(G733), .O(G757) );
nand2 gate245( .a(G248), .b(G736), .O(G758) );
nand2 gate246( .a(G724), .b(G736), .O(G759) );

  xor2  gate2787(.a(G739), .b(G251), .O(gate247inter0));
  nand2 gate2788(.a(gate247inter0), .b(s_320), .O(gate247inter1));
  and2  gate2789(.a(G739), .b(G251), .O(gate247inter2));
  inv1  gate2790(.a(s_320), .O(gate247inter3));
  inv1  gate2791(.a(s_321), .O(gate247inter4));
  nand2 gate2792(.a(gate247inter4), .b(gate247inter3), .O(gate247inter5));
  nor2  gate2793(.a(gate247inter5), .b(gate247inter2), .O(gate247inter6));
  inv1  gate2794(.a(G251), .O(gate247inter7));
  inv1  gate2795(.a(G739), .O(gate247inter8));
  nand2 gate2796(.a(gate247inter8), .b(gate247inter7), .O(gate247inter9));
  nand2 gate2797(.a(s_321), .b(gate247inter3), .O(gate247inter10));
  nor2  gate2798(.a(gate247inter10), .b(gate247inter9), .O(gate247inter11));
  nor2  gate2799(.a(gate247inter11), .b(gate247inter6), .O(gate247inter12));
  nand2 gate2800(.a(gate247inter12), .b(gate247inter1), .O(G760));
nand2 gate248( .a(G727), .b(G739), .O(G761) );

  xor2  gate2983(.a(G742), .b(G254), .O(gate249inter0));
  nand2 gate2984(.a(gate249inter0), .b(s_348), .O(gate249inter1));
  and2  gate2985(.a(G742), .b(G254), .O(gate249inter2));
  inv1  gate2986(.a(s_348), .O(gate249inter3));
  inv1  gate2987(.a(s_349), .O(gate249inter4));
  nand2 gate2988(.a(gate249inter4), .b(gate249inter3), .O(gate249inter5));
  nor2  gate2989(.a(gate249inter5), .b(gate249inter2), .O(gate249inter6));
  inv1  gate2990(.a(G254), .O(gate249inter7));
  inv1  gate2991(.a(G742), .O(gate249inter8));
  nand2 gate2992(.a(gate249inter8), .b(gate249inter7), .O(gate249inter9));
  nand2 gate2993(.a(s_349), .b(gate249inter3), .O(gate249inter10));
  nor2  gate2994(.a(gate249inter10), .b(gate249inter9), .O(gate249inter11));
  nor2  gate2995(.a(gate249inter11), .b(gate249inter6), .O(gate249inter12));
  nand2 gate2996(.a(gate249inter12), .b(gate249inter1), .O(G762));
nand2 gate250( .a(G706), .b(G742), .O(G763) );
nand2 gate251( .a(G257), .b(G745), .O(G764) );
nand2 gate252( .a(G709), .b(G745), .O(G765) );

  xor2  gate1765(.a(G748), .b(G260), .O(gate253inter0));
  nand2 gate1766(.a(gate253inter0), .b(s_174), .O(gate253inter1));
  and2  gate1767(.a(G748), .b(G260), .O(gate253inter2));
  inv1  gate1768(.a(s_174), .O(gate253inter3));
  inv1  gate1769(.a(s_175), .O(gate253inter4));
  nand2 gate1770(.a(gate253inter4), .b(gate253inter3), .O(gate253inter5));
  nor2  gate1771(.a(gate253inter5), .b(gate253inter2), .O(gate253inter6));
  inv1  gate1772(.a(G260), .O(gate253inter7));
  inv1  gate1773(.a(G748), .O(gate253inter8));
  nand2 gate1774(.a(gate253inter8), .b(gate253inter7), .O(gate253inter9));
  nand2 gate1775(.a(s_175), .b(gate253inter3), .O(gate253inter10));
  nor2  gate1776(.a(gate253inter10), .b(gate253inter9), .O(gate253inter11));
  nor2  gate1777(.a(gate253inter11), .b(gate253inter6), .O(gate253inter12));
  nand2 gate1778(.a(gate253inter12), .b(gate253inter1), .O(G766));

  xor2  gate2507(.a(G748), .b(G712), .O(gate254inter0));
  nand2 gate2508(.a(gate254inter0), .b(s_280), .O(gate254inter1));
  and2  gate2509(.a(G748), .b(G712), .O(gate254inter2));
  inv1  gate2510(.a(s_280), .O(gate254inter3));
  inv1  gate2511(.a(s_281), .O(gate254inter4));
  nand2 gate2512(.a(gate254inter4), .b(gate254inter3), .O(gate254inter5));
  nor2  gate2513(.a(gate254inter5), .b(gate254inter2), .O(gate254inter6));
  inv1  gate2514(.a(G712), .O(gate254inter7));
  inv1  gate2515(.a(G748), .O(gate254inter8));
  nand2 gate2516(.a(gate254inter8), .b(gate254inter7), .O(gate254inter9));
  nand2 gate2517(.a(s_281), .b(gate254inter3), .O(gate254inter10));
  nor2  gate2518(.a(gate254inter10), .b(gate254inter9), .O(gate254inter11));
  nor2  gate2519(.a(gate254inter11), .b(gate254inter6), .O(gate254inter12));
  nand2 gate2520(.a(gate254inter12), .b(gate254inter1), .O(G767));
nand2 gate255( .a(G263), .b(G751), .O(G768) );

  xor2  gate1807(.a(G751), .b(G715), .O(gate256inter0));
  nand2 gate1808(.a(gate256inter0), .b(s_180), .O(gate256inter1));
  and2  gate1809(.a(G751), .b(G715), .O(gate256inter2));
  inv1  gate1810(.a(s_180), .O(gate256inter3));
  inv1  gate1811(.a(s_181), .O(gate256inter4));
  nand2 gate1812(.a(gate256inter4), .b(gate256inter3), .O(gate256inter5));
  nor2  gate1813(.a(gate256inter5), .b(gate256inter2), .O(gate256inter6));
  inv1  gate1814(.a(G715), .O(gate256inter7));
  inv1  gate1815(.a(G751), .O(gate256inter8));
  nand2 gate1816(.a(gate256inter8), .b(gate256inter7), .O(gate256inter9));
  nand2 gate1817(.a(s_181), .b(gate256inter3), .O(gate256inter10));
  nor2  gate1818(.a(gate256inter10), .b(gate256inter9), .O(gate256inter11));
  nor2  gate1819(.a(gate256inter11), .b(gate256inter6), .O(gate256inter12));
  nand2 gate1820(.a(gate256inter12), .b(gate256inter1), .O(G769));
nand2 gate257( .a(G754), .b(G755), .O(G770) );

  xor2  gate2017(.a(G757), .b(G756), .O(gate258inter0));
  nand2 gate2018(.a(gate258inter0), .b(s_210), .O(gate258inter1));
  and2  gate2019(.a(G757), .b(G756), .O(gate258inter2));
  inv1  gate2020(.a(s_210), .O(gate258inter3));
  inv1  gate2021(.a(s_211), .O(gate258inter4));
  nand2 gate2022(.a(gate258inter4), .b(gate258inter3), .O(gate258inter5));
  nor2  gate2023(.a(gate258inter5), .b(gate258inter2), .O(gate258inter6));
  inv1  gate2024(.a(G756), .O(gate258inter7));
  inv1  gate2025(.a(G757), .O(gate258inter8));
  nand2 gate2026(.a(gate258inter8), .b(gate258inter7), .O(gate258inter9));
  nand2 gate2027(.a(s_211), .b(gate258inter3), .O(gate258inter10));
  nor2  gate2028(.a(gate258inter10), .b(gate258inter9), .O(gate258inter11));
  nor2  gate2029(.a(gate258inter11), .b(gate258inter6), .O(gate258inter12));
  nand2 gate2030(.a(gate258inter12), .b(gate258inter1), .O(G773));
nand2 gate259( .a(G758), .b(G759), .O(G776) );
nand2 gate260( .a(G760), .b(G761), .O(G779) );
nand2 gate261( .a(G762), .b(G763), .O(G782) );
nand2 gate262( .a(G764), .b(G765), .O(G785) );
nand2 gate263( .a(G766), .b(G767), .O(G788) );

  xor2  gate2955(.a(G769), .b(G768), .O(gate264inter0));
  nand2 gate2956(.a(gate264inter0), .b(s_344), .O(gate264inter1));
  and2  gate2957(.a(G769), .b(G768), .O(gate264inter2));
  inv1  gate2958(.a(s_344), .O(gate264inter3));
  inv1  gate2959(.a(s_345), .O(gate264inter4));
  nand2 gate2960(.a(gate264inter4), .b(gate264inter3), .O(gate264inter5));
  nor2  gate2961(.a(gate264inter5), .b(gate264inter2), .O(gate264inter6));
  inv1  gate2962(.a(G768), .O(gate264inter7));
  inv1  gate2963(.a(G769), .O(gate264inter8));
  nand2 gate2964(.a(gate264inter8), .b(gate264inter7), .O(gate264inter9));
  nand2 gate2965(.a(s_345), .b(gate264inter3), .O(gate264inter10));
  nor2  gate2966(.a(gate264inter10), .b(gate264inter9), .O(gate264inter11));
  nor2  gate2967(.a(gate264inter11), .b(gate264inter6), .O(gate264inter12));
  nand2 gate2968(.a(gate264inter12), .b(gate264inter1), .O(G791));
nand2 gate265( .a(G642), .b(G770), .O(G794) );

  xor2  gate855(.a(G773), .b(G645), .O(gate266inter0));
  nand2 gate856(.a(gate266inter0), .b(s_44), .O(gate266inter1));
  and2  gate857(.a(G773), .b(G645), .O(gate266inter2));
  inv1  gate858(.a(s_44), .O(gate266inter3));
  inv1  gate859(.a(s_45), .O(gate266inter4));
  nand2 gate860(.a(gate266inter4), .b(gate266inter3), .O(gate266inter5));
  nor2  gate861(.a(gate266inter5), .b(gate266inter2), .O(gate266inter6));
  inv1  gate862(.a(G645), .O(gate266inter7));
  inv1  gate863(.a(G773), .O(gate266inter8));
  nand2 gate864(.a(gate266inter8), .b(gate266inter7), .O(gate266inter9));
  nand2 gate865(.a(s_45), .b(gate266inter3), .O(gate266inter10));
  nor2  gate866(.a(gate266inter10), .b(gate266inter9), .O(gate266inter11));
  nor2  gate867(.a(gate266inter11), .b(gate266inter6), .O(gate266inter12));
  nand2 gate868(.a(gate266inter12), .b(gate266inter1), .O(G797));

  xor2  gate2885(.a(G776), .b(G648), .O(gate267inter0));
  nand2 gate2886(.a(gate267inter0), .b(s_334), .O(gate267inter1));
  and2  gate2887(.a(G776), .b(G648), .O(gate267inter2));
  inv1  gate2888(.a(s_334), .O(gate267inter3));
  inv1  gate2889(.a(s_335), .O(gate267inter4));
  nand2 gate2890(.a(gate267inter4), .b(gate267inter3), .O(gate267inter5));
  nor2  gate2891(.a(gate267inter5), .b(gate267inter2), .O(gate267inter6));
  inv1  gate2892(.a(G648), .O(gate267inter7));
  inv1  gate2893(.a(G776), .O(gate267inter8));
  nand2 gate2894(.a(gate267inter8), .b(gate267inter7), .O(gate267inter9));
  nand2 gate2895(.a(s_335), .b(gate267inter3), .O(gate267inter10));
  nor2  gate2896(.a(gate267inter10), .b(gate267inter9), .O(gate267inter11));
  nor2  gate2897(.a(gate267inter11), .b(gate267inter6), .O(gate267inter12));
  nand2 gate2898(.a(gate267inter12), .b(gate267inter1), .O(G800));
nand2 gate268( .a(G651), .b(G779), .O(G803) );
nand2 gate269( .a(G654), .b(G782), .O(G806) );
nand2 gate270( .a(G657), .b(G785), .O(G809) );

  xor2  gate785(.a(G788), .b(G660), .O(gate271inter0));
  nand2 gate786(.a(gate271inter0), .b(s_34), .O(gate271inter1));
  and2  gate787(.a(G788), .b(G660), .O(gate271inter2));
  inv1  gate788(.a(s_34), .O(gate271inter3));
  inv1  gate789(.a(s_35), .O(gate271inter4));
  nand2 gate790(.a(gate271inter4), .b(gate271inter3), .O(gate271inter5));
  nor2  gate791(.a(gate271inter5), .b(gate271inter2), .O(gate271inter6));
  inv1  gate792(.a(G660), .O(gate271inter7));
  inv1  gate793(.a(G788), .O(gate271inter8));
  nand2 gate794(.a(gate271inter8), .b(gate271inter7), .O(gate271inter9));
  nand2 gate795(.a(s_35), .b(gate271inter3), .O(gate271inter10));
  nor2  gate796(.a(gate271inter10), .b(gate271inter9), .O(gate271inter11));
  nor2  gate797(.a(gate271inter11), .b(gate271inter6), .O(gate271inter12));
  nand2 gate798(.a(gate271inter12), .b(gate271inter1), .O(G812));
nand2 gate272( .a(G663), .b(G791), .O(G815) );
nand2 gate273( .a(G642), .b(G794), .O(G818) );
nand2 gate274( .a(G770), .b(G794), .O(G819) );

  xor2  gate1177(.a(G797), .b(G645), .O(gate275inter0));
  nand2 gate1178(.a(gate275inter0), .b(s_90), .O(gate275inter1));
  and2  gate1179(.a(G797), .b(G645), .O(gate275inter2));
  inv1  gate1180(.a(s_90), .O(gate275inter3));
  inv1  gate1181(.a(s_91), .O(gate275inter4));
  nand2 gate1182(.a(gate275inter4), .b(gate275inter3), .O(gate275inter5));
  nor2  gate1183(.a(gate275inter5), .b(gate275inter2), .O(gate275inter6));
  inv1  gate1184(.a(G645), .O(gate275inter7));
  inv1  gate1185(.a(G797), .O(gate275inter8));
  nand2 gate1186(.a(gate275inter8), .b(gate275inter7), .O(gate275inter9));
  nand2 gate1187(.a(s_91), .b(gate275inter3), .O(gate275inter10));
  nor2  gate1188(.a(gate275inter10), .b(gate275inter9), .O(gate275inter11));
  nor2  gate1189(.a(gate275inter11), .b(gate275inter6), .O(gate275inter12));
  nand2 gate1190(.a(gate275inter12), .b(gate275inter1), .O(G820));
nand2 gate276( .a(G773), .b(G797), .O(G821) );
nand2 gate277( .a(G648), .b(G800), .O(G822) );
nand2 gate278( .a(G776), .b(G800), .O(G823) );
nand2 gate279( .a(G651), .b(G803), .O(G824) );

  xor2  gate1737(.a(G803), .b(G779), .O(gate280inter0));
  nand2 gate1738(.a(gate280inter0), .b(s_170), .O(gate280inter1));
  and2  gate1739(.a(G803), .b(G779), .O(gate280inter2));
  inv1  gate1740(.a(s_170), .O(gate280inter3));
  inv1  gate1741(.a(s_171), .O(gate280inter4));
  nand2 gate1742(.a(gate280inter4), .b(gate280inter3), .O(gate280inter5));
  nor2  gate1743(.a(gate280inter5), .b(gate280inter2), .O(gate280inter6));
  inv1  gate1744(.a(G779), .O(gate280inter7));
  inv1  gate1745(.a(G803), .O(gate280inter8));
  nand2 gate1746(.a(gate280inter8), .b(gate280inter7), .O(gate280inter9));
  nand2 gate1747(.a(s_171), .b(gate280inter3), .O(gate280inter10));
  nor2  gate1748(.a(gate280inter10), .b(gate280inter9), .O(gate280inter11));
  nor2  gate1749(.a(gate280inter11), .b(gate280inter6), .O(gate280inter12));
  nand2 gate1750(.a(gate280inter12), .b(gate280inter1), .O(G825));
nand2 gate281( .a(G654), .b(G806), .O(G826) );
nand2 gate282( .a(G782), .b(G806), .O(G827) );

  xor2  gate1429(.a(G809), .b(G657), .O(gate283inter0));
  nand2 gate1430(.a(gate283inter0), .b(s_126), .O(gate283inter1));
  and2  gate1431(.a(G809), .b(G657), .O(gate283inter2));
  inv1  gate1432(.a(s_126), .O(gate283inter3));
  inv1  gate1433(.a(s_127), .O(gate283inter4));
  nand2 gate1434(.a(gate283inter4), .b(gate283inter3), .O(gate283inter5));
  nor2  gate1435(.a(gate283inter5), .b(gate283inter2), .O(gate283inter6));
  inv1  gate1436(.a(G657), .O(gate283inter7));
  inv1  gate1437(.a(G809), .O(gate283inter8));
  nand2 gate1438(.a(gate283inter8), .b(gate283inter7), .O(gate283inter9));
  nand2 gate1439(.a(s_127), .b(gate283inter3), .O(gate283inter10));
  nor2  gate1440(.a(gate283inter10), .b(gate283inter9), .O(gate283inter11));
  nor2  gate1441(.a(gate283inter11), .b(gate283inter6), .O(gate283inter12));
  nand2 gate1442(.a(gate283inter12), .b(gate283inter1), .O(G828));

  xor2  gate687(.a(G809), .b(G785), .O(gate284inter0));
  nand2 gate688(.a(gate284inter0), .b(s_20), .O(gate284inter1));
  and2  gate689(.a(G809), .b(G785), .O(gate284inter2));
  inv1  gate690(.a(s_20), .O(gate284inter3));
  inv1  gate691(.a(s_21), .O(gate284inter4));
  nand2 gate692(.a(gate284inter4), .b(gate284inter3), .O(gate284inter5));
  nor2  gate693(.a(gate284inter5), .b(gate284inter2), .O(gate284inter6));
  inv1  gate694(.a(G785), .O(gate284inter7));
  inv1  gate695(.a(G809), .O(gate284inter8));
  nand2 gate696(.a(gate284inter8), .b(gate284inter7), .O(gate284inter9));
  nand2 gate697(.a(s_21), .b(gate284inter3), .O(gate284inter10));
  nor2  gate698(.a(gate284inter10), .b(gate284inter9), .O(gate284inter11));
  nor2  gate699(.a(gate284inter11), .b(gate284inter6), .O(gate284inter12));
  nand2 gate700(.a(gate284inter12), .b(gate284inter1), .O(G829));
nand2 gate285( .a(G660), .b(G812), .O(G830) );

  xor2  gate645(.a(G812), .b(G788), .O(gate286inter0));
  nand2 gate646(.a(gate286inter0), .b(s_14), .O(gate286inter1));
  and2  gate647(.a(G812), .b(G788), .O(gate286inter2));
  inv1  gate648(.a(s_14), .O(gate286inter3));
  inv1  gate649(.a(s_15), .O(gate286inter4));
  nand2 gate650(.a(gate286inter4), .b(gate286inter3), .O(gate286inter5));
  nor2  gate651(.a(gate286inter5), .b(gate286inter2), .O(gate286inter6));
  inv1  gate652(.a(G788), .O(gate286inter7));
  inv1  gate653(.a(G812), .O(gate286inter8));
  nand2 gate654(.a(gate286inter8), .b(gate286inter7), .O(gate286inter9));
  nand2 gate655(.a(s_15), .b(gate286inter3), .O(gate286inter10));
  nor2  gate656(.a(gate286inter10), .b(gate286inter9), .O(gate286inter11));
  nor2  gate657(.a(gate286inter11), .b(gate286inter6), .O(gate286inter12));
  nand2 gate658(.a(gate286inter12), .b(gate286inter1), .O(G831));
nand2 gate287( .a(G663), .b(G815), .O(G832) );

  xor2  gate1499(.a(G815), .b(G791), .O(gate288inter0));
  nand2 gate1500(.a(gate288inter0), .b(s_136), .O(gate288inter1));
  and2  gate1501(.a(G815), .b(G791), .O(gate288inter2));
  inv1  gate1502(.a(s_136), .O(gate288inter3));
  inv1  gate1503(.a(s_137), .O(gate288inter4));
  nand2 gate1504(.a(gate288inter4), .b(gate288inter3), .O(gate288inter5));
  nor2  gate1505(.a(gate288inter5), .b(gate288inter2), .O(gate288inter6));
  inv1  gate1506(.a(G791), .O(gate288inter7));
  inv1  gate1507(.a(G815), .O(gate288inter8));
  nand2 gate1508(.a(gate288inter8), .b(gate288inter7), .O(gate288inter9));
  nand2 gate1509(.a(s_137), .b(gate288inter3), .O(gate288inter10));
  nor2  gate1510(.a(gate288inter10), .b(gate288inter9), .O(gate288inter11));
  nor2  gate1511(.a(gate288inter11), .b(gate288inter6), .O(gate288inter12));
  nand2 gate1512(.a(gate288inter12), .b(gate288inter1), .O(G833));
nand2 gate289( .a(G818), .b(G819), .O(G834) );

  xor2  gate2213(.a(G821), .b(G820), .O(gate290inter0));
  nand2 gate2214(.a(gate290inter0), .b(s_238), .O(gate290inter1));
  and2  gate2215(.a(G821), .b(G820), .O(gate290inter2));
  inv1  gate2216(.a(s_238), .O(gate290inter3));
  inv1  gate2217(.a(s_239), .O(gate290inter4));
  nand2 gate2218(.a(gate290inter4), .b(gate290inter3), .O(gate290inter5));
  nor2  gate2219(.a(gate290inter5), .b(gate290inter2), .O(gate290inter6));
  inv1  gate2220(.a(G820), .O(gate290inter7));
  inv1  gate2221(.a(G821), .O(gate290inter8));
  nand2 gate2222(.a(gate290inter8), .b(gate290inter7), .O(gate290inter9));
  nand2 gate2223(.a(s_239), .b(gate290inter3), .O(gate290inter10));
  nor2  gate2224(.a(gate290inter10), .b(gate290inter9), .O(gate290inter11));
  nor2  gate2225(.a(gate290inter11), .b(gate290inter6), .O(gate290inter12));
  nand2 gate2226(.a(gate290inter12), .b(gate290inter1), .O(G847));
nand2 gate291( .a(G822), .b(G823), .O(G860) );
nand2 gate292( .a(G824), .b(G825), .O(G873) );
nand2 gate293( .a(G828), .b(G829), .O(G886) );

  xor2  gate729(.a(G833), .b(G832), .O(gate294inter0));
  nand2 gate730(.a(gate294inter0), .b(s_26), .O(gate294inter1));
  and2  gate731(.a(G833), .b(G832), .O(gate294inter2));
  inv1  gate732(.a(s_26), .O(gate294inter3));
  inv1  gate733(.a(s_27), .O(gate294inter4));
  nand2 gate734(.a(gate294inter4), .b(gate294inter3), .O(gate294inter5));
  nor2  gate735(.a(gate294inter5), .b(gate294inter2), .O(gate294inter6));
  inv1  gate736(.a(G832), .O(gate294inter7));
  inv1  gate737(.a(G833), .O(gate294inter8));
  nand2 gate738(.a(gate294inter8), .b(gate294inter7), .O(gate294inter9));
  nand2 gate739(.a(s_27), .b(gate294inter3), .O(gate294inter10));
  nor2  gate740(.a(gate294inter10), .b(gate294inter9), .O(gate294inter11));
  nor2  gate741(.a(gate294inter11), .b(gate294inter6), .O(gate294inter12));
  nand2 gate742(.a(gate294inter12), .b(gate294inter1), .O(G899));
nand2 gate295( .a(G830), .b(G831), .O(G912) );
nand2 gate296( .a(G826), .b(G827), .O(G925) );
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );
nand2 gate387( .a(G1), .b(G1036), .O(G1132) );
nand2 gate388( .a(G2), .b(G1039), .O(G1135) );
nand2 gate389( .a(G3), .b(G1042), .O(G1138) );
nand2 gate390( .a(G4), .b(G1045), .O(G1141) );

  xor2  gate1905(.a(G1048), .b(G5), .O(gate391inter0));
  nand2 gate1906(.a(gate391inter0), .b(s_194), .O(gate391inter1));
  and2  gate1907(.a(G1048), .b(G5), .O(gate391inter2));
  inv1  gate1908(.a(s_194), .O(gate391inter3));
  inv1  gate1909(.a(s_195), .O(gate391inter4));
  nand2 gate1910(.a(gate391inter4), .b(gate391inter3), .O(gate391inter5));
  nor2  gate1911(.a(gate391inter5), .b(gate391inter2), .O(gate391inter6));
  inv1  gate1912(.a(G5), .O(gate391inter7));
  inv1  gate1913(.a(G1048), .O(gate391inter8));
  nand2 gate1914(.a(gate391inter8), .b(gate391inter7), .O(gate391inter9));
  nand2 gate1915(.a(s_195), .b(gate391inter3), .O(gate391inter10));
  nor2  gate1916(.a(gate391inter10), .b(gate391inter9), .O(gate391inter11));
  nor2  gate1917(.a(gate391inter11), .b(gate391inter6), .O(gate391inter12));
  nand2 gate1918(.a(gate391inter12), .b(gate391inter1), .O(G1144));
nand2 gate392( .a(G6), .b(G1051), .O(G1147) );
nand2 gate393( .a(G7), .b(G1054), .O(G1150) );

  xor2  gate1387(.a(G1057), .b(G8), .O(gate394inter0));
  nand2 gate1388(.a(gate394inter0), .b(s_120), .O(gate394inter1));
  and2  gate1389(.a(G1057), .b(G8), .O(gate394inter2));
  inv1  gate1390(.a(s_120), .O(gate394inter3));
  inv1  gate1391(.a(s_121), .O(gate394inter4));
  nand2 gate1392(.a(gate394inter4), .b(gate394inter3), .O(gate394inter5));
  nor2  gate1393(.a(gate394inter5), .b(gate394inter2), .O(gate394inter6));
  inv1  gate1394(.a(G8), .O(gate394inter7));
  inv1  gate1395(.a(G1057), .O(gate394inter8));
  nand2 gate1396(.a(gate394inter8), .b(gate394inter7), .O(gate394inter9));
  nand2 gate1397(.a(s_121), .b(gate394inter3), .O(gate394inter10));
  nor2  gate1398(.a(gate394inter10), .b(gate394inter9), .O(gate394inter11));
  nor2  gate1399(.a(gate394inter11), .b(gate394inter6), .O(gate394inter12));
  nand2 gate1400(.a(gate394inter12), .b(gate394inter1), .O(G1153));

  xor2  gate3137(.a(G1060), .b(G9), .O(gate395inter0));
  nand2 gate3138(.a(gate395inter0), .b(s_370), .O(gate395inter1));
  and2  gate3139(.a(G1060), .b(G9), .O(gate395inter2));
  inv1  gate3140(.a(s_370), .O(gate395inter3));
  inv1  gate3141(.a(s_371), .O(gate395inter4));
  nand2 gate3142(.a(gate395inter4), .b(gate395inter3), .O(gate395inter5));
  nor2  gate3143(.a(gate395inter5), .b(gate395inter2), .O(gate395inter6));
  inv1  gate3144(.a(G9), .O(gate395inter7));
  inv1  gate3145(.a(G1060), .O(gate395inter8));
  nand2 gate3146(.a(gate395inter8), .b(gate395inter7), .O(gate395inter9));
  nand2 gate3147(.a(s_371), .b(gate395inter3), .O(gate395inter10));
  nor2  gate3148(.a(gate395inter10), .b(gate395inter9), .O(gate395inter11));
  nor2  gate3149(.a(gate395inter11), .b(gate395inter6), .O(gate395inter12));
  nand2 gate3150(.a(gate395inter12), .b(gate395inter1), .O(G1156));
nand2 gate396( .a(G10), .b(G1063), .O(G1159) );

  xor2  gate3053(.a(G1066), .b(G11), .O(gate397inter0));
  nand2 gate3054(.a(gate397inter0), .b(s_358), .O(gate397inter1));
  and2  gate3055(.a(G1066), .b(G11), .O(gate397inter2));
  inv1  gate3056(.a(s_358), .O(gate397inter3));
  inv1  gate3057(.a(s_359), .O(gate397inter4));
  nand2 gate3058(.a(gate397inter4), .b(gate397inter3), .O(gate397inter5));
  nor2  gate3059(.a(gate397inter5), .b(gate397inter2), .O(gate397inter6));
  inv1  gate3060(.a(G11), .O(gate397inter7));
  inv1  gate3061(.a(G1066), .O(gate397inter8));
  nand2 gate3062(.a(gate397inter8), .b(gate397inter7), .O(gate397inter9));
  nand2 gate3063(.a(s_359), .b(gate397inter3), .O(gate397inter10));
  nor2  gate3064(.a(gate397inter10), .b(gate397inter9), .O(gate397inter11));
  nor2  gate3065(.a(gate397inter11), .b(gate397inter6), .O(gate397inter12));
  nand2 gate3066(.a(gate397inter12), .b(gate397inter1), .O(G1162));
nand2 gate398( .a(G12), .b(G1069), .O(G1165) );
nand2 gate399( .a(G13), .b(G1072), .O(G1168) );

  xor2  gate813(.a(G1075), .b(G14), .O(gate400inter0));
  nand2 gate814(.a(gate400inter0), .b(s_38), .O(gate400inter1));
  and2  gate815(.a(G1075), .b(G14), .O(gate400inter2));
  inv1  gate816(.a(s_38), .O(gate400inter3));
  inv1  gate817(.a(s_39), .O(gate400inter4));
  nand2 gate818(.a(gate400inter4), .b(gate400inter3), .O(gate400inter5));
  nor2  gate819(.a(gate400inter5), .b(gate400inter2), .O(gate400inter6));
  inv1  gate820(.a(G14), .O(gate400inter7));
  inv1  gate821(.a(G1075), .O(gate400inter8));
  nand2 gate822(.a(gate400inter8), .b(gate400inter7), .O(gate400inter9));
  nand2 gate823(.a(s_39), .b(gate400inter3), .O(gate400inter10));
  nor2  gate824(.a(gate400inter10), .b(gate400inter9), .O(gate400inter11));
  nor2  gate825(.a(gate400inter11), .b(gate400inter6), .O(gate400inter12));
  nand2 gate826(.a(gate400inter12), .b(gate400inter1), .O(G1171));
nand2 gate401( .a(G15), .b(G1078), .O(G1174) );

  xor2  gate1835(.a(G1081), .b(G16), .O(gate402inter0));
  nand2 gate1836(.a(gate402inter0), .b(s_184), .O(gate402inter1));
  and2  gate1837(.a(G1081), .b(G16), .O(gate402inter2));
  inv1  gate1838(.a(s_184), .O(gate402inter3));
  inv1  gate1839(.a(s_185), .O(gate402inter4));
  nand2 gate1840(.a(gate402inter4), .b(gate402inter3), .O(gate402inter5));
  nor2  gate1841(.a(gate402inter5), .b(gate402inter2), .O(gate402inter6));
  inv1  gate1842(.a(G16), .O(gate402inter7));
  inv1  gate1843(.a(G1081), .O(gate402inter8));
  nand2 gate1844(.a(gate402inter8), .b(gate402inter7), .O(gate402inter9));
  nand2 gate1845(.a(s_185), .b(gate402inter3), .O(gate402inter10));
  nor2  gate1846(.a(gate402inter10), .b(gate402inter9), .O(gate402inter11));
  nor2  gate1847(.a(gate402inter11), .b(gate402inter6), .O(gate402inter12));
  nand2 gate1848(.a(gate402inter12), .b(gate402inter1), .O(G1177));

  xor2  gate2297(.a(G1084), .b(G17), .O(gate403inter0));
  nand2 gate2298(.a(gate403inter0), .b(s_250), .O(gate403inter1));
  and2  gate2299(.a(G1084), .b(G17), .O(gate403inter2));
  inv1  gate2300(.a(s_250), .O(gate403inter3));
  inv1  gate2301(.a(s_251), .O(gate403inter4));
  nand2 gate2302(.a(gate403inter4), .b(gate403inter3), .O(gate403inter5));
  nor2  gate2303(.a(gate403inter5), .b(gate403inter2), .O(gate403inter6));
  inv1  gate2304(.a(G17), .O(gate403inter7));
  inv1  gate2305(.a(G1084), .O(gate403inter8));
  nand2 gate2306(.a(gate403inter8), .b(gate403inter7), .O(gate403inter9));
  nand2 gate2307(.a(s_251), .b(gate403inter3), .O(gate403inter10));
  nor2  gate2308(.a(gate403inter10), .b(gate403inter9), .O(gate403inter11));
  nor2  gate2309(.a(gate403inter11), .b(gate403inter6), .O(gate403inter12));
  nand2 gate2310(.a(gate403inter12), .b(gate403inter1), .O(G1180));

  xor2  gate2493(.a(G1087), .b(G18), .O(gate404inter0));
  nand2 gate2494(.a(gate404inter0), .b(s_278), .O(gate404inter1));
  and2  gate2495(.a(G1087), .b(G18), .O(gate404inter2));
  inv1  gate2496(.a(s_278), .O(gate404inter3));
  inv1  gate2497(.a(s_279), .O(gate404inter4));
  nand2 gate2498(.a(gate404inter4), .b(gate404inter3), .O(gate404inter5));
  nor2  gate2499(.a(gate404inter5), .b(gate404inter2), .O(gate404inter6));
  inv1  gate2500(.a(G18), .O(gate404inter7));
  inv1  gate2501(.a(G1087), .O(gate404inter8));
  nand2 gate2502(.a(gate404inter8), .b(gate404inter7), .O(gate404inter9));
  nand2 gate2503(.a(s_279), .b(gate404inter3), .O(gate404inter10));
  nor2  gate2504(.a(gate404inter10), .b(gate404inter9), .O(gate404inter11));
  nor2  gate2505(.a(gate404inter11), .b(gate404inter6), .O(gate404inter12));
  nand2 gate2506(.a(gate404inter12), .b(gate404inter1), .O(G1183));

  xor2  gate603(.a(G1090), .b(G19), .O(gate405inter0));
  nand2 gate604(.a(gate405inter0), .b(s_8), .O(gate405inter1));
  and2  gate605(.a(G1090), .b(G19), .O(gate405inter2));
  inv1  gate606(.a(s_8), .O(gate405inter3));
  inv1  gate607(.a(s_9), .O(gate405inter4));
  nand2 gate608(.a(gate405inter4), .b(gate405inter3), .O(gate405inter5));
  nor2  gate609(.a(gate405inter5), .b(gate405inter2), .O(gate405inter6));
  inv1  gate610(.a(G19), .O(gate405inter7));
  inv1  gate611(.a(G1090), .O(gate405inter8));
  nand2 gate612(.a(gate405inter8), .b(gate405inter7), .O(gate405inter9));
  nand2 gate613(.a(s_9), .b(gate405inter3), .O(gate405inter10));
  nor2  gate614(.a(gate405inter10), .b(gate405inter9), .O(gate405inter11));
  nor2  gate615(.a(gate405inter11), .b(gate405inter6), .O(gate405inter12));
  nand2 gate616(.a(gate405inter12), .b(gate405inter1), .O(G1186));

  xor2  gate715(.a(G1093), .b(G20), .O(gate406inter0));
  nand2 gate716(.a(gate406inter0), .b(s_24), .O(gate406inter1));
  and2  gate717(.a(G1093), .b(G20), .O(gate406inter2));
  inv1  gate718(.a(s_24), .O(gate406inter3));
  inv1  gate719(.a(s_25), .O(gate406inter4));
  nand2 gate720(.a(gate406inter4), .b(gate406inter3), .O(gate406inter5));
  nor2  gate721(.a(gate406inter5), .b(gate406inter2), .O(gate406inter6));
  inv1  gate722(.a(G20), .O(gate406inter7));
  inv1  gate723(.a(G1093), .O(gate406inter8));
  nand2 gate724(.a(gate406inter8), .b(gate406inter7), .O(gate406inter9));
  nand2 gate725(.a(s_25), .b(gate406inter3), .O(gate406inter10));
  nor2  gate726(.a(gate406inter10), .b(gate406inter9), .O(gate406inter11));
  nor2  gate727(.a(gate406inter11), .b(gate406inter6), .O(gate406inter12));
  nand2 gate728(.a(gate406inter12), .b(gate406inter1), .O(G1189));

  xor2  gate2283(.a(G1096), .b(G21), .O(gate407inter0));
  nand2 gate2284(.a(gate407inter0), .b(s_248), .O(gate407inter1));
  and2  gate2285(.a(G1096), .b(G21), .O(gate407inter2));
  inv1  gate2286(.a(s_248), .O(gate407inter3));
  inv1  gate2287(.a(s_249), .O(gate407inter4));
  nand2 gate2288(.a(gate407inter4), .b(gate407inter3), .O(gate407inter5));
  nor2  gate2289(.a(gate407inter5), .b(gate407inter2), .O(gate407inter6));
  inv1  gate2290(.a(G21), .O(gate407inter7));
  inv1  gate2291(.a(G1096), .O(gate407inter8));
  nand2 gate2292(.a(gate407inter8), .b(gate407inter7), .O(gate407inter9));
  nand2 gate2293(.a(s_249), .b(gate407inter3), .O(gate407inter10));
  nor2  gate2294(.a(gate407inter10), .b(gate407inter9), .O(gate407inter11));
  nor2  gate2295(.a(gate407inter11), .b(gate407inter6), .O(gate407inter12));
  nand2 gate2296(.a(gate407inter12), .b(gate407inter1), .O(G1192));

  xor2  gate1219(.a(G1099), .b(G22), .O(gate408inter0));
  nand2 gate1220(.a(gate408inter0), .b(s_96), .O(gate408inter1));
  and2  gate1221(.a(G1099), .b(G22), .O(gate408inter2));
  inv1  gate1222(.a(s_96), .O(gate408inter3));
  inv1  gate1223(.a(s_97), .O(gate408inter4));
  nand2 gate1224(.a(gate408inter4), .b(gate408inter3), .O(gate408inter5));
  nor2  gate1225(.a(gate408inter5), .b(gate408inter2), .O(gate408inter6));
  inv1  gate1226(.a(G22), .O(gate408inter7));
  inv1  gate1227(.a(G1099), .O(gate408inter8));
  nand2 gate1228(.a(gate408inter8), .b(gate408inter7), .O(gate408inter9));
  nand2 gate1229(.a(s_97), .b(gate408inter3), .O(gate408inter10));
  nor2  gate1230(.a(gate408inter10), .b(gate408inter9), .O(gate408inter11));
  nor2  gate1231(.a(gate408inter11), .b(gate408inter6), .O(gate408inter12));
  nand2 gate1232(.a(gate408inter12), .b(gate408inter1), .O(G1195));
nand2 gate409( .a(G23), .b(G1102), .O(G1198) );
nand2 gate410( .a(G24), .b(G1105), .O(G1201) );
nand2 gate411( .a(G25), .b(G1108), .O(G1204) );
nand2 gate412( .a(G26), .b(G1111), .O(G1207) );
nand2 gate413( .a(G27), .b(G1114), .O(G1210) );

  xor2  gate1345(.a(G1117), .b(G28), .O(gate414inter0));
  nand2 gate1346(.a(gate414inter0), .b(s_114), .O(gate414inter1));
  and2  gate1347(.a(G1117), .b(G28), .O(gate414inter2));
  inv1  gate1348(.a(s_114), .O(gate414inter3));
  inv1  gate1349(.a(s_115), .O(gate414inter4));
  nand2 gate1350(.a(gate414inter4), .b(gate414inter3), .O(gate414inter5));
  nor2  gate1351(.a(gate414inter5), .b(gate414inter2), .O(gate414inter6));
  inv1  gate1352(.a(G28), .O(gate414inter7));
  inv1  gate1353(.a(G1117), .O(gate414inter8));
  nand2 gate1354(.a(gate414inter8), .b(gate414inter7), .O(gate414inter9));
  nand2 gate1355(.a(s_115), .b(gate414inter3), .O(gate414inter10));
  nor2  gate1356(.a(gate414inter10), .b(gate414inter9), .O(gate414inter11));
  nor2  gate1357(.a(gate414inter11), .b(gate414inter6), .O(gate414inter12));
  nand2 gate1358(.a(gate414inter12), .b(gate414inter1), .O(G1213));

  xor2  gate1485(.a(G1120), .b(G29), .O(gate415inter0));
  nand2 gate1486(.a(gate415inter0), .b(s_134), .O(gate415inter1));
  and2  gate1487(.a(G1120), .b(G29), .O(gate415inter2));
  inv1  gate1488(.a(s_134), .O(gate415inter3));
  inv1  gate1489(.a(s_135), .O(gate415inter4));
  nand2 gate1490(.a(gate415inter4), .b(gate415inter3), .O(gate415inter5));
  nor2  gate1491(.a(gate415inter5), .b(gate415inter2), .O(gate415inter6));
  inv1  gate1492(.a(G29), .O(gate415inter7));
  inv1  gate1493(.a(G1120), .O(gate415inter8));
  nand2 gate1494(.a(gate415inter8), .b(gate415inter7), .O(gate415inter9));
  nand2 gate1495(.a(s_135), .b(gate415inter3), .O(gate415inter10));
  nor2  gate1496(.a(gate415inter10), .b(gate415inter9), .O(gate415inter11));
  nor2  gate1497(.a(gate415inter11), .b(gate415inter6), .O(gate415inter12));
  nand2 gate1498(.a(gate415inter12), .b(gate415inter1), .O(G1216));

  xor2  gate1527(.a(G1123), .b(G30), .O(gate416inter0));
  nand2 gate1528(.a(gate416inter0), .b(s_140), .O(gate416inter1));
  and2  gate1529(.a(G1123), .b(G30), .O(gate416inter2));
  inv1  gate1530(.a(s_140), .O(gate416inter3));
  inv1  gate1531(.a(s_141), .O(gate416inter4));
  nand2 gate1532(.a(gate416inter4), .b(gate416inter3), .O(gate416inter5));
  nor2  gate1533(.a(gate416inter5), .b(gate416inter2), .O(gate416inter6));
  inv1  gate1534(.a(G30), .O(gate416inter7));
  inv1  gate1535(.a(G1123), .O(gate416inter8));
  nand2 gate1536(.a(gate416inter8), .b(gate416inter7), .O(gate416inter9));
  nand2 gate1537(.a(s_141), .b(gate416inter3), .O(gate416inter10));
  nor2  gate1538(.a(gate416inter10), .b(gate416inter9), .O(gate416inter11));
  nor2  gate1539(.a(gate416inter11), .b(gate416inter6), .O(gate416inter12));
  nand2 gate1540(.a(gate416inter12), .b(gate416inter1), .O(G1219));
nand2 gate417( .a(G31), .b(G1126), .O(G1222) );

  xor2  gate911(.a(G1129), .b(G32), .O(gate418inter0));
  nand2 gate912(.a(gate418inter0), .b(s_52), .O(gate418inter1));
  and2  gate913(.a(G1129), .b(G32), .O(gate418inter2));
  inv1  gate914(.a(s_52), .O(gate418inter3));
  inv1  gate915(.a(s_53), .O(gate418inter4));
  nand2 gate916(.a(gate418inter4), .b(gate418inter3), .O(gate418inter5));
  nor2  gate917(.a(gate418inter5), .b(gate418inter2), .O(gate418inter6));
  inv1  gate918(.a(G32), .O(gate418inter7));
  inv1  gate919(.a(G1129), .O(gate418inter8));
  nand2 gate920(.a(gate418inter8), .b(gate418inter7), .O(gate418inter9));
  nand2 gate921(.a(s_53), .b(gate418inter3), .O(gate418inter10));
  nor2  gate922(.a(gate418inter10), .b(gate418inter9), .O(gate418inter11));
  nor2  gate923(.a(gate418inter11), .b(gate418inter6), .O(gate418inter12));
  nand2 gate924(.a(gate418inter12), .b(gate418inter1), .O(G1225));

  xor2  gate2969(.a(G1132), .b(G1), .O(gate419inter0));
  nand2 gate2970(.a(gate419inter0), .b(s_346), .O(gate419inter1));
  and2  gate2971(.a(G1132), .b(G1), .O(gate419inter2));
  inv1  gate2972(.a(s_346), .O(gate419inter3));
  inv1  gate2973(.a(s_347), .O(gate419inter4));
  nand2 gate2974(.a(gate419inter4), .b(gate419inter3), .O(gate419inter5));
  nor2  gate2975(.a(gate419inter5), .b(gate419inter2), .O(gate419inter6));
  inv1  gate2976(.a(G1), .O(gate419inter7));
  inv1  gate2977(.a(G1132), .O(gate419inter8));
  nand2 gate2978(.a(gate419inter8), .b(gate419inter7), .O(gate419inter9));
  nand2 gate2979(.a(s_347), .b(gate419inter3), .O(gate419inter10));
  nor2  gate2980(.a(gate419inter10), .b(gate419inter9), .O(gate419inter11));
  nor2  gate2981(.a(gate419inter11), .b(gate419inter6), .O(gate419inter12));
  nand2 gate2982(.a(gate419inter12), .b(gate419inter1), .O(G1228));
nand2 gate420( .a(G1036), .b(G1132), .O(G1229) );

  xor2  gate953(.a(G1135), .b(G2), .O(gate421inter0));
  nand2 gate954(.a(gate421inter0), .b(s_58), .O(gate421inter1));
  and2  gate955(.a(G1135), .b(G2), .O(gate421inter2));
  inv1  gate956(.a(s_58), .O(gate421inter3));
  inv1  gate957(.a(s_59), .O(gate421inter4));
  nand2 gate958(.a(gate421inter4), .b(gate421inter3), .O(gate421inter5));
  nor2  gate959(.a(gate421inter5), .b(gate421inter2), .O(gate421inter6));
  inv1  gate960(.a(G2), .O(gate421inter7));
  inv1  gate961(.a(G1135), .O(gate421inter8));
  nand2 gate962(.a(gate421inter8), .b(gate421inter7), .O(gate421inter9));
  nand2 gate963(.a(s_59), .b(gate421inter3), .O(gate421inter10));
  nor2  gate964(.a(gate421inter10), .b(gate421inter9), .O(gate421inter11));
  nor2  gate965(.a(gate421inter11), .b(gate421inter6), .O(gate421inter12));
  nand2 gate966(.a(gate421inter12), .b(gate421inter1), .O(G1230));
nand2 gate422( .a(G1039), .b(G1135), .O(G1231) );
nand2 gate423( .a(G3), .b(G1138), .O(G1232) );
nand2 gate424( .a(G1042), .b(G1138), .O(G1233) );
nand2 gate425( .a(G4), .b(G1141), .O(G1234) );
nand2 gate426( .a(G1045), .b(G1141), .O(G1235) );
nand2 gate427( .a(G5), .b(G1144), .O(G1236) );

  xor2  gate1457(.a(G1144), .b(G1048), .O(gate428inter0));
  nand2 gate1458(.a(gate428inter0), .b(s_130), .O(gate428inter1));
  and2  gate1459(.a(G1144), .b(G1048), .O(gate428inter2));
  inv1  gate1460(.a(s_130), .O(gate428inter3));
  inv1  gate1461(.a(s_131), .O(gate428inter4));
  nand2 gate1462(.a(gate428inter4), .b(gate428inter3), .O(gate428inter5));
  nor2  gate1463(.a(gate428inter5), .b(gate428inter2), .O(gate428inter6));
  inv1  gate1464(.a(G1048), .O(gate428inter7));
  inv1  gate1465(.a(G1144), .O(gate428inter8));
  nand2 gate1466(.a(gate428inter8), .b(gate428inter7), .O(gate428inter9));
  nand2 gate1467(.a(s_131), .b(gate428inter3), .O(gate428inter10));
  nor2  gate1468(.a(gate428inter10), .b(gate428inter9), .O(gate428inter11));
  nor2  gate1469(.a(gate428inter11), .b(gate428inter6), .O(gate428inter12));
  nand2 gate1470(.a(gate428inter12), .b(gate428inter1), .O(G1237));

  xor2  gate1751(.a(G1147), .b(G6), .O(gate429inter0));
  nand2 gate1752(.a(gate429inter0), .b(s_172), .O(gate429inter1));
  and2  gate1753(.a(G1147), .b(G6), .O(gate429inter2));
  inv1  gate1754(.a(s_172), .O(gate429inter3));
  inv1  gate1755(.a(s_173), .O(gate429inter4));
  nand2 gate1756(.a(gate429inter4), .b(gate429inter3), .O(gate429inter5));
  nor2  gate1757(.a(gate429inter5), .b(gate429inter2), .O(gate429inter6));
  inv1  gate1758(.a(G6), .O(gate429inter7));
  inv1  gate1759(.a(G1147), .O(gate429inter8));
  nand2 gate1760(.a(gate429inter8), .b(gate429inter7), .O(gate429inter9));
  nand2 gate1761(.a(s_173), .b(gate429inter3), .O(gate429inter10));
  nor2  gate1762(.a(gate429inter10), .b(gate429inter9), .O(gate429inter11));
  nor2  gate1763(.a(gate429inter11), .b(gate429inter6), .O(gate429inter12));
  nand2 gate1764(.a(gate429inter12), .b(gate429inter1), .O(G1238));

  xor2  gate2325(.a(G1147), .b(G1051), .O(gate430inter0));
  nand2 gate2326(.a(gate430inter0), .b(s_254), .O(gate430inter1));
  and2  gate2327(.a(G1147), .b(G1051), .O(gate430inter2));
  inv1  gate2328(.a(s_254), .O(gate430inter3));
  inv1  gate2329(.a(s_255), .O(gate430inter4));
  nand2 gate2330(.a(gate430inter4), .b(gate430inter3), .O(gate430inter5));
  nor2  gate2331(.a(gate430inter5), .b(gate430inter2), .O(gate430inter6));
  inv1  gate2332(.a(G1051), .O(gate430inter7));
  inv1  gate2333(.a(G1147), .O(gate430inter8));
  nand2 gate2334(.a(gate430inter8), .b(gate430inter7), .O(gate430inter9));
  nand2 gate2335(.a(s_255), .b(gate430inter3), .O(gate430inter10));
  nor2  gate2336(.a(gate430inter10), .b(gate430inter9), .O(gate430inter11));
  nor2  gate2337(.a(gate430inter11), .b(gate430inter6), .O(gate430inter12));
  nand2 gate2338(.a(gate430inter12), .b(gate430inter1), .O(G1239));
nand2 gate431( .a(G7), .b(G1150), .O(G1240) );
nand2 gate432( .a(G1054), .b(G1150), .O(G1241) );

  xor2  gate925(.a(G1153), .b(G8), .O(gate433inter0));
  nand2 gate926(.a(gate433inter0), .b(s_54), .O(gate433inter1));
  and2  gate927(.a(G1153), .b(G8), .O(gate433inter2));
  inv1  gate928(.a(s_54), .O(gate433inter3));
  inv1  gate929(.a(s_55), .O(gate433inter4));
  nand2 gate930(.a(gate433inter4), .b(gate433inter3), .O(gate433inter5));
  nor2  gate931(.a(gate433inter5), .b(gate433inter2), .O(gate433inter6));
  inv1  gate932(.a(G8), .O(gate433inter7));
  inv1  gate933(.a(G1153), .O(gate433inter8));
  nand2 gate934(.a(gate433inter8), .b(gate433inter7), .O(gate433inter9));
  nand2 gate935(.a(s_55), .b(gate433inter3), .O(gate433inter10));
  nor2  gate936(.a(gate433inter10), .b(gate433inter9), .O(gate433inter11));
  nor2  gate937(.a(gate433inter11), .b(gate433inter6), .O(gate433inter12));
  nand2 gate938(.a(gate433inter12), .b(gate433inter1), .O(G1242));
nand2 gate434( .a(G1057), .b(G1153), .O(G1243) );

  xor2  gate589(.a(G1156), .b(G9), .O(gate435inter0));
  nand2 gate590(.a(gate435inter0), .b(s_6), .O(gate435inter1));
  and2  gate591(.a(G1156), .b(G9), .O(gate435inter2));
  inv1  gate592(.a(s_6), .O(gate435inter3));
  inv1  gate593(.a(s_7), .O(gate435inter4));
  nand2 gate594(.a(gate435inter4), .b(gate435inter3), .O(gate435inter5));
  nor2  gate595(.a(gate435inter5), .b(gate435inter2), .O(gate435inter6));
  inv1  gate596(.a(G9), .O(gate435inter7));
  inv1  gate597(.a(G1156), .O(gate435inter8));
  nand2 gate598(.a(gate435inter8), .b(gate435inter7), .O(gate435inter9));
  nand2 gate599(.a(s_7), .b(gate435inter3), .O(gate435inter10));
  nor2  gate600(.a(gate435inter10), .b(gate435inter9), .O(gate435inter11));
  nor2  gate601(.a(gate435inter11), .b(gate435inter6), .O(gate435inter12));
  nand2 gate602(.a(gate435inter12), .b(gate435inter1), .O(G1244));

  xor2  gate1891(.a(G1156), .b(G1060), .O(gate436inter0));
  nand2 gate1892(.a(gate436inter0), .b(s_192), .O(gate436inter1));
  and2  gate1893(.a(G1156), .b(G1060), .O(gate436inter2));
  inv1  gate1894(.a(s_192), .O(gate436inter3));
  inv1  gate1895(.a(s_193), .O(gate436inter4));
  nand2 gate1896(.a(gate436inter4), .b(gate436inter3), .O(gate436inter5));
  nor2  gate1897(.a(gate436inter5), .b(gate436inter2), .O(gate436inter6));
  inv1  gate1898(.a(G1060), .O(gate436inter7));
  inv1  gate1899(.a(G1156), .O(gate436inter8));
  nand2 gate1900(.a(gate436inter8), .b(gate436inter7), .O(gate436inter9));
  nand2 gate1901(.a(s_193), .b(gate436inter3), .O(gate436inter10));
  nor2  gate1902(.a(gate436inter10), .b(gate436inter9), .O(gate436inter11));
  nor2  gate1903(.a(gate436inter11), .b(gate436inter6), .O(gate436inter12));
  nand2 gate1904(.a(gate436inter12), .b(gate436inter1), .O(G1245));
nand2 gate437( .a(G10), .b(G1159), .O(G1246) );
nand2 gate438( .a(G1063), .b(G1159), .O(G1247) );

  xor2  gate2479(.a(G1162), .b(G11), .O(gate439inter0));
  nand2 gate2480(.a(gate439inter0), .b(s_276), .O(gate439inter1));
  and2  gate2481(.a(G1162), .b(G11), .O(gate439inter2));
  inv1  gate2482(.a(s_276), .O(gate439inter3));
  inv1  gate2483(.a(s_277), .O(gate439inter4));
  nand2 gate2484(.a(gate439inter4), .b(gate439inter3), .O(gate439inter5));
  nor2  gate2485(.a(gate439inter5), .b(gate439inter2), .O(gate439inter6));
  inv1  gate2486(.a(G11), .O(gate439inter7));
  inv1  gate2487(.a(G1162), .O(gate439inter8));
  nand2 gate2488(.a(gate439inter8), .b(gate439inter7), .O(gate439inter9));
  nand2 gate2489(.a(s_277), .b(gate439inter3), .O(gate439inter10));
  nor2  gate2490(.a(gate439inter10), .b(gate439inter9), .O(gate439inter11));
  nor2  gate2491(.a(gate439inter11), .b(gate439inter6), .O(gate439inter12));
  nand2 gate2492(.a(gate439inter12), .b(gate439inter1), .O(G1248));
nand2 gate440( .a(G1066), .b(G1162), .O(G1249) );

  xor2  gate1443(.a(G1165), .b(G12), .O(gate441inter0));
  nand2 gate1444(.a(gate441inter0), .b(s_128), .O(gate441inter1));
  and2  gate1445(.a(G1165), .b(G12), .O(gate441inter2));
  inv1  gate1446(.a(s_128), .O(gate441inter3));
  inv1  gate1447(.a(s_129), .O(gate441inter4));
  nand2 gate1448(.a(gate441inter4), .b(gate441inter3), .O(gate441inter5));
  nor2  gate1449(.a(gate441inter5), .b(gate441inter2), .O(gate441inter6));
  inv1  gate1450(.a(G12), .O(gate441inter7));
  inv1  gate1451(.a(G1165), .O(gate441inter8));
  nand2 gate1452(.a(gate441inter8), .b(gate441inter7), .O(gate441inter9));
  nand2 gate1453(.a(s_129), .b(gate441inter3), .O(gate441inter10));
  nor2  gate1454(.a(gate441inter10), .b(gate441inter9), .O(gate441inter11));
  nor2  gate1455(.a(gate441inter11), .b(gate441inter6), .O(gate441inter12));
  nand2 gate1456(.a(gate441inter12), .b(gate441inter1), .O(G1250));
nand2 gate442( .a(G1069), .b(G1165), .O(G1251) );
nand2 gate443( .a(G13), .b(G1168), .O(G1252) );
nand2 gate444( .a(G1072), .b(G1168), .O(G1253) );
nand2 gate445( .a(G14), .b(G1171), .O(G1254) );
nand2 gate446( .a(G1075), .b(G1171), .O(G1255) );

  xor2  gate3095(.a(G1174), .b(G15), .O(gate447inter0));
  nand2 gate3096(.a(gate447inter0), .b(s_364), .O(gate447inter1));
  and2  gate3097(.a(G1174), .b(G15), .O(gate447inter2));
  inv1  gate3098(.a(s_364), .O(gate447inter3));
  inv1  gate3099(.a(s_365), .O(gate447inter4));
  nand2 gate3100(.a(gate447inter4), .b(gate447inter3), .O(gate447inter5));
  nor2  gate3101(.a(gate447inter5), .b(gate447inter2), .O(gate447inter6));
  inv1  gate3102(.a(G15), .O(gate447inter7));
  inv1  gate3103(.a(G1174), .O(gate447inter8));
  nand2 gate3104(.a(gate447inter8), .b(gate447inter7), .O(gate447inter9));
  nand2 gate3105(.a(s_365), .b(gate447inter3), .O(gate447inter10));
  nor2  gate3106(.a(gate447inter10), .b(gate447inter9), .O(gate447inter11));
  nor2  gate3107(.a(gate447inter11), .b(gate447inter6), .O(gate447inter12));
  nand2 gate3108(.a(gate447inter12), .b(gate447inter1), .O(G1256));

  xor2  gate1037(.a(G1174), .b(G1078), .O(gate448inter0));
  nand2 gate1038(.a(gate448inter0), .b(s_70), .O(gate448inter1));
  and2  gate1039(.a(G1174), .b(G1078), .O(gate448inter2));
  inv1  gate1040(.a(s_70), .O(gate448inter3));
  inv1  gate1041(.a(s_71), .O(gate448inter4));
  nand2 gate1042(.a(gate448inter4), .b(gate448inter3), .O(gate448inter5));
  nor2  gate1043(.a(gate448inter5), .b(gate448inter2), .O(gate448inter6));
  inv1  gate1044(.a(G1078), .O(gate448inter7));
  inv1  gate1045(.a(G1174), .O(gate448inter8));
  nand2 gate1046(.a(gate448inter8), .b(gate448inter7), .O(gate448inter9));
  nand2 gate1047(.a(s_71), .b(gate448inter3), .O(gate448inter10));
  nor2  gate1048(.a(gate448inter10), .b(gate448inter9), .O(gate448inter11));
  nor2  gate1049(.a(gate448inter11), .b(gate448inter6), .O(gate448inter12));
  nand2 gate1050(.a(gate448inter12), .b(gate448inter1), .O(G1257));

  xor2  gate3109(.a(G1177), .b(G16), .O(gate449inter0));
  nand2 gate3110(.a(gate449inter0), .b(s_366), .O(gate449inter1));
  and2  gate3111(.a(G1177), .b(G16), .O(gate449inter2));
  inv1  gate3112(.a(s_366), .O(gate449inter3));
  inv1  gate3113(.a(s_367), .O(gate449inter4));
  nand2 gate3114(.a(gate449inter4), .b(gate449inter3), .O(gate449inter5));
  nor2  gate3115(.a(gate449inter5), .b(gate449inter2), .O(gate449inter6));
  inv1  gate3116(.a(G16), .O(gate449inter7));
  inv1  gate3117(.a(G1177), .O(gate449inter8));
  nand2 gate3118(.a(gate449inter8), .b(gate449inter7), .O(gate449inter9));
  nand2 gate3119(.a(s_367), .b(gate449inter3), .O(gate449inter10));
  nor2  gate3120(.a(gate449inter10), .b(gate449inter9), .O(gate449inter11));
  nor2  gate3121(.a(gate449inter11), .b(gate449inter6), .O(gate449inter12));
  nand2 gate3122(.a(gate449inter12), .b(gate449inter1), .O(G1258));
nand2 gate450( .a(G1081), .b(G1177), .O(G1259) );
nand2 gate451( .a(G17), .b(G1180), .O(G1260) );
nand2 gate452( .a(G1084), .b(G1180), .O(G1261) );

  xor2  gate2913(.a(G1183), .b(G18), .O(gate453inter0));
  nand2 gate2914(.a(gate453inter0), .b(s_338), .O(gate453inter1));
  and2  gate2915(.a(G1183), .b(G18), .O(gate453inter2));
  inv1  gate2916(.a(s_338), .O(gate453inter3));
  inv1  gate2917(.a(s_339), .O(gate453inter4));
  nand2 gate2918(.a(gate453inter4), .b(gate453inter3), .O(gate453inter5));
  nor2  gate2919(.a(gate453inter5), .b(gate453inter2), .O(gate453inter6));
  inv1  gate2920(.a(G18), .O(gate453inter7));
  inv1  gate2921(.a(G1183), .O(gate453inter8));
  nand2 gate2922(.a(gate453inter8), .b(gate453inter7), .O(gate453inter9));
  nand2 gate2923(.a(s_339), .b(gate453inter3), .O(gate453inter10));
  nor2  gate2924(.a(gate453inter10), .b(gate453inter9), .O(gate453inter11));
  nor2  gate2925(.a(gate453inter11), .b(gate453inter6), .O(gate453inter12));
  nand2 gate2926(.a(gate453inter12), .b(gate453inter1), .O(G1262));
nand2 gate454( .a(G1087), .b(G1183), .O(G1263) );
nand2 gate455( .a(G19), .b(G1186), .O(G1264) );

  xor2  gate1933(.a(G1186), .b(G1090), .O(gate456inter0));
  nand2 gate1934(.a(gate456inter0), .b(s_198), .O(gate456inter1));
  and2  gate1935(.a(G1186), .b(G1090), .O(gate456inter2));
  inv1  gate1936(.a(s_198), .O(gate456inter3));
  inv1  gate1937(.a(s_199), .O(gate456inter4));
  nand2 gate1938(.a(gate456inter4), .b(gate456inter3), .O(gate456inter5));
  nor2  gate1939(.a(gate456inter5), .b(gate456inter2), .O(gate456inter6));
  inv1  gate1940(.a(G1090), .O(gate456inter7));
  inv1  gate1941(.a(G1186), .O(gate456inter8));
  nand2 gate1942(.a(gate456inter8), .b(gate456inter7), .O(gate456inter9));
  nand2 gate1943(.a(s_199), .b(gate456inter3), .O(gate456inter10));
  nor2  gate1944(.a(gate456inter10), .b(gate456inter9), .O(gate456inter11));
  nor2  gate1945(.a(gate456inter11), .b(gate456inter6), .O(gate456inter12));
  nand2 gate1946(.a(gate456inter12), .b(gate456inter1), .O(G1265));

  xor2  gate1163(.a(G1189), .b(G20), .O(gate457inter0));
  nand2 gate1164(.a(gate457inter0), .b(s_88), .O(gate457inter1));
  and2  gate1165(.a(G1189), .b(G20), .O(gate457inter2));
  inv1  gate1166(.a(s_88), .O(gate457inter3));
  inv1  gate1167(.a(s_89), .O(gate457inter4));
  nand2 gate1168(.a(gate457inter4), .b(gate457inter3), .O(gate457inter5));
  nor2  gate1169(.a(gate457inter5), .b(gate457inter2), .O(gate457inter6));
  inv1  gate1170(.a(G20), .O(gate457inter7));
  inv1  gate1171(.a(G1189), .O(gate457inter8));
  nand2 gate1172(.a(gate457inter8), .b(gate457inter7), .O(gate457inter9));
  nand2 gate1173(.a(s_89), .b(gate457inter3), .O(gate457inter10));
  nor2  gate1174(.a(gate457inter10), .b(gate457inter9), .O(gate457inter11));
  nor2  gate1175(.a(gate457inter11), .b(gate457inter6), .O(gate457inter12));
  nand2 gate1176(.a(gate457inter12), .b(gate457inter1), .O(G1266));
nand2 gate458( .a(G1093), .b(G1189), .O(G1267) );

  xor2  gate1317(.a(G1192), .b(G21), .O(gate459inter0));
  nand2 gate1318(.a(gate459inter0), .b(s_110), .O(gate459inter1));
  and2  gate1319(.a(G1192), .b(G21), .O(gate459inter2));
  inv1  gate1320(.a(s_110), .O(gate459inter3));
  inv1  gate1321(.a(s_111), .O(gate459inter4));
  nand2 gate1322(.a(gate459inter4), .b(gate459inter3), .O(gate459inter5));
  nor2  gate1323(.a(gate459inter5), .b(gate459inter2), .O(gate459inter6));
  inv1  gate1324(.a(G21), .O(gate459inter7));
  inv1  gate1325(.a(G1192), .O(gate459inter8));
  nand2 gate1326(.a(gate459inter8), .b(gate459inter7), .O(gate459inter9));
  nand2 gate1327(.a(s_111), .b(gate459inter3), .O(gate459inter10));
  nor2  gate1328(.a(gate459inter10), .b(gate459inter9), .O(gate459inter11));
  nor2  gate1329(.a(gate459inter11), .b(gate459inter6), .O(gate459inter12));
  nand2 gate1330(.a(gate459inter12), .b(gate459inter1), .O(G1268));

  xor2  gate2059(.a(G1192), .b(G1096), .O(gate460inter0));
  nand2 gate2060(.a(gate460inter0), .b(s_216), .O(gate460inter1));
  and2  gate2061(.a(G1192), .b(G1096), .O(gate460inter2));
  inv1  gate2062(.a(s_216), .O(gate460inter3));
  inv1  gate2063(.a(s_217), .O(gate460inter4));
  nand2 gate2064(.a(gate460inter4), .b(gate460inter3), .O(gate460inter5));
  nor2  gate2065(.a(gate460inter5), .b(gate460inter2), .O(gate460inter6));
  inv1  gate2066(.a(G1096), .O(gate460inter7));
  inv1  gate2067(.a(G1192), .O(gate460inter8));
  nand2 gate2068(.a(gate460inter8), .b(gate460inter7), .O(gate460inter9));
  nand2 gate2069(.a(s_217), .b(gate460inter3), .O(gate460inter10));
  nor2  gate2070(.a(gate460inter10), .b(gate460inter9), .O(gate460inter11));
  nor2  gate2071(.a(gate460inter11), .b(gate460inter6), .O(gate460inter12));
  nand2 gate2072(.a(gate460inter12), .b(gate460inter1), .O(G1269));
nand2 gate461( .a(G22), .b(G1195), .O(G1270) );
nand2 gate462( .a(G1099), .b(G1195), .O(G1271) );
nand2 gate463( .a(G23), .b(G1198), .O(G1272) );
nand2 gate464( .a(G1102), .b(G1198), .O(G1273) );
nand2 gate465( .a(G24), .b(G1201), .O(G1274) );
nand2 gate466( .a(G1105), .b(G1201), .O(G1275) );

  xor2  gate2521(.a(G1204), .b(G25), .O(gate467inter0));
  nand2 gate2522(.a(gate467inter0), .b(s_282), .O(gate467inter1));
  and2  gate2523(.a(G1204), .b(G25), .O(gate467inter2));
  inv1  gate2524(.a(s_282), .O(gate467inter3));
  inv1  gate2525(.a(s_283), .O(gate467inter4));
  nand2 gate2526(.a(gate467inter4), .b(gate467inter3), .O(gate467inter5));
  nor2  gate2527(.a(gate467inter5), .b(gate467inter2), .O(gate467inter6));
  inv1  gate2528(.a(G25), .O(gate467inter7));
  inv1  gate2529(.a(G1204), .O(gate467inter8));
  nand2 gate2530(.a(gate467inter8), .b(gate467inter7), .O(gate467inter9));
  nand2 gate2531(.a(s_283), .b(gate467inter3), .O(gate467inter10));
  nor2  gate2532(.a(gate467inter10), .b(gate467inter9), .O(gate467inter11));
  nor2  gate2533(.a(gate467inter11), .b(gate467inter6), .O(gate467inter12));
  nand2 gate2534(.a(gate467inter12), .b(gate467inter1), .O(G1276));
nand2 gate468( .a(G1108), .b(G1204), .O(G1277) );

  xor2  gate2871(.a(G1207), .b(G26), .O(gate469inter0));
  nand2 gate2872(.a(gate469inter0), .b(s_332), .O(gate469inter1));
  and2  gate2873(.a(G1207), .b(G26), .O(gate469inter2));
  inv1  gate2874(.a(s_332), .O(gate469inter3));
  inv1  gate2875(.a(s_333), .O(gate469inter4));
  nand2 gate2876(.a(gate469inter4), .b(gate469inter3), .O(gate469inter5));
  nor2  gate2877(.a(gate469inter5), .b(gate469inter2), .O(gate469inter6));
  inv1  gate2878(.a(G26), .O(gate469inter7));
  inv1  gate2879(.a(G1207), .O(gate469inter8));
  nand2 gate2880(.a(gate469inter8), .b(gate469inter7), .O(gate469inter9));
  nand2 gate2881(.a(s_333), .b(gate469inter3), .O(gate469inter10));
  nor2  gate2882(.a(gate469inter10), .b(gate469inter9), .O(gate469inter11));
  nor2  gate2883(.a(gate469inter11), .b(gate469inter6), .O(gate469inter12));
  nand2 gate2884(.a(gate469inter12), .b(gate469inter1), .O(G1278));

  xor2  gate2185(.a(G1207), .b(G1111), .O(gate470inter0));
  nand2 gate2186(.a(gate470inter0), .b(s_234), .O(gate470inter1));
  and2  gate2187(.a(G1207), .b(G1111), .O(gate470inter2));
  inv1  gate2188(.a(s_234), .O(gate470inter3));
  inv1  gate2189(.a(s_235), .O(gate470inter4));
  nand2 gate2190(.a(gate470inter4), .b(gate470inter3), .O(gate470inter5));
  nor2  gate2191(.a(gate470inter5), .b(gate470inter2), .O(gate470inter6));
  inv1  gate2192(.a(G1111), .O(gate470inter7));
  inv1  gate2193(.a(G1207), .O(gate470inter8));
  nand2 gate2194(.a(gate470inter8), .b(gate470inter7), .O(gate470inter9));
  nand2 gate2195(.a(s_235), .b(gate470inter3), .O(gate470inter10));
  nor2  gate2196(.a(gate470inter10), .b(gate470inter9), .O(gate470inter11));
  nor2  gate2197(.a(gate470inter11), .b(gate470inter6), .O(gate470inter12));
  nand2 gate2198(.a(gate470inter12), .b(gate470inter1), .O(G1279));
nand2 gate471( .a(G27), .b(G1210), .O(G1280) );
nand2 gate472( .a(G1114), .b(G1210), .O(G1281) );

  xor2  gate2759(.a(G1213), .b(G28), .O(gate473inter0));
  nand2 gate2760(.a(gate473inter0), .b(s_316), .O(gate473inter1));
  and2  gate2761(.a(G1213), .b(G28), .O(gate473inter2));
  inv1  gate2762(.a(s_316), .O(gate473inter3));
  inv1  gate2763(.a(s_317), .O(gate473inter4));
  nand2 gate2764(.a(gate473inter4), .b(gate473inter3), .O(gate473inter5));
  nor2  gate2765(.a(gate473inter5), .b(gate473inter2), .O(gate473inter6));
  inv1  gate2766(.a(G28), .O(gate473inter7));
  inv1  gate2767(.a(G1213), .O(gate473inter8));
  nand2 gate2768(.a(gate473inter8), .b(gate473inter7), .O(gate473inter9));
  nand2 gate2769(.a(s_317), .b(gate473inter3), .O(gate473inter10));
  nor2  gate2770(.a(gate473inter10), .b(gate473inter9), .O(gate473inter11));
  nor2  gate2771(.a(gate473inter11), .b(gate473inter6), .O(gate473inter12));
  nand2 gate2772(.a(gate473inter12), .b(gate473inter1), .O(G1282));
nand2 gate474( .a(G1117), .b(G1213), .O(G1283) );
nand2 gate475( .a(G29), .b(G1216), .O(G1284) );
nand2 gate476( .a(G1120), .b(G1216), .O(G1285) );

  xor2  gate1695(.a(G1219), .b(G30), .O(gate477inter0));
  nand2 gate1696(.a(gate477inter0), .b(s_164), .O(gate477inter1));
  and2  gate1697(.a(G1219), .b(G30), .O(gate477inter2));
  inv1  gate1698(.a(s_164), .O(gate477inter3));
  inv1  gate1699(.a(s_165), .O(gate477inter4));
  nand2 gate1700(.a(gate477inter4), .b(gate477inter3), .O(gate477inter5));
  nor2  gate1701(.a(gate477inter5), .b(gate477inter2), .O(gate477inter6));
  inv1  gate1702(.a(G30), .O(gate477inter7));
  inv1  gate1703(.a(G1219), .O(gate477inter8));
  nand2 gate1704(.a(gate477inter8), .b(gate477inter7), .O(gate477inter9));
  nand2 gate1705(.a(s_165), .b(gate477inter3), .O(gate477inter10));
  nor2  gate1706(.a(gate477inter10), .b(gate477inter9), .O(gate477inter11));
  nor2  gate1707(.a(gate477inter11), .b(gate477inter6), .O(gate477inter12));
  nand2 gate1708(.a(gate477inter12), .b(gate477inter1), .O(G1286));
nand2 gate478( .a(G1123), .b(G1219), .O(G1287) );

  xor2  gate2227(.a(G1222), .b(G31), .O(gate479inter0));
  nand2 gate2228(.a(gate479inter0), .b(s_240), .O(gate479inter1));
  and2  gate2229(.a(G1222), .b(G31), .O(gate479inter2));
  inv1  gate2230(.a(s_240), .O(gate479inter3));
  inv1  gate2231(.a(s_241), .O(gate479inter4));
  nand2 gate2232(.a(gate479inter4), .b(gate479inter3), .O(gate479inter5));
  nor2  gate2233(.a(gate479inter5), .b(gate479inter2), .O(gate479inter6));
  inv1  gate2234(.a(G31), .O(gate479inter7));
  inv1  gate2235(.a(G1222), .O(gate479inter8));
  nand2 gate2236(.a(gate479inter8), .b(gate479inter7), .O(gate479inter9));
  nand2 gate2237(.a(s_241), .b(gate479inter3), .O(gate479inter10));
  nor2  gate2238(.a(gate479inter10), .b(gate479inter9), .O(gate479inter11));
  nor2  gate2239(.a(gate479inter11), .b(gate479inter6), .O(gate479inter12));
  nand2 gate2240(.a(gate479inter12), .b(gate479inter1), .O(G1288));

  xor2  gate2661(.a(G1222), .b(G1126), .O(gate480inter0));
  nand2 gate2662(.a(gate480inter0), .b(s_302), .O(gate480inter1));
  and2  gate2663(.a(G1222), .b(G1126), .O(gate480inter2));
  inv1  gate2664(.a(s_302), .O(gate480inter3));
  inv1  gate2665(.a(s_303), .O(gate480inter4));
  nand2 gate2666(.a(gate480inter4), .b(gate480inter3), .O(gate480inter5));
  nor2  gate2667(.a(gate480inter5), .b(gate480inter2), .O(gate480inter6));
  inv1  gate2668(.a(G1126), .O(gate480inter7));
  inv1  gate2669(.a(G1222), .O(gate480inter8));
  nand2 gate2670(.a(gate480inter8), .b(gate480inter7), .O(gate480inter9));
  nand2 gate2671(.a(s_303), .b(gate480inter3), .O(gate480inter10));
  nor2  gate2672(.a(gate480inter10), .b(gate480inter9), .O(gate480inter11));
  nor2  gate2673(.a(gate480inter11), .b(gate480inter6), .O(gate480inter12));
  nand2 gate2674(.a(gate480inter12), .b(gate480inter1), .O(G1289));
nand2 gate481( .a(G32), .b(G1225), .O(G1290) );

  xor2  gate869(.a(G1225), .b(G1129), .O(gate482inter0));
  nand2 gate870(.a(gate482inter0), .b(s_46), .O(gate482inter1));
  and2  gate871(.a(G1225), .b(G1129), .O(gate482inter2));
  inv1  gate872(.a(s_46), .O(gate482inter3));
  inv1  gate873(.a(s_47), .O(gate482inter4));
  nand2 gate874(.a(gate482inter4), .b(gate482inter3), .O(gate482inter5));
  nor2  gate875(.a(gate482inter5), .b(gate482inter2), .O(gate482inter6));
  inv1  gate876(.a(G1129), .O(gate482inter7));
  inv1  gate877(.a(G1225), .O(gate482inter8));
  nand2 gate878(.a(gate482inter8), .b(gate482inter7), .O(gate482inter9));
  nand2 gate879(.a(s_47), .b(gate482inter3), .O(gate482inter10));
  nor2  gate880(.a(gate482inter10), .b(gate482inter9), .O(gate482inter11));
  nor2  gate881(.a(gate482inter11), .b(gate482inter6), .O(gate482inter12));
  nand2 gate882(.a(gate482inter12), .b(gate482inter1), .O(G1291));

  xor2  gate2157(.a(G1229), .b(G1228), .O(gate483inter0));
  nand2 gate2158(.a(gate483inter0), .b(s_230), .O(gate483inter1));
  and2  gate2159(.a(G1229), .b(G1228), .O(gate483inter2));
  inv1  gate2160(.a(s_230), .O(gate483inter3));
  inv1  gate2161(.a(s_231), .O(gate483inter4));
  nand2 gate2162(.a(gate483inter4), .b(gate483inter3), .O(gate483inter5));
  nor2  gate2163(.a(gate483inter5), .b(gate483inter2), .O(gate483inter6));
  inv1  gate2164(.a(G1228), .O(gate483inter7));
  inv1  gate2165(.a(G1229), .O(gate483inter8));
  nand2 gate2166(.a(gate483inter8), .b(gate483inter7), .O(gate483inter9));
  nand2 gate2167(.a(s_231), .b(gate483inter3), .O(gate483inter10));
  nor2  gate2168(.a(gate483inter10), .b(gate483inter9), .O(gate483inter11));
  nor2  gate2169(.a(gate483inter11), .b(gate483inter6), .O(gate483inter12));
  nand2 gate2170(.a(gate483inter12), .b(gate483inter1), .O(G1292));
nand2 gate484( .a(G1230), .b(G1231), .O(G1293) );

  xor2  gate2619(.a(G1233), .b(G1232), .O(gate485inter0));
  nand2 gate2620(.a(gate485inter0), .b(s_296), .O(gate485inter1));
  and2  gate2621(.a(G1233), .b(G1232), .O(gate485inter2));
  inv1  gate2622(.a(s_296), .O(gate485inter3));
  inv1  gate2623(.a(s_297), .O(gate485inter4));
  nand2 gate2624(.a(gate485inter4), .b(gate485inter3), .O(gate485inter5));
  nor2  gate2625(.a(gate485inter5), .b(gate485inter2), .O(gate485inter6));
  inv1  gate2626(.a(G1232), .O(gate485inter7));
  inv1  gate2627(.a(G1233), .O(gate485inter8));
  nand2 gate2628(.a(gate485inter8), .b(gate485inter7), .O(gate485inter9));
  nand2 gate2629(.a(s_297), .b(gate485inter3), .O(gate485inter10));
  nor2  gate2630(.a(gate485inter10), .b(gate485inter9), .O(gate485inter11));
  nor2  gate2631(.a(gate485inter11), .b(gate485inter6), .O(gate485inter12));
  nand2 gate2632(.a(gate485inter12), .b(gate485inter1), .O(G1294));
nand2 gate486( .a(G1234), .b(G1235), .O(G1295) );

  xor2  gate1051(.a(G1237), .b(G1236), .O(gate487inter0));
  nand2 gate1052(.a(gate487inter0), .b(s_72), .O(gate487inter1));
  and2  gate1053(.a(G1237), .b(G1236), .O(gate487inter2));
  inv1  gate1054(.a(s_72), .O(gate487inter3));
  inv1  gate1055(.a(s_73), .O(gate487inter4));
  nand2 gate1056(.a(gate487inter4), .b(gate487inter3), .O(gate487inter5));
  nor2  gate1057(.a(gate487inter5), .b(gate487inter2), .O(gate487inter6));
  inv1  gate1058(.a(G1236), .O(gate487inter7));
  inv1  gate1059(.a(G1237), .O(gate487inter8));
  nand2 gate1060(.a(gate487inter8), .b(gate487inter7), .O(gate487inter9));
  nand2 gate1061(.a(s_73), .b(gate487inter3), .O(gate487inter10));
  nor2  gate1062(.a(gate487inter10), .b(gate487inter9), .O(gate487inter11));
  nor2  gate1063(.a(gate487inter11), .b(gate487inter6), .O(gate487inter12));
  nand2 gate1064(.a(gate487inter12), .b(gate487inter1), .O(G1296));
nand2 gate488( .a(G1238), .b(G1239), .O(G1297) );

  xor2  gate617(.a(G1241), .b(G1240), .O(gate489inter0));
  nand2 gate618(.a(gate489inter0), .b(s_10), .O(gate489inter1));
  and2  gate619(.a(G1241), .b(G1240), .O(gate489inter2));
  inv1  gate620(.a(s_10), .O(gate489inter3));
  inv1  gate621(.a(s_11), .O(gate489inter4));
  nand2 gate622(.a(gate489inter4), .b(gate489inter3), .O(gate489inter5));
  nor2  gate623(.a(gate489inter5), .b(gate489inter2), .O(gate489inter6));
  inv1  gate624(.a(G1240), .O(gate489inter7));
  inv1  gate625(.a(G1241), .O(gate489inter8));
  nand2 gate626(.a(gate489inter8), .b(gate489inter7), .O(gate489inter9));
  nand2 gate627(.a(s_11), .b(gate489inter3), .O(gate489inter10));
  nor2  gate628(.a(gate489inter10), .b(gate489inter9), .O(gate489inter11));
  nor2  gate629(.a(gate489inter11), .b(gate489inter6), .O(gate489inter12));
  nand2 gate630(.a(gate489inter12), .b(gate489inter1), .O(G1298));
nand2 gate490( .a(G1242), .b(G1243), .O(G1299) );
nand2 gate491( .a(G1244), .b(G1245), .O(G1300) );
nand2 gate492( .a(G1246), .b(G1247), .O(G1301) );
nand2 gate493( .a(G1248), .b(G1249), .O(G1302) );
nand2 gate494( .a(G1250), .b(G1251), .O(G1303) );

  xor2  gate1779(.a(G1253), .b(G1252), .O(gate495inter0));
  nand2 gate1780(.a(gate495inter0), .b(s_176), .O(gate495inter1));
  and2  gate1781(.a(G1253), .b(G1252), .O(gate495inter2));
  inv1  gate1782(.a(s_176), .O(gate495inter3));
  inv1  gate1783(.a(s_177), .O(gate495inter4));
  nand2 gate1784(.a(gate495inter4), .b(gate495inter3), .O(gate495inter5));
  nor2  gate1785(.a(gate495inter5), .b(gate495inter2), .O(gate495inter6));
  inv1  gate1786(.a(G1252), .O(gate495inter7));
  inv1  gate1787(.a(G1253), .O(gate495inter8));
  nand2 gate1788(.a(gate495inter8), .b(gate495inter7), .O(gate495inter9));
  nand2 gate1789(.a(s_177), .b(gate495inter3), .O(gate495inter10));
  nor2  gate1790(.a(gate495inter10), .b(gate495inter9), .O(gate495inter11));
  nor2  gate1791(.a(gate495inter11), .b(gate495inter6), .O(gate495inter12));
  nand2 gate1792(.a(gate495inter12), .b(gate495inter1), .O(G1304));
nand2 gate496( .a(G1254), .b(G1255), .O(G1305) );

  xor2  gate1303(.a(G1257), .b(G1256), .O(gate497inter0));
  nand2 gate1304(.a(gate497inter0), .b(s_108), .O(gate497inter1));
  and2  gate1305(.a(G1257), .b(G1256), .O(gate497inter2));
  inv1  gate1306(.a(s_108), .O(gate497inter3));
  inv1  gate1307(.a(s_109), .O(gate497inter4));
  nand2 gate1308(.a(gate497inter4), .b(gate497inter3), .O(gate497inter5));
  nor2  gate1309(.a(gate497inter5), .b(gate497inter2), .O(gate497inter6));
  inv1  gate1310(.a(G1256), .O(gate497inter7));
  inv1  gate1311(.a(G1257), .O(gate497inter8));
  nand2 gate1312(.a(gate497inter8), .b(gate497inter7), .O(gate497inter9));
  nand2 gate1313(.a(s_109), .b(gate497inter3), .O(gate497inter10));
  nor2  gate1314(.a(gate497inter10), .b(gate497inter9), .O(gate497inter11));
  nor2  gate1315(.a(gate497inter11), .b(gate497inter6), .O(gate497inter12));
  nand2 gate1316(.a(gate497inter12), .b(gate497inter1), .O(G1306));
nand2 gate498( .a(G1258), .b(G1259), .O(G1307) );

  xor2  gate1639(.a(G1261), .b(G1260), .O(gate499inter0));
  nand2 gate1640(.a(gate499inter0), .b(s_156), .O(gate499inter1));
  and2  gate1641(.a(G1261), .b(G1260), .O(gate499inter2));
  inv1  gate1642(.a(s_156), .O(gate499inter3));
  inv1  gate1643(.a(s_157), .O(gate499inter4));
  nand2 gate1644(.a(gate499inter4), .b(gate499inter3), .O(gate499inter5));
  nor2  gate1645(.a(gate499inter5), .b(gate499inter2), .O(gate499inter6));
  inv1  gate1646(.a(G1260), .O(gate499inter7));
  inv1  gate1647(.a(G1261), .O(gate499inter8));
  nand2 gate1648(.a(gate499inter8), .b(gate499inter7), .O(gate499inter9));
  nand2 gate1649(.a(s_157), .b(gate499inter3), .O(gate499inter10));
  nor2  gate1650(.a(gate499inter10), .b(gate499inter9), .O(gate499inter11));
  nor2  gate1651(.a(gate499inter11), .b(gate499inter6), .O(gate499inter12));
  nand2 gate1652(.a(gate499inter12), .b(gate499inter1), .O(G1308));
nand2 gate500( .a(G1262), .b(G1263), .O(G1309) );
nand2 gate501( .a(G1264), .b(G1265), .O(G1310) );

  xor2  gate841(.a(G1267), .b(G1266), .O(gate502inter0));
  nand2 gate842(.a(gate502inter0), .b(s_42), .O(gate502inter1));
  and2  gate843(.a(G1267), .b(G1266), .O(gate502inter2));
  inv1  gate844(.a(s_42), .O(gate502inter3));
  inv1  gate845(.a(s_43), .O(gate502inter4));
  nand2 gate846(.a(gate502inter4), .b(gate502inter3), .O(gate502inter5));
  nor2  gate847(.a(gate502inter5), .b(gate502inter2), .O(gate502inter6));
  inv1  gate848(.a(G1266), .O(gate502inter7));
  inv1  gate849(.a(G1267), .O(gate502inter8));
  nand2 gate850(.a(gate502inter8), .b(gate502inter7), .O(gate502inter9));
  nand2 gate851(.a(s_43), .b(gate502inter3), .O(gate502inter10));
  nor2  gate852(.a(gate502inter10), .b(gate502inter9), .O(gate502inter11));
  nor2  gate853(.a(gate502inter11), .b(gate502inter6), .O(gate502inter12));
  nand2 gate854(.a(gate502inter12), .b(gate502inter1), .O(G1311));
nand2 gate503( .a(G1268), .b(G1269), .O(G1312) );

  xor2  gate1611(.a(G1271), .b(G1270), .O(gate504inter0));
  nand2 gate1612(.a(gate504inter0), .b(s_152), .O(gate504inter1));
  and2  gate1613(.a(G1271), .b(G1270), .O(gate504inter2));
  inv1  gate1614(.a(s_152), .O(gate504inter3));
  inv1  gate1615(.a(s_153), .O(gate504inter4));
  nand2 gate1616(.a(gate504inter4), .b(gate504inter3), .O(gate504inter5));
  nor2  gate1617(.a(gate504inter5), .b(gate504inter2), .O(gate504inter6));
  inv1  gate1618(.a(G1270), .O(gate504inter7));
  inv1  gate1619(.a(G1271), .O(gate504inter8));
  nand2 gate1620(.a(gate504inter8), .b(gate504inter7), .O(gate504inter9));
  nand2 gate1621(.a(s_153), .b(gate504inter3), .O(gate504inter10));
  nor2  gate1622(.a(gate504inter10), .b(gate504inter9), .O(gate504inter11));
  nor2  gate1623(.a(gate504inter11), .b(gate504inter6), .O(gate504inter12));
  nand2 gate1624(.a(gate504inter12), .b(gate504inter1), .O(G1313));

  xor2  gate3067(.a(G1273), .b(G1272), .O(gate505inter0));
  nand2 gate3068(.a(gate505inter0), .b(s_360), .O(gate505inter1));
  and2  gate3069(.a(G1273), .b(G1272), .O(gate505inter2));
  inv1  gate3070(.a(s_360), .O(gate505inter3));
  inv1  gate3071(.a(s_361), .O(gate505inter4));
  nand2 gate3072(.a(gate505inter4), .b(gate505inter3), .O(gate505inter5));
  nor2  gate3073(.a(gate505inter5), .b(gate505inter2), .O(gate505inter6));
  inv1  gate3074(.a(G1272), .O(gate505inter7));
  inv1  gate3075(.a(G1273), .O(gate505inter8));
  nand2 gate3076(.a(gate505inter8), .b(gate505inter7), .O(gate505inter9));
  nand2 gate3077(.a(s_361), .b(gate505inter3), .O(gate505inter10));
  nor2  gate3078(.a(gate505inter10), .b(gate505inter9), .O(gate505inter11));
  nor2  gate3079(.a(gate505inter11), .b(gate505inter6), .O(gate505inter12));
  nand2 gate3080(.a(gate505inter12), .b(gate505inter1), .O(G1314));
nand2 gate506( .a(G1274), .b(G1275), .O(G1315) );
nand2 gate507( .a(G1276), .b(G1277), .O(G1316) );

  xor2  gate827(.a(G1279), .b(G1278), .O(gate508inter0));
  nand2 gate828(.a(gate508inter0), .b(s_40), .O(gate508inter1));
  and2  gate829(.a(G1279), .b(G1278), .O(gate508inter2));
  inv1  gate830(.a(s_40), .O(gate508inter3));
  inv1  gate831(.a(s_41), .O(gate508inter4));
  nand2 gate832(.a(gate508inter4), .b(gate508inter3), .O(gate508inter5));
  nor2  gate833(.a(gate508inter5), .b(gate508inter2), .O(gate508inter6));
  inv1  gate834(.a(G1278), .O(gate508inter7));
  inv1  gate835(.a(G1279), .O(gate508inter8));
  nand2 gate836(.a(gate508inter8), .b(gate508inter7), .O(gate508inter9));
  nand2 gate837(.a(s_41), .b(gate508inter3), .O(gate508inter10));
  nor2  gate838(.a(gate508inter10), .b(gate508inter9), .O(gate508inter11));
  nor2  gate839(.a(gate508inter11), .b(gate508inter6), .O(gate508inter12));
  nand2 gate840(.a(gate508inter12), .b(gate508inter1), .O(G1317));
nand2 gate509( .a(G1280), .b(G1281), .O(G1318) );

  xor2  gate2689(.a(G1283), .b(G1282), .O(gate510inter0));
  nand2 gate2690(.a(gate510inter0), .b(s_306), .O(gate510inter1));
  and2  gate2691(.a(G1283), .b(G1282), .O(gate510inter2));
  inv1  gate2692(.a(s_306), .O(gate510inter3));
  inv1  gate2693(.a(s_307), .O(gate510inter4));
  nand2 gate2694(.a(gate510inter4), .b(gate510inter3), .O(gate510inter5));
  nor2  gate2695(.a(gate510inter5), .b(gate510inter2), .O(gate510inter6));
  inv1  gate2696(.a(G1282), .O(gate510inter7));
  inv1  gate2697(.a(G1283), .O(gate510inter8));
  nand2 gate2698(.a(gate510inter8), .b(gate510inter7), .O(gate510inter9));
  nand2 gate2699(.a(s_307), .b(gate510inter3), .O(gate510inter10));
  nor2  gate2700(.a(gate510inter10), .b(gate510inter9), .O(gate510inter11));
  nor2  gate2701(.a(gate510inter11), .b(gate510inter6), .O(gate510inter12));
  nand2 gate2702(.a(gate510inter12), .b(gate510inter1), .O(G1319));

  xor2  gate2143(.a(G1285), .b(G1284), .O(gate511inter0));
  nand2 gate2144(.a(gate511inter0), .b(s_228), .O(gate511inter1));
  and2  gate2145(.a(G1285), .b(G1284), .O(gate511inter2));
  inv1  gate2146(.a(s_228), .O(gate511inter3));
  inv1  gate2147(.a(s_229), .O(gate511inter4));
  nand2 gate2148(.a(gate511inter4), .b(gate511inter3), .O(gate511inter5));
  nor2  gate2149(.a(gate511inter5), .b(gate511inter2), .O(gate511inter6));
  inv1  gate2150(.a(G1284), .O(gate511inter7));
  inv1  gate2151(.a(G1285), .O(gate511inter8));
  nand2 gate2152(.a(gate511inter8), .b(gate511inter7), .O(gate511inter9));
  nand2 gate2153(.a(s_229), .b(gate511inter3), .O(gate511inter10));
  nor2  gate2154(.a(gate511inter10), .b(gate511inter9), .O(gate511inter11));
  nor2  gate2155(.a(gate511inter11), .b(gate511inter6), .O(gate511inter12));
  nand2 gate2156(.a(gate511inter12), .b(gate511inter1), .O(G1320));
nand2 gate512( .a(G1286), .b(G1287), .O(G1321) );

  xor2  gate2899(.a(G1289), .b(G1288), .O(gate513inter0));
  nand2 gate2900(.a(gate513inter0), .b(s_336), .O(gate513inter1));
  and2  gate2901(.a(G1289), .b(G1288), .O(gate513inter2));
  inv1  gate2902(.a(s_336), .O(gate513inter3));
  inv1  gate2903(.a(s_337), .O(gate513inter4));
  nand2 gate2904(.a(gate513inter4), .b(gate513inter3), .O(gate513inter5));
  nor2  gate2905(.a(gate513inter5), .b(gate513inter2), .O(gate513inter6));
  inv1  gate2906(.a(G1288), .O(gate513inter7));
  inv1  gate2907(.a(G1289), .O(gate513inter8));
  nand2 gate2908(.a(gate513inter8), .b(gate513inter7), .O(gate513inter9));
  nand2 gate2909(.a(s_337), .b(gate513inter3), .O(gate513inter10));
  nor2  gate2910(.a(gate513inter10), .b(gate513inter9), .O(gate513inter11));
  nor2  gate2911(.a(gate513inter11), .b(gate513inter6), .O(gate513inter12));
  nand2 gate2912(.a(gate513inter12), .b(gate513inter1), .O(G1322));

  xor2  gate3123(.a(G1291), .b(G1290), .O(gate514inter0));
  nand2 gate3124(.a(gate514inter0), .b(s_368), .O(gate514inter1));
  and2  gate3125(.a(G1291), .b(G1290), .O(gate514inter2));
  inv1  gate3126(.a(s_368), .O(gate514inter3));
  inv1  gate3127(.a(s_369), .O(gate514inter4));
  nand2 gate3128(.a(gate514inter4), .b(gate514inter3), .O(gate514inter5));
  nor2  gate3129(.a(gate514inter5), .b(gate514inter2), .O(gate514inter6));
  inv1  gate3130(.a(G1290), .O(gate514inter7));
  inv1  gate3131(.a(G1291), .O(gate514inter8));
  nand2 gate3132(.a(gate514inter8), .b(gate514inter7), .O(gate514inter9));
  nand2 gate3133(.a(s_369), .b(gate514inter3), .O(gate514inter10));
  nor2  gate3134(.a(gate514inter10), .b(gate514inter9), .O(gate514inter11));
  nor2  gate3135(.a(gate514inter11), .b(gate514inter6), .O(gate514inter12));
  nand2 gate3136(.a(gate514inter12), .b(gate514inter1), .O(G1323));
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule