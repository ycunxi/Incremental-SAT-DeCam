module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);

input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;//RE__PI;

input s_0,s_1;//RE__ALLOW(00,01,10,11);
input s_2,s_3;//RE__ALLOW(00,01,10,11);
input s_4,s_5;//RE__ALLOW(00,01,10,11);
input s_6,s_7;//RE__ALLOW(00,01,10,11);
input s_8,s_9;//RE__ALLOW(00,01,10,11);
input s_10,s_11;//RE__ALLOW(00,01,10,11);
input s_12,s_13;//RE__ALLOW(00,01,10,11);
input s_14,s_15;//RE__ALLOW(00,01,10,11);
input s_16,s_17;//RE__ALLOW(00,01,10,11);
input s_18,s_19;//RE__ALLOW(00,01,10,11);
input s_20,s_21;//RE__ALLOW(00,01,10,11);
input s_22,s_23;//RE__ALLOW(00,01,10,11);
input s_24,s_25;//RE__ALLOW(00,01,10,11);
input s_26,s_27;//RE__ALLOW(00,01,10,11);
input s_28,s_29;//RE__ALLOW(00,01,10,11);
input s_30,s_31;//RE__ALLOW(00,01,10,11);
input s_32,s_33;//RE__ALLOW(00,01,10,11);
input s_34,s_35;//RE__ALLOW(00,01,10,11);
input s_36,s_37;//RE__ALLOW(00,01,10,11);
input s_38,s_39;//RE__ALLOW(00,01,10,11);
input s_40,s_41;//RE__ALLOW(00,01,10,11);
input s_42,s_43;//RE__ALLOW(00,01,10,11);
input s_44,s_45;//RE__ALLOW(00,01,10,11);
input s_46,s_47;//RE__ALLOW(00,01,10,11);
input s_48,s_49;//RE__ALLOW(00,01,10,11);
input s_50,s_51;//RE__ALLOW(00,01,10,11);
input s_52,s_53;//RE__ALLOW(00,01,10,11);
input s_54,s_55;//RE__ALLOW(00,01,10,11);
input s_56,s_57;//RE__ALLOW(00,01,10,11);
input s_58,s_59;//RE__ALLOW(00,01,10,11);
input s_60,s_61;//RE__ALLOW(00,01,10,11);
input s_62,s_63;//RE__ALLOW(00,01,10,11);
input s_64,s_65;//RE__ALLOW(00,01,10,11);
input s_66,s_67;//RE__ALLOW(00,01,10,11);
input s_68,s_69;//RE__ALLOW(00,01,10,11);
input s_70,s_71;//RE__ALLOW(00,01,10,11);
input s_72,s_73;//RE__ALLOW(00,01,10,11);
input s_74,s_75;//RE__ALLOW(00,01,10,11);
input s_76,s_77;//RE__ALLOW(00,01,10,11);
input s_78,s_79;//RE__ALLOW(00,01,10,11);
input s_80,s_81;//RE__ALLOW(00,01,10,11);
input s_82,s_83;//RE__ALLOW(00,01,10,11);
input s_84,s_85;//RE__ALLOW(00,01,10,11);
input s_86,s_87;//RE__ALLOW(00,01,10,11);
input s_88,s_89;//RE__ALLOW(00,01,10,11);
input s_90,s_91;//RE__ALLOW(00,01,10,11);
input s_92,s_93;//RE__ALLOW(00,01,10,11);
input s_94,s_95;//RE__ALLOW(00,01,10,11);
input s_96,s_97;//RE__ALLOW(00,01,10,11);
input s_98,s_99;//RE__ALLOW(00,01,10,11);
input s_100,s_101;//RE__ALLOW(00,01,10,11);
input s_102,s_103;//RE__ALLOW(00,01,10,11);
input s_104,s_105;//RE__ALLOW(00,01,10,11);
input s_106,s_107;//RE__ALLOW(00,01,10,11);
input s_108,s_109;//RE__ALLOW(00,01,10,11);
input s_110,s_111;//RE__ALLOW(00,01,10,11);
input s_112,s_113;//RE__ALLOW(00,01,10,11);
input s_114,s_115;//RE__ALLOW(00,01,10,11);
input s_116,s_117;//RE__ALLOW(00,01,10,11);
input s_118,s_119;//RE__ALLOW(00,01,10,11);
input s_120,s_121;//RE__ALLOW(00,01,10,11);
input s_122,s_123;//RE__ALLOW(00,01,10,11);
input s_124,s_125;//RE__ALLOW(00,01,10,11);
input s_126,s_127;//RE__ALLOW(00,01,10,11);
input s_128,s_129;//RE__ALLOW(00,01,10,11);
input s_130,s_131;//RE__ALLOW(00,01,10,11);
input s_132,s_133;//RE__ALLOW(00,01,10,11);
input s_134,s_135;//RE__ALLOW(00,01,10,11);
input s_136,s_137;//RE__ALLOW(00,01,10,11);
input s_138,s_139;//RE__ALLOW(00,01,10,11);
input s_140,s_141;//RE__ALLOW(00,01,10,11);
input s_142,s_143;//RE__ALLOW(00,01,10,11);
input s_144,s_145;//RE__ALLOW(00,01,10,11);
input s_146,s_147;//RE__ALLOW(00,01,10,11);
input s_148,s_149;//RE__ALLOW(00,01,10,11);
input s_150,s_151;//RE__ALLOW(00,01,10,11);
input s_152,s_153;//RE__ALLOW(00,01,10,11);
input s_154,s_155;//RE__ALLOW(00,01,10,11);
input s_156,s_157;//RE__ALLOW(00,01,10,11);
input s_158,s_159;//RE__ALLOW(00,01,10,11);
input s_160,s_161;//RE__ALLOW(00,01,10,11);
input s_162,s_163;//RE__ALLOW(00,01,10,11);
input s_164,s_165;//RE__ALLOW(00,01,10,11);
input s_166,s_167;//RE__ALLOW(00,01,10,11);
input s_168,s_169;//RE__ALLOW(00,01,10,11);
input s_170,s_171;//RE__ALLOW(00,01,10,11);
input s_172,s_173;//RE__ALLOW(00,01,10,11);
input s_174,s_175;//RE__ALLOW(00,01,10,11);
input s_176,s_177;//RE__ALLOW(00,01,10,11);
input s_178,s_179;//RE__ALLOW(00,01,10,11);
input s_180,s_181;//RE__ALLOW(00,01,10,11);
input s_182,s_183;//RE__ALLOW(00,01,10,11);
input s_184,s_185;//RE__ALLOW(00,01,10,11);
input s_186,s_187;//RE__ALLOW(00,01,10,11);
input s_188,s_189;//RE__ALLOW(00,01,10,11);
input s_190,s_191;//RE__ALLOW(00,01,10,11);
input s_192,s_193;//RE__ALLOW(00,01,10,11);
input s_194,s_195;//RE__ALLOW(00,01,10,11);
input s_196,s_197;//RE__ALLOW(00,01,10,11);
input s_198,s_199;//RE__ALLOW(00,01,10,11);
input s_200,s_201;//RE__ALLOW(00,01,10,11);
input s_202,s_203;//RE__ALLOW(00,01,10,11);
input s_204,s_205;//RE__ALLOW(00,01,10,11);
input s_206,s_207;//RE__ALLOW(00,01,10,11);
input s_208,s_209;//RE__ALLOW(00,01,10,11);
input s_210,s_211;//RE__ALLOW(00,01,10,11);
input s_212,s_213;//RE__ALLOW(00,01,10,11);
input s_214,s_215;//RE__ALLOW(00,01,10,11);
input s_216,s_217;//RE__ALLOW(00,01,10,11);
input s_218,s_219;//RE__ALLOW(00,01,10,11);
input s_220,s_221;//RE__ALLOW(00,01,10,11);
input s_222,s_223;//RE__ALLOW(00,01,10,11);
input s_224,s_225;//RE__ALLOW(00,01,10,11);
input s_226,s_227;//RE__ALLOW(00,01,10,11);
input s_228,s_229;//RE__ALLOW(00,01,10,11);
input s_230,s_231;//RE__ALLOW(00,01,10,11);
input s_232,s_233;//RE__ALLOW(00,01,10,11);
input s_234,s_235;//RE__ALLOW(00,01,10,11);
input s_236,s_237;//RE__ALLOW(00,01,10,11);
input s_238,s_239;//RE__ALLOW(00,01,10,11);
input s_240,s_241;//RE__ALLOW(00,01,10,11);
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;

  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate215inter0, gate215inter1, gate215inter2, gate215inter3, gate215inter4, gate215inter5, gate215inter6, gate215inter7, gate215inter8, gate215inter9, gate215inter10, gate215inter11, gate215inter12, gate289inter0, gate289inter1, gate289inter2, gate289inter3, gate289inter4, gate289inter5, gate289inter6, gate289inter7, gate289inter8, gate289inter9, gate289inter10, gate289inter11, gate289inter12, gate110inter0, gate110inter1, gate110inter2, gate110inter3, gate110inter4, gate110inter5, gate110inter6, gate110inter7, gate110inter8, gate110inter9, gate110inter10, gate110inter11, gate110inter12, gate196inter0, gate196inter1, gate196inter2, gate196inter3, gate196inter4, gate196inter5, gate196inter6, gate196inter7, gate196inter8, gate196inter9, gate196inter10, gate196inter11, gate196inter12, gate485inter0, gate485inter1, gate485inter2, gate485inter3, gate485inter4, gate485inter5, gate485inter6, gate485inter7, gate485inter8, gate485inter9, gate485inter10, gate485inter11, gate485inter12, gate112inter0, gate112inter1, gate112inter2, gate112inter3, gate112inter4, gate112inter5, gate112inter6, gate112inter7, gate112inter8, gate112inter9, gate112inter10, gate112inter11, gate112inter12, gate439inter0, gate439inter1, gate439inter2, gate439inter3, gate439inter4, gate439inter5, gate439inter6, gate439inter7, gate439inter8, gate439inter9, gate439inter10, gate439inter11, gate439inter12, gate134inter0, gate134inter1, gate134inter2, gate134inter3, gate134inter4, gate134inter5, gate134inter6, gate134inter7, gate134inter8, gate134inter9, gate134inter10, gate134inter11, gate134inter12, gate474inter0, gate474inter1, gate474inter2, gate474inter3, gate474inter4, gate474inter5, gate474inter6, gate474inter7, gate474inter8, gate474inter9, gate474inter10, gate474inter11, gate474inter12, gate453inter0, gate453inter1, gate453inter2, gate453inter3, gate453inter4, gate453inter5, gate453inter6, gate453inter7, gate453inter8, gate453inter9, gate453inter10, gate453inter11, gate453inter12, gate114inter0, gate114inter1, gate114inter2, gate114inter3, gate114inter4, gate114inter5, gate114inter6, gate114inter7, gate114inter8, gate114inter9, gate114inter10, gate114inter11, gate114inter12, gate18inter0, gate18inter1, gate18inter2, gate18inter3, gate18inter4, gate18inter5, gate18inter6, gate18inter7, gate18inter8, gate18inter9, gate18inter10, gate18inter11, gate18inter12, gate262inter0, gate262inter1, gate262inter2, gate262inter3, gate262inter4, gate262inter5, gate262inter6, gate262inter7, gate262inter8, gate262inter9, gate262inter10, gate262inter11, gate262inter12, gate14inter0, gate14inter1, gate14inter2, gate14inter3, gate14inter4, gate14inter5, gate14inter6, gate14inter7, gate14inter8, gate14inter9, gate14inter10, gate14inter11, gate14inter12, gate82inter0, gate82inter1, gate82inter2, gate82inter3, gate82inter4, gate82inter5, gate82inter6, gate82inter7, gate82inter8, gate82inter9, gate82inter10, gate82inter11, gate82inter12, gate125inter0, gate125inter1, gate125inter2, gate125inter3, gate125inter4, gate125inter5, gate125inter6, gate125inter7, gate125inter8, gate125inter9, gate125inter10, gate125inter11, gate125inter12, gate280inter0, gate280inter1, gate280inter2, gate280inter3, gate280inter4, gate280inter5, gate280inter6, gate280inter7, gate280inter8, gate280inter9, gate280inter10, gate280inter11, gate280inter12, gate444inter0, gate444inter1, gate444inter2, gate444inter3, gate444inter4, gate444inter5, gate444inter6, gate444inter7, gate444inter8, gate444inter9, gate444inter10, gate444inter11, gate444inter12, gate443inter0, gate443inter1, gate443inter2, gate443inter3, gate443inter4, gate443inter5, gate443inter6, gate443inter7, gate443inter8, gate443inter9, gate443inter10, gate443inter11, gate443inter12, gate29inter0, gate29inter1, gate29inter2, gate29inter3, gate29inter4, gate29inter5, gate29inter6, gate29inter7, gate29inter8, gate29inter9, gate29inter10, gate29inter11, gate29inter12, gate165inter0, gate165inter1, gate165inter2, gate165inter3, gate165inter4, gate165inter5, gate165inter6, gate165inter7, gate165inter8, gate165inter9, gate165inter10, gate165inter11, gate165inter12, gate87inter0, gate87inter1, gate87inter2, gate87inter3, gate87inter4, gate87inter5, gate87inter6, gate87inter7, gate87inter8, gate87inter9, gate87inter10, gate87inter11, gate87inter12, gate410inter0, gate410inter1, gate410inter2, gate410inter3, gate410inter4, gate410inter5, gate410inter6, gate410inter7, gate410inter8, gate410inter9, gate410inter10, gate410inter11, gate410inter12, gate164inter0, gate164inter1, gate164inter2, gate164inter3, gate164inter4, gate164inter5, gate164inter6, gate164inter7, gate164inter8, gate164inter9, gate164inter10, gate164inter11, gate164inter12, gate12inter0, gate12inter1, gate12inter2, gate12inter3, gate12inter4, gate12inter5, gate12inter6, gate12inter7, gate12inter8, gate12inter9, gate12inter10, gate12inter11, gate12inter12, gate217inter0, gate217inter1, gate217inter2, gate217inter3, gate217inter4, gate217inter5, gate217inter6, gate217inter7, gate217inter8, gate217inter9, gate217inter10, gate217inter11, gate217inter12, gate104inter0, gate104inter1, gate104inter2, gate104inter3, gate104inter4, gate104inter5, gate104inter6, gate104inter7, gate104inter8, gate104inter9, gate104inter10, gate104inter11, gate104inter12, gate184inter0, gate184inter1, gate184inter2, gate184inter3, gate184inter4, gate184inter5, gate184inter6, gate184inter7, gate184inter8, gate184inter9, gate184inter10, gate184inter11, gate184inter12, gate287inter0, gate287inter1, gate287inter2, gate287inter3, gate287inter4, gate287inter5, gate287inter6, gate287inter7, gate287inter8, gate287inter9, gate287inter10, gate287inter11, gate287inter12, gate175inter0, gate175inter1, gate175inter2, gate175inter3, gate175inter4, gate175inter5, gate175inter6, gate175inter7, gate175inter8, gate175inter9, gate175inter10, gate175inter11, gate175inter12, gate235inter0, gate235inter1, gate235inter2, gate235inter3, gate235inter4, gate235inter5, gate235inter6, gate235inter7, gate235inter8, gate235inter9, gate235inter10, gate235inter11, gate235inter12, gate268inter0, gate268inter1, gate268inter2, gate268inter3, gate268inter4, gate268inter5, gate268inter6, gate268inter7, gate268inter8, gate268inter9, gate268inter10, gate268inter11, gate268inter12, gate23inter0, gate23inter1, gate23inter2, gate23inter3, gate23inter4, gate23inter5, gate23inter6, gate23inter7, gate23inter8, gate23inter9, gate23inter10, gate23inter11, gate23inter12, gate98inter0, gate98inter1, gate98inter2, gate98inter3, gate98inter4, gate98inter5, gate98inter6, gate98inter7, gate98inter8, gate98inter9, gate98inter10, gate98inter11, gate98inter12, gate154inter0, gate154inter1, gate154inter2, gate154inter3, gate154inter4, gate154inter5, gate154inter6, gate154inter7, gate154inter8, gate154inter9, gate154inter10, gate154inter11, gate154inter12, gate407inter0, gate407inter1, gate407inter2, gate407inter3, gate407inter4, gate407inter5, gate407inter6, gate407inter7, gate407inter8, gate407inter9, gate407inter10, gate407inter11, gate407inter12, gate28inter0, gate28inter1, gate28inter2, gate28inter3, gate28inter4, gate28inter5, gate28inter6, gate28inter7, gate28inter8, gate28inter9, gate28inter10, gate28inter11, gate28inter12, gate90inter0, gate90inter1, gate90inter2, gate90inter3, gate90inter4, gate90inter5, gate90inter6, gate90inter7, gate90inter8, gate90inter9, gate90inter10, gate90inter11, gate90inter12, gate185inter0, gate185inter1, gate185inter2, gate185inter3, gate185inter4, gate185inter5, gate185inter6, gate185inter7, gate185inter8, gate185inter9, gate185inter10, gate185inter11, gate185inter12, gate480inter0, gate480inter1, gate480inter2, gate480inter3, gate480inter4, gate480inter5, gate480inter6, gate480inter7, gate480inter8, gate480inter9, gate480inter10, gate480inter11, gate480inter12, gate210inter0, gate210inter1, gate210inter2, gate210inter3, gate210inter4, gate210inter5, gate210inter6, gate210inter7, gate210inter8, gate210inter9, gate210inter10, gate210inter11, gate210inter12, gate488inter0, gate488inter1, gate488inter2, gate488inter3, gate488inter4, gate488inter5, gate488inter6, gate488inter7, gate488inter8, gate488inter9, gate488inter10, gate488inter11, gate488inter12, gate44inter0, gate44inter1, gate44inter2, gate44inter3, gate44inter4, gate44inter5, gate44inter6, gate44inter7, gate44inter8, gate44inter9, gate44inter10, gate44inter11, gate44inter12, gate413inter0, gate413inter1, gate413inter2, gate413inter3, gate413inter4, gate413inter5, gate413inter6, gate413inter7, gate413inter8, gate413inter9, gate413inter10, gate413inter11, gate413inter12, gate115inter0, gate115inter1, gate115inter2, gate115inter3, gate115inter4, gate115inter5, gate115inter6, gate115inter7, gate115inter8, gate115inter9, gate115inter10, gate115inter11, gate115inter12, gate121inter0, gate121inter1, gate121inter2, gate121inter3, gate121inter4, gate121inter5, gate121inter6, gate121inter7, gate121inter8, gate121inter9, gate121inter10, gate121inter11, gate121inter12, gate92inter0, gate92inter1, gate92inter2, gate92inter3, gate92inter4, gate92inter5, gate92inter6, gate92inter7, gate92inter8, gate92inter9, gate92inter10, gate92inter11, gate92inter12, gate391inter0, gate391inter1, gate391inter2, gate391inter3, gate391inter4, gate391inter5, gate391inter6, gate391inter7, gate391inter8, gate391inter9, gate391inter10, gate391inter11, gate391inter12, gate27inter0, gate27inter1, gate27inter2, gate27inter3, gate27inter4, gate27inter5, gate27inter6, gate27inter7, gate27inter8, gate27inter9, gate27inter10, gate27inter11, gate27inter12, gate501inter0, gate501inter1, gate501inter2, gate501inter3, gate501inter4, gate501inter5, gate501inter6, gate501inter7, gate501inter8, gate501inter9, gate501inter10, gate501inter11, gate501inter12, gate414inter0, gate414inter1, gate414inter2, gate414inter3, gate414inter4, gate414inter5, gate414inter6, gate414inter7, gate414inter8, gate414inter9, gate414inter10, gate414inter11, gate414inter12, gate397inter0, gate397inter1, gate397inter2, gate397inter3, gate397inter4, gate397inter5, gate397inter6, gate397inter7, gate397inter8, gate397inter9, gate397inter10, gate397inter11, gate397inter12, gate435inter0, gate435inter1, gate435inter2, gate435inter3, gate435inter4, gate435inter5, gate435inter6, gate435inter7, gate435inter8, gate435inter9, gate435inter10, gate435inter11, gate435inter12, gate194inter0, gate194inter1, gate194inter2, gate194inter3, gate194inter4, gate194inter5, gate194inter6, gate194inter7, gate194inter8, gate194inter9, gate194inter10, gate194inter11, gate194inter12, gate511inter0, gate511inter1, gate511inter2, gate511inter3, gate511inter4, gate511inter5, gate511inter6, gate511inter7, gate511inter8, gate511inter9, gate511inter10, gate511inter11, gate511inter12, gate89inter0, gate89inter1, gate89inter2, gate89inter3, gate89inter4, gate89inter5, gate89inter6, gate89inter7, gate89inter8, gate89inter9, gate89inter10, gate89inter11, gate89inter12, gate79inter0, gate79inter1, gate79inter2, gate79inter3, gate79inter4, gate79inter5, gate79inter6, gate79inter7, gate79inter8, gate79inter9, gate79inter10, gate79inter11, gate79inter12, gate495inter0, gate495inter1, gate495inter2, gate495inter3, gate495inter4, gate495inter5, gate495inter6, gate495inter7, gate495inter8, gate495inter9, gate495inter10, gate495inter11, gate495inter12, gate67inter0, gate67inter1, gate67inter2, gate67inter3, gate67inter4, gate67inter5, gate67inter6, gate67inter7, gate67inter8, gate67inter9, gate67inter10, gate67inter11, gate67inter12, gate230inter0, gate230inter1, gate230inter2, gate230inter3, gate230inter4, gate230inter5, gate230inter6, gate230inter7, gate230inter8, gate230inter9, gate230inter10, gate230inter11, gate230inter12, gate469inter0, gate469inter1, gate469inter2, gate469inter3, gate469inter4, gate469inter5, gate469inter6, gate469inter7, gate469inter8, gate469inter9, gate469inter10, gate469inter11, gate469inter12, gate206inter0, gate206inter1, gate206inter2, gate206inter3, gate206inter4, gate206inter5, gate206inter6, gate206inter7, gate206inter8, gate206inter9, gate206inter10, gate206inter11, gate206inter12, gate246inter0, gate246inter1, gate246inter2, gate246inter3, gate246inter4, gate246inter5, gate246inter6, gate246inter7, gate246inter8, gate246inter9, gate246inter10, gate246inter11, gate246inter12, gate45inter0, gate45inter1, gate45inter2, gate45inter3, gate45inter4, gate45inter5, gate45inter6, gate45inter7, gate45inter8, gate45inter9, gate45inter10, gate45inter11, gate45inter12, gate133inter0, gate133inter1, gate133inter2, gate133inter3, gate133inter4, gate133inter5, gate133inter6, gate133inter7, gate133inter8, gate133inter9, gate133inter10, gate133inter11, gate133inter12, gate272inter0, gate272inter1, gate272inter2, gate272inter3, gate272inter4, gate272inter5, gate272inter6, gate272inter7, gate272inter8, gate272inter9, gate272inter10, gate272inter11, gate272inter12, gate425inter0, gate425inter1, gate425inter2, gate425inter3, gate425inter4, gate425inter5, gate425inter6, gate425inter7, gate425inter8, gate425inter9, gate425inter10, gate425inter11, gate425inter12, gate465inter0, gate465inter1, gate465inter2, gate465inter3, gate465inter4, gate465inter5, gate465inter6, gate465inter7, gate465inter8, gate465inter9, gate465inter10, gate465inter11, gate465inter12, gate283inter0, gate283inter1, gate283inter2, gate283inter3, gate283inter4, gate283inter5, gate283inter6, gate283inter7, gate283inter8, gate283inter9, gate283inter10, gate283inter11, gate283inter12, gate403inter0, gate403inter1, gate403inter2, gate403inter3, gate403inter4, gate403inter5, gate403inter6, gate403inter7, gate403inter8, gate403inter9, gate403inter10, gate403inter11, gate403inter12, gate105inter0, gate105inter1, gate105inter2, gate105inter3, gate105inter4, gate105inter5, gate105inter6, gate105inter7, gate105inter8, gate105inter9, gate105inter10, gate105inter11, gate105inter12, gate240inter0, gate240inter1, gate240inter2, gate240inter3, gate240inter4, gate240inter5, gate240inter6, gate240inter7, gate240inter8, gate240inter9, gate240inter10, gate240inter11, gate240inter12, gate108inter0, gate108inter1, gate108inter2, gate108inter3, gate108inter4, gate108inter5, gate108inter6, gate108inter7, gate108inter8, gate108inter9, gate108inter10, gate108inter11, gate108inter12, gate220inter0, gate220inter1, gate220inter2, gate220inter3, gate220inter4, gate220inter5, gate220inter6, gate220inter7, gate220inter8, gate220inter9, gate220inter10, gate220inter11, gate220inter12, gate17inter0, gate17inter1, gate17inter2, gate17inter3, gate17inter4, gate17inter5, gate17inter6, gate17inter7, gate17inter8, gate17inter9, gate17inter10, gate17inter11, gate17inter12, gate503inter0, gate503inter1, gate503inter2, gate503inter3, gate503inter4, gate503inter5, gate503inter6, gate503inter7, gate503inter8, gate503inter9, gate503inter10, gate503inter11, gate503inter12, gate253inter0, gate253inter1, gate253inter2, gate253inter3, gate253inter4, gate253inter5, gate253inter6, gate253inter7, gate253inter8, gate253inter9, gate253inter10, gate253inter11, gate253inter12, gate159inter0, gate159inter1, gate159inter2, gate159inter3, gate159inter4, gate159inter5, gate159inter6, gate159inter7, gate159inter8, gate159inter9, gate159inter10, gate159inter11, gate159inter12, gate442inter0, gate442inter1, gate442inter2, gate442inter3, gate442inter4, gate442inter5, gate442inter6, gate442inter7, gate442inter8, gate442inter9, gate442inter10, gate442inter11, gate442inter12, gate214inter0, gate214inter1, gate214inter2, gate214inter3, gate214inter4, gate214inter5, gate214inter6, gate214inter7, gate214inter8, gate214inter9, gate214inter10, gate214inter11, gate214inter12, gate254inter0, gate254inter1, gate254inter2, gate254inter3, gate254inter4, gate254inter5, gate254inter6, gate254inter7, gate254inter8, gate254inter9, gate254inter10, gate254inter11, gate254inter12, gate392inter0, gate392inter1, gate392inter2, gate392inter3, gate392inter4, gate392inter5, gate392inter6, gate392inter7, gate392inter8, gate392inter9, gate392inter10, gate392inter11, gate392inter12, gate514inter0, gate514inter1, gate514inter2, gate514inter3, gate514inter4, gate514inter5, gate514inter6, gate514inter7, gate514inter8, gate514inter9, gate514inter10, gate514inter11, gate514inter12, gate117inter0, gate117inter1, gate117inter2, gate117inter3, gate117inter4, gate117inter5, gate117inter6, gate117inter7, gate117inter8, gate117inter9, gate117inter10, gate117inter11, gate117inter12, gate256inter0, gate256inter1, gate256inter2, gate256inter3, gate256inter4, gate256inter5, gate256inter6, gate256inter7, gate256inter8, gate256inter9, gate256inter10, gate256inter11, gate256inter12, gate234inter0, gate234inter1, gate234inter2, gate234inter3, gate234inter4, gate234inter5, gate234inter6, gate234inter7, gate234inter8, gate234inter9, gate234inter10, gate234inter11, gate234inter12, gate212inter0, gate212inter1, gate212inter2, gate212inter3, gate212inter4, gate212inter5, gate212inter6, gate212inter7, gate212inter8, gate212inter9, gate212inter10, gate212inter11, gate212inter12, gate492inter0, gate492inter1, gate492inter2, gate492inter3, gate492inter4, gate492inter5, gate492inter6, gate492inter7, gate492inter8, gate492inter9, gate492inter10, gate492inter11, gate492inter12, gate266inter0, gate266inter1, gate266inter2, gate266inter3, gate266inter4, gate266inter5, gate266inter6, gate266inter7, gate266inter8, gate266inter9, gate266inter10, gate266inter11, gate266inter12, gate116inter0, gate116inter1, gate116inter2, gate116inter3, gate116inter4, gate116inter5, gate116inter6, gate116inter7, gate116inter8, gate116inter9, gate116inter10, gate116inter11, gate116inter12, gate11inter0, gate11inter1, gate11inter2, gate11inter3, gate11inter4, gate11inter5, gate11inter6, gate11inter7, gate11inter8, gate11inter9, gate11inter10, gate11inter11, gate11inter12, gate257inter0, gate257inter1, gate257inter2, gate257inter3, gate257inter4, gate257inter5, gate257inter6, gate257inter7, gate257inter8, gate257inter9, gate257inter10, gate257inter11, gate257inter12, gate489inter0, gate489inter1, gate489inter2, gate489inter3, gate489inter4, gate489inter5, gate489inter6, gate489inter7, gate489inter8, gate489inter9, gate489inter10, gate489inter11, gate489inter12, gate193inter0, gate193inter1, gate193inter2, gate193inter3, gate193inter4, gate193inter5, gate193inter6, gate193inter7, gate193inter8, gate193inter9, gate193inter10, gate193inter11, gate193inter12, gate491inter0, gate491inter1, gate491inter2, gate491inter3, gate491inter4, gate491inter5, gate491inter6, gate491inter7, gate491inter8, gate491inter9, gate491inter10, gate491inter11, gate491inter12, gate279inter0, gate279inter1, gate279inter2, gate279inter3, gate279inter4, gate279inter5, gate279inter6, gate279inter7, gate279inter8, gate279inter9, gate279inter10, gate279inter11, gate279inter12, gate139inter0, gate139inter1, gate139inter2, gate139inter3, gate139inter4, gate139inter5, gate139inter6, gate139inter7, gate139inter8, gate139inter9, gate139inter10, gate139inter11, gate139inter12, gate441inter0, gate441inter1, gate441inter2, gate441inter3, gate441inter4, gate441inter5, gate441inter6, gate441inter7, gate441inter8, gate441inter9, gate441inter10, gate441inter11, gate441inter12, gate229inter0, gate229inter1, gate229inter2, gate229inter3, gate229inter4, gate229inter5, gate229inter6, gate229inter7, gate229inter8, gate229inter9, gate229inter10, gate229inter11, gate229inter12, gate400inter0, gate400inter1, gate400inter2, gate400inter3, gate400inter4, gate400inter5, gate400inter6, gate400inter7, gate400inter8, gate400inter9, gate400inter10, gate400inter11, gate400inter12, gate72inter0, gate72inter1, gate72inter2, gate72inter3, gate72inter4, gate72inter5, gate72inter6, gate72inter7, gate72inter8, gate72inter9, gate72inter10, gate72inter11, gate72inter12, gate487inter0, gate487inter1, gate487inter2, gate487inter3, gate487inter4, gate487inter5, gate487inter6, gate487inter7, gate487inter8, gate487inter9, gate487inter10, gate487inter11, gate487inter12, gate232inter0, gate232inter1, gate232inter2, gate232inter3, gate232inter4, gate232inter5, gate232inter6, gate232inter7, gate232inter8, gate232inter9, gate232inter10, gate232inter11, gate232inter12, gate77inter0, gate77inter1, gate77inter2, gate77inter3, gate77inter4, gate77inter5, gate77inter6, gate77inter7, gate77inter8, gate77inter9, gate77inter10, gate77inter11, gate77inter12, gate223inter0, gate223inter1, gate223inter2, gate223inter3, gate223inter4, gate223inter5, gate223inter6, gate223inter7, gate223inter8, gate223inter9, gate223inter10, gate223inter11, gate223inter12, gate431inter0, gate431inter1, gate431inter2, gate431inter3, gate431inter4, gate431inter5, gate431inter6, gate431inter7, gate431inter8, gate431inter9, gate431inter10, gate431inter11, gate431inter12, gate454inter0, gate454inter1, gate454inter2, gate454inter3, gate454inter4, gate454inter5, gate454inter6, gate454inter7, gate454inter8, gate454inter9, gate454inter10, gate454inter11, gate454inter12, gate459inter0, gate459inter1, gate459inter2, gate459inter3, gate459inter4, gate459inter5, gate459inter6, gate459inter7, gate459inter8, gate459inter9, gate459inter10, gate459inter11, gate459inter12, gate39inter0, gate39inter1, gate39inter2, gate39inter3, gate39inter4, gate39inter5, gate39inter6, gate39inter7, gate39inter8, gate39inter9, gate39inter10, gate39inter11, gate39inter12, gate396inter0, gate396inter1, gate396inter2, gate396inter3, gate396inter4, gate396inter5, gate396inter6, gate396inter7, gate396inter8, gate396inter9, gate396inter10, gate396inter11, gate396inter12, gate505inter0, gate505inter1, gate505inter2, gate505inter3, gate505inter4, gate505inter5, gate505inter6, gate505inter7, gate505inter8, gate505inter9, gate505inter10, gate505inter11, gate505inter12, gate53inter0, gate53inter1, gate53inter2, gate53inter3, gate53inter4, gate53inter5, gate53inter6, gate53inter7, gate53inter8, gate53inter9, gate53inter10, gate53inter11, gate53inter12, gate123inter0, gate123inter1, gate123inter2, gate123inter3, gate123inter4, gate123inter5, gate123inter6, gate123inter7, gate123inter8, gate123inter9, gate123inter10, gate123inter11, gate123inter12, gate288inter0, gate288inter1, gate288inter2, gate288inter3, gate288inter4, gate288inter5, gate288inter6, gate288inter7, gate288inter8, gate288inter9, gate288inter10, gate288inter11, gate288inter12, gate162inter0, gate162inter1, gate162inter2, gate162inter3, gate162inter4, gate162inter5, gate162inter6, gate162inter7, gate162inter8, gate162inter9, gate162inter10, gate162inter11, gate162inter12, gate415inter0, gate415inter1, gate415inter2, gate415inter3, gate415inter4, gate415inter5, gate415inter6, gate415inter7, gate415inter8, gate415inter9, gate415inter10, gate415inter11, gate415inter12, gate434inter0, gate434inter1, gate434inter2, gate434inter3, gate434inter4, gate434inter5, gate434inter6, gate434inter7, gate434inter8, gate434inter9, gate434inter10, gate434inter11, gate434inter12, gate446inter0, gate446inter1, gate446inter2, gate446inter3, gate446inter4, gate446inter5, gate446inter6, gate446inter7, gate446inter8, gate446inter9, gate446inter10, gate446inter11, gate446inter12, gate142inter0, gate142inter1, gate142inter2, gate142inter3, gate142inter4, gate142inter5, gate142inter6, gate142inter7, gate142inter8, gate142inter9, gate142inter10, gate142inter11, gate142inter12, gate9inter0, gate9inter1, gate9inter2, gate9inter3, gate9inter4, gate9inter5, gate9inter6, gate9inter7, gate9inter8, gate9inter9, gate9inter10, gate9inter11, gate9inter12, gate394inter0, gate394inter1, gate394inter2, gate394inter3, gate394inter4, gate394inter5, gate394inter6, gate394inter7, gate394inter8, gate394inter9, gate394inter10, gate394inter11, gate394inter12;



and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );

  xor2  gate2213(.a(G2), .b(G1), .O(gate9inter0));
  nand2 gate2214(.a(gate9inter0), .b(s_238), .O(gate9inter1));
  and2  gate2215(.a(G2), .b(G1), .O(gate9inter2));
  inv1  gate2216(.a(s_238), .O(gate9inter3));
  inv1  gate2217(.a(s_239), .O(gate9inter4));
  nand2 gate2218(.a(gate9inter4), .b(gate9inter3), .O(gate9inter5));
  nor2  gate2219(.a(gate9inter5), .b(gate9inter2), .O(gate9inter6));
  inv1  gate2220(.a(G1), .O(gate9inter7));
  inv1  gate2221(.a(G2), .O(gate9inter8));
  nand2 gate2222(.a(gate9inter8), .b(gate9inter7), .O(gate9inter9));
  nand2 gate2223(.a(s_239), .b(gate9inter3), .O(gate9inter10));
  nor2  gate2224(.a(gate9inter10), .b(gate9inter9), .O(gate9inter11));
  nor2  gate2225(.a(gate9inter11), .b(gate9inter6), .O(gate9inter12));
  nand2 gate2226(.a(gate9inter12), .b(gate9inter1), .O(G266));
nand2 gate10( .a(G3), .b(G4), .O(G269) );

  xor2  gate1807(.a(G6), .b(G5), .O(gate11inter0));
  nand2 gate1808(.a(gate11inter0), .b(s_180), .O(gate11inter1));
  and2  gate1809(.a(G6), .b(G5), .O(gate11inter2));
  inv1  gate1810(.a(s_180), .O(gate11inter3));
  inv1  gate1811(.a(s_181), .O(gate11inter4));
  nand2 gate1812(.a(gate11inter4), .b(gate11inter3), .O(gate11inter5));
  nor2  gate1813(.a(gate11inter5), .b(gate11inter2), .O(gate11inter6));
  inv1  gate1814(.a(G5), .O(gate11inter7));
  inv1  gate1815(.a(G6), .O(gate11inter8));
  nand2 gate1816(.a(gate11inter8), .b(gate11inter7), .O(gate11inter9));
  nand2 gate1817(.a(s_181), .b(gate11inter3), .O(gate11inter10));
  nor2  gate1818(.a(gate11inter10), .b(gate11inter9), .O(gate11inter11));
  nor2  gate1819(.a(gate11inter11), .b(gate11inter6), .O(gate11inter12));
  nand2 gate1820(.a(gate11inter12), .b(gate11inter1), .O(G272));

  xor2  gate883(.a(G8), .b(G7), .O(gate12inter0));
  nand2 gate884(.a(gate12inter0), .b(s_48), .O(gate12inter1));
  and2  gate885(.a(G8), .b(G7), .O(gate12inter2));
  inv1  gate886(.a(s_48), .O(gate12inter3));
  inv1  gate887(.a(s_49), .O(gate12inter4));
  nand2 gate888(.a(gate12inter4), .b(gate12inter3), .O(gate12inter5));
  nor2  gate889(.a(gate12inter5), .b(gate12inter2), .O(gate12inter6));
  inv1  gate890(.a(G7), .O(gate12inter7));
  inv1  gate891(.a(G8), .O(gate12inter8));
  nand2 gate892(.a(gate12inter8), .b(gate12inter7), .O(gate12inter9));
  nand2 gate893(.a(s_49), .b(gate12inter3), .O(gate12inter10));
  nor2  gate894(.a(gate12inter10), .b(gate12inter9), .O(gate12inter11));
  nor2  gate895(.a(gate12inter11), .b(gate12inter6), .O(gate12inter12));
  nand2 gate896(.a(gate12inter12), .b(gate12inter1), .O(G275));
nand2 gate13( .a(G9), .b(G10), .O(G278) );

  xor2  gate729(.a(G12), .b(G11), .O(gate14inter0));
  nand2 gate730(.a(gate14inter0), .b(s_26), .O(gate14inter1));
  and2  gate731(.a(G12), .b(G11), .O(gate14inter2));
  inv1  gate732(.a(s_26), .O(gate14inter3));
  inv1  gate733(.a(s_27), .O(gate14inter4));
  nand2 gate734(.a(gate14inter4), .b(gate14inter3), .O(gate14inter5));
  nor2  gate735(.a(gate14inter5), .b(gate14inter2), .O(gate14inter6));
  inv1  gate736(.a(G11), .O(gate14inter7));
  inv1  gate737(.a(G12), .O(gate14inter8));
  nand2 gate738(.a(gate14inter8), .b(gate14inter7), .O(gate14inter9));
  nand2 gate739(.a(s_27), .b(gate14inter3), .O(gate14inter10));
  nor2  gate740(.a(gate14inter10), .b(gate14inter9), .O(gate14inter11));
  nor2  gate741(.a(gate14inter11), .b(gate14inter6), .O(gate14inter12));
  nand2 gate742(.a(gate14inter12), .b(gate14inter1), .O(G281));
nand2 gate15( .a(G13), .b(G14), .O(G284) );
nand2 gate16( .a(G15), .b(G16), .O(G287) );

  xor2  gate1583(.a(G18), .b(G17), .O(gate17inter0));
  nand2 gate1584(.a(gate17inter0), .b(s_148), .O(gate17inter1));
  and2  gate1585(.a(G18), .b(G17), .O(gate17inter2));
  inv1  gate1586(.a(s_148), .O(gate17inter3));
  inv1  gate1587(.a(s_149), .O(gate17inter4));
  nand2 gate1588(.a(gate17inter4), .b(gate17inter3), .O(gate17inter5));
  nor2  gate1589(.a(gate17inter5), .b(gate17inter2), .O(gate17inter6));
  inv1  gate1590(.a(G17), .O(gate17inter7));
  inv1  gate1591(.a(G18), .O(gate17inter8));
  nand2 gate1592(.a(gate17inter8), .b(gate17inter7), .O(gate17inter9));
  nand2 gate1593(.a(s_149), .b(gate17inter3), .O(gate17inter10));
  nor2  gate1594(.a(gate17inter10), .b(gate17inter9), .O(gate17inter11));
  nor2  gate1595(.a(gate17inter11), .b(gate17inter6), .O(gate17inter12));
  nand2 gate1596(.a(gate17inter12), .b(gate17inter1), .O(G290));

  xor2  gate701(.a(G20), .b(G19), .O(gate18inter0));
  nand2 gate702(.a(gate18inter0), .b(s_22), .O(gate18inter1));
  and2  gate703(.a(G20), .b(G19), .O(gate18inter2));
  inv1  gate704(.a(s_22), .O(gate18inter3));
  inv1  gate705(.a(s_23), .O(gate18inter4));
  nand2 gate706(.a(gate18inter4), .b(gate18inter3), .O(gate18inter5));
  nor2  gate707(.a(gate18inter5), .b(gate18inter2), .O(gate18inter6));
  inv1  gate708(.a(G19), .O(gate18inter7));
  inv1  gate709(.a(G20), .O(gate18inter8));
  nand2 gate710(.a(gate18inter8), .b(gate18inter7), .O(gate18inter9));
  nand2 gate711(.a(s_23), .b(gate18inter3), .O(gate18inter10));
  nor2  gate712(.a(gate18inter10), .b(gate18inter9), .O(gate18inter11));
  nor2  gate713(.a(gate18inter11), .b(gate18inter6), .O(gate18inter12));
  nand2 gate714(.a(gate18inter12), .b(gate18inter1), .O(G293));
nand2 gate19( .a(G21), .b(G22), .O(G296) );
nand2 gate20( .a(G23), .b(G24), .O(G299) );
nand2 gate21( .a(G25), .b(G26), .O(G302) );
nand2 gate22( .a(G27), .b(G28), .O(G305) );

  xor2  gate995(.a(G30), .b(G29), .O(gate23inter0));
  nand2 gate996(.a(gate23inter0), .b(s_64), .O(gate23inter1));
  and2  gate997(.a(G30), .b(G29), .O(gate23inter2));
  inv1  gate998(.a(s_64), .O(gate23inter3));
  inv1  gate999(.a(s_65), .O(gate23inter4));
  nand2 gate1000(.a(gate23inter4), .b(gate23inter3), .O(gate23inter5));
  nor2  gate1001(.a(gate23inter5), .b(gate23inter2), .O(gate23inter6));
  inv1  gate1002(.a(G29), .O(gate23inter7));
  inv1  gate1003(.a(G30), .O(gate23inter8));
  nand2 gate1004(.a(gate23inter8), .b(gate23inter7), .O(gate23inter9));
  nand2 gate1005(.a(s_65), .b(gate23inter3), .O(gate23inter10));
  nor2  gate1006(.a(gate23inter10), .b(gate23inter9), .O(gate23inter11));
  nor2  gate1007(.a(gate23inter11), .b(gate23inter6), .O(gate23inter12));
  nand2 gate1008(.a(gate23inter12), .b(gate23inter1), .O(G308));
nand2 gate24( .a(G31), .b(G32), .O(G311) );
nand2 gate25( .a(G1), .b(G5), .O(G314) );
nand2 gate26( .a(G9), .b(G13), .O(G317) );

  xor2  gate1219(.a(G6), .b(G2), .O(gate27inter0));
  nand2 gate1220(.a(gate27inter0), .b(s_96), .O(gate27inter1));
  and2  gate1221(.a(G6), .b(G2), .O(gate27inter2));
  inv1  gate1222(.a(s_96), .O(gate27inter3));
  inv1  gate1223(.a(s_97), .O(gate27inter4));
  nand2 gate1224(.a(gate27inter4), .b(gate27inter3), .O(gate27inter5));
  nor2  gate1225(.a(gate27inter5), .b(gate27inter2), .O(gate27inter6));
  inv1  gate1226(.a(G2), .O(gate27inter7));
  inv1  gate1227(.a(G6), .O(gate27inter8));
  nand2 gate1228(.a(gate27inter8), .b(gate27inter7), .O(gate27inter9));
  nand2 gate1229(.a(s_97), .b(gate27inter3), .O(gate27inter10));
  nor2  gate1230(.a(gate27inter10), .b(gate27inter9), .O(gate27inter11));
  nor2  gate1231(.a(gate27inter11), .b(gate27inter6), .O(gate27inter12));
  nand2 gate1232(.a(gate27inter12), .b(gate27inter1), .O(G320));

  xor2  gate1051(.a(G14), .b(G10), .O(gate28inter0));
  nand2 gate1052(.a(gate28inter0), .b(s_72), .O(gate28inter1));
  and2  gate1053(.a(G14), .b(G10), .O(gate28inter2));
  inv1  gate1054(.a(s_72), .O(gate28inter3));
  inv1  gate1055(.a(s_73), .O(gate28inter4));
  nand2 gate1056(.a(gate28inter4), .b(gate28inter3), .O(gate28inter5));
  nor2  gate1057(.a(gate28inter5), .b(gate28inter2), .O(gate28inter6));
  inv1  gate1058(.a(G10), .O(gate28inter7));
  inv1  gate1059(.a(G14), .O(gate28inter8));
  nand2 gate1060(.a(gate28inter8), .b(gate28inter7), .O(gate28inter9));
  nand2 gate1061(.a(s_73), .b(gate28inter3), .O(gate28inter10));
  nor2  gate1062(.a(gate28inter10), .b(gate28inter9), .O(gate28inter11));
  nor2  gate1063(.a(gate28inter11), .b(gate28inter6), .O(gate28inter12));
  nand2 gate1064(.a(gate28inter12), .b(gate28inter1), .O(G323));

  xor2  gate813(.a(G7), .b(G3), .O(gate29inter0));
  nand2 gate814(.a(gate29inter0), .b(s_38), .O(gate29inter1));
  and2  gate815(.a(G7), .b(G3), .O(gate29inter2));
  inv1  gate816(.a(s_38), .O(gate29inter3));
  inv1  gate817(.a(s_39), .O(gate29inter4));
  nand2 gate818(.a(gate29inter4), .b(gate29inter3), .O(gate29inter5));
  nor2  gate819(.a(gate29inter5), .b(gate29inter2), .O(gate29inter6));
  inv1  gate820(.a(G3), .O(gate29inter7));
  inv1  gate821(.a(G7), .O(gate29inter8));
  nand2 gate822(.a(gate29inter8), .b(gate29inter7), .O(gate29inter9));
  nand2 gate823(.a(s_39), .b(gate29inter3), .O(gate29inter10));
  nor2  gate824(.a(gate29inter10), .b(gate29inter9), .O(gate29inter11));
  nor2  gate825(.a(gate29inter11), .b(gate29inter6), .O(gate29inter12));
  nand2 gate826(.a(gate29inter12), .b(gate29inter1), .O(G326));
nand2 gate30( .a(G11), .b(G15), .O(G329) );
nand2 gate31( .a(G4), .b(G8), .O(G332) );
nand2 gate32( .a(G12), .b(G16), .O(G335) );
nand2 gate33( .a(G17), .b(G21), .O(G338) );
nand2 gate34( .a(G25), .b(G29), .O(G341) );
nand2 gate35( .a(G18), .b(G22), .O(G344) );
nand2 gate36( .a(G26), .b(G30), .O(G347) );
nand2 gate37( .a(G19), .b(G23), .O(G350) );
nand2 gate38( .a(G27), .b(G31), .O(G353) );

  xor2  gate2059(.a(G24), .b(G20), .O(gate39inter0));
  nand2 gate2060(.a(gate39inter0), .b(s_216), .O(gate39inter1));
  and2  gate2061(.a(G24), .b(G20), .O(gate39inter2));
  inv1  gate2062(.a(s_216), .O(gate39inter3));
  inv1  gate2063(.a(s_217), .O(gate39inter4));
  nand2 gate2064(.a(gate39inter4), .b(gate39inter3), .O(gate39inter5));
  nor2  gate2065(.a(gate39inter5), .b(gate39inter2), .O(gate39inter6));
  inv1  gate2066(.a(G20), .O(gate39inter7));
  inv1  gate2067(.a(G24), .O(gate39inter8));
  nand2 gate2068(.a(gate39inter8), .b(gate39inter7), .O(gate39inter9));
  nand2 gate2069(.a(s_217), .b(gate39inter3), .O(gate39inter10));
  nor2  gate2070(.a(gate39inter10), .b(gate39inter9), .O(gate39inter11));
  nor2  gate2071(.a(gate39inter11), .b(gate39inter6), .O(gate39inter12));
  nand2 gate2072(.a(gate39inter12), .b(gate39inter1), .O(G356));
nand2 gate40( .a(G28), .b(G32), .O(G359) );
nand2 gate41( .a(G1), .b(G266), .O(G362) );
nand2 gate42( .a(G2), .b(G266), .O(G363) );
nand2 gate43( .a(G3), .b(G269), .O(G364) );

  xor2  gate1135(.a(G269), .b(G4), .O(gate44inter0));
  nand2 gate1136(.a(gate44inter0), .b(s_84), .O(gate44inter1));
  and2  gate1137(.a(G269), .b(G4), .O(gate44inter2));
  inv1  gate1138(.a(s_84), .O(gate44inter3));
  inv1  gate1139(.a(s_85), .O(gate44inter4));
  nand2 gate1140(.a(gate44inter4), .b(gate44inter3), .O(gate44inter5));
  nor2  gate1141(.a(gate44inter5), .b(gate44inter2), .O(gate44inter6));
  inv1  gate1142(.a(G4), .O(gate44inter7));
  inv1  gate1143(.a(G269), .O(gate44inter8));
  nand2 gate1144(.a(gate44inter8), .b(gate44inter7), .O(gate44inter9));
  nand2 gate1145(.a(s_85), .b(gate44inter3), .O(gate44inter10));
  nor2  gate1146(.a(gate44inter10), .b(gate44inter9), .O(gate44inter11));
  nor2  gate1147(.a(gate44inter11), .b(gate44inter6), .O(gate44inter12));
  nand2 gate1148(.a(gate44inter12), .b(gate44inter1), .O(G365));

  xor2  gate1429(.a(G272), .b(G5), .O(gate45inter0));
  nand2 gate1430(.a(gate45inter0), .b(s_126), .O(gate45inter1));
  and2  gate1431(.a(G272), .b(G5), .O(gate45inter2));
  inv1  gate1432(.a(s_126), .O(gate45inter3));
  inv1  gate1433(.a(s_127), .O(gate45inter4));
  nand2 gate1434(.a(gate45inter4), .b(gate45inter3), .O(gate45inter5));
  nor2  gate1435(.a(gate45inter5), .b(gate45inter2), .O(gate45inter6));
  inv1  gate1436(.a(G5), .O(gate45inter7));
  inv1  gate1437(.a(G272), .O(gate45inter8));
  nand2 gate1438(.a(gate45inter8), .b(gate45inter7), .O(gate45inter9));
  nand2 gate1439(.a(s_127), .b(gate45inter3), .O(gate45inter10));
  nor2  gate1440(.a(gate45inter10), .b(gate45inter9), .O(gate45inter11));
  nor2  gate1441(.a(gate45inter11), .b(gate45inter6), .O(gate45inter12));
  nand2 gate1442(.a(gate45inter12), .b(gate45inter1), .O(G366));
nand2 gate46( .a(G6), .b(G272), .O(G367) );
nand2 gate47( .a(G7), .b(G275), .O(G368) );
nand2 gate48( .a(G8), .b(G275), .O(G369) );
nand2 gate49( .a(G9), .b(G278), .O(G370) );
nand2 gate50( .a(G10), .b(G278), .O(G371) );
nand2 gate51( .a(G11), .b(G281), .O(G372) );
nand2 gate52( .a(G12), .b(G281), .O(G373) );

  xor2  gate2101(.a(G284), .b(G13), .O(gate53inter0));
  nand2 gate2102(.a(gate53inter0), .b(s_222), .O(gate53inter1));
  and2  gate2103(.a(G284), .b(G13), .O(gate53inter2));
  inv1  gate2104(.a(s_222), .O(gate53inter3));
  inv1  gate2105(.a(s_223), .O(gate53inter4));
  nand2 gate2106(.a(gate53inter4), .b(gate53inter3), .O(gate53inter5));
  nor2  gate2107(.a(gate53inter5), .b(gate53inter2), .O(gate53inter6));
  inv1  gate2108(.a(G13), .O(gate53inter7));
  inv1  gate2109(.a(G284), .O(gate53inter8));
  nand2 gate2110(.a(gate53inter8), .b(gate53inter7), .O(gate53inter9));
  nand2 gate2111(.a(s_223), .b(gate53inter3), .O(gate53inter10));
  nor2  gate2112(.a(gate53inter10), .b(gate53inter9), .O(gate53inter11));
  nor2  gate2113(.a(gate53inter11), .b(gate53inter6), .O(gate53inter12));
  nand2 gate2114(.a(gate53inter12), .b(gate53inter1), .O(G374));
nand2 gate54( .a(G14), .b(G284), .O(G375) );
nand2 gate55( .a(G15), .b(G287), .O(G376) );
nand2 gate56( .a(G16), .b(G287), .O(G377) );
nand2 gate57( .a(G17), .b(G290), .O(G378) );
nand2 gate58( .a(G18), .b(G290), .O(G379) );
nand2 gate59( .a(G19), .b(G293), .O(G380) );
nand2 gate60( .a(G20), .b(G293), .O(G381) );
nand2 gate61( .a(G21), .b(G296), .O(G382) );
nand2 gate62( .a(G22), .b(G296), .O(G383) );
nand2 gate63( .a(G23), .b(G299), .O(G384) );
nand2 gate64( .a(G24), .b(G299), .O(G385) );
nand2 gate65( .a(G25), .b(G302), .O(G386) );
nand2 gate66( .a(G26), .b(G302), .O(G387) );

  xor2  gate1359(.a(G305), .b(G27), .O(gate67inter0));
  nand2 gate1360(.a(gate67inter0), .b(s_116), .O(gate67inter1));
  and2  gate1361(.a(G305), .b(G27), .O(gate67inter2));
  inv1  gate1362(.a(s_116), .O(gate67inter3));
  inv1  gate1363(.a(s_117), .O(gate67inter4));
  nand2 gate1364(.a(gate67inter4), .b(gate67inter3), .O(gate67inter5));
  nor2  gate1365(.a(gate67inter5), .b(gate67inter2), .O(gate67inter6));
  inv1  gate1366(.a(G27), .O(gate67inter7));
  inv1  gate1367(.a(G305), .O(gate67inter8));
  nand2 gate1368(.a(gate67inter8), .b(gate67inter7), .O(gate67inter9));
  nand2 gate1369(.a(s_117), .b(gate67inter3), .O(gate67inter10));
  nor2  gate1370(.a(gate67inter10), .b(gate67inter9), .O(gate67inter11));
  nor2  gate1371(.a(gate67inter11), .b(gate67inter6), .O(gate67inter12));
  nand2 gate1372(.a(gate67inter12), .b(gate67inter1), .O(G388));
nand2 gate68( .a(G28), .b(G305), .O(G389) );
nand2 gate69( .a(G29), .b(G308), .O(G390) );
nand2 gate70( .a(G30), .b(G308), .O(G391) );
nand2 gate71( .a(G31), .b(G311), .O(G392) );

  xor2  gate1947(.a(G311), .b(G32), .O(gate72inter0));
  nand2 gate1948(.a(gate72inter0), .b(s_200), .O(gate72inter1));
  and2  gate1949(.a(G311), .b(G32), .O(gate72inter2));
  inv1  gate1950(.a(s_200), .O(gate72inter3));
  inv1  gate1951(.a(s_201), .O(gate72inter4));
  nand2 gate1952(.a(gate72inter4), .b(gate72inter3), .O(gate72inter5));
  nor2  gate1953(.a(gate72inter5), .b(gate72inter2), .O(gate72inter6));
  inv1  gate1954(.a(G32), .O(gate72inter7));
  inv1  gate1955(.a(G311), .O(gate72inter8));
  nand2 gate1956(.a(gate72inter8), .b(gate72inter7), .O(gate72inter9));
  nand2 gate1957(.a(s_201), .b(gate72inter3), .O(gate72inter10));
  nor2  gate1958(.a(gate72inter10), .b(gate72inter9), .O(gate72inter11));
  nor2  gate1959(.a(gate72inter11), .b(gate72inter6), .O(gate72inter12));
  nand2 gate1960(.a(gate72inter12), .b(gate72inter1), .O(G393));
nand2 gate73( .a(G1), .b(G314), .O(G394) );
nand2 gate74( .a(G5), .b(G314), .O(G395) );
nand2 gate75( .a(G9), .b(G317), .O(G396) );
nand2 gate76( .a(G13), .b(G317), .O(G397) );

  xor2  gate1989(.a(G320), .b(G2), .O(gate77inter0));
  nand2 gate1990(.a(gate77inter0), .b(s_206), .O(gate77inter1));
  and2  gate1991(.a(G320), .b(G2), .O(gate77inter2));
  inv1  gate1992(.a(s_206), .O(gate77inter3));
  inv1  gate1993(.a(s_207), .O(gate77inter4));
  nand2 gate1994(.a(gate77inter4), .b(gate77inter3), .O(gate77inter5));
  nor2  gate1995(.a(gate77inter5), .b(gate77inter2), .O(gate77inter6));
  inv1  gate1996(.a(G2), .O(gate77inter7));
  inv1  gate1997(.a(G320), .O(gate77inter8));
  nand2 gate1998(.a(gate77inter8), .b(gate77inter7), .O(gate77inter9));
  nand2 gate1999(.a(s_207), .b(gate77inter3), .O(gate77inter10));
  nor2  gate2000(.a(gate77inter10), .b(gate77inter9), .O(gate77inter11));
  nor2  gate2001(.a(gate77inter11), .b(gate77inter6), .O(gate77inter12));
  nand2 gate2002(.a(gate77inter12), .b(gate77inter1), .O(G398));
nand2 gate78( .a(G6), .b(G320), .O(G399) );

  xor2  gate1331(.a(G323), .b(G10), .O(gate79inter0));
  nand2 gate1332(.a(gate79inter0), .b(s_112), .O(gate79inter1));
  and2  gate1333(.a(G323), .b(G10), .O(gate79inter2));
  inv1  gate1334(.a(s_112), .O(gate79inter3));
  inv1  gate1335(.a(s_113), .O(gate79inter4));
  nand2 gate1336(.a(gate79inter4), .b(gate79inter3), .O(gate79inter5));
  nor2  gate1337(.a(gate79inter5), .b(gate79inter2), .O(gate79inter6));
  inv1  gate1338(.a(G10), .O(gate79inter7));
  inv1  gate1339(.a(G323), .O(gate79inter8));
  nand2 gate1340(.a(gate79inter8), .b(gate79inter7), .O(gate79inter9));
  nand2 gate1341(.a(s_113), .b(gate79inter3), .O(gate79inter10));
  nor2  gate1342(.a(gate79inter10), .b(gate79inter9), .O(gate79inter11));
  nor2  gate1343(.a(gate79inter11), .b(gate79inter6), .O(gate79inter12));
  nand2 gate1344(.a(gate79inter12), .b(gate79inter1), .O(G400));
nand2 gate80( .a(G14), .b(G323), .O(G401) );
nand2 gate81( .a(G3), .b(G326), .O(G402) );

  xor2  gate743(.a(G326), .b(G7), .O(gate82inter0));
  nand2 gate744(.a(gate82inter0), .b(s_28), .O(gate82inter1));
  and2  gate745(.a(G326), .b(G7), .O(gate82inter2));
  inv1  gate746(.a(s_28), .O(gate82inter3));
  inv1  gate747(.a(s_29), .O(gate82inter4));
  nand2 gate748(.a(gate82inter4), .b(gate82inter3), .O(gate82inter5));
  nor2  gate749(.a(gate82inter5), .b(gate82inter2), .O(gate82inter6));
  inv1  gate750(.a(G7), .O(gate82inter7));
  inv1  gate751(.a(G326), .O(gate82inter8));
  nand2 gate752(.a(gate82inter8), .b(gate82inter7), .O(gate82inter9));
  nand2 gate753(.a(s_29), .b(gate82inter3), .O(gate82inter10));
  nor2  gate754(.a(gate82inter10), .b(gate82inter9), .O(gate82inter11));
  nor2  gate755(.a(gate82inter11), .b(gate82inter6), .O(gate82inter12));
  nand2 gate756(.a(gate82inter12), .b(gate82inter1), .O(G403));
nand2 gate83( .a(G11), .b(G329), .O(G404) );
nand2 gate84( .a(G15), .b(G329), .O(G405) );
nand2 gate85( .a(G4), .b(G332), .O(G406) );
nand2 gate86( .a(G8), .b(G332), .O(G407) );

  xor2  gate841(.a(G335), .b(G12), .O(gate87inter0));
  nand2 gate842(.a(gate87inter0), .b(s_42), .O(gate87inter1));
  and2  gate843(.a(G335), .b(G12), .O(gate87inter2));
  inv1  gate844(.a(s_42), .O(gate87inter3));
  inv1  gate845(.a(s_43), .O(gate87inter4));
  nand2 gate846(.a(gate87inter4), .b(gate87inter3), .O(gate87inter5));
  nor2  gate847(.a(gate87inter5), .b(gate87inter2), .O(gate87inter6));
  inv1  gate848(.a(G12), .O(gate87inter7));
  inv1  gate849(.a(G335), .O(gate87inter8));
  nand2 gate850(.a(gate87inter8), .b(gate87inter7), .O(gate87inter9));
  nand2 gate851(.a(s_43), .b(gate87inter3), .O(gate87inter10));
  nor2  gate852(.a(gate87inter10), .b(gate87inter9), .O(gate87inter11));
  nor2  gate853(.a(gate87inter11), .b(gate87inter6), .O(gate87inter12));
  nand2 gate854(.a(gate87inter12), .b(gate87inter1), .O(G408));
nand2 gate88( .a(G16), .b(G335), .O(G409) );

  xor2  gate1317(.a(G338), .b(G17), .O(gate89inter0));
  nand2 gate1318(.a(gate89inter0), .b(s_110), .O(gate89inter1));
  and2  gate1319(.a(G338), .b(G17), .O(gate89inter2));
  inv1  gate1320(.a(s_110), .O(gate89inter3));
  inv1  gate1321(.a(s_111), .O(gate89inter4));
  nand2 gate1322(.a(gate89inter4), .b(gate89inter3), .O(gate89inter5));
  nor2  gate1323(.a(gate89inter5), .b(gate89inter2), .O(gate89inter6));
  inv1  gate1324(.a(G17), .O(gate89inter7));
  inv1  gate1325(.a(G338), .O(gate89inter8));
  nand2 gate1326(.a(gate89inter8), .b(gate89inter7), .O(gate89inter9));
  nand2 gate1327(.a(s_111), .b(gate89inter3), .O(gate89inter10));
  nor2  gate1328(.a(gate89inter10), .b(gate89inter9), .O(gate89inter11));
  nor2  gate1329(.a(gate89inter11), .b(gate89inter6), .O(gate89inter12));
  nand2 gate1330(.a(gate89inter12), .b(gate89inter1), .O(G410));

  xor2  gate1065(.a(G338), .b(G21), .O(gate90inter0));
  nand2 gate1066(.a(gate90inter0), .b(s_74), .O(gate90inter1));
  and2  gate1067(.a(G338), .b(G21), .O(gate90inter2));
  inv1  gate1068(.a(s_74), .O(gate90inter3));
  inv1  gate1069(.a(s_75), .O(gate90inter4));
  nand2 gate1070(.a(gate90inter4), .b(gate90inter3), .O(gate90inter5));
  nor2  gate1071(.a(gate90inter5), .b(gate90inter2), .O(gate90inter6));
  inv1  gate1072(.a(G21), .O(gate90inter7));
  inv1  gate1073(.a(G338), .O(gate90inter8));
  nand2 gate1074(.a(gate90inter8), .b(gate90inter7), .O(gate90inter9));
  nand2 gate1075(.a(s_75), .b(gate90inter3), .O(gate90inter10));
  nor2  gate1076(.a(gate90inter10), .b(gate90inter9), .O(gate90inter11));
  nor2  gate1077(.a(gate90inter11), .b(gate90inter6), .O(gate90inter12));
  nand2 gate1078(.a(gate90inter12), .b(gate90inter1), .O(G411));
nand2 gate91( .a(G25), .b(G341), .O(G412) );

  xor2  gate1191(.a(G341), .b(G29), .O(gate92inter0));
  nand2 gate1192(.a(gate92inter0), .b(s_92), .O(gate92inter1));
  and2  gate1193(.a(G341), .b(G29), .O(gate92inter2));
  inv1  gate1194(.a(s_92), .O(gate92inter3));
  inv1  gate1195(.a(s_93), .O(gate92inter4));
  nand2 gate1196(.a(gate92inter4), .b(gate92inter3), .O(gate92inter5));
  nor2  gate1197(.a(gate92inter5), .b(gate92inter2), .O(gate92inter6));
  inv1  gate1198(.a(G29), .O(gate92inter7));
  inv1  gate1199(.a(G341), .O(gate92inter8));
  nand2 gate1200(.a(gate92inter8), .b(gate92inter7), .O(gate92inter9));
  nand2 gate1201(.a(s_93), .b(gate92inter3), .O(gate92inter10));
  nor2  gate1202(.a(gate92inter10), .b(gate92inter9), .O(gate92inter11));
  nor2  gate1203(.a(gate92inter11), .b(gate92inter6), .O(gate92inter12));
  nand2 gate1204(.a(gate92inter12), .b(gate92inter1), .O(G413));
nand2 gate93( .a(G18), .b(G344), .O(G414) );
nand2 gate94( .a(G22), .b(G344), .O(G415) );
nand2 gate95( .a(G26), .b(G347), .O(G416) );
nand2 gate96( .a(G30), .b(G347), .O(G417) );
nand2 gate97( .a(G19), .b(G350), .O(G418) );

  xor2  gate1009(.a(G350), .b(G23), .O(gate98inter0));
  nand2 gate1010(.a(gate98inter0), .b(s_66), .O(gate98inter1));
  and2  gate1011(.a(G350), .b(G23), .O(gate98inter2));
  inv1  gate1012(.a(s_66), .O(gate98inter3));
  inv1  gate1013(.a(s_67), .O(gate98inter4));
  nand2 gate1014(.a(gate98inter4), .b(gate98inter3), .O(gate98inter5));
  nor2  gate1015(.a(gate98inter5), .b(gate98inter2), .O(gate98inter6));
  inv1  gate1016(.a(G23), .O(gate98inter7));
  inv1  gate1017(.a(G350), .O(gate98inter8));
  nand2 gate1018(.a(gate98inter8), .b(gate98inter7), .O(gate98inter9));
  nand2 gate1019(.a(s_67), .b(gate98inter3), .O(gate98inter10));
  nor2  gate1020(.a(gate98inter10), .b(gate98inter9), .O(gate98inter11));
  nor2  gate1021(.a(gate98inter11), .b(gate98inter6), .O(gate98inter12));
  nand2 gate1022(.a(gate98inter12), .b(gate98inter1), .O(G419));
nand2 gate99( .a(G27), .b(G353), .O(G420) );
nand2 gate100( .a(G31), .b(G353), .O(G421) );
nand2 gate101( .a(G20), .b(G356), .O(G422) );
nand2 gate102( .a(G24), .b(G356), .O(G423) );
nand2 gate103( .a(G28), .b(G359), .O(G424) );

  xor2  gate911(.a(G359), .b(G32), .O(gate104inter0));
  nand2 gate912(.a(gate104inter0), .b(s_52), .O(gate104inter1));
  and2  gate913(.a(G359), .b(G32), .O(gate104inter2));
  inv1  gate914(.a(s_52), .O(gate104inter3));
  inv1  gate915(.a(s_53), .O(gate104inter4));
  nand2 gate916(.a(gate104inter4), .b(gate104inter3), .O(gate104inter5));
  nor2  gate917(.a(gate104inter5), .b(gate104inter2), .O(gate104inter6));
  inv1  gate918(.a(G32), .O(gate104inter7));
  inv1  gate919(.a(G359), .O(gate104inter8));
  nand2 gate920(.a(gate104inter8), .b(gate104inter7), .O(gate104inter9));
  nand2 gate921(.a(s_53), .b(gate104inter3), .O(gate104inter10));
  nor2  gate922(.a(gate104inter10), .b(gate104inter9), .O(gate104inter11));
  nor2  gate923(.a(gate104inter11), .b(gate104inter6), .O(gate104inter12));
  nand2 gate924(.a(gate104inter12), .b(gate104inter1), .O(G425));

  xor2  gate1527(.a(G363), .b(G362), .O(gate105inter0));
  nand2 gate1528(.a(gate105inter0), .b(s_140), .O(gate105inter1));
  and2  gate1529(.a(G363), .b(G362), .O(gate105inter2));
  inv1  gate1530(.a(s_140), .O(gate105inter3));
  inv1  gate1531(.a(s_141), .O(gate105inter4));
  nand2 gate1532(.a(gate105inter4), .b(gate105inter3), .O(gate105inter5));
  nor2  gate1533(.a(gate105inter5), .b(gate105inter2), .O(gate105inter6));
  inv1  gate1534(.a(G362), .O(gate105inter7));
  inv1  gate1535(.a(G363), .O(gate105inter8));
  nand2 gate1536(.a(gate105inter8), .b(gate105inter7), .O(gate105inter9));
  nand2 gate1537(.a(s_141), .b(gate105inter3), .O(gate105inter10));
  nor2  gate1538(.a(gate105inter10), .b(gate105inter9), .O(gate105inter11));
  nor2  gate1539(.a(gate105inter11), .b(gate105inter6), .O(gate105inter12));
  nand2 gate1540(.a(gate105inter12), .b(gate105inter1), .O(G426));
nand2 gate106( .a(G364), .b(G365), .O(G429) );
nand2 gate107( .a(G366), .b(G367), .O(G432) );

  xor2  gate1555(.a(G369), .b(G368), .O(gate108inter0));
  nand2 gate1556(.a(gate108inter0), .b(s_144), .O(gate108inter1));
  and2  gate1557(.a(G369), .b(G368), .O(gate108inter2));
  inv1  gate1558(.a(s_144), .O(gate108inter3));
  inv1  gate1559(.a(s_145), .O(gate108inter4));
  nand2 gate1560(.a(gate108inter4), .b(gate108inter3), .O(gate108inter5));
  nor2  gate1561(.a(gate108inter5), .b(gate108inter2), .O(gate108inter6));
  inv1  gate1562(.a(G368), .O(gate108inter7));
  inv1  gate1563(.a(G369), .O(gate108inter8));
  nand2 gate1564(.a(gate108inter8), .b(gate108inter7), .O(gate108inter9));
  nand2 gate1565(.a(s_145), .b(gate108inter3), .O(gate108inter10));
  nor2  gate1566(.a(gate108inter10), .b(gate108inter9), .O(gate108inter11));
  nor2  gate1567(.a(gate108inter11), .b(gate108inter6), .O(gate108inter12));
  nand2 gate1568(.a(gate108inter12), .b(gate108inter1), .O(G435));
nand2 gate109( .a(G370), .b(G371), .O(G438) );

  xor2  gate575(.a(G373), .b(G372), .O(gate110inter0));
  nand2 gate576(.a(gate110inter0), .b(s_4), .O(gate110inter1));
  and2  gate577(.a(G373), .b(G372), .O(gate110inter2));
  inv1  gate578(.a(s_4), .O(gate110inter3));
  inv1  gate579(.a(s_5), .O(gate110inter4));
  nand2 gate580(.a(gate110inter4), .b(gate110inter3), .O(gate110inter5));
  nor2  gate581(.a(gate110inter5), .b(gate110inter2), .O(gate110inter6));
  inv1  gate582(.a(G372), .O(gate110inter7));
  inv1  gate583(.a(G373), .O(gate110inter8));
  nand2 gate584(.a(gate110inter8), .b(gate110inter7), .O(gate110inter9));
  nand2 gate585(.a(s_5), .b(gate110inter3), .O(gate110inter10));
  nor2  gate586(.a(gate110inter10), .b(gate110inter9), .O(gate110inter11));
  nor2  gate587(.a(gate110inter11), .b(gate110inter6), .O(gate110inter12));
  nand2 gate588(.a(gate110inter12), .b(gate110inter1), .O(G441));
nand2 gate111( .a(G374), .b(G375), .O(G444) );

  xor2  gate617(.a(G377), .b(G376), .O(gate112inter0));
  nand2 gate618(.a(gate112inter0), .b(s_10), .O(gate112inter1));
  and2  gate619(.a(G377), .b(G376), .O(gate112inter2));
  inv1  gate620(.a(s_10), .O(gate112inter3));
  inv1  gate621(.a(s_11), .O(gate112inter4));
  nand2 gate622(.a(gate112inter4), .b(gate112inter3), .O(gate112inter5));
  nor2  gate623(.a(gate112inter5), .b(gate112inter2), .O(gate112inter6));
  inv1  gate624(.a(G376), .O(gate112inter7));
  inv1  gate625(.a(G377), .O(gate112inter8));
  nand2 gate626(.a(gate112inter8), .b(gate112inter7), .O(gate112inter9));
  nand2 gate627(.a(s_11), .b(gate112inter3), .O(gate112inter10));
  nor2  gate628(.a(gate112inter10), .b(gate112inter9), .O(gate112inter11));
  nor2  gate629(.a(gate112inter11), .b(gate112inter6), .O(gate112inter12));
  nand2 gate630(.a(gate112inter12), .b(gate112inter1), .O(G447));
nand2 gate113( .a(G378), .b(G379), .O(G450) );

  xor2  gate687(.a(G381), .b(G380), .O(gate114inter0));
  nand2 gate688(.a(gate114inter0), .b(s_20), .O(gate114inter1));
  and2  gate689(.a(G381), .b(G380), .O(gate114inter2));
  inv1  gate690(.a(s_20), .O(gate114inter3));
  inv1  gate691(.a(s_21), .O(gate114inter4));
  nand2 gate692(.a(gate114inter4), .b(gate114inter3), .O(gate114inter5));
  nor2  gate693(.a(gate114inter5), .b(gate114inter2), .O(gate114inter6));
  inv1  gate694(.a(G380), .O(gate114inter7));
  inv1  gate695(.a(G381), .O(gate114inter8));
  nand2 gate696(.a(gate114inter8), .b(gate114inter7), .O(gate114inter9));
  nand2 gate697(.a(s_21), .b(gate114inter3), .O(gate114inter10));
  nor2  gate698(.a(gate114inter10), .b(gate114inter9), .O(gate114inter11));
  nor2  gate699(.a(gate114inter11), .b(gate114inter6), .O(gate114inter12));
  nand2 gate700(.a(gate114inter12), .b(gate114inter1), .O(G453));

  xor2  gate1163(.a(G383), .b(G382), .O(gate115inter0));
  nand2 gate1164(.a(gate115inter0), .b(s_88), .O(gate115inter1));
  and2  gate1165(.a(G383), .b(G382), .O(gate115inter2));
  inv1  gate1166(.a(s_88), .O(gate115inter3));
  inv1  gate1167(.a(s_89), .O(gate115inter4));
  nand2 gate1168(.a(gate115inter4), .b(gate115inter3), .O(gate115inter5));
  nor2  gate1169(.a(gate115inter5), .b(gate115inter2), .O(gate115inter6));
  inv1  gate1170(.a(G382), .O(gate115inter7));
  inv1  gate1171(.a(G383), .O(gate115inter8));
  nand2 gate1172(.a(gate115inter8), .b(gate115inter7), .O(gate115inter9));
  nand2 gate1173(.a(s_89), .b(gate115inter3), .O(gate115inter10));
  nor2  gate1174(.a(gate115inter10), .b(gate115inter9), .O(gate115inter11));
  nor2  gate1175(.a(gate115inter11), .b(gate115inter6), .O(gate115inter12));
  nand2 gate1176(.a(gate115inter12), .b(gate115inter1), .O(G456));

  xor2  gate1793(.a(G385), .b(G384), .O(gate116inter0));
  nand2 gate1794(.a(gate116inter0), .b(s_178), .O(gate116inter1));
  and2  gate1795(.a(G385), .b(G384), .O(gate116inter2));
  inv1  gate1796(.a(s_178), .O(gate116inter3));
  inv1  gate1797(.a(s_179), .O(gate116inter4));
  nand2 gate1798(.a(gate116inter4), .b(gate116inter3), .O(gate116inter5));
  nor2  gate1799(.a(gate116inter5), .b(gate116inter2), .O(gate116inter6));
  inv1  gate1800(.a(G384), .O(gate116inter7));
  inv1  gate1801(.a(G385), .O(gate116inter8));
  nand2 gate1802(.a(gate116inter8), .b(gate116inter7), .O(gate116inter9));
  nand2 gate1803(.a(s_179), .b(gate116inter3), .O(gate116inter10));
  nor2  gate1804(.a(gate116inter10), .b(gate116inter9), .O(gate116inter11));
  nor2  gate1805(.a(gate116inter11), .b(gate116inter6), .O(gate116inter12));
  nand2 gate1806(.a(gate116inter12), .b(gate116inter1), .O(G459));

  xor2  gate1709(.a(G387), .b(G386), .O(gate117inter0));
  nand2 gate1710(.a(gate117inter0), .b(s_166), .O(gate117inter1));
  and2  gate1711(.a(G387), .b(G386), .O(gate117inter2));
  inv1  gate1712(.a(s_166), .O(gate117inter3));
  inv1  gate1713(.a(s_167), .O(gate117inter4));
  nand2 gate1714(.a(gate117inter4), .b(gate117inter3), .O(gate117inter5));
  nor2  gate1715(.a(gate117inter5), .b(gate117inter2), .O(gate117inter6));
  inv1  gate1716(.a(G386), .O(gate117inter7));
  inv1  gate1717(.a(G387), .O(gate117inter8));
  nand2 gate1718(.a(gate117inter8), .b(gate117inter7), .O(gate117inter9));
  nand2 gate1719(.a(s_167), .b(gate117inter3), .O(gate117inter10));
  nor2  gate1720(.a(gate117inter10), .b(gate117inter9), .O(gate117inter11));
  nor2  gate1721(.a(gate117inter11), .b(gate117inter6), .O(gate117inter12));
  nand2 gate1722(.a(gate117inter12), .b(gate117inter1), .O(G462));
nand2 gate118( .a(G388), .b(G389), .O(G465) );
nand2 gate119( .a(G390), .b(G391), .O(G468) );
nand2 gate120( .a(G392), .b(G393), .O(G471) );

  xor2  gate1177(.a(G395), .b(G394), .O(gate121inter0));
  nand2 gate1178(.a(gate121inter0), .b(s_90), .O(gate121inter1));
  and2  gate1179(.a(G395), .b(G394), .O(gate121inter2));
  inv1  gate1180(.a(s_90), .O(gate121inter3));
  inv1  gate1181(.a(s_91), .O(gate121inter4));
  nand2 gate1182(.a(gate121inter4), .b(gate121inter3), .O(gate121inter5));
  nor2  gate1183(.a(gate121inter5), .b(gate121inter2), .O(gate121inter6));
  inv1  gate1184(.a(G394), .O(gate121inter7));
  inv1  gate1185(.a(G395), .O(gate121inter8));
  nand2 gate1186(.a(gate121inter8), .b(gate121inter7), .O(gate121inter9));
  nand2 gate1187(.a(s_91), .b(gate121inter3), .O(gate121inter10));
  nor2  gate1188(.a(gate121inter10), .b(gate121inter9), .O(gate121inter11));
  nor2  gate1189(.a(gate121inter11), .b(gate121inter6), .O(gate121inter12));
  nand2 gate1190(.a(gate121inter12), .b(gate121inter1), .O(G474));
nand2 gate122( .a(G396), .b(G397), .O(G477) );

  xor2  gate2115(.a(G399), .b(G398), .O(gate123inter0));
  nand2 gate2116(.a(gate123inter0), .b(s_224), .O(gate123inter1));
  and2  gate2117(.a(G399), .b(G398), .O(gate123inter2));
  inv1  gate2118(.a(s_224), .O(gate123inter3));
  inv1  gate2119(.a(s_225), .O(gate123inter4));
  nand2 gate2120(.a(gate123inter4), .b(gate123inter3), .O(gate123inter5));
  nor2  gate2121(.a(gate123inter5), .b(gate123inter2), .O(gate123inter6));
  inv1  gate2122(.a(G398), .O(gate123inter7));
  inv1  gate2123(.a(G399), .O(gate123inter8));
  nand2 gate2124(.a(gate123inter8), .b(gate123inter7), .O(gate123inter9));
  nand2 gate2125(.a(s_225), .b(gate123inter3), .O(gate123inter10));
  nor2  gate2126(.a(gate123inter10), .b(gate123inter9), .O(gate123inter11));
  nor2  gate2127(.a(gate123inter11), .b(gate123inter6), .O(gate123inter12));
  nand2 gate2128(.a(gate123inter12), .b(gate123inter1), .O(G480));
nand2 gate124( .a(G400), .b(G401), .O(G483) );

  xor2  gate757(.a(G403), .b(G402), .O(gate125inter0));
  nand2 gate758(.a(gate125inter0), .b(s_30), .O(gate125inter1));
  and2  gate759(.a(G403), .b(G402), .O(gate125inter2));
  inv1  gate760(.a(s_30), .O(gate125inter3));
  inv1  gate761(.a(s_31), .O(gate125inter4));
  nand2 gate762(.a(gate125inter4), .b(gate125inter3), .O(gate125inter5));
  nor2  gate763(.a(gate125inter5), .b(gate125inter2), .O(gate125inter6));
  inv1  gate764(.a(G402), .O(gate125inter7));
  inv1  gate765(.a(G403), .O(gate125inter8));
  nand2 gate766(.a(gate125inter8), .b(gate125inter7), .O(gate125inter9));
  nand2 gate767(.a(s_31), .b(gate125inter3), .O(gate125inter10));
  nor2  gate768(.a(gate125inter10), .b(gate125inter9), .O(gate125inter11));
  nor2  gate769(.a(gate125inter11), .b(gate125inter6), .O(gate125inter12));
  nand2 gate770(.a(gate125inter12), .b(gate125inter1), .O(G486));
nand2 gate126( .a(G404), .b(G405), .O(G489) );
nand2 gate127( .a(G406), .b(G407), .O(G492) );
nand2 gate128( .a(G408), .b(G409), .O(G495) );
nand2 gate129( .a(G410), .b(G411), .O(G498) );
nand2 gate130( .a(G412), .b(G413), .O(G501) );
nand2 gate131( .a(G414), .b(G415), .O(G504) );
nand2 gate132( .a(G416), .b(G417), .O(G507) );

  xor2  gate1443(.a(G419), .b(G418), .O(gate133inter0));
  nand2 gate1444(.a(gate133inter0), .b(s_128), .O(gate133inter1));
  and2  gate1445(.a(G419), .b(G418), .O(gate133inter2));
  inv1  gate1446(.a(s_128), .O(gate133inter3));
  inv1  gate1447(.a(s_129), .O(gate133inter4));
  nand2 gate1448(.a(gate133inter4), .b(gate133inter3), .O(gate133inter5));
  nor2  gate1449(.a(gate133inter5), .b(gate133inter2), .O(gate133inter6));
  inv1  gate1450(.a(G418), .O(gate133inter7));
  inv1  gate1451(.a(G419), .O(gate133inter8));
  nand2 gate1452(.a(gate133inter8), .b(gate133inter7), .O(gate133inter9));
  nand2 gate1453(.a(s_129), .b(gate133inter3), .O(gate133inter10));
  nor2  gate1454(.a(gate133inter10), .b(gate133inter9), .O(gate133inter11));
  nor2  gate1455(.a(gate133inter11), .b(gate133inter6), .O(gate133inter12));
  nand2 gate1456(.a(gate133inter12), .b(gate133inter1), .O(G510));

  xor2  gate645(.a(G421), .b(G420), .O(gate134inter0));
  nand2 gate646(.a(gate134inter0), .b(s_14), .O(gate134inter1));
  and2  gate647(.a(G421), .b(G420), .O(gate134inter2));
  inv1  gate648(.a(s_14), .O(gate134inter3));
  inv1  gate649(.a(s_15), .O(gate134inter4));
  nand2 gate650(.a(gate134inter4), .b(gate134inter3), .O(gate134inter5));
  nor2  gate651(.a(gate134inter5), .b(gate134inter2), .O(gate134inter6));
  inv1  gate652(.a(G420), .O(gate134inter7));
  inv1  gate653(.a(G421), .O(gate134inter8));
  nand2 gate654(.a(gate134inter8), .b(gate134inter7), .O(gate134inter9));
  nand2 gate655(.a(s_15), .b(gate134inter3), .O(gate134inter10));
  nor2  gate656(.a(gate134inter10), .b(gate134inter9), .O(gate134inter11));
  nor2  gate657(.a(gate134inter11), .b(gate134inter6), .O(gate134inter12));
  nand2 gate658(.a(gate134inter12), .b(gate134inter1), .O(G513));
nand2 gate135( .a(G422), .b(G423), .O(G516) );
nand2 gate136( .a(G424), .b(G425), .O(G519) );
nand2 gate137( .a(G426), .b(G429), .O(G522) );
nand2 gate138( .a(G432), .b(G435), .O(G525) );

  xor2  gate1891(.a(G441), .b(G438), .O(gate139inter0));
  nand2 gate1892(.a(gate139inter0), .b(s_192), .O(gate139inter1));
  and2  gate1893(.a(G441), .b(G438), .O(gate139inter2));
  inv1  gate1894(.a(s_192), .O(gate139inter3));
  inv1  gate1895(.a(s_193), .O(gate139inter4));
  nand2 gate1896(.a(gate139inter4), .b(gate139inter3), .O(gate139inter5));
  nor2  gate1897(.a(gate139inter5), .b(gate139inter2), .O(gate139inter6));
  inv1  gate1898(.a(G438), .O(gate139inter7));
  inv1  gate1899(.a(G441), .O(gate139inter8));
  nand2 gate1900(.a(gate139inter8), .b(gate139inter7), .O(gate139inter9));
  nand2 gate1901(.a(s_193), .b(gate139inter3), .O(gate139inter10));
  nor2  gate1902(.a(gate139inter10), .b(gate139inter9), .O(gate139inter11));
  nor2  gate1903(.a(gate139inter11), .b(gate139inter6), .O(gate139inter12));
  nand2 gate1904(.a(gate139inter12), .b(gate139inter1), .O(G528));
nand2 gate140( .a(G444), .b(G447), .O(G531) );
nand2 gate141( .a(G450), .b(G453), .O(G534) );

  xor2  gate2199(.a(G459), .b(G456), .O(gate142inter0));
  nand2 gate2200(.a(gate142inter0), .b(s_236), .O(gate142inter1));
  and2  gate2201(.a(G459), .b(G456), .O(gate142inter2));
  inv1  gate2202(.a(s_236), .O(gate142inter3));
  inv1  gate2203(.a(s_237), .O(gate142inter4));
  nand2 gate2204(.a(gate142inter4), .b(gate142inter3), .O(gate142inter5));
  nor2  gate2205(.a(gate142inter5), .b(gate142inter2), .O(gate142inter6));
  inv1  gate2206(.a(G456), .O(gate142inter7));
  inv1  gate2207(.a(G459), .O(gate142inter8));
  nand2 gate2208(.a(gate142inter8), .b(gate142inter7), .O(gate142inter9));
  nand2 gate2209(.a(s_237), .b(gate142inter3), .O(gate142inter10));
  nor2  gate2210(.a(gate142inter10), .b(gate142inter9), .O(gate142inter11));
  nor2  gate2211(.a(gate142inter11), .b(gate142inter6), .O(gate142inter12));
  nand2 gate2212(.a(gate142inter12), .b(gate142inter1), .O(G537));
nand2 gate143( .a(G462), .b(G465), .O(G540) );
nand2 gate144( .a(G468), .b(G471), .O(G543) );
nand2 gate145( .a(G474), .b(G477), .O(G546) );
nand2 gate146( .a(G480), .b(G483), .O(G549) );
nand2 gate147( .a(G486), .b(G489), .O(G552) );
nand2 gate148( .a(G492), .b(G495), .O(G555) );
nand2 gate149( .a(G498), .b(G501), .O(G558) );
nand2 gate150( .a(G504), .b(G507), .O(G561) );
nand2 gate151( .a(G510), .b(G513), .O(G564) );
nand2 gate152( .a(G516), .b(G519), .O(G567) );
nand2 gate153( .a(G426), .b(G522), .O(G570) );

  xor2  gate1023(.a(G522), .b(G429), .O(gate154inter0));
  nand2 gate1024(.a(gate154inter0), .b(s_68), .O(gate154inter1));
  and2  gate1025(.a(G522), .b(G429), .O(gate154inter2));
  inv1  gate1026(.a(s_68), .O(gate154inter3));
  inv1  gate1027(.a(s_69), .O(gate154inter4));
  nand2 gate1028(.a(gate154inter4), .b(gate154inter3), .O(gate154inter5));
  nor2  gate1029(.a(gate154inter5), .b(gate154inter2), .O(gate154inter6));
  inv1  gate1030(.a(G429), .O(gate154inter7));
  inv1  gate1031(.a(G522), .O(gate154inter8));
  nand2 gate1032(.a(gate154inter8), .b(gate154inter7), .O(gate154inter9));
  nand2 gate1033(.a(s_69), .b(gate154inter3), .O(gate154inter10));
  nor2  gate1034(.a(gate154inter10), .b(gate154inter9), .O(gate154inter11));
  nor2  gate1035(.a(gate154inter11), .b(gate154inter6), .O(gate154inter12));
  nand2 gate1036(.a(gate154inter12), .b(gate154inter1), .O(G571));
nand2 gate155( .a(G432), .b(G525), .O(G572) );
nand2 gate156( .a(G435), .b(G525), .O(G573) );
nand2 gate157( .a(G438), .b(G528), .O(G574) );
nand2 gate158( .a(G441), .b(G528), .O(G575) );

  xor2  gate1625(.a(G531), .b(G444), .O(gate159inter0));
  nand2 gate1626(.a(gate159inter0), .b(s_154), .O(gate159inter1));
  and2  gate1627(.a(G531), .b(G444), .O(gate159inter2));
  inv1  gate1628(.a(s_154), .O(gate159inter3));
  inv1  gate1629(.a(s_155), .O(gate159inter4));
  nand2 gate1630(.a(gate159inter4), .b(gate159inter3), .O(gate159inter5));
  nor2  gate1631(.a(gate159inter5), .b(gate159inter2), .O(gate159inter6));
  inv1  gate1632(.a(G444), .O(gate159inter7));
  inv1  gate1633(.a(G531), .O(gate159inter8));
  nand2 gate1634(.a(gate159inter8), .b(gate159inter7), .O(gate159inter9));
  nand2 gate1635(.a(s_155), .b(gate159inter3), .O(gate159inter10));
  nor2  gate1636(.a(gate159inter10), .b(gate159inter9), .O(gate159inter11));
  nor2  gate1637(.a(gate159inter11), .b(gate159inter6), .O(gate159inter12));
  nand2 gate1638(.a(gate159inter12), .b(gate159inter1), .O(G576));
nand2 gate160( .a(G447), .b(G531), .O(G577) );
nand2 gate161( .a(G450), .b(G534), .O(G578) );

  xor2  gate2143(.a(G534), .b(G453), .O(gate162inter0));
  nand2 gate2144(.a(gate162inter0), .b(s_228), .O(gate162inter1));
  and2  gate2145(.a(G534), .b(G453), .O(gate162inter2));
  inv1  gate2146(.a(s_228), .O(gate162inter3));
  inv1  gate2147(.a(s_229), .O(gate162inter4));
  nand2 gate2148(.a(gate162inter4), .b(gate162inter3), .O(gate162inter5));
  nor2  gate2149(.a(gate162inter5), .b(gate162inter2), .O(gate162inter6));
  inv1  gate2150(.a(G453), .O(gate162inter7));
  inv1  gate2151(.a(G534), .O(gate162inter8));
  nand2 gate2152(.a(gate162inter8), .b(gate162inter7), .O(gate162inter9));
  nand2 gate2153(.a(s_229), .b(gate162inter3), .O(gate162inter10));
  nor2  gate2154(.a(gate162inter10), .b(gate162inter9), .O(gate162inter11));
  nor2  gate2155(.a(gate162inter11), .b(gate162inter6), .O(gate162inter12));
  nand2 gate2156(.a(gate162inter12), .b(gate162inter1), .O(G579));
nand2 gate163( .a(G456), .b(G537), .O(G580) );

  xor2  gate869(.a(G537), .b(G459), .O(gate164inter0));
  nand2 gate870(.a(gate164inter0), .b(s_46), .O(gate164inter1));
  and2  gate871(.a(G537), .b(G459), .O(gate164inter2));
  inv1  gate872(.a(s_46), .O(gate164inter3));
  inv1  gate873(.a(s_47), .O(gate164inter4));
  nand2 gate874(.a(gate164inter4), .b(gate164inter3), .O(gate164inter5));
  nor2  gate875(.a(gate164inter5), .b(gate164inter2), .O(gate164inter6));
  inv1  gate876(.a(G459), .O(gate164inter7));
  inv1  gate877(.a(G537), .O(gate164inter8));
  nand2 gate878(.a(gate164inter8), .b(gate164inter7), .O(gate164inter9));
  nand2 gate879(.a(s_47), .b(gate164inter3), .O(gate164inter10));
  nor2  gate880(.a(gate164inter10), .b(gate164inter9), .O(gate164inter11));
  nor2  gate881(.a(gate164inter11), .b(gate164inter6), .O(gate164inter12));
  nand2 gate882(.a(gate164inter12), .b(gate164inter1), .O(G581));

  xor2  gate827(.a(G540), .b(G462), .O(gate165inter0));
  nand2 gate828(.a(gate165inter0), .b(s_40), .O(gate165inter1));
  and2  gate829(.a(G540), .b(G462), .O(gate165inter2));
  inv1  gate830(.a(s_40), .O(gate165inter3));
  inv1  gate831(.a(s_41), .O(gate165inter4));
  nand2 gate832(.a(gate165inter4), .b(gate165inter3), .O(gate165inter5));
  nor2  gate833(.a(gate165inter5), .b(gate165inter2), .O(gate165inter6));
  inv1  gate834(.a(G462), .O(gate165inter7));
  inv1  gate835(.a(G540), .O(gate165inter8));
  nand2 gate836(.a(gate165inter8), .b(gate165inter7), .O(gate165inter9));
  nand2 gate837(.a(s_41), .b(gate165inter3), .O(gate165inter10));
  nor2  gate838(.a(gate165inter10), .b(gate165inter9), .O(gate165inter11));
  nor2  gate839(.a(gate165inter11), .b(gate165inter6), .O(gate165inter12));
  nand2 gate840(.a(gate165inter12), .b(gate165inter1), .O(G582));
nand2 gate166( .a(G465), .b(G540), .O(G583) );
nand2 gate167( .a(G468), .b(G543), .O(G584) );
nand2 gate168( .a(G471), .b(G543), .O(G585) );
nand2 gate169( .a(G474), .b(G546), .O(G586) );
nand2 gate170( .a(G477), .b(G546), .O(G587) );
nand2 gate171( .a(G480), .b(G549), .O(G588) );
nand2 gate172( .a(G483), .b(G549), .O(G589) );
nand2 gate173( .a(G486), .b(G552), .O(G590) );
nand2 gate174( .a(G489), .b(G552), .O(G591) );

  xor2  gate953(.a(G555), .b(G492), .O(gate175inter0));
  nand2 gate954(.a(gate175inter0), .b(s_58), .O(gate175inter1));
  and2  gate955(.a(G555), .b(G492), .O(gate175inter2));
  inv1  gate956(.a(s_58), .O(gate175inter3));
  inv1  gate957(.a(s_59), .O(gate175inter4));
  nand2 gate958(.a(gate175inter4), .b(gate175inter3), .O(gate175inter5));
  nor2  gate959(.a(gate175inter5), .b(gate175inter2), .O(gate175inter6));
  inv1  gate960(.a(G492), .O(gate175inter7));
  inv1  gate961(.a(G555), .O(gate175inter8));
  nand2 gate962(.a(gate175inter8), .b(gate175inter7), .O(gate175inter9));
  nand2 gate963(.a(s_59), .b(gate175inter3), .O(gate175inter10));
  nor2  gate964(.a(gate175inter10), .b(gate175inter9), .O(gate175inter11));
  nor2  gate965(.a(gate175inter11), .b(gate175inter6), .O(gate175inter12));
  nand2 gate966(.a(gate175inter12), .b(gate175inter1), .O(G592));
nand2 gate176( .a(G495), .b(G555), .O(G593) );
nand2 gate177( .a(G498), .b(G558), .O(G594) );
nand2 gate178( .a(G501), .b(G558), .O(G595) );
nand2 gate179( .a(G504), .b(G561), .O(G596) );
nand2 gate180( .a(G507), .b(G561), .O(G597) );
nand2 gate181( .a(G510), .b(G564), .O(G598) );
nand2 gate182( .a(G513), .b(G564), .O(G599) );
nand2 gate183( .a(G516), .b(G567), .O(G600) );

  xor2  gate925(.a(G567), .b(G519), .O(gate184inter0));
  nand2 gate926(.a(gate184inter0), .b(s_54), .O(gate184inter1));
  and2  gate927(.a(G567), .b(G519), .O(gate184inter2));
  inv1  gate928(.a(s_54), .O(gate184inter3));
  inv1  gate929(.a(s_55), .O(gate184inter4));
  nand2 gate930(.a(gate184inter4), .b(gate184inter3), .O(gate184inter5));
  nor2  gate931(.a(gate184inter5), .b(gate184inter2), .O(gate184inter6));
  inv1  gate932(.a(G519), .O(gate184inter7));
  inv1  gate933(.a(G567), .O(gate184inter8));
  nand2 gate934(.a(gate184inter8), .b(gate184inter7), .O(gate184inter9));
  nand2 gate935(.a(s_55), .b(gate184inter3), .O(gate184inter10));
  nor2  gate936(.a(gate184inter10), .b(gate184inter9), .O(gate184inter11));
  nor2  gate937(.a(gate184inter11), .b(gate184inter6), .O(gate184inter12));
  nand2 gate938(.a(gate184inter12), .b(gate184inter1), .O(G601));

  xor2  gate1079(.a(G571), .b(G570), .O(gate185inter0));
  nand2 gate1080(.a(gate185inter0), .b(s_76), .O(gate185inter1));
  and2  gate1081(.a(G571), .b(G570), .O(gate185inter2));
  inv1  gate1082(.a(s_76), .O(gate185inter3));
  inv1  gate1083(.a(s_77), .O(gate185inter4));
  nand2 gate1084(.a(gate185inter4), .b(gate185inter3), .O(gate185inter5));
  nor2  gate1085(.a(gate185inter5), .b(gate185inter2), .O(gate185inter6));
  inv1  gate1086(.a(G570), .O(gate185inter7));
  inv1  gate1087(.a(G571), .O(gate185inter8));
  nand2 gate1088(.a(gate185inter8), .b(gate185inter7), .O(gate185inter9));
  nand2 gate1089(.a(s_77), .b(gate185inter3), .O(gate185inter10));
  nor2  gate1090(.a(gate185inter10), .b(gate185inter9), .O(gate185inter11));
  nor2  gate1091(.a(gate185inter11), .b(gate185inter6), .O(gate185inter12));
  nand2 gate1092(.a(gate185inter12), .b(gate185inter1), .O(G602));
nand2 gate186( .a(G572), .b(G573), .O(G607) );
nand2 gate187( .a(G574), .b(G575), .O(G612) );
nand2 gate188( .a(G576), .b(G577), .O(G617) );
nand2 gate189( .a(G578), .b(G579), .O(G622) );
nand2 gate190( .a(G580), .b(G581), .O(G627) );
nand2 gate191( .a(G582), .b(G583), .O(G632) );
nand2 gate192( .a(G584), .b(G585), .O(G637) );

  xor2  gate1849(.a(G587), .b(G586), .O(gate193inter0));
  nand2 gate1850(.a(gate193inter0), .b(s_186), .O(gate193inter1));
  and2  gate1851(.a(G587), .b(G586), .O(gate193inter2));
  inv1  gate1852(.a(s_186), .O(gate193inter3));
  inv1  gate1853(.a(s_187), .O(gate193inter4));
  nand2 gate1854(.a(gate193inter4), .b(gate193inter3), .O(gate193inter5));
  nor2  gate1855(.a(gate193inter5), .b(gate193inter2), .O(gate193inter6));
  inv1  gate1856(.a(G586), .O(gate193inter7));
  inv1  gate1857(.a(G587), .O(gate193inter8));
  nand2 gate1858(.a(gate193inter8), .b(gate193inter7), .O(gate193inter9));
  nand2 gate1859(.a(s_187), .b(gate193inter3), .O(gate193inter10));
  nor2  gate1860(.a(gate193inter10), .b(gate193inter9), .O(gate193inter11));
  nor2  gate1861(.a(gate193inter11), .b(gate193inter6), .O(gate193inter12));
  nand2 gate1862(.a(gate193inter12), .b(gate193inter1), .O(G642));

  xor2  gate1289(.a(G589), .b(G588), .O(gate194inter0));
  nand2 gate1290(.a(gate194inter0), .b(s_106), .O(gate194inter1));
  and2  gate1291(.a(G589), .b(G588), .O(gate194inter2));
  inv1  gate1292(.a(s_106), .O(gate194inter3));
  inv1  gate1293(.a(s_107), .O(gate194inter4));
  nand2 gate1294(.a(gate194inter4), .b(gate194inter3), .O(gate194inter5));
  nor2  gate1295(.a(gate194inter5), .b(gate194inter2), .O(gate194inter6));
  inv1  gate1296(.a(G588), .O(gate194inter7));
  inv1  gate1297(.a(G589), .O(gate194inter8));
  nand2 gate1298(.a(gate194inter8), .b(gate194inter7), .O(gate194inter9));
  nand2 gate1299(.a(s_107), .b(gate194inter3), .O(gate194inter10));
  nor2  gate1300(.a(gate194inter10), .b(gate194inter9), .O(gate194inter11));
  nor2  gate1301(.a(gate194inter11), .b(gate194inter6), .O(gate194inter12));
  nand2 gate1302(.a(gate194inter12), .b(gate194inter1), .O(G645));
nand2 gate195( .a(G590), .b(G591), .O(G648) );

  xor2  gate589(.a(G593), .b(G592), .O(gate196inter0));
  nand2 gate590(.a(gate196inter0), .b(s_6), .O(gate196inter1));
  and2  gate591(.a(G593), .b(G592), .O(gate196inter2));
  inv1  gate592(.a(s_6), .O(gate196inter3));
  inv1  gate593(.a(s_7), .O(gate196inter4));
  nand2 gate594(.a(gate196inter4), .b(gate196inter3), .O(gate196inter5));
  nor2  gate595(.a(gate196inter5), .b(gate196inter2), .O(gate196inter6));
  inv1  gate596(.a(G592), .O(gate196inter7));
  inv1  gate597(.a(G593), .O(gate196inter8));
  nand2 gate598(.a(gate196inter8), .b(gate196inter7), .O(gate196inter9));
  nand2 gate599(.a(s_7), .b(gate196inter3), .O(gate196inter10));
  nor2  gate600(.a(gate196inter10), .b(gate196inter9), .O(gate196inter11));
  nor2  gate601(.a(gate196inter11), .b(gate196inter6), .O(gate196inter12));
  nand2 gate602(.a(gate196inter12), .b(gate196inter1), .O(G651));
nand2 gate197( .a(G594), .b(G595), .O(G654) );
nand2 gate198( .a(G596), .b(G597), .O(G657) );
nand2 gate199( .a(G598), .b(G599), .O(G660) );
nand2 gate200( .a(G600), .b(G601), .O(G663) );
nand2 gate201( .a(G602), .b(G607), .O(G666) );
nand2 gate202( .a(G612), .b(G617), .O(G669) );
nand2 gate203( .a(G602), .b(G612), .O(G672) );
nand2 gate204( .a(G607), .b(G617), .O(G675) );
nand2 gate205( .a(G622), .b(G627), .O(G678) );

  xor2  gate1401(.a(G637), .b(G632), .O(gate206inter0));
  nand2 gate1402(.a(gate206inter0), .b(s_122), .O(gate206inter1));
  and2  gate1403(.a(G637), .b(G632), .O(gate206inter2));
  inv1  gate1404(.a(s_122), .O(gate206inter3));
  inv1  gate1405(.a(s_123), .O(gate206inter4));
  nand2 gate1406(.a(gate206inter4), .b(gate206inter3), .O(gate206inter5));
  nor2  gate1407(.a(gate206inter5), .b(gate206inter2), .O(gate206inter6));
  inv1  gate1408(.a(G632), .O(gate206inter7));
  inv1  gate1409(.a(G637), .O(gate206inter8));
  nand2 gate1410(.a(gate206inter8), .b(gate206inter7), .O(gate206inter9));
  nand2 gate1411(.a(s_123), .b(gate206inter3), .O(gate206inter10));
  nor2  gate1412(.a(gate206inter10), .b(gate206inter9), .O(gate206inter11));
  nor2  gate1413(.a(gate206inter11), .b(gate206inter6), .O(gate206inter12));
  nand2 gate1414(.a(gate206inter12), .b(gate206inter1), .O(G681));
nand2 gate207( .a(G622), .b(G632), .O(G684) );
nand2 gate208( .a(G627), .b(G637), .O(G687) );
nand2 gate209( .a(G602), .b(G666), .O(G690) );

  xor2  gate1107(.a(G666), .b(G607), .O(gate210inter0));
  nand2 gate1108(.a(gate210inter0), .b(s_80), .O(gate210inter1));
  and2  gate1109(.a(G666), .b(G607), .O(gate210inter2));
  inv1  gate1110(.a(s_80), .O(gate210inter3));
  inv1  gate1111(.a(s_81), .O(gate210inter4));
  nand2 gate1112(.a(gate210inter4), .b(gate210inter3), .O(gate210inter5));
  nor2  gate1113(.a(gate210inter5), .b(gate210inter2), .O(gate210inter6));
  inv1  gate1114(.a(G607), .O(gate210inter7));
  inv1  gate1115(.a(G666), .O(gate210inter8));
  nand2 gate1116(.a(gate210inter8), .b(gate210inter7), .O(gate210inter9));
  nand2 gate1117(.a(s_81), .b(gate210inter3), .O(gate210inter10));
  nor2  gate1118(.a(gate210inter10), .b(gate210inter9), .O(gate210inter11));
  nor2  gate1119(.a(gate210inter11), .b(gate210inter6), .O(gate210inter12));
  nand2 gate1120(.a(gate210inter12), .b(gate210inter1), .O(G691));
nand2 gate211( .a(G612), .b(G669), .O(G692) );

  xor2  gate1751(.a(G669), .b(G617), .O(gate212inter0));
  nand2 gate1752(.a(gate212inter0), .b(s_172), .O(gate212inter1));
  and2  gate1753(.a(G669), .b(G617), .O(gate212inter2));
  inv1  gate1754(.a(s_172), .O(gate212inter3));
  inv1  gate1755(.a(s_173), .O(gate212inter4));
  nand2 gate1756(.a(gate212inter4), .b(gate212inter3), .O(gate212inter5));
  nor2  gate1757(.a(gate212inter5), .b(gate212inter2), .O(gate212inter6));
  inv1  gate1758(.a(G617), .O(gate212inter7));
  inv1  gate1759(.a(G669), .O(gate212inter8));
  nand2 gate1760(.a(gate212inter8), .b(gate212inter7), .O(gate212inter9));
  nand2 gate1761(.a(s_173), .b(gate212inter3), .O(gate212inter10));
  nor2  gate1762(.a(gate212inter10), .b(gate212inter9), .O(gate212inter11));
  nor2  gate1763(.a(gate212inter11), .b(gate212inter6), .O(gate212inter12));
  nand2 gate1764(.a(gate212inter12), .b(gate212inter1), .O(G693));
nand2 gate213( .a(G602), .b(G672), .O(G694) );

  xor2  gate1653(.a(G672), .b(G612), .O(gate214inter0));
  nand2 gate1654(.a(gate214inter0), .b(s_158), .O(gate214inter1));
  and2  gate1655(.a(G672), .b(G612), .O(gate214inter2));
  inv1  gate1656(.a(s_158), .O(gate214inter3));
  inv1  gate1657(.a(s_159), .O(gate214inter4));
  nand2 gate1658(.a(gate214inter4), .b(gate214inter3), .O(gate214inter5));
  nor2  gate1659(.a(gate214inter5), .b(gate214inter2), .O(gate214inter6));
  inv1  gate1660(.a(G612), .O(gate214inter7));
  inv1  gate1661(.a(G672), .O(gate214inter8));
  nand2 gate1662(.a(gate214inter8), .b(gate214inter7), .O(gate214inter9));
  nand2 gate1663(.a(s_159), .b(gate214inter3), .O(gate214inter10));
  nor2  gate1664(.a(gate214inter10), .b(gate214inter9), .O(gate214inter11));
  nor2  gate1665(.a(gate214inter11), .b(gate214inter6), .O(gate214inter12));
  nand2 gate1666(.a(gate214inter12), .b(gate214inter1), .O(G695));

  xor2  gate547(.a(G675), .b(G607), .O(gate215inter0));
  nand2 gate548(.a(gate215inter0), .b(s_0), .O(gate215inter1));
  and2  gate549(.a(G675), .b(G607), .O(gate215inter2));
  inv1  gate550(.a(s_0), .O(gate215inter3));
  inv1  gate551(.a(s_1), .O(gate215inter4));
  nand2 gate552(.a(gate215inter4), .b(gate215inter3), .O(gate215inter5));
  nor2  gate553(.a(gate215inter5), .b(gate215inter2), .O(gate215inter6));
  inv1  gate554(.a(G607), .O(gate215inter7));
  inv1  gate555(.a(G675), .O(gate215inter8));
  nand2 gate556(.a(gate215inter8), .b(gate215inter7), .O(gate215inter9));
  nand2 gate557(.a(s_1), .b(gate215inter3), .O(gate215inter10));
  nor2  gate558(.a(gate215inter10), .b(gate215inter9), .O(gate215inter11));
  nor2  gate559(.a(gate215inter11), .b(gate215inter6), .O(gate215inter12));
  nand2 gate560(.a(gate215inter12), .b(gate215inter1), .O(G696));
nand2 gate216( .a(G617), .b(G675), .O(G697) );

  xor2  gate897(.a(G678), .b(G622), .O(gate217inter0));
  nand2 gate898(.a(gate217inter0), .b(s_50), .O(gate217inter1));
  and2  gate899(.a(G678), .b(G622), .O(gate217inter2));
  inv1  gate900(.a(s_50), .O(gate217inter3));
  inv1  gate901(.a(s_51), .O(gate217inter4));
  nand2 gate902(.a(gate217inter4), .b(gate217inter3), .O(gate217inter5));
  nor2  gate903(.a(gate217inter5), .b(gate217inter2), .O(gate217inter6));
  inv1  gate904(.a(G622), .O(gate217inter7));
  inv1  gate905(.a(G678), .O(gate217inter8));
  nand2 gate906(.a(gate217inter8), .b(gate217inter7), .O(gate217inter9));
  nand2 gate907(.a(s_51), .b(gate217inter3), .O(gate217inter10));
  nor2  gate908(.a(gate217inter10), .b(gate217inter9), .O(gate217inter11));
  nor2  gate909(.a(gate217inter11), .b(gate217inter6), .O(gate217inter12));
  nand2 gate910(.a(gate217inter12), .b(gate217inter1), .O(G698));
nand2 gate218( .a(G627), .b(G678), .O(G699) );
nand2 gate219( .a(G632), .b(G681), .O(G700) );

  xor2  gate1569(.a(G681), .b(G637), .O(gate220inter0));
  nand2 gate1570(.a(gate220inter0), .b(s_146), .O(gate220inter1));
  and2  gate1571(.a(G681), .b(G637), .O(gate220inter2));
  inv1  gate1572(.a(s_146), .O(gate220inter3));
  inv1  gate1573(.a(s_147), .O(gate220inter4));
  nand2 gate1574(.a(gate220inter4), .b(gate220inter3), .O(gate220inter5));
  nor2  gate1575(.a(gate220inter5), .b(gate220inter2), .O(gate220inter6));
  inv1  gate1576(.a(G637), .O(gate220inter7));
  inv1  gate1577(.a(G681), .O(gate220inter8));
  nand2 gate1578(.a(gate220inter8), .b(gate220inter7), .O(gate220inter9));
  nand2 gate1579(.a(s_147), .b(gate220inter3), .O(gate220inter10));
  nor2  gate1580(.a(gate220inter10), .b(gate220inter9), .O(gate220inter11));
  nor2  gate1581(.a(gate220inter11), .b(gate220inter6), .O(gate220inter12));
  nand2 gate1582(.a(gate220inter12), .b(gate220inter1), .O(G701));
nand2 gate221( .a(G622), .b(G684), .O(G702) );
nand2 gate222( .a(G632), .b(G684), .O(G703) );

  xor2  gate2003(.a(G687), .b(G627), .O(gate223inter0));
  nand2 gate2004(.a(gate223inter0), .b(s_208), .O(gate223inter1));
  and2  gate2005(.a(G687), .b(G627), .O(gate223inter2));
  inv1  gate2006(.a(s_208), .O(gate223inter3));
  inv1  gate2007(.a(s_209), .O(gate223inter4));
  nand2 gate2008(.a(gate223inter4), .b(gate223inter3), .O(gate223inter5));
  nor2  gate2009(.a(gate223inter5), .b(gate223inter2), .O(gate223inter6));
  inv1  gate2010(.a(G627), .O(gate223inter7));
  inv1  gate2011(.a(G687), .O(gate223inter8));
  nand2 gate2012(.a(gate223inter8), .b(gate223inter7), .O(gate223inter9));
  nand2 gate2013(.a(s_209), .b(gate223inter3), .O(gate223inter10));
  nor2  gate2014(.a(gate223inter10), .b(gate223inter9), .O(gate223inter11));
  nor2  gate2015(.a(gate223inter11), .b(gate223inter6), .O(gate223inter12));
  nand2 gate2016(.a(gate223inter12), .b(gate223inter1), .O(G704));
nand2 gate224( .a(G637), .b(G687), .O(G705) );
nand2 gate225( .a(G690), .b(G691), .O(G706) );
nand2 gate226( .a(G692), .b(G693), .O(G709) );
nand2 gate227( .a(G694), .b(G695), .O(G712) );
nand2 gate228( .a(G696), .b(G697), .O(G715) );

  xor2  gate1919(.a(G699), .b(G698), .O(gate229inter0));
  nand2 gate1920(.a(gate229inter0), .b(s_196), .O(gate229inter1));
  and2  gate1921(.a(G699), .b(G698), .O(gate229inter2));
  inv1  gate1922(.a(s_196), .O(gate229inter3));
  inv1  gate1923(.a(s_197), .O(gate229inter4));
  nand2 gate1924(.a(gate229inter4), .b(gate229inter3), .O(gate229inter5));
  nor2  gate1925(.a(gate229inter5), .b(gate229inter2), .O(gate229inter6));
  inv1  gate1926(.a(G698), .O(gate229inter7));
  inv1  gate1927(.a(G699), .O(gate229inter8));
  nand2 gate1928(.a(gate229inter8), .b(gate229inter7), .O(gate229inter9));
  nand2 gate1929(.a(s_197), .b(gate229inter3), .O(gate229inter10));
  nor2  gate1930(.a(gate229inter10), .b(gate229inter9), .O(gate229inter11));
  nor2  gate1931(.a(gate229inter11), .b(gate229inter6), .O(gate229inter12));
  nand2 gate1932(.a(gate229inter12), .b(gate229inter1), .O(G718));

  xor2  gate1373(.a(G701), .b(G700), .O(gate230inter0));
  nand2 gate1374(.a(gate230inter0), .b(s_118), .O(gate230inter1));
  and2  gate1375(.a(G701), .b(G700), .O(gate230inter2));
  inv1  gate1376(.a(s_118), .O(gate230inter3));
  inv1  gate1377(.a(s_119), .O(gate230inter4));
  nand2 gate1378(.a(gate230inter4), .b(gate230inter3), .O(gate230inter5));
  nor2  gate1379(.a(gate230inter5), .b(gate230inter2), .O(gate230inter6));
  inv1  gate1380(.a(G700), .O(gate230inter7));
  inv1  gate1381(.a(G701), .O(gate230inter8));
  nand2 gate1382(.a(gate230inter8), .b(gate230inter7), .O(gate230inter9));
  nand2 gate1383(.a(s_119), .b(gate230inter3), .O(gate230inter10));
  nor2  gate1384(.a(gate230inter10), .b(gate230inter9), .O(gate230inter11));
  nor2  gate1385(.a(gate230inter11), .b(gate230inter6), .O(gate230inter12));
  nand2 gate1386(.a(gate230inter12), .b(gate230inter1), .O(G721));
nand2 gate231( .a(G702), .b(G703), .O(G724) );

  xor2  gate1975(.a(G705), .b(G704), .O(gate232inter0));
  nand2 gate1976(.a(gate232inter0), .b(s_204), .O(gate232inter1));
  and2  gate1977(.a(G705), .b(G704), .O(gate232inter2));
  inv1  gate1978(.a(s_204), .O(gate232inter3));
  inv1  gate1979(.a(s_205), .O(gate232inter4));
  nand2 gate1980(.a(gate232inter4), .b(gate232inter3), .O(gate232inter5));
  nor2  gate1981(.a(gate232inter5), .b(gate232inter2), .O(gate232inter6));
  inv1  gate1982(.a(G704), .O(gate232inter7));
  inv1  gate1983(.a(G705), .O(gate232inter8));
  nand2 gate1984(.a(gate232inter8), .b(gate232inter7), .O(gate232inter9));
  nand2 gate1985(.a(s_205), .b(gate232inter3), .O(gate232inter10));
  nor2  gate1986(.a(gate232inter10), .b(gate232inter9), .O(gate232inter11));
  nor2  gate1987(.a(gate232inter11), .b(gate232inter6), .O(gate232inter12));
  nand2 gate1988(.a(gate232inter12), .b(gate232inter1), .O(G727));
nand2 gate233( .a(G242), .b(G718), .O(G730) );

  xor2  gate1737(.a(G721), .b(G245), .O(gate234inter0));
  nand2 gate1738(.a(gate234inter0), .b(s_170), .O(gate234inter1));
  and2  gate1739(.a(G721), .b(G245), .O(gate234inter2));
  inv1  gate1740(.a(s_170), .O(gate234inter3));
  inv1  gate1741(.a(s_171), .O(gate234inter4));
  nand2 gate1742(.a(gate234inter4), .b(gate234inter3), .O(gate234inter5));
  nor2  gate1743(.a(gate234inter5), .b(gate234inter2), .O(gate234inter6));
  inv1  gate1744(.a(G245), .O(gate234inter7));
  inv1  gate1745(.a(G721), .O(gate234inter8));
  nand2 gate1746(.a(gate234inter8), .b(gate234inter7), .O(gate234inter9));
  nand2 gate1747(.a(s_171), .b(gate234inter3), .O(gate234inter10));
  nor2  gate1748(.a(gate234inter10), .b(gate234inter9), .O(gate234inter11));
  nor2  gate1749(.a(gate234inter11), .b(gate234inter6), .O(gate234inter12));
  nand2 gate1750(.a(gate234inter12), .b(gate234inter1), .O(G733));

  xor2  gate967(.a(G724), .b(G248), .O(gate235inter0));
  nand2 gate968(.a(gate235inter0), .b(s_60), .O(gate235inter1));
  and2  gate969(.a(G724), .b(G248), .O(gate235inter2));
  inv1  gate970(.a(s_60), .O(gate235inter3));
  inv1  gate971(.a(s_61), .O(gate235inter4));
  nand2 gate972(.a(gate235inter4), .b(gate235inter3), .O(gate235inter5));
  nor2  gate973(.a(gate235inter5), .b(gate235inter2), .O(gate235inter6));
  inv1  gate974(.a(G248), .O(gate235inter7));
  inv1  gate975(.a(G724), .O(gate235inter8));
  nand2 gate976(.a(gate235inter8), .b(gate235inter7), .O(gate235inter9));
  nand2 gate977(.a(s_61), .b(gate235inter3), .O(gate235inter10));
  nor2  gate978(.a(gate235inter10), .b(gate235inter9), .O(gate235inter11));
  nor2  gate979(.a(gate235inter11), .b(gate235inter6), .O(gate235inter12));
  nand2 gate980(.a(gate235inter12), .b(gate235inter1), .O(G736));
nand2 gate236( .a(G251), .b(G727), .O(G739) );
nand2 gate237( .a(G254), .b(G706), .O(G742) );
nand2 gate238( .a(G257), .b(G709), .O(G745) );
nand2 gate239( .a(G260), .b(G712), .O(G748) );

  xor2  gate1541(.a(G715), .b(G263), .O(gate240inter0));
  nand2 gate1542(.a(gate240inter0), .b(s_142), .O(gate240inter1));
  and2  gate1543(.a(G715), .b(G263), .O(gate240inter2));
  inv1  gate1544(.a(s_142), .O(gate240inter3));
  inv1  gate1545(.a(s_143), .O(gate240inter4));
  nand2 gate1546(.a(gate240inter4), .b(gate240inter3), .O(gate240inter5));
  nor2  gate1547(.a(gate240inter5), .b(gate240inter2), .O(gate240inter6));
  inv1  gate1548(.a(G263), .O(gate240inter7));
  inv1  gate1549(.a(G715), .O(gate240inter8));
  nand2 gate1550(.a(gate240inter8), .b(gate240inter7), .O(gate240inter9));
  nand2 gate1551(.a(s_143), .b(gate240inter3), .O(gate240inter10));
  nor2  gate1552(.a(gate240inter10), .b(gate240inter9), .O(gate240inter11));
  nor2  gate1553(.a(gate240inter11), .b(gate240inter6), .O(gate240inter12));
  nand2 gate1554(.a(gate240inter12), .b(gate240inter1), .O(G751));
nand2 gate241( .a(G242), .b(G730), .O(G754) );
nand2 gate242( .a(G718), .b(G730), .O(G755) );
nand2 gate243( .a(G245), .b(G733), .O(G756) );
nand2 gate244( .a(G721), .b(G733), .O(G757) );
nand2 gate245( .a(G248), .b(G736), .O(G758) );

  xor2  gate1415(.a(G736), .b(G724), .O(gate246inter0));
  nand2 gate1416(.a(gate246inter0), .b(s_124), .O(gate246inter1));
  and2  gate1417(.a(G736), .b(G724), .O(gate246inter2));
  inv1  gate1418(.a(s_124), .O(gate246inter3));
  inv1  gate1419(.a(s_125), .O(gate246inter4));
  nand2 gate1420(.a(gate246inter4), .b(gate246inter3), .O(gate246inter5));
  nor2  gate1421(.a(gate246inter5), .b(gate246inter2), .O(gate246inter6));
  inv1  gate1422(.a(G724), .O(gate246inter7));
  inv1  gate1423(.a(G736), .O(gate246inter8));
  nand2 gate1424(.a(gate246inter8), .b(gate246inter7), .O(gate246inter9));
  nand2 gate1425(.a(s_125), .b(gate246inter3), .O(gate246inter10));
  nor2  gate1426(.a(gate246inter10), .b(gate246inter9), .O(gate246inter11));
  nor2  gate1427(.a(gate246inter11), .b(gate246inter6), .O(gate246inter12));
  nand2 gate1428(.a(gate246inter12), .b(gate246inter1), .O(G759));
nand2 gate247( .a(G251), .b(G739), .O(G760) );
nand2 gate248( .a(G727), .b(G739), .O(G761) );
nand2 gate249( .a(G254), .b(G742), .O(G762) );
nand2 gate250( .a(G706), .b(G742), .O(G763) );
nand2 gate251( .a(G257), .b(G745), .O(G764) );
nand2 gate252( .a(G709), .b(G745), .O(G765) );

  xor2  gate1611(.a(G748), .b(G260), .O(gate253inter0));
  nand2 gate1612(.a(gate253inter0), .b(s_152), .O(gate253inter1));
  and2  gate1613(.a(G748), .b(G260), .O(gate253inter2));
  inv1  gate1614(.a(s_152), .O(gate253inter3));
  inv1  gate1615(.a(s_153), .O(gate253inter4));
  nand2 gate1616(.a(gate253inter4), .b(gate253inter3), .O(gate253inter5));
  nor2  gate1617(.a(gate253inter5), .b(gate253inter2), .O(gate253inter6));
  inv1  gate1618(.a(G260), .O(gate253inter7));
  inv1  gate1619(.a(G748), .O(gate253inter8));
  nand2 gate1620(.a(gate253inter8), .b(gate253inter7), .O(gate253inter9));
  nand2 gate1621(.a(s_153), .b(gate253inter3), .O(gate253inter10));
  nor2  gate1622(.a(gate253inter10), .b(gate253inter9), .O(gate253inter11));
  nor2  gate1623(.a(gate253inter11), .b(gate253inter6), .O(gate253inter12));
  nand2 gate1624(.a(gate253inter12), .b(gate253inter1), .O(G766));

  xor2  gate1667(.a(G748), .b(G712), .O(gate254inter0));
  nand2 gate1668(.a(gate254inter0), .b(s_160), .O(gate254inter1));
  and2  gate1669(.a(G748), .b(G712), .O(gate254inter2));
  inv1  gate1670(.a(s_160), .O(gate254inter3));
  inv1  gate1671(.a(s_161), .O(gate254inter4));
  nand2 gate1672(.a(gate254inter4), .b(gate254inter3), .O(gate254inter5));
  nor2  gate1673(.a(gate254inter5), .b(gate254inter2), .O(gate254inter6));
  inv1  gate1674(.a(G712), .O(gate254inter7));
  inv1  gate1675(.a(G748), .O(gate254inter8));
  nand2 gate1676(.a(gate254inter8), .b(gate254inter7), .O(gate254inter9));
  nand2 gate1677(.a(s_161), .b(gate254inter3), .O(gate254inter10));
  nor2  gate1678(.a(gate254inter10), .b(gate254inter9), .O(gate254inter11));
  nor2  gate1679(.a(gate254inter11), .b(gate254inter6), .O(gate254inter12));
  nand2 gate1680(.a(gate254inter12), .b(gate254inter1), .O(G767));
nand2 gate255( .a(G263), .b(G751), .O(G768) );

  xor2  gate1723(.a(G751), .b(G715), .O(gate256inter0));
  nand2 gate1724(.a(gate256inter0), .b(s_168), .O(gate256inter1));
  and2  gate1725(.a(G751), .b(G715), .O(gate256inter2));
  inv1  gate1726(.a(s_168), .O(gate256inter3));
  inv1  gate1727(.a(s_169), .O(gate256inter4));
  nand2 gate1728(.a(gate256inter4), .b(gate256inter3), .O(gate256inter5));
  nor2  gate1729(.a(gate256inter5), .b(gate256inter2), .O(gate256inter6));
  inv1  gate1730(.a(G715), .O(gate256inter7));
  inv1  gate1731(.a(G751), .O(gate256inter8));
  nand2 gate1732(.a(gate256inter8), .b(gate256inter7), .O(gate256inter9));
  nand2 gate1733(.a(s_169), .b(gate256inter3), .O(gate256inter10));
  nor2  gate1734(.a(gate256inter10), .b(gate256inter9), .O(gate256inter11));
  nor2  gate1735(.a(gate256inter11), .b(gate256inter6), .O(gate256inter12));
  nand2 gate1736(.a(gate256inter12), .b(gate256inter1), .O(G769));

  xor2  gate1821(.a(G755), .b(G754), .O(gate257inter0));
  nand2 gate1822(.a(gate257inter0), .b(s_182), .O(gate257inter1));
  and2  gate1823(.a(G755), .b(G754), .O(gate257inter2));
  inv1  gate1824(.a(s_182), .O(gate257inter3));
  inv1  gate1825(.a(s_183), .O(gate257inter4));
  nand2 gate1826(.a(gate257inter4), .b(gate257inter3), .O(gate257inter5));
  nor2  gate1827(.a(gate257inter5), .b(gate257inter2), .O(gate257inter6));
  inv1  gate1828(.a(G754), .O(gate257inter7));
  inv1  gate1829(.a(G755), .O(gate257inter8));
  nand2 gate1830(.a(gate257inter8), .b(gate257inter7), .O(gate257inter9));
  nand2 gate1831(.a(s_183), .b(gate257inter3), .O(gate257inter10));
  nor2  gate1832(.a(gate257inter10), .b(gate257inter9), .O(gate257inter11));
  nor2  gate1833(.a(gate257inter11), .b(gate257inter6), .O(gate257inter12));
  nand2 gate1834(.a(gate257inter12), .b(gate257inter1), .O(G770));
nand2 gate258( .a(G756), .b(G757), .O(G773) );
nand2 gate259( .a(G758), .b(G759), .O(G776) );
nand2 gate260( .a(G760), .b(G761), .O(G779) );
nand2 gate261( .a(G762), .b(G763), .O(G782) );

  xor2  gate715(.a(G765), .b(G764), .O(gate262inter0));
  nand2 gate716(.a(gate262inter0), .b(s_24), .O(gate262inter1));
  and2  gate717(.a(G765), .b(G764), .O(gate262inter2));
  inv1  gate718(.a(s_24), .O(gate262inter3));
  inv1  gate719(.a(s_25), .O(gate262inter4));
  nand2 gate720(.a(gate262inter4), .b(gate262inter3), .O(gate262inter5));
  nor2  gate721(.a(gate262inter5), .b(gate262inter2), .O(gate262inter6));
  inv1  gate722(.a(G764), .O(gate262inter7));
  inv1  gate723(.a(G765), .O(gate262inter8));
  nand2 gate724(.a(gate262inter8), .b(gate262inter7), .O(gate262inter9));
  nand2 gate725(.a(s_25), .b(gate262inter3), .O(gate262inter10));
  nor2  gate726(.a(gate262inter10), .b(gate262inter9), .O(gate262inter11));
  nor2  gate727(.a(gate262inter11), .b(gate262inter6), .O(gate262inter12));
  nand2 gate728(.a(gate262inter12), .b(gate262inter1), .O(G785));
nand2 gate263( .a(G766), .b(G767), .O(G788) );
nand2 gate264( .a(G768), .b(G769), .O(G791) );
nand2 gate265( .a(G642), .b(G770), .O(G794) );

  xor2  gate1779(.a(G773), .b(G645), .O(gate266inter0));
  nand2 gate1780(.a(gate266inter0), .b(s_176), .O(gate266inter1));
  and2  gate1781(.a(G773), .b(G645), .O(gate266inter2));
  inv1  gate1782(.a(s_176), .O(gate266inter3));
  inv1  gate1783(.a(s_177), .O(gate266inter4));
  nand2 gate1784(.a(gate266inter4), .b(gate266inter3), .O(gate266inter5));
  nor2  gate1785(.a(gate266inter5), .b(gate266inter2), .O(gate266inter6));
  inv1  gate1786(.a(G645), .O(gate266inter7));
  inv1  gate1787(.a(G773), .O(gate266inter8));
  nand2 gate1788(.a(gate266inter8), .b(gate266inter7), .O(gate266inter9));
  nand2 gate1789(.a(s_177), .b(gate266inter3), .O(gate266inter10));
  nor2  gate1790(.a(gate266inter10), .b(gate266inter9), .O(gate266inter11));
  nor2  gate1791(.a(gate266inter11), .b(gate266inter6), .O(gate266inter12));
  nand2 gate1792(.a(gate266inter12), .b(gate266inter1), .O(G797));
nand2 gate267( .a(G648), .b(G776), .O(G800) );

  xor2  gate981(.a(G779), .b(G651), .O(gate268inter0));
  nand2 gate982(.a(gate268inter0), .b(s_62), .O(gate268inter1));
  and2  gate983(.a(G779), .b(G651), .O(gate268inter2));
  inv1  gate984(.a(s_62), .O(gate268inter3));
  inv1  gate985(.a(s_63), .O(gate268inter4));
  nand2 gate986(.a(gate268inter4), .b(gate268inter3), .O(gate268inter5));
  nor2  gate987(.a(gate268inter5), .b(gate268inter2), .O(gate268inter6));
  inv1  gate988(.a(G651), .O(gate268inter7));
  inv1  gate989(.a(G779), .O(gate268inter8));
  nand2 gate990(.a(gate268inter8), .b(gate268inter7), .O(gate268inter9));
  nand2 gate991(.a(s_63), .b(gate268inter3), .O(gate268inter10));
  nor2  gate992(.a(gate268inter10), .b(gate268inter9), .O(gate268inter11));
  nor2  gate993(.a(gate268inter11), .b(gate268inter6), .O(gate268inter12));
  nand2 gate994(.a(gate268inter12), .b(gate268inter1), .O(G803));
nand2 gate269( .a(G654), .b(G782), .O(G806) );
nand2 gate270( .a(G657), .b(G785), .O(G809) );
nand2 gate271( .a(G660), .b(G788), .O(G812) );

  xor2  gate1457(.a(G791), .b(G663), .O(gate272inter0));
  nand2 gate1458(.a(gate272inter0), .b(s_130), .O(gate272inter1));
  and2  gate1459(.a(G791), .b(G663), .O(gate272inter2));
  inv1  gate1460(.a(s_130), .O(gate272inter3));
  inv1  gate1461(.a(s_131), .O(gate272inter4));
  nand2 gate1462(.a(gate272inter4), .b(gate272inter3), .O(gate272inter5));
  nor2  gate1463(.a(gate272inter5), .b(gate272inter2), .O(gate272inter6));
  inv1  gate1464(.a(G663), .O(gate272inter7));
  inv1  gate1465(.a(G791), .O(gate272inter8));
  nand2 gate1466(.a(gate272inter8), .b(gate272inter7), .O(gate272inter9));
  nand2 gate1467(.a(s_131), .b(gate272inter3), .O(gate272inter10));
  nor2  gate1468(.a(gate272inter10), .b(gate272inter9), .O(gate272inter11));
  nor2  gate1469(.a(gate272inter11), .b(gate272inter6), .O(gate272inter12));
  nand2 gate1470(.a(gate272inter12), .b(gate272inter1), .O(G815));
nand2 gate273( .a(G642), .b(G794), .O(G818) );
nand2 gate274( .a(G770), .b(G794), .O(G819) );
nand2 gate275( .a(G645), .b(G797), .O(G820) );
nand2 gate276( .a(G773), .b(G797), .O(G821) );
nand2 gate277( .a(G648), .b(G800), .O(G822) );
nand2 gate278( .a(G776), .b(G800), .O(G823) );

  xor2  gate1877(.a(G803), .b(G651), .O(gate279inter0));
  nand2 gate1878(.a(gate279inter0), .b(s_190), .O(gate279inter1));
  and2  gate1879(.a(G803), .b(G651), .O(gate279inter2));
  inv1  gate1880(.a(s_190), .O(gate279inter3));
  inv1  gate1881(.a(s_191), .O(gate279inter4));
  nand2 gate1882(.a(gate279inter4), .b(gate279inter3), .O(gate279inter5));
  nor2  gate1883(.a(gate279inter5), .b(gate279inter2), .O(gate279inter6));
  inv1  gate1884(.a(G651), .O(gate279inter7));
  inv1  gate1885(.a(G803), .O(gate279inter8));
  nand2 gate1886(.a(gate279inter8), .b(gate279inter7), .O(gate279inter9));
  nand2 gate1887(.a(s_191), .b(gate279inter3), .O(gate279inter10));
  nor2  gate1888(.a(gate279inter10), .b(gate279inter9), .O(gate279inter11));
  nor2  gate1889(.a(gate279inter11), .b(gate279inter6), .O(gate279inter12));
  nand2 gate1890(.a(gate279inter12), .b(gate279inter1), .O(G824));

  xor2  gate771(.a(G803), .b(G779), .O(gate280inter0));
  nand2 gate772(.a(gate280inter0), .b(s_32), .O(gate280inter1));
  and2  gate773(.a(G803), .b(G779), .O(gate280inter2));
  inv1  gate774(.a(s_32), .O(gate280inter3));
  inv1  gate775(.a(s_33), .O(gate280inter4));
  nand2 gate776(.a(gate280inter4), .b(gate280inter3), .O(gate280inter5));
  nor2  gate777(.a(gate280inter5), .b(gate280inter2), .O(gate280inter6));
  inv1  gate778(.a(G779), .O(gate280inter7));
  inv1  gate779(.a(G803), .O(gate280inter8));
  nand2 gate780(.a(gate280inter8), .b(gate280inter7), .O(gate280inter9));
  nand2 gate781(.a(s_33), .b(gate280inter3), .O(gate280inter10));
  nor2  gate782(.a(gate280inter10), .b(gate280inter9), .O(gate280inter11));
  nor2  gate783(.a(gate280inter11), .b(gate280inter6), .O(gate280inter12));
  nand2 gate784(.a(gate280inter12), .b(gate280inter1), .O(G825));
nand2 gate281( .a(G654), .b(G806), .O(G826) );
nand2 gate282( .a(G782), .b(G806), .O(G827) );

  xor2  gate1499(.a(G809), .b(G657), .O(gate283inter0));
  nand2 gate1500(.a(gate283inter0), .b(s_136), .O(gate283inter1));
  and2  gate1501(.a(G809), .b(G657), .O(gate283inter2));
  inv1  gate1502(.a(s_136), .O(gate283inter3));
  inv1  gate1503(.a(s_137), .O(gate283inter4));
  nand2 gate1504(.a(gate283inter4), .b(gate283inter3), .O(gate283inter5));
  nor2  gate1505(.a(gate283inter5), .b(gate283inter2), .O(gate283inter6));
  inv1  gate1506(.a(G657), .O(gate283inter7));
  inv1  gate1507(.a(G809), .O(gate283inter8));
  nand2 gate1508(.a(gate283inter8), .b(gate283inter7), .O(gate283inter9));
  nand2 gate1509(.a(s_137), .b(gate283inter3), .O(gate283inter10));
  nor2  gate1510(.a(gate283inter10), .b(gate283inter9), .O(gate283inter11));
  nor2  gate1511(.a(gate283inter11), .b(gate283inter6), .O(gate283inter12));
  nand2 gate1512(.a(gate283inter12), .b(gate283inter1), .O(G828));
nand2 gate284( .a(G785), .b(G809), .O(G829) );
nand2 gate285( .a(G660), .b(G812), .O(G830) );
nand2 gate286( .a(G788), .b(G812), .O(G831) );

  xor2  gate939(.a(G815), .b(G663), .O(gate287inter0));
  nand2 gate940(.a(gate287inter0), .b(s_56), .O(gate287inter1));
  and2  gate941(.a(G815), .b(G663), .O(gate287inter2));
  inv1  gate942(.a(s_56), .O(gate287inter3));
  inv1  gate943(.a(s_57), .O(gate287inter4));
  nand2 gate944(.a(gate287inter4), .b(gate287inter3), .O(gate287inter5));
  nor2  gate945(.a(gate287inter5), .b(gate287inter2), .O(gate287inter6));
  inv1  gate946(.a(G663), .O(gate287inter7));
  inv1  gate947(.a(G815), .O(gate287inter8));
  nand2 gate948(.a(gate287inter8), .b(gate287inter7), .O(gate287inter9));
  nand2 gate949(.a(s_57), .b(gate287inter3), .O(gate287inter10));
  nor2  gate950(.a(gate287inter10), .b(gate287inter9), .O(gate287inter11));
  nor2  gate951(.a(gate287inter11), .b(gate287inter6), .O(gate287inter12));
  nand2 gate952(.a(gate287inter12), .b(gate287inter1), .O(G832));

  xor2  gate2129(.a(G815), .b(G791), .O(gate288inter0));
  nand2 gate2130(.a(gate288inter0), .b(s_226), .O(gate288inter1));
  and2  gate2131(.a(G815), .b(G791), .O(gate288inter2));
  inv1  gate2132(.a(s_226), .O(gate288inter3));
  inv1  gate2133(.a(s_227), .O(gate288inter4));
  nand2 gate2134(.a(gate288inter4), .b(gate288inter3), .O(gate288inter5));
  nor2  gate2135(.a(gate288inter5), .b(gate288inter2), .O(gate288inter6));
  inv1  gate2136(.a(G791), .O(gate288inter7));
  inv1  gate2137(.a(G815), .O(gate288inter8));
  nand2 gate2138(.a(gate288inter8), .b(gate288inter7), .O(gate288inter9));
  nand2 gate2139(.a(s_227), .b(gate288inter3), .O(gate288inter10));
  nor2  gate2140(.a(gate288inter10), .b(gate288inter9), .O(gate288inter11));
  nor2  gate2141(.a(gate288inter11), .b(gate288inter6), .O(gate288inter12));
  nand2 gate2142(.a(gate288inter12), .b(gate288inter1), .O(G833));

  xor2  gate561(.a(G819), .b(G818), .O(gate289inter0));
  nand2 gate562(.a(gate289inter0), .b(s_2), .O(gate289inter1));
  and2  gate563(.a(G819), .b(G818), .O(gate289inter2));
  inv1  gate564(.a(s_2), .O(gate289inter3));
  inv1  gate565(.a(s_3), .O(gate289inter4));
  nand2 gate566(.a(gate289inter4), .b(gate289inter3), .O(gate289inter5));
  nor2  gate567(.a(gate289inter5), .b(gate289inter2), .O(gate289inter6));
  inv1  gate568(.a(G818), .O(gate289inter7));
  inv1  gate569(.a(G819), .O(gate289inter8));
  nand2 gate570(.a(gate289inter8), .b(gate289inter7), .O(gate289inter9));
  nand2 gate571(.a(s_3), .b(gate289inter3), .O(gate289inter10));
  nor2  gate572(.a(gate289inter10), .b(gate289inter9), .O(gate289inter11));
  nor2  gate573(.a(gate289inter11), .b(gate289inter6), .O(gate289inter12));
  nand2 gate574(.a(gate289inter12), .b(gate289inter1), .O(G834));
nand2 gate290( .a(G820), .b(G821), .O(G847) );
nand2 gate291( .a(G822), .b(G823), .O(G860) );
nand2 gate292( .a(G824), .b(G825), .O(G873) );
nand2 gate293( .a(G828), .b(G829), .O(G886) );
nand2 gate294( .a(G832), .b(G833), .O(G899) );
nand2 gate295( .a(G830), .b(G831), .O(G912) );
nand2 gate296( .a(G826), .b(G827), .O(G925) );
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );
nand2 gate387( .a(G1), .b(G1036), .O(G1132) );
nand2 gate388( .a(G2), .b(G1039), .O(G1135) );
nand2 gate389( .a(G3), .b(G1042), .O(G1138) );
nand2 gate390( .a(G4), .b(G1045), .O(G1141) );

  xor2  gate1205(.a(G1048), .b(G5), .O(gate391inter0));
  nand2 gate1206(.a(gate391inter0), .b(s_94), .O(gate391inter1));
  and2  gate1207(.a(G1048), .b(G5), .O(gate391inter2));
  inv1  gate1208(.a(s_94), .O(gate391inter3));
  inv1  gate1209(.a(s_95), .O(gate391inter4));
  nand2 gate1210(.a(gate391inter4), .b(gate391inter3), .O(gate391inter5));
  nor2  gate1211(.a(gate391inter5), .b(gate391inter2), .O(gate391inter6));
  inv1  gate1212(.a(G5), .O(gate391inter7));
  inv1  gate1213(.a(G1048), .O(gate391inter8));
  nand2 gate1214(.a(gate391inter8), .b(gate391inter7), .O(gate391inter9));
  nand2 gate1215(.a(s_95), .b(gate391inter3), .O(gate391inter10));
  nor2  gate1216(.a(gate391inter10), .b(gate391inter9), .O(gate391inter11));
  nor2  gate1217(.a(gate391inter11), .b(gate391inter6), .O(gate391inter12));
  nand2 gate1218(.a(gate391inter12), .b(gate391inter1), .O(G1144));

  xor2  gate1681(.a(G1051), .b(G6), .O(gate392inter0));
  nand2 gate1682(.a(gate392inter0), .b(s_162), .O(gate392inter1));
  and2  gate1683(.a(G1051), .b(G6), .O(gate392inter2));
  inv1  gate1684(.a(s_162), .O(gate392inter3));
  inv1  gate1685(.a(s_163), .O(gate392inter4));
  nand2 gate1686(.a(gate392inter4), .b(gate392inter3), .O(gate392inter5));
  nor2  gate1687(.a(gate392inter5), .b(gate392inter2), .O(gate392inter6));
  inv1  gate1688(.a(G6), .O(gate392inter7));
  inv1  gate1689(.a(G1051), .O(gate392inter8));
  nand2 gate1690(.a(gate392inter8), .b(gate392inter7), .O(gate392inter9));
  nand2 gate1691(.a(s_163), .b(gate392inter3), .O(gate392inter10));
  nor2  gate1692(.a(gate392inter10), .b(gate392inter9), .O(gate392inter11));
  nor2  gate1693(.a(gate392inter11), .b(gate392inter6), .O(gate392inter12));
  nand2 gate1694(.a(gate392inter12), .b(gate392inter1), .O(G1147));
nand2 gate393( .a(G7), .b(G1054), .O(G1150) );

  xor2  gate2227(.a(G1057), .b(G8), .O(gate394inter0));
  nand2 gate2228(.a(gate394inter0), .b(s_240), .O(gate394inter1));
  and2  gate2229(.a(G1057), .b(G8), .O(gate394inter2));
  inv1  gate2230(.a(s_240), .O(gate394inter3));
  inv1  gate2231(.a(s_241), .O(gate394inter4));
  nand2 gate2232(.a(gate394inter4), .b(gate394inter3), .O(gate394inter5));
  nor2  gate2233(.a(gate394inter5), .b(gate394inter2), .O(gate394inter6));
  inv1  gate2234(.a(G8), .O(gate394inter7));
  inv1  gate2235(.a(G1057), .O(gate394inter8));
  nand2 gate2236(.a(gate394inter8), .b(gate394inter7), .O(gate394inter9));
  nand2 gate2237(.a(s_241), .b(gate394inter3), .O(gate394inter10));
  nor2  gate2238(.a(gate394inter10), .b(gate394inter9), .O(gate394inter11));
  nor2  gate2239(.a(gate394inter11), .b(gate394inter6), .O(gate394inter12));
  nand2 gate2240(.a(gate394inter12), .b(gate394inter1), .O(G1153));
nand2 gate395( .a(G9), .b(G1060), .O(G1156) );

  xor2  gate2073(.a(G1063), .b(G10), .O(gate396inter0));
  nand2 gate2074(.a(gate396inter0), .b(s_218), .O(gate396inter1));
  and2  gate2075(.a(G1063), .b(G10), .O(gate396inter2));
  inv1  gate2076(.a(s_218), .O(gate396inter3));
  inv1  gate2077(.a(s_219), .O(gate396inter4));
  nand2 gate2078(.a(gate396inter4), .b(gate396inter3), .O(gate396inter5));
  nor2  gate2079(.a(gate396inter5), .b(gate396inter2), .O(gate396inter6));
  inv1  gate2080(.a(G10), .O(gate396inter7));
  inv1  gate2081(.a(G1063), .O(gate396inter8));
  nand2 gate2082(.a(gate396inter8), .b(gate396inter7), .O(gate396inter9));
  nand2 gate2083(.a(s_219), .b(gate396inter3), .O(gate396inter10));
  nor2  gate2084(.a(gate396inter10), .b(gate396inter9), .O(gate396inter11));
  nor2  gate2085(.a(gate396inter11), .b(gate396inter6), .O(gate396inter12));
  nand2 gate2086(.a(gate396inter12), .b(gate396inter1), .O(G1159));

  xor2  gate1261(.a(G1066), .b(G11), .O(gate397inter0));
  nand2 gate1262(.a(gate397inter0), .b(s_102), .O(gate397inter1));
  and2  gate1263(.a(G1066), .b(G11), .O(gate397inter2));
  inv1  gate1264(.a(s_102), .O(gate397inter3));
  inv1  gate1265(.a(s_103), .O(gate397inter4));
  nand2 gate1266(.a(gate397inter4), .b(gate397inter3), .O(gate397inter5));
  nor2  gate1267(.a(gate397inter5), .b(gate397inter2), .O(gate397inter6));
  inv1  gate1268(.a(G11), .O(gate397inter7));
  inv1  gate1269(.a(G1066), .O(gate397inter8));
  nand2 gate1270(.a(gate397inter8), .b(gate397inter7), .O(gate397inter9));
  nand2 gate1271(.a(s_103), .b(gate397inter3), .O(gate397inter10));
  nor2  gate1272(.a(gate397inter10), .b(gate397inter9), .O(gate397inter11));
  nor2  gate1273(.a(gate397inter11), .b(gate397inter6), .O(gate397inter12));
  nand2 gate1274(.a(gate397inter12), .b(gate397inter1), .O(G1162));
nand2 gate398( .a(G12), .b(G1069), .O(G1165) );
nand2 gate399( .a(G13), .b(G1072), .O(G1168) );

  xor2  gate1933(.a(G1075), .b(G14), .O(gate400inter0));
  nand2 gate1934(.a(gate400inter0), .b(s_198), .O(gate400inter1));
  and2  gate1935(.a(G1075), .b(G14), .O(gate400inter2));
  inv1  gate1936(.a(s_198), .O(gate400inter3));
  inv1  gate1937(.a(s_199), .O(gate400inter4));
  nand2 gate1938(.a(gate400inter4), .b(gate400inter3), .O(gate400inter5));
  nor2  gate1939(.a(gate400inter5), .b(gate400inter2), .O(gate400inter6));
  inv1  gate1940(.a(G14), .O(gate400inter7));
  inv1  gate1941(.a(G1075), .O(gate400inter8));
  nand2 gate1942(.a(gate400inter8), .b(gate400inter7), .O(gate400inter9));
  nand2 gate1943(.a(s_199), .b(gate400inter3), .O(gate400inter10));
  nor2  gate1944(.a(gate400inter10), .b(gate400inter9), .O(gate400inter11));
  nor2  gate1945(.a(gate400inter11), .b(gate400inter6), .O(gate400inter12));
  nand2 gate1946(.a(gate400inter12), .b(gate400inter1), .O(G1171));
nand2 gate401( .a(G15), .b(G1078), .O(G1174) );
nand2 gate402( .a(G16), .b(G1081), .O(G1177) );

  xor2  gate1513(.a(G1084), .b(G17), .O(gate403inter0));
  nand2 gate1514(.a(gate403inter0), .b(s_138), .O(gate403inter1));
  and2  gate1515(.a(G1084), .b(G17), .O(gate403inter2));
  inv1  gate1516(.a(s_138), .O(gate403inter3));
  inv1  gate1517(.a(s_139), .O(gate403inter4));
  nand2 gate1518(.a(gate403inter4), .b(gate403inter3), .O(gate403inter5));
  nor2  gate1519(.a(gate403inter5), .b(gate403inter2), .O(gate403inter6));
  inv1  gate1520(.a(G17), .O(gate403inter7));
  inv1  gate1521(.a(G1084), .O(gate403inter8));
  nand2 gate1522(.a(gate403inter8), .b(gate403inter7), .O(gate403inter9));
  nand2 gate1523(.a(s_139), .b(gate403inter3), .O(gate403inter10));
  nor2  gate1524(.a(gate403inter10), .b(gate403inter9), .O(gate403inter11));
  nor2  gate1525(.a(gate403inter11), .b(gate403inter6), .O(gate403inter12));
  nand2 gate1526(.a(gate403inter12), .b(gate403inter1), .O(G1180));
nand2 gate404( .a(G18), .b(G1087), .O(G1183) );
nand2 gate405( .a(G19), .b(G1090), .O(G1186) );
nand2 gate406( .a(G20), .b(G1093), .O(G1189) );

  xor2  gate1037(.a(G1096), .b(G21), .O(gate407inter0));
  nand2 gate1038(.a(gate407inter0), .b(s_70), .O(gate407inter1));
  and2  gate1039(.a(G1096), .b(G21), .O(gate407inter2));
  inv1  gate1040(.a(s_70), .O(gate407inter3));
  inv1  gate1041(.a(s_71), .O(gate407inter4));
  nand2 gate1042(.a(gate407inter4), .b(gate407inter3), .O(gate407inter5));
  nor2  gate1043(.a(gate407inter5), .b(gate407inter2), .O(gate407inter6));
  inv1  gate1044(.a(G21), .O(gate407inter7));
  inv1  gate1045(.a(G1096), .O(gate407inter8));
  nand2 gate1046(.a(gate407inter8), .b(gate407inter7), .O(gate407inter9));
  nand2 gate1047(.a(s_71), .b(gate407inter3), .O(gate407inter10));
  nor2  gate1048(.a(gate407inter10), .b(gate407inter9), .O(gate407inter11));
  nor2  gate1049(.a(gate407inter11), .b(gate407inter6), .O(gate407inter12));
  nand2 gate1050(.a(gate407inter12), .b(gate407inter1), .O(G1192));
nand2 gate408( .a(G22), .b(G1099), .O(G1195) );
nand2 gate409( .a(G23), .b(G1102), .O(G1198) );

  xor2  gate855(.a(G1105), .b(G24), .O(gate410inter0));
  nand2 gate856(.a(gate410inter0), .b(s_44), .O(gate410inter1));
  and2  gate857(.a(G1105), .b(G24), .O(gate410inter2));
  inv1  gate858(.a(s_44), .O(gate410inter3));
  inv1  gate859(.a(s_45), .O(gate410inter4));
  nand2 gate860(.a(gate410inter4), .b(gate410inter3), .O(gate410inter5));
  nor2  gate861(.a(gate410inter5), .b(gate410inter2), .O(gate410inter6));
  inv1  gate862(.a(G24), .O(gate410inter7));
  inv1  gate863(.a(G1105), .O(gate410inter8));
  nand2 gate864(.a(gate410inter8), .b(gate410inter7), .O(gate410inter9));
  nand2 gate865(.a(s_45), .b(gate410inter3), .O(gate410inter10));
  nor2  gate866(.a(gate410inter10), .b(gate410inter9), .O(gate410inter11));
  nor2  gate867(.a(gate410inter11), .b(gate410inter6), .O(gate410inter12));
  nand2 gate868(.a(gate410inter12), .b(gate410inter1), .O(G1201));
nand2 gate411( .a(G25), .b(G1108), .O(G1204) );
nand2 gate412( .a(G26), .b(G1111), .O(G1207) );

  xor2  gate1149(.a(G1114), .b(G27), .O(gate413inter0));
  nand2 gate1150(.a(gate413inter0), .b(s_86), .O(gate413inter1));
  and2  gate1151(.a(G1114), .b(G27), .O(gate413inter2));
  inv1  gate1152(.a(s_86), .O(gate413inter3));
  inv1  gate1153(.a(s_87), .O(gate413inter4));
  nand2 gate1154(.a(gate413inter4), .b(gate413inter3), .O(gate413inter5));
  nor2  gate1155(.a(gate413inter5), .b(gate413inter2), .O(gate413inter6));
  inv1  gate1156(.a(G27), .O(gate413inter7));
  inv1  gate1157(.a(G1114), .O(gate413inter8));
  nand2 gate1158(.a(gate413inter8), .b(gate413inter7), .O(gate413inter9));
  nand2 gate1159(.a(s_87), .b(gate413inter3), .O(gate413inter10));
  nor2  gate1160(.a(gate413inter10), .b(gate413inter9), .O(gate413inter11));
  nor2  gate1161(.a(gate413inter11), .b(gate413inter6), .O(gate413inter12));
  nand2 gate1162(.a(gate413inter12), .b(gate413inter1), .O(G1210));

  xor2  gate1247(.a(G1117), .b(G28), .O(gate414inter0));
  nand2 gate1248(.a(gate414inter0), .b(s_100), .O(gate414inter1));
  and2  gate1249(.a(G1117), .b(G28), .O(gate414inter2));
  inv1  gate1250(.a(s_100), .O(gate414inter3));
  inv1  gate1251(.a(s_101), .O(gate414inter4));
  nand2 gate1252(.a(gate414inter4), .b(gate414inter3), .O(gate414inter5));
  nor2  gate1253(.a(gate414inter5), .b(gate414inter2), .O(gate414inter6));
  inv1  gate1254(.a(G28), .O(gate414inter7));
  inv1  gate1255(.a(G1117), .O(gate414inter8));
  nand2 gate1256(.a(gate414inter8), .b(gate414inter7), .O(gate414inter9));
  nand2 gate1257(.a(s_101), .b(gate414inter3), .O(gate414inter10));
  nor2  gate1258(.a(gate414inter10), .b(gate414inter9), .O(gate414inter11));
  nor2  gate1259(.a(gate414inter11), .b(gate414inter6), .O(gate414inter12));
  nand2 gate1260(.a(gate414inter12), .b(gate414inter1), .O(G1213));

  xor2  gate2157(.a(G1120), .b(G29), .O(gate415inter0));
  nand2 gate2158(.a(gate415inter0), .b(s_230), .O(gate415inter1));
  and2  gate2159(.a(G1120), .b(G29), .O(gate415inter2));
  inv1  gate2160(.a(s_230), .O(gate415inter3));
  inv1  gate2161(.a(s_231), .O(gate415inter4));
  nand2 gate2162(.a(gate415inter4), .b(gate415inter3), .O(gate415inter5));
  nor2  gate2163(.a(gate415inter5), .b(gate415inter2), .O(gate415inter6));
  inv1  gate2164(.a(G29), .O(gate415inter7));
  inv1  gate2165(.a(G1120), .O(gate415inter8));
  nand2 gate2166(.a(gate415inter8), .b(gate415inter7), .O(gate415inter9));
  nand2 gate2167(.a(s_231), .b(gate415inter3), .O(gate415inter10));
  nor2  gate2168(.a(gate415inter10), .b(gate415inter9), .O(gate415inter11));
  nor2  gate2169(.a(gate415inter11), .b(gate415inter6), .O(gate415inter12));
  nand2 gate2170(.a(gate415inter12), .b(gate415inter1), .O(G1216));
nand2 gate416( .a(G30), .b(G1123), .O(G1219) );
nand2 gate417( .a(G31), .b(G1126), .O(G1222) );
nand2 gate418( .a(G32), .b(G1129), .O(G1225) );
nand2 gate419( .a(G1), .b(G1132), .O(G1228) );
nand2 gate420( .a(G1036), .b(G1132), .O(G1229) );
nand2 gate421( .a(G2), .b(G1135), .O(G1230) );
nand2 gate422( .a(G1039), .b(G1135), .O(G1231) );
nand2 gate423( .a(G3), .b(G1138), .O(G1232) );
nand2 gate424( .a(G1042), .b(G1138), .O(G1233) );

  xor2  gate1471(.a(G1141), .b(G4), .O(gate425inter0));
  nand2 gate1472(.a(gate425inter0), .b(s_132), .O(gate425inter1));
  and2  gate1473(.a(G1141), .b(G4), .O(gate425inter2));
  inv1  gate1474(.a(s_132), .O(gate425inter3));
  inv1  gate1475(.a(s_133), .O(gate425inter4));
  nand2 gate1476(.a(gate425inter4), .b(gate425inter3), .O(gate425inter5));
  nor2  gate1477(.a(gate425inter5), .b(gate425inter2), .O(gate425inter6));
  inv1  gate1478(.a(G4), .O(gate425inter7));
  inv1  gate1479(.a(G1141), .O(gate425inter8));
  nand2 gate1480(.a(gate425inter8), .b(gate425inter7), .O(gate425inter9));
  nand2 gate1481(.a(s_133), .b(gate425inter3), .O(gate425inter10));
  nor2  gate1482(.a(gate425inter10), .b(gate425inter9), .O(gate425inter11));
  nor2  gate1483(.a(gate425inter11), .b(gate425inter6), .O(gate425inter12));
  nand2 gate1484(.a(gate425inter12), .b(gate425inter1), .O(G1234));
nand2 gate426( .a(G1045), .b(G1141), .O(G1235) );
nand2 gate427( .a(G5), .b(G1144), .O(G1236) );
nand2 gate428( .a(G1048), .b(G1144), .O(G1237) );
nand2 gate429( .a(G6), .b(G1147), .O(G1238) );
nand2 gate430( .a(G1051), .b(G1147), .O(G1239) );

  xor2  gate2017(.a(G1150), .b(G7), .O(gate431inter0));
  nand2 gate2018(.a(gate431inter0), .b(s_210), .O(gate431inter1));
  and2  gate2019(.a(G1150), .b(G7), .O(gate431inter2));
  inv1  gate2020(.a(s_210), .O(gate431inter3));
  inv1  gate2021(.a(s_211), .O(gate431inter4));
  nand2 gate2022(.a(gate431inter4), .b(gate431inter3), .O(gate431inter5));
  nor2  gate2023(.a(gate431inter5), .b(gate431inter2), .O(gate431inter6));
  inv1  gate2024(.a(G7), .O(gate431inter7));
  inv1  gate2025(.a(G1150), .O(gate431inter8));
  nand2 gate2026(.a(gate431inter8), .b(gate431inter7), .O(gate431inter9));
  nand2 gate2027(.a(s_211), .b(gate431inter3), .O(gate431inter10));
  nor2  gate2028(.a(gate431inter10), .b(gate431inter9), .O(gate431inter11));
  nor2  gate2029(.a(gate431inter11), .b(gate431inter6), .O(gate431inter12));
  nand2 gate2030(.a(gate431inter12), .b(gate431inter1), .O(G1240));
nand2 gate432( .a(G1054), .b(G1150), .O(G1241) );
nand2 gate433( .a(G8), .b(G1153), .O(G1242) );

  xor2  gate2171(.a(G1153), .b(G1057), .O(gate434inter0));
  nand2 gate2172(.a(gate434inter0), .b(s_232), .O(gate434inter1));
  and2  gate2173(.a(G1153), .b(G1057), .O(gate434inter2));
  inv1  gate2174(.a(s_232), .O(gate434inter3));
  inv1  gate2175(.a(s_233), .O(gate434inter4));
  nand2 gate2176(.a(gate434inter4), .b(gate434inter3), .O(gate434inter5));
  nor2  gate2177(.a(gate434inter5), .b(gate434inter2), .O(gate434inter6));
  inv1  gate2178(.a(G1057), .O(gate434inter7));
  inv1  gate2179(.a(G1153), .O(gate434inter8));
  nand2 gate2180(.a(gate434inter8), .b(gate434inter7), .O(gate434inter9));
  nand2 gate2181(.a(s_233), .b(gate434inter3), .O(gate434inter10));
  nor2  gate2182(.a(gate434inter10), .b(gate434inter9), .O(gate434inter11));
  nor2  gate2183(.a(gate434inter11), .b(gate434inter6), .O(gate434inter12));
  nand2 gate2184(.a(gate434inter12), .b(gate434inter1), .O(G1243));

  xor2  gate1275(.a(G1156), .b(G9), .O(gate435inter0));
  nand2 gate1276(.a(gate435inter0), .b(s_104), .O(gate435inter1));
  and2  gate1277(.a(G1156), .b(G9), .O(gate435inter2));
  inv1  gate1278(.a(s_104), .O(gate435inter3));
  inv1  gate1279(.a(s_105), .O(gate435inter4));
  nand2 gate1280(.a(gate435inter4), .b(gate435inter3), .O(gate435inter5));
  nor2  gate1281(.a(gate435inter5), .b(gate435inter2), .O(gate435inter6));
  inv1  gate1282(.a(G9), .O(gate435inter7));
  inv1  gate1283(.a(G1156), .O(gate435inter8));
  nand2 gate1284(.a(gate435inter8), .b(gate435inter7), .O(gate435inter9));
  nand2 gate1285(.a(s_105), .b(gate435inter3), .O(gate435inter10));
  nor2  gate1286(.a(gate435inter10), .b(gate435inter9), .O(gate435inter11));
  nor2  gate1287(.a(gate435inter11), .b(gate435inter6), .O(gate435inter12));
  nand2 gate1288(.a(gate435inter12), .b(gate435inter1), .O(G1244));
nand2 gate436( .a(G1060), .b(G1156), .O(G1245) );
nand2 gate437( .a(G10), .b(G1159), .O(G1246) );
nand2 gate438( .a(G1063), .b(G1159), .O(G1247) );

  xor2  gate631(.a(G1162), .b(G11), .O(gate439inter0));
  nand2 gate632(.a(gate439inter0), .b(s_12), .O(gate439inter1));
  and2  gate633(.a(G1162), .b(G11), .O(gate439inter2));
  inv1  gate634(.a(s_12), .O(gate439inter3));
  inv1  gate635(.a(s_13), .O(gate439inter4));
  nand2 gate636(.a(gate439inter4), .b(gate439inter3), .O(gate439inter5));
  nor2  gate637(.a(gate439inter5), .b(gate439inter2), .O(gate439inter6));
  inv1  gate638(.a(G11), .O(gate439inter7));
  inv1  gate639(.a(G1162), .O(gate439inter8));
  nand2 gate640(.a(gate439inter8), .b(gate439inter7), .O(gate439inter9));
  nand2 gate641(.a(s_13), .b(gate439inter3), .O(gate439inter10));
  nor2  gate642(.a(gate439inter10), .b(gate439inter9), .O(gate439inter11));
  nor2  gate643(.a(gate439inter11), .b(gate439inter6), .O(gate439inter12));
  nand2 gate644(.a(gate439inter12), .b(gate439inter1), .O(G1248));
nand2 gate440( .a(G1066), .b(G1162), .O(G1249) );

  xor2  gate1905(.a(G1165), .b(G12), .O(gate441inter0));
  nand2 gate1906(.a(gate441inter0), .b(s_194), .O(gate441inter1));
  and2  gate1907(.a(G1165), .b(G12), .O(gate441inter2));
  inv1  gate1908(.a(s_194), .O(gate441inter3));
  inv1  gate1909(.a(s_195), .O(gate441inter4));
  nand2 gate1910(.a(gate441inter4), .b(gate441inter3), .O(gate441inter5));
  nor2  gate1911(.a(gate441inter5), .b(gate441inter2), .O(gate441inter6));
  inv1  gate1912(.a(G12), .O(gate441inter7));
  inv1  gate1913(.a(G1165), .O(gate441inter8));
  nand2 gate1914(.a(gate441inter8), .b(gate441inter7), .O(gate441inter9));
  nand2 gate1915(.a(s_195), .b(gate441inter3), .O(gate441inter10));
  nor2  gate1916(.a(gate441inter10), .b(gate441inter9), .O(gate441inter11));
  nor2  gate1917(.a(gate441inter11), .b(gate441inter6), .O(gate441inter12));
  nand2 gate1918(.a(gate441inter12), .b(gate441inter1), .O(G1250));

  xor2  gate1639(.a(G1165), .b(G1069), .O(gate442inter0));
  nand2 gate1640(.a(gate442inter0), .b(s_156), .O(gate442inter1));
  and2  gate1641(.a(G1165), .b(G1069), .O(gate442inter2));
  inv1  gate1642(.a(s_156), .O(gate442inter3));
  inv1  gate1643(.a(s_157), .O(gate442inter4));
  nand2 gate1644(.a(gate442inter4), .b(gate442inter3), .O(gate442inter5));
  nor2  gate1645(.a(gate442inter5), .b(gate442inter2), .O(gate442inter6));
  inv1  gate1646(.a(G1069), .O(gate442inter7));
  inv1  gate1647(.a(G1165), .O(gate442inter8));
  nand2 gate1648(.a(gate442inter8), .b(gate442inter7), .O(gate442inter9));
  nand2 gate1649(.a(s_157), .b(gate442inter3), .O(gate442inter10));
  nor2  gate1650(.a(gate442inter10), .b(gate442inter9), .O(gate442inter11));
  nor2  gate1651(.a(gate442inter11), .b(gate442inter6), .O(gate442inter12));
  nand2 gate1652(.a(gate442inter12), .b(gate442inter1), .O(G1251));

  xor2  gate799(.a(G1168), .b(G13), .O(gate443inter0));
  nand2 gate800(.a(gate443inter0), .b(s_36), .O(gate443inter1));
  and2  gate801(.a(G1168), .b(G13), .O(gate443inter2));
  inv1  gate802(.a(s_36), .O(gate443inter3));
  inv1  gate803(.a(s_37), .O(gate443inter4));
  nand2 gate804(.a(gate443inter4), .b(gate443inter3), .O(gate443inter5));
  nor2  gate805(.a(gate443inter5), .b(gate443inter2), .O(gate443inter6));
  inv1  gate806(.a(G13), .O(gate443inter7));
  inv1  gate807(.a(G1168), .O(gate443inter8));
  nand2 gate808(.a(gate443inter8), .b(gate443inter7), .O(gate443inter9));
  nand2 gate809(.a(s_37), .b(gate443inter3), .O(gate443inter10));
  nor2  gate810(.a(gate443inter10), .b(gate443inter9), .O(gate443inter11));
  nor2  gate811(.a(gate443inter11), .b(gate443inter6), .O(gate443inter12));
  nand2 gate812(.a(gate443inter12), .b(gate443inter1), .O(G1252));

  xor2  gate785(.a(G1168), .b(G1072), .O(gate444inter0));
  nand2 gate786(.a(gate444inter0), .b(s_34), .O(gate444inter1));
  and2  gate787(.a(G1168), .b(G1072), .O(gate444inter2));
  inv1  gate788(.a(s_34), .O(gate444inter3));
  inv1  gate789(.a(s_35), .O(gate444inter4));
  nand2 gate790(.a(gate444inter4), .b(gate444inter3), .O(gate444inter5));
  nor2  gate791(.a(gate444inter5), .b(gate444inter2), .O(gate444inter6));
  inv1  gate792(.a(G1072), .O(gate444inter7));
  inv1  gate793(.a(G1168), .O(gate444inter8));
  nand2 gate794(.a(gate444inter8), .b(gate444inter7), .O(gate444inter9));
  nand2 gate795(.a(s_35), .b(gate444inter3), .O(gate444inter10));
  nor2  gate796(.a(gate444inter10), .b(gate444inter9), .O(gate444inter11));
  nor2  gate797(.a(gate444inter11), .b(gate444inter6), .O(gate444inter12));
  nand2 gate798(.a(gate444inter12), .b(gate444inter1), .O(G1253));
nand2 gate445( .a(G14), .b(G1171), .O(G1254) );

  xor2  gate2185(.a(G1171), .b(G1075), .O(gate446inter0));
  nand2 gate2186(.a(gate446inter0), .b(s_234), .O(gate446inter1));
  and2  gate2187(.a(G1171), .b(G1075), .O(gate446inter2));
  inv1  gate2188(.a(s_234), .O(gate446inter3));
  inv1  gate2189(.a(s_235), .O(gate446inter4));
  nand2 gate2190(.a(gate446inter4), .b(gate446inter3), .O(gate446inter5));
  nor2  gate2191(.a(gate446inter5), .b(gate446inter2), .O(gate446inter6));
  inv1  gate2192(.a(G1075), .O(gate446inter7));
  inv1  gate2193(.a(G1171), .O(gate446inter8));
  nand2 gate2194(.a(gate446inter8), .b(gate446inter7), .O(gate446inter9));
  nand2 gate2195(.a(s_235), .b(gate446inter3), .O(gate446inter10));
  nor2  gate2196(.a(gate446inter10), .b(gate446inter9), .O(gate446inter11));
  nor2  gate2197(.a(gate446inter11), .b(gate446inter6), .O(gate446inter12));
  nand2 gate2198(.a(gate446inter12), .b(gate446inter1), .O(G1255));
nand2 gate447( .a(G15), .b(G1174), .O(G1256) );
nand2 gate448( .a(G1078), .b(G1174), .O(G1257) );
nand2 gate449( .a(G16), .b(G1177), .O(G1258) );
nand2 gate450( .a(G1081), .b(G1177), .O(G1259) );
nand2 gate451( .a(G17), .b(G1180), .O(G1260) );
nand2 gate452( .a(G1084), .b(G1180), .O(G1261) );

  xor2  gate673(.a(G1183), .b(G18), .O(gate453inter0));
  nand2 gate674(.a(gate453inter0), .b(s_18), .O(gate453inter1));
  and2  gate675(.a(G1183), .b(G18), .O(gate453inter2));
  inv1  gate676(.a(s_18), .O(gate453inter3));
  inv1  gate677(.a(s_19), .O(gate453inter4));
  nand2 gate678(.a(gate453inter4), .b(gate453inter3), .O(gate453inter5));
  nor2  gate679(.a(gate453inter5), .b(gate453inter2), .O(gate453inter6));
  inv1  gate680(.a(G18), .O(gate453inter7));
  inv1  gate681(.a(G1183), .O(gate453inter8));
  nand2 gate682(.a(gate453inter8), .b(gate453inter7), .O(gate453inter9));
  nand2 gate683(.a(s_19), .b(gate453inter3), .O(gate453inter10));
  nor2  gate684(.a(gate453inter10), .b(gate453inter9), .O(gate453inter11));
  nor2  gate685(.a(gate453inter11), .b(gate453inter6), .O(gate453inter12));
  nand2 gate686(.a(gate453inter12), .b(gate453inter1), .O(G1262));

  xor2  gate2031(.a(G1183), .b(G1087), .O(gate454inter0));
  nand2 gate2032(.a(gate454inter0), .b(s_212), .O(gate454inter1));
  and2  gate2033(.a(G1183), .b(G1087), .O(gate454inter2));
  inv1  gate2034(.a(s_212), .O(gate454inter3));
  inv1  gate2035(.a(s_213), .O(gate454inter4));
  nand2 gate2036(.a(gate454inter4), .b(gate454inter3), .O(gate454inter5));
  nor2  gate2037(.a(gate454inter5), .b(gate454inter2), .O(gate454inter6));
  inv1  gate2038(.a(G1087), .O(gate454inter7));
  inv1  gate2039(.a(G1183), .O(gate454inter8));
  nand2 gate2040(.a(gate454inter8), .b(gate454inter7), .O(gate454inter9));
  nand2 gate2041(.a(s_213), .b(gate454inter3), .O(gate454inter10));
  nor2  gate2042(.a(gate454inter10), .b(gate454inter9), .O(gate454inter11));
  nor2  gate2043(.a(gate454inter11), .b(gate454inter6), .O(gate454inter12));
  nand2 gate2044(.a(gate454inter12), .b(gate454inter1), .O(G1263));
nand2 gate455( .a(G19), .b(G1186), .O(G1264) );
nand2 gate456( .a(G1090), .b(G1186), .O(G1265) );
nand2 gate457( .a(G20), .b(G1189), .O(G1266) );
nand2 gate458( .a(G1093), .b(G1189), .O(G1267) );

  xor2  gate2045(.a(G1192), .b(G21), .O(gate459inter0));
  nand2 gate2046(.a(gate459inter0), .b(s_214), .O(gate459inter1));
  and2  gate2047(.a(G1192), .b(G21), .O(gate459inter2));
  inv1  gate2048(.a(s_214), .O(gate459inter3));
  inv1  gate2049(.a(s_215), .O(gate459inter4));
  nand2 gate2050(.a(gate459inter4), .b(gate459inter3), .O(gate459inter5));
  nor2  gate2051(.a(gate459inter5), .b(gate459inter2), .O(gate459inter6));
  inv1  gate2052(.a(G21), .O(gate459inter7));
  inv1  gate2053(.a(G1192), .O(gate459inter8));
  nand2 gate2054(.a(gate459inter8), .b(gate459inter7), .O(gate459inter9));
  nand2 gate2055(.a(s_215), .b(gate459inter3), .O(gate459inter10));
  nor2  gate2056(.a(gate459inter10), .b(gate459inter9), .O(gate459inter11));
  nor2  gate2057(.a(gate459inter11), .b(gate459inter6), .O(gate459inter12));
  nand2 gate2058(.a(gate459inter12), .b(gate459inter1), .O(G1268));
nand2 gate460( .a(G1096), .b(G1192), .O(G1269) );
nand2 gate461( .a(G22), .b(G1195), .O(G1270) );
nand2 gate462( .a(G1099), .b(G1195), .O(G1271) );
nand2 gate463( .a(G23), .b(G1198), .O(G1272) );
nand2 gate464( .a(G1102), .b(G1198), .O(G1273) );

  xor2  gate1485(.a(G1201), .b(G24), .O(gate465inter0));
  nand2 gate1486(.a(gate465inter0), .b(s_134), .O(gate465inter1));
  and2  gate1487(.a(G1201), .b(G24), .O(gate465inter2));
  inv1  gate1488(.a(s_134), .O(gate465inter3));
  inv1  gate1489(.a(s_135), .O(gate465inter4));
  nand2 gate1490(.a(gate465inter4), .b(gate465inter3), .O(gate465inter5));
  nor2  gate1491(.a(gate465inter5), .b(gate465inter2), .O(gate465inter6));
  inv1  gate1492(.a(G24), .O(gate465inter7));
  inv1  gate1493(.a(G1201), .O(gate465inter8));
  nand2 gate1494(.a(gate465inter8), .b(gate465inter7), .O(gate465inter9));
  nand2 gate1495(.a(s_135), .b(gate465inter3), .O(gate465inter10));
  nor2  gate1496(.a(gate465inter10), .b(gate465inter9), .O(gate465inter11));
  nor2  gate1497(.a(gate465inter11), .b(gate465inter6), .O(gate465inter12));
  nand2 gate1498(.a(gate465inter12), .b(gate465inter1), .O(G1274));
nand2 gate466( .a(G1105), .b(G1201), .O(G1275) );
nand2 gate467( .a(G25), .b(G1204), .O(G1276) );
nand2 gate468( .a(G1108), .b(G1204), .O(G1277) );

  xor2  gate1387(.a(G1207), .b(G26), .O(gate469inter0));
  nand2 gate1388(.a(gate469inter0), .b(s_120), .O(gate469inter1));
  and2  gate1389(.a(G1207), .b(G26), .O(gate469inter2));
  inv1  gate1390(.a(s_120), .O(gate469inter3));
  inv1  gate1391(.a(s_121), .O(gate469inter4));
  nand2 gate1392(.a(gate469inter4), .b(gate469inter3), .O(gate469inter5));
  nor2  gate1393(.a(gate469inter5), .b(gate469inter2), .O(gate469inter6));
  inv1  gate1394(.a(G26), .O(gate469inter7));
  inv1  gate1395(.a(G1207), .O(gate469inter8));
  nand2 gate1396(.a(gate469inter8), .b(gate469inter7), .O(gate469inter9));
  nand2 gate1397(.a(s_121), .b(gate469inter3), .O(gate469inter10));
  nor2  gate1398(.a(gate469inter10), .b(gate469inter9), .O(gate469inter11));
  nor2  gate1399(.a(gate469inter11), .b(gate469inter6), .O(gate469inter12));
  nand2 gate1400(.a(gate469inter12), .b(gate469inter1), .O(G1278));
nand2 gate470( .a(G1111), .b(G1207), .O(G1279) );
nand2 gate471( .a(G27), .b(G1210), .O(G1280) );
nand2 gate472( .a(G1114), .b(G1210), .O(G1281) );
nand2 gate473( .a(G28), .b(G1213), .O(G1282) );

  xor2  gate659(.a(G1213), .b(G1117), .O(gate474inter0));
  nand2 gate660(.a(gate474inter0), .b(s_16), .O(gate474inter1));
  and2  gate661(.a(G1213), .b(G1117), .O(gate474inter2));
  inv1  gate662(.a(s_16), .O(gate474inter3));
  inv1  gate663(.a(s_17), .O(gate474inter4));
  nand2 gate664(.a(gate474inter4), .b(gate474inter3), .O(gate474inter5));
  nor2  gate665(.a(gate474inter5), .b(gate474inter2), .O(gate474inter6));
  inv1  gate666(.a(G1117), .O(gate474inter7));
  inv1  gate667(.a(G1213), .O(gate474inter8));
  nand2 gate668(.a(gate474inter8), .b(gate474inter7), .O(gate474inter9));
  nand2 gate669(.a(s_17), .b(gate474inter3), .O(gate474inter10));
  nor2  gate670(.a(gate474inter10), .b(gate474inter9), .O(gate474inter11));
  nor2  gate671(.a(gate474inter11), .b(gate474inter6), .O(gate474inter12));
  nand2 gate672(.a(gate474inter12), .b(gate474inter1), .O(G1283));
nand2 gate475( .a(G29), .b(G1216), .O(G1284) );
nand2 gate476( .a(G1120), .b(G1216), .O(G1285) );
nand2 gate477( .a(G30), .b(G1219), .O(G1286) );
nand2 gate478( .a(G1123), .b(G1219), .O(G1287) );
nand2 gate479( .a(G31), .b(G1222), .O(G1288) );

  xor2  gate1093(.a(G1222), .b(G1126), .O(gate480inter0));
  nand2 gate1094(.a(gate480inter0), .b(s_78), .O(gate480inter1));
  and2  gate1095(.a(G1222), .b(G1126), .O(gate480inter2));
  inv1  gate1096(.a(s_78), .O(gate480inter3));
  inv1  gate1097(.a(s_79), .O(gate480inter4));
  nand2 gate1098(.a(gate480inter4), .b(gate480inter3), .O(gate480inter5));
  nor2  gate1099(.a(gate480inter5), .b(gate480inter2), .O(gate480inter6));
  inv1  gate1100(.a(G1126), .O(gate480inter7));
  inv1  gate1101(.a(G1222), .O(gate480inter8));
  nand2 gate1102(.a(gate480inter8), .b(gate480inter7), .O(gate480inter9));
  nand2 gate1103(.a(s_79), .b(gate480inter3), .O(gate480inter10));
  nor2  gate1104(.a(gate480inter10), .b(gate480inter9), .O(gate480inter11));
  nor2  gate1105(.a(gate480inter11), .b(gate480inter6), .O(gate480inter12));
  nand2 gate1106(.a(gate480inter12), .b(gate480inter1), .O(G1289));
nand2 gate481( .a(G32), .b(G1225), .O(G1290) );
nand2 gate482( .a(G1129), .b(G1225), .O(G1291) );
nand2 gate483( .a(G1228), .b(G1229), .O(G1292) );
nand2 gate484( .a(G1230), .b(G1231), .O(G1293) );

  xor2  gate603(.a(G1233), .b(G1232), .O(gate485inter0));
  nand2 gate604(.a(gate485inter0), .b(s_8), .O(gate485inter1));
  and2  gate605(.a(G1233), .b(G1232), .O(gate485inter2));
  inv1  gate606(.a(s_8), .O(gate485inter3));
  inv1  gate607(.a(s_9), .O(gate485inter4));
  nand2 gate608(.a(gate485inter4), .b(gate485inter3), .O(gate485inter5));
  nor2  gate609(.a(gate485inter5), .b(gate485inter2), .O(gate485inter6));
  inv1  gate610(.a(G1232), .O(gate485inter7));
  inv1  gate611(.a(G1233), .O(gate485inter8));
  nand2 gate612(.a(gate485inter8), .b(gate485inter7), .O(gate485inter9));
  nand2 gate613(.a(s_9), .b(gate485inter3), .O(gate485inter10));
  nor2  gate614(.a(gate485inter10), .b(gate485inter9), .O(gate485inter11));
  nor2  gate615(.a(gate485inter11), .b(gate485inter6), .O(gate485inter12));
  nand2 gate616(.a(gate485inter12), .b(gate485inter1), .O(G1294));
nand2 gate486( .a(G1234), .b(G1235), .O(G1295) );

  xor2  gate1961(.a(G1237), .b(G1236), .O(gate487inter0));
  nand2 gate1962(.a(gate487inter0), .b(s_202), .O(gate487inter1));
  and2  gate1963(.a(G1237), .b(G1236), .O(gate487inter2));
  inv1  gate1964(.a(s_202), .O(gate487inter3));
  inv1  gate1965(.a(s_203), .O(gate487inter4));
  nand2 gate1966(.a(gate487inter4), .b(gate487inter3), .O(gate487inter5));
  nor2  gate1967(.a(gate487inter5), .b(gate487inter2), .O(gate487inter6));
  inv1  gate1968(.a(G1236), .O(gate487inter7));
  inv1  gate1969(.a(G1237), .O(gate487inter8));
  nand2 gate1970(.a(gate487inter8), .b(gate487inter7), .O(gate487inter9));
  nand2 gate1971(.a(s_203), .b(gate487inter3), .O(gate487inter10));
  nor2  gate1972(.a(gate487inter10), .b(gate487inter9), .O(gate487inter11));
  nor2  gate1973(.a(gate487inter11), .b(gate487inter6), .O(gate487inter12));
  nand2 gate1974(.a(gate487inter12), .b(gate487inter1), .O(G1296));

  xor2  gate1121(.a(G1239), .b(G1238), .O(gate488inter0));
  nand2 gate1122(.a(gate488inter0), .b(s_82), .O(gate488inter1));
  and2  gate1123(.a(G1239), .b(G1238), .O(gate488inter2));
  inv1  gate1124(.a(s_82), .O(gate488inter3));
  inv1  gate1125(.a(s_83), .O(gate488inter4));
  nand2 gate1126(.a(gate488inter4), .b(gate488inter3), .O(gate488inter5));
  nor2  gate1127(.a(gate488inter5), .b(gate488inter2), .O(gate488inter6));
  inv1  gate1128(.a(G1238), .O(gate488inter7));
  inv1  gate1129(.a(G1239), .O(gate488inter8));
  nand2 gate1130(.a(gate488inter8), .b(gate488inter7), .O(gate488inter9));
  nand2 gate1131(.a(s_83), .b(gate488inter3), .O(gate488inter10));
  nor2  gate1132(.a(gate488inter10), .b(gate488inter9), .O(gate488inter11));
  nor2  gate1133(.a(gate488inter11), .b(gate488inter6), .O(gate488inter12));
  nand2 gate1134(.a(gate488inter12), .b(gate488inter1), .O(G1297));

  xor2  gate1835(.a(G1241), .b(G1240), .O(gate489inter0));
  nand2 gate1836(.a(gate489inter0), .b(s_184), .O(gate489inter1));
  and2  gate1837(.a(G1241), .b(G1240), .O(gate489inter2));
  inv1  gate1838(.a(s_184), .O(gate489inter3));
  inv1  gate1839(.a(s_185), .O(gate489inter4));
  nand2 gate1840(.a(gate489inter4), .b(gate489inter3), .O(gate489inter5));
  nor2  gate1841(.a(gate489inter5), .b(gate489inter2), .O(gate489inter6));
  inv1  gate1842(.a(G1240), .O(gate489inter7));
  inv1  gate1843(.a(G1241), .O(gate489inter8));
  nand2 gate1844(.a(gate489inter8), .b(gate489inter7), .O(gate489inter9));
  nand2 gate1845(.a(s_185), .b(gate489inter3), .O(gate489inter10));
  nor2  gate1846(.a(gate489inter10), .b(gate489inter9), .O(gate489inter11));
  nor2  gate1847(.a(gate489inter11), .b(gate489inter6), .O(gate489inter12));
  nand2 gate1848(.a(gate489inter12), .b(gate489inter1), .O(G1298));
nand2 gate490( .a(G1242), .b(G1243), .O(G1299) );

  xor2  gate1863(.a(G1245), .b(G1244), .O(gate491inter0));
  nand2 gate1864(.a(gate491inter0), .b(s_188), .O(gate491inter1));
  and2  gate1865(.a(G1245), .b(G1244), .O(gate491inter2));
  inv1  gate1866(.a(s_188), .O(gate491inter3));
  inv1  gate1867(.a(s_189), .O(gate491inter4));
  nand2 gate1868(.a(gate491inter4), .b(gate491inter3), .O(gate491inter5));
  nor2  gate1869(.a(gate491inter5), .b(gate491inter2), .O(gate491inter6));
  inv1  gate1870(.a(G1244), .O(gate491inter7));
  inv1  gate1871(.a(G1245), .O(gate491inter8));
  nand2 gate1872(.a(gate491inter8), .b(gate491inter7), .O(gate491inter9));
  nand2 gate1873(.a(s_189), .b(gate491inter3), .O(gate491inter10));
  nor2  gate1874(.a(gate491inter10), .b(gate491inter9), .O(gate491inter11));
  nor2  gate1875(.a(gate491inter11), .b(gate491inter6), .O(gate491inter12));
  nand2 gate1876(.a(gate491inter12), .b(gate491inter1), .O(G1300));

  xor2  gate1765(.a(G1247), .b(G1246), .O(gate492inter0));
  nand2 gate1766(.a(gate492inter0), .b(s_174), .O(gate492inter1));
  and2  gate1767(.a(G1247), .b(G1246), .O(gate492inter2));
  inv1  gate1768(.a(s_174), .O(gate492inter3));
  inv1  gate1769(.a(s_175), .O(gate492inter4));
  nand2 gate1770(.a(gate492inter4), .b(gate492inter3), .O(gate492inter5));
  nor2  gate1771(.a(gate492inter5), .b(gate492inter2), .O(gate492inter6));
  inv1  gate1772(.a(G1246), .O(gate492inter7));
  inv1  gate1773(.a(G1247), .O(gate492inter8));
  nand2 gate1774(.a(gate492inter8), .b(gate492inter7), .O(gate492inter9));
  nand2 gate1775(.a(s_175), .b(gate492inter3), .O(gate492inter10));
  nor2  gate1776(.a(gate492inter10), .b(gate492inter9), .O(gate492inter11));
  nor2  gate1777(.a(gate492inter11), .b(gate492inter6), .O(gate492inter12));
  nand2 gate1778(.a(gate492inter12), .b(gate492inter1), .O(G1301));
nand2 gate493( .a(G1248), .b(G1249), .O(G1302) );
nand2 gate494( .a(G1250), .b(G1251), .O(G1303) );

  xor2  gate1345(.a(G1253), .b(G1252), .O(gate495inter0));
  nand2 gate1346(.a(gate495inter0), .b(s_114), .O(gate495inter1));
  and2  gate1347(.a(G1253), .b(G1252), .O(gate495inter2));
  inv1  gate1348(.a(s_114), .O(gate495inter3));
  inv1  gate1349(.a(s_115), .O(gate495inter4));
  nand2 gate1350(.a(gate495inter4), .b(gate495inter3), .O(gate495inter5));
  nor2  gate1351(.a(gate495inter5), .b(gate495inter2), .O(gate495inter6));
  inv1  gate1352(.a(G1252), .O(gate495inter7));
  inv1  gate1353(.a(G1253), .O(gate495inter8));
  nand2 gate1354(.a(gate495inter8), .b(gate495inter7), .O(gate495inter9));
  nand2 gate1355(.a(s_115), .b(gate495inter3), .O(gate495inter10));
  nor2  gate1356(.a(gate495inter10), .b(gate495inter9), .O(gate495inter11));
  nor2  gate1357(.a(gate495inter11), .b(gate495inter6), .O(gate495inter12));
  nand2 gate1358(.a(gate495inter12), .b(gate495inter1), .O(G1304));
nand2 gate496( .a(G1254), .b(G1255), .O(G1305) );
nand2 gate497( .a(G1256), .b(G1257), .O(G1306) );
nand2 gate498( .a(G1258), .b(G1259), .O(G1307) );
nand2 gate499( .a(G1260), .b(G1261), .O(G1308) );
nand2 gate500( .a(G1262), .b(G1263), .O(G1309) );

  xor2  gate1233(.a(G1265), .b(G1264), .O(gate501inter0));
  nand2 gate1234(.a(gate501inter0), .b(s_98), .O(gate501inter1));
  and2  gate1235(.a(G1265), .b(G1264), .O(gate501inter2));
  inv1  gate1236(.a(s_98), .O(gate501inter3));
  inv1  gate1237(.a(s_99), .O(gate501inter4));
  nand2 gate1238(.a(gate501inter4), .b(gate501inter3), .O(gate501inter5));
  nor2  gate1239(.a(gate501inter5), .b(gate501inter2), .O(gate501inter6));
  inv1  gate1240(.a(G1264), .O(gate501inter7));
  inv1  gate1241(.a(G1265), .O(gate501inter8));
  nand2 gate1242(.a(gate501inter8), .b(gate501inter7), .O(gate501inter9));
  nand2 gate1243(.a(s_99), .b(gate501inter3), .O(gate501inter10));
  nor2  gate1244(.a(gate501inter10), .b(gate501inter9), .O(gate501inter11));
  nor2  gate1245(.a(gate501inter11), .b(gate501inter6), .O(gate501inter12));
  nand2 gate1246(.a(gate501inter12), .b(gate501inter1), .O(G1310));
nand2 gate502( .a(G1266), .b(G1267), .O(G1311) );

  xor2  gate1597(.a(G1269), .b(G1268), .O(gate503inter0));
  nand2 gate1598(.a(gate503inter0), .b(s_150), .O(gate503inter1));
  and2  gate1599(.a(G1269), .b(G1268), .O(gate503inter2));
  inv1  gate1600(.a(s_150), .O(gate503inter3));
  inv1  gate1601(.a(s_151), .O(gate503inter4));
  nand2 gate1602(.a(gate503inter4), .b(gate503inter3), .O(gate503inter5));
  nor2  gate1603(.a(gate503inter5), .b(gate503inter2), .O(gate503inter6));
  inv1  gate1604(.a(G1268), .O(gate503inter7));
  inv1  gate1605(.a(G1269), .O(gate503inter8));
  nand2 gate1606(.a(gate503inter8), .b(gate503inter7), .O(gate503inter9));
  nand2 gate1607(.a(s_151), .b(gate503inter3), .O(gate503inter10));
  nor2  gate1608(.a(gate503inter10), .b(gate503inter9), .O(gate503inter11));
  nor2  gate1609(.a(gate503inter11), .b(gate503inter6), .O(gate503inter12));
  nand2 gate1610(.a(gate503inter12), .b(gate503inter1), .O(G1312));
nand2 gate504( .a(G1270), .b(G1271), .O(G1313) );

  xor2  gate2087(.a(G1273), .b(G1272), .O(gate505inter0));
  nand2 gate2088(.a(gate505inter0), .b(s_220), .O(gate505inter1));
  and2  gate2089(.a(G1273), .b(G1272), .O(gate505inter2));
  inv1  gate2090(.a(s_220), .O(gate505inter3));
  inv1  gate2091(.a(s_221), .O(gate505inter4));
  nand2 gate2092(.a(gate505inter4), .b(gate505inter3), .O(gate505inter5));
  nor2  gate2093(.a(gate505inter5), .b(gate505inter2), .O(gate505inter6));
  inv1  gate2094(.a(G1272), .O(gate505inter7));
  inv1  gate2095(.a(G1273), .O(gate505inter8));
  nand2 gate2096(.a(gate505inter8), .b(gate505inter7), .O(gate505inter9));
  nand2 gate2097(.a(s_221), .b(gate505inter3), .O(gate505inter10));
  nor2  gate2098(.a(gate505inter10), .b(gate505inter9), .O(gate505inter11));
  nor2  gate2099(.a(gate505inter11), .b(gate505inter6), .O(gate505inter12));
  nand2 gate2100(.a(gate505inter12), .b(gate505inter1), .O(G1314));
nand2 gate506( .a(G1274), .b(G1275), .O(G1315) );
nand2 gate507( .a(G1276), .b(G1277), .O(G1316) );
nand2 gate508( .a(G1278), .b(G1279), .O(G1317) );
nand2 gate509( .a(G1280), .b(G1281), .O(G1318) );
nand2 gate510( .a(G1282), .b(G1283), .O(G1319) );

  xor2  gate1303(.a(G1285), .b(G1284), .O(gate511inter0));
  nand2 gate1304(.a(gate511inter0), .b(s_108), .O(gate511inter1));
  and2  gate1305(.a(G1285), .b(G1284), .O(gate511inter2));
  inv1  gate1306(.a(s_108), .O(gate511inter3));
  inv1  gate1307(.a(s_109), .O(gate511inter4));
  nand2 gate1308(.a(gate511inter4), .b(gate511inter3), .O(gate511inter5));
  nor2  gate1309(.a(gate511inter5), .b(gate511inter2), .O(gate511inter6));
  inv1  gate1310(.a(G1284), .O(gate511inter7));
  inv1  gate1311(.a(G1285), .O(gate511inter8));
  nand2 gate1312(.a(gate511inter8), .b(gate511inter7), .O(gate511inter9));
  nand2 gate1313(.a(s_109), .b(gate511inter3), .O(gate511inter10));
  nor2  gate1314(.a(gate511inter10), .b(gate511inter9), .O(gate511inter11));
  nor2  gate1315(.a(gate511inter11), .b(gate511inter6), .O(gate511inter12));
  nand2 gate1316(.a(gate511inter12), .b(gate511inter1), .O(G1320));
nand2 gate512( .a(G1286), .b(G1287), .O(G1321) );
nand2 gate513( .a(G1288), .b(G1289), .O(G1322) );

  xor2  gate1695(.a(G1291), .b(G1290), .O(gate514inter0));
  nand2 gate1696(.a(gate514inter0), .b(s_164), .O(gate514inter1));
  and2  gate1697(.a(G1291), .b(G1290), .O(gate514inter2));
  inv1  gate1698(.a(s_164), .O(gate514inter3));
  inv1  gate1699(.a(s_165), .O(gate514inter4));
  nand2 gate1700(.a(gate514inter4), .b(gate514inter3), .O(gate514inter5));
  nor2  gate1701(.a(gate514inter5), .b(gate514inter2), .O(gate514inter6));
  inv1  gate1702(.a(G1290), .O(gate514inter7));
  inv1  gate1703(.a(G1291), .O(gate514inter8));
  nand2 gate1704(.a(gate514inter8), .b(gate514inter7), .O(gate514inter9));
  nand2 gate1705(.a(s_165), .b(gate514inter3), .O(gate514inter10));
  nor2  gate1706(.a(gate514inter10), .b(gate514inter9), .O(gate514inter11));
  nor2  gate1707(.a(gate514inter11), .b(gate514inter6), .O(gate514inter12));
  nand2 gate1708(.a(gate514inter12), .b(gate514inter1), .O(G1323));
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule