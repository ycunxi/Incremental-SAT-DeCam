module c499 (N1,N5,N9,N13,N17,N21,N25,N29,N33,N37,
             N41,N45,N49,N53,N57,N61,N65,N69,N73,N77,
             N81,N85,N89,N93,N97,N101,N105,N109,N113,N117,
             N121,N125,N129,N130,N131,N132,N133,N134,N135,N136,
             N137,N724,N725,N726,N727,N728,N729,N730,N731,N732,
             N733,N734,N735,N736,N737,N738,N739,N740,N741,N742,
             N743,N744,N745,N746,N747,N748,N749,N750,N751,N752,
             N753,N754,N755);

input N1,N5,N9,N13,N17,N21,N25,N29,N33,N37,
      N41,N45,N49,N53,N57,N61,N65,N69,N73,N77,
      N81,N85,N89,N93,N97,N101,N105,N109,N113,N117,
      N121,N125,N129,N130,N131,N132,N133,N134,N135,N136,
      N137;//RE__PI;

input s_0,s_1;//RE__ALLOW(00,01,10,11);
input s_2,s_3;//RE__ALLOW(00,01,10,11);
input s_4,s_5;//RE__ALLOW(00,01,10,11);
input s_6,s_7;//RE__ALLOW(00,01,10,11);
input s_8,s_9;//RE__ALLOW(00,01,10,11);
input s_10,s_11;//RE__ALLOW(00,01,10,11);
input s_12,s_13;//RE__ALLOW(00,01,10,11);
input s_14,s_15;//RE__ALLOW(00,01,10,11);
input s_16,s_17;//RE__ALLOW(00,01,10,11);
input s_18,s_19;//RE__ALLOW(00,01,10,11);
input s_20,s_21;//RE__ALLOW(00,01,10,11);
input s_22,s_23;//RE__ALLOW(00,01,10,11);
input s_24,s_25;//RE__ALLOW(00,01,10,11);
input s_26,s_27;//RE__ALLOW(00,01,10,11);
input s_28,s_29;//RE__ALLOW(00,01,10,11);
input s_30,s_31;//RE__ALLOW(00,01,10,11);
input s_32,s_33;//RE__ALLOW(00,01,10,11);
input s_34,s_35;//RE__ALLOW(00,01,10,11);
input s_36,s_37;//RE__ALLOW(00,01,10,11);
input s_38,s_39;//RE__ALLOW(00,01,10,11);
input s_40,s_41;//RE__ALLOW(00,01,10,11);
input s_42,s_43;//RE__ALLOW(00,01,10,11);
input s_44,s_45;//RE__ALLOW(00,01,10,11);
input s_46,s_47;//RE__ALLOW(00,01,10,11);
input s_48,s_49;//RE__ALLOW(00,01,10,11);
input s_50,s_51;//RE__ALLOW(00,01,10,11);
input s_52,s_53;//RE__ALLOW(00,01,10,11);
input s_54,s_55;//RE__ALLOW(00,01,10,11);
input s_56,s_57;//RE__ALLOW(00,01,10,11);
input s_58,s_59;//RE__ALLOW(00,01,10,11);
input s_60,s_61;//RE__ALLOW(00,01,10,11);
input s_62,s_63;//RE__ALLOW(00,01,10,11);
input s_64,s_65;//RE__ALLOW(00,01,10,11);
input s_66,s_67;//RE__ALLOW(00,01,10,11);
input s_68,s_69;//RE__ALLOW(00,01,10,11);
input s_70,s_71;//RE__ALLOW(00,01,10,11);
input s_72,s_73;//RE__ALLOW(00,01,10,11);
input s_74,s_75;//RE__ALLOW(00,01,10,11);
input s_76,s_77;//RE__ALLOW(00,01,10,11);
input s_78,s_79;//RE__ALLOW(00,01,10,11);
input s_80,s_81;//RE__ALLOW(00,01,10,11);
input s_82,s_83;//RE__ALLOW(00,01,10,11);
input s_84,s_85;//RE__ALLOW(00,01,10,11);
input s_86,s_87;//RE__ALLOW(00,01,10,11);
input s_88,s_89;//RE__ALLOW(00,01,10,11);
input s_90,s_91;//RE__ALLOW(00,01,10,11);
output N724,N725,N726,N727,N728,N729,N730,N731,N732,N733,
       N734,N735,N736,N737,N738,N739,N740,N741,N742,N743,
       N744,N745,N746,N747,N748,N749,N750,N751,N752,N753,
       N754,N755;

wire N250,N251,N252,N253,N254,N255,N256,N257,N258,N259,
     N260,N261,N262,N263,N264,N265,N266,N267,N268,N269,
     N270,N271,N272,N273,N274,N275,N276,N277,N278,N279,
     N280,N281,N282,N283,N284,N285,N286,N287,N288,N289,
     N290,N293,N296,N299,N302,N305,N308,N311,N314,N315,
     N316,N317,N318,N319,N320,N321,N338,N339,N340,N341,
     N342,N343,N344,N345,N346,N347,N348,N349,N350,N351,
     N352,N353,N354,N367,N380,N393,N406,N419,N432,N445,
     N554,N555,N556,N557,N558,N559,N560,N561,N562,N563,
     N564,N565,N566,N567,N568,N569,N570,N571,N572,N573,
     N574,N575,N576,N577,N578,N579,N580,N581,N582,N583,
     N584,N585,N586,N587,N588,N589,N590,N591,N592,N593,
     N594,N595,N596,N597,N598,N599,N600,N601,N602,N607,
     N620,N625,N630,N635,N640,N645,N650,N655,N692,N693,
     N694,N695,N696,N697,N698,N699,N700,N701,N702,N703,
     N704,N705,N706,N707,N708,N709,N710,N711,N712,N713,
     N714,N715,N716,N717,N718,N719,N720,N721,N722,N723, gate57inter0, gate57inter1, gate57inter2, gate57inter3, gate57inter4, gate57inter5, gate57inter6, gate57inter7, gate57inter8, gate57inter9, gate57inter10, gate57inter11, gate57inter12, gate37inter0, gate37inter1, gate37inter2, gate37inter3, gate37inter4, gate37inter5, gate37inter6, gate37inter7, gate37inter8, gate37inter9, gate37inter10, gate37inter11, gate37inter12, gate179inter0, gate179inter1, gate179inter2, gate179inter3, gate179inter4, gate179inter5, gate179inter6, gate179inter7, gate179inter8, gate179inter9, gate179inter10, gate179inter11, gate179inter12, gate75inter0, gate75inter1, gate75inter2, gate75inter3, gate75inter4, gate75inter5, gate75inter6, gate75inter7, gate75inter8, gate75inter9, gate75inter10, gate75inter11, gate75inter12, gate50inter0, gate50inter1, gate50inter2, gate50inter3, gate50inter4, gate50inter5, gate50inter6, gate50inter7, gate50inter8, gate50inter9, gate50inter10, gate50inter11, gate50inter12, gate56inter0, gate56inter1, gate56inter2, gate56inter3, gate56inter4, gate56inter5, gate56inter6, gate56inter7, gate56inter8, gate56inter9, gate56inter10, gate56inter11, gate56inter12, gate197inter0, gate197inter1, gate197inter2, gate197inter3, gate197inter4, gate197inter5, gate197inter6, gate197inter7, gate197inter8, gate197inter9, gate197inter10, gate197inter11, gate197inter12, gate33inter0, gate33inter1, gate33inter2, gate33inter3, gate33inter4, gate33inter5, gate33inter6, gate33inter7, gate33inter8, gate33inter9, gate33inter10, gate33inter11, gate33inter12, gate80inter0, gate80inter1, gate80inter2, gate80inter3, gate80inter4, gate80inter5, gate80inter6, gate80inter7, gate80inter8, gate80inter9, gate80inter10, gate80inter11, gate80inter12, gate26inter0, gate26inter1, gate26inter2, gate26inter3, gate26inter4, gate26inter5, gate26inter6, gate26inter7, gate26inter8, gate26inter9, gate26inter10, gate26inter11, gate26inter12, gate13inter0, gate13inter1, gate13inter2, gate13inter3, gate13inter4, gate13inter5, gate13inter6, gate13inter7, gate13inter8, gate13inter9, gate13inter10, gate13inter11, gate13inter12, gate65inter0, gate65inter1, gate65inter2, gate65inter3, gate65inter4, gate65inter5, gate65inter6, gate65inter7, gate65inter8, gate65inter9, gate65inter10, gate65inter11, gate65inter12, gate198inter0, gate198inter1, gate198inter2, gate198inter3, gate198inter4, gate198inter5, gate198inter6, gate198inter7, gate198inter8, gate198inter9, gate198inter10, gate198inter11, gate198inter12, gate42inter0, gate42inter1, gate42inter2, gate42inter3, gate42inter4, gate42inter5, gate42inter6, gate42inter7, gate42inter8, gate42inter9, gate42inter10, gate42inter11, gate42inter12, gate196inter0, gate196inter1, gate196inter2, gate196inter3, gate196inter4, gate196inter5, gate196inter6, gate196inter7, gate196inter8, gate196inter9, gate196inter10, gate196inter11, gate196inter12, gate176inter0, gate176inter1, gate176inter2, gate176inter3, gate176inter4, gate176inter5, gate176inter6, gate176inter7, gate176inter8, gate176inter9, gate176inter10, gate176inter11, gate176inter12, gate52inter0, gate52inter1, gate52inter2, gate52inter3, gate52inter4, gate52inter5, gate52inter6, gate52inter7, gate52inter8, gate52inter9, gate52inter10, gate52inter11, gate52inter12, gate178inter0, gate178inter1, gate178inter2, gate178inter3, gate178inter4, gate178inter5, gate178inter6, gate178inter7, gate178inter8, gate178inter9, gate178inter10, gate178inter11, gate178inter12, gate202inter0, gate202inter1, gate202inter2, gate202inter3, gate202inter4, gate202inter5, gate202inter6, gate202inter7, gate202inter8, gate202inter9, gate202inter10, gate202inter11, gate202inter12, gate199inter0, gate199inter1, gate199inter2, gate199inter3, gate199inter4, gate199inter5, gate199inter6, gate199inter7, gate199inter8, gate199inter9, gate199inter10, gate199inter11, gate199inter12, gate186inter0, gate186inter1, gate186inter2, gate186inter3, gate186inter4, gate186inter5, gate186inter6, gate186inter7, gate186inter8, gate186inter9, gate186inter10, gate186inter11, gate186inter12, gate200inter0, gate200inter1, gate200inter2, gate200inter3, gate200inter4, gate200inter5, gate200inter6, gate200inter7, gate200inter8, gate200inter9, gate200inter10, gate200inter11, gate200inter12, gate58inter0, gate58inter1, gate58inter2, gate58inter3, gate58inter4, gate58inter5, gate58inter6, gate58inter7, gate58inter8, gate58inter9, gate58inter10, gate58inter11, gate58inter12, gate27inter0, gate27inter1, gate27inter2, gate27inter3, gate27inter4, gate27inter5, gate27inter6, gate27inter7, gate27inter8, gate27inter9, gate27inter10, gate27inter11, gate27inter12, gate194inter0, gate194inter1, gate194inter2, gate194inter3, gate194inter4, gate194inter5, gate194inter6, gate194inter7, gate194inter8, gate194inter9, gate194inter10, gate194inter11, gate194inter12, gate16inter0, gate16inter1, gate16inter2, gate16inter3, gate16inter4, gate16inter5, gate16inter6, gate16inter7, gate16inter8, gate16inter9, gate16inter10, gate16inter11, gate16inter12, gate187inter0, gate187inter1, gate187inter2, gate187inter3, gate187inter4, gate187inter5, gate187inter6, gate187inter7, gate187inter8, gate187inter9, gate187inter10, gate187inter11, gate187inter12, gate15inter0, gate15inter1, gate15inter2, gate15inter3, gate15inter4, gate15inter5, gate15inter6, gate15inter7, gate15inter8, gate15inter9, gate15inter10, gate15inter11, gate15inter12, gate25inter0, gate25inter1, gate25inter2, gate25inter3, gate25inter4, gate25inter5, gate25inter6, gate25inter7, gate25inter8, gate25inter9, gate25inter10, gate25inter11, gate25inter12, gate73inter0, gate73inter1, gate73inter2, gate73inter3, gate73inter4, gate73inter5, gate73inter6, gate73inter7, gate73inter8, gate73inter9, gate73inter10, gate73inter11, gate73inter12, gate29inter0, gate29inter1, gate29inter2, gate29inter3, gate29inter4, gate29inter5, gate29inter6, gate29inter7, gate29inter8, gate29inter9, gate29inter10, gate29inter11, gate29inter12, gate38inter0, gate38inter1, gate38inter2, gate38inter3, gate38inter4, gate38inter5, gate38inter6, gate38inter7, gate38inter8, gate38inter9, gate38inter10, gate38inter11, gate38inter12, gate74inter0, gate74inter1, gate74inter2, gate74inter3, gate74inter4, gate74inter5, gate74inter6, gate74inter7, gate74inter8, gate74inter9, gate74inter10, gate74inter11, gate74inter12, gate1inter0, gate1inter1, gate1inter2, gate1inter3, gate1inter4, gate1inter5, gate1inter6, gate1inter7, gate1inter8, gate1inter9, gate1inter10, gate1inter11, gate1inter12, gate4inter0, gate4inter1, gate4inter2, gate4inter3, gate4inter4, gate4inter5, gate4inter6, gate4inter7, gate4inter8, gate4inter9, gate4inter10, gate4inter11, gate4inter12, gate195inter0, gate195inter1, gate195inter2, gate195inter3, gate195inter4, gate195inter5, gate195inter6, gate195inter7, gate195inter8, gate195inter9, gate195inter10, gate195inter11, gate195inter12, gate46inter0, gate46inter1, gate46inter2, gate46inter3, gate46inter4, gate46inter5, gate46inter6, gate46inter7, gate46inter8, gate46inter9, gate46inter10, gate46inter11, gate46inter12, gate177inter0, gate177inter1, gate177inter2, gate177inter3, gate177inter4, gate177inter5, gate177inter6, gate177inter7, gate177inter8, gate177inter9, gate177inter10, gate177inter11, gate177inter12, gate45inter0, gate45inter1, gate45inter2, gate45inter3, gate45inter4, gate45inter5, gate45inter6, gate45inter7, gate45inter8, gate45inter9, gate45inter10, gate45inter11, gate45inter12, gate34inter0, gate34inter1, gate34inter2, gate34inter3, gate34inter4, gate34inter5, gate34inter6, gate34inter7, gate34inter8, gate34inter9, gate34inter10, gate34inter11, gate34inter12, gate62inter0, gate62inter1, gate62inter2, gate62inter3, gate62inter4, gate62inter5, gate62inter6, gate62inter7, gate62inter8, gate62inter9, gate62inter10, gate62inter11, gate62inter12, gate9inter0, gate9inter1, gate9inter2, gate9inter3, gate9inter4, gate9inter5, gate9inter6, gate9inter7, gate9inter8, gate9inter9, gate9inter10, gate9inter11, gate9inter12, gate43inter0, gate43inter1, gate43inter2, gate43inter3, gate43inter4, gate43inter5, gate43inter6, gate43inter7, gate43inter8, gate43inter9, gate43inter10, gate43inter11, gate43inter12, gate14inter0, gate14inter1, gate14inter2, gate14inter3, gate14inter4, gate14inter5, gate14inter6, gate14inter7, gate14inter8, gate14inter9, gate14inter10, gate14inter11, gate14inter12, gate78inter0, gate78inter1, gate78inter2, gate78inter3, gate78inter4, gate78inter5, gate78inter6, gate78inter7, gate78inter8, gate78inter9, gate78inter10, gate78inter11, gate78inter12, gate11inter0, gate11inter1, gate11inter2, gate11inter3, gate11inter4, gate11inter5, gate11inter6, gate11inter7, gate11inter8, gate11inter9, gate11inter10, gate11inter11, gate11inter12;


  xor2  gate665(.a(N5), .b(N1), .O(gate1inter0));
  nand2 gate666(.a(gate1inter0), .b(s_66), .O(gate1inter1));
  and2  gate667(.a(N5), .b(N1), .O(gate1inter2));
  inv1  gate668(.a(s_66), .O(gate1inter3));
  inv1  gate669(.a(s_67), .O(gate1inter4));
  nand2 gate670(.a(gate1inter4), .b(gate1inter3), .O(gate1inter5));
  nor2  gate671(.a(gate1inter5), .b(gate1inter2), .O(gate1inter6));
  inv1  gate672(.a(N1), .O(gate1inter7));
  inv1  gate673(.a(N5), .O(gate1inter8));
  nand2 gate674(.a(gate1inter8), .b(gate1inter7), .O(gate1inter9));
  nand2 gate675(.a(s_67), .b(gate1inter3), .O(gate1inter10));
  nor2  gate676(.a(gate1inter10), .b(gate1inter9), .O(gate1inter11));
  nor2  gate677(.a(gate1inter11), .b(gate1inter6), .O(gate1inter12));
  nand2 gate678(.a(gate1inter12), .b(gate1inter1), .O(N250));
xor2 gate2( .a(N9), .b(N13), .O(N251) );
xor2 gate3( .a(N17), .b(N21), .O(N252) );

  xor2  gate679(.a(N29), .b(N25), .O(gate4inter0));
  nand2 gate680(.a(gate4inter0), .b(s_68), .O(gate4inter1));
  and2  gate681(.a(N29), .b(N25), .O(gate4inter2));
  inv1  gate682(.a(s_68), .O(gate4inter3));
  inv1  gate683(.a(s_69), .O(gate4inter4));
  nand2 gate684(.a(gate4inter4), .b(gate4inter3), .O(gate4inter5));
  nor2  gate685(.a(gate4inter5), .b(gate4inter2), .O(gate4inter6));
  inv1  gate686(.a(N25), .O(gate4inter7));
  inv1  gate687(.a(N29), .O(gate4inter8));
  nand2 gate688(.a(gate4inter8), .b(gate4inter7), .O(gate4inter9));
  nand2 gate689(.a(s_69), .b(gate4inter3), .O(gate4inter10));
  nor2  gate690(.a(gate4inter10), .b(gate4inter9), .O(gate4inter11));
  nor2  gate691(.a(gate4inter11), .b(gate4inter6), .O(gate4inter12));
  nand2 gate692(.a(gate4inter12), .b(gate4inter1), .O(N253));
xor2 gate5( .a(N33), .b(N37), .O(N254) );
xor2 gate6( .a(N41), .b(N45), .O(N255) );
xor2 gate7( .a(N49), .b(N53), .O(N256) );
xor2 gate8( .a(N57), .b(N61), .O(N257) );

  xor2  gate777(.a(N69), .b(N65), .O(gate9inter0));
  nand2 gate778(.a(gate9inter0), .b(s_82), .O(gate9inter1));
  and2  gate779(.a(N69), .b(N65), .O(gate9inter2));
  inv1  gate780(.a(s_82), .O(gate9inter3));
  inv1  gate781(.a(s_83), .O(gate9inter4));
  nand2 gate782(.a(gate9inter4), .b(gate9inter3), .O(gate9inter5));
  nor2  gate783(.a(gate9inter5), .b(gate9inter2), .O(gate9inter6));
  inv1  gate784(.a(N65), .O(gate9inter7));
  inv1  gate785(.a(N69), .O(gate9inter8));
  nand2 gate786(.a(gate9inter8), .b(gate9inter7), .O(gate9inter9));
  nand2 gate787(.a(s_83), .b(gate9inter3), .O(gate9inter10));
  nor2  gate788(.a(gate9inter10), .b(gate9inter9), .O(gate9inter11));
  nor2  gate789(.a(gate9inter11), .b(gate9inter6), .O(gate9inter12));
  nand2 gate790(.a(gate9inter12), .b(gate9inter1), .O(N258));
xor2 gate10( .a(N73), .b(N77), .O(N259) );

  xor2  gate833(.a(N85), .b(N81), .O(gate11inter0));
  nand2 gate834(.a(gate11inter0), .b(s_90), .O(gate11inter1));
  and2  gate835(.a(N85), .b(N81), .O(gate11inter2));
  inv1  gate836(.a(s_90), .O(gate11inter3));
  inv1  gate837(.a(s_91), .O(gate11inter4));
  nand2 gate838(.a(gate11inter4), .b(gate11inter3), .O(gate11inter5));
  nor2  gate839(.a(gate11inter5), .b(gate11inter2), .O(gate11inter6));
  inv1  gate840(.a(N81), .O(gate11inter7));
  inv1  gate841(.a(N85), .O(gate11inter8));
  nand2 gate842(.a(gate11inter8), .b(gate11inter7), .O(gate11inter9));
  nand2 gate843(.a(s_91), .b(gate11inter3), .O(gate11inter10));
  nor2  gate844(.a(gate11inter10), .b(gate11inter9), .O(gate11inter11));
  nor2  gate845(.a(gate11inter11), .b(gate11inter6), .O(gate11inter12));
  nand2 gate846(.a(gate11inter12), .b(gate11inter1), .O(N260));
xor2 gate12( .a(N89), .b(N93), .O(N261) );

  xor2  gate343(.a(N101), .b(N97), .O(gate13inter0));
  nand2 gate344(.a(gate13inter0), .b(s_20), .O(gate13inter1));
  and2  gate345(.a(N101), .b(N97), .O(gate13inter2));
  inv1  gate346(.a(s_20), .O(gate13inter3));
  inv1  gate347(.a(s_21), .O(gate13inter4));
  nand2 gate348(.a(gate13inter4), .b(gate13inter3), .O(gate13inter5));
  nor2  gate349(.a(gate13inter5), .b(gate13inter2), .O(gate13inter6));
  inv1  gate350(.a(N97), .O(gate13inter7));
  inv1  gate351(.a(N101), .O(gate13inter8));
  nand2 gate352(.a(gate13inter8), .b(gate13inter7), .O(gate13inter9));
  nand2 gate353(.a(s_21), .b(gate13inter3), .O(gate13inter10));
  nor2  gate354(.a(gate13inter10), .b(gate13inter9), .O(gate13inter11));
  nor2  gate355(.a(gate13inter11), .b(gate13inter6), .O(gate13inter12));
  nand2 gate356(.a(gate13inter12), .b(gate13inter1), .O(N262));

  xor2  gate805(.a(N109), .b(N105), .O(gate14inter0));
  nand2 gate806(.a(gate14inter0), .b(s_86), .O(gate14inter1));
  and2  gate807(.a(N109), .b(N105), .O(gate14inter2));
  inv1  gate808(.a(s_86), .O(gate14inter3));
  inv1  gate809(.a(s_87), .O(gate14inter4));
  nand2 gate810(.a(gate14inter4), .b(gate14inter3), .O(gate14inter5));
  nor2  gate811(.a(gate14inter5), .b(gate14inter2), .O(gate14inter6));
  inv1  gate812(.a(N105), .O(gate14inter7));
  inv1  gate813(.a(N109), .O(gate14inter8));
  nand2 gate814(.a(gate14inter8), .b(gate14inter7), .O(gate14inter9));
  nand2 gate815(.a(s_87), .b(gate14inter3), .O(gate14inter10));
  nor2  gate816(.a(gate14inter10), .b(gate14inter9), .O(gate14inter11));
  nor2  gate817(.a(gate14inter11), .b(gate14inter6), .O(gate14inter12));
  nand2 gate818(.a(gate14inter12), .b(gate14inter1), .O(N263));

  xor2  gate581(.a(N117), .b(N113), .O(gate15inter0));
  nand2 gate582(.a(gate15inter0), .b(s_54), .O(gate15inter1));
  and2  gate583(.a(N117), .b(N113), .O(gate15inter2));
  inv1  gate584(.a(s_54), .O(gate15inter3));
  inv1  gate585(.a(s_55), .O(gate15inter4));
  nand2 gate586(.a(gate15inter4), .b(gate15inter3), .O(gate15inter5));
  nor2  gate587(.a(gate15inter5), .b(gate15inter2), .O(gate15inter6));
  inv1  gate588(.a(N113), .O(gate15inter7));
  inv1  gate589(.a(N117), .O(gate15inter8));
  nand2 gate590(.a(gate15inter8), .b(gate15inter7), .O(gate15inter9));
  nand2 gate591(.a(s_55), .b(gate15inter3), .O(gate15inter10));
  nor2  gate592(.a(gate15inter10), .b(gate15inter9), .O(gate15inter11));
  nor2  gate593(.a(gate15inter11), .b(gate15inter6), .O(gate15inter12));
  nand2 gate594(.a(gate15inter12), .b(gate15inter1), .O(N264));

  xor2  gate553(.a(N125), .b(N121), .O(gate16inter0));
  nand2 gate554(.a(gate16inter0), .b(s_50), .O(gate16inter1));
  and2  gate555(.a(N125), .b(N121), .O(gate16inter2));
  inv1  gate556(.a(s_50), .O(gate16inter3));
  inv1  gate557(.a(s_51), .O(gate16inter4));
  nand2 gate558(.a(gate16inter4), .b(gate16inter3), .O(gate16inter5));
  nor2  gate559(.a(gate16inter5), .b(gate16inter2), .O(gate16inter6));
  inv1  gate560(.a(N121), .O(gate16inter7));
  inv1  gate561(.a(N125), .O(gate16inter8));
  nand2 gate562(.a(gate16inter8), .b(gate16inter7), .O(gate16inter9));
  nand2 gate563(.a(s_51), .b(gate16inter3), .O(gate16inter10));
  nor2  gate564(.a(gate16inter10), .b(gate16inter9), .O(gate16inter11));
  nor2  gate565(.a(gate16inter11), .b(gate16inter6), .O(gate16inter12));
  nand2 gate566(.a(gate16inter12), .b(gate16inter1), .O(N265));
and2 gate17( .a(N129), .b(N137), .O(N266) );
and2 gate18( .a(N130), .b(N137), .O(N267) );
and2 gate19( .a(N131), .b(N137), .O(N268) );
and2 gate20( .a(N132), .b(N137), .O(N269) );
and2 gate21( .a(N133), .b(N137), .O(N270) );
and2 gate22( .a(N134), .b(N137), .O(N271) );
and2 gate23( .a(N135), .b(N137), .O(N272) );
and2 gate24( .a(N136), .b(N137), .O(N273) );

  xor2  gate595(.a(N17), .b(N1), .O(gate25inter0));
  nand2 gate596(.a(gate25inter0), .b(s_56), .O(gate25inter1));
  and2  gate597(.a(N17), .b(N1), .O(gate25inter2));
  inv1  gate598(.a(s_56), .O(gate25inter3));
  inv1  gate599(.a(s_57), .O(gate25inter4));
  nand2 gate600(.a(gate25inter4), .b(gate25inter3), .O(gate25inter5));
  nor2  gate601(.a(gate25inter5), .b(gate25inter2), .O(gate25inter6));
  inv1  gate602(.a(N1), .O(gate25inter7));
  inv1  gate603(.a(N17), .O(gate25inter8));
  nand2 gate604(.a(gate25inter8), .b(gate25inter7), .O(gate25inter9));
  nand2 gate605(.a(s_57), .b(gate25inter3), .O(gate25inter10));
  nor2  gate606(.a(gate25inter10), .b(gate25inter9), .O(gate25inter11));
  nor2  gate607(.a(gate25inter11), .b(gate25inter6), .O(gate25inter12));
  nand2 gate608(.a(gate25inter12), .b(gate25inter1), .O(N274));

  xor2  gate329(.a(N49), .b(N33), .O(gate26inter0));
  nand2 gate330(.a(gate26inter0), .b(s_18), .O(gate26inter1));
  and2  gate331(.a(N49), .b(N33), .O(gate26inter2));
  inv1  gate332(.a(s_18), .O(gate26inter3));
  inv1  gate333(.a(s_19), .O(gate26inter4));
  nand2 gate334(.a(gate26inter4), .b(gate26inter3), .O(gate26inter5));
  nor2  gate335(.a(gate26inter5), .b(gate26inter2), .O(gate26inter6));
  inv1  gate336(.a(N33), .O(gate26inter7));
  inv1  gate337(.a(N49), .O(gate26inter8));
  nand2 gate338(.a(gate26inter8), .b(gate26inter7), .O(gate26inter9));
  nand2 gate339(.a(s_19), .b(gate26inter3), .O(gate26inter10));
  nor2  gate340(.a(gate26inter10), .b(gate26inter9), .O(gate26inter11));
  nor2  gate341(.a(gate26inter11), .b(gate26inter6), .O(gate26inter12));
  nand2 gate342(.a(gate26inter12), .b(gate26inter1), .O(N275));

  xor2  gate525(.a(N21), .b(N5), .O(gate27inter0));
  nand2 gate526(.a(gate27inter0), .b(s_46), .O(gate27inter1));
  and2  gate527(.a(N21), .b(N5), .O(gate27inter2));
  inv1  gate528(.a(s_46), .O(gate27inter3));
  inv1  gate529(.a(s_47), .O(gate27inter4));
  nand2 gate530(.a(gate27inter4), .b(gate27inter3), .O(gate27inter5));
  nor2  gate531(.a(gate27inter5), .b(gate27inter2), .O(gate27inter6));
  inv1  gate532(.a(N5), .O(gate27inter7));
  inv1  gate533(.a(N21), .O(gate27inter8));
  nand2 gate534(.a(gate27inter8), .b(gate27inter7), .O(gate27inter9));
  nand2 gate535(.a(s_47), .b(gate27inter3), .O(gate27inter10));
  nor2  gate536(.a(gate27inter10), .b(gate27inter9), .O(gate27inter11));
  nor2  gate537(.a(gate27inter11), .b(gate27inter6), .O(gate27inter12));
  nand2 gate538(.a(gate27inter12), .b(gate27inter1), .O(N276));
xor2 gate28( .a(N37), .b(N53), .O(N277) );

  xor2  gate623(.a(N25), .b(N9), .O(gate29inter0));
  nand2 gate624(.a(gate29inter0), .b(s_60), .O(gate29inter1));
  and2  gate625(.a(N25), .b(N9), .O(gate29inter2));
  inv1  gate626(.a(s_60), .O(gate29inter3));
  inv1  gate627(.a(s_61), .O(gate29inter4));
  nand2 gate628(.a(gate29inter4), .b(gate29inter3), .O(gate29inter5));
  nor2  gate629(.a(gate29inter5), .b(gate29inter2), .O(gate29inter6));
  inv1  gate630(.a(N9), .O(gate29inter7));
  inv1  gate631(.a(N25), .O(gate29inter8));
  nand2 gate632(.a(gate29inter8), .b(gate29inter7), .O(gate29inter9));
  nand2 gate633(.a(s_61), .b(gate29inter3), .O(gate29inter10));
  nor2  gate634(.a(gate29inter10), .b(gate29inter9), .O(gate29inter11));
  nor2  gate635(.a(gate29inter11), .b(gate29inter6), .O(gate29inter12));
  nand2 gate636(.a(gate29inter12), .b(gate29inter1), .O(N278));
xor2 gate30( .a(N41), .b(N57), .O(N279) );
xor2 gate31( .a(N13), .b(N29), .O(N280) );
xor2 gate32( .a(N45), .b(N61), .O(N281) );

  xor2  gate301(.a(N81), .b(N65), .O(gate33inter0));
  nand2 gate302(.a(gate33inter0), .b(s_14), .O(gate33inter1));
  and2  gate303(.a(N81), .b(N65), .O(gate33inter2));
  inv1  gate304(.a(s_14), .O(gate33inter3));
  inv1  gate305(.a(s_15), .O(gate33inter4));
  nand2 gate306(.a(gate33inter4), .b(gate33inter3), .O(gate33inter5));
  nor2  gate307(.a(gate33inter5), .b(gate33inter2), .O(gate33inter6));
  inv1  gate308(.a(N65), .O(gate33inter7));
  inv1  gate309(.a(N81), .O(gate33inter8));
  nand2 gate310(.a(gate33inter8), .b(gate33inter7), .O(gate33inter9));
  nand2 gate311(.a(s_15), .b(gate33inter3), .O(gate33inter10));
  nor2  gate312(.a(gate33inter10), .b(gate33inter9), .O(gate33inter11));
  nor2  gate313(.a(gate33inter11), .b(gate33inter6), .O(gate33inter12));
  nand2 gate314(.a(gate33inter12), .b(gate33inter1), .O(N282));

  xor2  gate749(.a(N113), .b(N97), .O(gate34inter0));
  nand2 gate750(.a(gate34inter0), .b(s_78), .O(gate34inter1));
  and2  gate751(.a(N113), .b(N97), .O(gate34inter2));
  inv1  gate752(.a(s_78), .O(gate34inter3));
  inv1  gate753(.a(s_79), .O(gate34inter4));
  nand2 gate754(.a(gate34inter4), .b(gate34inter3), .O(gate34inter5));
  nor2  gate755(.a(gate34inter5), .b(gate34inter2), .O(gate34inter6));
  inv1  gate756(.a(N97), .O(gate34inter7));
  inv1  gate757(.a(N113), .O(gate34inter8));
  nand2 gate758(.a(gate34inter8), .b(gate34inter7), .O(gate34inter9));
  nand2 gate759(.a(s_79), .b(gate34inter3), .O(gate34inter10));
  nor2  gate760(.a(gate34inter10), .b(gate34inter9), .O(gate34inter11));
  nor2  gate761(.a(gate34inter11), .b(gate34inter6), .O(gate34inter12));
  nand2 gate762(.a(gate34inter12), .b(gate34inter1), .O(N283));
xor2 gate35( .a(N69), .b(N85), .O(N284) );
xor2 gate36( .a(N101), .b(N117), .O(N285) );

  xor2  gate217(.a(N89), .b(N73), .O(gate37inter0));
  nand2 gate218(.a(gate37inter0), .b(s_2), .O(gate37inter1));
  and2  gate219(.a(N89), .b(N73), .O(gate37inter2));
  inv1  gate220(.a(s_2), .O(gate37inter3));
  inv1  gate221(.a(s_3), .O(gate37inter4));
  nand2 gate222(.a(gate37inter4), .b(gate37inter3), .O(gate37inter5));
  nor2  gate223(.a(gate37inter5), .b(gate37inter2), .O(gate37inter6));
  inv1  gate224(.a(N73), .O(gate37inter7));
  inv1  gate225(.a(N89), .O(gate37inter8));
  nand2 gate226(.a(gate37inter8), .b(gate37inter7), .O(gate37inter9));
  nand2 gate227(.a(s_3), .b(gate37inter3), .O(gate37inter10));
  nor2  gate228(.a(gate37inter10), .b(gate37inter9), .O(gate37inter11));
  nor2  gate229(.a(gate37inter11), .b(gate37inter6), .O(gate37inter12));
  nand2 gate230(.a(gate37inter12), .b(gate37inter1), .O(N286));

  xor2  gate637(.a(N121), .b(N105), .O(gate38inter0));
  nand2 gate638(.a(gate38inter0), .b(s_62), .O(gate38inter1));
  and2  gate639(.a(N121), .b(N105), .O(gate38inter2));
  inv1  gate640(.a(s_62), .O(gate38inter3));
  inv1  gate641(.a(s_63), .O(gate38inter4));
  nand2 gate642(.a(gate38inter4), .b(gate38inter3), .O(gate38inter5));
  nor2  gate643(.a(gate38inter5), .b(gate38inter2), .O(gate38inter6));
  inv1  gate644(.a(N105), .O(gate38inter7));
  inv1  gate645(.a(N121), .O(gate38inter8));
  nand2 gate646(.a(gate38inter8), .b(gate38inter7), .O(gate38inter9));
  nand2 gate647(.a(s_63), .b(gate38inter3), .O(gate38inter10));
  nor2  gate648(.a(gate38inter10), .b(gate38inter9), .O(gate38inter11));
  nor2  gate649(.a(gate38inter11), .b(gate38inter6), .O(gate38inter12));
  nand2 gate650(.a(gate38inter12), .b(gate38inter1), .O(N287));
xor2 gate39( .a(N77), .b(N93), .O(N288) );
xor2 gate40( .a(N109), .b(N125), .O(N289) );
xor2 gate41( .a(N250), .b(N251), .O(N290) );

  xor2  gate385(.a(N253), .b(N252), .O(gate42inter0));
  nand2 gate386(.a(gate42inter0), .b(s_26), .O(gate42inter1));
  and2  gate387(.a(N253), .b(N252), .O(gate42inter2));
  inv1  gate388(.a(s_26), .O(gate42inter3));
  inv1  gate389(.a(s_27), .O(gate42inter4));
  nand2 gate390(.a(gate42inter4), .b(gate42inter3), .O(gate42inter5));
  nor2  gate391(.a(gate42inter5), .b(gate42inter2), .O(gate42inter6));
  inv1  gate392(.a(N252), .O(gate42inter7));
  inv1  gate393(.a(N253), .O(gate42inter8));
  nand2 gate394(.a(gate42inter8), .b(gate42inter7), .O(gate42inter9));
  nand2 gate395(.a(s_27), .b(gate42inter3), .O(gate42inter10));
  nor2  gate396(.a(gate42inter10), .b(gate42inter9), .O(gate42inter11));
  nor2  gate397(.a(gate42inter11), .b(gate42inter6), .O(gate42inter12));
  nand2 gate398(.a(gate42inter12), .b(gate42inter1), .O(N293));

  xor2  gate791(.a(N255), .b(N254), .O(gate43inter0));
  nand2 gate792(.a(gate43inter0), .b(s_84), .O(gate43inter1));
  and2  gate793(.a(N255), .b(N254), .O(gate43inter2));
  inv1  gate794(.a(s_84), .O(gate43inter3));
  inv1  gate795(.a(s_85), .O(gate43inter4));
  nand2 gate796(.a(gate43inter4), .b(gate43inter3), .O(gate43inter5));
  nor2  gate797(.a(gate43inter5), .b(gate43inter2), .O(gate43inter6));
  inv1  gate798(.a(N254), .O(gate43inter7));
  inv1  gate799(.a(N255), .O(gate43inter8));
  nand2 gate800(.a(gate43inter8), .b(gate43inter7), .O(gate43inter9));
  nand2 gate801(.a(s_85), .b(gate43inter3), .O(gate43inter10));
  nor2  gate802(.a(gate43inter10), .b(gate43inter9), .O(gate43inter11));
  nor2  gate803(.a(gate43inter11), .b(gate43inter6), .O(gate43inter12));
  nand2 gate804(.a(gate43inter12), .b(gate43inter1), .O(N296));
xor2 gate44( .a(N256), .b(N257), .O(N299) );

  xor2  gate735(.a(N259), .b(N258), .O(gate45inter0));
  nand2 gate736(.a(gate45inter0), .b(s_76), .O(gate45inter1));
  and2  gate737(.a(N259), .b(N258), .O(gate45inter2));
  inv1  gate738(.a(s_76), .O(gate45inter3));
  inv1  gate739(.a(s_77), .O(gate45inter4));
  nand2 gate740(.a(gate45inter4), .b(gate45inter3), .O(gate45inter5));
  nor2  gate741(.a(gate45inter5), .b(gate45inter2), .O(gate45inter6));
  inv1  gate742(.a(N258), .O(gate45inter7));
  inv1  gate743(.a(N259), .O(gate45inter8));
  nand2 gate744(.a(gate45inter8), .b(gate45inter7), .O(gate45inter9));
  nand2 gate745(.a(s_77), .b(gate45inter3), .O(gate45inter10));
  nor2  gate746(.a(gate45inter10), .b(gate45inter9), .O(gate45inter11));
  nor2  gate747(.a(gate45inter11), .b(gate45inter6), .O(gate45inter12));
  nand2 gate748(.a(gate45inter12), .b(gate45inter1), .O(N302));

  xor2  gate707(.a(N261), .b(N260), .O(gate46inter0));
  nand2 gate708(.a(gate46inter0), .b(s_72), .O(gate46inter1));
  and2  gate709(.a(N261), .b(N260), .O(gate46inter2));
  inv1  gate710(.a(s_72), .O(gate46inter3));
  inv1  gate711(.a(s_73), .O(gate46inter4));
  nand2 gate712(.a(gate46inter4), .b(gate46inter3), .O(gate46inter5));
  nor2  gate713(.a(gate46inter5), .b(gate46inter2), .O(gate46inter6));
  inv1  gate714(.a(N260), .O(gate46inter7));
  inv1  gate715(.a(N261), .O(gate46inter8));
  nand2 gate716(.a(gate46inter8), .b(gate46inter7), .O(gate46inter9));
  nand2 gate717(.a(s_73), .b(gate46inter3), .O(gate46inter10));
  nor2  gate718(.a(gate46inter10), .b(gate46inter9), .O(gate46inter11));
  nor2  gate719(.a(gate46inter11), .b(gate46inter6), .O(gate46inter12));
  nand2 gate720(.a(gate46inter12), .b(gate46inter1), .O(N305));
xor2 gate47( .a(N262), .b(N263), .O(N308) );
xor2 gate48( .a(N264), .b(N265), .O(N311) );
xor2 gate49( .a(N274), .b(N275), .O(N314) );

  xor2  gate259(.a(N277), .b(N276), .O(gate50inter0));
  nand2 gate260(.a(gate50inter0), .b(s_8), .O(gate50inter1));
  and2  gate261(.a(N277), .b(N276), .O(gate50inter2));
  inv1  gate262(.a(s_8), .O(gate50inter3));
  inv1  gate263(.a(s_9), .O(gate50inter4));
  nand2 gate264(.a(gate50inter4), .b(gate50inter3), .O(gate50inter5));
  nor2  gate265(.a(gate50inter5), .b(gate50inter2), .O(gate50inter6));
  inv1  gate266(.a(N276), .O(gate50inter7));
  inv1  gate267(.a(N277), .O(gate50inter8));
  nand2 gate268(.a(gate50inter8), .b(gate50inter7), .O(gate50inter9));
  nand2 gate269(.a(s_9), .b(gate50inter3), .O(gate50inter10));
  nor2  gate270(.a(gate50inter10), .b(gate50inter9), .O(gate50inter11));
  nor2  gate271(.a(gate50inter11), .b(gate50inter6), .O(gate50inter12));
  nand2 gate272(.a(gate50inter12), .b(gate50inter1), .O(N315));
xor2 gate51( .a(N278), .b(N279), .O(N316) );

  xor2  gate427(.a(N281), .b(N280), .O(gate52inter0));
  nand2 gate428(.a(gate52inter0), .b(s_32), .O(gate52inter1));
  and2  gate429(.a(N281), .b(N280), .O(gate52inter2));
  inv1  gate430(.a(s_32), .O(gate52inter3));
  inv1  gate431(.a(s_33), .O(gate52inter4));
  nand2 gate432(.a(gate52inter4), .b(gate52inter3), .O(gate52inter5));
  nor2  gate433(.a(gate52inter5), .b(gate52inter2), .O(gate52inter6));
  inv1  gate434(.a(N280), .O(gate52inter7));
  inv1  gate435(.a(N281), .O(gate52inter8));
  nand2 gate436(.a(gate52inter8), .b(gate52inter7), .O(gate52inter9));
  nand2 gate437(.a(s_33), .b(gate52inter3), .O(gate52inter10));
  nor2  gate438(.a(gate52inter10), .b(gate52inter9), .O(gate52inter11));
  nor2  gate439(.a(gate52inter11), .b(gate52inter6), .O(gate52inter12));
  nand2 gate440(.a(gate52inter12), .b(gate52inter1), .O(N317));
xor2 gate53( .a(N282), .b(N283), .O(N318) );
xor2 gate54( .a(N284), .b(N285), .O(N319) );
xor2 gate55( .a(N286), .b(N287), .O(N320) );

  xor2  gate273(.a(N289), .b(N288), .O(gate56inter0));
  nand2 gate274(.a(gate56inter0), .b(s_10), .O(gate56inter1));
  and2  gate275(.a(N289), .b(N288), .O(gate56inter2));
  inv1  gate276(.a(s_10), .O(gate56inter3));
  inv1  gate277(.a(s_11), .O(gate56inter4));
  nand2 gate278(.a(gate56inter4), .b(gate56inter3), .O(gate56inter5));
  nor2  gate279(.a(gate56inter5), .b(gate56inter2), .O(gate56inter6));
  inv1  gate280(.a(N288), .O(gate56inter7));
  inv1  gate281(.a(N289), .O(gate56inter8));
  nand2 gate282(.a(gate56inter8), .b(gate56inter7), .O(gate56inter9));
  nand2 gate283(.a(s_11), .b(gate56inter3), .O(gate56inter10));
  nor2  gate284(.a(gate56inter10), .b(gate56inter9), .O(gate56inter11));
  nor2  gate285(.a(gate56inter11), .b(gate56inter6), .O(gate56inter12));
  nand2 gate286(.a(gate56inter12), .b(gate56inter1), .O(N321));

  xor2  gate203(.a(N293), .b(N290), .O(gate57inter0));
  nand2 gate204(.a(gate57inter0), .b(s_0), .O(gate57inter1));
  and2  gate205(.a(N293), .b(N290), .O(gate57inter2));
  inv1  gate206(.a(s_0), .O(gate57inter3));
  inv1  gate207(.a(s_1), .O(gate57inter4));
  nand2 gate208(.a(gate57inter4), .b(gate57inter3), .O(gate57inter5));
  nor2  gate209(.a(gate57inter5), .b(gate57inter2), .O(gate57inter6));
  inv1  gate210(.a(N290), .O(gate57inter7));
  inv1  gate211(.a(N293), .O(gate57inter8));
  nand2 gate212(.a(gate57inter8), .b(gate57inter7), .O(gate57inter9));
  nand2 gate213(.a(s_1), .b(gate57inter3), .O(gate57inter10));
  nor2  gate214(.a(gate57inter10), .b(gate57inter9), .O(gate57inter11));
  nor2  gate215(.a(gate57inter11), .b(gate57inter6), .O(gate57inter12));
  nand2 gate216(.a(gate57inter12), .b(gate57inter1), .O(N338));

  xor2  gate511(.a(N299), .b(N296), .O(gate58inter0));
  nand2 gate512(.a(gate58inter0), .b(s_44), .O(gate58inter1));
  and2  gate513(.a(N299), .b(N296), .O(gate58inter2));
  inv1  gate514(.a(s_44), .O(gate58inter3));
  inv1  gate515(.a(s_45), .O(gate58inter4));
  nand2 gate516(.a(gate58inter4), .b(gate58inter3), .O(gate58inter5));
  nor2  gate517(.a(gate58inter5), .b(gate58inter2), .O(gate58inter6));
  inv1  gate518(.a(N296), .O(gate58inter7));
  inv1  gate519(.a(N299), .O(gate58inter8));
  nand2 gate520(.a(gate58inter8), .b(gate58inter7), .O(gate58inter9));
  nand2 gate521(.a(s_45), .b(gate58inter3), .O(gate58inter10));
  nor2  gate522(.a(gate58inter10), .b(gate58inter9), .O(gate58inter11));
  nor2  gate523(.a(gate58inter11), .b(gate58inter6), .O(gate58inter12));
  nand2 gate524(.a(gate58inter12), .b(gate58inter1), .O(N339));
xor2 gate59( .a(N290), .b(N296), .O(N340) );
xor2 gate60( .a(N293), .b(N299), .O(N341) );
xor2 gate61( .a(N302), .b(N305), .O(N342) );

  xor2  gate763(.a(N311), .b(N308), .O(gate62inter0));
  nand2 gate764(.a(gate62inter0), .b(s_80), .O(gate62inter1));
  and2  gate765(.a(N311), .b(N308), .O(gate62inter2));
  inv1  gate766(.a(s_80), .O(gate62inter3));
  inv1  gate767(.a(s_81), .O(gate62inter4));
  nand2 gate768(.a(gate62inter4), .b(gate62inter3), .O(gate62inter5));
  nor2  gate769(.a(gate62inter5), .b(gate62inter2), .O(gate62inter6));
  inv1  gate770(.a(N308), .O(gate62inter7));
  inv1  gate771(.a(N311), .O(gate62inter8));
  nand2 gate772(.a(gate62inter8), .b(gate62inter7), .O(gate62inter9));
  nand2 gate773(.a(s_81), .b(gate62inter3), .O(gate62inter10));
  nor2  gate774(.a(gate62inter10), .b(gate62inter9), .O(gate62inter11));
  nor2  gate775(.a(gate62inter11), .b(gate62inter6), .O(gate62inter12));
  nand2 gate776(.a(gate62inter12), .b(gate62inter1), .O(N343));
xor2 gate63( .a(N302), .b(N308), .O(N344) );
xor2 gate64( .a(N305), .b(N311), .O(N345) );

  xor2  gate357(.a(N342), .b(N266), .O(gate65inter0));
  nand2 gate358(.a(gate65inter0), .b(s_22), .O(gate65inter1));
  and2  gate359(.a(N342), .b(N266), .O(gate65inter2));
  inv1  gate360(.a(s_22), .O(gate65inter3));
  inv1  gate361(.a(s_23), .O(gate65inter4));
  nand2 gate362(.a(gate65inter4), .b(gate65inter3), .O(gate65inter5));
  nor2  gate363(.a(gate65inter5), .b(gate65inter2), .O(gate65inter6));
  inv1  gate364(.a(N266), .O(gate65inter7));
  inv1  gate365(.a(N342), .O(gate65inter8));
  nand2 gate366(.a(gate65inter8), .b(gate65inter7), .O(gate65inter9));
  nand2 gate367(.a(s_23), .b(gate65inter3), .O(gate65inter10));
  nor2  gate368(.a(gate65inter10), .b(gate65inter9), .O(gate65inter11));
  nor2  gate369(.a(gate65inter11), .b(gate65inter6), .O(gate65inter12));
  nand2 gate370(.a(gate65inter12), .b(gate65inter1), .O(N346));
xor2 gate66( .a(N267), .b(N343), .O(N347) );
xor2 gate67( .a(N268), .b(N344), .O(N348) );
xor2 gate68( .a(N269), .b(N345), .O(N349) );
xor2 gate69( .a(N270), .b(N338), .O(N350) );
xor2 gate70( .a(N271), .b(N339), .O(N351) );
xor2 gate71( .a(N272), .b(N340), .O(N352) );
xor2 gate72( .a(N273), .b(N341), .O(N353) );

  xor2  gate609(.a(N346), .b(N314), .O(gate73inter0));
  nand2 gate610(.a(gate73inter0), .b(s_58), .O(gate73inter1));
  and2  gate611(.a(N346), .b(N314), .O(gate73inter2));
  inv1  gate612(.a(s_58), .O(gate73inter3));
  inv1  gate613(.a(s_59), .O(gate73inter4));
  nand2 gate614(.a(gate73inter4), .b(gate73inter3), .O(gate73inter5));
  nor2  gate615(.a(gate73inter5), .b(gate73inter2), .O(gate73inter6));
  inv1  gate616(.a(N314), .O(gate73inter7));
  inv1  gate617(.a(N346), .O(gate73inter8));
  nand2 gate618(.a(gate73inter8), .b(gate73inter7), .O(gate73inter9));
  nand2 gate619(.a(s_59), .b(gate73inter3), .O(gate73inter10));
  nor2  gate620(.a(gate73inter10), .b(gate73inter9), .O(gate73inter11));
  nor2  gate621(.a(gate73inter11), .b(gate73inter6), .O(gate73inter12));
  nand2 gate622(.a(gate73inter12), .b(gate73inter1), .O(N354));

  xor2  gate651(.a(N347), .b(N315), .O(gate74inter0));
  nand2 gate652(.a(gate74inter0), .b(s_64), .O(gate74inter1));
  and2  gate653(.a(N347), .b(N315), .O(gate74inter2));
  inv1  gate654(.a(s_64), .O(gate74inter3));
  inv1  gate655(.a(s_65), .O(gate74inter4));
  nand2 gate656(.a(gate74inter4), .b(gate74inter3), .O(gate74inter5));
  nor2  gate657(.a(gate74inter5), .b(gate74inter2), .O(gate74inter6));
  inv1  gate658(.a(N315), .O(gate74inter7));
  inv1  gate659(.a(N347), .O(gate74inter8));
  nand2 gate660(.a(gate74inter8), .b(gate74inter7), .O(gate74inter9));
  nand2 gate661(.a(s_65), .b(gate74inter3), .O(gate74inter10));
  nor2  gate662(.a(gate74inter10), .b(gate74inter9), .O(gate74inter11));
  nor2  gate663(.a(gate74inter11), .b(gate74inter6), .O(gate74inter12));
  nand2 gate664(.a(gate74inter12), .b(gate74inter1), .O(N367));

  xor2  gate245(.a(N348), .b(N316), .O(gate75inter0));
  nand2 gate246(.a(gate75inter0), .b(s_6), .O(gate75inter1));
  and2  gate247(.a(N348), .b(N316), .O(gate75inter2));
  inv1  gate248(.a(s_6), .O(gate75inter3));
  inv1  gate249(.a(s_7), .O(gate75inter4));
  nand2 gate250(.a(gate75inter4), .b(gate75inter3), .O(gate75inter5));
  nor2  gate251(.a(gate75inter5), .b(gate75inter2), .O(gate75inter6));
  inv1  gate252(.a(N316), .O(gate75inter7));
  inv1  gate253(.a(N348), .O(gate75inter8));
  nand2 gate254(.a(gate75inter8), .b(gate75inter7), .O(gate75inter9));
  nand2 gate255(.a(s_7), .b(gate75inter3), .O(gate75inter10));
  nor2  gate256(.a(gate75inter10), .b(gate75inter9), .O(gate75inter11));
  nor2  gate257(.a(gate75inter11), .b(gate75inter6), .O(gate75inter12));
  nand2 gate258(.a(gate75inter12), .b(gate75inter1), .O(N380));
xor2 gate76( .a(N317), .b(N349), .O(N393) );
xor2 gate77( .a(N318), .b(N350), .O(N406) );

  xor2  gate819(.a(N351), .b(N319), .O(gate78inter0));
  nand2 gate820(.a(gate78inter0), .b(s_88), .O(gate78inter1));
  and2  gate821(.a(N351), .b(N319), .O(gate78inter2));
  inv1  gate822(.a(s_88), .O(gate78inter3));
  inv1  gate823(.a(s_89), .O(gate78inter4));
  nand2 gate824(.a(gate78inter4), .b(gate78inter3), .O(gate78inter5));
  nor2  gate825(.a(gate78inter5), .b(gate78inter2), .O(gate78inter6));
  inv1  gate826(.a(N319), .O(gate78inter7));
  inv1  gate827(.a(N351), .O(gate78inter8));
  nand2 gate828(.a(gate78inter8), .b(gate78inter7), .O(gate78inter9));
  nand2 gate829(.a(s_89), .b(gate78inter3), .O(gate78inter10));
  nor2  gate830(.a(gate78inter10), .b(gate78inter9), .O(gate78inter11));
  nor2  gate831(.a(gate78inter11), .b(gate78inter6), .O(gate78inter12));
  nand2 gate832(.a(gate78inter12), .b(gate78inter1), .O(N419));
xor2 gate79( .a(N320), .b(N352), .O(N432) );

  xor2  gate315(.a(N353), .b(N321), .O(gate80inter0));
  nand2 gate316(.a(gate80inter0), .b(s_16), .O(gate80inter1));
  and2  gate317(.a(N353), .b(N321), .O(gate80inter2));
  inv1  gate318(.a(s_16), .O(gate80inter3));
  inv1  gate319(.a(s_17), .O(gate80inter4));
  nand2 gate320(.a(gate80inter4), .b(gate80inter3), .O(gate80inter5));
  nor2  gate321(.a(gate80inter5), .b(gate80inter2), .O(gate80inter6));
  inv1  gate322(.a(N321), .O(gate80inter7));
  inv1  gate323(.a(N353), .O(gate80inter8));
  nand2 gate324(.a(gate80inter8), .b(gate80inter7), .O(gate80inter9));
  nand2 gate325(.a(s_17), .b(gate80inter3), .O(gate80inter10));
  nor2  gate326(.a(gate80inter10), .b(gate80inter9), .O(gate80inter11));
  nor2  gate327(.a(gate80inter11), .b(gate80inter6), .O(gate80inter12));
  nand2 gate328(.a(gate80inter12), .b(gate80inter1), .O(N445));
inv1 gate81( .a(N354), .O(N554) );
inv1 gate82( .a(N367), .O(N555) );
inv1 gate83( .a(N380), .O(N556) );
inv1 gate84( .a(N354), .O(N557) );
inv1 gate85( .a(N367), .O(N558) );
inv1 gate86( .a(N393), .O(N559) );
inv1 gate87( .a(N354), .O(N560) );
inv1 gate88( .a(N380), .O(N561) );
inv1 gate89( .a(N393), .O(N562) );
inv1 gate90( .a(N367), .O(N563) );
inv1 gate91( .a(N380), .O(N564) );
inv1 gate92( .a(N393), .O(N565) );
inv1 gate93( .a(N419), .O(N566) );
inv1 gate94( .a(N445), .O(N567) );
inv1 gate95( .a(N419), .O(N568) );
inv1 gate96( .a(N432), .O(N569) );
inv1 gate97( .a(N406), .O(N570) );
inv1 gate98( .a(N445), .O(N571) );
inv1 gate99( .a(N406), .O(N572) );
inv1 gate100( .a(N432), .O(N573) );
inv1 gate101( .a(N406), .O(N574) );
inv1 gate102( .a(N419), .O(N575) );
inv1 gate103( .a(N432), .O(N576) );
inv1 gate104( .a(N406), .O(N577) );
inv1 gate105( .a(N419), .O(N578) );
inv1 gate106( .a(N445), .O(N579) );
inv1 gate107( .a(N406), .O(N580) );
inv1 gate108( .a(N432), .O(N581) );
inv1 gate109( .a(N445), .O(N582) );
inv1 gate110( .a(N419), .O(N583) );
inv1 gate111( .a(N432), .O(N584) );
inv1 gate112( .a(N445), .O(N585) );
inv1 gate113( .a(N367), .O(N586) );
inv1 gate114( .a(N393), .O(N587) );
inv1 gate115( .a(N367), .O(N588) );
inv1 gate116( .a(N380), .O(N589) );
inv1 gate117( .a(N354), .O(N590) );
inv1 gate118( .a(N393), .O(N591) );
inv1 gate119( .a(N354), .O(N592) );
inv1 gate120( .a(N380), .O(N593) );
and4 gate121( .a(N554), .b(N555), .c(N556), .d(N393), .O(N594) );
and4 gate122( .a(N557), .b(N558), .c(N380), .d(N559), .O(N595) );
and4 gate123( .a(N560), .b(N367), .c(N561), .d(N562), .O(N596) );
and4 gate124( .a(N354), .b(N563), .c(N564), .d(N565), .O(N597) );
and4 gate125( .a(N574), .b(N575), .c(N576), .d(N445), .O(N598) );
and4 gate126( .a(N577), .b(N578), .c(N432), .d(N579), .O(N599) );
and4 gate127( .a(N580), .b(N419), .c(N581), .d(N582), .O(N600) );
and4 gate128( .a(N406), .b(N583), .c(N584), .d(N585), .O(N601) );
or4 gate129( .a(N594), .b(N595), .c(N596), .d(N597), .O(N602) );
or4 gate130( .a(N598), .b(N599), .c(N600), .d(N601), .O(N607) );
and5 gate131( .a(N406), .b(N566), .c(N432), .d(N567), .e(N602), .O(N620) );
and5 gate132( .a(N406), .b(N568), .c(N569), .d(N445), .e(N602), .O(N625) );
and5 gate133( .a(N570), .b(N419), .c(N432), .d(N571), .e(N602), .O(N630) );
and5 gate134( .a(N572), .b(N419), .c(N573), .d(N445), .e(N602), .O(N635) );
and5 gate135( .a(N354), .b(N586), .c(N380), .d(N587), .e(N607), .O(N640) );
and5 gate136( .a(N354), .b(N588), .c(N589), .d(N393), .e(N607), .O(N645) );
and5 gate137( .a(N590), .b(N367), .c(N380), .d(N591), .e(N607), .O(N650) );
and5 gate138( .a(N592), .b(N367), .c(N593), .d(N393), .e(N607), .O(N655) );
and2 gate139( .a(N354), .b(N620), .O(N692) );
and2 gate140( .a(N367), .b(N620), .O(N693) );
and2 gate141( .a(N380), .b(N620), .O(N694) );
and2 gate142( .a(N393), .b(N620), .O(N695) );
and2 gate143( .a(N354), .b(N625), .O(N696) );
and2 gate144( .a(N367), .b(N625), .O(N697) );
and2 gate145( .a(N380), .b(N625), .O(N698) );
and2 gate146( .a(N393), .b(N625), .O(N699) );
and2 gate147( .a(N354), .b(N630), .O(N700) );
and2 gate148( .a(N367), .b(N630), .O(N701) );
and2 gate149( .a(N380), .b(N630), .O(N702) );
and2 gate150( .a(N393), .b(N630), .O(N703) );
and2 gate151( .a(N354), .b(N635), .O(N704) );
and2 gate152( .a(N367), .b(N635), .O(N705) );
and2 gate153( .a(N380), .b(N635), .O(N706) );
and2 gate154( .a(N393), .b(N635), .O(N707) );
and2 gate155( .a(N406), .b(N640), .O(N708) );
and2 gate156( .a(N419), .b(N640), .O(N709) );
and2 gate157( .a(N432), .b(N640), .O(N710) );
and2 gate158( .a(N445), .b(N640), .O(N711) );
and2 gate159( .a(N406), .b(N645), .O(N712) );
and2 gate160( .a(N419), .b(N645), .O(N713) );
and2 gate161( .a(N432), .b(N645), .O(N714) );
and2 gate162( .a(N445), .b(N645), .O(N715) );
and2 gate163( .a(N406), .b(N650), .O(N716) );
and2 gate164( .a(N419), .b(N650), .O(N717) );
and2 gate165( .a(N432), .b(N650), .O(N718) );
and2 gate166( .a(N445), .b(N650), .O(N719) );
and2 gate167( .a(N406), .b(N655), .O(N720) );
and2 gate168( .a(N419), .b(N655), .O(N721) );
and2 gate169( .a(N432), .b(N655), .O(N722) );
and2 gate170( .a(N445), .b(N655), .O(N723) );
xor2 gate171( .a(N1), .b(N692), .O(N724) );
xor2 gate172( .a(N5), .b(N693), .O(N725) );
xor2 gate173( .a(N9), .b(N694), .O(N726) );
xor2 gate174( .a(N13), .b(N695), .O(N727) );
xor2 gate175( .a(N17), .b(N696), .O(N728) );

  xor2  gate413(.a(N697), .b(N21), .O(gate176inter0));
  nand2 gate414(.a(gate176inter0), .b(s_30), .O(gate176inter1));
  and2  gate415(.a(N697), .b(N21), .O(gate176inter2));
  inv1  gate416(.a(s_30), .O(gate176inter3));
  inv1  gate417(.a(s_31), .O(gate176inter4));
  nand2 gate418(.a(gate176inter4), .b(gate176inter3), .O(gate176inter5));
  nor2  gate419(.a(gate176inter5), .b(gate176inter2), .O(gate176inter6));
  inv1  gate420(.a(N21), .O(gate176inter7));
  inv1  gate421(.a(N697), .O(gate176inter8));
  nand2 gate422(.a(gate176inter8), .b(gate176inter7), .O(gate176inter9));
  nand2 gate423(.a(s_31), .b(gate176inter3), .O(gate176inter10));
  nor2  gate424(.a(gate176inter10), .b(gate176inter9), .O(gate176inter11));
  nor2  gate425(.a(gate176inter11), .b(gate176inter6), .O(gate176inter12));
  nand2 gate426(.a(gate176inter12), .b(gate176inter1), .O(N729));

  xor2  gate721(.a(N698), .b(N25), .O(gate177inter0));
  nand2 gate722(.a(gate177inter0), .b(s_74), .O(gate177inter1));
  and2  gate723(.a(N698), .b(N25), .O(gate177inter2));
  inv1  gate724(.a(s_74), .O(gate177inter3));
  inv1  gate725(.a(s_75), .O(gate177inter4));
  nand2 gate726(.a(gate177inter4), .b(gate177inter3), .O(gate177inter5));
  nor2  gate727(.a(gate177inter5), .b(gate177inter2), .O(gate177inter6));
  inv1  gate728(.a(N25), .O(gate177inter7));
  inv1  gate729(.a(N698), .O(gate177inter8));
  nand2 gate730(.a(gate177inter8), .b(gate177inter7), .O(gate177inter9));
  nand2 gate731(.a(s_75), .b(gate177inter3), .O(gate177inter10));
  nor2  gate732(.a(gate177inter10), .b(gate177inter9), .O(gate177inter11));
  nor2  gate733(.a(gate177inter11), .b(gate177inter6), .O(gate177inter12));
  nand2 gate734(.a(gate177inter12), .b(gate177inter1), .O(N730));

  xor2  gate441(.a(N699), .b(N29), .O(gate178inter0));
  nand2 gate442(.a(gate178inter0), .b(s_34), .O(gate178inter1));
  and2  gate443(.a(N699), .b(N29), .O(gate178inter2));
  inv1  gate444(.a(s_34), .O(gate178inter3));
  inv1  gate445(.a(s_35), .O(gate178inter4));
  nand2 gate446(.a(gate178inter4), .b(gate178inter3), .O(gate178inter5));
  nor2  gate447(.a(gate178inter5), .b(gate178inter2), .O(gate178inter6));
  inv1  gate448(.a(N29), .O(gate178inter7));
  inv1  gate449(.a(N699), .O(gate178inter8));
  nand2 gate450(.a(gate178inter8), .b(gate178inter7), .O(gate178inter9));
  nand2 gate451(.a(s_35), .b(gate178inter3), .O(gate178inter10));
  nor2  gate452(.a(gate178inter10), .b(gate178inter9), .O(gate178inter11));
  nor2  gate453(.a(gate178inter11), .b(gate178inter6), .O(gate178inter12));
  nand2 gate454(.a(gate178inter12), .b(gate178inter1), .O(N731));

  xor2  gate231(.a(N700), .b(N33), .O(gate179inter0));
  nand2 gate232(.a(gate179inter0), .b(s_4), .O(gate179inter1));
  and2  gate233(.a(N700), .b(N33), .O(gate179inter2));
  inv1  gate234(.a(s_4), .O(gate179inter3));
  inv1  gate235(.a(s_5), .O(gate179inter4));
  nand2 gate236(.a(gate179inter4), .b(gate179inter3), .O(gate179inter5));
  nor2  gate237(.a(gate179inter5), .b(gate179inter2), .O(gate179inter6));
  inv1  gate238(.a(N33), .O(gate179inter7));
  inv1  gate239(.a(N700), .O(gate179inter8));
  nand2 gate240(.a(gate179inter8), .b(gate179inter7), .O(gate179inter9));
  nand2 gate241(.a(s_5), .b(gate179inter3), .O(gate179inter10));
  nor2  gate242(.a(gate179inter10), .b(gate179inter9), .O(gate179inter11));
  nor2  gate243(.a(gate179inter11), .b(gate179inter6), .O(gate179inter12));
  nand2 gate244(.a(gate179inter12), .b(gate179inter1), .O(N732));
xor2 gate180( .a(N37), .b(N701), .O(N733) );
xor2 gate181( .a(N41), .b(N702), .O(N734) );
xor2 gate182( .a(N45), .b(N703), .O(N735) );
xor2 gate183( .a(N49), .b(N704), .O(N736) );
xor2 gate184( .a(N53), .b(N705), .O(N737) );
xor2 gate185( .a(N57), .b(N706), .O(N738) );

  xor2  gate483(.a(N707), .b(N61), .O(gate186inter0));
  nand2 gate484(.a(gate186inter0), .b(s_40), .O(gate186inter1));
  and2  gate485(.a(N707), .b(N61), .O(gate186inter2));
  inv1  gate486(.a(s_40), .O(gate186inter3));
  inv1  gate487(.a(s_41), .O(gate186inter4));
  nand2 gate488(.a(gate186inter4), .b(gate186inter3), .O(gate186inter5));
  nor2  gate489(.a(gate186inter5), .b(gate186inter2), .O(gate186inter6));
  inv1  gate490(.a(N61), .O(gate186inter7));
  inv1  gate491(.a(N707), .O(gate186inter8));
  nand2 gate492(.a(gate186inter8), .b(gate186inter7), .O(gate186inter9));
  nand2 gate493(.a(s_41), .b(gate186inter3), .O(gate186inter10));
  nor2  gate494(.a(gate186inter10), .b(gate186inter9), .O(gate186inter11));
  nor2  gate495(.a(gate186inter11), .b(gate186inter6), .O(gate186inter12));
  nand2 gate496(.a(gate186inter12), .b(gate186inter1), .O(N739));

  xor2  gate567(.a(N708), .b(N65), .O(gate187inter0));
  nand2 gate568(.a(gate187inter0), .b(s_52), .O(gate187inter1));
  and2  gate569(.a(N708), .b(N65), .O(gate187inter2));
  inv1  gate570(.a(s_52), .O(gate187inter3));
  inv1  gate571(.a(s_53), .O(gate187inter4));
  nand2 gate572(.a(gate187inter4), .b(gate187inter3), .O(gate187inter5));
  nor2  gate573(.a(gate187inter5), .b(gate187inter2), .O(gate187inter6));
  inv1  gate574(.a(N65), .O(gate187inter7));
  inv1  gate575(.a(N708), .O(gate187inter8));
  nand2 gate576(.a(gate187inter8), .b(gate187inter7), .O(gate187inter9));
  nand2 gate577(.a(s_53), .b(gate187inter3), .O(gate187inter10));
  nor2  gate578(.a(gate187inter10), .b(gate187inter9), .O(gate187inter11));
  nor2  gate579(.a(gate187inter11), .b(gate187inter6), .O(gate187inter12));
  nand2 gate580(.a(gate187inter12), .b(gate187inter1), .O(N740));
xor2 gate188( .a(N69), .b(N709), .O(N741) );
xor2 gate189( .a(N73), .b(N710), .O(N742) );
xor2 gate190( .a(N77), .b(N711), .O(N743) );
xor2 gate191( .a(N81), .b(N712), .O(N744) );
xor2 gate192( .a(N85), .b(N713), .O(N745) );
xor2 gate193( .a(N89), .b(N714), .O(N746) );

  xor2  gate539(.a(N715), .b(N93), .O(gate194inter0));
  nand2 gate540(.a(gate194inter0), .b(s_48), .O(gate194inter1));
  and2  gate541(.a(N715), .b(N93), .O(gate194inter2));
  inv1  gate542(.a(s_48), .O(gate194inter3));
  inv1  gate543(.a(s_49), .O(gate194inter4));
  nand2 gate544(.a(gate194inter4), .b(gate194inter3), .O(gate194inter5));
  nor2  gate545(.a(gate194inter5), .b(gate194inter2), .O(gate194inter6));
  inv1  gate546(.a(N93), .O(gate194inter7));
  inv1  gate547(.a(N715), .O(gate194inter8));
  nand2 gate548(.a(gate194inter8), .b(gate194inter7), .O(gate194inter9));
  nand2 gate549(.a(s_49), .b(gate194inter3), .O(gate194inter10));
  nor2  gate550(.a(gate194inter10), .b(gate194inter9), .O(gate194inter11));
  nor2  gate551(.a(gate194inter11), .b(gate194inter6), .O(gate194inter12));
  nand2 gate552(.a(gate194inter12), .b(gate194inter1), .O(N747));

  xor2  gate693(.a(N716), .b(N97), .O(gate195inter0));
  nand2 gate694(.a(gate195inter0), .b(s_70), .O(gate195inter1));
  and2  gate695(.a(N716), .b(N97), .O(gate195inter2));
  inv1  gate696(.a(s_70), .O(gate195inter3));
  inv1  gate697(.a(s_71), .O(gate195inter4));
  nand2 gate698(.a(gate195inter4), .b(gate195inter3), .O(gate195inter5));
  nor2  gate699(.a(gate195inter5), .b(gate195inter2), .O(gate195inter6));
  inv1  gate700(.a(N97), .O(gate195inter7));
  inv1  gate701(.a(N716), .O(gate195inter8));
  nand2 gate702(.a(gate195inter8), .b(gate195inter7), .O(gate195inter9));
  nand2 gate703(.a(s_71), .b(gate195inter3), .O(gate195inter10));
  nor2  gate704(.a(gate195inter10), .b(gate195inter9), .O(gate195inter11));
  nor2  gate705(.a(gate195inter11), .b(gate195inter6), .O(gate195inter12));
  nand2 gate706(.a(gate195inter12), .b(gate195inter1), .O(N748));

  xor2  gate399(.a(N717), .b(N101), .O(gate196inter0));
  nand2 gate400(.a(gate196inter0), .b(s_28), .O(gate196inter1));
  and2  gate401(.a(N717), .b(N101), .O(gate196inter2));
  inv1  gate402(.a(s_28), .O(gate196inter3));
  inv1  gate403(.a(s_29), .O(gate196inter4));
  nand2 gate404(.a(gate196inter4), .b(gate196inter3), .O(gate196inter5));
  nor2  gate405(.a(gate196inter5), .b(gate196inter2), .O(gate196inter6));
  inv1  gate406(.a(N101), .O(gate196inter7));
  inv1  gate407(.a(N717), .O(gate196inter8));
  nand2 gate408(.a(gate196inter8), .b(gate196inter7), .O(gate196inter9));
  nand2 gate409(.a(s_29), .b(gate196inter3), .O(gate196inter10));
  nor2  gate410(.a(gate196inter10), .b(gate196inter9), .O(gate196inter11));
  nor2  gate411(.a(gate196inter11), .b(gate196inter6), .O(gate196inter12));
  nand2 gate412(.a(gate196inter12), .b(gate196inter1), .O(N749));

  xor2  gate287(.a(N718), .b(N105), .O(gate197inter0));
  nand2 gate288(.a(gate197inter0), .b(s_12), .O(gate197inter1));
  and2  gate289(.a(N718), .b(N105), .O(gate197inter2));
  inv1  gate290(.a(s_12), .O(gate197inter3));
  inv1  gate291(.a(s_13), .O(gate197inter4));
  nand2 gate292(.a(gate197inter4), .b(gate197inter3), .O(gate197inter5));
  nor2  gate293(.a(gate197inter5), .b(gate197inter2), .O(gate197inter6));
  inv1  gate294(.a(N105), .O(gate197inter7));
  inv1  gate295(.a(N718), .O(gate197inter8));
  nand2 gate296(.a(gate197inter8), .b(gate197inter7), .O(gate197inter9));
  nand2 gate297(.a(s_13), .b(gate197inter3), .O(gate197inter10));
  nor2  gate298(.a(gate197inter10), .b(gate197inter9), .O(gate197inter11));
  nor2  gate299(.a(gate197inter11), .b(gate197inter6), .O(gate197inter12));
  nand2 gate300(.a(gate197inter12), .b(gate197inter1), .O(N750));

  xor2  gate371(.a(N719), .b(N109), .O(gate198inter0));
  nand2 gate372(.a(gate198inter0), .b(s_24), .O(gate198inter1));
  and2  gate373(.a(N719), .b(N109), .O(gate198inter2));
  inv1  gate374(.a(s_24), .O(gate198inter3));
  inv1  gate375(.a(s_25), .O(gate198inter4));
  nand2 gate376(.a(gate198inter4), .b(gate198inter3), .O(gate198inter5));
  nor2  gate377(.a(gate198inter5), .b(gate198inter2), .O(gate198inter6));
  inv1  gate378(.a(N109), .O(gate198inter7));
  inv1  gate379(.a(N719), .O(gate198inter8));
  nand2 gate380(.a(gate198inter8), .b(gate198inter7), .O(gate198inter9));
  nand2 gate381(.a(s_25), .b(gate198inter3), .O(gate198inter10));
  nor2  gate382(.a(gate198inter10), .b(gate198inter9), .O(gate198inter11));
  nor2  gate383(.a(gate198inter11), .b(gate198inter6), .O(gate198inter12));
  nand2 gate384(.a(gate198inter12), .b(gate198inter1), .O(N751));

  xor2  gate469(.a(N720), .b(N113), .O(gate199inter0));
  nand2 gate470(.a(gate199inter0), .b(s_38), .O(gate199inter1));
  and2  gate471(.a(N720), .b(N113), .O(gate199inter2));
  inv1  gate472(.a(s_38), .O(gate199inter3));
  inv1  gate473(.a(s_39), .O(gate199inter4));
  nand2 gate474(.a(gate199inter4), .b(gate199inter3), .O(gate199inter5));
  nor2  gate475(.a(gate199inter5), .b(gate199inter2), .O(gate199inter6));
  inv1  gate476(.a(N113), .O(gate199inter7));
  inv1  gate477(.a(N720), .O(gate199inter8));
  nand2 gate478(.a(gate199inter8), .b(gate199inter7), .O(gate199inter9));
  nand2 gate479(.a(s_39), .b(gate199inter3), .O(gate199inter10));
  nor2  gate480(.a(gate199inter10), .b(gate199inter9), .O(gate199inter11));
  nor2  gate481(.a(gate199inter11), .b(gate199inter6), .O(gate199inter12));
  nand2 gate482(.a(gate199inter12), .b(gate199inter1), .O(N752));

  xor2  gate497(.a(N721), .b(N117), .O(gate200inter0));
  nand2 gate498(.a(gate200inter0), .b(s_42), .O(gate200inter1));
  and2  gate499(.a(N721), .b(N117), .O(gate200inter2));
  inv1  gate500(.a(s_42), .O(gate200inter3));
  inv1  gate501(.a(s_43), .O(gate200inter4));
  nand2 gate502(.a(gate200inter4), .b(gate200inter3), .O(gate200inter5));
  nor2  gate503(.a(gate200inter5), .b(gate200inter2), .O(gate200inter6));
  inv1  gate504(.a(N117), .O(gate200inter7));
  inv1  gate505(.a(N721), .O(gate200inter8));
  nand2 gate506(.a(gate200inter8), .b(gate200inter7), .O(gate200inter9));
  nand2 gate507(.a(s_43), .b(gate200inter3), .O(gate200inter10));
  nor2  gate508(.a(gate200inter10), .b(gate200inter9), .O(gate200inter11));
  nor2  gate509(.a(gate200inter11), .b(gate200inter6), .O(gate200inter12));
  nand2 gate510(.a(gate200inter12), .b(gate200inter1), .O(N753));
xor2 gate201( .a(N121), .b(N722), .O(N754) );

  xor2  gate455(.a(N723), .b(N125), .O(gate202inter0));
  nand2 gate456(.a(gate202inter0), .b(s_36), .O(gate202inter1));
  and2  gate457(.a(N723), .b(N125), .O(gate202inter2));
  inv1  gate458(.a(s_36), .O(gate202inter3));
  inv1  gate459(.a(s_37), .O(gate202inter4));
  nand2 gate460(.a(gate202inter4), .b(gate202inter3), .O(gate202inter5));
  nor2  gate461(.a(gate202inter5), .b(gate202inter2), .O(gate202inter6));
  inv1  gate462(.a(N125), .O(gate202inter7));
  inv1  gate463(.a(N723), .O(gate202inter8));
  nand2 gate464(.a(gate202inter8), .b(gate202inter7), .O(gate202inter9));
  nand2 gate465(.a(s_37), .b(gate202inter3), .O(gate202inter10));
  nor2  gate466(.a(gate202inter10), .b(gate202inter9), .O(gate202inter11));
  nor2  gate467(.a(gate202inter11), .b(gate202inter6), .O(gate202inter12));
  nand2 gate468(.a(gate202inter12), .b(gate202inter1), .O(N755));

endmodule