module c432 (N1,N4,N8,N11,N14,N17,N21,N24,N27,N30,
             N34,N37,N40,N43,N47,N50,N53,N56,N60,N63,
             N66,N69,N73,N76,N79,N82,N86,N89,N92,N95,
             N99,N102,N105,N108,N112,N115,N223,N329,N370,N421,
             N430,N431,N432);

input N1,N4,N8,N11,N14,N17,N21,N24,N27,N30,
      N34,N37,N40,N43,N47,N50,N53,N56,N60,N63,
      N66,N69,N73,N76,N79,N82,N86,N89,N92,N95,
      N99,N102,N105,N108,N112,N115;//RE__PI;

input s_0,s_1;//RE__ALLOW(00,01,10,11);
input s_2,s_3;//RE__ALLOW(00,01,10,11);
input s_4,s_5;//RE__ALLOW(00,01,10,11);
input s_6,s_7;//RE__ALLOW(00,01,10,11);
input s_8,s_9;//RE__ALLOW(00,01,10,11);
input s_10,s_11;//RE__ALLOW(00,01,10,11);
input s_12,s_13;//RE__ALLOW(00,01,10,11);
input s_14,s_15;//RE__ALLOW(00,01,10,11);
input s_16,s_17;//RE__ALLOW(00,01,10,11);
input s_18,s_19;//RE__ALLOW(00,01,10,11);
input s_20,s_21;//RE__ALLOW(00,01,10,11);
input s_22,s_23;//RE__ALLOW(00,01,10,11);
input s_24,s_25;//RE__ALLOW(00,01,10,11);
input s_26,s_27;//RE__ALLOW(00,01,10,11);
input s_28,s_29;//RE__ALLOW(00,01,10,11);
input s_30,s_31;//RE__ALLOW(00,01,10,11);
input s_32,s_33;//RE__ALLOW(00,01,10,11);
input s_34,s_35;//RE__ALLOW(00,01,10,11);
input s_36,s_37;//RE__ALLOW(00,01,10,11);
input s_38,s_39;//RE__ALLOW(00,01,10,11);
input s_40,s_41;//RE__ALLOW(00,01,10,11);
input s_42,s_43;//RE__ALLOW(00,01,10,11);
input s_44,s_45;//RE__ALLOW(00,01,10,11);
input s_46,s_47;//RE__ALLOW(00,01,10,11);
input s_48,s_49;//RE__ALLOW(00,01,10,11);
input s_50,s_51;//RE__ALLOW(00,01,10,11);
input s_52,s_53;//RE__ALLOW(00,01,10,11);
input s_54,s_55;//RE__ALLOW(00,01,10,11);
input s_56,s_57;//RE__ALLOW(00,01,10,11);
input s_58,s_59;//RE__ALLOW(00,01,10,11);
input s_60,s_61;//RE__ALLOW(00,01,10,11);
input s_62,s_63;//RE__ALLOW(00,01,10,11);
input s_64,s_65;//RE__ALLOW(00,01,10,11);
input s_66,s_67;//RE__ALLOW(00,01,10,11);
input s_68,s_69;//RE__ALLOW(00,01,10,11);
input s_70,s_71;//RE__ALLOW(00,01,10,11);
output N223,N329,N370,N421,N430,N431,N432;

wire N118,N119,N122,N123,N126,N127,N130,N131,N134,N135,
     N138,N139,N142,N143,N146,N147,N150,N151,N154,N157,
     N158,N159,N162,N165,N168,N171,N174,N177,N180,N183,
     N184,N185,N186,N187,N188,N189,N190,N191,N192,N193,
     N194,N195,N196,N197,N198,N199,N203,N213,N224,N227,
     N230,N233,N236,N239,N242,N243,N246,N247,N250,N251,
     N254,N255,N256,N257,N258,N259,N260,N263,N264,N267,
     N270,N273,N276,N279,N282,N285,N288,N289,N290,N291,
     N292,N293,N294,N295,N296,N300,N301,N302,N303,N304,
     N305,N306,N307,N308,N309,N319,N330,N331,N332,N333,
     N334,N335,N336,N337,N338,N339,N340,N341,N342,N343,
     N344,N345,N346,N347,N348,N349,N350,N351,N352,N353,
     N354,N355,N356,N357,N360,N371,N372,N373,N374,N375,
     N376,N377,N378,N379,N380,N381,N386,N393,N399,N404,
     N407,N411,N414,N415,N416,N417,N418,N419,N420,N422,
     N425,N428,N429, gate67inter0, gate67inter1, gate67inter2, gate67inter3, gate67inter4, gate67inter5, gate67inter6, gate67inter7, gate67inter8, gate67inter9, gate67inter10, gate67inter11, gate67inter12, gate134inter0, gate134inter1, gate134inter2, gate134inter3, gate134inter4, gate134inter5, gate134inter6, gate134inter7, gate134inter8, gate134inter9, gate134inter10, gate134inter11, gate134inter12, gate113inter0, gate113inter1, gate113inter2, gate113inter3, gate113inter4, gate113inter5, gate113inter6, gate113inter7, gate113inter8, gate113inter9, gate113inter10, gate113inter11, gate113inter12, gate71inter0, gate71inter1, gate71inter2, gate71inter3, gate71inter4, gate71inter5, gate71inter6, gate71inter7, gate71inter8, gate71inter9, gate71inter10, gate71inter11, gate71inter12, gate78inter0, gate78inter1, gate78inter2, gate78inter3, gate78inter4, gate78inter5, gate78inter6, gate78inter7, gate78inter8, gate78inter9, gate78inter10, gate78inter11, gate78inter12, gate19inter0, gate19inter1, gate19inter2, gate19inter3, gate19inter4, gate19inter5, gate19inter6, gate19inter7, gate19inter8, gate19inter9, gate19inter10, gate19inter11, gate19inter12, gate69inter0, gate69inter1, gate69inter2, gate69inter3, gate69inter4, gate69inter5, gate69inter6, gate69inter7, gate69inter8, gate69inter9, gate69inter10, gate69inter11, gate69inter12, gate121inter0, gate121inter1, gate121inter2, gate121inter3, gate121inter4, gate121inter5, gate121inter6, gate121inter7, gate121inter8, gate121inter9, gate121inter10, gate121inter11, gate121inter12, gate41inter0, gate41inter1, gate41inter2, gate41inter3, gate41inter4, gate41inter5, gate41inter6, gate41inter7, gate41inter8, gate41inter9, gate41inter10, gate41inter11, gate41inter12, gate116inter0, gate116inter1, gate116inter2, gate116inter3, gate116inter4, gate116inter5, gate116inter6, gate116inter7, gate116inter8, gate116inter9, gate116inter10, gate116inter11, gate116inter12, gate37inter0, gate37inter1, gate37inter2, gate37inter3, gate37inter4, gate37inter5, gate37inter6, gate37inter7, gate37inter8, gate37inter9, gate37inter10, gate37inter11, gate37inter12, gate29inter0, gate29inter1, gate29inter2, gate29inter3, gate29inter4, gate29inter5, gate29inter6, gate29inter7, gate29inter8, gate29inter9, gate29inter10, gate29inter11, gate29inter12, gate107inter0, gate107inter1, gate107inter2, gate107inter3, gate107inter4, gate107inter5, gate107inter6, gate107inter7, gate107inter8, gate107inter9, gate107inter10, gate107inter11, gate107inter12, gate103inter0, gate103inter1, gate103inter2, gate103inter3, gate103inter4, gate103inter5, gate103inter6, gate103inter7, gate103inter8, gate103inter9, gate103inter10, gate103inter11, gate103inter12, gate44inter0, gate44inter1, gate44inter2, gate44inter3, gate44inter4, gate44inter5, gate44inter6, gate44inter7, gate44inter8, gate44inter9, gate44inter10, gate44inter11, gate44inter12, gate39inter0, gate39inter1, gate39inter2, gate39inter3, gate39inter4, gate39inter5, gate39inter6, gate39inter7, gate39inter8, gate39inter9, gate39inter10, gate39inter11, gate39inter12, gate108inter0, gate108inter1, gate108inter2, gate108inter3, gate108inter4, gate108inter5, gate108inter6, gate108inter7, gate108inter8, gate108inter9, gate108inter10, gate108inter11, gate108inter12, gate119inter0, gate119inter1, gate119inter2, gate119inter3, gate119inter4, gate119inter5, gate119inter6, gate119inter7, gate119inter8, gate119inter9, gate119inter10, gate119inter11, gate119inter12, gate60inter0, gate60inter1, gate60inter2, gate60inter3, gate60inter4, gate60inter5, gate60inter6, gate60inter7, gate60inter8, gate60inter9, gate60inter10, gate60inter11, gate60inter12, gate136inter0, gate136inter1, gate136inter2, gate136inter3, gate136inter4, gate136inter5, gate136inter6, gate136inter7, gate136inter8, gate136inter9, gate136inter10, gate136inter11, gate136inter12, gate24inter0, gate24inter1, gate24inter2, gate24inter3, gate24inter4, gate24inter5, gate24inter6, gate24inter7, gate24inter8, gate24inter9, gate24inter10, gate24inter11, gate24inter12, gate133inter0, gate133inter1, gate133inter2, gate133inter3, gate133inter4, gate133inter5, gate133inter6, gate133inter7, gate133inter8, gate133inter9, gate133inter10, gate133inter11, gate133inter12, gate51inter0, gate51inter1, gate51inter2, gate51inter3, gate51inter4, gate51inter5, gate51inter6, gate51inter7, gate51inter8, gate51inter9, gate51inter10, gate51inter11, gate51inter12, gate137inter0, gate137inter1, gate137inter2, gate137inter3, gate137inter4, gate137inter5, gate137inter6, gate137inter7, gate137inter8, gate137inter9, gate137inter10, gate137inter11, gate137inter12, gate35inter0, gate35inter1, gate35inter2, gate35inter3, gate35inter4, gate35inter5, gate35inter6, gate35inter7, gate35inter8, gate35inter9, gate35inter10, gate35inter11, gate35inter12, gate122inter0, gate122inter1, gate122inter2, gate122inter3, gate122inter4, gate122inter5, gate122inter6, gate122inter7, gate122inter8, gate122inter9, gate122inter10, gate122inter11, gate122inter12, gate130inter0, gate130inter1, gate130inter2, gate130inter3, gate130inter4, gate130inter5, gate130inter6, gate130inter7, gate130inter8, gate130inter9, gate130inter10, gate130inter11, gate130inter12, gate54inter0, gate54inter1, gate54inter2, gate54inter3, gate54inter4, gate54inter5, gate54inter6, gate54inter7, gate54inter8, gate54inter9, gate54inter10, gate54inter11, gate54inter12, gate20inter0, gate20inter1, gate20inter2, gate20inter3, gate20inter4, gate20inter5, gate20inter6, gate20inter7, gate20inter8, gate20inter9, gate20inter10, gate20inter11, gate20inter12, gate50inter0, gate50inter1, gate50inter2, gate50inter3, gate50inter4, gate50inter5, gate50inter6, gate50inter7, gate50inter8, gate50inter9, gate50inter10, gate50inter11, gate50inter12, gate115inter0, gate115inter1, gate115inter2, gate115inter3, gate115inter4, gate115inter5, gate115inter6, gate115inter7, gate115inter8, gate115inter9, gate115inter10, gate115inter11, gate115inter12, gate34inter0, gate34inter1, gate34inter2, gate34inter3, gate34inter4, gate34inter5, gate34inter6, gate34inter7, gate34inter8, gate34inter9, gate34inter10, gate34inter11, gate34inter12, gate59inter0, gate59inter1, gate59inter2, gate59inter3, gate59inter4, gate59inter5, gate59inter6, gate59inter7, gate59inter8, gate59inter9, gate59inter10, gate59inter11, gate59inter12, gate109inter0, gate109inter1, gate109inter2, gate109inter3, gate109inter4, gate109inter5, gate109inter6, gate109inter7, gate109inter8, gate109inter9, gate109inter10, gate109inter11, gate109inter12, gate64inter0, gate64inter1, gate64inter2, gate64inter3, gate64inter4, gate64inter5, gate64inter6, gate64inter7, gate64inter8, gate64inter9, gate64inter10, gate64inter11, gate64inter12, gate40inter0, gate40inter1, gate40inter2, gate40inter3, gate40inter4, gate40inter5, gate40inter6, gate40inter7, gate40inter8, gate40inter9, gate40inter10, gate40inter11, gate40inter12;



inv1 gate1( .a(N1), .O(N118) );
inv1 gate2( .a(N4), .O(N119) );
inv1 gate3( .a(N11), .O(N122) );
inv1 gate4( .a(N17), .O(N123) );
inv1 gate5( .a(N24), .O(N126) );
inv1 gate6( .a(N30), .O(N127) );
inv1 gate7( .a(N37), .O(N130) );
inv1 gate8( .a(N43), .O(N131) );
inv1 gate9( .a(N50), .O(N134) );
inv1 gate10( .a(N56), .O(N135) );
inv1 gate11( .a(N63), .O(N138) );
inv1 gate12( .a(N69), .O(N139) );
inv1 gate13( .a(N76), .O(N142) );
inv1 gate14( .a(N82), .O(N143) );
inv1 gate15( .a(N89), .O(N146) );
inv1 gate16( .a(N95), .O(N147) );
inv1 gate17( .a(N102), .O(N150) );
inv1 gate18( .a(N108), .O(N151) );

  xor2  gate231(.a(N4), .b(N118), .O(gate19inter0));
  nand2 gate232(.a(gate19inter0), .b(s_10), .O(gate19inter1));
  and2  gate233(.a(N4), .b(N118), .O(gate19inter2));
  inv1  gate234(.a(s_10), .O(gate19inter3));
  inv1  gate235(.a(s_11), .O(gate19inter4));
  nand2 gate236(.a(gate19inter4), .b(gate19inter3), .O(gate19inter5));
  nor2  gate237(.a(gate19inter5), .b(gate19inter2), .O(gate19inter6));
  inv1  gate238(.a(N118), .O(gate19inter7));
  inv1  gate239(.a(N4), .O(gate19inter8));
  nand2 gate240(.a(gate19inter8), .b(gate19inter7), .O(gate19inter9));
  nand2 gate241(.a(s_11), .b(gate19inter3), .O(gate19inter10));
  nor2  gate242(.a(gate19inter10), .b(gate19inter9), .O(gate19inter11));
  nor2  gate243(.a(gate19inter11), .b(gate19inter6), .O(gate19inter12));
  nand2 gate244(.a(gate19inter12), .b(gate19inter1), .O(N154));

  xor2  gate553(.a(N119), .b(N8), .O(gate20inter0));
  nand2 gate554(.a(gate20inter0), .b(s_56), .O(gate20inter1));
  and2  gate555(.a(N119), .b(N8), .O(gate20inter2));
  inv1  gate556(.a(s_56), .O(gate20inter3));
  inv1  gate557(.a(s_57), .O(gate20inter4));
  nand2 gate558(.a(gate20inter4), .b(gate20inter3), .O(gate20inter5));
  nor2  gate559(.a(gate20inter5), .b(gate20inter2), .O(gate20inter6));
  inv1  gate560(.a(N8), .O(gate20inter7));
  inv1  gate561(.a(N119), .O(gate20inter8));
  nand2 gate562(.a(gate20inter8), .b(gate20inter7), .O(gate20inter9));
  nand2 gate563(.a(s_57), .b(gate20inter3), .O(gate20inter10));
  nor2  gate564(.a(gate20inter10), .b(gate20inter9), .O(gate20inter11));
  nor2  gate565(.a(gate20inter11), .b(gate20inter6), .O(gate20inter12));
  nand2 gate566(.a(gate20inter12), .b(gate20inter1), .O(N157));
nor2 gate21( .a(N14), .b(N119), .O(N158) );
nand2 gate22( .a(N122), .b(N17), .O(N159) );
nand2 gate23( .a(N126), .b(N30), .O(N162) );

  xor2  gate441(.a(N43), .b(N130), .O(gate24inter0));
  nand2 gate442(.a(gate24inter0), .b(s_40), .O(gate24inter1));
  and2  gate443(.a(N43), .b(N130), .O(gate24inter2));
  inv1  gate444(.a(s_40), .O(gate24inter3));
  inv1  gate445(.a(s_41), .O(gate24inter4));
  nand2 gate446(.a(gate24inter4), .b(gate24inter3), .O(gate24inter5));
  nor2  gate447(.a(gate24inter5), .b(gate24inter2), .O(gate24inter6));
  inv1  gate448(.a(N130), .O(gate24inter7));
  inv1  gate449(.a(N43), .O(gate24inter8));
  nand2 gate450(.a(gate24inter8), .b(gate24inter7), .O(gate24inter9));
  nand2 gate451(.a(s_41), .b(gate24inter3), .O(gate24inter10));
  nor2  gate452(.a(gate24inter10), .b(gate24inter9), .O(gate24inter11));
  nor2  gate453(.a(gate24inter11), .b(gate24inter6), .O(gate24inter12));
  nand2 gate454(.a(gate24inter12), .b(gate24inter1), .O(N165));
nand2 gate25( .a(N134), .b(N56), .O(N168) );
nand2 gate26( .a(N138), .b(N69), .O(N171) );
nand2 gate27( .a(N142), .b(N82), .O(N174) );
nand2 gate28( .a(N146), .b(N95), .O(N177) );

  xor2  gate315(.a(N108), .b(N150), .O(gate29inter0));
  nand2 gate316(.a(gate29inter0), .b(s_22), .O(gate29inter1));
  and2  gate317(.a(N108), .b(N150), .O(gate29inter2));
  inv1  gate318(.a(s_22), .O(gate29inter3));
  inv1  gate319(.a(s_23), .O(gate29inter4));
  nand2 gate320(.a(gate29inter4), .b(gate29inter3), .O(gate29inter5));
  nor2  gate321(.a(gate29inter5), .b(gate29inter2), .O(gate29inter6));
  inv1  gate322(.a(N150), .O(gate29inter7));
  inv1  gate323(.a(N108), .O(gate29inter8));
  nand2 gate324(.a(gate29inter8), .b(gate29inter7), .O(gate29inter9));
  nand2 gate325(.a(s_23), .b(gate29inter3), .O(gate29inter10));
  nor2  gate326(.a(gate29inter10), .b(gate29inter9), .O(gate29inter11));
  nor2  gate327(.a(gate29inter11), .b(gate29inter6), .O(gate29inter12));
  nand2 gate328(.a(gate29inter12), .b(gate29inter1), .O(N180));
nor2 gate30( .a(N21), .b(N123), .O(N183) );
nor2 gate31( .a(N27), .b(N123), .O(N184) );
nor2 gate32( .a(N34), .b(N127), .O(N185) );
nor2 gate33( .a(N40), .b(N127), .O(N186) );

  xor2  gate595(.a(N131), .b(N47), .O(gate34inter0));
  nand2 gate596(.a(gate34inter0), .b(s_62), .O(gate34inter1));
  and2  gate597(.a(N131), .b(N47), .O(gate34inter2));
  inv1  gate598(.a(s_62), .O(gate34inter3));
  inv1  gate599(.a(s_63), .O(gate34inter4));
  nand2 gate600(.a(gate34inter4), .b(gate34inter3), .O(gate34inter5));
  nor2  gate601(.a(gate34inter5), .b(gate34inter2), .O(gate34inter6));
  inv1  gate602(.a(N47), .O(gate34inter7));
  inv1  gate603(.a(N131), .O(gate34inter8));
  nand2 gate604(.a(gate34inter8), .b(gate34inter7), .O(gate34inter9));
  nand2 gate605(.a(s_63), .b(gate34inter3), .O(gate34inter10));
  nor2  gate606(.a(gate34inter10), .b(gate34inter9), .O(gate34inter11));
  nor2  gate607(.a(gate34inter11), .b(gate34inter6), .O(gate34inter12));
  nand2 gate608(.a(gate34inter12), .b(gate34inter1), .O(N187));

  xor2  gate497(.a(N131), .b(N53), .O(gate35inter0));
  nand2 gate498(.a(gate35inter0), .b(s_48), .O(gate35inter1));
  and2  gate499(.a(N131), .b(N53), .O(gate35inter2));
  inv1  gate500(.a(s_48), .O(gate35inter3));
  inv1  gate501(.a(s_49), .O(gate35inter4));
  nand2 gate502(.a(gate35inter4), .b(gate35inter3), .O(gate35inter5));
  nor2  gate503(.a(gate35inter5), .b(gate35inter2), .O(gate35inter6));
  inv1  gate504(.a(N53), .O(gate35inter7));
  inv1  gate505(.a(N131), .O(gate35inter8));
  nand2 gate506(.a(gate35inter8), .b(gate35inter7), .O(gate35inter9));
  nand2 gate507(.a(s_49), .b(gate35inter3), .O(gate35inter10));
  nor2  gate508(.a(gate35inter10), .b(gate35inter9), .O(gate35inter11));
  nor2  gate509(.a(gate35inter11), .b(gate35inter6), .O(gate35inter12));
  nand2 gate510(.a(gate35inter12), .b(gate35inter1), .O(N188));
nor2 gate36( .a(N60), .b(N135), .O(N189) );

  xor2  gate301(.a(N135), .b(N66), .O(gate37inter0));
  nand2 gate302(.a(gate37inter0), .b(s_20), .O(gate37inter1));
  and2  gate303(.a(N135), .b(N66), .O(gate37inter2));
  inv1  gate304(.a(s_20), .O(gate37inter3));
  inv1  gate305(.a(s_21), .O(gate37inter4));
  nand2 gate306(.a(gate37inter4), .b(gate37inter3), .O(gate37inter5));
  nor2  gate307(.a(gate37inter5), .b(gate37inter2), .O(gate37inter6));
  inv1  gate308(.a(N66), .O(gate37inter7));
  inv1  gate309(.a(N135), .O(gate37inter8));
  nand2 gate310(.a(gate37inter8), .b(gate37inter7), .O(gate37inter9));
  nand2 gate311(.a(s_21), .b(gate37inter3), .O(gate37inter10));
  nor2  gate312(.a(gate37inter10), .b(gate37inter9), .O(gate37inter11));
  nor2  gate313(.a(gate37inter11), .b(gate37inter6), .O(gate37inter12));
  nand2 gate314(.a(gate37inter12), .b(gate37inter1), .O(N190));
nor2 gate38( .a(N73), .b(N139), .O(N191) );

  xor2  gate371(.a(N139), .b(N79), .O(gate39inter0));
  nand2 gate372(.a(gate39inter0), .b(s_30), .O(gate39inter1));
  and2  gate373(.a(N139), .b(N79), .O(gate39inter2));
  inv1  gate374(.a(s_30), .O(gate39inter3));
  inv1  gate375(.a(s_31), .O(gate39inter4));
  nand2 gate376(.a(gate39inter4), .b(gate39inter3), .O(gate39inter5));
  nor2  gate377(.a(gate39inter5), .b(gate39inter2), .O(gate39inter6));
  inv1  gate378(.a(N79), .O(gate39inter7));
  inv1  gate379(.a(N139), .O(gate39inter8));
  nand2 gate380(.a(gate39inter8), .b(gate39inter7), .O(gate39inter9));
  nand2 gate381(.a(s_31), .b(gate39inter3), .O(gate39inter10));
  nor2  gate382(.a(gate39inter10), .b(gate39inter9), .O(gate39inter11));
  nor2  gate383(.a(gate39inter11), .b(gate39inter6), .O(gate39inter12));
  nand2 gate384(.a(gate39inter12), .b(gate39inter1), .O(N192));

  xor2  gate651(.a(N143), .b(N86), .O(gate40inter0));
  nand2 gate652(.a(gate40inter0), .b(s_70), .O(gate40inter1));
  and2  gate653(.a(N143), .b(N86), .O(gate40inter2));
  inv1  gate654(.a(s_70), .O(gate40inter3));
  inv1  gate655(.a(s_71), .O(gate40inter4));
  nand2 gate656(.a(gate40inter4), .b(gate40inter3), .O(gate40inter5));
  nor2  gate657(.a(gate40inter5), .b(gate40inter2), .O(gate40inter6));
  inv1  gate658(.a(N86), .O(gate40inter7));
  inv1  gate659(.a(N143), .O(gate40inter8));
  nand2 gate660(.a(gate40inter8), .b(gate40inter7), .O(gate40inter9));
  nand2 gate661(.a(s_71), .b(gate40inter3), .O(gate40inter10));
  nor2  gate662(.a(gate40inter10), .b(gate40inter9), .O(gate40inter11));
  nor2  gate663(.a(gate40inter11), .b(gate40inter6), .O(gate40inter12));
  nand2 gate664(.a(gate40inter12), .b(gate40inter1), .O(N193));

  xor2  gate273(.a(N143), .b(N92), .O(gate41inter0));
  nand2 gate274(.a(gate41inter0), .b(s_16), .O(gate41inter1));
  and2  gate275(.a(N143), .b(N92), .O(gate41inter2));
  inv1  gate276(.a(s_16), .O(gate41inter3));
  inv1  gate277(.a(s_17), .O(gate41inter4));
  nand2 gate278(.a(gate41inter4), .b(gate41inter3), .O(gate41inter5));
  nor2  gate279(.a(gate41inter5), .b(gate41inter2), .O(gate41inter6));
  inv1  gate280(.a(N92), .O(gate41inter7));
  inv1  gate281(.a(N143), .O(gate41inter8));
  nand2 gate282(.a(gate41inter8), .b(gate41inter7), .O(gate41inter9));
  nand2 gate283(.a(s_17), .b(gate41inter3), .O(gate41inter10));
  nor2  gate284(.a(gate41inter10), .b(gate41inter9), .O(gate41inter11));
  nor2  gate285(.a(gate41inter11), .b(gate41inter6), .O(gate41inter12));
  nand2 gate286(.a(gate41inter12), .b(gate41inter1), .O(N194));
nor2 gate42( .a(N99), .b(N147), .O(N195) );
nor2 gate43( .a(N105), .b(N147), .O(N196) );

  xor2  gate357(.a(N151), .b(N112), .O(gate44inter0));
  nand2 gate358(.a(gate44inter0), .b(s_28), .O(gate44inter1));
  and2  gate359(.a(N151), .b(N112), .O(gate44inter2));
  inv1  gate360(.a(s_28), .O(gate44inter3));
  inv1  gate361(.a(s_29), .O(gate44inter4));
  nand2 gate362(.a(gate44inter4), .b(gate44inter3), .O(gate44inter5));
  nor2  gate363(.a(gate44inter5), .b(gate44inter2), .O(gate44inter6));
  inv1  gate364(.a(N112), .O(gate44inter7));
  inv1  gate365(.a(N151), .O(gate44inter8));
  nand2 gate366(.a(gate44inter8), .b(gate44inter7), .O(gate44inter9));
  nand2 gate367(.a(s_29), .b(gate44inter3), .O(gate44inter10));
  nor2  gate368(.a(gate44inter10), .b(gate44inter9), .O(gate44inter11));
  nor2  gate369(.a(gate44inter11), .b(gate44inter6), .O(gate44inter12));
  nand2 gate370(.a(gate44inter12), .b(gate44inter1), .O(N197));
nor2 gate45( .a(N115), .b(N151), .O(N198) );
and9 gate46( .a(N154), .b(N159), .c(N162), .d(N165), .e(N168), .f(N171), .g(N174), .h(N177), .i(N180), .O(N199) );
inv1 gate47( .a(N199), .O(N203) );
inv1 gate48( .a(N199), .O(N213) );
inv1 gate49( .a(N199), .O(N223) );

  xor2  gate567(.a(N154), .b(N203), .O(gate50inter0));
  nand2 gate568(.a(gate50inter0), .b(s_58), .O(gate50inter1));
  and2  gate569(.a(N154), .b(N203), .O(gate50inter2));
  inv1  gate570(.a(s_58), .O(gate50inter3));
  inv1  gate571(.a(s_59), .O(gate50inter4));
  nand2 gate572(.a(gate50inter4), .b(gate50inter3), .O(gate50inter5));
  nor2  gate573(.a(gate50inter5), .b(gate50inter2), .O(gate50inter6));
  inv1  gate574(.a(N203), .O(gate50inter7));
  inv1  gate575(.a(N154), .O(gate50inter8));
  nand2 gate576(.a(gate50inter8), .b(gate50inter7), .O(gate50inter9));
  nand2 gate577(.a(s_59), .b(gate50inter3), .O(gate50inter10));
  nor2  gate578(.a(gate50inter10), .b(gate50inter9), .O(gate50inter11));
  nor2  gate579(.a(gate50inter11), .b(gate50inter6), .O(gate50inter12));
  nand2 gate580(.a(gate50inter12), .b(gate50inter1), .O(N224));

  xor2  gate469(.a(N159), .b(N203), .O(gate51inter0));
  nand2 gate470(.a(gate51inter0), .b(s_44), .O(gate51inter1));
  and2  gate471(.a(N159), .b(N203), .O(gate51inter2));
  inv1  gate472(.a(s_44), .O(gate51inter3));
  inv1  gate473(.a(s_45), .O(gate51inter4));
  nand2 gate474(.a(gate51inter4), .b(gate51inter3), .O(gate51inter5));
  nor2  gate475(.a(gate51inter5), .b(gate51inter2), .O(gate51inter6));
  inv1  gate476(.a(N203), .O(gate51inter7));
  inv1  gate477(.a(N159), .O(gate51inter8));
  nand2 gate478(.a(gate51inter8), .b(gate51inter7), .O(gate51inter9));
  nand2 gate479(.a(s_45), .b(gate51inter3), .O(gate51inter10));
  nor2  gate480(.a(gate51inter10), .b(gate51inter9), .O(gate51inter11));
  nor2  gate481(.a(gate51inter11), .b(gate51inter6), .O(gate51inter12));
  nand2 gate482(.a(gate51inter12), .b(gate51inter1), .O(N227));
xor2 gate52( .a(N203), .b(N162), .O(N230) );
xor2 gate53( .a(N203), .b(N165), .O(N233) );

  xor2  gate539(.a(N168), .b(N203), .O(gate54inter0));
  nand2 gate540(.a(gate54inter0), .b(s_54), .O(gate54inter1));
  and2  gate541(.a(N168), .b(N203), .O(gate54inter2));
  inv1  gate542(.a(s_54), .O(gate54inter3));
  inv1  gate543(.a(s_55), .O(gate54inter4));
  nand2 gate544(.a(gate54inter4), .b(gate54inter3), .O(gate54inter5));
  nor2  gate545(.a(gate54inter5), .b(gate54inter2), .O(gate54inter6));
  inv1  gate546(.a(N203), .O(gate54inter7));
  inv1  gate547(.a(N168), .O(gate54inter8));
  nand2 gate548(.a(gate54inter8), .b(gate54inter7), .O(gate54inter9));
  nand2 gate549(.a(s_55), .b(gate54inter3), .O(gate54inter10));
  nor2  gate550(.a(gate54inter10), .b(gate54inter9), .O(gate54inter11));
  nor2  gate551(.a(gate54inter11), .b(gate54inter6), .O(gate54inter12));
  nand2 gate552(.a(gate54inter12), .b(gate54inter1), .O(N236));
xor2 gate55( .a(N203), .b(N171), .O(N239) );
nand2 gate56( .a(N1), .b(N213), .O(N242) );
xor2 gate57( .a(N203), .b(N174), .O(N243) );
nand2 gate58( .a(N213), .b(N11), .O(N246) );

  xor2  gate609(.a(N177), .b(N203), .O(gate59inter0));
  nand2 gate610(.a(gate59inter0), .b(s_64), .O(gate59inter1));
  and2  gate611(.a(N177), .b(N203), .O(gate59inter2));
  inv1  gate612(.a(s_64), .O(gate59inter3));
  inv1  gate613(.a(s_65), .O(gate59inter4));
  nand2 gate614(.a(gate59inter4), .b(gate59inter3), .O(gate59inter5));
  nor2  gate615(.a(gate59inter5), .b(gate59inter2), .O(gate59inter6));
  inv1  gate616(.a(N203), .O(gate59inter7));
  inv1  gate617(.a(N177), .O(gate59inter8));
  nand2 gate618(.a(gate59inter8), .b(gate59inter7), .O(gate59inter9));
  nand2 gate619(.a(s_65), .b(gate59inter3), .O(gate59inter10));
  nor2  gate620(.a(gate59inter10), .b(gate59inter9), .O(gate59inter11));
  nor2  gate621(.a(gate59inter11), .b(gate59inter6), .O(gate59inter12));
  nand2 gate622(.a(gate59inter12), .b(gate59inter1), .O(N247));

  xor2  gate413(.a(N24), .b(N213), .O(gate60inter0));
  nand2 gate414(.a(gate60inter0), .b(s_36), .O(gate60inter1));
  and2  gate415(.a(N24), .b(N213), .O(gate60inter2));
  inv1  gate416(.a(s_36), .O(gate60inter3));
  inv1  gate417(.a(s_37), .O(gate60inter4));
  nand2 gate418(.a(gate60inter4), .b(gate60inter3), .O(gate60inter5));
  nor2  gate419(.a(gate60inter5), .b(gate60inter2), .O(gate60inter6));
  inv1  gate420(.a(N213), .O(gate60inter7));
  inv1  gate421(.a(N24), .O(gate60inter8));
  nand2 gate422(.a(gate60inter8), .b(gate60inter7), .O(gate60inter9));
  nand2 gate423(.a(s_37), .b(gate60inter3), .O(gate60inter10));
  nor2  gate424(.a(gate60inter10), .b(gate60inter9), .O(gate60inter11));
  nor2  gate425(.a(gate60inter11), .b(gate60inter6), .O(gate60inter12));
  nand2 gate426(.a(gate60inter12), .b(gate60inter1), .O(N250));
xor2 gate61( .a(N203), .b(N180), .O(N251) );
nand2 gate62( .a(N213), .b(N37), .O(N254) );
nand2 gate63( .a(N213), .b(N50), .O(N255) );

  xor2  gate637(.a(N63), .b(N213), .O(gate64inter0));
  nand2 gate638(.a(gate64inter0), .b(s_68), .O(gate64inter1));
  and2  gate639(.a(N63), .b(N213), .O(gate64inter2));
  inv1  gate640(.a(s_68), .O(gate64inter3));
  inv1  gate641(.a(s_69), .O(gate64inter4));
  nand2 gate642(.a(gate64inter4), .b(gate64inter3), .O(gate64inter5));
  nor2  gate643(.a(gate64inter5), .b(gate64inter2), .O(gate64inter6));
  inv1  gate644(.a(N213), .O(gate64inter7));
  inv1  gate645(.a(N63), .O(gate64inter8));
  nand2 gate646(.a(gate64inter8), .b(gate64inter7), .O(gate64inter9));
  nand2 gate647(.a(s_69), .b(gate64inter3), .O(gate64inter10));
  nor2  gate648(.a(gate64inter10), .b(gate64inter9), .O(gate64inter11));
  nor2  gate649(.a(gate64inter11), .b(gate64inter6), .O(gate64inter12));
  nand2 gate650(.a(gate64inter12), .b(gate64inter1), .O(N256));
nand2 gate65( .a(N213), .b(N76), .O(N257) );
nand2 gate66( .a(N213), .b(N89), .O(N258) );

  xor2  gate161(.a(N102), .b(N213), .O(gate67inter0));
  nand2 gate162(.a(gate67inter0), .b(s_0), .O(gate67inter1));
  and2  gate163(.a(N102), .b(N213), .O(gate67inter2));
  inv1  gate164(.a(s_0), .O(gate67inter3));
  inv1  gate165(.a(s_1), .O(gate67inter4));
  nand2 gate166(.a(gate67inter4), .b(gate67inter3), .O(gate67inter5));
  nor2  gate167(.a(gate67inter5), .b(gate67inter2), .O(gate67inter6));
  inv1  gate168(.a(N213), .O(gate67inter7));
  inv1  gate169(.a(N102), .O(gate67inter8));
  nand2 gate170(.a(gate67inter8), .b(gate67inter7), .O(gate67inter9));
  nand2 gate171(.a(s_1), .b(gate67inter3), .O(gate67inter10));
  nor2  gate172(.a(gate67inter10), .b(gate67inter9), .O(gate67inter11));
  nor2  gate173(.a(gate67inter11), .b(gate67inter6), .O(gate67inter12));
  nand2 gate174(.a(gate67inter12), .b(gate67inter1), .O(N259));
nand2 gate68( .a(N224), .b(N157), .O(N260) );

  xor2  gate245(.a(N158), .b(N224), .O(gate69inter0));
  nand2 gate246(.a(gate69inter0), .b(s_12), .O(gate69inter1));
  and2  gate247(.a(N158), .b(N224), .O(gate69inter2));
  inv1  gate248(.a(s_12), .O(gate69inter3));
  inv1  gate249(.a(s_13), .O(gate69inter4));
  nand2 gate250(.a(gate69inter4), .b(gate69inter3), .O(gate69inter5));
  nor2  gate251(.a(gate69inter5), .b(gate69inter2), .O(gate69inter6));
  inv1  gate252(.a(N224), .O(gate69inter7));
  inv1  gate253(.a(N158), .O(gate69inter8));
  nand2 gate254(.a(gate69inter8), .b(gate69inter7), .O(gate69inter9));
  nand2 gate255(.a(s_13), .b(gate69inter3), .O(gate69inter10));
  nor2  gate256(.a(gate69inter10), .b(gate69inter9), .O(gate69inter11));
  nor2  gate257(.a(gate69inter11), .b(gate69inter6), .O(gate69inter12));
  nand2 gate258(.a(gate69inter12), .b(gate69inter1), .O(N263));
nand2 gate70( .a(N227), .b(N183), .O(N264) );

  xor2  gate203(.a(N185), .b(N230), .O(gate71inter0));
  nand2 gate204(.a(gate71inter0), .b(s_6), .O(gate71inter1));
  and2  gate205(.a(N185), .b(N230), .O(gate71inter2));
  inv1  gate206(.a(s_6), .O(gate71inter3));
  inv1  gate207(.a(s_7), .O(gate71inter4));
  nand2 gate208(.a(gate71inter4), .b(gate71inter3), .O(gate71inter5));
  nor2  gate209(.a(gate71inter5), .b(gate71inter2), .O(gate71inter6));
  inv1  gate210(.a(N230), .O(gate71inter7));
  inv1  gate211(.a(N185), .O(gate71inter8));
  nand2 gate212(.a(gate71inter8), .b(gate71inter7), .O(gate71inter9));
  nand2 gate213(.a(s_7), .b(gate71inter3), .O(gate71inter10));
  nor2  gate214(.a(gate71inter10), .b(gate71inter9), .O(gate71inter11));
  nor2  gate215(.a(gate71inter11), .b(gate71inter6), .O(gate71inter12));
  nand2 gate216(.a(gate71inter12), .b(gate71inter1), .O(N267));
nand2 gate72( .a(N233), .b(N187), .O(N270) );
nand2 gate73( .a(N236), .b(N189), .O(N273) );
nand2 gate74( .a(N239), .b(N191), .O(N276) );
nand2 gate75( .a(N243), .b(N193), .O(N279) );
nand2 gate76( .a(N247), .b(N195), .O(N282) );
nand2 gate77( .a(N251), .b(N197), .O(N285) );

  xor2  gate217(.a(N184), .b(N227), .O(gate78inter0));
  nand2 gate218(.a(gate78inter0), .b(s_8), .O(gate78inter1));
  and2  gate219(.a(N184), .b(N227), .O(gate78inter2));
  inv1  gate220(.a(s_8), .O(gate78inter3));
  inv1  gate221(.a(s_9), .O(gate78inter4));
  nand2 gate222(.a(gate78inter4), .b(gate78inter3), .O(gate78inter5));
  nor2  gate223(.a(gate78inter5), .b(gate78inter2), .O(gate78inter6));
  inv1  gate224(.a(N227), .O(gate78inter7));
  inv1  gate225(.a(N184), .O(gate78inter8));
  nand2 gate226(.a(gate78inter8), .b(gate78inter7), .O(gate78inter9));
  nand2 gate227(.a(s_9), .b(gate78inter3), .O(gate78inter10));
  nor2  gate228(.a(gate78inter10), .b(gate78inter9), .O(gate78inter11));
  nor2  gate229(.a(gate78inter11), .b(gate78inter6), .O(gate78inter12));
  nand2 gate230(.a(gate78inter12), .b(gate78inter1), .O(N288));
nand2 gate79( .a(N230), .b(N186), .O(N289) );
nand2 gate80( .a(N233), .b(N188), .O(N290) );
nand2 gate81( .a(N236), .b(N190), .O(N291) );
nand2 gate82( .a(N239), .b(N192), .O(N292) );
nand2 gate83( .a(N243), .b(N194), .O(N293) );
nand2 gate84( .a(N247), .b(N196), .O(N294) );
nand2 gate85( .a(N251), .b(N198), .O(N295) );
and9 gate86( .a(N260), .b(N264), .c(N267), .d(N270), .e(N273), .f(N276), .g(N279), .h(N282), .i(N285), .O(N296) );
inv1 gate87( .a(N263), .O(N300) );
inv1 gate88( .a(N288), .O(N301) );
inv1 gate89( .a(N289), .O(N302) );
inv1 gate90( .a(N290), .O(N303) );
inv1 gate91( .a(N291), .O(N304) );
inv1 gate92( .a(N292), .O(N305) );
inv1 gate93( .a(N293), .O(N306) );
inv1 gate94( .a(N294), .O(N307) );
inv1 gate95( .a(N295), .O(N308) );
inv1 gate96( .a(N296), .O(N309) );
inv1 gate97( .a(N296), .O(N319) );
inv1 gate98( .a(N296), .O(N329) );
xor2 gate99( .a(N309), .b(N260), .O(N330) );
xor2 gate100( .a(N309), .b(N264), .O(N331) );
xor2 gate101( .a(N309), .b(N267), .O(N332) );
xor2 gate102( .a(N309), .b(N270), .O(N333) );

  xor2  gate343(.a(N319), .b(N8), .O(gate103inter0));
  nand2 gate344(.a(gate103inter0), .b(s_26), .O(gate103inter1));
  and2  gate345(.a(N319), .b(N8), .O(gate103inter2));
  inv1  gate346(.a(s_26), .O(gate103inter3));
  inv1  gate347(.a(s_27), .O(gate103inter4));
  nand2 gate348(.a(gate103inter4), .b(gate103inter3), .O(gate103inter5));
  nor2  gate349(.a(gate103inter5), .b(gate103inter2), .O(gate103inter6));
  inv1  gate350(.a(N8), .O(gate103inter7));
  inv1  gate351(.a(N319), .O(gate103inter8));
  nand2 gate352(.a(gate103inter8), .b(gate103inter7), .O(gate103inter9));
  nand2 gate353(.a(s_27), .b(gate103inter3), .O(gate103inter10));
  nor2  gate354(.a(gate103inter10), .b(gate103inter9), .O(gate103inter11));
  nor2  gate355(.a(gate103inter11), .b(gate103inter6), .O(gate103inter12));
  nand2 gate356(.a(gate103inter12), .b(gate103inter1), .O(N334));
xor2 gate104( .a(N309), .b(N273), .O(N335) );
nand2 gate105( .a(N319), .b(N21), .O(N336) );
xor2 gate106( .a(N309), .b(N276), .O(N337) );

  xor2  gate329(.a(N34), .b(N319), .O(gate107inter0));
  nand2 gate330(.a(gate107inter0), .b(s_24), .O(gate107inter1));
  and2  gate331(.a(N34), .b(N319), .O(gate107inter2));
  inv1  gate332(.a(s_24), .O(gate107inter3));
  inv1  gate333(.a(s_25), .O(gate107inter4));
  nand2 gate334(.a(gate107inter4), .b(gate107inter3), .O(gate107inter5));
  nor2  gate335(.a(gate107inter5), .b(gate107inter2), .O(gate107inter6));
  inv1  gate336(.a(N319), .O(gate107inter7));
  inv1  gate337(.a(N34), .O(gate107inter8));
  nand2 gate338(.a(gate107inter8), .b(gate107inter7), .O(gate107inter9));
  nand2 gate339(.a(s_25), .b(gate107inter3), .O(gate107inter10));
  nor2  gate340(.a(gate107inter10), .b(gate107inter9), .O(gate107inter11));
  nor2  gate341(.a(gate107inter11), .b(gate107inter6), .O(gate107inter12));
  nand2 gate342(.a(gate107inter12), .b(gate107inter1), .O(N338));

  xor2  gate385(.a(N279), .b(N309), .O(gate108inter0));
  nand2 gate386(.a(gate108inter0), .b(s_32), .O(gate108inter1));
  and2  gate387(.a(N279), .b(N309), .O(gate108inter2));
  inv1  gate388(.a(s_32), .O(gate108inter3));
  inv1  gate389(.a(s_33), .O(gate108inter4));
  nand2 gate390(.a(gate108inter4), .b(gate108inter3), .O(gate108inter5));
  nor2  gate391(.a(gate108inter5), .b(gate108inter2), .O(gate108inter6));
  inv1  gate392(.a(N309), .O(gate108inter7));
  inv1  gate393(.a(N279), .O(gate108inter8));
  nand2 gate394(.a(gate108inter8), .b(gate108inter7), .O(gate108inter9));
  nand2 gate395(.a(s_33), .b(gate108inter3), .O(gate108inter10));
  nor2  gate396(.a(gate108inter10), .b(gate108inter9), .O(gate108inter11));
  nor2  gate397(.a(gate108inter11), .b(gate108inter6), .O(gate108inter12));
  nand2 gate398(.a(gate108inter12), .b(gate108inter1), .O(N339));

  xor2  gate623(.a(N47), .b(N319), .O(gate109inter0));
  nand2 gate624(.a(gate109inter0), .b(s_66), .O(gate109inter1));
  and2  gate625(.a(N47), .b(N319), .O(gate109inter2));
  inv1  gate626(.a(s_66), .O(gate109inter3));
  inv1  gate627(.a(s_67), .O(gate109inter4));
  nand2 gate628(.a(gate109inter4), .b(gate109inter3), .O(gate109inter5));
  nor2  gate629(.a(gate109inter5), .b(gate109inter2), .O(gate109inter6));
  inv1  gate630(.a(N319), .O(gate109inter7));
  inv1  gate631(.a(N47), .O(gate109inter8));
  nand2 gate632(.a(gate109inter8), .b(gate109inter7), .O(gate109inter9));
  nand2 gate633(.a(s_67), .b(gate109inter3), .O(gate109inter10));
  nor2  gate634(.a(gate109inter10), .b(gate109inter9), .O(gate109inter11));
  nor2  gate635(.a(gate109inter11), .b(gate109inter6), .O(gate109inter12));
  nand2 gate636(.a(gate109inter12), .b(gate109inter1), .O(N340));
xor2 gate110( .a(N309), .b(N282), .O(N341) );
nand2 gate111( .a(N319), .b(N60), .O(N342) );
xor2 gate112( .a(N309), .b(N285), .O(N343) );

  xor2  gate189(.a(N73), .b(N319), .O(gate113inter0));
  nand2 gate190(.a(gate113inter0), .b(s_4), .O(gate113inter1));
  and2  gate191(.a(N73), .b(N319), .O(gate113inter2));
  inv1  gate192(.a(s_4), .O(gate113inter3));
  inv1  gate193(.a(s_5), .O(gate113inter4));
  nand2 gate194(.a(gate113inter4), .b(gate113inter3), .O(gate113inter5));
  nor2  gate195(.a(gate113inter5), .b(gate113inter2), .O(gate113inter6));
  inv1  gate196(.a(N319), .O(gate113inter7));
  inv1  gate197(.a(N73), .O(gate113inter8));
  nand2 gate198(.a(gate113inter8), .b(gate113inter7), .O(gate113inter9));
  nand2 gate199(.a(s_5), .b(gate113inter3), .O(gate113inter10));
  nor2  gate200(.a(gate113inter10), .b(gate113inter9), .O(gate113inter11));
  nor2  gate201(.a(gate113inter11), .b(gate113inter6), .O(gate113inter12));
  nand2 gate202(.a(gate113inter12), .b(gate113inter1), .O(N344));
nand2 gate114( .a(N319), .b(N86), .O(N345) );

  xor2  gate581(.a(N99), .b(N319), .O(gate115inter0));
  nand2 gate582(.a(gate115inter0), .b(s_60), .O(gate115inter1));
  and2  gate583(.a(N99), .b(N319), .O(gate115inter2));
  inv1  gate584(.a(s_60), .O(gate115inter3));
  inv1  gate585(.a(s_61), .O(gate115inter4));
  nand2 gate586(.a(gate115inter4), .b(gate115inter3), .O(gate115inter5));
  nor2  gate587(.a(gate115inter5), .b(gate115inter2), .O(gate115inter6));
  inv1  gate588(.a(N319), .O(gate115inter7));
  inv1  gate589(.a(N99), .O(gate115inter8));
  nand2 gate590(.a(gate115inter8), .b(gate115inter7), .O(gate115inter9));
  nand2 gate591(.a(s_61), .b(gate115inter3), .O(gate115inter10));
  nor2  gate592(.a(gate115inter10), .b(gate115inter9), .O(gate115inter11));
  nor2  gate593(.a(gate115inter11), .b(gate115inter6), .O(gate115inter12));
  nand2 gate594(.a(gate115inter12), .b(gate115inter1), .O(N346));

  xor2  gate287(.a(N112), .b(N319), .O(gate116inter0));
  nand2 gate288(.a(gate116inter0), .b(s_18), .O(gate116inter1));
  and2  gate289(.a(N112), .b(N319), .O(gate116inter2));
  inv1  gate290(.a(s_18), .O(gate116inter3));
  inv1  gate291(.a(s_19), .O(gate116inter4));
  nand2 gate292(.a(gate116inter4), .b(gate116inter3), .O(gate116inter5));
  nor2  gate293(.a(gate116inter5), .b(gate116inter2), .O(gate116inter6));
  inv1  gate294(.a(N319), .O(gate116inter7));
  inv1  gate295(.a(N112), .O(gate116inter8));
  nand2 gate296(.a(gate116inter8), .b(gate116inter7), .O(gate116inter9));
  nand2 gate297(.a(s_19), .b(gate116inter3), .O(gate116inter10));
  nor2  gate298(.a(gate116inter10), .b(gate116inter9), .O(gate116inter11));
  nor2  gate299(.a(gate116inter11), .b(gate116inter6), .O(gate116inter12));
  nand2 gate300(.a(gate116inter12), .b(gate116inter1), .O(N347));
nand2 gate117( .a(N330), .b(N300), .O(N348) );
nand2 gate118( .a(N331), .b(N301), .O(N349) );

  xor2  gate399(.a(N302), .b(N332), .O(gate119inter0));
  nand2 gate400(.a(gate119inter0), .b(s_34), .O(gate119inter1));
  and2  gate401(.a(N302), .b(N332), .O(gate119inter2));
  inv1  gate402(.a(s_34), .O(gate119inter3));
  inv1  gate403(.a(s_35), .O(gate119inter4));
  nand2 gate404(.a(gate119inter4), .b(gate119inter3), .O(gate119inter5));
  nor2  gate405(.a(gate119inter5), .b(gate119inter2), .O(gate119inter6));
  inv1  gate406(.a(N332), .O(gate119inter7));
  inv1  gate407(.a(N302), .O(gate119inter8));
  nand2 gate408(.a(gate119inter8), .b(gate119inter7), .O(gate119inter9));
  nand2 gate409(.a(s_35), .b(gate119inter3), .O(gate119inter10));
  nor2  gate410(.a(gate119inter10), .b(gate119inter9), .O(gate119inter11));
  nor2  gate411(.a(gate119inter11), .b(gate119inter6), .O(gate119inter12));
  nand2 gate412(.a(gate119inter12), .b(gate119inter1), .O(N350));
nand2 gate120( .a(N333), .b(N303), .O(N351) );

  xor2  gate259(.a(N304), .b(N335), .O(gate121inter0));
  nand2 gate260(.a(gate121inter0), .b(s_14), .O(gate121inter1));
  and2  gate261(.a(N304), .b(N335), .O(gate121inter2));
  inv1  gate262(.a(s_14), .O(gate121inter3));
  inv1  gate263(.a(s_15), .O(gate121inter4));
  nand2 gate264(.a(gate121inter4), .b(gate121inter3), .O(gate121inter5));
  nor2  gate265(.a(gate121inter5), .b(gate121inter2), .O(gate121inter6));
  inv1  gate266(.a(N335), .O(gate121inter7));
  inv1  gate267(.a(N304), .O(gate121inter8));
  nand2 gate268(.a(gate121inter8), .b(gate121inter7), .O(gate121inter9));
  nand2 gate269(.a(s_15), .b(gate121inter3), .O(gate121inter10));
  nor2  gate270(.a(gate121inter10), .b(gate121inter9), .O(gate121inter11));
  nor2  gate271(.a(gate121inter11), .b(gate121inter6), .O(gate121inter12));
  nand2 gate272(.a(gate121inter12), .b(gate121inter1), .O(N352));

  xor2  gate511(.a(N305), .b(N337), .O(gate122inter0));
  nand2 gate512(.a(gate122inter0), .b(s_50), .O(gate122inter1));
  and2  gate513(.a(N305), .b(N337), .O(gate122inter2));
  inv1  gate514(.a(s_50), .O(gate122inter3));
  inv1  gate515(.a(s_51), .O(gate122inter4));
  nand2 gate516(.a(gate122inter4), .b(gate122inter3), .O(gate122inter5));
  nor2  gate517(.a(gate122inter5), .b(gate122inter2), .O(gate122inter6));
  inv1  gate518(.a(N337), .O(gate122inter7));
  inv1  gate519(.a(N305), .O(gate122inter8));
  nand2 gate520(.a(gate122inter8), .b(gate122inter7), .O(gate122inter9));
  nand2 gate521(.a(s_51), .b(gate122inter3), .O(gate122inter10));
  nor2  gate522(.a(gate122inter10), .b(gate122inter9), .O(gate122inter11));
  nor2  gate523(.a(gate122inter11), .b(gate122inter6), .O(gate122inter12));
  nand2 gate524(.a(gate122inter12), .b(gate122inter1), .O(N353));
nand2 gate123( .a(N339), .b(N306), .O(N354) );
nand2 gate124( .a(N341), .b(N307), .O(N355) );
nand2 gate125( .a(N343), .b(N308), .O(N356) );
and9 gate126( .a(N348), .b(N349), .c(N350), .d(N351), .e(N352), .f(N353), .g(N354), .h(N355), .i(N356), .O(N357) );
inv1 gate127( .a(N357), .O(N360) );
inv1 gate128( .a(N357), .O(N370) );
nand2 gate129( .a(N14), .b(N360), .O(N371) );

  xor2  gate525(.a(N27), .b(N360), .O(gate130inter0));
  nand2 gate526(.a(gate130inter0), .b(s_52), .O(gate130inter1));
  and2  gate527(.a(N27), .b(N360), .O(gate130inter2));
  inv1  gate528(.a(s_52), .O(gate130inter3));
  inv1  gate529(.a(s_53), .O(gate130inter4));
  nand2 gate530(.a(gate130inter4), .b(gate130inter3), .O(gate130inter5));
  nor2  gate531(.a(gate130inter5), .b(gate130inter2), .O(gate130inter6));
  inv1  gate532(.a(N360), .O(gate130inter7));
  inv1  gate533(.a(N27), .O(gate130inter8));
  nand2 gate534(.a(gate130inter8), .b(gate130inter7), .O(gate130inter9));
  nand2 gate535(.a(s_53), .b(gate130inter3), .O(gate130inter10));
  nor2  gate536(.a(gate130inter10), .b(gate130inter9), .O(gate130inter11));
  nor2  gate537(.a(gate130inter11), .b(gate130inter6), .O(gate130inter12));
  nand2 gate538(.a(gate130inter12), .b(gate130inter1), .O(N372));
nand2 gate131( .a(N360), .b(N40), .O(N373) );
nand2 gate132( .a(N360), .b(N53), .O(N374) );

  xor2  gate455(.a(N66), .b(N360), .O(gate133inter0));
  nand2 gate456(.a(gate133inter0), .b(s_42), .O(gate133inter1));
  and2  gate457(.a(N66), .b(N360), .O(gate133inter2));
  inv1  gate458(.a(s_42), .O(gate133inter3));
  inv1  gate459(.a(s_43), .O(gate133inter4));
  nand2 gate460(.a(gate133inter4), .b(gate133inter3), .O(gate133inter5));
  nor2  gate461(.a(gate133inter5), .b(gate133inter2), .O(gate133inter6));
  inv1  gate462(.a(N360), .O(gate133inter7));
  inv1  gate463(.a(N66), .O(gate133inter8));
  nand2 gate464(.a(gate133inter8), .b(gate133inter7), .O(gate133inter9));
  nand2 gate465(.a(s_43), .b(gate133inter3), .O(gate133inter10));
  nor2  gate466(.a(gate133inter10), .b(gate133inter9), .O(gate133inter11));
  nor2  gate467(.a(gate133inter11), .b(gate133inter6), .O(gate133inter12));
  nand2 gate468(.a(gate133inter12), .b(gate133inter1), .O(N375));

  xor2  gate175(.a(N79), .b(N360), .O(gate134inter0));
  nand2 gate176(.a(gate134inter0), .b(s_2), .O(gate134inter1));
  and2  gate177(.a(N79), .b(N360), .O(gate134inter2));
  inv1  gate178(.a(s_2), .O(gate134inter3));
  inv1  gate179(.a(s_3), .O(gate134inter4));
  nand2 gate180(.a(gate134inter4), .b(gate134inter3), .O(gate134inter5));
  nor2  gate181(.a(gate134inter5), .b(gate134inter2), .O(gate134inter6));
  inv1  gate182(.a(N360), .O(gate134inter7));
  inv1  gate183(.a(N79), .O(gate134inter8));
  nand2 gate184(.a(gate134inter8), .b(gate134inter7), .O(gate134inter9));
  nand2 gate185(.a(s_3), .b(gate134inter3), .O(gate134inter10));
  nor2  gate186(.a(gate134inter10), .b(gate134inter9), .O(gate134inter11));
  nor2  gate187(.a(gate134inter11), .b(gate134inter6), .O(gate134inter12));
  nand2 gate188(.a(gate134inter12), .b(gate134inter1), .O(N376));
nand2 gate135( .a(N360), .b(N92), .O(N377) );

  xor2  gate427(.a(N105), .b(N360), .O(gate136inter0));
  nand2 gate428(.a(gate136inter0), .b(s_38), .O(gate136inter1));
  and2  gate429(.a(N105), .b(N360), .O(gate136inter2));
  inv1  gate430(.a(s_38), .O(gate136inter3));
  inv1  gate431(.a(s_39), .O(gate136inter4));
  nand2 gate432(.a(gate136inter4), .b(gate136inter3), .O(gate136inter5));
  nor2  gate433(.a(gate136inter5), .b(gate136inter2), .O(gate136inter6));
  inv1  gate434(.a(N360), .O(gate136inter7));
  inv1  gate435(.a(N105), .O(gate136inter8));
  nand2 gate436(.a(gate136inter8), .b(gate136inter7), .O(gate136inter9));
  nand2 gate437(.a(s_39), .b(gate136inter3), .O(gate136inter10));
  nor2  gate438(.a(gate136inter10), .b(gate136inter9), .O(gate136inter11));
  nor2  gate439(.a(gate136inter11), .b(gate136inter6), .O(gate136inter12));
  nand2 gate440(.a(gate136inter12), .b(gate136inter1), .O(N378));

  xor2  gate483(.a(N115), .b(N360), .O(gate137inter0));
  nand2 gate484(.a(gate137inter0), .b(s_46), .O(gate137inter1));
  and2  gate485(.a(N115), .b(N360), .O(gate137inter2));
  inv1  gate486(.a(s_46), .O(gate137inter3));
  inv1  gate487(.a(s_47), .O(gate137inter4));
  nand2 gate488(.a(gate137inter4), .b(gate137inter3), .O(gate137inter5));
  nor2  gate489(.a(gate137inter5), .b(gate137inter2), .O(gate137inter6));
  inv1  gate490(.a(N360), .O(gate137inter7));
  inv1  gate491(.a(N115), .O(gate137inter8));
  nand2 gate492(.a(gate137inter8), .b(gate137inter7), .O(gate137inter9));
  nand2 gate493(.a(s_47), .b(gate137inter3), .O(gate137inter10));
  nor2  gate494(.a(gate137inter10), .b(gate137inter9), .O(gate137inter11));
  nor2  gate495(.a(gate137inter11), .b(gate137inter6), .O(gate137inter12));
  nand2 gate496(.a(gate137inter12), .b(gate137inter1), .O(N379));
nand4 gate138( .a(N4), .b(N242), .c(N334), .d(N371), .O(N380) );
nand4 gate139( .a(N246), .b(N336), .c(N372), .d(N17), .O(N381) );
nand4 gate140( .a(N250), .b(N338), .c(N373), .d(N30), .O(N386) );
nand4 gate141( .a(N254), .b(N340), .c(N374), .d(N43), .O(N393) );
nand4 gate142( .a(N255), .b(N342), .c(N375), .d(N56), .O(N399) );
nand4 gate143( .a(N256), .b(N344), .c(N376), .d(N69), .O(N404) );
nand4 gate144( .a(N257), .b(N345), .c(N377), .d(N82), .O(N407) );
nand4 gate145( .a(N258), .b(N346), .c(N378), .d(N95), .O(N411) );
nand4 gate146( .a(N259), .b(N347), .c(N379), .d(N108), .O(N414) );
inv1 gate147( .a(N380), .O(N415) );
and8 gate148( .a(N381), .b(N386), .c(N393), .d(N399), .e(N404), .f(N407), .g(N411), .h(N414), .O(N416) );
inv1 gate149( .a(N393), .O(N417) );
inv1 gate150( .a(N404), .O(N418) );
inv1 gate151( .a(N407), .O(N419) );
inv1 gate152( .a(N411), .O(N420) );
nor2 gate153( .a(N415), .b(N416), .O(N421) );
nand2 gate154( .a(N386), .b(N417), .O(N422) );
nand4 gate155( .a(N386), .b(N393), .c(N418), .d(N399), .O(N425) );
nand3 gate156( .a(N399), .b(N393), .c(N419), .O(N428) );
nand4 gate157( .a(N386), .b(N393), .c(N407), .d(N420), .O(N429) );
nand4 gate158( .a(N381), .b(N386), .c(N422), .d(N399), .O(N430) );
nand4 gate159( .a(N381), .b(N386), .c(N425), .d(N428), .O(N431) );
nand4 gate160( .a(N381), .b(N422), .c(N425), .d(N429), .O(N432) );

endmodule