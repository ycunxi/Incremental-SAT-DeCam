module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);

input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;//RE__PI;

input s_0,s_1;//RE__ALLOW(00,01,10,11);
input s_2,s_3;//RE__ALLOW(00,01,10,11);
input s_4,s_5;//RE__ALLOW(00,01,10,11);
input s_6,s_7;//RE__ALLOW(00,01,10,11);
input s_8,s_9;//RE__ALLOW(00,01,10,11);
input s_10,s_11;//RE__ALLOW(00,01,10,11);
input s_12,s_13;//RE__ALLOW(00,01,10,11);
input s_14,s_15;//RE__ALLOW(00,01,10,11);
input s_16,s_17;//RE__ALLOW(00,01,10,11);
input s_18,s_19;//RE__ALLOW(00,01,10,11);
input s_20,s_21;//RE__ALLOW(00,01,10,11);
input s_22,s_23;//RE__ALLOW(00,01,10,11);
input s_24,s_25;//RE__ALLOW(00,01,10,11);
input s_26,s_27;//RE__ALLOW(00,01,10,11);
input s_28,s_29;//RE__ALLOW(00,01,10,11);
input s_30,s_31;//RE__ALLOW(00,01,10,11);
input s_32,s_33;//RE__ALLOW(00,01,10,11);
input s_34,s_35;//RE__ALLOW(00,01,10,11);
input s_36,s_37;//RE__ALLOW(00,01,10,11);
input s_38,s_39;//RE__ALLOW(00,01,10,11);
input s_40,s_41;//RE__ALLOW(00,01,10,11);
input s_42,s_43;//RE__ALLOW(00,01,10,11);
input s_44,s_45;//RE__ALLOW(00,01,10,11);
input s_46,s_47;//RE__ALLOW(00,01,10,11);
input s_48,s_49;//RE__ALLOW(00,01,10,11);
input s_50,s_51;//RE__ALLOW(00,01,10,11);
input s_52,s_53;//RE__ALLOW(00,01,10,11);
input s_54,s_55;//RE__ALLOW(00,01,10,11);
input s_56,s_57;//RE__ALLOW(00,01,10,11);
input s_58,s_59;//RE__ALLOW(00,01,10,11);
input s_60,s_61;//RE__ALLOW(00,01,10,11);
input s_62,s_63;//RE__ALLOW(00,01,10,11);
input s_64,s_65;//RE__ALLOW(00,01,10,11);
input s_66,s_67;//RE__ALLOW(00,01,10,11);
input s_68,s_69;//RE__ALLOW(00,01,10,11);
input s_70,s_71;//RE__ALLOW(00,01,10,11);
input s_72,s_73;//RE__ALLOW(00,01,10,11);
input s_74,s_75;//RE__ALLOW(00,01,10,11);
input s_76,s_77;//RE__ALLOW(00,01,10,11);
input s_78,s_79;//RE__ALLOW(00,01,10,11);
input s_80,s_81;//RE__ALLOW(00,01,10,11);
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;

  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate63inter0, gate63inter1, gate63inter2, gate63inter3, gate63inter4, gate63inter5, gate63inter6, gate63inter7, gate63inter8, gate63inter9, gate63inter10, gate63inter11, gate63inter12, gate420inter0, gate420inter1, gate420inter2, gate420inter3, gate420inter4, gate420inter5, gate420inter6, gate420inter7, gate420inter8, gate420inter9, gate420inter10, gate420inter11, gate420inter12, gate81inter0, gate81inter1, gate81inter2, gate81inter3, gate81inter4, gate81inter5, gate81inter6, gate81inter7, gate81inter8, gate81inter9, gate81inter10, gate81inter11, gate81inter12, gate188inter0, gate188inter1, gate188inter2, gate188inter3, gate188inter4, gate188inter5, gate188inter6, gate188inter7, gate188inter8, gate188inter9, gate188inter10, gate188inter11, gate188inter12, gate112inter0, gate112inter1, gate112inter2, gate112inter3, gate112inter4, gate112inter5, gate112inter6, gate112inter7, gate112inter8, gate112inter9, gate112inter10, gate112inter11, gate112inter12, gate260inter0, gate260inter1, gate260inter2, gate260inter3, gate260inter4, gate260inter5, gate260inter6, gate260inter7, gate260inter8, gate260inter9, gate260inter10, gate260inter11, gate260inter12, gate237inter0, gate237inter1, gate237inter2, gate237inter3, gate237inter4, gate237inter5, gate237inter6, gate237inter7, gate237inter8, gate237inter9, gate237inter10, gate237inter11, gate237inter12, gate110inter0, gate110inter1, gate110inter2, gate110inter3, gate110inter4, gate110inter5, gate110inter6, gate110inter7, gate110inter8, gate110inter9, gate110inter10, gate110inter11, gate110inter12, gate129inter0, gate129inter1, gate129inter2, gate129inter3, gate129inter4, gate129inter5, gate129inter6, gate129inter7, gate129inter8, gate129inter9, gate129inter10, gate129inter11, gate129inter12, gate134inter0, gate134inter1, gate134inter2, gate134inter3, gate134inter4, gate134inter5, gate134inter6, gate134inter7, gate134inter8, gate134inter9, gate134inter10, gate134inter11, gate134inter12, gate50inter0, gate50inter1, gate50inter2, gate50inter3, gate50inter4, gate50inter5, gate50inter6, gate50inter7, gate50inter8, gate50inter9, gate50inter10, gate50inter11, gate50inter12, gate34inter0, gate34inter1, gate34inter2, gate34inter3, gate34inter4, gate34inter5, gate34inter6, gate34inter7, gate34inter8, gate34inter9, gate34inter10, gate34inter11, gate34inter12, gate265inter0, gate265inter1, gate265inter2, gate265inter3, gate265inter4, gate265inter5, gate265inter6, gate265inter7, gate265inter8, gate265inter9, gate265inter10, gate265inter11, gate265inter12, gate36inter0, gate36inter1, gate36inter2, gate36inter3, gate36inter4, gate36inter5, gate36inter6, gate36inter7, gate36inter8, gate36inter9, gate36inter10, gate36inter11, gate36inter12, gate409inter0, gate409inter1, gate409inter2, gate409inter3, gate409inter4, gate409inter5, gate409inter6, gate409inter7, gate409inter8, gate409inter9, gate409inter10, gate409inter11, gate409inter12, gate119inter0, gate119inter1, gate119inter2, gate119inter3, gate119inter4, gate119inter5, gate119inter6, gate119inter7, gate119inter8, gate119inter9, gate119inter10, gate119inter11, gate119inter12, gate219inter0, gate219inter1, gate219inter2, gate219inter3, gate219inter4, gate219inter5, gate219inter6, gate219inter7, gate219inter8, gate219inter9, gate219inter10, gate219inter11, gate219inter12, gate121inter0, gate121inter1, gate121inter2, gate121inter3, gate121inter4, gate121inter5, gate121inter6, gate121inter7, gate121inter8, gate121inter9, gate121inter10, gate121inter11, gate121inter12, gate91inter0, gate91inter1, gate91inter2, gate91inter3, gate91inter4, gate91inter5, gate91inter6, gate91inter7, gate91inter8, gate91inter9, gate91inter10, gate91inter11, gate91inter12, gate225inter0, gate225inter1, gate225inter2, gate225inter3, gate225inter4, gate225inter5, gate225inter6, gate225inter7, gate225inter8, gate225inter9, gate225inter10, gate225inter11, gate225inter12, gate150inter0, gate150inter1, gate150inter2, gate150inter3, gate150inter4, gate150inter5, gate150inter6, gate150inter7, gate150inter8, gate150inter9, gate150inter10, gate150inter11, gate150inter12, gate42inter0, gate42inter1, gate42inter2, gate42inter3, gate42inter4, gate42inter5, gate42inter6, gate42inter7, gate42inter8, gate42inter9, gate42inter10, gate42inter11, gate42inter12, gate29inter0, gate29inter1, gate29inter2, gate29inter3, gate29inter4, gate29inter5, gate29inter6, gate29inter7, gate29inter8, gate29inter9, gate29inter10, gate29inter11, gate29inter12, gate13inter0, gate13inter1, gate13inter2, gate13inter3, gate13inter4, gate13inter5, gate13inter6, gate13inter7, gate13inter8, gate13inter9, gate13inter10, gate13inter11, gate13inter12, gate198inter0, gate198inter1, gate198inter2, gate198inter3, gate198inter4, gate198inter5, gate198inter6, gate198inter7, gate198inter8, gate198inter9, gate198inter10, gate198inter11, gate198inter12, gate20inter0, gate20inter1, gate20inter2, gate20inter3, gate20inter4, gate20inter5, gate20inter6, gate20inter7, gate20inter8, gate20inter9, gate20inter10, gate20inter11, gate20inter12, gate457inter0, gate457inter1, gate457inter2, gate457inter3, gate457inter4, gate457inter5, gate457inter6, gate457inter7, gate457inter8, gate457inter9, gate457inter10, gate457inter11, gate457inter12, gate170inter0, gate170inter1, gate170inter2, gate170inter3, gate170inter4, gate170inter5, gate170inter6, gate170inter7, gate170inter8, gate170inter9, gate170inter10, gate170inter11, gate170inter12, gate228inter0, gate228inter1, gate228inter2, gate228inter3, gate228inter4, gate228inter5, gate228inter6, gate228inter7, gate228inter8, gate228inter9, gate228inter10, gate228inter11, gate228inter12, gate100inter0, gate100inter1, gate100inter2, gate100inter3, gate100inter4, gate100inter5, gate100inter6, gate100inter7, gate100inter8, gate100inter9, gate100inter10, gate100inter11, gate100inter12, gate78inter0, gate78inter1, gate78inter2, gate78inter3, gate78inter4, gate78inter5, gate78inter6, gate78inter7, gate78inter8, gate78inter9, gate78inter10, gate78inter11, gate78inter12, gate396inter0, gate396inter1, gate396inter2, gate396inter3, gate396inter4, gate396inter5, gate396inter6, gate396inter7, gate396inter8, gate396inter9, gate396inter10, gate396inter11, gate396inter12, gate270inter0, gate270inter1, gate270inter2, gate270inter3, gate270inter4, gate270inter5, gate270inter6, gate270inter7, gate270inter8, gate270inter9, gate270inter10, gate270inter11, gate270inter12, gate505inter0, gate505inter1, gate505inter2, gate505inter3, gate505inter4, gate505inter5, gate505inter6, gate505inter7, gate505inter8, gate505inter9, gate505inter10, gate505inter11, gate505inter12, gate469inter0, gate469inter1, gate469inter2, gate469inter3, gate469inter4, gate469inter5, gate469inter6, gate469inter7, gate469inter8, gate469inter9, gate469inter10, gate469inter11, gate469inter12, gate64inter0, gate64inter1, gate64inter2, gate64inter3, gate64inter4, gate64inter5, gate64inter6, gate64inter7, gate64inter8, gate64inter9, gate64inter10, gate64inter11, gate64inter12, gate54inter0, gate54inter1, gate54inter2, gate54inter3, gate54inter4, gate54inter5, gate54inter6, gate54inter7, gate54inter8, gate54inter9, gate54inter10, gate54inter11, gate54inter12, gate468inter0, gate468inter1, gate468inter2, gate468inter3, gate468inter4, gate468inter5, gate468inter6, gate468inter7, gate468inter8, gate468inter9, gate468inter10, gate468inter11, gate468inter12, gate58inter0, gate58inter1, gate58inter2, gate58inter3, gate58inter4, gate58inter5, gate58inter6, gate58inter7, gate58inter8, gate58inter9, gate58inter10, gate58inter11, gate58inter12, gate111inter0, gate111inter1, gate111inter2, gate111inter3, gate111inter4, gate111inter5, gate111inter6, gate111inter7, gate111inter8, gate111inter9, gate111inter10, gate111inter11, gate111inter12, gate441inter0, gate441inter1, gate441inter2, gate441inter3, gate441inter4, gate441inter5, gate441inter6, gate441inter7, gate441inter8, gate441inter9, gate441inter10, gate441inter11, gate441inter12;



and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );
nand2 gate9( .a(G1), .b(G2), .O(G266) );
nand2 gate10( .a(G3), .b(G4), .O(G269) );
nand2 gate11( .a(G5), .b(G6), .O(G272) );
nand2 gate12( .a(G7), .b(G8), .O(G275) );

  xor2  gate869(.a(G10), .b(G9), .O(gate13inter0));
  nand2 gate870(.a(gate13inter0), .b(s_46), .O(gate13inter1));
  and2  gate871(.a(G10), .b(G9), .O(gate13inter2));
  inv1  gate872(.a(s_46), .O(gate13inter3));
  inv1  gate873(.a(s_47), .O(gate13inter4));
  nand2 gate874(.a(gate13inter4), .b(gate13inter3), .O(gate13inter5));
  nor2  gate875(.a(gate13inter5), .b(gate13inter2), .O(gate13inter6));
  inv1  gate876(.a(G9), .O(gate13inter7));
  inv1  gate877(.a(G10), .O(gate13inter8));
  nand2 gate878(.a(gate13inter8), .b(gate13inter7), .O(gate13inter9));
  nand2 gate879(.a(s_47), .b(gate13inter3), .O(gate13inter10));
  nor2  gate880(.a(gate13inter10), .b(gate13inter9), .O(gate13inter11));
  nor2  gate881(.a(gate13inter11), .b(gate13inter6), .O(gate13inter12));
  nand2 gate882(.a(gate13inter12), .b(gate13inter1), .O(G278));
nand2 gate14( .a(G11), .b(G12), .O(G281) );
nand2 gate15( .a(G13), .b(G14), .O(G284) );
nand2 gate16( .a(G15), .b(G16), .O(G287) );
nand2 gate17( .a(G17), .b(G18), .O(G290) );
nand2 gate18( .a(G19), .b(G20), .O(G293) );
nand2 gate19( .a(G21), .b(G22), .O(G296) );

  xor2  gate897(.a(G24), .b(G23), .O(gate20inter0));
  nand2 gate898(.a(gate20inter0), .b(s_50), .O(gate20inter1));
  and2  gate899(.a(G24), .b(G23), .O(gate20inter2));
  inv1  gate900(.a(s_50), .O(gate20inter3));
  inv1  gate901(.a(s_51), .O(gate20inter4));
  nand2 gate902(.a(gate20inter4), .b(gate20inter3), .O(gate20inter5));
  nor2  gate903(.a(gate20inter5), .b(gate20inter2), .O(gate20inter6));
  inv1  gate904(.a(G23), .O(gate20inter7));
  inv1  gate905(.a(G24), .O(gate20inter8));
  nand2 gate906(.a(gate20inter8), .b(gate20inter7), .O(gate20inter9));
  nand2 gate907(.a(s_51), .b(gate20inter3), .O(gate20inter10));
  nor2  gate908(.a(gate20inter10), .b(gate20inter9), .O(gate20inter11));
  nor2  gate909(.a(gate20inter11), .b(gate20inter6), .O(gate20inter12));
  nand2 gate910(.a(gate20inter12), .b(gate20inter1), .O(G299));
nand2 gate21( .a(G25), .b(G26), .O(G302) );
nand2 gate22( .a(G27), .b(G28), .O(G305) );
nand2 gate23( .a(G29), .b(G30), .O(G308) );
nand2 gate24( .a(G31), .b(G32), .O(G311) );
nand2 gate25( .a(G1), .b(G5), .O(G314) );
nand2 gate26( .a(G9), .b(G13), .O(G317) );
nand2 gate27( .a(G2), .b(G6), .O(G320) );
nand2 gate28( .a(G10), .b(G14), .O(G323) );

  xor2  gate855(.a(G7), .b(G3), .O(gate29inter0));
  nand2 gate856(.a(gate29inter0), .b(s_44), .O(gate29inter1));
  and2  gate857(.a(G7), .b(G3), .O(gate29inter2));
  inv1  gate858(.a(s_44), .O(gate29inter3));
  inv1  gate859(.a(s_45), .O(gate29inter4));
  nand2 gate860(.a(gate29inter4), .b(gate29inter3), .O(gate29inter5));
  nor2  gate861(.a(gate29inter5), .b(gate29inter2), .O(gate29inter6));
  inv1  gate862(.a(G3), .O(gate29inter7));
  inv1  gate863(.a(G7), .O(gate29inter8));
  nand2 gate864(.a(gate29inter8), .b(gate29inter7), .O(gate29inter9));
  nand2 gate865(.a(s_45), .b(gate29inter3), .O(gate29inter10));
  nor2  gate866(.a(gate29inter10), .b(gate29inter9), .O(gate29inter11));
  nor2  gate867(.a(gate29inter11), .b(gate29inter6), .O(gate29inter12));
  nand2 gate868(.a(gate29inter12), .b(gate29inter1), .O(G326));
nand2 gate30( .a(G11), .b(G15), .O(G329) );
nand2 gate31( .a(G4), .b(G8), .O(G332) );
nand2 gate32( .a(G12), .b(G16), .O(G335) );
nand2 gate33( .a(G17), .b(G21), .O(G338) );

  xor2  gate701(.a(G29), .b(G25), .O(gate34inter0));
  nand2 gate702(.a(gate34inter0), .b(s_22), .O(gate34inter1));
  and2  gate703(.a(G29), .b(G25), .O(gate34inter2));
  inv1  gate704(.a(s_22), .O(gate34inter3));
  inv1  gate705(.a(s_23), .O(gate34inter4));
  nand2 gate706(.a(gate34inter4), .b(gate34inter3), .O(gate34inter5));
  nor2  gate707(.a(gate34inter5), .b(gate34inter2), .O(gate34inter6));
  inv1  gate708(.a(G25), .O(gate34inter7));
  inv1  gate709(.a(G29), .O(gate34inter8));
  nand2 gate710(.a(gate34inter8), .b(gate34inter7), .O(gate34inter9));
  nand2 gate711(.a(s_23), .b(gate34inter3), .O(gate34inter10));
  nor2  gate712(.a(gate34inter10), .b(gate34inter9), .O(gate34inter11));
  nor2  gate713(.a(gate34inter11), .b(gate34inter6), .O(gate34inter12));
  nand2 gate714(.a(gate34inter12), .b(gate34inter1), .O(G341));
nand2 gate35( .a(G18), .b(G22), .O(G344) );

  xor2  gate729(.a(G30), .b(G26), .O(gate36inter0));
  nand2 gate730(.a(gate36inter0), .b(s_26), .O(gate36inter1));
  and2  gate731(.a(G30), .b(G26), .O(gate36inter2));
  inv1  gate732(.a(s_26), .O(gate36inter3));
  inv1  gate733(.a(s_27), .O(gate36inter4));
  nand2 gate734(.a(gate36inter4), .b(gate36inter3), .O(gate36inter5));
  nor2  gate735(.a(gate36inter5), .b(gate36inter2), .O(gate36inter6));
  inv1  gate736(.a(G26), .O(gate36inter7));
  inv1  gate737(.a(G30), .O(gate36inter8));
  nand2 gate738(.a(gate36inter8), .b(gate36inter7), .O(gate36inter9));
  nand2 gate739(.a(s_27), .b(gate36inter3), .O(gate36inter10));
  nor2  gate740(.a(gate36inter10), .b(gate36inter9), .O(gate36inter11));
  nor2  gate741(.a(gate36inter11), .b(gate36inter6), .O(gate36inter12));
  nand2 gate742(.a(gate36inter12), .b(gate36inter1), .O(G347));
nand2 gate37( .a(G19), .b(G23), .O(G350) );
nand2 gate38( .a(G27), .b(G31), .O(G353) );
nand2 gate39( .a(G20), .b(G24), .O(G356) );
nand2 gate40( .a(G28), .b(G32), .O(G359) );
nand2 gate41( .a(G1), .b(G266), .O(G362) );

  xor2  gate841(.a(G266), .b(G2), .O(gate42inter0));
  nand2 gate842(.a(gate42inter0), .b(s_42), .O(gate42inter1));
  and2  gate843(.a(G266), .b(G2), .O(gate42inter2));
  inv1  gate844(.a(s_42), .O(gate42inter3));
  inv1  gate845(.a(s_43), .O(gate42inter4));
  nand2 gate846(.a(gate42inter4), .b(gate42inter3), .O(gate42inter5));
  nor2  gate847(.a(gate42inter5), .b(gate42inter2), .O(gate42inter6));
  inv1  gate848(.a(G2), .O(gate42inter7));
  inv1  gate849(.a(G266), .O(gate42inter8));
  nand2 gate850(.a(gate42inter8), .b(gate42inter7), .O(gate42inter9));
  nand2 gate851(.a(s_43), .b(gate42inter3), .O(gate42inter10));
  nor2  gate852(.a(gate42inter10), .b(gate42inter9), .O(gate42inter11));
  nor2  gate853(.a(gate42inter11), .b(gate42inter6), .O(gate42inter12));
  nand2 gate854(.a(gate42inter12), .b(gate42inter1), .O(G363));
nand2 gate43( .a(G3), .b(G269), .O(G364) );
nand2 gate44( .a(G4), .b(G269), .O(G365) );
nand2 gate45( .a(G5), .b(G272), .O(G366) );
nand2 gate46( .a(G6), .b(G272), .O(G367) );
nand2 gate47( .a(G7), .b(G275), .O(G368) );
nand2 gate48( .a(G8), .b(G275), .O(G369) );
nand2 gate49( .a(G9), .b(G278), .O(G370) );

  xor2  gate687(.a(G278), .b(G10), .O(gate50inter0));
  nand2 gate688(.a(gate50inter0), .b(s_20), .O(gate50inter1));
  and2  gate689(.a(G278), .b(G10), .O(gate50inter2));
  inv1  gate690(.a(s_20), .O(gate50inter3));
  inv1  gate691(.a(s_21), .O(gate50inter4));
  nand2 gate692(.a(gate50inter4), .b(gate50inter3), .O(gate50inter5));
  nor2  gate693(.a(gate50inter5), .b(gate50inter2), .O(gate50inter6));
  inv1  gate694(.a(G10), .O(gate50inter7));
  inv1  gate695(.a(G278), .O(gate50inter8));
  nand2 gate696(.a(gate50inter8), .b(gate50inter7), .O(gate50inter9));
  nand2 gate697(.a(s_21), .b(gate50inter3), .O(gate50inter10));
  nor2  gate698(.a(gate50inter10), .b(gate50inter9), .O(gate50inter11));
  nor2  gate699(.a(gate50inter11), .b(gate50inter6), .O(gate50inter12));
  nand2 gate700(.a(gate50inter12), .b(gate50inter1), .O(G371));
nand2 gate51( .a(G11), .b(G281), .O(G372) );
nand2 gate52( .a(G12), .b(G281), .O(G373) );
nand2 gate53( .a(G13), .b(G284), .O(G374) );

  xor2  gate1051(.a(G284), .b(G14), .O(gate54inter0));
  nand2 gate1052(.a(gate54inter0), .b(s_72), .O(gate54inter1));
  and2  gate1053(.a(G284), .b(G14), .O(gate54inter2));
  inv1  gate1054(.a(s_72), .O(gate54inter3));
  inv1  gate1055(.a(s_73), .O(gate54inter4));
  nand2 gate1056(.a(gate54inter4), .b(gate54inter3), .O(gate54inter5));
  nor2  gate1057(.a(gate54inter5), .b(gate54inter2), .O(gate54inter6));
  inv1  gate1058(.a(G14), .O(gate54inter7));
  inv1  gate1059(.a(G284), .O(gate54inter8));
  nand2 gate1060(.a(gate54inter8), .b(gate54inter7), .O(gate54inter9));
  nand2 gate1061(.a(s_73), .b(gate54inter3), .O(gate54inter10));
  nor2  gate1062(.a(gate54inter10), .b(gate54inter9), .O(gate54inter11));
  nor2  gate1063(.a(gate54inter11), .b(gate54inter6), .O(gate54inter12));
  nand2 gate1064(.a(gate54inter12), .b(gate54inter1), .O(G375));
nand2 gate55( .a(G15), .b(G287), .O(G376) );
nand2 gate56( .a(G16), .b(G287), .O(G377) );
nand2 gate57( .a(G17), .b(G290), .O(G378) );

  xor2  gate1079(.a(G290), .b(G18), .O(gate58inter0));
  nand2 gate1080(.a(gate58inter0), .b(s_76), .O(gate58inter1));
  and2  gate1081(.a(G290), .b(G18), .O(gate58inter2));
  inv1  gate1082(.a(s_76), .O(gate58inter3));
  inv1  gate1083(.a(s_77), .O(gate58inter4));
  nand2 gate1084(.a(gate58inter4), .b(gate58inter3), .O(gate58inter5));
  nor2  gate1085(.a(gate58inter5), .b(gate58inter2), .O(gate58inter6));
  inv1  gate1086(.a(G18), .O(gate58inter7));
  inv1  gate1087(.a(G290), .O(gate58inter8));
  nand2 gate1088(.a(gate58inter8), .b(gate58inter7), .O(gate58inter9));
  nand2 gate1089(.a(s_77), .b(gate58inter3), .O(gate58inter10));
  nor2  gate1090(.a(gate58inter10), .b(gate58inter9), .O(gate58inter11));
  nor2  gate1091(.a(gate58inter11), .b(gate58inter6), .O(gate58inter12));
  nand2 gate1092(.a(gate58inter12), .b(gate58inter1), .O(G379));
nand2 gate59( .a(G19), .b(G293), .O(G380) );
nand2 gate60( .a(G20), .b(G293), .O(G381) );
nand2 gate61( .a(G21), .b(G296), .O(G382) );
nand2 gate62( .a(G22), .b(G296), .O(G383) );

  xor2  gate547(.a(G299), .b(G23), .O(gate63inter0));
  nand2 gate548(.a(gate63inter0), .b(s_0), .O(gate63inter1));
  and2  gate549(.a(G299), .b(G23), .O(gate63inter2));
  inv1  gate550(.a(s_0), .O(gate63inter3));
  inv1  gate551(.a(s_1), .O(gate63inter4));
  nand2 gate552(.a(gate63inter4), .b(gate63inter3), .O(gate63inter5));
  nor2  gate553(.a(gate63inter5), .b(gate63inter2), .O(gate63inter6));
  inv1  gate554(.a(G23), .O(gate63inter7));
  inv1  gate555(.a(G299), .O(gate63inter8));
  nand2 gate556(.a(gate63inter8), .b(gate63inter7), .O(gate63inter9));
  nand2 gate557(.a(s_1), .b(gate63inter3), .O(gate63inter10));
  nor2  gate558(.a(gate63inter10), .b(gate63inter9), .O(gate63inter11));
  nor2  gate559(.a(gate63inter11), .b(gate63inter6), .O(gate63inter12));
  nand2 gate560(.a(gate63inter12), .b(gate63inter1), .O(G384));

  xor2  gate1037(.a(G299), .b(G24), .O(gate64inter0));
  nand2 gate1038(.a(gate64inter0), .b(s_70), .O(gate64inter1));
  and2  gate1039(.a(G299), .b(G24), .O(gate64inter2));
  inv1  gate1040(.a(s_70), .O(gate64inter3));
  inv1  gate1041(.a(s_71), .O(gate64inter4));
  nand2 gate1042(.a(gate64inter4), .b(gate64inter3), .O(gate64inter5));
  nor2  gate1043(.a(gate64inter5), .b(gate64inter2), .O(gate64inter6));
  inv1  gate1044(.a(G24), .O(gate64inter7));
  inv1  gate1045(.a(G299), .O(gate64inter8));
  nand2 gate1046(.a(gate64inter8), .b(gate64inter7), .O(gate64inter9));
  nand2 gate1047(.a(s_71), .b(gate64inter3), .O(gate64inter10));
  nor2  gate1048(.a(gate64inter10), .b(gate64inter9), .O(gate64inter11));
  nor2  gate1049(.a(gate64inter11), .b(gate64inter6), .O(gate64inter12));
  nand2 gate1050(.a(gate64inter12), .b(gate64inter1), .O(G385));
nand2 gate65( .a(G25), .b(G302), .O(G386) );
nand2 gate66( .a(G26), .b(G302), .O(G387) );
nand2 gate67( .a(G27), .b(G305), .O(G388) );
nand2 gate68( .a(G28), .b(G305), .O(G389) );
nand2 gate69( .a(G29), .b(G308), .O(G390) );
nand2 gate70( .a(G30), .b(G308), .O(G391) );
nand2 gate71( .a(G31), .b(G311), .O(G392) );
nand2 gate72( .a(G32), .b(G311), .O(G393) );
nand2 gate73( .a(G1), .b(G314), .O(G394) );
nand2 gate74( .a(G5), .b(G314), .O(G395) );
nand2 gate75( .a(G9), .b(G317), .O(G396) );
nand2 gate76( .a(G13), .b(G317), .O(G397) );
nand2 gate77( .a(G2), .b(G320), .O(G398) );

  xor2  gate967(.a(G320), .b(G6), .O(gate78inter0));
  nand2 gate968(.a(gate78inter0), .b(s_60), .O(gate78inter1));
  and2  gate969(.a(G320), .b(G6), .O(gate78inter2));
  inv1  gate970(.a(s_60), .O(gate78inter3));
  inv1  gate971(.a(s_61), .O(gate78inter4));
  nand2 gate972(.a(gate78inter4), .b(gate78inter3), .O(gate78inter5));
  nor2  gate973(.a(gate78inter5), .b(gate78inter2), .O(gate78inter6));
  inv1  gate974(.a(G6), .O(gate78inter7));
  inv1  gate975(.a(G320), .O(gate78inter8));
  nand2 gate976(.a(gate78inter8), .b(gate78inter7), .O(gate78inter9));
  nand2 gate977(.a(s_61), .b(gate78inter3), .O(gate78inter10));
  nor2  gate978(.a(gate78inter10), .b(gate78inter9), .O(gate78inter11));
  nor2  gate979(.a(gate78inter11), .b(gate78inter6), .O(gate78inter12));
  nand2 gate980(.a(gate78inter12), .b(gate78inter1), .O(G399));
nand2 gate79( .a(G10), .b(G323), .O(G400) );
nand2 gate80( .a(G14), .b(G323), .O(G401) );

  xor2  gate575(.a(G326), .b(G3), .O(gate81inter0));
  nand2 gate576(.a(gate81inter0), .b(s_4), .O(gate81inter1));
  and2  gate577(.a(G326), .b(G3), .O(gate81inter2));
  inv1  gate578(.a(s_4), .O(gate81inter3));
  inv1  gate579(.a(s_5), .O(gate81inter4));
  nand2 gate580(.a(gate81inter4), .b(gate81inter3), .O(gate81inter5));
  nor2  gate581(.a(gate81inter5), .b(gate81inter2), .O(gate81inter6));
  inv1  gate582(.a(G3), .O(gate81inter7));
  inv1  gate583(.a(G326), .O(gate81inter8));
  nand2 gate584(.a(gate81inter8), .b(gate81inter7), .O(gate81inter9));
  nand2 gate585(.a(s_5), .b(gate81inter3), .O(gate81inter10));
  nor2  gate586(.a(gate81inter10), .b(gate81inter9), .O(gate81inter11));
  nor2  gate587(.a(gate81inter11), .b(gate81inter6), .O(gate81inter12));
  nand2 gate588(.a(gate81inter12), .b(gate81inter1), .O(G402));
nand2 gate82( .a(G7), .b(G326), .O(G403) );
nand2 gate83( .a(G11), .b(G329), .O(G404) );
nand2 gate84( .a(G15), .b(G329), .O(G405) );
nand2 gate85( .a(G4), .b(G332), .O(G406) );
nand2 gate86( .a(G8), .b(G332), .O(G407) );
nand2 gate87( .a(G12), .b(G335), .O(G408) );
nand2 gate88( .a(G16), .b(G335), .O(G409) );
nand2 gate89( .a(G17), .b(G338), .O(G410) );
nand2 gate90( .a(G21), .b(G338), .O(G411) );

  xor2  gate799(.a(G341), .b(G25), .O(gate91inter0));
  nand2 gate800(.a(gate91inter0), .b(s_36), .O(gate91inter1));
  and2  gate801(.a(G341), .b(G25), .O(gate91inter2));
  inv1  gate802(.a(s_36), .O(gate91inter3));
  inv1  gate803(.a(s_37), .O(gate91inter4));
  nand2 gate804(.a(gate91inter4), .b(gate91inter3), .O(gate91inter5));
  nor2  gate805(.a(gate91inter5), .b(gate91inter2), .O(gate91inter6));
  inv1  gate806(.a(G25), .O(gate91inter7));
  inv1  gate807(.a(G341), .O(gate91inter8));
  nand2 gate808(.a(gate91inter8), .b(gate91inter7), .O(gate91inter9));
  nand2 gate809(.a(s_37), .b(gate91inter3), .O(gate91inter10));
  nor2  gate810(.a(gate91inter10), .b(gate91inter9), .O(gate91inter11));
  nor2  gate811(.a(gate91inter11), .b(gate91inter6), .O(gate91inter12));
  nand2 gate812(.a(gate91inter12), .b(gate91inter1), .O(G412));
nand2 gate92( .a(G29), .b(G341), .O(G413) );
nand2 gate93( .a(G18), .b(G344), .O(G414) );
nand2 gate94( .a(G22), .b(G344), .O(G415) );
nand2 gate95( .a(G26), .b(G347), .O(G416) );
nand2 gate96( .a(G30), .b(G347), .O(G417) );
nand2 gate97( .a(G19), .b(G350), .O(G418) );
nand2 gate98( .a(G23), .b(G350), .O(G419) );
nand2 gate99( .a(G27), .b(G353), .O(G420) );

  xor2  gate953(.a(G353), .b(G31), .O(gate100inter0));
  nand2 gate954(.a(gate100inter0), .b(s_58), .O(gate100inter1));
  and2  gate955(.a(G353), .b(G31), .O(gate100inter2));
  inv1  gate956(.a(s_58), .O(gate100inter3));
  inv1  gate957(.a(s_59), .O(gate100inter4));
  nand2 gate958(.a(gate100inter4), .b(gate100inter3), .O(gate100inter5));
  nor2  gate959(.a(gate100inter5), .b(gate100inter2), .O(gate100inter6));
  inv1  gate960(.a(G31), .O(gate100inter7));
  inv1  gate961(.a(G353), .O(gate100inter8));
  nand2 gate962(.a(gate100inter8), .b(gate100inter7), .O(gate100inter9));
  nand2 gate963(.a(s_59), .b(gate100inter3), .O(gate100inter10));
  nor2  gate964(.a(gate100inter10), .b(gate100inter9), .O(gate100inter11));
  nor2  gate965(.a(gate100inter11), .b(gate100inter6), .O(gate100inter12));
  nand2 gate966(.a(gate100inter12), .b(gate100inter1), .O(G421));
nand2 gate101( .a(G20), .b(G356), .O(G422) );
nand2 gate102( .a(G24), .b(G356), .O(G423) );
nand2 gate103( .a(G28), .b(G359), .O(G424) );
nand2 gate104( .a(G32), .b(G359), .O(G425) );
nand2 gate105( .a(G362), .b(G363), .O(G426) );
nand2 gate106( .a(G364), .b(G365), .O(G429) );
nand2 gate107( .a(G366), .b(G367), .O(G432) );
nand2 gate108( .a(G368), .b(G369), .O(G435) );
nand2 gate109( .a(G370), .b(G371), .O(G438) );

  xor2  gate645(.a(G373), .b(G372), .O(gate110inter0));
  nand2 gate646(.a(gate110inter0), .b(s_14), .O(gate110inter1));
  and2  gate647(.a(G373), .b(G372), .O(gate110inter2));
  inv1  gate648(.a(s_14), .O(gate110inter3));
  inv1  gate649(.a(s_15), .O(gate110inter4));
  nand2 gate650(.a(gate110inter4), .b(gate110inter3), .O(gate110inter5));
  nor2  gate651(.a(gate110inter5), .b(gate110inter2), .O(gate110inter6));
  inv1  gate652(.a(G372), .O(gate110inter7));
  inv1  gate653(.a(G373), .O(gate110inter8));
  nand2 gate654(.a(gate110inter8), .b(gate110inter7), .O(gate110inter9));
  nand2 gate655(.a(s_15), .b(gate110inter3), .O(gate110inter10));
  nor2  gate656(.a(gate110inter10), .b(gate110inter9), .O(gate110inter11));
  nor2  gate657(.a(gate110inter11), .b(gate110inter6), .O(gate110inter12));
  nand2 gate658(.a(gate110inter12), .b(gate110inter1), .O(G441));

  xor2  gate1093(.a(G375), .b(G374), .O(gate111inter0));
  nand2 gate1094(.a(gate111inter0), .b(s_78), .O(gate111inter1));
  and2  gate1095(.a(G375), .b(G374), .O(gate111inter2));
  inv1  gate1096(.a(s_78), .O(gate111inter3));
  inv1  gate1097(.a(s_79), .O(gate111inter4));
  nand2 gate1098(.a(gate111inter4), .b(gate111inter3), .O(gate111inter5));
  nor2  gate1099(.a(gate111inter5), .b(gate111inter2), .O(gate111inter6));
  inv1  gate1100(.a(G374), .O(gate111inter7));
  inv1  gate1101(.a(G375), .O(gate111inter8));
  nand2 gate1102(.a(gate111inter8), .b(gate111inter7), .O(gate111inter9));
  nand2 gate1103(.a(s_79), .b(gate111inter3), .O(gate111inter10));
  nor2  gate1104(.a(gate111inter10), .b(gate111inter9), .O(gate111inter11));
  nor2  gate1105(.a(gate111inter11), .b(gate111inter6), .O(gate111inter12));
  nand2 gate1106(.a(gate111inter12), .b(gate111inter1), .O(G444));

  xor2  gate603(.a(G377), .b(G376), .O(gate112inter0));
  nand2 gate604(.a(gate112inter0), .b(s_8), .O(gate112inter1));
  and2  gate605(.a(G377), .b(G376), .O(gate112inter2));
  inv1  gate606(.a(s_8), .O(gate112inter3));
  inv1  gate607(.a(s_9), .O(gate112inter4));
  nand2 gate608(.a(gate112inter4), .b(gate112inter3), .O(gate112inter5));
  nor2  gate609(.a(gate112inter5), .b(gate112inter2), .O(gate112inter6));
  inv1  gate610(.a(G376), .O(gate112inter7));
  inv1  gate611(.a(G377), .O(gate112inter8));
  nand2 gate612(.a(gate112inter8), .b(gate112inter7), .O(gate112inter9));
  nand2 gate613(.a(s_9), .b(gate112inter3), .O(gate112inter10));
  nor2  gate614(.a(gate112inter10), .b(gate112inter9), .O(gate112inter11));
  nor2  gate615(.a(gate112inter11), .b(gate112inter6), .O(gate112inter12));
  nand2 gate616(.a(gate112inter12), .b(gate112inter1), .O(G447));
nand2 gate113( .a(G378), .b(G379), .O(G450) );
nand2 gate114( .a(G380), .b(G381), .O(G453) );
nand2 gate115( .a(G382), .b(G383), .O(G456) );
nand2 gate116( .a(G384), .b(G385), .O(G459) );
nand2 gate117( .a(G386), .b(G387), .O(G462) );
nand2 gate118( .a(G388), .b(G389), .O(G465) );

  xor2  gate757(.a(G391), .b(G390), .O(gate119inter0));
  nand2 gate758(.a(gate119inter0), .b(s_30), .O(gate119inter1));
  and2  gate759(.a(G391), .b(G390), .O(gate119inter2));
  inv1  gate760(.a(s_30), .O(gate119inter3));
  inv1  gate761(.a(s_31), .O(gate119inter4));
  nand2 gate762(.a(gate119inter4), .b(gate119inter3), .O(gate119inter5));
  nor2  gate763(.a(gate119inter5), .b(gate119inter2), .O(gate119inter6));
  inv1  gate764(.a(G390), .O(gate119inter7));
  inv1  gate765(.a(G391), .O(gate119inter8));
  nand2 gate766(.a(gate119inter8), .b(gate119inter7), .O(gate119inter9));
  nand2 gate767(.a(s_31), .b(gate119inter3), .O(gate119inter10));
  nor2  gate768(.a(gate119inter10), .b(gate119inter9), .O(gate119inter11));
  nor2  gate769(.a(gate119inter11), .b(gate119inter6), .O(gate119inter12));
  nand2 gate770(.a(gate119inter12), .b(gate119inter1), .O(G468));
nand2 gate120( .a(G392), .b(G393), .O(G471) );

  xor2  gate785(.a(G395), .b(G394), .O(gate121inter0));
  nand2 gate786(.a(gate121inter0), .b(s_34), .O(gate121inter1));
  and2  gate787(.a(G395), .b(G394), .O(gate121inter2));
  inv1  gate788(.a(s_34), .O(gate121inter3));
  inv1  gate789(.a(s_35), .O(gate121inter4));
  nand2 gate790(.a(gate121inter4), .b(gate121inter3), .O(gate121inter5));
  nor2  gate791(.a(gate121inter5), .b(gate121inter2), .O(gate121inter6));
  inv1  gate792(.a(G394), .O(gate121inter7));
  inv1  gate793(.a(G395), .O(gate121inter8));
  nand2 gate794(.a(gate121inter8), .b(gate121inter7), .O(gate121inter9));
  nand2 gate795(.a(s_35), .b(gate121inter3), .O(gate121inter10));
  nor2  gate796(.a(gate121inter10), .b(gate121inter9), .O(gate121inter11));
  nor2  gate797(.a(gate121inter11), .b(gate121inter6), .O(gate121inter12));
  nand2 gate798(.a(gate121inter12), .b(gate121inter1), .O(G474));
nand2 gate122( .a(G396), .b(G397), .O(G477) );
nand2 gate123( .a(G398), .b(G399), .O(G480) );
nand2 gate124( .a(G400), .b(G401), .O(G483) );
nand2 gate125( .a(G402), .b(G403), .O(G486) );
nand2 gate126( .a(G404), .b(G405), .O(G489) );
nand2 gate127( .a(G406), .b(G407), .O(G492) );
nand2 gate128( .a(G408), .b(G409), .O(G495) );

  xor2  gate659(.a(G411), .b(G410), .O(gate129inter0));
  nand2 gate660(.a(gate129inter0), .b(s_16), .O(gate129inter1));
  and2  gate661(.a(G411), .b(G410), .O(gate129inter2));
  inv1  gate662(.a(s_16), .O(gate129inter3));
  inv1  gate663(.a(s_17), .O(gate129inter4));
  nand2 gate664(.a(gate129inter4), .b(gate129inter3), .O(gate129inter5));
  nor2  gate665(.a(gate129inter5), .b(gate129inter2), .O(gate129inter6));
  inv1  gate666(.a(G410), .O(gate129inter7));
  inv1  gate667(.a(G411), .O(gate129inter8));
  nand2 gate668(.a(gate129inter8), .b(gate129inter7), .O(gate129inter9));
  nand2 gate669(.a(s_17), .b(gate129inter3), .O(gate129inter10));
  nor2  gate670(.a(gate129inter10), .b(gate129inter9), .O(gate129inter11));
  nor2  gate671(.a(gate129inter11), .b(gate129inter6), .O(gate129inter12));
  nand2 gate672(.a(gate129inter12), .b(gate129inter1), .O(G498));
nand2 gate130( .a(G412), .b(G413), .O(G501) );
nand2 gate131( .a(G414), .b(G415), .O(G504) );
nand2 gate132( .a(G416), .b(G417), .O(G507) );
nand2 gate133( .a(G418), .b(G419), .O(G510) );

  xor2  gate673(.a(G421), .b(G420), .O(gate134inter0));
  nand2 gate674(.a(gate134inter0), .b(s_18), .O(gate134inter1));
  and2  gate675(.a(G421), .b(G420), .O(gate134inter2));
  inv1  gate676(.a(s_18), .O(gate134inter3));
  inv1  gate677(.a(s_19), .O(gate134inter4));
  nand2 gate678(.a(gate134inter4), .b(gate134inter3), .O(gate134inter5));
  nor2  gate679(.a(gate134inter5), .b(gate134inter2), .O(gate134inter6));
  inv1  gate680(.a(G420), .O(gate134inter7));
  inv1  gate681(.a(G421), .O(gate134inter8));
  nand2 gate682(.a(gate134inter8), .b(gate134inter7), .O(gate134inter9));
  nand2 gate683(.a(s_19), .b(gate134inter3), .O(gate134inter10));
  nor2  gate684(.a(gate134inter10), .b(gate134inter9), .O(gate134inter11));
  nor2  gate685(.a(gate134inter11), .b(gate134inter6), .O(gate134inter12));
  nand2 gate686(.a(gate134inter12), .b(gate134inter1), .O(G513));
nand2 gate135( .a(G422), .b(G423), .O(G516) );
nand2 gate136( .a(G424), .b(G425), .O(G519) );
nand2 gate137( .a(G426), .b(G429), .O(G522) );
nand2 gate138( .a(G432), .b(G435), .O(G525) );
nand2 gate139( .a(G438), .b(G441), .O(G528) );
nand2 gate140( .a(G444), .b(G447), .O(G531) );
nand2 gate141( .a(G450), .b(G453), .O(G534) );
nand2 gate142( .a(G456), .b(G459), .O(G537) );
nand2 gate143( .a(G462), .b(G465), .O(G540) );
nand2 gate144( .a(G468), .b(G471), .O(G543) );
nand2 gate145( .a(G474), .b(G477), .O(G546) );
nand2 gate146( .a(G480), .b(G483), .O(G549) );
nand2 gate147( .a(G486), .b(G489), .O(G552) );
nand2 gate148( .a(G492), .b(G495), .O(G555) );
nand2 gate149( .a(G498), .b(G501), .O(G558) );

  xor2  gate827(.a(G507), .b(G504), .O(gate150inter0));
  nand2 gate828(.a(gate150inter0), .b(s_40), .O(gate150inter1));
  and2  gate829(.a(G507), .b(G504), .O(gate150inter2));
  inv1  gate830(.a(s_40), .O(gate150inter3));
  inv1  gate831(.a(s_41), .O(gate150inter4));
  nand2 gate832(.a(gate150inter4), .b(gate150inter3), .O(gate150inter5));
  nor2  gate833(.a(gate150inter5), .b(gate150inter2), .O(gate150inter6));
  inv1  gate834(.a(G504), .O(gate150inter7));
  inv1  gate835(.a(G507), .O(gate150inter8));
  nand2 gate836(.a(gate150inter8), .b(gate150inter7), .O(gate150inter9));
  nand2 gate837(.a(s_41), .b(gate150inter3), .O(gate150inter10));
  nor2  gate838(.a(gate150inter10), .b(gate150inter9), .O(gate150inter11));
  nor2  gate839(.a(gate150inter11), .b(gate150inter6), .O(gate150inter12));
  nand2 gate840(.a(gate150inter12), .b(gate150inter1), .O(G561));
nand2 gate151( .a(G510), .b(G513), .O(G564) );
nand2 gate152( .a(G516), .b(G519), .O(G567) );
nand2 gate153( .a(G426), .b(G522), .O(G570) );
nand2 gate154( .a(G429), .b(G522), .O(G571) );
nand2 gate155( .a(G432), .b(G525), .O(G572) );
nand2 gate156( .a(G435), .b(G525), .O(G573) );
nand2 gate157( .a(G438), .b(G528), .O(G574) );
nand2 gate158( .a(G441), .b(G528), .O(G575) );
nand2 gate159( .a(G444), .b(G531), .O(G576) );
nand2 gate160( .a(G447), .b(G531), .O(G577) );
nand2 gate161( .a(G450), .b(G534), .O(G578) );
nand2 gate162( .a(G453), .b(G534), .O(G579) );
nand2 gate163( .a(G456), .b(G537), .O(G580) );
nand2 gate164( .a(G459), .b(G537), .O(G581) );
nand2 gate165( .a(G462), .b(G540), .O(G582) );
nand2 gate166( .a(G465), .b(G540), .O(G583) );
nand2 gate167( .a(G468), .b(G543), .O(G584) );
nand2 gate168( .a(G471), .b(G543), .O(G585) );
nand2 gate169( .a(G474), .b(G546), .O(G586) );

  xor2  gate925(.a(G546), .b(G477), .O(gate170inter0));
  nand2 gate926(.a(gate170inter0), .b(s_54), .O(gate170inter1));
  and2  gate927(.a(G546), .b(G477), .O(gate170inter2));
  inv1  gate928(.a(s_54), .O(gate170inter3));
  inv1  gate929(.a(s_55), .O(gate170inter4));
  nand2 gate930(.a(gate170inter4), .b(gate170inter3), .O(gate170inter5));
  nor2  gate931(.a(gate170inter5), .b(gate170inter2), .O(gate170inter6));
  inv1  gate932(.a(G477), .O(gate170inter7));
  inv1  gate933(.a(G546), .O(gate170inter8));
  nand2 gate934(.a(gate170inter8), .b(gate170inter7), .O(gate170inter9));
  nand2 gate935(.a(s_55), .b(gate170inter3), .O(gate170inter10));
  nor2  gate936(.a(gate170inter10), .b(gate170inter9), .O(gate170inter11));
  nor2  gate937(.a(gate170inter11), .b(gate170inter6), .O(gate170inter12));
  nand2 gate938(.a(gate170inter12), .b(gate170inter1), .O(G587));
nand2 gate171( .a(G480), .b(G549), .O(G588) );
nand2 gate172( .a(G483), .b(G549), .O(G589) );
nand2 gate173( .a(G486), .b(G552), .O(G590) );
nand2 gate174( .a(G489), .b(G552), .O(G591) );
nand2 gate175( .a(G492), .b(G555), .O(G592) );
nand2 gate176( .a(G495), .b(G555), .O(G593) );
nand2 gate177( .a(G498), .b(G558), .O(G594) );
nand2 gate178( .a(G501), .b(G558), .O(G595) );
nand2 gate179( .a(G504), .b(G561), .O(G596) );
nand2 gate180( .a(G507), .b(G561), .O(G597) );
nand2 gate181( .a(G510), .b(G564), .O(G598) );
nand2 gate182( .a(G513), .b(G564), .O(G599) );
nand2 gate183( .a(G516), .b(G567), .O(G600) );
nand2 gate184( .a(G519), .b(G567), .O(G601) );
nand2 gate185( .a(G570), .b(G571), .O(G602) );
nand2 gate186( .a(G572), .b(G573), .O(G607) );
nand2 gate187( .a(G574), .b(G575), .O(G612) );

  xor2  gate589(.a(G577), .b(G576), .O(gate188inter0));
  nand2 gate590(.a(gate188inter0), .b(s_6), .O(gate188inter1));
  and2  gate591(.a(G577), .b(G576), .O(gate188inter2));
  inv1  gate592(.a(s_6), .O(gate188inter3));
  inv1  gate593(.a(s_7), .O(gate188inter4));
  nand2 gate594(.a(gate188inter4), .b(gate188inter3), .O(gate188inter5));
  nor2  gate595(.a(gate188inter5), .b(gate188inter2), .O(gate188inter6));
  inv1  gate596(.a(G576), .O(gate188inter7));
  inv1  gate597(.a(G577), .O(gate188inter8));
  nand2 gate598(.a(gate188inter8), .b(gate188inter7), .O(gate188inter9));
  nand2 gate599(.a(s_7), .b(gate188inter3), .O(gate188inter10));
  nor2  gate600(.a(gate188inter10), .b(gate188inter9), .O(gate188inter11));
  nor2  gate601(.a(gate188inter11), .b(gate188inter6), .O(gate188inter12));
  nand2 gate602(.a(gate188inter12), .b(gate188inter1), .O(G617));
nand2 gate189( .a(G578), .b(G579), .O(G622) );
nand2 gate190( .a(G580), .b(G581), .O(G627) );
nand2 gate191( .a(G582), .b(G583), .O(G632) );
nand2 gate192( .a(G584), .b(G585), .O(G637) );
nand2 gate193( .a(G586), .b(G587), .O(G642) );
nand2 gate194( .a(G588), .b(G589), .O(G645) );
nand2 gate195( .a(G590), .b(G591), .O(G648) );
nand2 gate196( .a(G592), .b(G593), .O(G651) );
nand2 gate197( .a(G594), .b(G595), .O(G654) );

  xor2  gate883(.a(G597), .b(G596), .O(gate198inter0));
  nand2 gate884(.a(gate198inter0), .b(s_48), .O(gate198inter1));
  and2  gate885(.a(G597), .b(G596), .O(gate198inter2));
  inv1  gate886(.a(s_48), .O(gate198inter3));
  inv1  gate887(.a(s_49), .O(gate198inter4));
  nand2 gate888(.a(gate198inter4), .b(gate198inter3), .O(gate198inter5));
  nor2  gate889(.a(gate198inter5), .b(gate198inter2), .O(gate198inter6));
  inv1  gate890(.a(G596), .O(gate198inter7));
  inv1  gate891(.a(G597), .O(gate198inter8));
  nand2 gate892(.a(gate198inter8), .b(gate198inter7), .O(gate198inter9));
  nand2 gate893(.a(s_49), .b(gate198inter3), .O(gate198inter10));
  nor2  gate894(.a(gate198inter10), .b(gate198inter9), .O(gate198inter11));
  nor2  gate895(.a(gate198inter11), .b(gate198inter6), .O(gate198inter12));
  nand2 gate896(.a(gate198inter12), .b(gate198inter1), .O(G657));
nand2 gate199( .a(G598), .b(G599), .O(G660) );
nand2 gate200( .a(G600), .b(G601), .O(G663) );
nand2 gate201( .a(G602), .b(G607), .O(G666) );
nand2 gate202( .a(G612), .b(G617), .O(G669) );
nand2 gate203( .a(G602), .b(G612), .O(G672) );
nand2 gate204( .a(G607), .b(G617), .O(G675) );
nand2 gate205( .a(G622), .b(G627), .O(G678) );
nand2 gate206( .a(G632), .b(G637), .O(G681) );
nand2 gate207( .a(G622), .b(G632), .O(G684) );
nand2 gate208( .a(G627), .b(G637), .O(G687) );
nand2 gate209( .a(G602), .b(G666), .O(G690) );
nand2 gate210( .a(G607), .b(G666), .O(G691) );
nand2 gate211( .a(G612), .b(G669), .O(G692) );
nand2 gate212( .a(G617), .b(G669), .O(G693) );
nand2 gate213( .a(G602), .b(G672), .O(G694) );
nand2 gate214( .a(G612), .b(G672), .O(G695) );
nand2 gate215( .a(G607), .b(G675), .O(G696) );
nand2 gate216( .a(G617), .b(G675), .O(G697) );
nand2 gate217( .a(G622), .b(G678), .O(G698) );
nand2 gate218( .a(G627), .b(G678), .O(G699) );

  xor2  gate771(.a(G681), .b(G632), .O(gate219inter0));
  nand2 gate772(.a(gate219inter0), .b(s_32), .O(gate219inter1));
  and2  gate773(.a(G681), .b(G632), .O(gate219inter2));
  inv1  gate774(.a(s_32), .O(gate219inter3));
  inv1  gate775(.a(s_33), .O(gate219inter4));
  nand2 gate776(.a(gate219inter4), .b(gate219inter3), .O(gate219inter5));
  nor2  gate777(.a(gate219inter5), .b(gate219inter2), .O(gate219inter6));
  inv1  gate778(.a(G632), .O(gate219inter7));
  inv1  gate779(.a(G681), .O(gate219inter8));
  nand2 gate780(.a(gate219inter8), .b(gate219inter7), .O(gate219inter9));
  nand2 gate781(.a(s_33), .b(gate219inter3), .O(gate219inter10));
  nor2  gate782(.a(gate219inter10), .b(gate219inter9), .O(gate219inter11));
  nor2  gate783(.a(gate219inter11), .b(gate219inter6), .O(gate219inter12));
  nand2 gate784(.a(gate219inter12), .b(gate219inter1), .O(G700));
nand2 gate220( .a(G637), .b(G681), .O(G701) );
nand2 gate221( .a(G622), .b(G684), .O(G702) );
nand2 gate222( .a(G632), .b(G684), .O(G703) );
nand2 gate223( .a(G627), .b(G687), .O(G704) );
nand2 gate224( .a(G637), .b(G687), .O(G705) );

  xor2  gate813(.a(G691), .b(G690), .O(gate225inter0));
  nand2 gate814(.a(gate225inter0), .b(s_38), .O(gate225inter1));
  and2  gate815(.a(G691), .b(G690), .O(gate225inter2));
  inv1  gate816(.a(s_38), .O(gate225inter3));
  inv1  gate817(.a(s_39), .O(gate225inter4));
  nand2 gate818(.a(gate225inter4), .b(gate225inter3), .O(gate225inter5));
  nor2  gate819(.a(gate225inter5), .b(gate225inter2), .O(gate225inter6));
  inv1  gate820(.a(G690), .O(gate225inter7));
  inv1  gate821(.a(G691), .O(gate225inter8));
  nand2 gate822(.a(gate225inter8), .b(gate225inter7), .O(gate225inter9));
  nand2 gate823(.a(s_39), .b(gate225inter3), .O(gate225inter10));
  nor2  gate824(.a(gate225inter10), .b(gate225inter9), .O(gate225inter11));
  nor2  gate825(.a(gate225inter11), .b(gate225inter6), .O(gate225inter12));
  nand2 gate826(.a(gate225inter12), .b(gate225inter1), .O(G706));
nand2 gate226( .a(G692), .b(G693), .O(G709) );
nand2 gate227( .a(G694), .b(G695), .O(G712) );

  xor2  gate939(.a(G697), .b(G696), .O(gate228inter0));
  nand2 gate940(.a(gate228inter0), .b(s_56), .O(gate228inter1));
  and2  gate941(.a(G697), .b(G696), .O(gate228inter2));
  inv1  gate942(.a(s_56), .O(gate228inter3));
  inv1  gate943(.a(s_57), .O(gate228inter4));
  nand2 gate944(.a(gate228inter4), .b(gate228inter3), .O(gate228inter5));
  nor2  gate945(.a(gate228inter5), .b(gate228inter2), .O(gate228inter6));
  inv1  gate946(.a(G696), .O(gate228inter7));
  inv1  gate947(.a(G697), .O(gate228inter8));
  nand2 gate948(.a(gate228inter8), .b(gate228inter7), .O(gate228inter9));
  nand2 gate949(.a(s_57), .b(gate228inter3), .O(gate228inter10));
  nor2  gate950(.a(gate228inter10), .b(gate228inter9), .O(gate228inter11));
  nor2  gate951(.a(gate228inter11), .b(gate228inter6), .O(gate228inter12));
  nand2 gate952(.a(gate228inter12), .b(gate228inter1), .O(G715));
nand2 gate229( .a(G698), .b(G699), .O(G718) );
nand2 gate230( .a(G700), .b(G701), .O(G721) );
nand2 gate231( .a(G702), .b(G703), .O(G724) );
nand2 gate232( .a(G704), .b(G705), .O(G727) );
nand2 gate233( .a(G242), .b(G718), .O(G730) );
nand2 gate234( .a(G245), .b(G721), .O(G733) );
nand2 gate235( .a(G248), .b(G724), .O(G736) );
nand2 gate236( .a(G251), .b(G727), .O(G739) );

  xor2  gate631(.a(G706), .b(G254), .O(gate237inter0));
  nand2 gate632(.a(gate237inter0), .b(s_12), .O(gate237inter1));
  and2  gate633(.a(G706), .b(G254), .O(gate237inter2));
  inv1  gate634(.a(s_12), .O(gate237inter3));
  inv1  gate635(.a(s_13), .O(gate237inter4));
  nand2 gate636(.a(gate237inter4), .b(gate237inter3), .O(gate237inter5));
  nor2  gate637(.a(gate237inter5), .b(gate237inter2), .O(gate237inter6));
  inv1  gate638(.a(G254), .O(gate237inter7));
  inv1  gate639(.a(G706), .O(gate237inter8));
  nand2 gate640(.a(gate237inter8), .b(gate237inter7), .O(gate237inter9));
  nand2 gate641(.a(s_13), .b(gate237inter3), .O(gate237inter10));
  nor2  gate642(.a(gate237inter10), .b(gate237inter9), .O(gate237inter11));
  nor2  gate643(.a(gate237inter11), .b(gate237inter6), .O(gate237inter12));
  nand2 gate644(.a(gate237inter12), .b(gate237inter1), .O(G742));
nand2 gate238( .a(G257), .b(G709), .O(G745) );
nand2 gate239( .a(G260), .b(G712), .O(G748) );
nand2 gate240( .a(G263), .b(G715), .O(G751) );
nand2 gate241( .a(G242), .b(G730), .O(G754) );
nand2 gate242( .a(G718), .b(G730), .O(G755) );
nand2 gate243( .a(G245), .b(G733), .O(G756) );
nand2 gate244( .a(G721), .b(G733), .O(G757) );
nand2 gate245( .a(G248), .b(G736), .O(G758) );
nand2 gate246( .a(G724), .b(G736), .O(G759) );
nand2 gate247( .a(G251), .b(G739), .O(G760) );
nand2 gate248( .a(G727), .b(G739), .O(G761) );
nand2 gate249( .a(G254), .b(G742), .O(G762) );
nand2 gate250( .a(G706), .b(G742), .O(G763) );
nand2 gate251( .a(G257), .b(G745), .O(G764) );
nand2 gate252( .a(G709), .b(G745), .O(G765) );
nand2 gate253( .a(G260), .b(G748), .O(G766) );
nand2 gate254( .a(G712), .b(G748), .O(G767) );
nand2 gate255( .a(G263), .b(G751), .O(G768) );
nand2 gate256( .a(G715), .b(G751), .O(G769) );
nand2 gate257( .a(G754), .b(G755), .O(G770) );
nand2 gate258( .a(G756), .b(G757), .O(G773) );
nand2 gate259( .a(G758), .b(G759), .O(G776) );

  xor2  gate617(.a(G761), .b(G760), .O(gate260inter0));
  nand2 gate618(.a(gate260inter0), .b(s_10), .O(gate260inter1));
  and2  gate619(.a(G761), .b(G760), .O(gate260inter2));
  inv1  gate620(.a(s_10), .O(gate260inter3));
  inv1  gate621(.a(s_11), .O(gate260inter4));
  nand2 gate622(.a(gate260inter4), .b(gate260inter3), .O(gate260inter5));
  nor2  gate623(.a(gate260inter5), .b(gate260inter2), .O(gate260inter6));
  inv1  gate624(.a(G760), .O(gate260inter7));
  inv1  gate625(.a(G761), .O(gate260inter8));
  nand2 gate626(.a(gate260inter8), .b(gate260inter7), .O(gate260inter9));
  nand2 gate627(.a(s_11), .b(gate260inter3), .O(gate260inter10));
  nor2  gate628(.a(gate260inter10), .b(gate260inter9), .O(gate260inter11));
  nor2  gate629(.a(gate260inter11), .b(gate260inter6), .O(gate260inter12));
  nand2 gate630(.a(gate260inter12), .b(gate260inter1), .O(G779));
nand2 gate261( .a(G762), .b(G763), .O(G782) );
nand2 gate262( .a(G764), .b(G765), .O(G785) );
nand2 gate263( .a(G766), .b(G767), .O(G788) );
nand2 gate264( .a(G768), .b(G769), .O(G791) );

  xor2  gate715(.a(G770), .b(G642), .O(gate265inter0));
  nand2 gate716(.a(gate265inter0), .b(s_24), .O(gate265inter1));
  and2  gate717(.a(G770), .b(G642), .O(gate265inter2));
  inv1  gate718(.a(s_24), .O(gate265inter3));
  inv1  gate719(.a(s_25), .O(gate265inter4));
  nand2 gate720(.a(gate265inter4), .b(gate265inter3), .O(gate265inter5));
  nor2  gate721(.a(gate265inter5), .b(gate265inter2), .O(gate265inter6));
  inv1  gate722(.a(G642), .O(gate265inter7));
  inv1  gate723(.a(G770), .O(gate265inter8));
  nand2 gate724(.a(gate265inter8), .b(gate265inter7), .O(gate265inter9));
  nand2 gate725(.a(s_25), .b(gate265inter3), .O(gate265inter10));
  nor2  gate726(.a(gate265inter10), .b(gate265inter9), .O(gate265inter11));
  nor2  gate727(.a(gate265inter11), .b(gate265inter6), .O(gate265inter12));
  nand2 gate728(.a(gate265inter12), .b(gate265inter1), .O(G794));
nand2 gate266( .a(G645), .b(G773), .O(G797) );
nand2 gate267( .a(G648), .b(G776), .O(G800) );
nand2 gate268( .a(G651), .b(G779), .O(G803) );
nand2 gate269( .a(G654), .b(G782), .O(G806) );

  xor2  gate995(.a(G785), .b(G657), .O(gate270inter0));
  nand2 gate996(.a(gate270inter0), .b(s_64), .O(gate270inter1));
  and2  gate997(.a(G785), .b(G657), .O(gate270inter2));
  inv1  gate998(.a(s_64), .O(gate270inter3));
  inv1  gate999(.a(s_65), .O(gate270inter4));
  nand2 gate1000(.a(gate270inter4), .b(gate270inter3), .O(gate270inter5));
  nor2  gate1001(.a(gate270inter5), .b(gate270inter2), .O(gate270inter6));
  inv1  gate1002(.a(G657), .O(gate270inter7));
  inv1  gate1003(.a(G785), .O(gate270inter8));
  nand2 gate1004(.a(gate270inter8), .b(gate270inter7), .O(gate270inter9));
  nand2 gate1005(.a(s_65), .b(gate270inter3), .O(gate270inter10));
  nor2  gate1006(.a(gate270inter10), .b(gate270inter9), .O(gate270inter11));
  nor2  gate1007(.a(gate270inter11), .b(gate270inter6), .O(gate270inter12));
  nand2 gate1008(.a(gate270inter12), .b(gate270inter1), .O(G809));
nand2 gate271( .a(G660), .b(G788), .O(G812) );
nand2 gate272( .a(G663), .b(G791), .O(G815) );
nand2 gate273( .a(G642), .b(G794), .O(G818) );
nand2 gate274( .a(G770), .b(G794), .O(G819) );
nand2 gate275( .a(G645), .b(G797), .O(G820) );
nand2 gate276( .a(G773), .b(G797), .O(G821) );
nand2 gate277( .a(G648), .b(G800), .O(G822) );
nand2 gate278( .a(G776), .b(G800), .O(G823) );
nand2 gate279( .a(G651), .b(G803), .O(G824) );
nand2 gate280( .a(G779), .b(G803), .O(G825) );
nand2 gate281( .a(G654), .b(G806), .O(G826) );
nand2 gate282( .a(G782), .b(G806), .O(G827) );
nand2 gate283( .a(G657), .b(G809), .O(G828) );
nand2 gate284( .a(G785), .b(G809), .O(G829) );
nand2 gate285( .a(G660), .b(G812), .O(G830) );
nand2 gate286( .a(G788), .b(G812), .O(G831) );
nand2 gate287( .a(G663), .b(G815), .O(G832) );
nand2 gate288( .a(G791), .b(G815), .O(G833) );
nand2 gate289( .a(G818), .b(G819), .O(G834) );
nand2 gate290( .a(G820), .b(G821), .O(G847) );
nand2 gate291( .a(G822), .b(G823), .O(G860) );
nand2 gate292( .a(G824), .b(G825), .O(G873) );
nand2 gate293( .a(G828), .b(G829), .O(G886) );
nand2 gate294( .a(G832), .b(G833), .O(G899) );
nand2 gate295( .a(G830), .b(G831), .O(G912) );
nand2 gate296( .a(G826), .b(G827), .O(G925) );
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );
nand2 gate387( .a(G1), .b(G1036), .O(G1132) );
nand2 gate388( .a(G2), .b(G1039), .O(G1135) );
nand2 gate389( .a(G3), .b(G1042), .O(G1138) );
nand2 gate390( .a(G4), .b(G1045), .O(G1141) );
nand2 gate391( .a(G5), .b(G1048), .O(G1144) );
nand2 gate392( .a(G6), .b(G1051), .O(G1147) );
nand2 gate393( .a(G7), .b(G1054), .O(G1150) );
nand2 gate394( .a(G8), .b(G1057), .O(G1153) );
nand2 gate395( .a(G9), .b(G1060), .O(G1156) );

  xor2  gate981(.a(G1063), .b(G10), .O(gate396inter0));
  nand2 gate982(.a(gate396inter0), .b(s_62), .O(gate396inter1));
  and2  gate983(.a(G1063), .b(G10), .O(gate396inter2));
  inv1  gate984(.a(s_62), .O(gate396inter3));
  inv1  gate985(.a(s_63), .O(gate396inter4));
  nand2 gate986(.a(gate396inter4), .b(gate396inter3), .O(gate396inter5));
  nor2  gate987(.a(gate396inter5), .b(gate396inter2), .O(gate396inter6));
  inv1  gate988(.a(G10), .O(gate396inter7));
  inv1  gate989(.a(G1063), .O(gate396inter8));
  nand2 gate990(.a(gate396inter8), .b(gate396inter7), .O(gate396inter9));
  nand2 gate991(.a(s_63), .b(gate396inter3), .O(gate396inter10));
  nor2  gate992(.a(gate396inter10), .b(gate396inter9), .O(gate396inter11));
  nor2  gate993(.a(gate396inter11), .b(gate396inter6), .O(gate396inter12));
  nand2 gate994(.a(gate396inter12), .b(gate396inter1), .O(G1159));
nand2 gate397( .a(G11), .b(G1066), .O(G1162) );
nand2 gate398( .a(G12), .b(G1069), .O(G1165) );
nand2 gate399( .a(G13), .b(G1072), .O(G1168) );
nand2 gate400( .a(G14), .b(G1075), .O(G1171) );
nand2 gate401( .a(G15), .b(G1078), .O(G1174) );
nand2 gate402( .a(G16), .b(G1081), .O(G1177) );
nand2 gate403( .a(G17), .b(G1084), .O(G1180) );
nand2 gate404( .a(G18), .b(G1087), .O(G1183) );
nand2 gate405( .a(G19), .b(G1090), .O(G1186) );
nand2 gate406( .a(G20), .b(G1093), .O(G1189) );
nand2 gate407( .a(G21), .b(G1096), .O(G1192) );
nand2 gate408( .a(G22), .b(G1099), .O(G1195) );

  xor2  gate743(.a(G1102), .b(G23), .O(gate409inter0));
  nand2 gate744(.a(gate409inter0), .b(s_28), .O(gate409inter1));
  and2  gate745(.a(G1102), .b(G23), .O(gate409inter2));
  inv1  gate746(.a(s_28), .O(gate409inter3));
  inv1  gate747(.a(s_29), .O(gate409inter4));
  nand2 gate748(.a(gate409inter4), .b(gate409inter3), .O(gate409inter5));
  nor2  gate749(.a(gate409inter5), .b(gate409inter2), .O(gate409inter6));
  inv1  gate750(.a(G23), .O(gate409inter7));
  inv1  gate751(.a(G1102), .O(gate409inter8));
  nand2 gate752(.a(gate409inter8), .b(gate409inter7), .O(gate409inter9));
  nand2 gate753(.a(s_29), .b(gate409inter3), .O(gate409inter10));
  nor2  gate754(.a(gate409inter10), .b(gate409inter9), .O(gate409inter11));
  nor2  gate755(.a(gate409inter11), .b(gate409inter6), .O(gate409inter12));
  nand2 gate756(.a(gate409inter12), .b(gate409inter1), .O(G1198));
nand2 gate410( .a(G24), .b(G1105), .O(G1201) );
nand2 gate411( .a(G25), .b(G1108), .O(G1204) );
nand2 gate412( .a(G26), .b(G1111), .O(G1207) );
nand2 gate413( .a(G27), .b(G1114), .O(G1210) );
nand2 gate414( .a(G28), .b(G1117), .O(G1213) );
nand2 gate415( .a(G29), .b(G1120), .O(G1216) );
nand2 gate416( .a(G30), .b(G1123), .O(G1219) );
nand2 gate417( .a(G31), .b(G1126), .O(G1222) );
nand2 gate418( .a(G32), .b(G1129), .O(G1225) );
nand2 gate419( .a(G1), .b(G1132), .O(G1228) );

  xor2  gate561(.a(G1132), .b(G1036), .O(gate420inter0));
  nand2 gate562(.a(gate420inter0), .b(s_2), .O(gate420inter1));
  and2  gate563(.a(G1132), .b(G1036), .O(gate420inter2));
  inv1  gate564(.a(s_2), .O(gate420inter3));
  inv1  gate565(.a(s_3), .O(gate420inter4));
  nand2 gate566(.a(gate420inter4), .b(gate420inter3), .O(gate420inter5));
  nor2  gate567(.a(gate420inter5), .b(gate420inter2), .O(gate420inter6));
  inv1  gate568(.a(G1036), .O(gate420inter7));
  inv1  gate569(.a(G1132), .O(gate420inter8));
  nand2 gate570(.a(gate420inter8), .b(gate420inter7), .O(gate420inter9));
  nand2 gate571(.a(s_3), .b(gate420inter3), .O(gate420inter10));
  nor2  gate572(.a(gate420inter10), .b(gate420inter9), .O(gate420inter11));
  nor2  gate573(.a(gate420inter11), .b(gate420inter6), .O(gate420inter12));
  nand2 gate574(.a(gate420inter12), .b(gate420inter1), .O(G1229));
nand2 gate421( .a(G2), .b(G1135), .O(G1230) );
nand2 gate422( .a(G1039), .b(G1135), .O(G1231) );
nand2 gate423( .a(G3), .b(G1138), .O(G1232) );
nand2 gate424( .a(G1042), .b(G1138), .O(G1233) );
nand2 gate425( .a(G4), .b(G1141), .O(G1234) );
nand2 gate426( .a(G1045), .b(G1141), .O(G1235) );
nand2 gate427( .a(G5), .b(G1144), .O(G1236) );
nand2 gate428( .a(G1048), .b(G1144), .O(G1237) );
nand2 gate429( .a(G6), .b(G1147), .O(G1238) );
nand2 gate430( .a(G1051), .b(G1147), .O(G1239) );
nand2 gate431( .a(G7), .b(G1150), .O(G1240) );
nand2 gate432( .a(G1054), .b(G1150), .O(G1241) );
nand2 gate433( .a(G8), .b(G1153), .O(G1242) );
nand2 gate434( .a(G1057), .b(G1153), .O(G1243) );
nand2 gate435( .a(G9), .b(G1156), .O(G1244) );
nand2 gate436( .a(G1060), .b(G1156), .O(G1245) );
nand2 gate437( .a(G10), .b(G1159), .O(G1246) );
nand2 gate438( .a(G1063), .b(G1159), .O(G1247) );
nand2 gate439( .a(G11), .b(G1162), .O(G1248) );
nand2 gate440( .a(G1066), .b(G1162), .O(G1249) );

  xor2  gate1107(.a(G1165), .b(G12), .O(gate441inter0));
  nand2 gate1108(.a(gate441inter0), .b(s_80), .O(gate441inter1));
  and2  gate1109(.a(G1165), .b(G12), .O(gate441inter2));
  inv1  gate1110(.a(s_80), .O(gate441inter3));
  inv1  gate1111(.a(s_81), .O(gate441inter4));
  nand2 gate1112(.a(gate441inter4), .b(gate441inter3), .O(gate441inter5));
  nor2  gate1113(.a(gate441inter5), .b(gate441inter2), .O(gate441inter6));
  inv1  gate1114(.a(G12), .O(gate441inter7));
  inv1  gate1115(.a(G1165), .O(gate441inter8));
  nand2 gate1116(.a(gate441inter8), .b(gate441inter7), .O(gate441inter9));
  nand2 gate1117(.a(s_81), .b(gate441inter3), .O(gate441inter10));
  nor2  gate1118(.a(gate441inter10), .b(gate441inter9), .O(gate441inter11));
  nor2  gate1119(.a(gate441inter11), .b(gate441inter6), .O(gate441inter12));
  nand2 gate1120(.a(gate441inter12), .b(gate441inter1), .O(G1250));
nand2 gate442( .a(G1069), .b(G1165), .O(G1251) );
nand2 gate443( .a(G13), .b(G1168), .O(G1252) );
nand2 gate444( .a(G1072), .b(G1168), .O(G1253) );
nand2 gate445( .a(G14), .b(G1171), .O(G1254) );
nand2 gate446( .a(G1075), .b(G1171), .O(G1255) );
nand2 gate447( .a(G15), .b(G1174), .O(G1256) );
nand2 gate448( .a(G1078), .b(G1174), .O(G1257) );
nand2 gate449( .a(G16), .b(G1177), .O(G1258) );
nand2 gate450( .a(G1081), .b(G1177), .O(G1259) );
nand2 gate451( .a(G17), .b(G1180), .O(G1260) );
nand2 gate452( .a(G1084), .b(G1180), .O(G1261) );
nand2 gate453( .a(G18), .b(G1183), .O(G1262) );
nand2 gate454( .a(G1087), .b(G1183), .O(G1263) );
nand2 gate455( .a(G19), .b(G1186), .O(G1264) );
nand2 gate456( .a(G1090), .b(G1186), .O(G1265) );

  xor2  gate911(.a(G1189), .b(G20), .O(gate457inter0));
  nand2 gate912(.a(gate457inter0), .b(s_52), .O(gate457inter1));
  and2  gate913(.a(G1189), .b(G20), .O(gate457inter2));
  inv1  gate914(.a(s_52), .O(gate457inter3));
  inv1  gate915(.a(s_53), .O(gate457inter4));
  nand2 gate916(.a(gate457inter4), .b(gate457inter3), .O(gate457inter5));
  nor2  gate917(.a(gate457inter5), .b(gate457inter2), .O(gate457inter6));
  inv1  gate918(.a(G20), .O(gate457inter7));
  inv1  gate919(.a(G1189), .O(gate457inter8));
  nand2 gate920(.a(gate457inter8), .b(gate457inter7), .O(gate457inter9));
  nand2 gate921(.a(s_53), .b(gate457inter3), .O(gate457inter10));
  nor2  gate922(.a(gate457inter10), .b(gate457inter9), .O(gate457inter11));
  nor2  gate923(.a(gate457inter11), .b(gate457inter6), .O(gate457inter12));
  nand2 gate924(.a(gate457inter12), .b(gate457inter1), .O(G1266));
nand2 gate458( .a(G1093), .b(G1189), .O(G1267) );
nand2 gate459( .a(G21), .b(G1192), .O(G1268) );
nand2 gate460( .a(G1096), .b(G1192), .O(G1269) );
nand2 gate461( .a(G22), .b(G1195), .O(G1270) );
nand2 gate462( .a(G1099), .b(G1195), .O(G1271) );
nand2 gate463( .a(G23), .b(G1198), .O(G1272) );
nand2 gate464( .a(G1102), .b(G1198), .O(G1273) );
nand2 gate465( .a(G24), .b(G1201), .O(G1274) );
nand2 gate466( .a(G1105), .b(G1201), .O(G1275) );
nand2 gate467( .a(G25), .b(G1204), .O(G1276) );

  xor2  gate1065(.a(G1204), .b(G1108), .O(gate468inter0));
  nand2 gate1066(.a(gate468inter0), .b(s_74), .O(gate468inter1));
  and2  gate1067(.a(G1204), .b(G1108), .O(gate468inter2));
  inv1  gate1068(.a(s_74), .O(gate468inter3));
  inv1  gate1069(.a(s_75), .O(gate468inter4));
  nand2 gate1070(.a(gate468inter4), .b(gate468inter3), .O(gate468inter5));
  nor2  gate1071(.a(gate468inter5), .b(gate468inter2), .O(gate468inter6));
  inv1  gate1072(.a(G1108), .O(gate468inter7));
  inv1  gate1073(.a(G1204), .O(gate468inter8));
  nand2 gate1074(.a(gate468inter8), .b(gate468inter7), .O(gate468inter9));
  nand2 gate1075(.a(s_75), .b(gate468inter3), .O(gate468inter10));
  nor2  gate1076(.a(gate468inter10), .b(gate468inter9), .O(gate468inter11));
  nor2  gate1077(.a(gate468inter11), .b(gate468inter6), .O(gate468inter12));
  nand2 gate1078(.a(gate468inter12), .b(gate468inter1), .O(G1277));

  xor2  gate1023(.a(G1207), .b(G26), .O(gate469inter0));
  nand2 gate1024(.a(gate469inter0), .b(s_68), .O(gate469inter1));
  and2  gate1025(.a(G1207), .b(G26), .O(gate469inter2));
  inv1  gate1026(.a(s_68), .O(gate469inter3));
  inv1  gate1027(.a(s_69), .O(gate469inter4));
  nand2 gate1028(.a(gate469inter4), .b(gate469inter3), .O(gate469inter5));
  nor2  gate1029(.a(gate469inter5), .b(gate469inter2), .O(gate469inter6));
  inv1  gate1030(.a(G26), .O(gate469inter7));
  inv1  gate1031(.a(G1207), .O(gate469inter8));
  nand2 gate1032(.a(gate469inter8), .b(gate469inter7), .O(gate469inter9));
  nand2 gate1033(.a(s_69), .b(gate469inter3), .O(gate469inter10));
  nor2  gate1034(.a(gate469inter10), .b(gate469inter9), .O(gate469inter11));
  nor2  gate1035(.a(gate469inter11), .b(gate469inter6), .O(gate469inter12));
  nand2 gate1036(.a(gate469inter12), .b(gate469inter1), .O(G1278));
nand2 gate470( .a(G1111), .b(G1207), .O(G1279) );
nand2 gate471( .a(G27), .b(G1210), .O(G1280) );
nand2 gate472( .a(G1114), .b(G1210), .O(G1281) );
nand2 gate473( .a(G28), .b(G1213), .O(G1282) );
nand2 gate474( .a(G1117), .b(G1213), .O(G1283) );
nand2 gate475( .a(G29), .b(G1216), .O(G1284) );
nand2 gate476( .a(G1120), .b(G1216), .O(G1285) );
nand2 gate477( .a(G30), .b(G1219), .O(G1286) );
nand2 gate478( .a(G1123), .b(G1219), .O(G1287) );
nand2 gate479( .a(G31), .b(G1222), .O(G1288) );
nand2 gate480( .a(G1126), .b(G1222), .O(G1289) );
nand2 gate481( .a(G32), .b(G1225), .O(G1290) );
nand2 gate482( .a(G1129), .b(G1225), .O(G1291) );
nand2 gate483( .a(G1228), .b(G1229), .O(G1292) );
nand2 gate484( .a(G1230), .b(G1231), .O(G1293) );
nand2 gate485( .a(G1232), .b(G1233), .O(G1294) );
nand2 gate486( .a(G1234), .b(G1235), .O(G1295) );
nand2 gate487( .a(G1236), .b(G1237), .O(G1296) );
nand2 gate488( .a(G1238), .b(G1239), .O(G1297) );
nand2 gate489( .a(G1240), .b(G1241), .O(G1298) );
nand2 gate490( .a(G1242), .b(G1243), .O(G1299) );
nand2 gate491( .a(G1244), .b(G1245), .O(G1300) );
nand2 gate492( .a(G1246), .b(G1247), .O(G1301) );
nand2 gate493( .a(G1248), .b(G1249), .O(G1302) );
nand2 gate494( .a(G1250), .b(G1251), .O(G1303) );
nand2 gate495( .a(G1252), .b(G1253), .O(G1304) );
nand2 gate496( .a(G1254), .b(G1255), .O(G1305) );
nand2 gate497( .a(G1256), .b(G1257), .O(G1306) );
nand2 gate498( .a(G1258), .b(G1259), .O(G1307) );
nand2 gate499( .a(G1260), .b(G1261), .O(G1308) );
nand2 gate500( .a(G1262), .b(G1263), .O(G1309) );
nand2 gate501( .a(G1264), .b(G1265), .O(G1310) );
nand2 gate502( .a(G1266), .b(G1267), .O(G1311) );
nand2 gate503( .a(G1268), .b(G1269), .O(G1312) );
nand2 gate504( .a(G1270), .b(G1271), .O(G1313) );

  xor2  gate1009(.a(G1273), .b(G1272), .O(gate505inter0));
  nand2 gate1010(.a(gate505inter0), .b(s_66), .O(gate505inter1));
  and2  gate1011(.a(G1273), .b(G1272), .O(gate505inter2));
  inv1  gate1012(.a(s_66), .O(gate505inter3));
  inv1  gate1013(.a(s_67), .O(gate505inter4));
  nand2 gate1014(.a(gate505inter4), .b(gate505inter3), .O(gate505inter5));
  nor2  gate1015(.a(gate505inter5), .b(gate505inter2), .O(gate505inter6));
  inv1  gate1016(.a(G1272), .O(gate505inter7));
  inv1  gate1017(.a(G1273), .O(gate505inter8));
  nand2 gate1018(.a(gate505inter8), .b(gate505inter7), .O(gate505inter9));
  nand2 gate1019(.a(s_67), .b(gate505inter3), .O(gate505inter10));
  nor2  gate1020(.a(gate505inter10), .b(gate505inter9), .O(gate505inter11));
  nor2  gate1021(.a(gate505inter11), .b(gate505inter6), .O(gate505inter12));
  nand2 gate1022(.a(gate505inter12), .b(gate505inter1), .O(G1314));
nand2 gate506( .a(G1274), .b(G1275), .O(G1315) );
nand2 gate507( .a(G1276), .b(G1277), .O(G1316) );
nand2 gate508( .a(G1278), .b(G1279), .O(G1317) );
nand2 gate509( .a(G1280), .b(G1281), .O(G1318) );
nand2 gate510( .a(G1282), .b(G1283), .O(G1319) );
nand2 gate511( .a(G1284), .b(G1285), .O(G1320) );
nand2 gate512( .a(G1286), .b(G1287), .O(G1321) );
nand2 gate513( .a(G1288), .b(G1289), .O(G1322) );
nand2 gate514( .a(G1290), .b(G1291), .O(G1323) );
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule