module c499 (N1,N5,N9,N13,N17,N21,N25,N29,N33,N37,
             N41,N45,N49,N53,N57,N61,N65,N69,N73,N77,
             N81,N85,N89,N93,N97,N101,N105,N109,N113,N117,
             N121,N125,N129,N130,N131,N132,N133,N134,N135,N136,
             N137,N724,N725,N726,N727,N728,N729,N730,N731,N732,
             N733,N734,N735,N736,N737,N738,N739,N740,N741,N742,
             N743,N744,N745,N746,N747,N748,N749,N750,N751,N752,
             N753,N754,N755);

input N1,N5,N9,N13,N17,N21,N25,N29,N33,N37,
      N41,N45,N49,N53,N57,N61,N65,N69,N73,N77,
      N81,N85,N89,N93,N97,N101,N105,N109,N113,N117,
      N121,N125,N129,N130,N131,N132,N133,N134,N135,N136,
      N137;//RE__PI;

input s_0,s_1;//RE__ALLOW(00,01,10,11);
input s_2,s_3;//RE__ALLOW(00,01,10,11);
input s_4,s_5;//RE__ALLOW(00,01,10,11);
input s_6,s_7;//RE__ALLOW(00,01,10,11);
input s_8,s_9;//RE__ALLOW(00,01,10,11);
input s_10,s_11;//RE__ALLOW(00,01,10,11);
input s_12,s_13;//RE__ALLOW(00,01,10,11);
input s_14,s_15;//RE__ALLOW(00,01,10,11);
input s_16,s_17;//RE__ALLOW(00,01,10,11);
input s_18,s_19;//RE__ALLOW(00,01,10,11);
input s_20,s_21;//RE__ALLOW(00,01,10,11);
input s_22,s_23;//RE__ALLOW(00,01,10,11);
input s_24,s_25;//RE__ALLOW(00,01,10,11);
input s_26,s_27;//RE__ALLOW(00,01,10,11);
input s_28,s_29;//RE__ALLOW(00,01,10,11);
input s_30,s_31;//RE__ALLOW(00,01,10,11);
input s_32,s_33;//RE__ALLOW(00,01,10,11);
input s_34,s_35;//RE__ALLOW(00,01,10,11);
input s_36,s_37;//RE__ALLOW(00,01,10,11);
input s_38,s_39;//RE__ALLOW(00,01,10,11);
input s_40,s_41;//RE__ALLOW(00,01,10,11);
output N724,N725,N726,N727,N728,N729,N730,N731,N732,N733,
       N734,N735,N736,N737,N738,N739,N740,N741,N742,N743,
       N744,N745,N746,N747,N748,N749,N750,N751,N752,N753,
       N754,N755;

wire N250,N251,N252,N253,N254,N255,N256,N257,N258,N259,
     N260,N261,N262,N263,N264,N265,N266,N267,N268,N269,
     N270,N271,N272,N273,N274,N275,N276,N277,N278,N279,
     N280,N281,N282,N283,N284,N285,N286,N287,N288,N289,
     N290,N293,N296,N299,N302,N305,N308,N311,N314,N315,
     N316,N317,N318,N319,N320,N321,N338,N339,N340,N341,
     N342,N343,N344,N345,N346,N347,N348,N349,N350,N351,
     N352,N353,N354,N367,N380,N393,N406,N419,N432,N445,
     N554,N555,N556,N557,N558,N559,N560,N561,N562,N563,
     N564,N565,N566,N567,N568,N569,N570,N571,N572,N573,
     N574,N575,N576,N577,N578,N579,N580,N581,N582,N583,
     N584,N585,N586,N587,N588,N589,N590,N591,N592,N593,
     N594,N595,N596,N597,N598,N599,N600,N601,N602,N607,
     N620,N625,N630,N635,N640,N645,N650,N655,N692,N693,
     N694,N695,N696,N697,N698,N699,N700,N701,N702,N703,
     N704,N705,N706,N707,N708,N709,N710,N711,N712,N713,
     N714,N715,N716,N717,N718,N719,N720,N721,N722,N723, gate14inter0, gate14inter1, gate14inter2, gate14inter3, gate14inter4, gate14inter5, gate14inter6, gate14inter7, gate14inter8, gate14inter9, gate14inter10, gate14inter11, gate14inter12, gate35inter0, gate35inter1, gate35inter2, gate35inter3, gate35inter4, gate35inter5, gate35inter6, gate35inter7, gate35inter8, gate35inter9, gate35inter10, gate35inter11, gate35inter12, gate188inter0, gate188inter1, gate188inter2, gate188inter3, gate188inter4, gate188inter5, gate188inter6, gate188inter7, gate188inter8, gate188inter9, gate188inter10, gate188inter11, gate188inter12, gate184inter0, gate184inter1, gate184inter2, gate184inter3, gate184inter4, gate184inter5, gate184inter6, gate184inter7, gate184inter8, gate184inter9, gate184inter10, gate184inter11, gate184inter12, gate193inter0, gate193inter1, gate193inter2, gate193inter3, gate193inter4, gate193inter5, gate193inter6, gate193inter7, gate193inter8, gate193inter9, gate193inter10, gate193inter11, gate193inter12, gate42inter0, gate42inter1, gate42inter2, gate42inter3, gate42inter4, gate42inter5, gate42inter6, gate42inter7, gate42inter8, gate42inter9, gate42inter10, gate42inter11, gate42inter12, gate45inter0, gate45inter1, gate45inter2, gate45inter3, gate45inter4, gate45inter5, gate45inter6, gate45inter7, gate45inter8, gate45inter9, gate45inter10, gate45inter11, gate45inter12, gate11inter0, gate11inter1, gate11inter2, gate11inter3, gate11inter4, gate11inter5, gate11inter6, gate11inter7, gate11inter8, gate11inter9, gate11inter10, gate11inter11, gate11inter12, gate29inter0, gate29inter1, gate29inter2, gate29inter3, gate29inter4, gate29inter5, gate29inter6, gate29inter7, gate29inter8, gate29inter9, gate29inter10, gate29inter11, gate29inter12, gate40inter0, gate40inter1, gate40inter2, gate40inter3, gate40inter4, gate40inter5, gate40inter6, gate40inter7, gate40inter8, gate40inter9, gate40inter10, gate40inter11, gate40inter12, gate197inter0, gate197inter1, gate197inter2, gate197inter3, gate197inter4, gate197inter5, gate197inter6, gate197inter7, gate197inter8, gate197inter9, gate197inter10, gate197inter11, gate197inter12, gate78inter0, gate78inter1, gate78inter2, gate78inter3, gate78inter4, gate78inter5, gate78inter6, gate78inter7, gate78inter8, gate78inter9, gate78inter10, gate78inter11, gate78inter12, gate80inter0, gate80inter1, gate80inter2, gate80inter3, gate80inter4, gate80inter5, gate80inter6, gate80inter7, gate80inter8, gate80inter9, gate80inter10, gate80inter11, gate80inter12, gate189inter0, gate189inter1, gate189inter2, gate189inter3, gate189inter4, gate189inter5, gate189inter6, gate189inter7, gate189inter8, gate189inter9, gate189inter10, gate189inter11, gate189inter12, gate36inter0, gate36inter1, gate36inter2, gate36inter3, gate36inter4, gate36inter5, gate36inter6, gate36inter7, gate36inter8, gate36inter9, gate36inter10, gate36inter11, gate36inter12, gate49inter0, gate49inter1, gate49inter2, gate49inter3, gate49inter4, gate49inter5, gate49inter6, gate49inter7, gate49inter8, gate49inter9, gate49inter10, gate49inter11, gate49inter12, gate192inter0, gate192inter1, gate192inter2, gate192inter3, gate192inter4, gate192inter5, gate192inter6, gate192inter7, gate192inter8, gate192inter9, gate192inter10, gate192inter11, gate192inter12, gate62inter0, gate62inter1, gate62inter2, gate62inter3, gate62inter4, gate62inter5, gate62inter6, gate62inter7, gate62inter8, gate62inter9, gate62inter10, gate62inter11, gate62inter12, gate198inter0, gate198inter1, gate198inter2, gate198inter3, gate198inter4, gate198inter5, gate198inter6, gate198inter7, gate198inter8, gate198inter9, gate198inter10, gate198inter11, gate198inter12, gate171inter0, gate171inter1, gate171inter2, gate171inter3, gate171inter4, gate171inter5, gate171inter6, gate171inter7, gate171inter8, gate171inter9, gate171inter10, gate171inter11, gate171inter12, gate3inter0, gate3inter1, gate3inter2, gate3inter3, gate3inter4, gate3inter5, gate3inter6, gate3inter7, gate3inter8, gate3inter9, gate3inter10, gate3inter11, gate3inter12;



xor2 gate1( .a(N1), .b(N5), .O(N250) );
xor2 gate2( .a(N9), .b(N13), .O(N251) );

  xor2  gate483(.a(N21), .b(N17), .O(gate3inter0));
  nand2 gate484(.a(gate3inter0), .b(s_40), .O(gate3inter1));
  and2  gate485(.a(N21), .b(N17), .O(gate3inter2));
  inv1  gate486(.a(s_40), .O(gate3inter3));
  inv1  gate487(.a(s_41), .O(gate3inter4));
  nand2 gate488(.a(gate3inter4), .b(gate3inter3), .O(gate3inter5));
  nor2  gate489(.a(gate3inter5), .b(gate3inter2), .O(gate3inter6));
  inv1  gate490(.a(N17), .O(gate3inter7));
  inv1  gate491(.a(N21), .O(gate3inter8));
  nand2 gate492(.a(gate3inter8), .b(gate3inter7), .O(gate3inter9));
  nand2 gate493(.a(s_41), .b(gate3inter3), .O(gate3inter10));
  nor2  gate494(.a(gate3inter10), .b(gate3inter9), .O(gate3inter11));
  nor2  gate495(.a(gate3inter11), .b(gate3inter6), .O(gate3inter12));
  nand2 gate496(.a(gate3inter12), .b(gate3inter1), .O(N252));
xor2 gate4( .a(N25), .b(N29), .O(N253) );
xor2 gate5( .a(N33), .b(N37), .O(N254) );
xor2 gate6( .a(N41), .b(N45), .O(N255) );
xor2 gate7( .a(N49), .b(N53), .O(N256) );
xor2 gate8( .a(N57), .b(N61), .O(N257) );
xor2 gate9( .a(N65), .b(N69), .O(N258) );
xor2 gate10( .a(N73), .b(N77), .O(N259) );

  xor2  gate301(.a(N85), .b(N81), .O(gate11inter0));
  nand2 gate302(.a(gate11inter0), .b(s_14), .O(gate11inter1));
  and2  gate303(.a(N85), .b(N81), .O(gate11inter2));
  inv1  gate304(.a(s_14), .O(gate11inter3));
  inv1  gate305(.a(s_15), .O(gate11inter4));
  nand2 gate306(.a(gate11inter4), .b(gate11inter3), .O(gate11inter5));
  nor2  gate307(.a(gate11inter5), .b(gate11inter2), .O(gate11inter6));
  inv1  gate308(.a(N81), .O(gate11inter7));
  inv1  gate309(.a(N85), .O(gate11inter8));
  nand2 gate310(.a(gate11inter8), .b(gate11inter7), .O(gate11inter9));
  nand2 gate311(.a(s_15), .b(gate11inter3), .O(gate11inter10));
  nor2  gate312(.a(gate11inter10), .b(gate11inter9), .O(gate11inter11));
  nor2  gate313(.a(gate11inter11), .b(gate11inter6), .O(gate11inter12));
  nand2 gate314(.a(gate11inter12), .b(gate11inter1), .O(N260));
xor2 gate12( .a(N89), .b(N93), .O(N261) );
xor2 gate13( .a(N97), .b(N101), .O(N262) );

  xor2  gate203(.a(N109), .b(N105), .O(gate14inter0));
  nand2 gate204(.a(gate14inter0), .b(s_0), .O(gate14inter1));
  and2  gate205(.a(N109), .b(N105), .O(gate14inter2));
  inv1  gate206(.a(s_0), .O(gate14inter3));
  inv1  gate207(.a(s_1), .O(gate14inter4));
  nand2 gate208(.a(gate14inter4), .b(gate14inter3), .O(gate14inter5));
  nor2  gate209(.a(gate14inter5), .b(gate14inter2), .O(gate14inter6));
  inv1  gate210(.a(N105), .O(gate14inter7));
  inv1  gate211(.a(N109), .O(gate14inter8));
  nand2 gate212(.a(gate14inter8), .b(gate14inter7), .O(gate14inter9));
  nand2 gate213(.a(s_1), .b(gate14inter3), .O(gate14inter10));
  nor2  gate214(.a(gate14inter10), .b(gate14inter9), .O(gate14inter11));
  nor2  gate215(.a(gate14inter11), .b(gate14inter6), .O(gate14inter12));
  nand2 gate216(.a(gate14inter12), .b(gate14inter1), .O(N263));
xor2 gate15( .a(N113), .b(N117), .O(N264) );
xor2 gate16( .a(N121), .b(N125), .O(N265) );
and2 gate17( .a(N129), .b(N137), .O(N266) );
and2 gate18( .a(N130), .b(N137), .O(N267) );
and2 gate19( .a(N131), .b(N137), .O(N268) );
and2 gate20( .a(N132), .b(N137), .O(N269) );
and2 gate21( .a(N133), .b(N137), .O(N270) );
and2 gate22( .a(N134), .b(N137), .O(N271) );
and2 gate23( .a(N135), .b(N137), .O(N272) );
and2 gate24( .a(N136), .b(N137), .O(N273) );
xor2 gate25( .a(N1), .b(N17), .O(N274) );
xor2 gate26( .a(N33), .b(N49), .O(N275) );
xor2 gate27( .a(N5), .b(N21), .O(N276) );
xor2 gate28( .a(N37), .b(N53), .O(N277) );

  xor2  gate315(.a(N25), .b(N9), .O(gate29inter0));
  nand2 gate316(.a(gate29inter0), .b(s_16), .O(gate29inter1));
  and2  gate317(.a(N25), .b(N9), .O(gate29inter2));
  inv1  gate318(.a(s_16), .O(gate29inter3));
  inv1  gate319(.a(s_17), .O(gate29inter4));
  nand2 gate320(.a(gate29inter4), .b(gate29inter3), .O(gate29inter5));
  nor2  gate321(.a(gate29inter5), .b(gate29inter2), .O(gate29inter6));
  inv1  gate322(.a(N9), .O(gate29inter7));
  inv1  gate323(.a(N25), .O(gate29inter8));
  nand2 gate324(.a(gate29inter8), .b(gate29inter7), .O(gate29inter9));
  nand2 gate325(.a(s_17), .b(gate29inter3), .O(gate29inter10));
  nor2  gate326(.a(gate29inter10), .b(gate29inter9), .O(gate29inter11));
  nor2  gate327(.a(gate29inter11), .b(gate29inter6), .O(gate29inter12));
  nand2 gate328(.a(gate29inter12), .b(gate29inter1), .O(N278));
xor2 gate30( .a(N41), .b(N57), .O(N279) );
xor2 gate31( .a(N13), .b(N29), .O(N280) );
xor2 gate32( .a(N45), .b(N61), .O(N281) );
xor2 gate33( .a(N65), .b(N81), .O(N282) );
xor2 gate34( .a(N97), .b(N113), .O(N283) );

  xor2  gate217(.a(N85), .b(N69), .O(gate35inter0));
  nand2 gate218(.a(gate35inter0), .b(s_2), .O(gate35inter1));
  and2  gate219(.a(N85), .b(N69), .O(gate35inter2));
  inv1  gate220(.a(s_2), .O(gate35inter3));
  inv1  gate221(.a(s_3), .O(gate35inter4));
  nand2 gate222(.a(gate35inter4), .b(gate35inter3), .O(gate35inter5));
  nor2  gate223(.a(gate35inter5), .b(gate35inter2), .O(gate35inter6));
  inv1  gate224(.a(N69), .O(gate35inter7));
  inv1  gate225(.a(N85), .O(gate35inter8));
  nand2 gate226(.a(gate35inter8), .b(gate35inter7), .O(gate35inter9));
  nand2 gate227(.a(s_3), .b(gate35inter3), .O(gate35inter10));
  nor2  gate228(.a(gate35inter10), .b(gate35inter9), .O(gate35inter11));
  nor2  gate229(.a(gate35inter11), .b(gate35inter6), .O(gate35inter12));
  nand2 gate230(.a(gate35inter12), .b(gate35inter1), .O(N284));

  xor2  gate399(.a(N117), .b(N101), .O(gate36inter0));
  nand2 gate400(.a(gate36inter0), .b(s_28), .O(gate36inter1));
  and2  gate401(.a(N117), .b(N101), .O(gate36inter2));
  inv1  gate402(.a(s_28), .O(gate36inter3));
  inv1  gate403(.a(s_29), .O(gate36inter4));
  nand2 gate404(.a(gate36inter4), .b(gate36inter3), .O(gate36inter5));
  nor2  gate405(.a(gate36inter5), .b(gate36inter2), .O(gate36inter6));
  inv1  gate406(.a(N101), .O(gate36inter7));
  inv1  gate407(.a(N117), .O(gate36inter8));
  nand2 gate408(.a(gate36inter8), .b(gate36inter7), .O(gate36inter9));
  nand2 gate409(.a(s_29), .b(gate36inter3), .O(gate36inter10));
  nor2  gate410(.a(gate36inter10), .b(gate36inter9), .O(gate36inter11));
  nor2  gate411(.a(gate36inter11), .b(gate36inter6), .O(gate36inter12));
  nand2 gate412(.a(gate36inter12), .b(gate36inter1), .O(N285));
xor2 gate37( .a(N73), .b(N89), .O(N286) );
xor2 gate38( .a(N105), .b(N121), .O(N287) );
xor2 gate39( .a(N77), .b(N93), .O(N288) );

  xor2  gate329(.a(N125), .b(N109), .O(gate40inter0));
  nand2 gate330(.a(gate40inter0), .b(s_18), .O(gate40inter1));
  and2  gate331(.a(N125), .b(N109), .O(gate40inter2));
  inv1  gate332(.a(s_18), .O(gate40inter3));
  inv1  gate333(.a(s_19), .O(gate40inter4));
  nand2 gate334(.a(gate40inter4), .b(gate40inter3), .O(gate40inter5));
  nor2  gate335(.a(gate40inter5), .b(gate40inter2), .O(gate40inter6));
  inv1  gate336(.a(N109), .O(gate40inter7));
  inv1  gate337(.a(N125), .O(gate40inter8));
  nand2 gate338(.a(gate40inter8), .b(gate40inter7), .O(gate40inter9));
  nand2 gate339(.a(s_19), .b(gate40inter3), .O(gate40inter10));
  nor2  gate340(.a(gate40inter10), .b(gate40inter9), .O(gate40inter11));
  nor2  gate341(.a(gate40inter11), .b(gate40inter6), .O(gate40inter12));
  nand2 gate342(.a(gate40inter12), .b(gate40inter1), .O(N289));
xor2 gate41( .a(N250), .b(N251), .O(N290) );

  xor2  gate273(.a(N253), .b(N252), .O(gate42inter0));
  nand2 gate274(.a(gate42inter0), .b(s_10), .O(gate42inter1));
  and2  gate275(.a(N253), .b(N252), .O(gate42inter2));
  inv1  gate276(.a(s_10), .O(gate42inter3));
  inv1  gate277(.a(s_11), .O(gate42inter4));
  nand2 gate278(.a(gate42inter4), .b(gate42inter3), .O(gate42inter5));
  nor2  gate279(.a(gate42inter5), .b(gate42inter2), .O(gate42inter6));
  inv1  gate280(.a(N252), .O(gate42inter7));
  inv1  gate281(.a(N253), .O(gate42inter8));
  nand2 gate282(.a(gate42inter8), .b(gate42inter7), .O(gate42inter9));
  nand2 gate283(.a(s_11), .b(gate42inter3), .O(gate42inter10));
  nor2  gate284(.a(gate42inter10), .b(gate42inter9), .O(gate42inter11));
  nor2  gate285(.a(gate42inter11), .b(gate42inter6), .O(gate42inter12));
  nand2 gate286(.a(gate42inter12), .b(gate42inter1), .O(N293));
xor2 gate43( .a(N254), .b(N255), .O(N296) );
xor2 gate44( .a(N256), .b(N257), .O(N299) );

  xor2  gate287(.a(N259), .b(N258), .O(gate45inter0));
  nand2 gate288(.a(gate45inter0), .b(s_12), .O(gate45inter1));
  and2  gate289(.a(N259), .b(N258), .O(gate45inter2));
  inv1  gate290(.a(s_12), .O(gate45inter3));
  inv1  gate291(.a(s_13), .O(gate45inter4));
  nand2 gate292(.a(gate45inter4), .b(gate45inter3), .O(gate45inter5));
  nor2  gate293(.a(gate45inter5), .b(gate45inter2), .O(gate45inter6));
  inv1  gate294(.a(N258), .O(gate45inter7));
  inv1  gate295(.a(N259), .O(gate45inter8));
  nand2 gate296(.a(gate45inter8), .b(gate45inter7), .O(gate45inter9));
  nand2 gate297(.a(s_13), .b(gate45inter3), .O(gate45inter10));
  nor2  gate298(.a(gate45inter10), .b(gate45inter9), .O(gate45inter11));
  nor2  gate299(.a(gate45inter11), .b(gate45inter6), .O(gate45inter12));
  nand2 gate300(.a(gate45inter12), .b(gate45inter1), .O(N302));
xor2 gate46( .a(N260), .b(N261), .O(N305) );
xor2 gate47( .a(N262), .b(N263), .O(N308) );
xor2 gate48( .a(N264), .b(N265), .O(N311) );

  xor2  gate413(.a(N275), .b(N274), .O(gate49inter0));
  nand2 gate414(.a(gate49inter0), .b(s_30), .O(gate49inter1));
  and2  gate415(.a(N275), .b(N274), .O(gate49inter2));
  inv1  gate416(.a(s_30), .O(gate49inter3));
  inv1  gate417(.a(s_31), .O(gate49inter4));
  nand2 gate418(.a(gate49inter4), .b(gate49inter3), .O(gate49inter5));
  nor2  gate419(.a(gate49inter5), .b(gate49inter2), .O(gate49inter6));
  inv1  gate420(.a(N274), .O(gate49inter7));
  inv1  gate421(.a(N275), .O(gate49inter8));
  nand2 gate422(.a(gate49inter8), .b(gate49inter7), .O(gate49inter9));
  nand2 gate423(.a(s_31), .b(gate49inter3), .O(gate49inter10));
  nor2  gate424(.a(gate49inter10), .b(gate49inter9), .O(gate49inter11));
  nor2  gate425(.a(gate49inter11), .b(gate49inter6), .O(gate49inter12));
  nand2 gate426(.a(gate49inter12), .b(gate49inter1), .O(N314));
xor2 gate50( .a(N276), .b(N277), .O(N315) );
xor2 gate51( .a(N278), .b(N279), .O(N316) );
xor2 gate52( .a(N280), .b(N281), .O(N317) );
xor2 gate53( .a(N282), .b(N283), .O(N318) );
xor2 gate54( .a(N284), .b(N285), .O(N319) );
xor2 gate55( .a(N286), .b(N287), .O(N320) );
xor2 gate56( .a(N288), .b(N289), .O(N321) );
xor2 gate57( .a(N290), .b(N293), .O(N338) );
xor2 gate58( .a(N296), .b(N299), .O(N339) );
xor2 gate59( .a(N290), .b(N296), .O(N340) );
xor2 gate60( .a(N293), .b(N299), .O(N341) );
xor2 gate61( .a(N302), .b(N305), .O(N342) );

  xor2  gate441(.a(N311), .b(N308), .O(gate62inter0));
  nand2 gate442(.a(gate62inter0), .b(s_34), .O(gate62inter1));
  and2  gate443(.a(N311), .b(N308), .O(gate62inter2));
  inv1  gate444(.a(s_34), .O(gate62inter3));
  inv1  gate445(.a(s_35), .O(gate62inter4));
  nand2 gate446(.a(gate62inter4), .b(gate62inter3), .O(gate62inter5));
  nor2  gate447(.a(gate62inter5), .b(gate62inter2), .O(gate62inter6));
  inv1  gate448(.a(N308), .O(gate62inter7));
  inv1  gate449(.a(N311), .O(gate62inter8));
  nand2 gate450(.a(gate62inter8), .b(gate62inter7), .O(gate62inter9));
  nand2 gate451(.a(s_35), .b(gate62inter3), .O(gate62inter10));
  nor2  gate452(.a(gate62inter10), .b(gate62inter9), .O(gate62inter11));
  nor2  gate453(.a(gate62inter11), .b(gate62inter6), .O(gate62inter12));
  nand2 gate454(.a(gate62inter12), .b(gate62inter1), .O(N343));
xor2 gate63( .a(N302), .b(N308), .O(N344) );
xor2 gate64( .a(N305), .b(N311), .O(N345) );
xor2 gate65( .a(N266), .b(N342), .O(N346) );
xor2 gate66( .a(N267), .b(N343), .O(N347) );
xor2 gate67( .a(N268), .b(N344), .O(N348) );
xor2 gate68( .a(N269), .b(N345), .O(N349) );
xor2 gate69( .a(N270), .b(N338), .O(N350) );
xor2 gate70( .a(N271), .b(N339), .O(N351) );
xor2 gate71( .a(N272), .b(N340), .O(N352) );
xor2 gate72( .a(N273), .b(N341), .O(N353) );
xor2 gate73( .a(N314), .b(N346), .O(N354) );
xor2 gate74( .a(N315), .b(N347), .O(N367) );
xor2 gate75( .a(N316), .b(N348), .O(N380) );
xor2 gate76( .a(N317), .b(N349), .O(N393) );
xor2 gate77( .a(N318), .b(N350), .O(N406) );

  xor2  gate357(.a(N351), .b(N319), .O(gate78inter0));
  nand2 gate358(.a(gate78inter0), .b(s_22), .O(gate78inter1));
  and2  gate359(.a(N351), .b(N319), .O(gate78inter2));
  inv1  gate360(.a(s_22), .O(gate78inter3));
  inv1  gate361(.a(s_23), .O(gate78inter4));
  nand2 gate362(.a(gate78inter4), .b(gate78inter3), .O(gate78inter5));
  nor2  gate363(.a(gate78inter5), .b(gate78inter2), .O(gate78inter6));
  inv1  gate364(.a(N319), .O(gate78inter7));
  inv1  gate365(.a(N351), .O(gate78inter8));
  nand2 gate366(.a(gate78inter8), .b(gate78inter7), .O(gate78inter9));
  nand2 gate367(.a(s_23), .b(gate78inter3), .O(gate78inter10));
  nor2  gate368(.a(gate78inter10), .b(gate78inter9), .O(gate78inter11));
  nor2  gate369(.a(gate78inter11), .b(gate78inter6), .O(gate78inter12));
  nand2 gate370(.a(gate78inter12), .b(gate78inter1), .O(N419));
xor2 gate79( .a(N320), .b(N352), .O(N432) );

  xor2  gate371(.a(N353), .b(N321), .O(gate80inter0));
  nand2 gate372(.a(gate80inter0), .b(s_24), .O(gate80inter1));
  and2  gate373(.a(N353), .b(N321), .O(gate80inter2));
  inv1  gate374(.a(s_24), .O(gate80inter3));
  inv1  gate375(.a(s_25), .O(gate80inter4));
  nand2 gate376(.a(gate80inter4), .b(gate80inter3), .O(gate80inter5));
  nor2  gate377(.a(gate80inter5), .b(gate80inter2), .O(gate80inter6));
  inv1  gate378(.a(N321), .O(gate80inter7));
  inv1  gate379(.a(N353), .O(gate80inter8));
  nand2 gate380(.a(gate80inter8), .b(gate80inter7), .O(gate80inter9));
  nand2 gate381(.a(s_25), .b(gate80inter3), .O(gate80inter10));
  nor2  gate382(.a(gate80inter10), .b(gate80inter9), .O(gate80inter11));
  nor2  gate383(.a(gate80inter11), .b(gate80inter6), .O(gate80inter12));
  nand2 gate384(.a(gate80inter12), .b(gate80inter1), .O(N445));
inv1 gate81( .a(N354), .O(N554) );
inv1 gate82( .a(N367), .O(N555) );
inv1 gate83( .a(N380), .O(N556) );
inv1 gate84( .a(N354), .O(N557) );
inv1 gate85( .a(N367), .O(N558) );
inv1 gate86( .a(N393), .O(N559) );
inv1 gate87( .a(N354), .O(N560) );
inv1 gate88( .a(N380), .O(N561) );
inv1 gate89( .a(N393), .O(N562) );
inv1 gate90( .a(N367), .O(N563) );
inv1 gate91( .a(N380), .O(N564) );
inv1 gate92( .a(N393), .O(N565) );
inv1 gate93( .a(N419), .O(N566) );
inv1 gate94( .a(N445), .O(N567) );
inv1 gate95( .a(N419), .O(N568) );
inv1 gate96( .a(N432), .O(N569) );
inv1 gate97( .a(N406), .O(N570) );
inv1 gate98( .a(N445), .O(N571) );
inv1 gate99( .a(N406), .O(N572) );
inv1 gate100( .a(N432), .O(N573) );
inv1 gate101( .a(N406), .O(N574) );
inv1 gate102( .a(N419), .O(N575) );
inv1 gate103( .a(N432), .O(N576) );
inv1 gate104( .a(N406), .O(N577) );
inv1 gate105( .a(N419), .O(N578) );
inv1 gate106( .a(N445), .O(N579) );
inv1 gate107( .a(N406), .O(N580) );
inv1 gate108( .a(N432), .O(N581) );
inv1 gate109( .a(N445), .O(N582) );
inv1 gate110( .a(N419), .O(N583) );
inv1 gate111( .a(N432), .O(N584) );
inv1 gate112( .a(N445), .O(N585) );
inv1 gate113( .a(N367), .O(N586) );
inv1 gate114( .a(N393), .O(N587) );
inv1 gate115( .a(N367), .O(N588) );
inv1 gate116( .a(N380), .O(N589) );
inv1 gate117( .a(N354), .O(N590) );
inv1 gate118( .a(N393), .O(N591) );
inv1 gate119( .a(N354), .O(N592) );
inv1 gate120( .a(N380), .O(N593) );
and4 gate121( .a(N554), .b(N555), .c(N556), .d(N393), .O(N594) );
and4 gate122( .a(N557), .b(N558), .c(N380), .d(N559), .O(N595) );
and4 gate123( .a(N560), .b(N367), .c(N561), .d(N562), .O(N596) );
and4 gate124( .a(N354), .b(N563), .c(N564), .d(N565), .O(N597) );
and4 gate125( .a(N574), .b(N575), .c(N576), .d(N445), .O(N598) );
and4 gate126( .a(N577), .b(N578), .c(N432), .d(N579), .O(N599) );
and4 gate127( .a(N580), .b(N419), .c(N581), .d(N582), .O(N600) );
and4 gate128( .a(N406), .b(N583), .c(N584), .d(N585), .O(N601) );
or4 gate129( .a(N594), .b(N595), .c(N596), .d(N597), .O(N602) );
or4 gate130( .a(N598), .b(N599), .c(N600), .d(N601), .O(N607) );
and5 gate131( .a(N406), .b(N566), .c(N432), .d(N567), .e(N602), .O(N620) );
and5 gate132( .a(N406), .b(N568), .c(N569), .d(N445), .e(N602), .O(N625) );
and5 gate133( .a(N570), .b(N419), .c(N432), .d(N571), .e(N602), .O(N630) );
and5 gate134( .a(N572), .b(N419), .c(N573), .d(N445), .e(N602), .O(N635) );
and5 gate135( .a(N354), .b(N586), .c(N380), .d(N587), .e(N607), .O(N640) );
and5 gate136( .a(N354), .b(N588), .c(N589), .d(N393), .e(N607), .O(N645) );
and5 gate137( .a(N590), .b(N367), .c(N380), .d(N591), .e(N607), .O(N650) );
and5 gate138( .a(N592), .b(N367), .c(N593), .d(N393), .e(N607), .O(N655) );
and2 gate139( .a(N354), .b(N620), .O(N692) );
and2 gate140( .a(N367), .b(N620), .O(N693) );
and2 gate141( .a(N380), .b(N620), .O(N694) );
and2 gate142( .a(N393), .b(N620), .O(N695) );
and2 gate143( .a(N354), .b(N625), .O(N696) );
and2 gate144( .a(N367), .b(N625), .O(N697) );
and2 gate145( .a(N380), .b(N625), .O(N698) );
and2 gate146( .a(N393), .b(N625), .O(N699) );
and2 gate147( .a(N354), .b(N630), .O(N700) );
and2 gate148( .a(N367), .b(N630), .O(N701) );
and2 gate149( .a(N380), .b(N630), .O(N702) );
and2 gate150( .a(N393), .b(N630), .O(N703) );
and2 gate151( .a(N354), .b(N635), .O(N704) );
and2 gate152( .a(N367), .b(N635), .O(N705) );
and2 gate153( .a(N380), .b(N635), .O(N706) );
and2 gate154( .a(N393), .b(N635), .O(N707) );
and2 gate155( .a(N406), .b(N640), .O(N708) );
and2 gate156( .a(N419), .b(N640), .O(N709) );
and2 gate157( .a(N432), .b(N640), .O(N710) );
and2 gate158( .a(N445), .b(N640), .O(N711) );
and2 gate159( .a(N406), .b(N645), .O(N712) );
and2 gate160( .a(N419), .b(N645), .O(N713) );
and2 gate161( .a(N432), .b(N645), .O(N714) );
and2 gate162( .a(N445), .b(N645), .O(N715) );
and2 gate163( .a(N406), .b(N650), .O(N716) );
and2 gate164( .a(N419), .b(N650), .O(N717) );
and2 gate165( .a(N432), .b(N650), .O(N718) );
and2 gate166( .a(N445), .b(N650), .O(N719) );
and2 gate167( .a(N406), .b(N655), .O(N720) );
and2 gate168( .a(N419), .b(N655), .O(N721) );
and2 gate169( .a(N432), .b(N655), .O(N722) );
and2 gate170( .a(N445), .b(N655), .O(N723) );

  xor2  gate469(.a(N692), .b(N1), .O(gate171inter0));
  nand2 gate470(.a(gate171inter0), .b(s_38), .O(gate171inter1));
  and2  gate471(.a(N692), .b(N1), .O(gate171inter2));
  inv1  gate472(.a(s_38), .O(gate171inter3));
  inv1  gate473(.a(s_39), .O(gate171inter4));
  nand2 gate474(.a(gate171inter4), .b(gate171inter3), .O(gate171inter5));
  nor2  gate475(.a(gate171inter5), .b(gate171inter2), .O(gate171inter6));
  inv1  gate476(.a(N1), .O(gate171inter7));
  inv1  gate477(.a(N692), .O(gate171inter8));
  nand2 gate478(.a(gate171inter8), .b(gate171inter7), .O(gate171inter9));
  nand2 gate479(.a(s_39), .b(gate171inter3), .O(gate171inter10));
  nor2  gate480(.a(gate171inter10), .b(gate171inter9), .O(gate171inter11));
  nor2  gate481(.a(gate171inter11), .b(gate171inter6), .O(gate171inter12));
  nand2 gate482(.a(gate171inter12), .b(gate171inter1), .O(N724));
xor2 gate172( .a(N5), .b(N693), .O(N725) );
xor2 gate173( .a(N9), .b(N694), .O(N726) );
xor2 gate174( .a(N13), .b(N695), .O(N727) );
xor2 gate175( .a(N17), .b(N696), .O(N728) );
xor2 gate176( .a(N21), .b(N697), .O(N729) );
xor2 gate177( .a(N25), .b(N698), .O(N730) );
xor2 gate178( .a(N29), .b(N699), .O(N731) );
xor2 gate179( .a(N33), .b(N700), .O(N732) );
xor2 gate180( .a(N37), .b(N701), .O(N733) );
xor2 gate181( .a(N41), .b(N702), .O(N734) );
xor2 gate182( .a(N45), .b(N703), .O(N735) );
xor2 gate183( .a(N49), .b(N704), .O(N736) );

  xor2  gate245(.a(N705), .b(N53), .O(gate184inter0));
  nand2 gate246(.a(gate184inter0), .b(s_6), .O(gate184inter1));
  and2  gate247(.a(N705), .b(N53), .O(gate184inter2));
  inv1  gate248(.a(s_6), .O(gate184inter3));
  inv1  gate249(.a(s_7), .O(gate184inter4));
  nand2 gate250(.a(gate184inter4), .b(gate184inter3), .O(gate184inter5));
  nor2  gate251(.a(gate184inter5), .b(gate184inter2), .O(gate184inter6));
  inv1  gate252(.a(N53), .O(gate184inter7));
  inv1  gate253(.a(N705), .O(gate184inter8));
  nand2 gate254(.a(gate184inter8), .b(gate184inter7), .O(gate184inter9));
  nand2 gate255(.a(s_7), .b(gate184inter3), .O(gate184inter10));
  nor2  gate256(.a(gate184inter10), .b(gate184inter9), .O(gate184inter11));
  nor2  gate257(.a(gate184inter11), .b(gate184inter6), .O(gate184inter12));
  nand2 gate258(.a(gate184inter12), .b(gate184inter1), .O(N737));
xor2 gate185( .a(N57), .b(N706), .O(N738) );
xor2 gate186( .a(N61), .b(N707), .O(N739) );
xor2 gate187( .a(N65), .b(N708), .O(N740) );

  xor2  gate231(.a(N709), .b(N69), .O(gate188inter0));
  nand2 gate232(.a(gate188inter0), .b(s_4), .O(gate188inter1));
  and2  gate233(.a(N709), .b(N69), .O(gate188inter2));
  inv1  gate234(.a(s_4), .O(gate188inter3));
  inv1  gate235(.a(s_5), .O(gate188inter4));
  nand2 gate236(.a(gate188inter4), .b(gate188inter3), .O(gate188inter5));
  nor2  gate237(.a(gate188inter5), .b(gate188inter2), .O(gate188inter6));
  inv1  gate238(.a(N69), .O(gate188inter7));
  inv1  gate239(.a(N709), .O(gate188inter8));
  nand2 gate240(.a(gate188inter8), .b(gate188inter7), .O(gate188inter9));
  nand2 gate241(.a(s_5), .b(gate188inter3), .O(gate188inter10));
  nor2  gate242(.a(gate188inter10), .b(gate188inter9), .O(gate188inter11));
  nor2  gate243(.a(gate188inter11), .b(gate188inter6), .O(gate188inter12));
  nand2 gate244(.a(gate188inter12), .b(gate188inter1), .O(N741));

  xor2  gate385(.a(N710), .b(N73), .O(gate189inter0));
  nand2 gate386(.a(gate189inter0), .b(s_26), .O(gate189inter1));
  and2  gate387(.a(N710), .b(N73), .O(gate189inter2));
  inv1  gate388(.a(s_26), .O(gate189inter3));
  inv1  gate389(.a(s_27), .O(gate189inter4));
  nand2 gate390(.a(gate189inter4), .b(gate189inter3), .O(gate189inter5));
  nor2  gate391(.a(gate189inter5), .b(gate189inter2), .O(gate189inter6));
  inv1  gate392(.a(N73), .O(gate189inter7));
  inv1  gate393(.a(N710), .O(gate189inter8));
  nand2 gate394(.a(gate189inter8), .b(gate189inter7), .O(gate189inter9));
  nand2 gate395(.a(s_27), .b(gate189inter3), .O(gate189inter10));
  nor2  gate396(.a(gate189inter10), .b(gate189inter9), .O(gate189inter11));
  nor2  gate397(.a(gate189inter11), .b(gate189inter6), .O(gate189inter12));
  nand2 gate398(.a(gate189inter12), .b(gate189inter1), .O(N742));
xor2 gate190( .a(N77), .b(N711), .O(N743) );
xor2 gate191( .a(N81), .b(N712), .O(N744) );

  xor2  gate427(.a(N713), .b(N85), .O(gate192inter0));
  nand2 gate428(.a(gate192inter0), .b(s_32), .O(gate192inter1));
  and2  gate429(.a(N713), .b(N85), .O(gate192inter2));
  inv1  gate430(.a(s_32), .O(gate192inter3));
  inv1  gate431(.a(s_33), .O(gate192inter4));
  nand2 gate432(.a(gate192inter4), .b(gate192inter3), .O(gate192inter5));
  nor2  gate433(.a(gate192inter5), .b(gate192inter2), .O(gate192inter6));
  inv1  gate434(.a(N85), .O(gate192inter7));
  inv1  gate435(.a(N713), .O(gate192inter8));
  nand2 gate436(.a(gate192inter8), .b(gate192inter7), .O(gate192inter9));
  nand2 gate437(.a(s_33), .b(gate192inter3), .O(gate192inter10));
  nor2  gate438(.a(gate192inter10), .b(gate192inter9), .O(gate192inter11));
  nor2  gate439(.a(gate192inter11), .b(gate192inter6), .O(gate192inter12));
  nand2 gate440(.a(gate192inter12), .b(gate192inter1), .O(N745));

  xor2  gate259(.a(N714), .b(N89), .O(gate193inter0));
  nand2 gate260(.a(gate193inter0), .b(s_8), .O(gate193inter1));
  and2  gate261(.a(N714), .b(N89), .O(gate193inter2));
  inv1  gate262(.a(s_8), .O(gate193inter3));
  inv1  gate263(.a(s_9), .O(gate193inter4));
  nand2 gate264(.a(gate193inter4), .b(gate193inter3), .O(gate193inter5));
  nor2  gate265(.a(gate193inter5), .b(gate193inter2), .O(gate193inter6));
  inv1  gate266(.a(N89), .O(gate193inter7));
  inv1  gate267(.a(N714), .O(gate193inter8));
  nand2 gate268(.a(gate193inter8), .b(gate193inter7), .O(gate193inter9));
  nand2 gate269(.a(s_9), .b(gate193inter3), .O(gate193inter10));
  nor2  gate270(.a(gate193inter10), .b(gate193inter9), .O(gate193inter11));
  nor2  gate271(.a(gate193inter11), .b(gate193inter6), .O(gate193inter12));
  nand2 gate272(.a(gate193inter12), .b(gate193inter1), .O(N746));
xor2 gate194( .a(N93), .b(N715), .O(N747) );
xor2 gate195( .a(N97), .b(N716), .O(N748) );
xor2 gate196( .a(N101), .b(N717), .O(N749) );

  xor2  gate343(.a(N718), .b(N105), .O(gate197inter0));
  nand2 gate344(.a(gate197inter0), .b(s_20), .O(gate197inter1));
  and2  gate345(.a(N718), .b(N105), .O(gate197inter2));
  inv1  gate346(.a(s_20), .O(gate197inter3));
  inv1  gate347(.a(s_21), .O(gate197inter4));
  nand2 gate348(.a(gate197inter4), .b(gate197inter3), .O(gate197inter5));
  nor2  gate349(.a(gate197inter5), .b(gate197inter2), .O(gate197inter6));
  inv1  gate350(.a(N105), .O(gate197inter7));
  inv1  gate351(.a(N718), .O(gate197inter8));
  nand2 gate352(.a(gate197inter8), .b(gate197inter7), .O(gate197inter9));
  nand2 gate353(.a(s_21), .b(gate197inter3), .O(gate197inter10));
  nor2  gate354(.a(gate197inter10), .b(gate197inter9), .O(gate197inter11));
  nor2  gate355(.a(gate197inter11), .b(gate197inter6), .O(gate197inter12));
  nand2 gate356(.a(gate197inter12), .b(gate197inter1), .O(N750));

  xor2  gate455(.a(N719), .b(N109), .O(gate198inter0));
  nand2 gate456(.a(gate198inter0), .b(s_36), .O(gate198inter1));
  and2  gate457(.a(N719), .b(N109), .O(gate198inter2));
  inv1  gate458(.a(s_36), .O(gate198inter3));
  inv1  gate459(.a(s_37), .O(gate198inter4));
  nand2 gate460(.a(gate198inter4), .b(gate198inter3), .O(gate198inter5));
  nor2  gate461(.a(gate198inter5), .b(gate198inter2), .O(gate198inter6));
  inv1  gate462(.a(N109), .O(gate198inter7));
  inv1  gate463(.a(N719), .O(gate198inter8));
  nand2 gate464(.a(gate198inter8), .b(gate198inter7), .O(gate198inter9));
  nand2 gate465(.a(s_37), .b(gate198inter3), .O(gate198inter10));
  nor2  gate466(.a(gate198inter10), .b(gate198inter9), .O(gate198inter11));
  nor2  gate467(.a(gate198inter11), .b(gate198inter6), .O(gate198inter12));
  nand2 gate468(.a(gate198inter12), .b(gate198inter1), .O(N751));
xor2 gate199( .a(N113), .b(N720), .O(N752) );
xor2 gate200( .a(N117), .b(N721), .O(N753) );
xor2 gate201( .a(N121), .b(N722), .O(N754) );
xor2 gate202( .a(N125), .b(N723), .O(N755) );

endmodule