module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);

input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;//RE__PI;

input s_0,s_1;//RE__ALLOW(00,01,10,11);
input s_2,s_3;//RE__ALLOW(00,01,10,11);
input s_4,s_5;//RE__ALLOW(00,01,10,11);
input s_6,s_7;//RE__ALLOW(00,01,10,11);
input s_8,s_9;//RE__ALLOW(00,01,10,11);
input s_10,s_11;//RE__ALLOW(00,01,10,11);
input s_12,s_13;//RE__ALLOW(00,01,10,11);
input s_14,s_15;//RE__ALLOW(00,01,10,11);
input s_16,s_17;//RE__ALLOW(00,01,10,11);
input s_18,s_19;//RE__ALLOW(00,01,10,11);
input s_20,s_21;//RE__ALLOW(00,01,10,11);
input s_22,s_23;//RE__ALLOW(00,01,10,11);
input s_24,s_25;//RE__ALLOW(00,01,10,11);
input s_26,s_27;//RE__ALLOW(00,01,10,11);
input s_28,s_29;//RE__ALLOW(00,01,10,11);
input s_30,s_31;//RE__ALLOW(00,01,10,11);
input s_32,s_33;//RE__ALLOW(00,01,10,11);
input s_34,s_35;//RE__ALLOW(00,01,10,11);
input s_36,s_37;//RE__ALLOW(00,01,10,11);
input s_38,s_39;//RE__ALLOW(00,01,10,11);
input s_40,s_41;//RE__ALLOW(00,01,10,11);
input s_42,s_43;//RE__ALLOW(00,01,10,11);
input s_44,s_45;//RE__ALLOW(00,01,10,11);
input s_46,s_47;//RE__ALLOW(00,01,10,11);
input s_48,s_49;//RE__ALLOW(00,01,10,11);
input s_50,s_51;//RE__ALLOW(00,01,10,11);
input s_52,s_53;//RE__ALLOW(00,01,10,11);
input s_54,s_55;//RE__ALLOW(00,01,10,11);
input s_56,s_57;//RE__ALLOW(00,01,10,11);
input s_58,s_59;//RE__ALLOW(00,01,10,11);
input s_60,s_61;//RE__ALLOW(00,01,10,11);
input s_62,s_63;//RE__ALLOW(00,01,10,11);
input s_64,s_65;//RE__ALLOW(00,01,10,11);
input s_66,s_67;//RE__ALLOW(00,01,10,11);
input s_68,s_69;//RE__ALLOW(00,01,10,11);
input s_70,s_71;//RE__ALLOW(00,01,10,11);
input s_72,s_73;//RE__ALLOW(00,01,10,11);
input s_74,s_75;//RE__ALLOW(00,01,10,11);
input s_76,s_77;//RE__ALLOW(00,01,10,11);
input s_78,s_79;//RE__ALLOW(00,01,10,11);
input s_80,s_81;//RE__ALLOW(00,01,10,11);
input s_82,s_83;//RE__ALLOW(00,01,10,11);
input s_84,s_85;//RE__ALLOW(00,01,10,11);
input s_86,s_87;//RE__ALLOW(00,01,10,11);
input s_88,s_89;//RE__ALLOW(00,01,10,11);
input s_90,s_91;//RE__ALLOW(00,01,10,11);
input s_92,s_93;//RE__ALLOW(00,01,10,11);
input s_94,s_95;//RE__ALLOW(00,01,10,11);
input s_96,s_97;//RE__ALLOW(00,01,10,11);
input s_98,s_99;//RE__ALLOW(00,01,10,11);
input s_100,s_101;//RE__ALLOW(00,01,10,11);
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;

  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate19inter0, gate19inter1, gate19inter2, gate19inter3, gate19inter4, gate19inter5, gate19inter6, gate19inter7, gate19inter8, gate19inter9, gate19inter10, gate19inter11, gate19inter12, gate431inter0, gate431inter1, gate431inter2, gate431inter3, gate431inter4, gate431inter5, gate431inter6, gate431inter7, gate431inter8, gate431inter9, gate431inter10, gate431inter11, gate431inter12, gate130inter0, gate130inter1, gate130inter2, gate130inter3, gate130inter4, gate130inter5, gate130inter6, gate130inter7, gate130inter8, gate130inter9, gate130inter10, gate130inter11, gate130inter12, gate218inter0, gate218inter1, gate218inter2, gate218inter3, gate218inter4, gate218inter5, gate218inter6, gate218inter7, gate218inter8, gate218inter9, gate218inter10, gate218inter11, gate218inter12, gate281inter0, gate281inter1, gate281inter2, gate281inter3, gate281inter4, gate281inter5, gate281inter6, gate281inter7, gate281inter8, gate281inter9, gate281inter10, gate281inter11, gate281inter12, gate89inter0, gate89inter1, gate89inter2, gate89inter3, gate89inter4, gate89inter5, gate89inter6, gate89inter7, gate89inter8, gate89inter9, gate89inter10, gate89inter11, gate89inter12, gate68inter0, gate68inter1, gate68inter2, gate68inter3, gate68inter4, gate68inter5, gate68inter6, gate68inter7, gate68inter8, gate68inter9, gate68inter10, gate68inter11, gate68inter12, gate396inter0, gate396inter1, gate396inter2, gate396inter3, gate396inter4, gate396inter5, gate396inter6, gate396inter7, gate396inter8, gate396inter9, gate396inter10, gate396inter11, gate396inter12, gate388inter0, gate388inter1, gate388inter2, gate388inter3, gate388inter4, gate388inter5, gate388inter6, gate388inter7, gate388inter8, gate388inter9, gate388inter10, gate388inter11, gate388inter12, gate453inter0, gate453inter1, gate453inter2, gate453inter3, gate453inter4, gate453inter5, gate453inter6, gate453inter7, gate453inter8, gate453inter9, gate453inter10, gate453inter11, gate453inter12, gate462inter0, gate462inter1, gate462inter2, gate462inter3, gate462inter4, gate462inter5, gate462inter6, gate462inter7, gate462inter8, gate462inter9, gate462inter10, gate462inter11, gate462inter12, gate454inter0, gate454inter1, gate454inter2, gate454inter3, gate454inter4, gate454inter5, gate454inter6, gate454inter7, gate454inter8, gate454inter9, gate454inter10, gate454inter11, gate454inter12, gate164inter0, gate164inter1, gate164inter2, gate164inter3, gate164inter4, gate164inter5, gate164inter6, gate164inter7, gate164inter8, gate164inter9, gate164inter10, gate164inter11, gate164inter12, gate10inter0, gate10inter1, gate10inter2, gate10inter3, gate10inter4, gate10inter5, gate10inter6, gate10inter7, gate10inter8, gate10inter9, gate10inter10, gate10inter11, gate10inter12, gate272inter0, gate272inter1, gate272inter2, gate272inter3, gate272inter4, gate272inter5, gate272inter6, gate272inter7, gate272inter8, gate272inter9, gate272inter10, gate272inter11, gate272inter12, gate223inter0, gate223inter1, gate223inter2, gate223inter3, gate223inter4, gate223inter5, gate223inter6, gate223inter7, gate223inter8, gate223inter9, gate223inter10, gate223inter11, gate223inter12, gate479inter0, gate479inter1, gate479inter2, gate479inter3, gate479inter4, gate479inter5, gate479inter6, gate479inter7, gate479inter8, gate479inter9, gate479inter10, gate479inter11, gate479inter12, gate291inter0, gate291inter1, gate291inter2, gate291inter3, gate291inter4, gate291inter5, gate291inter6, gate291inter7, gate291inter8, gate291inter9, gate291inter10, gate291inter11, gate291inter12, gate390inter0, gate390inter1, gate390inter2, gate390inter3, gate390inter4, gate390inter5, gate390inter6, gate390inter7, gate390inter8, gate390inter9, gate390inter10, gate390inter11, gate390inter12, gate501inter0, gate501inter1, gate501inter2, gate501inter3, gate501inter4, gate501inter5, gate501inter6, gate501inter7, gate501inter8, gate501inter9, gate501inter10, gate501inter11, gate501inter12, gate439inter0, gate439inter1, gate439inter2, gate439inter3, gate439inter4, gate439inter5, gate439inter6, gate439inter7, gate439inter8, gate439inter9, gate439inter10, gate439inter11, gate439inter12, gate77inter0, gate77inter1, gate77inter2, gate77inter3, gate77inter4, gate77inter5, gate77inter6, gate77inter7, gate77inter8, gate77inter9, gate77inter10, gate77inter11, gate77inter12, gate103inter0, gate103inter1, gate103inter2, gate103inter3, gate103inter4, gate103inter5, gate103inter6, gate103inter7, gate103inter8, gate103inter9, gate103inter10, gate103inter11, gate103inter12, gate94inter0, gate94inter1, gate94inter2, gate94inter3, gate94inter4, gate94inter5, gate94inter6, gate94inter7, gate94inter8, gate94inter9, gate94inter10, gate94inter11, gate94inter12, gate25inter0, gate25inter1, gate25inter2, gate25inter3, gate25inter4, gate25inter5, gate25inter6, gate25inter7, gate25inter8, gate25inter9, gate25inter10, gate25inter11, gate25inter12, gate170inter0, gate170inter1, gate170inter2, gate170inter3, gate170inter4, gate170inter5, gate170inter6, gate170inter7, gate170inter8, gate170inter9, gate170inter10, gate170inter11, gate170inter12, gate243inter0, gate243inter1, gate243inter2, gate243inter3, gate243inter4, gate243inter5, gate243inter6, gate243inter7, gate243inter8, gate243inter9, gate243inter10, gate243inter11, gate243inter12, gate163inter0, gate163inter1, gate163inter2, gate163inter3, gate163inter4, gate163inter5, gate163inter6, gate163inter7, gate163inter8, gate163inter9, gate163inter10, gate163inter11, gate163inter12, gate75inter0, gate75inter1, gate75inter2, gate75inter3, gate75inter4, gate75inter5, gate75inter6, gate75inter7, gate75inter8, gate75inter9, gate75inter10, gate75inter11, gate75inter12, gate246inter0, gate246inter1, gate246inter2, gate246inter3, gate246inter4, gate246inter5, gate246inter6, gate246inter7, gate246inter8, gate246inter9, gate246inter10, gate246inter11, gate246inter12, gate438inter0, gate438inter1, gate438inter2, gate438inter3, gate438inter4, gate438inter5, gate438inter6, gate438inter7, gate438inter8, gate438inter9, gate438inter10, gate438inter11, gate438inter12, gate514inter0, gate514inter1, gate514inter2, gate514inter3, gate514inter4, gate514inter5, gate514inter6, gate514inter7, gate514inter8, gate514inter9, gate514inter10, gate514inter11, gate514inter12, gate98inter0, gate98inter1, gate98inter2, gate98inter3, gate98inter4, gate98inter5, gate98inter6, gate98inter7, gate98inter8, gate98inter9, gate98inter10, gate98inter11, gate98inter12, gate265inter0, gate265inter1, gate265inter2, gate265inter3, gate265inter4, gate265inter5, gate265inter6, gate265inter7, gate265inter8, gate265inter9, gate265inter10, gate265inter11, gate265inter12, gate220inter0, gate220inter1, gate220inter2, gate220inter3, gate220inter4, gate220inter5, gate220inter6, gate220inter7, gate220inter8, gate220inter9, gate220inter10, gate220inter11, gate220inter12, gate175inter0, gate175inter1, gate175inter2, gate175inter3, gate175inter4, gate175inter5, gate175inter6, gate175inter7, gate175inter8, gate175inter9, gate175inter10, gate175inter11, gate175inter12, gate102inter0, gate102inter1, gate102inter2, gate102inter3, gate102inter4, gate102inter5, gate102inter6, gate102inter7, gate102inter8, gate102inter9, gate102inter10, gate102inter11, gate102inter12, gate231inter0, gate231inter1, gate231inter2, gate231inter3, gate231inter4, gate231inter5, gate231inter6, gate231inter7, gate231inter8, gate231inter9, gate231inter10, gate231inter11, gate231inter12, gate510inter0, gate510inter1, gate510inter2, gate510inter3, gate510inter4, gate510inter5, gate510inter6, gate510inter7, gate510inter8, gate510inter9, gate510inter10, gate510inter11, gate510inter12, gate470inter0, gate470inter1, gate470inter2, gate470inter3, gate470inter4, gate470inter5, gate470inter6, gate470inter7, gate470inter8, gate470inter9, gate470inter10, gate470inter11, gate470inter12, gate179inter0, gate179inter1, gate179inter2, gate179inter3, gate179inter4, gate179inter5, gate179inter6, gate179inter7, gate179inter8, gate179inter9, gate179inter10, gate179inter11, gate179inter12, gate495inter0, gate495inter1, gate495inter2, gate495inter3, gate495inter4, gate495inter5, gate495inter6, gate495inter7, gate495inter8, gate495inter9, gate495inter10, gate495inter11, gate495inter12, gate508inter0, gate508inter1, gate508inter2, gate508inter3, gate508inter4, gate508inter5, gate508inter6, gate508inter7, gate508inter8, gate508inter9, gate508inter10, gate508inter11, gate508inter12, gate232inter0, gate232inter1, gate232inter2, gate232inter3, gate232inter4, gate232inter5, gate232inter6, gate232inter7, gate232inter8, gate232inter9, gate232inter10, gate232inter11, gate232inter12, gate200inter0, gate200inter1, gate200inter2, gate200inter3, gate200inter4, gate200inter5, gate200inter6, gate200inter7, gate200inter8, gate200inter9, gate200inter10, gate200inter11, gate200inter12, gate234inter0, gate234inter1, gate234inter2, gate234inter3, gate234inter4, gate234inter5, gate234inter6, gate234inter7, gate234inter8, gate234inter9, gate234inter10, gate234inter11, gate234inter12, gate140inter0, gate140inter1, gate140inter2, gate140inter3, gate140inter4, gate140inter5, gate140inter6, gate140inter7, gate140inter8, gate140inter9, gate140inter10, gate140inter11, gate140inter12, gate209inter0, gate209inter1, gate209inter2, gate209inter3, gate209inter4, gate209inter5, gate209inter6, gate209inter7, gate209inter8, gate209inter9, gate209inter10, gate209inter11, gate209inter12, gate441inter0, gate441inter1, gate441inter2, gate441inter3, gate441inter4, gate441inter5, gate441inter6, gate441inter7, gate441inter8, gate441inter9, gate441inter10, gate441inter11, gate441inter12, gate187inter0, gate187inter1, gate187inter2, gate187inter3, gate187inter4, gate187inter5, gate187inter6, gate187inter7, gate187inter8, gate187inter9, gate187inter10, gate187inter11, gate187inter12, gate256inter0, gate256inter1, gate256inter2, gate256inter3, gate256inter4, gate256inter5, gate256inter6, gate256inter7, gate256inter8, gate256inter9, gate256inter10, gate256inter11, gate256inter12;



and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );
nand2 gate9( .a(G1), .b(G2), .O(G266) );

  xor2  gate729(.a(G4), .b(G3), .O(gate10inter0));
  nand2 gate730(.a(gate10inter0), .b(s_26), .O(gate10inter1));
  and2  gate731(.a(G4), .b(G3), .O(gate10inter2));
  inv1  gate732(.a(s_26), .O(gate10inter3));
  inv1  gate733(.a(s_27), .O(gate10inter4));
  nand2 gate734(.a(gate10inter4), .b(gate10inter3), .O(gate10inter5));
  nor2  gate735(.a(gate10inter5), .b(gate10inter2), .O(gate10inter6));
  inv1  gate736(.a(G3), .O(gate10inter7));
  inv1  gate737(.a(G4), .O(gate10inter8));
  nand2 gate738(.a(gate10inter8), .b(gate10inter7), .O(gate10inter9));
  nand2 gate739(.a(s_27), .b(gate10inter3), .O(gate10inter10));
  nor2  gate740(.a(gate10inter10), .b(gate10inter9), .O(gate10inter11));
  nor2  gate741(.a(gate10inter11), .b(gate10inter6), .O(gate10inter12));
  nand2 gate742(.a(gate10inter12), .b(gate10inter1), .O(G269));
nand2 gate11( .a(G5), .b(G6), .O(G272) );
nand2 gate12( .a(G7), .b(G8), .O(G275) );
nand2 gate13( .a(G9), .b(G10), .O(G278) );
nand2 gate14( .a(G11), .b(G12), .O(G281) );
nand2 gate15( .a(G13), .b(G14), .O(G284) );
nand2 gate16( .a(G15), .b(G16), .O(G287) );
nand2 gate17( .a(G17), .b(G18), .O(G290) );
nand2 gate18( .a(G19), .b(G20), .O(G293) );

  xor2  gate547(.a(G22), .b(G21), .O(gate19inter0));
  nand2 gate548(.a(gate19inter0), .b(s_0), .O(gate19inter1));
  and2  gate549(.a(G22), .b(G21), .O(gate19inter2));
  inv1  gate550(.a(s_0), .O(gate19inter3));
  inv1  gate551(.a(s_1), .O(gate19inter4));
  nand2 gate552(.a(gate19inter4), .b(gate19inter3), .O(gate19inter5));
  nor2  gate553(.a(gate19inter5), .b(gate19inter2), .O(gate19inter6));
  inv1  gate554(.a(G21), .O(gate19inter7));
  inv1  gate555(.a(G22), .O(gate19inter8));
  nand2 gate556(.a(gate19inter8), .b(gate19inter7), .O(gate19inter9));
  nand2 gate557(.a(s_1), .b(gate19inter3), .O(gate19inter10));
  nor2  gate558(.a(gate19inter10), .b(gate19inter9), .O(gate19inter11));
  nor2  gate559(.a(gate19inter11), .b(gate19inter6), .O(gate19inter12));
  nand2 gate560(.a(gate19inter12), .b(gate19inter1), .O(G296));
nand2 gate20( .a(G23), .b(G24), .O(G299) );
nand2 gate21( .a(G25), .b(G26), .O(G302) );
nand2 gate22( .a(G27), .b(G28), .O(G305) );
nand2 gate23( .a(G29), .b(G30), .O(G308) );
nand2 gate24( .a(G31), .b(G32), .O(G311) );

  xor2  gate883(.a(G5), .b(G1), .O(gate25inter0));
  nand2 gate884(.a(gate25inter0), .b(s_48), .O(gate25inter1));
  and2  gate885(.a(G5), .b(G1), .O(gate25inter2));
  inv1  gate886(.a(s_48), .O(gate25inter3));
  inv1  gate887(.a(s_49), .O(gate25inter4));
  nand2 gate888(.a(gate25inter4), .b(gate25inter3), .O(gate25inter5));
  nor2  gate889(.a(gate25inter5), .b(gate25inter2), .O(gate25inter6));
  inv1  gate890(.a(G1), .O(gate25inter7));
  inv1  gate891(.a(G5), .O(gate25inter8));
  nand2 gate892(.a(gate25inter8), .b(gate25inter7), .O(gate25inter9));
  nand2 gate893(.a(s_49), .b(gate25inter3), .O(gate25inter10));
  nor2  gate894(.a(gate25inter10), .b(gate25inter9), .O(gate25inter11));
  nor2  gate895(.a(gate25inter11), .b(gate25inter6), .O(gate25inter12));
  nand2 gate896(.a(gate25inter12), .b(gate25inter1), .O(G314));
nand2 gate26( .a(G9), .b(G13), .O(G317) );
nand2 gate27( .a(G2), .b(G6), .O(G320) );
nand2 gate28( .a(G10), .b(G14), .O(G323) );
nand2 gate29( .a(G3), .b(G7), .O(G326) );
nand2 gate30( .a(G11), .b(G15), .O(G329) );
nand2 gate31( .a(G4), .b(G8), .O(G332) );
nand2 gate32( .a(G12), .b(G16), .O(G335) );
nand2 gate33( .a(G17), .b(G21), .O(G338) );
nand2 gate34( .a(G25), .b(G29), .O(G341) );
nand2 gate35( .a(G18), .b(G22), .O(G344) );
nand2 gate36( .a(G26), .b(G30), .O(G347) );
nand2 gate37( .a(G19), .b(G23), .O(G350) );
nand2 gate38( .a(G27), .b(G31), .O(G353) );
nand2 gate39( .a(G20), .b(G24), .O(G356) );
nand2 gate40( .a(G28), .b(G32), .O(G359) );
nand2 gate41( .a(G1), .b(G266), .O(G362) );
nand2 gate42( .a(G2), .b(G266), .O(G363) );
nand2 gate43( .a(G3), .b(G269), .O(G364) );
nand2 gate44( .a(G4), .b(G269), .O(G365) );
nand2 gate45( .a(G5), .b(G272), .O(G366) );
nand2 gate46( .a(G6), .b(G272), .O(G367) );
nand2 gate47( .a(G7), .b(G275), .O(G368) );
nand2 gate48( .a(G8), .b(G275), .O(G369) );
nand2 gate49( .a(G9), .b(G278), .O(G370) );
nand2 gate50( .a(G10), .b(G278), .O(G371) );
nand2 gate51( .a(G11), .b(G281), .O(G372) );
nand2 gate52( .a(G12), .b(G281), .O(G373) );
nand2 gate53( .a(G13), .b(G284), .O(G374) );
nand2 gate54( .a(G14), .b(G284), .O(G375) );
nand2 gate55( .a(G15), .b(G287), .O(G376) );
nand2 gate56( .a(G16), .b(G287), .O(G377) );
nand2 gate57( .a(G17), .b(G290), .O(G378) );
nand2 gate58( .a(G18), .b(G290), .O(G379) );
nand2 gate59( .a(G19), .b(G293), .O(G380) );
nand2 gate60( .a(G20), .b(G293), .O(G381) );
nand2 gate61( .a(G21), .b(G296), .O(G382) );
nand2 gate62( .a(G22), .b(G296), .O(G383) );
nand2 gate63( .a(G23), .b(G299), .O(G384) );
nand2 gate64( .a(G24), .b(G299), .O(G385) );
nand2 gate65( .a(G25), .b(G302), .O(G386) );
nand2 gate66( .a(G26), .b(G302), .O(G387) );
nand2 gate67( .a(G27), .b(G305), .O(G388) );

  xor2  gate631(.a(G305), .b(G28), .O(gate68inter0));
  nand2 gate632(.a(gate68inter0), .b(s_12), .O(gate68inter1));
  and2  gate633(.a(G305), .b(G28), .O(gate68inter2));
  inv1  gate634(.a(s_12), .O(gate68inter3));
  inv1  gate635(.a(s_13), .O(gate68inter4));
  nand2 gate636(.a(gate68inter4), .b(gate68inter3), .O(gate68inter5));
  nor2  gate637(.a(gate68inter5), .b(gate68inter2), .O(gate68inter6));
  inv1  gate638(.a(G28), .O(gate68inter7));
  inv1  gate639(.a(G305), .O(gate68inter8));
  nand2 gate640(.a(gate68inter8), .b(gate68inter7), .O(gate68inter9));
  nand2 gate641(.a(s_13), .b(gate68inter3), .O(gate68inter10));
  nor2  gate642(.a(gate68inter10), .b(gate68inter9), .O(gate68inter11));
  nor2  gate643(.a(gate68inter11), .b(gate68inter6), .O(gate68inter12));
  nand2 gate644(.a(gate68inter12), .b(gate68inter1), .O(G389));
nand2 gate69( .a(G29), .b(G308), .O(G390) );
nand2 gate70( .a(G30), .b(G308), .O(G391) );
nand2 gate71( .a(G31), .b(G311), .O(G392) );
nand2 gate72( .a(G32), .b(G311), .O(G393) );
nand2 gate73( .a(G1), .b(G314), .O(G394) );
nand2 gate74( .a(G5), .b(G314), .O(G395) );

  xor2  gate939(.a(G317), .b(G9), .O(gate75inter0));
  nand2 gate940(.a(gate75inter0), .b(s_56), .O(gate75inter1));
  and2  gate941(.a(G317), .b(G9), .O(gate75inter2));
  inv1  gate942(.a(s_56), .O(gate75inter3));
  inv1  gate943(.a(s_57), .O(gate75inter4));
  nand2 gate944(.a(gate75inter4), .b(gate75inter3), .O(gate75inter5));
  nor2  gate945(.a(gate75inter5), .b(gate75inter2), .O(gate75inter6));
  inv1  gate946(.a(G9), .O(gate75inter7));
  inv1  gate947(.a(G317), .O(gate75inter8));
  nand2 gate948(.a(gate75inter8), .b(gate75inter7), .O(gate75inter9));
  nand2 gate949(.a(s_57), .b(gate75inter3), .O(gate75inter10));
  nor2  gate950(.a(gate75inter10), .b(gate75inter9), .O(gate75inter11));
  nor2  gate951(.a(gate75inter11), .b(gate75inter6), .O(gate75inter12));
  nand2 gate952(.a(gate75inter12), .b(gate75inter1), .O(G396));
nand2 gate76( .a(G13), .b(G317), .O(G397) );

  xor2  gate841(.a(G320), .b(G2), .O(gate77inter0));
  nand2 gate842(.a(gate77inter0), .b(s_42), .O(gate77inter1));
  and2  gate843(.a(G320), .b(G2), .O(gate77inter2));
  inv1  gate844(.a(s_42), .O(gate77inter3));
  inv1  gate845(.a(s_43), .O(gate77inter4));
  nand2 gate846(.a(gate77inter4), .b(gate77inter3), .O(gate77inter5));
  nor2  gate847(.a(gate77inter5), .b(gate77inter2), .O(gate77inter6));
  inv1  gate848(.a(G2), .O(gate77inter7));
  inv1  gate849(.a(G320), .O(gate77inter8));
  nand2 gate850(.a(gate77inter8), .b(gate77inter7), .O(gate77inter9));
  nand2 gate851(.a(s_43), .b(gate77inter3), .O(gate77inter10));
  nor2  gate852(.a(gate77inter10), .b(gate77inter9), .O(gate77inter11));
  nor2  gate853(.a(gate77inter11), .b(gate77inter6), .O(gate77inter12));
  nand2 gate854(.a(gate77inter12), .b(gate77inter1), .O(G398));
nand2 gate78( .a(G6), .b(G320), .O(G399) );
nand2 gate79( .a(G10), .b(G323), .O(G400) );
nand2 gate80( .a(G14), .b(G323), .O(G401) );
nand2 gate81( .a(G3), .b(G326), .O(G402) );
nand2 gate82( .a(G7), .b(G326), .O(G403) );
nand2 gate83( .a(G11), .b(G329), .O(G404) );
nand2 gate84( .a(G15), .b(G329), .O(G405) );
nand2 gate85( .a(G4), .b(G332), .O(G406) );
nand2 gate86( .a(G8), .b(G332), .O(G407) );
nand2 gate87( .a(G12), .b(G335), .O(G408) );
nand2 gate88( .a(G16), .b(G335), .O(G409) );

  xor2  gate617(.a(G338), .b(G17), .O(gate89inter0));
  nand2 gate618(.a(gate89inter0), .b(s_10), .O(gate89inter1));
  and2  gate619(.a(G338), .b(G17), .O(gate89inter2));
  inv1  gate620(.a(s_10), .O(gate89inter3));
  inv1  gate621(.a(s_11), .O(gate89inter4));
  nand2 gate622(.a(gate89inter4), .b(gate89inter3), .O(gate89inter5));
  nor2  gate623(.a(gate89inter5), .b(gate89inter2), .O(gate89inter6));
  inv1  gate624(.a(G17), .O(gate89inter7));
  inv1  gate625(.a(G338), .O(gate89inter8));
  nand2 gate626(.a(gate89inter8), .b(gate89inter7), .O(gate89inter9));
  nand2 gate627(.a(s_11), .b(gate89inter3), .O(gate89inter10));
  nor2  gate628(.a(gate89inter10), .b(gate89inter9), .O(gate89inter11));
  nor2  gate629(.a(gate89inter11), .b(gate89inter6), .O(gate89inter12));
  nand2 gate630(.a(gate89inter12), .b(gate89inter1), .O(G410));
nand2 gate90( .a(G21), .b(G338), .O(G411) );
nand2 gate91( .a(G25), .b(G341), .O(G412) );
nand2 gate92( .a(G29), .b(G341), .O(G413) );
nand2 gate93( .a(G18), .b(G344), .O(G414) );

  xor2  gate869(.a(G344), .b(G22), .O(gate94inter0));
  nand2 gate870(.a(gate94inter0), .b(s_46), .O(gate94inter1));
  and2  gate871(.a(G344), .b(G22), .O(gate94inter2));
  inv1  gate872(.a(s_46), .O(gate94inter3));
  inv1  gate873(.a(s_47), .O(gate94inter4));
  nand2 gate874(.a(gate94inter4), .b(gate94inter3), .O(gate94inter5));
  nor2  gate875(.a(gate94inter5), .b(gate94inter2), .O(gate94inter6));
  inv1  gate876(.a(G22), .O(gate94inter7));
  inv1  gate877(.a(G344), .O(gate94inter8));
  nand2 gate878(.a(gate94inter8), .b(gate94inter7), .O(gate94inter9));
  nand2 gate879(.a(s_47), .b(gate94inter3), .O(gate94inter10));
  nor2  gate880(.a(gate94inter10), .b(gate94inter9), .O(gate94inter11));
  nor2  gate881(.a(gate94inter11), .b(gate94inter6), .O(gate94inter12));
  nand2 gate882(.a(gate94inter12), .b(gate94inter1), .O(G415));
nand2 gate95( .a(G26), .b(G347), .O(G416) );
nand2 gate96( .a(G30), .b(G347), .O(G417) );
nand2 gate97( .a(G19), .b(G350), .O(G418) );

  xor2  gate995(.a(G350), .b(G23), .O(gate98inter0));
  nand2 gate996(.a(gate98inter0), .b(s_64), .O(gate98inter1));
  and2  gate997(.a(G350), .b(G23), .O(gate98inter2));
  inv1  gate998(.a(s_64), .O(gate98inter3));
  inv1  gate999(.a(s_65), .O(gate98inter4));
  nand2 gate1000(.a(gate98inter4), .b(gate98inter3), .O(gate98inter5));
  nor2  gate1001(.a(gate98inter5), .b(gate98inter2), .O(gate98inter6));
  inv1  gate1002(.a(G23), .O(gate98inter7));
  inv1  gate1003(.a(G350), .O(gate98inter8));
  nand2 gate1004(.a(gate98inter8), .b(gate98inter7), .O(gate98inter9));
  nand2 gate1005(.a(s_65), .b(gate98inter3), .O(gate98inter10));
  nor2  gate1006(.a(gate98inter10), .b(gate98inter9), .O(gate98inter11));
  nor2  gate1007(.a(gate98inter11), .b(gate98inter6), .O(gate98inter12));
  nand2 gate1008(.a(gate98inter12), .b(gate98inter1), .O(G419));
nand2 gate99( .a(G27), .b(G353), .O(G420) );
nand2 gate100( .a(G31), .b(G353), .O(G421) );
nand2 gate101( .a(G20), .b(G356), .O(G422) );

  xor2  gate1051(.a(G356), .b(G24), .O(gate102inter0));
  nand2 gate1052(.a(gate102inter0), .b(s_72), .O(gate102inter1));
  and2  gate1053(.a(G356), .b(G24), .O(gate102inter2));
  inv1  gate1054(.a(s_72), .O(gate102inter3));
  inv1  gate1055(.a(s_73), .O(gate102inter4));
  nand2 gate1056(.a(gate102inter4), .b(gate102inter3), .O(gate102inter5));
  nor2  gate1057(.a(gate102inter5), .b(gate102inter2), .O(gate102inter6));
  inv1  gate1058(.a(G24), .O(gate102inter7));
  inv1  gate1059(.a(G356), .O(gate102inter8));
  nand2 gate1060(.a(gate102inter8), .b(gate102inter7), .O(gate102inter9));
  nand2 gate1061(.a(s_73), .b(gate102inter3), .O(gate102inter10));
  nor2  gate1062(.a(gate102inter10), .b(gate102inter9), .O(gate102inter11));
  nor2  gate1063(.a(gate102inter11), .b(gate102inter6), .O(gate102inter12));
  nand2 gate1064(.a(gate102inter12), .b(gate102inter1), .O(G423));

  xor2  gate855(.a(G359), .b(G28), .O(gate103inter0));
  nand2 gate856(.a(gate103inter0), .b(s_44), .O(gate103inter1));
  and2  gate857(.a(G359), .b(G28), .O(gate103inter2));
  inv1  gate858(.a(s_44), .O(gate103inter3));
  inv1  gate859(.a(s_45), .O(gate103inter4));
  nand2 gate860(.a(gate103inter4), .b(gate103inter3), .O(gate103inter5));
  nor2  gate861(.a(gate103inter5), .b(gate103inter2), .O(gate103inter6));
  inv1  gate862(.a(G28), .O(gate103inter7));
  inv1  gate863(.a(G359), .O(gate103inter8));
  nand2 gate864(.a(gate103inter8), .b(gate103inter7), .O(gate103inter9));
  nand2 gate865(.a(s_45), .b(gate103inter3), .O(gate103inter10));
  nor2  gate866(.a(gate103inter10), .b(gate103inter9), .O(gate103inter11));
  nor2  gate867(.a(gate103inter11), .b(gate103inter6), .O(gate103inter12));
  nand2 gate868(.a(gate103inter12), .b(gate103inter1), .O(G424));
nand2 gate104( .a(G32), .b(G359), .O(G425) );
nand2 gate105( .a(G362), .b(G363), .O(G426) );
nand2 gate106( .a(G364), .b(G365), .O(G429) );
nand2 gate107( .a(G366), .b(G367), .O(G432) );
nand2 gate108( .a(G368), .b(G369), .O(G435) );
nand2 gate109( .a(G370), .b(G371), .O(G438) );
nand2 gate110( .a(G372), .b(G373), .O(G441) );
nand2 gate111( .a(G374), .b(G375), .O(G444) );
nand2 gate112( .a(G376), .b(G377), .O(G447) );
nand2 gate113( .a(G378), .b(G379), .O(G450) );
nand2 gate114( .a(G380), .b(G381), .O(G453) );
nand2 gate115( .a(G382), .b(G383), .O(G456) );
nand2 gate116( .a(G384), .b(G385), .O(G459) );
nand2 gate117( .a(G386), .b(G387), .O(G462) );
nand2 gate118( .a(G388), .b(G389), .O(G465) );
nand2 gate119( .a(G390), .b(G391), .O(G468) );
nand2 gate120( .a(G392), .b(G393), .O(G471) );
nand2 gate121( .a(G394), .b(G395), .O(G474) );
nand2 gate122( .a(G396), .b(G397), .O(G477) );
nand2 gate123( .a(G398), .b(G399), .O(G480) );
nand2 gate124( .a(G400), .b(G401), .O(G483) );
nand2 gate125( .a(G402), .b(G403), .O(G486) );
nand2 gate126( .a(G404), .b(G405), .O(G489) );
nand2 gate127( .a(G406), .b(G407), .O(G492) );
nand2 gate128( .a(G408), .b(G409), .O(G495) );
nand2 gate129( .a(G410), .b(G411), .O(G498) );

  xor2  gate575(.a(G413), .b(G412), .O(gate130inter0));
  nand2 gate576(.a(gate130inter0), .b(s_4), .O(gate130inter1));
  and2  gate577(.a(G413), .b(G412), .O(gate130inter2));
  inv1  gate578(.a(s_4), .O(gate130inter3));
  inv1  gate579(.a(s_5), .O(gate130inter4));
  nand2 gate580(.a(gate130inter4), .b(gate130inter3), .O(gate130inter5));
  nor2  gate581(.a(gate130inter5), .b(gate130inter2), .O(gate130inter6));
  inv1  gate582(.a(G412), .O(gate130inter7));
  inv1  gate583(.a(G413), .O(gate130inter8));
  nand2 gate584(.a(gate130inter8), .b(gate130inter7), .O(gate130inter9));
  nand2 gate585(.a(s_5), .b(gate130inter3), .O(gate130inter10));
  nor2  gate586(.a(gate130inter10), .b(gate130inter9), .O(gate130inter11));
  nor2  gate587(.a(gate130inter11), .b(gate130inter6), .O(gate130inter12));
  nand2 gate588(.a(gate130inter12), .b(gate130inter1), .O(G501));
nand2 gate131( .a(G414), .b(G415), .O(G504) );
nand2 gate132( .a(G416), .b(G417), .O(G507) );
nand2 gate133( .a(G418), .b(G419), .O(G510) );
nand2 gate134( .a(G420), .b(G421), .O(G513) );
nand2 gate135( .a(G422), .b(G423), .O(G516) );
nand2 gate136( .a(G424), .b(G425), .O(G519) );
nand2 gate137( .a(G426), .b(G429), .O(G522) );
nand2 gate138( .a(G432), .b(G435), .O(G525) );
nand2 gate139( .a(G438), .b(G441), .O(G528) );

  xor2  gate1191(.a(G447), .b(G444), .O(gate140inter0));
  nand2 gate1192(.a(gate140inter0), .b(s_92), .O(gate140inter1));
  and2  gate1193(.a(G447), .b(G444), .O(gate140inter2));
  inv1  gate1194(.a(s_92), .O(gate140inter3));
  inv1  gate1195(.a(s_93), .O(gate140inter4));
  nand2 gate1196(.a(gate140inter4), .b(gate140inter3), .O(gate140inter5));
  nor2  gate1197(.a(gate140inter5), .b(gate140inter2), .O(gate140inter6));
  inv1  gate1198(.a(G444), .O(gate140inter7));
  inv1  gate1199(.a(G447), .O(gate140inter8));
  nand2 gate1200(.a(gate140inter8), .b(gate140inter7), .O(gate140inter9));
  nand2 gate1201(.a(s_93), .b(gate140inter3), .O(gate140inter10));
  nor2  gate1202(.a(gate140inter10), .b(gate140inter9), .O(gate140inter11));
  nor2  gate1203(.a(gate140inter11), .b(gate140inter6), .O(gate140inter12));
  nand2 gate1204(.a(gate140inter12), .b(gate140inter1), .O(G531));
nand2 gate141( .a(G450), .b(G453), .O(G534) );
nand2 gate142( .a(G456), .b(G459), .O(G537) );
nand2 gate143( .a(G462), .b(G465), .O(G540) );
nand2 gate144( .a(G468), .b(G471), .O(G543) );
nand2 gate145( .a(G474), .b(G477), .O(G546) );
nand2 gate146( .a(G480), .b(G483), .O(G549) );
nand2 gate147( .a(G486), .b(G489), .O(G552) );
nand2 gate148( .a(G492), .b(G495), .O(G555) );
nand2 gate149( .a(G498), .b(G501), .O(G558) );
nand2 gate150( .a(G504), .b(G507), .O(G561) );
nand2 gate151( .a(G510), .b(G513), .O(G564) );
nand2 gate152( .a(G516), .b(G519), .O(G567) );
nand2 gate153( .a(G426), .b(G522), .O(G570) );
nand2 gate154( .a(G429), .b(G522), .O(G571) );
nand2 gate155( .a(G432), .b(G525), .O(G572) );
nand2 gate156( .a(G435), .b(G525), .O(G573) );
nand2 gate157( .a(G438), .b(G528), .O(G574) );
nand2 gate158( .a(G441), .b(G528), .O(G575) );
nand2 gate159( .a(G444), .b(G531), .O(G576) );
nand2 gate160( .a(G447), .b(G531), .O(G577) );
nand2 gate161( .a(G450), .b(G534), .O(G578) );
nand2 gate162( .a(G453), .b(G534), .O(G579) );

  xor2  gate925(.a(G537), .b(G456), .O(gate163inter0));
  nand2 gate926(.a(gate163inter0), .b(s_54), .O(gate163inter1));
  and2  gate927(.a(G537), .b(G456), .O(gate163inter2));
  inv1  gate928(.a(s_54), .O(gate163inter3));
  inv1  gate929(.a(s_55), .O(gate163inter4));
  nand2 gate930(.a(gate163inter4), .b(gate163inter3), .O(gate163inter5));
  nor2  gate931(.a(gate163inter5), .b(gate163inter2), .O(gate163inter6));
  inv1  gate932(.a(G456), .O(gate163inter7));
  inv1  gate933(.a(G537), .O(gate163inter8));
  nand2 gate934(.a(gate163inter8), .b(gate163inter7), .O(gate163inter9));
  nand2 gate935(.a(s_55), .b(gate163inter3), .O(gate163inter10));
  nor2  gate936(.a(gate163inter10), .b(gate163inter9), .O(gate163inter11));
  nor2  gate937(.a(gate163inter11), .b(gate163inter6), .O(gate163inter12));
  nand2 gate938(.a(gate163inter12), .b(gate163inter1), .O(G580));

  xor2  gate715(.a(G537), .b(G459), .O(gate164inter0));
  nand2 gate716(.a(gate164inter0), .b(s_24), .O(gate164inter1));
  and2  gate717(.a(G537), .b(G459), .O(gate164inter2));
  inv1  gate718(.a(s_24), .O(gate164inter3));
  inv1  gate719(.a(s_25), .O(gate164inter4));
  nand2 gate720(.a(gate164inter4), .b(gate164inter3), .O(gate164inter5));
  nor2  gate721(.a(gate164inter5), .b(gate164inter2), .O(gate164inter6));
  inv1  gate722(.a(G459), .O(gate164inter7));
  inv1  gate723(.a(G537), .O(gate164inter8));
  nand2 gate724(.a(gate164inter8), .b(gate164inter7), .O(gate164inter9));
  nand2 gate725(.a(s_25), .b(gate164inter3), .O(gate164inter10));
  nor2  gate726(.a(gate164inter10), .b(gate164inter9), .O(gate164inter11));
  nor2  gate727(.a(gate164inter11), .b(gate164inter6), .O(gate164inter12));
  nand2 gate728(.a(gate164inter12), .b(gate164inter1), .O(G581));
nand2 gate165( .a(G462), .b(G540), .O(G582) );
nand2 gate166( .a(G465), .b(G540), .O(G583) );
nand2 gate167( .a(G468), .b(G543), .O(G584) );
nand2 gate168( .a(G471), .b(G543), .O(G585) );
nand2 gate169( .a(G474), .b(G546), .O(G586) );

  xor2  gate897(.a(G546), .b(G477), .O(gate170inter0));
  nand2 gate898(.a(gate170inter0), .b(s_50), .O(gate170inter1));
  and2  gate899(.a(G546), .b(G477), .O(gate170inter2));
  inv1  gate900(.a(s_50), .O(gate170inter3));
  inv1  gate901(.a(s_51), .O(gate170inter4));
  nand2 gate902(.a(gate170inter4), .b(gate170inter3), .O(gate170inter5));
  nor2  gate903(.a(gate170inter5), .b(gate170inter2), .O(gate170inter6));
  inv1  gate904(.a(G477), .O(gate170inter7));
  inv1  gate905(.a(G546), .O(gate170inter8));
  nand2 gate906(.a(gate170inter8), .b(gate170inter7), .O(gate170inter9));
  nand2 gate907(.a(s_51), .b(gate170inter3), .O(gate170inter10));
  nor2  gate908(.a(gate170inter10), .b(gate170inter9), .O(gate170inter11));
  nor2  gate909(.a(gate170inter11), .b(gate170inter6), .O(gate170inter12));
  nand2 gate910(.a(gate170inter12), .b(gate170inter1), .O(G587));
nand2 gate171( .a(G480), .b(G549), .O(G588) );
nand2 gate172( .a(G483), .b(G549), .O(G589) );
nand2 gate173( .a(G486), .b(G552), .O(G590) );
nand2 gate174( .a(G489), .b(G552), .O(G591) );

  xor2  gate1037(.a(G555), .b(G492), .O(gate175inter0));
  nand2 gate1038(.a(gate175inter0), .b(s_70), .O(gate175inter1));
  and2  gate1039(.a(G555), .b(G492), .O(gate175inter2));
  inv1  gate1040(.a(s_70), .O(gate175inter3));
  inv1  gate1041(.a(s_71), .O(gate175inter4));
  nand2 gate1042(.a(gate175inter4), .b(gate175inter3), .O(gate175inter5));
  nor2  gate1043(.a(gate175inter5), .b(gate175inter2), .O(gate175inter6));
  inv1  gate1044(.a(G492), .O(gate175inter7));
  inv1  gate1045(.a(G555), .O(gate175inter8));
  nand2 gate1046(.a(gate175inter8), .b(gate175inter7), .O(gate175inter9));
  nand2 gate1047(.a(s_71), .b(gate175inter3), .O(gate175inter10));
  nor2  gate1048(.a(gate175inter10), .b(gate175inter9), .O(gate175inter11));
  nor2  gate1049(.a(gate175inter11), .b(gate175inter6), .O(gate175inter12));
  nand2 gate1050(.a(gate175inter12), .b(gate175inter1), .O(G592));
nand2 gate176( .a(G495), .b(G555), .O(G593) );
nand2 gate177( .a(G498), .b(G558), .O(G594) );
nand2 gate178( .a(G501), .b(G558), .O(G595) );

  xor2  gate1107(.a(G561), .b(G504), .O(gate179inter0));
  nand2 gate1108(.a(gate179inter0), .b(s_80), .O(gate179inter1));
  and2  gate1109(.a(G561), .b(G504), .O(gate179inter2));
  inv1  gate1110(.a(s_80), .O(gate179inter3));
  inv1  gate1111(.a(s_81), .O(gate179inter4));
  nand2 gate1112(.a(gate179inter4), .b(gate179inter3), .O(gate179inter5));
  nor2  gate1113(.a(gate179inter5), .b(gate179inter2), .O(gate179inter6));
  inv1  gate1114(.a(G504), .O(gate179inter7));
  inv1  gate1115(.a(G561), .O(gate179inter8));
  nand2 gate1116(.a(gate179inter8), .b(gate179inter7), .O(gate179inter9));
  nand2 gate1117(.a(s_81), .b(gate179inter3), .O(gate179inter10));
  nor2  gate1118(.a(gate179inter10), .b(gate179inter9), .O(gate179inter11));
  nor2  gate1119(.a(gate179inter11), .b(gate179inter6), .O(gate179inter12));
  nand2 gate1120(.a(gate179inter12), .b(gate179inter1), .O(G596));
nand2 gate180( .a(G507), .b(G561), .O(G597) );
nand2 gate181( .a(G510), .b(G564), .O(G598) );
nand2 gate182( .a(G513), .b(G564), .O(G599) );
nand2 gate183( .a(G516), .b(G567), .O(G600) );
nand2 gate184( .a(G519), .b(G567), .O(G601) );
nand2 gate185( .a(G570), .b(G571), .O(G602) );
nand2 gate186( .a(G572), .b(G573), .O(G607) );

  xor2  gate1233(.a(G575), .b(G574), .O(gate187inter0));
  nand2 gate1234(.a(gate187inter0), .b(s_98), .O(gate187inter1));
  and2  gate1235(.a(G575), .b(G574), .O(gate187inter2));
  inv1  gate1236(.a(s_98), .O(gate187inter3));
  inv1  gate1237(.a(s_99), .O(gate187inter4));
  nand2 gate1238(.a(gate187inter4), .b(gate187inter3), .O(gate187inter5));
  nor2  gate1239(.a(gate187inter5), .b(gate187inter2), .O(gate187inter6));
  inv1  gate1240(.a(G574), .O(gate187inter7));
  inv1  gate1241(.a(G575), .O(gate187inter8));
  nand2 gate1242(.a(gate187inter8), .b(gate187inter7), .O(gate187inter9));
  nand2 gate1243(.a(s_99), .b(gate187inter3), .O(gate187inter10));
  nor2  gate1244(.a(gate187inter10), .b(gate187inter9), .O(gate187inter11));
  nor2  gate1245(.a(gate187inter11), .b(gate187inter6), .O(gate187inter12));
  nand2 gate1246(.a(gate187inter12), .b(gate187inter1), .O(G612));
nand2 gate188( .a(G576), .b(G577), .O(G617) );
nand2 gate189( .a(G578), .b(G579), .O(G622) );
nand2 gate190( .a(G580), .b(G581), .O(G627) );
nand2 gate191( .a(G582), .b(G583), .O(G632) );
nand2 gate192( .a(G584), .b(G585), .O(G637) );
nand2 gate193( .a(G586), .b(G587), .O(G642) );
nand2 gate194( .a(G588), .b(G589), .O(G645) );
nand2 gate195( .a(G590), .b(G591), .O(G648) );
nand2 gate196( .a(G592), .b(G593), .O(G651) );
nand2 gate197( .a(G594), .b(G595), .O(G654) );
nand2 gate198( .a(G596), .b(G597), .O(G657) );
nand2 gate199( .a(G598), .b(G599), .O(G660) );

  xor2  gate1163(.a(G601), .b(G600), .O(gate200inter0));
  nand2 gate1164(.a(gate200inter0), .b(s_88), .O(gate200inter1));
  and2  gate1165(.a(G601), .b(G600), .O(gate200inter2));
  inv1  gate1166(.a(s_88), .O(gate200inter3));
  inv1  gate1167(.a(s_89), .O(gate200inter4));
  nand2 gate1168(.a(gate200inter4), .b(gate200inter3), .O(gate200inter5));
  nor2  gate1169(.a(gate200inter5), .b(gate200inter2), .O(gate200inter6));
  inv1  gate1170(.a(G600), .O(gate200inter7));
  inv1  gate1171(.a(G601), .O(gate200inter8));
  nand2 gate1172(.a(gate200inter8), .b(gate200inter7), .O(gate200inter9));
  nand2 gate1173(.a(s_89), .b(gate200inter3), .O(gate200inter10));
  nor2  gate1174(.a(gate200inter10), .b(gate200inter9), .O(gate200inter11));
  nor2  gate1175(.a(gate200inter11), .b(gate200inter6), .O(gate200inter12));
  nand2 gate1176(.a(gate200inter12), .b(gate200inter1), .O(G663));
nand2 gate201( .a(G602), .b(G607), .O(G666) );
nand2 gate202( .a(G612), .b(G617), .O(G669) );
nand2 gate203( .a(G602), .b(G612), .O(G672) );
nand2 gate204( .a(G607), .b(G617), .O(G675) );
nand2 gate205( .a(G622), .b(G627), .O(G678) );
nand2 gate206( .a(G632), .b(G637), .O(G681) );
nand2 gate207( .a(G622), .b(G632), .O(G684) );
nand2 gate208( .a(G627), .b(G637), .O(G687) );

  xor2  gate1205(.a(G666), .b(G602), .O(gate209inter0));
  nand2 gate1206(.a(gate209inter0), .b(s_94), .O(gate209inter1));
  and2  gate1207(.a(G666), .b(G602), .O(gate209inter2));
  inv1  gate1208(.a(s_94), .O(gate209inter3));
  inv1  gate1209(.a(s_95), .O(gate209inter4));
  nand2 gate1210(.a(gate209inter4), .b(gate209inter3), .O(gate209inter5));
  nor2  gate1211(.a(gate209inter5), .b(gate209inter2), .O(gate209inter6));
  inv1  gate1212(.a(G602), .O(gate209inter7));
  inv1  gate1213(.a(G666), .O(gate209inter8));
  nand2 gate1214(.a(gate209inter8), .b(gate209inter7), .O(gate209inter9));
  nand2 gate1215(.a(s_95), .b(gate209inter3), .O(gate209inter10));
  nor2  gate1216(.a(gate209inter10), .b(gate209inter9), .O(gate209inter11));
  nor2  gate1217(.a(gate209inter11), .b(gate209inter6), .O(gate209inter12));
  nand2 gate1218(.a(gate209inter12), .b(gate209inter1), .O(G690));
nand2 gate210( .a(G607), .b(G666), .O(G691) );
nand2 gate211( .a(G612), .b(G669), .O(G692) );
nand2 gate212( .a(G617), .b(G669), .O(G693) );
nand2 gate213( .a(G602), .b(G672), .O(G694) );
nand2 gate214( .a(G612), .b(G672), .O(G695) );
nand2 gate215( .a(G607), .b(G675), .O(G696) );
nand2 gate216( .a(G617), .b(G675), .O(G697) );
nand2 gate217( .a(G622), .b(G678), .O(G698) );

  xor2  gate589(.a(G678), .b(G627), .O(gate218inter0));
  nand2 gate590(.a(gate218inter0), .b(s_6), .O(gate218inter1));
  and2  gate591(.a(G678), .b(G627), .O(gate218inter2));
  inv1  gate592(.a(s_6), .O(gate218inter3));
  inv1  gate593(.a(s_7), .O(gate218inter4));
  nand2 gate594(.a(gate218inter4), .b(gate218inter3), .O(gate218inter5));
  nor2  gate595(.a(gate218inter5), .b(gate218inter2), .O(gate218inter6));
  inv1  gate596(.a(G627), .O(gate218inter7));
  inv1  gate597(.a(G678), .O(gate218inter8));
  nand2 gate598(.a(gate218inter8), .b(gate218inter7), .O(gate218inter9));
  nand2 gate599(.a(s_7), .b(gate218inter3), .O(gate218inter10));
  nor2  gate600(.a(gate218inter10), .b(gate218inter9), .O(gate218inter11));
  nor2  gate601(.a(gate218inter11), .b(gate218inter6), .O(gate218inter12));
  nand2 gate602(.a(gate218inter12), .b(gate218inter1), .O(G699));
nand2 gate219( .a(G632), .b(G681), .O(G700) );

  xor2  gate1023(.a(G681), .b(G637), .O(gate220inter0));
  nand2 gate1024(.a(gate220inter0), .b(s_68), .O(gate220inter1));
  and2  gate1025(.a(G681), .b(G637), .O(gate220inter2));
  inv1  gate1026(.a(s_68), .O(gate220inter3));
  inv1  gate1027(.a(s_69), .O(gate220inter4));
  nand2 gate1028(.a(gate220inter4), .b(gate220inter3), .O(gate220inter5));
  nor2  gate1029(.a(gate220inter5), .b(gate220inter2), .O(gate220inter6));
  inv1  gate1030(.a(G637), .O(gate220inter7));
  inv1  gate1031(.a(G681), .O(gate220inter8));
  nand2 gate1032(.a(gate220inter8), .b(gate220inter7), .O(gate220inter9));
  nand2 gate1033(.a(s_69), .b(gate220inter3), .O(gate220inter10));
  nor2  gate1034(.a(gate220inter10), .b(gate220inter9), .O(gate220inter11));
  nor2  gate1035(.a(gate220inter11), .b(gate220inter6), .O(gate220inter12));
  nand2 gate1036(.a(gate220inter12), .b(gate220inter1), .O(G701));
nand2 gate221( .a(G622), .b(G684), .O(G702) );
nand2 gate222( .a(G632), .b(G684), .O(G703) );

  xor2  gate757(.a(G687), .b(G627), .O(gate223inter0));
  nand2 gate758(.a(gate223inter0), .b(s_30), .O(gate223inter1));
  and2  gate759(.a(G687), .b(G627), .O(gate223inter2));
  inv1  gate760(.a(s_30), .O(gate223inter3));
  inv1  gate761(.a(s_31), .O(gate223inter4));
  nand2 gate762(.a(gate223inter4), .b(gate223inter3), .O(gate223inter5));
  nor2  gate763(.a(gate223inter5), .b(gate223inter2), .O(gate223inter6));
  inv1  gate764(.a(G627), .O(gate223inter7));
  inv1  gate765(.a(G687), .O(gate223inter8));
  nand2 gate766(.a(gate223inter8), .b(gate223inter7), .O(gate223inter9));
  nand2 gate767(.a(s_31), .b(gate223inter3), .O(gate223inter10));
  nor2  gate768(.a(gate223inter10), .b(gate223inter9), .O(gate223inter11));
  nor2  gate769(.a(gate223inter11), .b(gate223inter6), .O(gate223inter12));
  nand2 gate770(.a(gate223inter12), .b(gate223inter1), .O(G704));
nand2 gate224( .a(G637), .b(G687), .O(G705) );
nand2 gate225( .a(G690), .b(G691), .O(G706) );
nand2 gate226( .a(G692), .b(G693), .O(G709) );
nand2 gate227( .a(G694), .b(G695), .O(G712) );
nand2 gate228( .a(G696), .b(G697), .O(G715) );
nand2 gate229( .a(G698), .b(G699), .O(G718) );
nand2 gate230( .a(G700), .b(G701), .O(G721) );

  xor2  gate1065(.a(G703), .b(G702), .O(gate231inter0));
  nand2 gate1066(.a(gate231inter0), .b(s_74), .O(gate231inter1));
  and2  gate1067(.a(G703), .b(G702), .O(gate231inter2));
  inv1  gate1068(.a(s_74), .O(gate231inter3));
  inv1  gate1069(.a(s_75), .O(gate231inter4));
  nand2 gate1070(.a(gate231inter4), .b(gate231inter3), .O(gate231inter5));
  nor2  gate1071(.a(gate231inter5), .b(gate231inter2), .O(gate231inter6));
  inv1  gate1072(.a(G702), .O(gate231inter7));
  inv1  gate1073(.a(G703), .O(gate231inter8));
  nand2 gate1074(.a(gate231inter8), .b(gate231inter7), .O(gate231inter9));
  nand2 gate1075(.a(s_75), .b(gate231inter3), .O(gate231inter10));
  nor2  gate1076(.a(gate231inter10), .b(gate231inter9), .O(gate231inter11));
  nor2  gate1077(.a(gate231inter11), .b(gate231inter6), .O(gate231inter12));
  nand2 gate1078(.a(gate231inter12), .b(gate231inter1), .O(G724));

  xor2  gate1149(.a(G705), .b(G704), .O(gate232inter0));
  nand2 gate1150(.a(gate232inter0), .b(s_86), .O(gate232inter1));
  and2  gate1151(.a(G705), .b(G704), .O(gate232inter2));
  inv1  gate1152(.a(s_86), .O(gate232inter3));
  inv1  gate1153(.a(s_87), .O(gate232inter4));
  nand2 gate1154(.a(gate232inter4), .b(gate232inter3), .O(gate232inter5));
  nor2  gate1155(.a(gate232inter5), .b(gate232inter2), .O(gate232inter6));
  inv1  gate1156(.a(G704), .O(gate232inter7));
  inv1  gate1157(.a(G705), .O(gate232inter8));
  nand2 gate1158(.a(gate232inter8), .b(gate232inter7), .O(gate232inter9));
  nand2 gate1159(.a(s_87), .b(gate232inter3), .O(gate232inter10));
  nor2  gate1160(.a(gate232inter10), .b(gate232inter9), .O(gate232inter11));
  nor2  gate1161(.a(gate232inter11), .b(gate232inter6), .O(gate232inter12));
  nand2 gate1162(.a(gate232inter12), .b(gate232inter1), .O(G727));
nand2 gate233( .a(G242), .b(G718), .O(G730) );

  xor2  gate1177(.a(G721), .b(G245), .O(gate234inter0));
  nand2 gate1178(.a(gate234inter0), .b(s_90), .O(gate234inter1));
  and2  gate1179(.a(G721), .b(G245), .O(gate234inter2));
  inv1  gate1180(.a(s_90), .O(gate234inter3));
  inv1  gate1181(.a(s_91), .O(gate234inter4));
  nand2 gate1182(.a(gate234inter4), .b(gate234inter3), .O(gate234inter5));
  nor2  gate1183(.a(gate234inter5), .b(gate234inter2), .O(gate234inter6));
  inv1  gate1184(.a(G245), .O(gate234inter7));
  inv1  gate1185(.a(G721), .O(gate234inter8));
  nand2 gate1186(.a(gate234inter8), .b(gate234inter7), .O(gate234inter9));
  nand2 gate1187(.a(s_91), .b(gate234inter3), .O(gate234inter10));
  nor2  gate1188(.a(gate234inter10), .b(gate234inter9), .O(gate234inter11));
  nor2  gate1189(.a(gate234inter11), .b(gate234inter6), .O(gate234inter12));
  nand2 gate1190(.a(gate234inter12), .b(gate234inter1), .O(G733));
nand2 gate235( .a(G248), .b(G724), .O(G736) );
nand2 gate236( .a(G251), .b(G727), .O(G739) );
nand2 gate237( .a(G254), .b(G706), .O(G742) );
nand2 gate238( .a(G257), .b(G709), .O(G745) );
nand2 gate239( .a(G260), .b(G712), .O(G748) );
nand2 gate240( .a(G263), .b(G715), .O(G751) );
nand2 gate241( .a(G242), .b(G730), .O(G754) );
nand2 gate242( .a(G718), .b(G730), .O(G755) );

  xor2  gate911(.a(G733), .b(G245), .O(gate243inter0));
  nand2 gate912(.a(gate243inter0), .b(s_52), .O(gate243inter1));
  and2  gate913(.a(G733), .b(G245), .O(gate243inter2));
  inv1  gate914(.a(s_52), .O(gate243inter3));
  inv1  gate915(.a(s_53), .O(gate243inter4));
  nand2 gate916(.a(gate243inter4), .b(gate243inter3), .O(gate243inter5));
  nor2  gate917(.a(gate243inter5), .b(gate243inter2), .O(gate243inter6));
  inv1  gate918(.a(G245), .O(gate243inter7));
  inv1  gate919(.a(G733), .O(gate243inter8));
  nand2 gate920(.a(gate243inter8), .b(gate243inter7), .O(gate243inter9));
  nand2 gate921(.a(s_53), .b(gate243inter3), .O(gate243inter10));
  nor2  gate922(.a(gate243inter10), .b(gate243inter9), .O(gate243inter11));
  nor2  gate923(.a(gate243inter11), .b(gate243inter6), .O(gate243inter12));
  nand2 gate924(.a(gate243inter12), .b(gate243inter1), .O(G756));
nand2 gate244( .a(G721), .b(G733), .O(G757) );
nand2 gate245( .a(G248), .b(G736), .O(G758) );

  xor2  gate953(.a(G736), .b(G724), .O(gate246inter0));
  nand2 gate954(.a(gate246inter0), .b(s_58), .O(gate246inter1));
  and2  gate955(.a(G736), .b(G724), .O(gate246inter2));
  inv1  gate956(.a(s_58), .O(gate246inter3));
  inv1  gate957(.a(s_59), .O(gate246inter4));
  nand2 gate958(.a(gate246inter4), .b(gate246inter3), .O(gate246inter5));
  nor2  gate959(.a(gate246inter5), .b(gate246inter2), .O(gate246inter6));
  inv1  gate960(.a(G724), .O(gate246inter7));
  inv1  gate961(.a(G736), .O(gate246inter8));
  nand2 gate962(.a(gate246inter8), .b(gate246inter7), .O(gate246inter9));
  nand2 gate963(.a(s_59), .b(gate246inter3), .O(gate246inter10));
  nor2  gate964(.a(gate246inter10), .b(gate246inter9), .O(gate246inter11));
  nor2  gate965(.a(gate246inter11), .b(gate246inter6), .O(gate246inter12));
  nand2 gate966(.a(gate246inter12), .b(gate246inter1), .O(G759));
nand2 gate247( .a(G251), .b(G739), .O(G760) );
nand2 gate248( .a(G727), .b(G739), .O(G761) );
nand2 gate249( .a(G254), .b(G742), .O(G762) );
nand2 gate250( .a(G706), .b(G742), .O(G763) );
nand2 gate251( .a(G257), .b(G745), .O(G764) );
nand2 gate252( .a(G709), .b(G745), .O(G765) );
nand2 gate253( .a(G260), .b(G748), .O(G766) );
nand2 gate254( .a(G712), .b(G748), .O(G767) );
nand2 gate255( .a(G263), .b(G751), .O(G768) );

  xor2  gate1247(.a(G751), .b(G715), .O(gate256inter0));
  nand2 gate1248(.a(gate256inter0), .b(s_100), .O(gate256inter1));
  and2  gate1249(.a(G751), .b(G715), .O(gate256inter2));
  inv1  gate1250(.a(s_100), .O(gate256inter3));
  inv1  gate1251(.a(s_101), .O(gate256inter4));
  nand2 gate1252(.a(gate256inter4), .b(gate256inter3), .O(gate256inter5));
  nor2  gate1253(.a(gate256inter5), .b(gate256inter2), .O(gate256inter6));
  inv1  gate1254(.a(G715), .O(gate256inter7));
  inv1  gate1255(.a(G751), .O(gate256inter8));
  nand2 gate1256(.a(gate256inter8), .b(gate256inter7), .O(gate256inter9));
  nand2 gate1257(.a(s_101), .b(gate256inter3), .O(gate256inter10));
  nor2  gate1258(.a(gate256inter10), .b(gate256inter9), .O(gate256inter11));
  nor2  gate1259(.a(gate256inter11), .b(gate256inter6), .O(gate256inter12));
  nand2 gate1260(.a(gate256inter12), .b(gate256inter1), .O(G769));
nand2 gate257( .a(G754), .b(G755), .O(G770) );
nand2 gate258( .a(G756), .b(G757), .O(G773) );
nand2 gate259( .a(G758), .b(G759), .O(G776) );
nand2 gate260( .a(G760), .b(G761), .O(G779) );
nand2 gate261( .a(G762), .b(G763), .O(G782) );
nand2 gate262( .a(G764), .b(G765), .O(G785) );
nand2 gate263( .a(G766), .b(G767), .O(G788) );
nand2 gate264( .a(G768), .b(G769), .O(G791) );

  xor2  gate1009(.a(G770), .b(G642), .O(gate265inter0));
  nand2 gate1010(.a(gate265inter0), .b(s_66), .O(gate265inter1));
  and2  gate1011(.a(G770), .b(G642), .O(gate265inter2));
  inv1  gate1012(.a(s_66), .O(gate265inter3));
  inv1  gate1013(.a(s_67), .O(gate265inter4));
  nand2 gate1014(.a(gate265inter4), .b(gate265inter3), .O(gate265inter5));
  nor2  gate1015(.a(gate265inter5), .b(gate265inter2), .O(gate265inter6));
  inv1  gate1016(.a(G642), .O(gate265inter7));
  inv1  gate1017(.a(G770), .O(gate265inter8));
  nand2 gate1018(.a(gate265inter8), .b(gate265inter7), .O(gate265inter9));
  nand2 gate1019(.a(s_67), .b(gate265inter3), .O(gate265inter10));
  nor2  gate1020(.a(gate265inter10), .b(gate265inter9), .O(gate265inter11));
  nor2  gate1021(.a(gate265inter11), .b(gate265inter6), .O(gate265inter12));
  nand2 gate1022(.a(gate265inter12), .b(gate265inter1), .O(G794));
nand2 gate266( .a(G645), .b(G773), .O(G797) );
nand2 gate267( .a(G648), .b(G776), .O(G800) );
nand2 gate268( .a(G651), .b(G779), .O(G803) );
nand2 gate269( .a(G654), .b(G782), .O(G806) );
nand2 gate270( .a(G657), .b(G785), .O(G809) );
nand2 gate271( .a(G660), .b(G788), .O(G812) );

  xor2  gate743(.a(G791), .b(G663), .O(gate272inter0));
  nand2 gate744(.a(gate272inter0), .b(s_28), .O(gate272inter1));
  and2  gate745(.a(G791), .b(G663), .O(gate272inter2));
  inv1  gate746(.a(s_28), .O(gate272inter3));
  inv1  gate747(.a(s_29), .O(gate272inter4));
  nand2 gate748(.a(gate272inter4), .b(gate272inter3), .O(gate272inter5));
  nor2  gate749(.a(gate272inter5), .b(gate272inter2), .O(gate272inter6));
  inv1  gate750(.a(G663), .O(gate272inter7));
  inv1  gate751(.a(G791), .O(gate272inter8));
  nand2 gate752(.a(gate272inter8), .b(gate272inter7), .O(gate272inter9));
  nand2 gate753(.a(s_29), .b(gate272inter3), .O(gate272inter10));
  nor2  gate754(.a(gate272inter10), .b(gate272inter9), .O(gate272inter11));
  nor2  gate755(.a(gate272inter11), .b(gate272inter6), .O(gate272inter12));
  nand2 gate756(.a(gate272inter12), .b(gate272inter1), .O(G815));
nand2 gate273( .a(G642), .b(G794), .O(G818) );
nand2 gate274( .a(G770), .b(G794), .O(G819) );
nand2 gate275( .a(G645), .b(G797), .O(G820) );
nand2 gate276( .a(G773), .b(G797), .O(G821) );
nand2 gate277( .a(G648), .b(G800), .O(G822) );
nand2 gate278( .a(G776), .b(G800), .O(G823) );
nand2 gate279( .a(G651), .b(G803), .O(G824) );
nand2 gate280( .a(G779), .b(G803), .O(G825) );

  xor2  gate603(.a(G806), .b(G654), .O(gate281inter0));
  nand2 gate604(.a(gate281inter0), .b(s_8), .O(gate281inter1));
  and2  gate605(.a(G806), .b(G654), .O(gate281inter2));
  inv1  gate606(.a(s_8), .O(gate281inter3));
  inv1  gate607(.a(s_9), .O(gate281inter4));
  nand2 gate608(.a(gate281inter4), .b(gate281inter3), .O(gate281inter5));
  nor2  gate609(.a(gate281inter5), .b(gate281inter2), .O(gate281inter6));
  inv1  gate610(.a(G654), .O(gate281inter7));
  inv1  gate611(.a(G806), .O(gate281inter8));
  nand2 gate612(.a(gate281inter8), .b(gate281inter7), .O(gate281inter9));
  nand2 gate613(.a(s_9), .b(gate281inter3), .O(gate281inter10));
  nor2  gate614(.a(gate281inter10), .b(gate281inter9), .O(gate281inter11));
  nor2  gate615(.a(gate281inter11), .b(gate281inter6), .O(gate281inter12));
  nand2 gate616(.a(gate281inter12), .b(gate281inter1), .O(G826));
nand2 gate282( .a(G782), .b(G806), .O(G827) );
nand2 gate283( .a(G657), .b(G809), .O(G828) );
nand2 gate284( .a(G785), .b(G809), .O(G829) );
nand2 gate285( .a(G660), .b(G812), .O(G830) );
nand2 gate286( .a(G788), .b(G812), .O(G831) );
nand2 gate287( .a(G663), .b(G815), .O(G832) );
nand2 gate288( .a(G791), .b(G815), .O(G833) );
nand2 gate289( .a(G818), .b(G819), .O(G834) );
nand2 gate290( .a(G820), .b(G821), .O(G847) );

  xor2  gate785(.a(G823), .b(G822), .O(gate291inter0));
  nand2 gate786(.a(gate291inter0), .b(s_34), .O(gate291inter1));
  and2  gate787(.a(G823), .b(G822), .O(gate291inter2));
  inv1  gate788(.a(s_34), .O(gate291inter3));
  inv1  gate789(.a(s_35), .O(gate291inter4));
  nand2 gate790(.a(gate291inter4), .b(gate291inter3), .O(gate291inter5));
  nor2  gate791(.a(gate291inter5), .b(gate291inter2), .O(gate291inter6));
  inv1  gate792(.a(G822), .O(gate291inter7));
  inv1  gate793(.a(G823), .O(gate291inter8));
  nand2 gate794(.a(gate291inter8), .b(gate291inter7), .O(gate291inter9));
  nand2 gate795(.a(s_35), .b(gate291inter3), .O(gate291inter10));
  nor2  gate796(.a(gate291inter10), .b(gate291inter9), .O(gate291inter11));
  nor2  gate797(.a(gate291inter11), .b(gate291inter6), .O(gate291inter12));
  nand2 gate798(.a(gate291inter12), .b(gate291inter1), .O(G860));
nand2 gate292( .a(G824), .b(G825), .O(G873) );
nand2 gate293( .a(G828), .b(G829), .O(G886) );
nand2 gate294( .a(G832), .b(G833), .O(G899) );
nand2 gate295( .a(G830), .b(G831), .O(G912) );
nand2 gate296( .a(G826), .b(G827), .O(G925) );
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );
nand2 gate387( .a(G1), .b(G1036), .O(G1132) );

  xor2  gate659(.a(G1039), .b(G2), .O(gate388inter0));
  nand2 gate660(.a(gate388inter0), .b(s_16), .O(gate388inter1));
  and2  gate661(.a(G1039), .b(G2), .O(gate388inter2));
  inv1  gate662(.a(s_16), .O(gate388inter3));
  inv1  gate663(.a(s_17), .O(gate388inter4));
  nand2 gate664(.a(gate388inter4), .b(gate388inter3), .O(gate388inter5));
  nor2  gate665(.a(gate388inter5), .b(gate388inter2), .O(gate388inter6));
  inv1  gate666(.a(G2), .O(gate388inter7));
  inv1  gate667(.a(G1039), .O(gate388inter8));
  nand2 gate668(.a(gate388inter8), .b(gate388inter7), .O(gate388inter9));
  nand2 gate669(.a(s_17), .b(gate388inter3), .O(gate388inter10));
  nor2  gate670(.a(gate388inter10), .b(gate388inter9), .O(gate388inter11));
  nor2  gate671(.a(gate388inter11), .b(gate388inter6), .O(gate388inter12));
  nand2 gate672(.a(gate388inter12), .b(gate388inter1), .O(G1135));
nand2 gate389( .a(G3), .b(G1042), .O(G1138) );

  xor2  gate799(.a(G1045), .b(G4), .O(gate390inter0));
  nand2 gate800(.a(gate390inter0), .b(s_36), .O(gate390inter1));
  and2  gate801(.a(G1045), .b(G4), .O(gate390inter2));
  inv1  gate802(.a(s_36), .O(gate390inter3));
  inv1  gate803(.a(s_37), .O(gate390inter4));
  nand2 gate804(.a(gate390inter4), .b(gate390inter3), .O(gate390inter5));
  nor2  gate805(.a(gate390inter5), .b(gate390inter2), .O(gate390inter6));
  inv1  gate806(.a(G4), .O(gate390inter7));
  inv1  gate807(.a(G1045), .O(gate390inter8));
  nand2 gate808(.a(gate390inter8), .b(gate390inter7), .O(gate390inter9));
  nand2 gate809(.a(s_37), .b(gate390inter3), .O(gate390inter10));
  nor2  gate810(.a(gate390inter10), .b(gate390inter9), .O(gate390inter11));
  nor2  gate811(.a(gate390inter11), .b(gate390inter6), .O(gate390inter12));
  nand2 gate812(.a(gate390inter12), .b(gate390inter1), .O(G1141));
nand2 gate391( .a(G5), .b(G1048), .O(G1144) );
nand2 gate392( .a(G6), .b(G1051), .O(G1147) );
nand2 gate393( .a(G7), .b(G1054), .O(G1150) );
nand2 gate394( .a(G8), .b(G1057), .O(G1153) );
nand2 gate395( .a(G9), .b(G1060), .O(G1156) );

  xor2  gate645(.a(G1063), .b(G10), .O(gate396inter0));
  nand2 gate646(.a(gate396inter0), .b(s_14), .O(gate396inter1));
  and2  gate647(.a(G1063), .b(G10), .O(gate396inter2));
  inv1  gate648(.a(s_14), .O(gate396inter3));
  inv1  gate649(.a(s_15), .O(gate396inter4));
  nand2 gate650(.a(gate396inter4), .b(gate396inter3), .O(gate396inter5));
  nor2  gate651(.a(gate396inter5), .b(gate396inter2), .O(gate396inter6));
  inv1  gate652(.a(G10), .O(gate396inter7));
  inv1  gate653(.a(G1063), .O(gate396inter8));
  nand2 gate654(.a(gate396inter8), .b(gate396inter7), .O(gate396inter9));
  nand2 gate655(.a(s_15), .b(gate396inter3), .O(gate396inter10));
  nor2  gate656(.a(gate396inter10), .b(gate396inter9), .O(gate396inter11));
  nor2  gate657(.a(gate396inter11), .b(gate396inter6), .O(gate396inter12));
  nand2 gate658(.a(gate396inter12), .b(gate396inter1), .O(G1159));
nand2 gate397( .a(G11), .b(G1066), .O(G1162) );
nand2 gate398( .a(G12), .b(G1069), .O(G1165) );
nand2 gate399( .a(G13), .b(G1072), .O(G1168) );
nand2 gate400( .a(G14), .b(G1075), .O(G1171) );
nand2 gate401( .a(G15), .b(G1078), .O(G1174) );
nand2 gate402( .a(G16), .b(G1081), .O(G1177) );
nand2 gate403( .a(G17), .b(G1084), .O(G1180) );
nand2 gate404( .a(G18), .b(G1087), .O(G1183) );
nand2 gate405( .a(G19), .b(G1090), .O(G1186) );
nand2 gate406( .a(G20), .b(G1093), .O(G1189) );
nand2 gate407( .a(G21), .b(G1096), .O(G1192) );
nand2 gate408( .a(G22), .b(G1099), .O(G1195) );
nand2 gate409( .a(G23), .b(G1102), .O(G1198) );
nand2 gate410( .a(G24), .b(G1105), .O(G1201) );
nand2 gate411( .a(G25), .b(G1108), .O(G1204) );
nand2 gate412( .a(G26), .b(G1111), .O(G1207) );
nand2 gate413( .a(G27), .b(G1114), .O(G1210) );
nand2 gate414( .a(G28), .b(G1117), .O(G1213) );
nand2 gate415( .a(G29), .b(G1120), .O(G1216) );
nand2 gate416( .a(G30), .b(G1123), .O(G1219) );
nand2 gate417( .a(G31), .b(G1126), .O(G1222) );
nand2 gate418( .a(G32), .b(G1129), .O(G1225) );
nand2 gate419( .a(G1), .b(G1132), .O(G1228) );
nand2 gate420( .a(G1036), .b(G1132), .O(G1229) );
nand2 gate421( .a(G2), .b(G1135), .O(G1230) );
nand2 gate422( .a(G1039), .b(G1135), .O(G1231) );
nand2 gate423( .a(G3), .b(G1138), .O(G1232) );
nand2 gate424( .a(G1042), .b(G1138), .O(G1233) );
nand2 gate425( .a(G4), .b(G1141), .O(G1234) );
nand2 gate426( .a(G1045), .b(G1141), .O(G1235) );
nand2 gate427( .a(G5), .b(G1144), .O(G1236) );
nand2 gate428( .a(G1048), .b(G1144), .O(G1237) );
nand2 gate429( .a(G6), .b(G1147), .O(G1238) );
nand2 gate430( .a(G1051), .b(G1147), .O(G1239) );

  xor2  gate561(.a(G1150), .b(G7), .O(gate431inter0));
  nand2 gate562(.a(gate431inter0), .b(s_2), .O(gate431inter1));
  and2  gate563(.a(G1150), .b(G7), .O(gate431inter2));
  inv1  gate564(.a(s_2), .O(gate431inter3));
  inv1  gate565(.a(s_3), .O(gate431inter4));
  nand2 gate566(.a(gate431inter4), .b(gate431inter3), .O(gate431inter5));
  nor2  gate567(.a(gate431inter5), .b(gate431inter2), .O(gate431inter6));
  inv1  gate568(.a(G7), .O(gate431inter7));
  inv1  gate569(.a(G1150), .O(gate431inter8));
  nand2 gate570(.a(gate431inter8), .b(gate431inter7), .O(gate431inter9));
  nand2 gate571(.a(s_3), .b(gate431inter3), .O(gate431inter10));
  nor2  gate572(.a(gate431inter10), .b(gate431inter9), .O(gate431inter11));
  nor2  gate573(.a(gate431inter11), .b(gate431inter6), .O(gate431inter12));
  nand2 gate574(.a(gate431inter12), .b(gate431inter1), .O(G1240));
nand2 gate432( .a(G1054), .b(G1150), .O(G1241) );
nand2 gate433( .a(G8), .b(G1153), .O(G1242) );
nand2 gate434( .a(G1057), .b(G1153), .O(G1243) );
nand2 gate435( .a(G9), .b(G1156), .O(G1244) );
nand2 gate436( .a(G1060), .b(G1156), .O(G1245) );
nand2 gate437( .a(G10), .b(G1159), .O(G1246) );

  xor2  gate967(.a(G1159), .b(G1063), .O(gate438inter0));
  nand2 gate968(.a(gate438inter0), .b(s_60), .O(gate438inter1));
  and2  gate969(.a(G1159), .b(G1063), .O(gate438inter2));
  inv1  gate970(.a(s_60), .O(gate438inter3));
  inv1  gate971(.a(s_61), .O(gate438inter4));
  nand2 gate972(.a(gate438inter4), .b(gate438inter3), .O(gate438inter5));
  nor2  gate973(.a(gate438inter5), .b(gate438inter2), .O(gate438inter6));
  inv1  gate974(.a(G1063), .O(gate438inter7));
  inv1  gate975(.a(G1159), .O(gate438inter8));
  nand2 gate976(.a(gate438inter8), .b(gate438inter7), .O(gate438inter9));
  nand2 gate977(.a(s_61), .b(gate438inter3), .O(gate438inter10));
  nor2  gate978(.a(gate438inter10), .b(gate438inter9), .O(gate438inter11));
  nor2  gate979(.a(gate438inter11), .b(gate438inter6), .O(gate438inter12));
  nand2 gate980(.a(gate438inter12), .b(gate438inter1), .O(G1247));

  xor2  gate827(.a(G1162), .b(G11), .O(gate439inter0));
  nand2 gate828(.a(gate439inter0), .b(s_40), .O(gate439inter1));
  and2  gate829(.a(G1162), .b(G11), .O(gate439inter2));
  inv1  gate830(.a(s_40), .O(gate439inter3));
  inv1  gate831(.a(s_41), .O(gate439inter4));
  nand2 gate832(.a(gate439inter4), .b(gate439inter3), .O(gate439inter5));
  nor2  gate833(.a(gate439inter5), .b(gate439inter2), .O(gate439inter6));
  inv1  gate834(.a(G11), .O(gate439inter7));
  inv1  gate835(.a(G1162), .O(gate439inter8));
  nand2 gate836(.a(gate439inter8), .b(gate439inter7), .O(gate439inter9));
  nand2 gate837(.a(s_41), .b(gate439inter3), .O(gate439inter10));
  nor2  gate838(.a(gate439inter10), .b(gate439inter9), .O(gate439inter11));
  nor2  gate839(.a(gate439inter11), .b(gate439inter6), .O(gate439inter12));
  nand2 gate840(.a(gate439inter12), .b(gate439inter1), .O(G1248));
nand2 gate440( .a(G1066), .b(G1162), .O(G1249) );

  xor2  gate1219(.a(G1165), .b(G12), .O(gate441inter0));
  nand2 gate1220(.a(gate441inter0), .b(s_96), .O(gate441inter1));
  and2  gate1221(.a(G1165), .b(G12), .O(gate441inter2));
  inv1  gate1222(.a(s_96), .O(gate441inter3));
  inv1  gate1223(.a(s_97), .O(gate441inter4));
  nand2 gate1224(.a(gate441inter4), .b(gate441inter3), .O(gate441inter5));
  nor2  gate1225(.a(gate441inter5), .b(gate441inter2), .O(gate441inter6));
  inv1  gate1226(.a(G12), .O(gate441inter7));
  inv1  gate1227(.a(G1165), .O(gate441inter8));
  nand2 gate1228(.a(gate441inter8), .b(gate441inter7), .O(gate441inter9));
  nand2 gate1229(.a(s_97), .b(gate441inter3), .O(gate441inter10));
  nor2  gate1230(.a(gate441inter10), .b(gate441inter9), .O(gate441inter11));
  nor2  gate1231(.a(gate441inter11), .b(gate441inter6), .O(gate441inter12));
  nand2 gate1232(.a(gate441inter12), .b(gate441inter1), .O(G1250));
nand2 gate442( .a(G1069), .b(G1165), .O(G1251) );
nand2 gate443( .a(G13), .b(G1168), .O(G1252) );
nand2 gate444( .a(G1072), .b(G1168), .O(G1253) );
nand2 gate445( .a(G14), .b(G1171), .O(G1254) );
nand2 gate446( .a(G1075), .b(G1171), .O(G1255) );
nand2 gate447( .a(G15), .b(G1174), .O(G1256) );
nand2 gate448( .a(G1078), .b(G1174), .O(G1257) );
nand2 gate449( .a(G16), .b(G1177), .O(G1258) );
nand2 gate450( .a(G1081), .b(G1177), .O(G1259) );
nand2 gate451( .a(G17), .b(G1180), .O(G1260) );
nand2 gate452( .a(G1084), .b(G1180), .O(G1261) );

  xor2  gate673(.a(G1183), .b(G18), .O(gate453inter0));
  nand2 gate674(.a(gate453inter0), .b(s_18), .O(gate453inter1));
  and2  gate675(.a(G1183), .b(G18), .O(gate453inter2));
  inv1  gate676(.a(s_18), .O(gate453inter3));
  inv1  gate677(.a(s_19), .O(gate453inter4));
  nand2 gate678(.a(gate453inter4), .b(gate453inter3), .O(gate453inter5));
  nor2  gate679(.a(gate453inter5), .b(gate453inter2), .O(gate453inter6));
  inv1  gate680(.a(G18), .O(gate453inter7));
  inv1  gate681(.a(G1183), .O(gate453inter8));
  nand2 gate682(.a(gate453inter8), .b(gate453inter7), .O(gate453inter9));
  nand2 gate683(.a(s_19), .b(gate453inter3), .O(gate453inter10));
  nor2  gate684(.a(gate453inter10), .b(gate453inter9), .O(gate453inter11));
  nor2  gate685(.a(gate453inter11), .b(gate453inter6), .O(gate453inter12));
  nand2 gate686(.a(gate453inter12), .b(gate453inter1), .O(G1262));

  xor2  gate701(.a(G1183), .b(G1087), .O(gate454inter0));
  nand2 gate702(.a(gate454inter0), .b(s_22), .O(gate454inter1));
  and2  gate703(.a(G1183), .b(G1087), .O(gate454inter2));
  inv1  gate704(.a(s_22), .O(gate454inter3));
  inv1  gate705(.a(s_23), .O(gate454inter4));
  nand2 gate706(.a(gate454inter4), .b(gate454inter3), .O(gate454inter5));
  nor2  gate707(.a(gate454inter5), .b(gate454inter2), .O(gate454inter6));
  inv1  gate708(.a(G1087), .O(gate454inter7));
  inv1  gate709(.a(G1183), .O(gate454inter8));
  nand2 gate710(.a(gate454inter8), .b(gate454inter7), .O(gate454inter9));
  nand2 gate711(.a(s_23), .b(gate454inter3), .O(gate454inter10));
  nor2  gate712(.a(gate454inter10), .b(gate454inter9), .O(gate454inter11));
  nor2  gate713(.a(gate454inter11), .b(gate454inter6), .O(gate454inter12));
  nand2 gate714(.a(gate454inter12), .b(gate454inter1), .O(G1263));
nand2 gate455( .a(G19), .b(G1186), .O(G1264) );
nand2 gate456( .a(G1090), .b(G1186), .O(G1265) );
nand2 gate457( .a(G20), .b(G1189), .O(G1266) );
nand2 gate458( .a(G1093), .b(G1189), .O(G1267) );
nand2 gate459( .a(G21), .b(G1192), .O(G1268) );
nand2 gate460( .a(G1096), .b(G1192), .O(G1269) );
nand2 gate461( .a(G22), .b(G1195), .O(G1270) );

  xor2  gate687(.a(G1195), .b(G1099), .O(gate462inter0));
  nand2 gate688(.a(gate462inter0), .b(s_20), .O(gate462inter1));
  and2  gate689(.a(G1195), .b(G1099), .O(gate462inter2));
  inv1  gate690(.a(s_20), .O(gate462inter3));
  inv1  gate691(.a(s_21), .O(gate462inter4));
  nand2 gate692(.a(gate462inter4), .b(gate462inter3), .O(gate462inter5));
  nor2  gate693(.a(gate462inter5), .b(gate462inter2), .O(gate462inter6));
  inv1  gate694(.a(G1099), .O(gate462inter7));
  inv1  gate695(.a(G1195), .O(gate462inter8));
  nand2 gate696(.a(gate462inter8), .b(gate462inter7), .O(gate462inter9));
  nand2 gate697(.a(s_21), .b(gate462inter3), .O(gate462inter10));
  nor2  gate698(.a(gate462inter10), .b(gate462inter9), .O(gate462inter11));
  nor2  gate699(.a(gate462inter11), .b(gate462inter6), .O(gate462inter12));
  nand2 gate700(.a(gate462inter12), .b(gate462inter1), .O(G1271));
nand2 gate463( .a(G23), .b(G1198), .O(G1272) );
nand2 gate464( .a(G1102), .b(G1198), .O(G1273) );
nand2 gate465( .a(G24), .b(G1201), .O(G1274) );
nand2 gate466( .a(G1105), .b(G1201), .O(G1275) );
nand2 gate467( .a(G25), .b(G1204), .O(G1276) );
nand2 gate468( .a(G1108), .b(G1204), .O(G1277) );
nand2 gate469( .a(G26), .b(G1207), .O(G1278) );

  xor2  gate1093(.a(G1207), .b(G1111), .O(gate470inter0));
  nand2 gate1094(.a(gate470inter0), .b(s_78), .O(gate470inter1));
  and2  gate1095(.a(G1207), .b(G1111), .O(gate470inter2));
  inv1  gate1096(.a(s_78), .O(gate470inter3));
  inv1  gate1097(.a(s_79), .O(gate470inter4));
  nand2 gate1098(.a(gate470inter4), .b(gate470inter3), .O(gate470inter5));
  nor2  gate1099(.a(gate470inter5), .b(gate470inter2), .O(gate470inter6));
  inv1  gate1100(.a(G1111), .O(gate470inter7));
  inv1  gate1101(.a(G1207), .O(gate470inter8));
  nand2 gate1102(.a(gate470inter8), .b(gate470inter7), .O(gate470inter9));
  nand2 gate1103(.a(s_79), .b(gate470inter3), .O(gate470inter10));
  nor2  gate1104(.a(gate470inter10), .b(gate470inter9), .O(gate470inter11));
  nor2  gate1105(.a(gate470inter11), .b(gate470inter6), .O(gate470inter12));
  nand2 gate1106(.a(gate470inter12), .b(gate470inter1), .O(G1279));
nand2 gate471( .a(G27), .b(G1210), .O(G1280) );
nand2 gate472( .a(G1114), .b(G1210), .O(G1281) );
nand2 gate473( .a(G28), .b(G1213), .O(G1282) );
nand2 gate474( .a(G1117), .b(G1213), .O(G1283) );
nand2 gate475( .a(G29), .b(G1216), .O(G1284) );
nand2 gate476( .a(G1120), .b(G1216), .O(G1285) );
nand2 gate477( .a(G30), .b(G1219), .O(G1286) );
nand2 gate478( .a(G1123), .b(G1219), .O(G1287) );

  xor2  gate771(.a(G1222), .b(G31), .O(gate479inter0));
  nand2 gate772(.a(gate479inter0), .b(s_32), .O(gate479inter1));
  and2  gate773(.a(G1222), .b(G31), .O(gate479inter2));
  inv1  gate774(.a(s_32), .O(gate479inter3));
  inv1  gate775(.a(s_33), .O(gate479inter4));
  nand2 gate776(.a(gate479inter4), .b(gate479inter3), .O(gate479inter5));
  nor2  gate777(.a(gate479inter5), .b(gate479inter2), .O(gate479inter6));
  inv1  gate778(.a(G31), .O(gate479inter7));
  inv1  gate779(.a(G1222), .O(gate479inter8));
  nand2 gate780(.a(gate479inter8), .b(gate479inter7), .O(gate479inter9));
  nand2 gate781(.a(s_33), .b(gate479inter3), .O(gate479inter10));
  nor2  gate782(.a(gate479inter10), .b(gate479inter9), .O(gate479inter11));
  nor2  gate783(.a(gate479inter11), .b(gate479inter6), .O(gate479inter12));
  nand2 gate784(.a(gate479inter12), .b(gate479inter1), .O(G1288));
nand2 gate480( .a(G1126), .b(G1222), .O(G1289) );
nand2 gate481( .a(G32), .b(G1225), .O(G1290) );
nand2 gate482( .a(G1129), .b(G1225), .O(G1291) );
nand2 gate483( .a(G1228), .b(G1229), .O(G1292) );
nand2 gate484( .a(G1230), .b(G1231), .O(G1293) );
nand2 gate485( .a(G1232), .b(G1233), .O(G1294) );
nand2 gate486( .a(G1234), .b(G1235), .O(G1295) );
nand2 gate487( .a(G1236), .b(G1237), .O(G1296) );
nand2 gate488( .a(G1238), .b(G1239), .O(G1297) );
nand2 gate489( .a(G1240), .b(G1241), .O(G1298) );
nand2 gate490( .a(G1242), .b(G1243), .O(G1299) );
nand2 gate491( .a(G1244), .b(G1245), .O(G1300) );
nand2 gate492( .a(G1246), .b(G1247), .O(G1301) );
nand2 gate493( .a(G1248), .b(G1249), .O(G1302) );
nand2 gate494( .a(G1250), .b(G1251), .O(G1303) );

  xor2  gate1121(.a(G1253), .b(G1252), .O(gate495inter0));
  nand2 gate1122(.a(gate495inter0), .b(s_82), .O(gate495inter1));
  and2  gate1123(.a(G1253), .b(G1252), .O(gate495inter2));
  inv1  gate1124(.a(s_82), .O(gate495inter3));
  inv1  gate1125(.a(s_83), .O(gate495inter4));
  nand2 gate1126(.a(gate495inter4), .b(gate495inter3), .O(gate495inter5));
  nor2  gate1127(.a(gate495inter5), .b(gate495inter2), .O(gate495inter6));
  inv1  gate1128(.a(G1252), .O(gate495inter7));
  inv1  gate1129(.a(G1253), .O(gate495inter8));
  nand2 gate1130(.a(gate495inter8), .b(gate495inter7), .O(gate495inter9));
  nand2 gate1131(.a(s_83), .b(gate495inter3), .O(gate495inter10));
  nor2  gate1132(.a(gate495inter10), .b(gate495inter9), .O(gate495inter11));
  nor2  gate1133(.a(gate495inter11), .b(gate495inter6), .O(gate495inter12));
  nand2 gate1134(.a(gate495inter12), .b(gate495inter1), .O(G1304));
nand2 gate496( .a(G1254), .b(G1255), .O(G1305) );
nand2 gate497( .a(G1256), .b(G1257), .O(G1306) );
nand2 gate498( .a(G1258), .b(G1259), .O(G1307) );
nand2 gate499( .a(G1260), .b(G1261), .O(G1308) );
nand2 gate500( .a(G1262), .b(G1263), .O(G1309) );

  xor2  gate813(.a(G1265), .b(G1264), .O(gate501inter0));
  nand2 gate814(.a(gate501inter0), .b(s_38), .O(gate501inter1));
  and2  gate815(.a(G1265), .b(G1264), .O(gate501inter2));
  inv1  gate816(.a(s_38), .O(gate501inter3));
  inv1  gate817(.a(s_39), .O(gate501inter4));
  nand2 gate818(.a(gate501inter4), .b(gate501inter3), .O(gate501inter5));
  nor2  gate819(.a(gate501inter5), .b(gate501inter2), .O(gate501inter6));
  inv1  gate820(.a(G1264), .O(gate501inter7));
  inv1  gate821(.a(G1265), .O(gate501inter8));
  nand2 gate822(.a(gate501inter8), .b(gate501inter7), .O(gate501inter9));
  nand2 gate823(.a(s_39), .b(gate501inter3), .O(gate501inter10));
  nor2  gate824(.a(gate501inter10), .b(gate501inter9), .O(gate501inter11));
  nor2  gate825(.a(gate501inter11), .b(gate501inter6), .O(gate501inter12));
  nand2 gate826(.a(gate501inter12), .b(gate501inter1), .O(G1310));
nand2 gate502( .a(G1266), .b(G1267), .O(G1311) );
nand2 gate503( .a(G1268), .b(G1269), .O(G1312) );
nand2 gate504( .a(G1270), .b(G1271), .O(G1313) );
nand2 gate505( .a(G1272), .b(G1273), .O(G1314) );
nand2 gate506( .a(G1274), .b(G1275), .O(G1315) );
nand2 gate507( .a(G1276), .b(G1277), .O(G1316) );

  xor2  gate1135(.a(G1279), .b(G1278), .O(gate508inter0));
  nand2 gate1136(.a(gate508inter0), .b(s_84), .O(gate508inter1));
  and2  gate1137(.a(G1279), .b(G1278), .O(gate508inter2));
  inv1  gate1138(.a(s_84), .O(gate508inter3));
  inv1  gate1139(.a(s_85), .O(gate508inter4));
  nand2 gate1140(.a(gate508inter4), .b(gate508inter3), .O(gate508inter5));
  nor2  gate1141(.a(gate508inter5), .b(gate508inter2), .O(gate508inter6));
  inv1  gate1142(.a(G1278), .O(gate508inter7));
  inv1  gate1143(.a(G1279), .O(gate508inter8));
  nand2 gate1144(.a(gate508inter8), .b(gate508inter7), .O(gate508inter9));
  nand2 gate1145(.a(s_85), .b(gate508inter3), .O(gate508inter10));
  nor2  gate1146(.a(gate508inter10), .b(gate508inter9), .O(gate508inter11));
  nor2  gate1147(.a(gate508inter11), .b(gate508inter6), .O(gate508inter12));
  nand2 gate1148(.a(gate508inter12), .b(gate508inter1), .O(G1317));
nand2 gate509( .a(G1280), .b(G1281), .O(G1318) );

  xor2  gate1079(.a(G1283), .b(G1282), .O(gate510inter0));
  nand2 gate1080(.a(gate510inter0), .b(s_76), .O(gate510inter1));
  and2  gate1081(.a(G1283), .b(G1282), .O(gate510inter2));
  inv1  gate1082(.a(s_76), .O(gate510inter3));
  inv1  gate1083(.a(s_77), .O(gate510inter4));
  nand2 gate1084(.a(gate510inter4), .b(gate510inter3), .O(gate510inter5));
  nor2  gate1085(.a(gate510inter5), .b(gate510inter2), .O(gate510inter6));
  inv1  gate1086(.a(G1282), .O(gate510inter7));
  inv1  gate1087(.a(G1283), .O(gate510inter8));
  nand2 gate1088(.a(gate510inter8), .b(gate510inter7), .O(gate510inter9));
  nand2 gate1089(.a(s_77), .b(gate510inter3), .O(gate510inter10));
  nor2  gate1090(.a(gate510inter10), .b(gate510inter9), .O(gate510inter11));
  nor2  gate1091(.a(gate510inter11), .b(gate510inter6), .O(gate510inter12));
  nand2 gate1092(.a(gate510inter12), .b(gate510inter1), .O(G1319));
nand2 gate511( .a(G1284), .b(G1285), .O(G1320) );
nand2 gate512( .a(G1286), .b(G1287), .O(G1321) );
nand2 gate513( .a(G1288), .b(G1289), .O(G1322) );

  xor2  gate981(.a(G1291), .b(G1290), .O(gate514inter0));
  nand2 gate982(.a(gate514inter0), .b(s_62), .O(gate514inter1));
  and2  gate983(.a(G1291), .b(G1290), .O(gate514inter2));
  inv1  gate984(.a(s_62), .O(gate514inter3));
  inv1  gate985(.a(s_63), .O(gate514inter4));
  nand2 gate986(.a(gate514inter4), .b(gate514inter3), .O(gate514inter5));
  nor2  gate987(.a(gate514inter5), .b(gate514inter2), .O(gate514inter6));
  inv1  gate988(.a(G1290), .O(gate514inter7));
  inv1  gate989(.a(G1291), .O(gate514inter8));
  nand2 gate990(.a(gate514inter8), .b(gate514inter7), .O(gate514inter9));
  nand2 gate991(.a(s_63), .b(gate514inter3), .O(gate514inter10));
  nor2  gate992(.a(gate514inter10), .b(gate514inter9), .O(gate514inter11));
  nor2  gate993(.a(gate514inter11), .b(gate514inter6), .O(gate514inter12));
  nand2 gate994(.a(gate514inter12), .b(gate514inter1), .O(G1323));
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule