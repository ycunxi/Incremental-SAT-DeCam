module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);

input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;//RE__PI;

input s_0,s_1;//RE__ALLOW(00,01,10,11);
input s_2,s_3;//RE__ALLOW(00,01,10,11);
input s_4,s_5;//RE__ALLOW(00,01,10,11);
input s_6,s_7;//RE__ALLOW(00,01,10,11);
input s_8,s_9;//RE__ALLOW(00,01,10,11);
input s_10,s_11;//RE__ALLOW(00,01,10,11);
input s_12,s_13;//RE__ALLOW(00,01,10,11);
input s_14,s_15;//RE__ALLOW(00,01,10,11);
input s_16,s_17;//RE__ALLOW(00,01,10,11);
input s_18,s_19;//RE__ALLOW(00,01,10,11);
input s_20,s_21;//RE__ALLOW(00,01,10,11);
input s_22,s_23;//RE__ALLOW(00,01,10,11);
input s_24,s_25;//RE__ALLOW(00,01,10,11);
input s_26,s_27;//RE__ALLOW(00,01,10,11);
input s_28,s_29;//RE__ALLOW(00,01,10,11);
input s_30,s_31;//RE__ALLOW(00,01,10,11);
input s_32,s_33;//RE__ALLOW(00,01,10,11);
input s_34,s_35;//RE__ALLOW(00,01,10,11);
input s_36,s_37;//RE__ALLOW(00,01,10,11);
input s_38,s_39;//RE__ALLOW(00,01,10,11);
input s_40,s_41;//RE__ALLOW(00,01,10,11);
input s_42,s_43;//RE__ALLOW(00,01,10,11);
input s_44,s_45;//RE__ALLOW(00,01,10,11);
input s_46,s_47;//RE__ALLOW(00,01,10,11);
input s_48,s_49;//RE__ALLOW(00,01,10,11);
input s_50,s_51;//RE__ALLOW(00,01,10,11);
input s_52,s_53;//RE__ALLOW(00,01,10,11);
input s_54,s_55;//RE__ALLOW(00,01,10,11);
input s_56,s_57;//RE__ALLOW(00,01,10,11);
input s_58,s_59;//RE__ALLOW(00,01,10,11);
input s_60,s_61;//RE__ALLOW(00,01,10,11);
input s_62,s_63;//RE__ALLOW(00,01,10,11);
input s_64,s_65;//RE__ALLOW(00,01,10,11);
input s_66,s_67;//RE__ALLOW(00,01,10,11);
input s_68,s_69;//RE__ALLOW(00,01,10,11);
input s_70,s_71;//RE__ALLOW(00,01,10,11);
input s_72,s_73;//RE__ALLOW(00,01,10,11);
input s_74,s_75;//RE__ALLOW(00,01,10,11);
input s_76,s_77;//RE__ALLOW(00,01,10,11);
input s_78,s_79;//RE__ALLOW(00,01,10,11);
input s_80,s_81;//RE__ALLOW(00,01,10,11);
input s_82,s_83;//RE__ALLOW(00,01,10,11);
input s_84,s_85;//RE__ALLOW(00,01,10,11);
input s_86,s_87;//RE__ALLOW(00,01,10,11);
input s_88,s_89;//RE__ALLOW(00,01,10,11);
input s_90,s_91;//RE__ALLOW(00,01,10,11);
input s_92,s_93;//RE__ALLOW(00,01,10,11);
input s_94,s_95;//RE__ALLOW(00,01,10,11);
input s_96,s_97;//RE__ALLOW(00,01,10,11);
input s_98,s_99;//RE__ALLOW(00,01,10,11);
input s_100,s_101;//RE__ALLOW(00,01,10,11);
input s_102,s_103;//RE__ALLOW(00,01,10,11);
input s_104,s_105;//RE__ALLOW(00,01,10,11);
input s_106,s_107;//RE__ALLOW(00,01,10,11);
input s_108,s_109;//RE__ALLOW(00,01,10,11);
input s_110,s_111;//RE__ALLOW(00,01,10,11);
input s_112,s_113;//RE__ALLOW(00,01,10,11);
input s_114,s_115;//RE__ALLOW(00,01,10,11);
input s_116,s_117;//RE__ALLOW(00,01,10,11);
input s_118,s_119;//RE__ALLOW(00,01,10,11);
input s_120,s_121;//RE__ALLOW(00,01,10,11);
input s_122,s_123;//RE__ALLOW(00,01,10,11);
input s_124,s_125;//RE__ALLOW(00,01,10,11);
input s_126,s_127;//RE__ALLOW(00,01,10,11);
input s_128,s_129;//RE__ALLOW(00,01,10,11);
input s_130,s_131;//RE__ALLOW(00,01,10,11);
input s_132,s_133;//RE__ALLOW(00,01,10,11);
input s_134,s_135;//RE__ALLOW(00,01,10,11);
input s_136,s_137;//RE__ALLOW(00,01,10,11);
input s_138,s_139;//RE__ALLOW(00,01,10,11);
input s_140,s_141;//RE__ALLOW(00,01,10,11);
input s_142,s_143;//RE__ALLOW(00,01,10,11);
input s_144,s_145;//RE__ALLOW(00,01,10,11);
input s_146,s_147;//RE__ALLOW(00,01,10,11);
input s_148,s_149;//RE__ALLOW(00,01,10,11);
input s_150,s_151;//RE__ALLOW(00,01,10,11);
input s_152,s_153;//RE__ALLOW(00,01,10,11);
input s_154,s_155;//RE__ALLOW(00,01,10,11);
input s_156,s_157;//RE__ALLOW(00,01,10,11);
input s_158,s_159;//RE__ALLOW(00,01,10,11);
input s_160,s_161;//RE__ALLOW(00,01,10,11);
input s_162,s_163;//RE__ALLOW(00,01,10,11);
input s_164,s_165;//RE__ALLOW(00,01,10,11);
input s_166,s_167;//RE__ALLOW(00,01,10,11);
input s_168,s_169;//RE__ALLOW(00,01,10,11);
input s_170,s_171;//RE__ALLOW(00,01,10,11);
input s_172,s_173;//RE__ALLOW(00,01,10,11);
input s_174,s_175;//RE__ALLOW(00,01,10,11);
input s_176,s_177;//RE__ALLOW(00,01,10,11);
input s_178,s_179;//RE__ALLOW(00,01,10,11);
input s_180,s_181;//RE__ALLOW(00,01,10,11);
input s_182,s_183;//RE__ALLOW(00,01,10,11);
input s_184,s_185;//RE__ALLOW(00,01,10,11);
input s_186,s_187;//RE__ALLOW(00,01,10,11);
input s_188,s_189;//RE__ALLOW(00,01,10,11);
input s_190,s_191;//RE__ALLOW(00,01,10,11);
input s_192,s_193;//RE__ALLOW(00,01,10,11);
input s_194,s_195;//RE__ALLOW(00,01,10,11);
input s_196,s_197;//RE__ALLOW(00,01,10,11);
input s_198,s_199;//RE__ALLOW(00,01,10,11);
input s_200,s_201;//RE__ALLOW(00,01,10,11);
input s_202,s_203;//RE__ALLOW(00,01,10,11);
input s_204,s_205;//RE__ALLOW(00,01,10,11);
input s_206,s_207;//RE__ALLOW(00,01,10,11);
input s_208,s_209;//RE__ALLOW(00,01,10,11);
input s_210,s_211;//RE__ALLOW(00,01,10,11);
input s_212,s_213;//RE__ALLOW(00,01,10,11);
input s_214,s_215;//RE__ALLOW(00,01,10,11);
input s_216,s_217;//RE__ALLOW(00,01,10,11);
input s_218,s_219;//RE__ALLOW(00,01,10,11);
input s_220,s_221;//RE__ALLOW(00,01,10,11);
input s_222,s_223;//RE__ALLOW(00,01,10,11);
input s_224,s_225;//RE__ALLOW(00,01,10,11);
input s_226,s_227;//RE__ALLOW(00,01,10,11);
input s_228,s_229;//RE__ALLOW(00,01,10,11);
input s_230,s_231;//RE__ALLOW(00,01,10,11);
input s_232,s_233;//RE__ALLOW(00,01,10,11);
input s_234,s_235;//RE__ALLOW(00,01,10,11);
input s_236,s_237;//RE__ALLOW(00,01,10,11);
input s_238,s_239;//RE__ALLOW(00,01,10,11);
input s_240,s_241;//RE__ALLOW(00,01,10,11);
input s_242,s_243;//RE__ALLOW(00,01,10,11);
input s_244,s_245;//RE__ALLOW(00,01,10,11);
input s_246,s_247;//RE__ALLOW(00,01,10,11);
input s_248,s_249;//RE__ALLOW(00,01,10,11);
input s_250,s_251;//RE__ALLOW(00,01,10,11);
input s_252,s_253;//RE__ALLOW(00,01,10,11);
input s_254,s_255;//RE__ALLOW(00,01,10,11);
input s_256,s_257;//RE__ALLOW(00,01,10,11);
input s_258,s_259;//RE__ALLOW(00,01,10,11);
input s_260,s_261;//RE__ALLOW(00,01,10,11);
input s_262,s_263;//RE__ALLOW(00,01,10,11);
input s_264,s_265;//RE__ALLOW(00,01,10,11);
input s_266,s_267;//RE__ALLOW(00,01,10,11);
input s_268,s_269;//RE__ALLOW(00,01,10,11);
input s_270,s_271;//RE__ALLOW(00,01,10,11);
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;

  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate453inter0, gate453inter1, gate453inter2, gate453inter3, gate453inter4, gate453inter5, gate453inter6, gate453inter7, gate453inter8, gate453inter9, gate453inter10, gate453inter11, gate453inter12, gate46inter0, gate46inter1, gate46inter2, gate46inter3, gate46inter4, gate46inter5, gate46inter6, gate46inter7, gate46inter8, gate46inter9, gate46inter10, gate46inter11, gate46inter12, gate78inter0, gate78inter1, gate78inter2, gate78inter3, gate78inter4, gate78inter5, gate78inter6, gate78inter7, gate78inter8, gate78inter9, gate78inter10, gate78inter11, gate78inter12, gate28inter0, gate28inter1, gate28inter2, gate28inter3, gate28inter4, gate28inter5, gate28inter6, gate28inter7, gate28inter8, gate28inter9, gate28inter10, gate28inter11, gate28inter12, gate228inter0, gate228inter1, gate228inter2, gate228inter3, gate228inter4, gate228inter5, gate228inter6, gate228inter7, gate228inter8, gate228inter9, gate228inter10, gate228inter11, gate228inter12, gate264inter0, gate264inter1, gate264inter2, gate264inter3, gate264inter4, gate264inter5, gate264inter6, gate264inter7, gate264inter8, gate264inter9, gate264inter10, gate264inter11, gate264inter12, gate147inter0, gate147inter1, gate147inter2, gate147inter3, gate147inter4, gate147inter5, gate147inter6, gate147inter7, gate147inter8, gate147inter9, gate147inter10, gate147inter11, gate147inter12, gate257inter0, gate257inter1, gate257inter2, gate257inter3, gate257inter4, gate257inter5, gate257inter6, gate257inter7, gate257inter8, gate257inter9, gate257inter10, gate257inter11, gate257inter12, gate490inter0, gate490inter1, gate490inter2, gate490inter3, gate490inter4, gate490inter5, gate490inter6, gate490inter7, gate490inter8, gate490inter9, gate490inter10, gate490inter11, gate490inter12, gate184inter0, gate184inter1, gate184inter2, gate184inter3, gate184inter4, gate184inter5, gate184inter6, gate184inter7, gate184inter8, gate184inter9, gate184inter10, gate184inter11, gate184inter12, gate77inter0, gate77inter1, gate77inter2, gate77inter3, gate77inter4, gate77inter5, gate77inter6, gate77inter7, gate77inter8, gate77inter9, gate77inter10, gate77inter11, gate77inter12, gate286inter0, gate286inter1, gate286inter2, gate286inter3, gate286inter4, gate286inter5, gate286inter6, gate286inter7, gate286inter8, gate286inter9, gate286inter10, gate286inter11, gate286inter12, gate278inter0, gate278inter1, gate278inter2, gate278inter3, gate278inter4, gate278inter5, gate278inter6, gate278inter7, gate278inter8, gate278inter9, gate278inter10, gate278inter11, gate278inter12, gate389inter0, gate389inter1, gate389inter2, gate389inter3, gate389inter4, gate389inter5, gate389inter6, gate389inter7, gate389inter8, gate389inter9, gate389inter10, gate389inter11, gate389inter12, gate112inter0, gate112inter1, gate112inter2, gate112inter3, gate112inter4, gate112inter5, gate112inter6, gate112inter7, gate112inter8, gate112inter9, gate112inter10, gate112inter11, gate112inter12, gate37inter0, gate37inter1, gate37inter2, gate37inter3, gate37inter4, gate37inter5, gate37inter6, gate37inter7, gate37inter8, gate37inter9, gate37inter10, gate37inter11, gate37inter12, gate135inter0, gate135inter1, gate135inter2, gate135inter3, gate135inter4, gate135inter5, gate135inter6, gate135inter7, gate135inter8, gate135inter9, gate135inter10, gate135inter11, gate135inter12, gate477inter0, gate477inter1, gate477inter2, gate477inter3, gate477inter4, gate477inter5, gate477inter6, gate477inter7, gate477inter8, gate477inter9, gate477inter10, gate477inter11, gate477inter12, gate89inter0, gate89inter1, gate89inter2, gate89inter3, gate89inter4, gate89inter5, gate89inter6, gate89inter7, gate89inter8, gate89inter9, gate89inter10, gate89inter11, gate89inter12, gate439inter0, gate439inter1, gate439inter2, gate439inter3, gate439inter4, gate439inter5, gate439inter6, gate439inter7, gate439inter8, gate439inter9, gate439inter10, gate439inter11, gate439inter12, gate416inter0, gate416inter1, gate416inter2, gate416inter3, gate416inter4, gate416inter5, gate416inter6, gate416inter7, gate416inter8, gate416inter9, gate416inter10, gate416inter11, gate416inter12, gate181inter0, gate181inter1, gate181inter2, gate181inter3, gate181inter4, gate181inter5, gate181inter6, gate181inter7, gate181inter8, gate181inter9, gate181inter10, gate181inter11, gate181inter12, gate397inter0, gate397inter1, gate397inter2, gate397inter3, gate397inter4, gate397inter5, gate397inter6, gate397inter7, gate397inter8, gate397inter9, gate397inter10, gate397inter11, gate397inter12, gate215inter0, gate215inter1, gate215inter2, gate215inter3, gate215inter4, gate215inter5, gate215inter6, gate215inter7, gate215inter8, gate215inter9, gate215inter10, gate215inter11, gate215inter12, gate101inter0, gate101inter1, gate101inter2, gate101inter3, gate101inter4, gate101inter5, gate101inter6, gate101inter7, gate101inter8, gate101inter9, gate101inter10, gate101inter11, gate101inter12, gate55inter0, gate55inter1, gate55inter2, gate55inter3, gate55inter4, gate55inter5, gate55inter6, gate55inter7, gate55inter8, gate55inter9, gate55inter10, gate55inter11, gate55inter12, gate458inter0, gate458inter1, gate458inter2, gate458inter3, gate458inter4, gate458inter5, gate458inter6, gate458inter7, gate458inter8, gate458inter9, gate458inter10, gate458inter11, gate458inter12, gate473inter0, gate473inter1, gate473inter2, gate473inter3, gate473inter4, gate473inter5, gate473inter6, gate473inter7, gate473inter8, gate473inter9, gate473inter10, gate473inter11, gate473inter12, gate440inter0, gate440inter1, gate440inter2, gate440inter3, gate440inter4, gate440inter5, gate440inter6, gate440inter7, gate440inter8, gate440inter9, gate440inter10, gate440inter11, gate440inter12, gate203inter0, gate203inter1, gate203inter2, gate203inter3, gate203inter4, gate203inter5, gate203inter6, gate203inter7, gate203inter8, gate203inter9, gate203inter10, gate203inter11, gate203inter12, gate258inter0, gate258inter1, gate258inter2, gate258inter3, gate258inter4, gate258inter5, gate258inter6, gate258inter7, gate258inter8, gate258inter9, gate258inter10, gate258inter11, gate258inter12, gate162inter0, gate162inter1, gate162inter2, gate162inter3, gate162inter4, gate162inter5, gate162inter6, gate162inter7, gate162inter8, gate162inter9, gate162inter10, gate162inter11, gate162inter12, gate294inter0, gate294inter1, gate294inter2, gate294inter3, gate294inter4, gate294inter5, gate294inter6, gate294inter7, gate294inter8, gate294inter9, gate294inter10, gate294inter11, gate294inter12, gate288inter0, gate288inter1, gate288inter2, gate288inter3, gate288inter4, gate288inter5, gate288inter6, gate288inter7, gate288inter8, gate288inter9, gate288inter10, gate288inter11, gate288inter12, gate237inter0, gate237inter1, gate237inter2, gate237inter3, gate237inter4, gate237inter5, gate237inter6, gate237inter7, gate237inter8, gate237inter9, gate237inter10, gate237inter11, gate237inter12, gate43inter0, gate43inter1, gate43inter2, gate43inter3, gate43inter4, gate43inter5, gate43inter6, gate43inter7, gate43inter8, gate43inter9, gate43inter10, gate43inter11, gate43inter12, gate472inter0, gate472inter1, gate472inter2, gate472inter3, gate472inter4, gate472inter5, gate472inter6, gate472inter7, gate472inter8, gate472inter9, gate472inter10, gate472inter11, gate472inter12, gate498inter0, gate498inter1, gate498inter2, gate498inter3, gate498inter4, gate498inter5, gate498inter6, gate498inter7, gate498inter8, gate498inter9, gate498inter10, gate498inter11, gate498inter12, gate276inter0, gate276inter1, gate276inter2, gate276inter3, gate276inter4, gate276inter5, gate276inter6, gate276inter7, gate276inter8, gate276inter9, gate276inter10, gate276inter11, gate276inter12, gate200inter0, gate200inter1, gate200inter2, gate200inter3, gate200inter4, gate200inter5, gate200inter6, gate200inter7, gate200inter8, gate200inter9, gate200inter10, gate200inter11, gate200inter12, gate510inter0, gate510inter1, gate510inter2, gate510inter3, gate510inter4, gate510inter5, gate510inter6, gate510inter7, gate510inter8, gate510inter9, gate510inter10, gate510inter11, gate510inter12, gate399inter0, gate399inter1, gate399inter2, gate399inter3, gate399inter4, gate399inter5, gate399inter6, gate399inter7, gate399inter8, gate399inter9, gate399inter10, gate399inter11, gate399inter12, gate507inter0, gate507inter1, gate507inter2, gate507inter3, gate507inter4, gate507inter5, gate507inter6, gate507inter7, gate507inter8, gate507inter9, gate507inter10, gate507inter11, gate507inter12, gate156inter0, gate156inter1, gate156inter2, gate156inter3, gate156inter4, gate156inter5, gate156inter6, gate156inter7, gate156inter8, gate156inter9, gate156inter10, gate156inter11, gate156inter12, gate98inter0, gate98inter1, gate98inter2, gate98inter3, gate98inter4, gate98inter5, gate98inter6, gate98inter7, gate98inter8, gate98inter9, gate98inter10, gate98inter11, gate98inter12, gate277inter0, gate277inter1, gate277inter2, gate277inter3, gate277inter4, gate277inter5, gate277inter6, gate277inter7, gate277inter8, gate277inter9, gate277inter10, gate277inter11, gate277inter12, gate82inter0, gate82inter1, gate82inter2, gate82inter3, gate82inter4, gate82inter5, gate82inter6, gate82inter7, gate82inter8, gate82inter9, gate82inter10, gate82inter11, gate82inter12, gate110inter0, gate110inter1, gate110inter2, gate110inter3, gate110inter4, gate110inter5, gate110inter6, gate110inter7, gate110inter8, gate110inter9, gate110inter10, gate110inter11, gate110inter12, gate103inter0, gate103inter1, gate103inter2, gate103inter3, gate103inter4, gate103inter5, gate103inter6, gate103inter7, gate103inter8, gate103inter9, gate103inter10, gate103inter11, gate103inter12, gate259inter0, gate259inter1, gate259inter2, gate259inter3, gate259inter4, gate259inter5, gate259inter6, gate259inter7, gate259inter8, gate259inter9, gate259inter10, gate259inter11, gate259inter12, gate480inter0, gate480inter1, gate480inter2, gate480inter3, gate480inter4, gate480inter5, gate480inter6, gate480inter7, gate480inter8, gate480inter9, gate480inter10, gate480inter11, gate480inter12, gate459inter0, gate459inter1, gate459inter2, gate459inter3, gate459inter4, gate459inter5, gate459inter6, gate459inter7, gate459inter8, gate459inter9, gate459inter10, gate459inter11, gate459inter12, gate30inter0, gate30inter1, gate30inter2, gate30inter3, gate30inter4, gate30inter5, gate30inter6, gate30inter7, gate30inter8, gate30inter9, gate30inter10, gate30inter11, gate30inter12, gate92inter0, gate92inter1, gate92inter2, gate92inter3, gate92inter4, gate92inter5, gate92inter6, gate92inter7, gate92inter8, gate92inter9, gate92inter10, gate92inter11, gate92inter12, gate482inter0, gate482inter1, gate482inter2, gate482inter3, gate482inter4, gate482inter5, gate482inter6, gate482inter7, gate482inter8, gate482inter9, gate482inter10, gate482inter11, gate482inter12, gate79inter0, gate79inter1, gate79inter2, gate79inter3, gate79inter4, gate79inter5, gate79inter6, gate79inter7, gate79inter8, gate79inter9, gate79inter10, gate79inter11, gate79inter12, gate206inter0, gate206inter1, gate206inter2, gate206inter3, gate206inter4, gate206inter5, gate206inter6, gate206inter7, gate206inter8, gate206inter9, gate206inter10, gate206inter11, gate206inter12, gate9inter0, gate9inter1, gate9inter2, gate9inter3, gate9inter4, gate9inter5, gate9inter6, gate9inter7, gate9inter8, gate9inter9, gate9inter10, gate9inter11, gate9inter12, gate478inter0, gate478inter1, gate478inter2, gate478inter3, gate478inter4, gate478inter5, gate478inter6, gate478inter7, gate478inter8, gate478inter9, gate478inter10, gate478inter11, gate478inter12, gate219inter0, gate219inter1, gate219inter2, gate219inter3, gate219inter4, gate219inter5, gate219inter6, gate219inter7, gate219inter8, gate219inter9, gate219inter10, gate219inter11, gate219inter12, gate422inter0, gate422inter1, gate422inter2, gate422inter3, gate422inter4, gate422inter5, gate422inter6, gate422inter7, gate422inter8, gate422inter9, gate422inter10, gate422inter11, gate422inter12, gate81inter0, gate81inter1, gate81inter2, gate81inter3, gate81inter4, gate81inter5, gate81inter6, gate81inter7, gate81inter8, gate81inter9, gate81inter10, gate81inter11, gate81inter12, gate171inter0, gate171inter1, gate171inter2, gate171inter3, gate171inter4, gate171inter5, gate171inter6, gate171inter7, gate171inter8, gate171inter9, gate171inter10, gate171inter11, gate171inter12, gate86inter0, gate86inter1, gate86inter2, gate86inter3, gate86inter4, gate86inter5, gate86inter6, gate86inter7, gate86inter8, gate86inter9, gate86inter10, gate86inter11, gate86inter12, gate113inter0, gate113inter1, gate113inter2, gate113inter3, gate113inter4, gate113inter5, gate113inter6, gate113inter7, gate113inter8, gate113inter9, gate113inter10, gate113inter11, gate113inter12, gate495inter0, gate495inter1, gate495inter2, gate495inter3, gate495inter4, gate495inter5, gate495inter6, gate495inter7, gate495inter8, gate495inter9, gate495inter10, gate495inter11, gate495inter12, gate239inter0, gate239inter1, gate239inter2, gate239inter3, gate239inter4, gate239inter5, gate239inter6, gate239inter7, gate239inter8, gate239inter9, gate239inter10, gate239inter11, gate239inter12, gate233inter0, gate233inter1, gate233inter2, gate233inter3, gate233inter4, gate233inter5, gate233inter6, gate233inter7, gate233inter8, gate233inter9, gate233inter10, gate233inter11, gate233inter12, gate186inter0, gate186inter1, gate186inter2, gate186inter3, gate186inter4, gate186inter5, gate186inter6, gate186inter7, gate186inter8, gate186inter9, gate186inter10, gate186inter11, gate186inter12, gate102inter0, gate102inter1, gate102inter2, gate102inter3, gate102inter4, gate102inter5, gate102inter6, gate102inter7, gate102inter8, gate102inter9, gate102inter10, gate102inter11, gate102inter12, gate467inter0, gate467inter1, gate467inter2, gate467inter3, gate467inter4, gate467inter5, gate467inter6, gate467inter7, gate467inter8, gate467inter9, gate467inter10, gate467inter11, gate467inter12, gate388inter0, gate388inter1, gate388inter2, gate388inter3, gate388inter4, gate388inter5, gate388inter6, gate388inter7, gate388inter8, gate388inter9, gate388inter10, gate388inter11, gate388inter12, gate244inter0, gate244inter1, gate244inter2, gate244inter3, gate244inter4, gate244inter5, gate244inter6, gate244inter7, gate244inter8, gate244inter9, gate244inter10, gate244inter11, gate244inter12, gate65inter0, gate65inter1, gate65inter2, gate65inter3, gate65inter4, gate65inter5, gate65inter6, gate65inter7, gate65inter8, gate65inter9, gate65inter10, gate65inter11, gate65inter12, gate35inter0, gate35inter1, gate35inter2, gate35inter3, gate35inter4, gate35inter5, gate35inter6, gate35inter7, gate35inter8, gate35inter9, gate35inter10, gate35inter11, gate35inter12, gate427inter0, gate427inter1, gate427inter2, gate427inter3, gate427inter4, gate427inter5, gate427inter6, gate427inter7, gate427inter8, gate427inter9, gate427inter10, gate427inter11, gate427inter12, gate107inter0, gate107inter1, gate107inter2, gate107inter3, gate107inter4, gate107inter5, gate107inter6, gate107inter7, gate107inter8, gate107inter9, gate107inter10, gate107inter11, gate107inter12, gate514inter0, gate514inter1, gate514inter2, gate514inter3, gate514inter4, gate514inter5, gate514inter6, gate514inter7, gate514inter8, gate514inter9, gate514inter10, gate514inter11, gate514inter12, gate132inter0, gate132inter1, gate132inter2, gate132inter3, gate132inter4, gate132inter5, gate132inter6, gate132inter7, gate132inter8, gate132inter9, gate132inter10, gate132inter11, gate132inter12, gate447inter0, gate447inter1, gate447inter2, gate447inter3, gate447inter4, gate447inter5, gate447inter6, gate447inter7, gate447inter8, gate447inter9, gate447inter10, gate447inter11, gate447inter12, gate404inter0, gate404inter1, gate404inter2, gate404inter3, gate404inter4, gate404inter5, gate404inter6, gate404inter7, gate404inter8, gate404inter9, gate404inter10, gate404inter11, gate404inter12, gate166inter0, gate166inter1, gate166inter2, gate166inter3, gate166inter4, gate166inter5, gate166inter6, gate166inter7, gate166inter8, gate166inter9, gate166inter10, gate166inter11, gate166inter12, gate84inter0, gate84inter1, gate84inter2, gate84inter3, gate84inter4, gate84inter5, gate84inter6, gate84inter7, gate84inter8, gate84inter9, gate84inter10, gate84inter11, gate84inter12, gate460inter0, gate460inter1, gate460inter2, gate460inter3, gate460inter4, gate460inter5, gate460inter6, gate460inter7, gate460inter8, gate460inter9, gate460inter10, gate460inter11, gate460inter12, gate122inter0, gate122inter1, gate122inter2, gate122inter3, gate122inter4, gate122inter5, gate122inter6, gate122inter7, gate122inter8, gate122inter9, gate122inter10, gate122inter11, gate122inter12, gate172inter0, gate172inter1, gate172inter2, gate172inter3, gate172inter4, gate172inter5, gate172inter6, gate172inter7, gate172inter8, gate172inter9, gate172inter10, gate172inter11, gate172inter12, gate25inter0, gate25inter1, gate25inter2, gate25inter3, gate25inter4, gate25inter5, gate25inter6, gate25inter7, gate25inter8, gate25inter9, gate25inter10, gate25inter11, gate25inter12, gate471inter0, gate471inter1, gate471inter2, gate471inter3, gate471inter4, gate471inter5, gate471inter6, gate471inter7, gate471inter8, gate471inter9, gate471inter10, gate471inter11, gate471inter12, gate234inter0, gate234inter1, gate234inter2, gate234inter3, gate234inter4, gate234inter5, gate234inter6, gate234inter7, gate234inter8, gate234inter9, gate234inter10, gate234inter11, gate234inter12, gate180inter0, gate180inter1, gate180inter2, gate180inter3, gate180inter4, gate180inter5, gate180inter6, gate180inter7, gate180inter8, gate180inter9, gate180inter10, gate180inter11, gate180inter12, gate223inter0, gate223inter1, gate223inter2, gate223inter3, gate223inter4, gate223inter5, gate223inter6, gate223inter7, gate223inter8, gate223inter9, gate223inter10, gate223inter11, gate223inter12, gate125inter0, gate125inter1, gate125inter2, gate125inter3, gate125inter4, gate125inter5, gate125inter6, gate125inter7, gate125inter8, gate125inter9, gate125inter10, gate125inter11, gate125inter12, gate83inter0, gate83inter1, gate83inter2, gate83inter3, gate83inter4, gate83inter5, gate83inter6, gate83inter7, gate83inter8, gate83inter9, gate83inter10, gate83inter11, gate83inter12, gate394inter0, gate394inter1, gate394inter2, gate394inter3, gate394inter4, gate394inter5, gate394inter6, gate394inter7, gate394inter8, gate394inter9, gate394inter10, gate394inter11, gate394inter12, gate500inter0, gate500inter1, gate500inter2, gate500inter3, gate500inter4, gate500inter5, gate500inter6, gate500inter7, gate500inter8, gate500inter9, gate500inter10, gate500inter11, gate500inter12, gate503inter0, gate503inter1, gate503inter2, gate503inter3, gate503inter4, gate503inter5, gate503inter6, gate503inter7, gate503inter8, gate503inter9, gate503inter10, gate503inter11, gate503inter12, gate185inter0, gate185inter1, gate185inter2, gate185inter3, gate185inter4, gate185inter5, gate185inter6, gate185inter7, gate185inter8, gate185inter9, gate185inter10, gate185inter11, gate185inter12, gate252inter0, gate252inter1, gate252inter2, gate252inter3, gate252inter4, gate252inter5, gate252inter6, gate252inter7, gate252inter8, gate252inter9, gate252inter10, gate252inter11, gate252inter12, gate33inter0, gate33inter1, gate33inter2, gate33inter3, gate33inter4, gate33inter5, gate33inter6, gate33inter7, gate33inter8, gate33inter9, gate33inter10, gate33inter11, gate33inter12, gate425inter0, gate425inter1, gate425inter2, gate425inter3, gate425inter4, gate425inter5, gate425inter6, gate425inter7, gate425inter8, gate425inter9, gate425inter10, gate425inter11, gate425inter12, gate445inter0, gate445inter1, gate445inter2, gate445inter3, gate445inter4, gate445inter5, gate445inter6, gate445inter7, gate445inter8, gate445inter9, gate445inter10, gate445inter11, gate445inter12, gate497inter0, gate497inter1, gate497inter2, gate497inter3, gate497inter4, gate497inter5, gate497inter6, gate497inter7, gate497inter8, gate497inter9, gate497inter10, gate497inter11, gate497inter12, gate444inter0, gate444inter1, gate444inter2, gate444inter3, gate444inter4, gate444inter5, gate444inter6, gate444inter7, gate444inter8, gate444inter9, gate444inter10, gate444inter11, gate444inter12, gate151inter0, gate151inter1, gate151inter2, gate151inter3, gate151inter4, gate151inter5, gate151inter6, gate151inter7, gate151inter8, gate151inter9, gate151inter10, gate151inter11, gate151inter12, gate251inter0, gate251inter1, gate251inter2, gate251inter3, gate251inter4, gate251inter5, gate251inter6, gate251inter7, gate251inter8, gate251inter9, gate251inter10, gate251inter11, gate251inter12, gate418inter0, gate418inter1, gate418inter2, gate418inter3, gate418inter4, gate418inter5, gate418inter6, gate418inter7, gate418inter8, gate418inter9, gate418inter10, gate418inter11, gate418inter12, gate36inter0, gate36inter1, gate36inter2, gate36inter3, gate36inter4, gate36inter5, gate36inter6, gate36inter7, gate36inter8, gate36inter9, gate36inter10, gate36inter11, gate36inter12, gate53inter0, gate53inter1, gate53inter2, gate53inter3, gate53inter4, gate53inter5, gate53inter6, gate53inter7, gate53inter8, gate53inter9, gate53inter10, gate53inter11, gate53inter12, gate133inter0, gate133inter1, gate133inter2, gate133inter3, gate133inter4, gate133inter5, gate133inter6, gate133inter7, gate133inter8, gate133inter9, gate133inter10, gate133inter11, gate133inter12, gate31inter0, gate31inter1, gate31inter2, gate31inter3, gate31inter4, gate31inter5, gate31inter6, gate31inter7, gate31inter8, gate31inter9, gate31inter10, gate31inter11, gate31inter12, gate144inter0, gate144inter1, gate144inter2, gate144inter3, gate144inter4, gate144inter5, gate144inter6, gate144inter7, gate144inter8, gate144inter9, gate144inter10, gate144inter11, gate144inter12, gate44inter0, gate44inter1, gate44inter2, gate44inter3, gate44inter4, gate44inter5, gate44inter6, gate44inter7, gate44inter8, gate44inter9, gate44inter10, gate44inter11, gate44inter12, gate443inter0, gate443inter1, gate443inter2, gate443inter3, gate443inter4, gate443inter5, gate443inter6, gate443inter7, gate443inter8, gate443inter9, gate443inter10, gate443inter11, gate443inter12, gate417inter0, gate417inter1, gate417inter2, gate417inter3, gate417inter4, gate417inter5, gate417inter6, gate417inter7, gate417inter8, gate417inter9, gate417inter10, gate417inter11, gate417inter12, gate229inter0, gate229inter1, gate229inter2, gate229inter3, gate229inter4, gate229inter5, gate229inter6, gate229inter7, gate229inter8, gate229inter9, gate229inter10, gate229inter11, gate229inter12, gate95inter0, gate95inter1, gate95inter2, gate95inter3, gate95inter4, gate95inter5, gate95inter6, gate95inter7, gate95inter8, gate95inter9, gate95inter10, gate95inter11, gate95inter12, gate167inter0, gate167inter1, gate167inter2, gate167inter3, gate167inter4, gate167inter5, gate167inter6, gate167inter7, gate167inter8, gate167inter9, gate167inter10, gate167inter11, gate167inter12, gate87inter0, gate87inter1, gate87inter2, gate87inter3, gate87inter4, gate87inter5, gate87inter6, gate87inter7, gate87inter8, gate87inter9, gate87inter10, gate87inter11, gate87inter12, gate192inter0, gate192inter1, gate192inter2, gate192inter3, gate192inter4, gate192inter5, gate192inter6, gate192inter7, gate192inter8, gate192inter9, gate192inter10, gate192inter11, gate192inter12, gate120inter0, gate120inter1, gate120inter2, gate120inter3, gate120inter4, gate120inter5, gate120inter6, gate120inter7, gate120inter8, gate120inter9, gate120inter10, gate120inter11, gate120inter12, gate485inter0, gate485inter1, gate485inter2, gate485inter3, gate485inter4, gate485inter5, gate485inter6, gate485inter7, gate485inter8, gate485inter9, gate485inter10, gate485inter11, gate485inter12, gate119inter0, gate119inter1, gate119inter2, gate119inter3, gate119inter4, gate119inter5, gate119inter6, gate119inter7, gate119inter8, gate119inter9, gate119inter10, gate119inter11, gate119inter12, gate66inter0, gate66inter1, gate66inter2, gate66inter3, gate66inter4, gate66inter5, gate66inter6, gate66inter7, gate66inter8, gate66inter9, gate66inter10, gate66inter11, gate66inter12, gate387inter0, gate387inter1, gate387inter2, gate387inter3, gate387inter4, gate387inter5, gate387inter6, gate387inter7, gate387inter8, gate387inter9, gate387inter10, gate387inter11, gate387inter12, gate138inter0, gate138inter1, gate138inter2, gate138inter3, gate138inter4, gate138inter5, gate138inter6, gate138inter7, gate138inter8, gate138inter9, gate138inter10, gate138inter11, gate138inter12, gate157inter0, gate157inter1, gate157inter2, gate157inter3, gate157inter4, gate157inter5, gate157inter6, gate157inter7, gate157inter8, gate157inter9, gate157inter10, gate157inter11, gate157inter12, gate91inter0, gate91inter1, gate91inter2, gate91inter3, gate91inter4, gate91inter5, gate91inter6, gate91inter7, gate91inter8, gate91inter9, gate91inter10, gate91inter11, gate91inter12, gate230inter0, gate230inter1, gate230inter2, gate230inter3, gate230inter4, gate230inter5, gate230inter6, gate230inter7, gate230inter8, gate230inter9, gate230inter10, gate230inter11, gate230inter12, gate152inter0, gate152inter1, gate152inter2, gate152inter3, gate152inter4, gate152inter5, gate152inter6, gate152inter7, gate152inter8, gate152inter9, gate152inter10, gate152inter11, gate152inter12, gate163inter0, gate163inter1, gate163inter2, gate163inter3, gate163inter4, gate163inter5, gate163inter6, gate163inter7, gate163inter8, gate163inter9, gate163inter10, gate163inter11, gate163inter12, gate290inter0, gate290inter1, gate290inter2, gate290inter3, gate290inter4, gate290inter5, gate290inter6, gate290inter7, gate290inter8, gate290inter9, gate290inter10, gate290inter11, gate290inter12, gate513inter0, gate513inter1, gate513inter2, gate513inter3, gate513inter4, gate513inter5, gate513inter6, gate513inter7, gate513inter8, gate513inter9, gate513inter10, gate513inter11, gate513inter12, gate249inter0, gate249inter1, gate249inter2, gate249inter3, gate249inter4, gate249inter5, gate249inter6, gate249inter7, gate249inter8, gate249inter9, gate249inter10, gate249inter11, gate249inter12, gate155inter0, gate155inter1, gate155inter2, gate155inter3, gate155inter4, gate155inter5, gate155inter6, gate155inter7, gate155inter8, gate155inter9, gate155inter10, gate155inter11, gate155inter12, gate414inter0, gate414inter1, gate414inter2, gate414inter3, gate414inter4, gate414inter5, gate414inter6, gate414inter7, gate414inter8, gate414inter9, gate414inter10, gate414inter11, gate414inter12, gate441inter0, gate441inter1, gate441inter2, gate441inter3, gate441inter4, gate441inter5, gate441inter6, gate441inter7, gate441inter8, gate441inter9, gate441inter10, gate441inter11, gate441inter12;



and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );

  xor2  gate1345(.a(G2), .b(G1), .O(gate9inter0));
  nand2 gate1346(.a(gate9inter0), .b(s_114), .O(gate9inter1));
  and2  gate1347(.a(G2), .b(G1), .O(gate9inter2));
  inv1  gate1348(.a(s_114), .O(gate9inter3));
  inv1  gate1349(.a(s_115), .O(gate9inter4));
  nand2 gate1350(.a(gate9inter4), .b(gate9inter3), .O(gate9inter5));
  nor2  gate1351(.a(gate9inter5), .b(gate9inter2), .O(gate9inter6));
  inv1  gate1352(.a(G1), .O(gate9inter7));
  inv1  gate1353(.a(G2), .O(gate9inter8));
  nand2 gate1354(.a(gate9inter8), .b(gate9inter7), .O(gate9inter9));
  nand2 gate1355(.a(s_115), .b(gate9inter3), .O(gate9inter10));
  nor2  gate1356(.a(gate9inter10), .b(gate9inter9), .O(gate9inter11));
  nor2  gate1357(.a(gate9inter11), .b(gate9inter6), .O(gate9inter12));
  nand2 gate1358(.a(gate9inter12), .b(gate9inter1), .O(G266));
nand2 gate10( .a(G3), .b(G4), .O(G269) );
nand2 gate11( .a(G5), .b(G6), .O(G272) );
nand2 gate12( .a(G7), .b(G8), .O(G275) );
nand2 gate13( .a(G9), .b(G10), .O(G278) );
nand2 gate14( .a(G11), .b(G12), .O(G281) );
nand2 gate15( .a(G13), .b(G14), .O(G284) );
nand2 gate16( .a(G15), .b(G16), .O(G287) );
nand2 gate17( .a(G17), .b(G18), .O(G290) );
nand2 gate18( .a(G19), .b(G20), .O(G293) );
nand2 gate19( .a(G21), .b(G22), .O(G296) );
nand2 gate20( .a(G23), .b(G24), .O(G299) );
nand2 gate21( .a(G25), .b(G26), .O(G302) );
nand2 gate22( .a(G27), .b(G28), .O(G305) );
nand2 gate23( .a(G29), .b(G30), .O(G308) );
nand2 gate24( .a(G31), .b(G32), .O(G311) );

  xor2  gate1751(.a(G5), .b(G1), .O(gate25inter0));
  nand2 gate1752(.a(gate25inter0), .b(s_172), .O(gate25inter1));
  and2  gate1753(.a(G5), .b(G1), .O(gate25inter2));
  inv1  gate1754(.a(s_172), .O(gate25inter3));
  inv1  gate1755(.a(s_173), .O(gate25inter4));
  nand2 gate1756(.a(gate25inter4), .b(gate25inter3), .O(gate25inter5));
  nor2  gate1757(.a(gate25inter5), .b(gate25inter2), .O(gate25inter6));
  inv1  gate1758(.a(G1), .O(gate25inter7));
  inv1  gate1759(.a(G5), .O(gate25inter8));
  nand2 gate1760(.a(gate25inter8), .b(gate25inter7), .O(gate25inter9));
  nand2 gate1761(.a(s_173), .b(gate25inter3), .O(gate25inter10));
  nor2  gate1762(.a(gate25inter10), .b(gate25inter9), .O(gate25inter11));
  nor2  gate1763(.a(gate25inter11), .b(gate25inter6), .O(gate25inter12));
  nand2 gate1764(.a(gate25inter12), .b(gate25inter1), .O(G314));
nand2 gate26( .a(G9), .b(G13), .O(G317) );
nand2 gate27( .a(G2), .b(G6), .O(G320) );

  xor2  gate589(.a(G14), .b(G10), .O(gate28inter0));
  nand2 gate590(.a(gate28inter0), .b(s_6), .O(gate28inter1));
  and2  gate591(.a(G14), .b(G10), .O(gate28inter2));
  inv1  gate592(.a(s_6), .O(gate28inter3));
  inv1  gate593(.a(s_7), .O(gate28inter4));
  nand2 gate594(.a(gate28inter4), .b(gate28inter3), .O(gate28inter5));
  nor2  gate595(.a(gate28inter5), .b(gate28inter2), .O(gate28inter6));
  inv1  gate596(.a(G10), .O(gate28inter7));
  inv1  gate597(.a(G14), .O(gate28inter8));
  nand2 gate598(.a(gate28inter8), .b(gate28inter7), .O(gate28inter9));
  nand2 gate599(.a(s_7), .b(gate28inter3), .O(gate28inter10));
  nor2  gate600(.a(gate28inter10), .b(gate28inter9), .O(gate28inter11));
  nor2  gate601(.a(gate28inter11), .b(gate28inter6), .O(gate28inter12));
  nand2 gate602(.a(gate28inter12), .b(gate28inter1), .O(G323));
nand2 gate29( .a(G3), .b(G7), .O(G326) );

  xor2  gate1275(.a(G15), .b(G11), .O(gate30inter0));
  nand2 gate1276(.a(gate30inter0), .b(s_104), .O(gate30inter1));
  and2  gate1277(.a(G15), .b(G11), .O(gate30inter2));
  inv1  gate1278(.a(s_104), .O(gate30inter3));
  inv1  gate1279(.a(s_105), .O(gate30inter4));
  nand2 gate1280(.a(gate30inter4), .b(gate30inter3), .O(gate30inter5));
  nor2  gate1281(.a(gate30inter5), .b(gate30inter2), .O(gate30inter6));
  inv1  gate1282(.a(G11), .O(gate30inter7));
  inv1  gate1283(.a(G15), .O(gate30inter8));
  nand2 gate1284(.a(gate30inter8), .b(gate30inter7), .O(gate30inter9));
  nand2 gate1285(.a(s_105), .b(gate30inter3), .O(gate30inter10));
  nor2  gate1286(.a(gate30inter10), .b(gate30inter9), .O(gate30inter11));
  nor2  gate1287(.a(gate30inter11), .b(gate30inter6), .O(gate30inter12));
  nand2 gate1288(.a(gate30inter12), .b(gate30inter1), .O(G329));

  xor2  gate2073(.a(G8), .b(G4), .O(gate31inter0));
  nand2 gate2074(.a(gate31inter0), .b(s_218), .O(gate31inter1));
  and2  gate2075(.a(G8), .b(G4), .O(gate31inter2));
  inv1  gate2076(.a(s_218), .O(gate31inter3));
  inv1  gate2077(.a(s_219), .O(gate31inter4));
  nand2 gate2078(.a(gate31inter4), .b(gate31inter3), .O(gate31inter5));
  nor2  gate2079(.a(gate31inter5), .b(gate31inter2), .O(gate31inter6));
  inv1  gate2080(.a(G4), .O(gate31inter7));
  inv1  gate2081(.a(G8), .O(gate31inter8));
  nand2 gate2082(.a(gate31inter8), .b(gate31inter7), .O(gate31inter9));
  nand2 gate2083(.a(s_219), .b(gate31inter3), .O(gate31inter10));
  nor2  gate2084(.a(gate31inter10), .b(gate31inter9), .O(gate31inter11));
  nor2  gate2085(.a(gate31inter11), .b(gate31inter6), .O(gate31inter12));
  nand2 gate2086(.a(gate31inter12), .b(gate31inter1), .O(G332));
nand2 gate32( .a(G12), .b(G16), .O(G335) );

  xor2  gate1919(.a(G21), .b(G17), .O(gate33inter0));
  nand2 gate1920(.a(gate33inter0), .b(s_196), .O(gate33inter1));
  and2  gate1921(.a(G21), .b(G17), .O(gate33inter2));
  inv1  gate1922(.a(s_196), .O(gate33inter3));
  inv1  gate1923(.a(s_197), .O(gate33inter4));
  nand2 gate1924(.a(gate33inter4), .b(gate33inter3), .O(gate33inter5));
  nor2  gate1925(.a(gate33inter5), .b(gate33inter2), .O(gate33inter6));
  inv1  gate1926(.a(G17), .O(gate33inter7));
  inv1  gate1927(.a(G21), .O(gate33inter8));
  nand2 gate1928(.a(gate33inter8), .b(gate33inter7), .O(gate33inter9));
  nand2 gate1929(.a(s_197), .b(gate33inter3), .O(gate33inter10));
  nor2  gate1930(.a(gate33inter10), .b(gate33inter9), .O(gate33inter11));
  nor2  gate1931(.a(gate33inter11), .b(gate33inter6), .O(gate33inter12));
  nand2 gate1932(.a(gate33inter12), .b(gate33inter1), .O(G338));
nand2 gate34( .a(G25), .b(G29), .O(G341) );

  xor2  gate1583(.a(G22), .b(G18), .O(gate35inter0));
  nand2 gate1584(.a(gate35inter0), .b(s_148), .O(gate35inter1));
  and2  gate1585(.a(G22), .b(G18), .O(gate35inter2));
  inv1  gate1586(.a(s_148), .O(gate35inter3));
  inv1  gate1587(.a(s_149), .O(gate35inter4));
  nand2 gate1588(.a(gate35inter4), .b(gate35inter3), .O(gate35inter5));
  nor2  gate1589(.a(gate35inter5), .b(gate35inter2), .O(gate35inter6));
  inv1  gate1590(.a(G18), .O(gate35inter7));
  inv1  gate1591(.a(G22), .O(gate35inter8));
  nand2 gate1592(.a(gate35inter8), .b(gate35inter7), .O(gate35inter9));
  nand2 gate1593(.a(s_149), .b(gate35inter3), .O(gate35inter10));
  nor2  gate1594(.a(gate35inter10), .b(gate35inter9), .O(gate35inter11));
  nor2  gate1595(.a(gate35inter11), .b(gate35inter6), .O(gate35inter12));
  nand2 gate1596(.a(gate35inter12), .b(gate35inter1), .O(G344));

  xor2  gate2031(.a(G30), .b(G26), .O(gate36inter0));
  nand2 gate2032(.a(gate36inter0), .b(s_212), .O(gate36inter1));
  and2  gate2033(.a(G30), .b(G26), .O(gate36inter2));
  inv1  gate2034(.a(s_212), .O(gate36inter3));
  inv1  gate2035(.a(s_213), .O(gate36inter4));
  nand2 gate2036(.a(gate36inter4), .b(gate36inter3), .O(gate36inter5));
  nor2  gate2037(.a(gate36inter5), .b(gate36inter2), .O(gate36inter6));
  inv1  gate2038(.a(G26), .O(gate36inter7));
  inv1  gate2039(.a(G30), .O(gate36inter8));
  nand2 gate2040(.a(gate36inter8), .b(gate36inter7), .O(gate36inter9));
  nand2 gate2041(.a(s_213), .b(gate36inter3), .O(gate36inter10));
  nor2  gate2042(.a(gate36inter10), .b(gate36inter9), .O(gate36inter11));
  nor2  gate2043(.a(gate36inter11), .b(gate36inter6), .O(gate36inter12));
  nand2 gate2044(.a(gate36inter12), .b(gate36inter1), .O(G347));

  xor2  gate757(.a(G23), .b(G19), .O(gate37inter0));
  nand2 gate758(.a(gate37inter0), .b(s_30), .O(gate37inter1));
  and2  gate759(.a(G23), .b(G19), .O(gate37inter2));
  inv1  gate760(.a(s_30), .O(gate37inter3));
  inv1  gate761(.a(s_31), .O(gate37inter4));
  nand2 gate762(.a(gate37inter4), .b(gate37inter3), .O(gate37inter5));
  nor2  gate763(.a(gate37inter5), .b(gate37inter2), .O(gate37inter6));
  inv1  gate764(.a(G19), .O(gate37inter7));
  inv1  gate765(.a(G23), .O(gate37inter8));
  nand2 gate766(.a(gate37inter8), .b(gate37inter7), .O(gate37inter9));
  nand2 gate767(.a(s_31), .b(gate37inter3), .O(gate37inter10));
  nor2  gate768(.a(gate37inter10), .b(gate37inter9), .O(gate37inter11));
  nor2  gate769(.a(gate37inter11), .b(gate37inter6), .O(gate37inter12));
  nand2 gate770(.a(gate37inter12), .b(gate37inter1), .O(G350));
nand2 gate38( .a(G27), .b(G31), .O(G353) );
nand2 gate39( .a(G20), .b(G24), .O(G356) );
nand2 gate40( .a(G28), .b(G32), .O(G359) );
nand2 gate41( .a(G1), .b(G266), .O(G362) );
nand2 gate42( .a(G2), .b(G266), .O(G363) );

  xor2  gate1037(.a(G269), .b(G3), .O(gate43inter0));
  nand2 gate1038(.a(gate43inter0), .b(s_70), .O(gate43inter1));
  and2  gate1039(.a(G269), .b(G3), .O(gate43inter2));
  inv1  gate1040(.a(s_70), .O(gate43inter3));
  inv1  gate1041(.a(s_71), .O(gate43inter4));
  nand2 gate1042(.a(gate43inter4), .b(gate43inter3), .O(gate43inter5));
  nor2  gate1043(.a(gate43inter5), .b(gate43inter2), .O(gate43inter6));
  inv1  gate1044(.a(G3), .O(gate43inter7));
  inv1  gate1045(.a(G269), .O(gate43inter8));
  nand2 gate1046(.a(gate43inter8), .b(gate43inter7), .O(gate43inter9));
  nand2 gate1047(.a(s_71), .b(gate43inter3), .O(gate43inter10));
  nor2  gate1048(.a(gate43inter10), .b(gate43inter9), .O(gate43inter11));
  nor2  gate1049(.a(gate43inter11), .b(gate43inter6), .O(gate43inter12));
  nand2 gate1050(.a(gate43inter12), .b(gate43inter1), .O(G364));

  xor2  gate2101(.a(G269), .b(G4), .O(gate44inter0));
  nand2 gate2102(.a(gate44inter0), .b(s_222), .O(gate44inter1));
  and2  gate2103(.a(G269), .b(G4), .O(gate44inter2));
  inv1  gate2104(.a(s_222), .O(gate44inter3));
  inv1  gate2105(.a(s_223), .O(gate44inter4));
  nand2 gate2106(.a(gate44inter4), .b(gate44inter3), .O(gate44inter5));
  nor2  gate2107(.a(gate44inter5), .b(gate44inter2), .O(gate44inter6));
  inv1  gate2108(.a(G4), .O(gate44inter7));
  inv1  gate2109(.a(G269), .O(gate44inter8));
  nand2 gate2110(.a(gate44inter8), .b(gate44inter7), .O(gate44inter9));
  nand2 gate2111(.a(s_223), .b(gate44inter3), .O(gate44inter10));
  nor2  gate2112(.a(gate44inter10), .b(gate44inter9), .O(gate44inter11));
  nor2  gate2113(.a(gate44inter11), .b(gate44inter6), .O(gate44inter12));
  nand2 gate2114(.a(gate44inter12), .b(gate44inter1), .O(G365));
nand2 gate45( .a(G5), .b(G272), .O(G366) );

  xor2  gate561(.a(G272), .b(G6), .O(gate46inter0));
  nand2 gate562(.a(gate46inter0), .b(s_2), .O(gate46inter1));
  and2  gate563(.a(G272), .b(G6), .O(gate46inter2));
  inv1  gate564(.a(s_2), .O(gate46inter3));
  inv1  gate565(.a(s_3), .O(gate46inter4));
  nand2 gate566(.a(gate46inter4), .b(gate46inter3), .O(gate46inter5));
  nor2  gate567(.a(gate46inter5), .b(gate46inter2), .O(gate46inter6));
  inv1  gate568(.a(G6), .O(gate46inter7));
  inv1  gate569(.a(G272), .O(gate46inter8));
  nand2 gate570(.a(gate46inter8), .b(gate46inter7), .O(gate46inter9));
  nand2 gate571(.a(s_3), .b(gate46inter3), .O(gate46inter10));
  nor2  gate572(.a(gate46inter10), .b(gate46inter9), .O(gate46inter11));
  nor2  gate573(.a(gate46inter11), .b(gate46inter6), .O(gate46inter12));
  nand2 gate574(.a(gate46inter12), .b(gate46inter1), .O(G367));
nand2 gate47( .a(G7), .b(G275), .O(G368) );
nand2 gate48( .a(G8), .b(G275), .O(G369) );
nand2 gate49( .a(G9), .b(G278), .O(G370) );
nand2 gate50( .a(G10), .b(G278), .O(G371) );
nand2 gate51( .a(G11), .b(G281), .O(G372) );
nand2 gate52( .a(G12), .b(G281), .O(G373) );

  xor2  gate2045(.a(G284), .b(G13), .O(gate53inter0));
  nand2 gate2046(.a(gate53inter0), .b(s_214), .O(gate53inter1));
  and2  gate2047(.a(G284), .b(G13), .O(gate53inter2));
  inv1  gate2048(.a(s_214), .O(gate53inter3));
  inv1  gate2049(.a(s_215), .O(gate53inter4));
  nand2 gate2050(.a(gate53inter4), .b(gate53inter3), .O(gate53inter5));
  nor2  gate2051(.a(gate53inter5), .b(gate53inter2), .O(gate53inter6));
  inv1  gate2052(.a(G13), .O(gate53inter7));
  inv1  gate2053(.a(G284), .O(gate53inter8));
  nand2 gate2054(.a(gate53inter8), .b(gate53inter7), .O(gate53inter9));
  nand2 gate2055(.a(s_215), .b(gate53inter3), .O(gate53inter10));
  nor2  gate2056(.a(gate53inter10), .b(gate53inter9), .O(gate53inter11));
  nor2  gate2057(.a(gate53inter11), .b(gate53inter6), .O(gate53inter12));
  nand2 gate2058(.a(gate53inter12), .b(gate53inter1), .O(G374));
nand2 gate54( .a(G14), .b(G284), .O(G375) );

  xor2  gate897(.a(G287), .b(G15), .O(gate55inter0));
  nand2 gate898(.a(gate55inter0), .b(s_50), .O(gate55inter1));
  and2  gate899(.a(G287), .b(G15), .O(gate55inter2));
  inv1  gate900(.a(s_50), .O(gate55inter3));
  inv1  gate901(.a(s_51), .O(gate55inter4));
  nand2 gate902(.a(gate55inter4), .b(gate55inter3), .O(gate55inter5));
  nor2  gate903(.a(gate55inter5), .b(gate55inter2), .O(gate55inter6));
  inv1  gate904(.a(G15), .O(gate55inter7));
  inv1  gate905(.a(G287), .O(gate55inter8));
  nand2 gate906(.a(gate55inter8), .b(gate55inter7), .O(gate55inter9));
  nand2 gate907(.a(s_51), .b(gate55inter3), .O(gate55inter10));
  nor2  gate908(.a(gate55inter10), .b(gate55inter9), .O(gate55inter11));
  nor2  gate909(.a(gate55inter11), .b(gate55inter6), .O(gate55inter12));
  nand2 gate910(.a(gate55inter12), .b(gate55inter1), .O(G376));
nand2 gate56( .a(G16), .b(G287), .O(G377) );
nand2 gate57( .a(G17), .b(G290), .O(G378) );
nand2 gate58( .a(G18), .b(G290), .O(G379) );
nand2 gate59( .a(G19), .b(G293), .O(G380) );
nand2 gate60( .a(G20), .b(G293), .O(G381) );
nand2 gate61( .a(G21), .b(G296), .O(G382) );
nand2 gate62( .a(G22), .b(G296), .O(G383) );
nand2 gate63( .a(G23), .b(G299), .O(G384) );
nand2 gate64( .a(G24), .b(G299), .O(G385) );

  xor2  gate1569(.a(G302), .b(G25), .O(gate65inter0));
  nand2 gate1570(.a(gate65inter0), .b(s_146), .O(gate65inter1));
  and2  gate1571(.a(G302), .b(G25), .O(gate65inter2));
  inv1  gate1572(.a(s_146), .O(gate65inter3));
  inv1  gate1573(.a(s_147), .O(gate65inter4));
  nand2 gate1574(.a(gate65inter4), .b(gate65inter3), .O(gate65inter5));
  nor2  gate1575(.a(gate65inter5), .b(gate65inter2), .O(gate65inter6));
  inv1  gate1576(.a(G25), .O(gate65inter7));
  inv1  gate1577(.a(G302), .O(gate65inter8));
  nand2 gate1578(.a(gate65inter8), .b(gate65inter7), .O(gate65inter9));
  nand2 gate1579(.a(s_147), .b(gate65inter3), .O(gate65inter10));
  nor2  gate1580(.a(gate65inter10), .b(gate65inter9), .O(gate65inter11));
  nor2  gate1581(.a(gate65inter11), .b(gate65inter6), .O(gate65inter12));
  nand2 gate1582(.a(gate65inter12), .b(gate65inter1), .O(G386));

  xor2  gate2255(.a(G302), .b(G26), .O(gate66inter0));
  nand2 gate2256(.a(gate66inter0), .b(s_244), .O(gate66inter1));
  and2  gate2257(.a(G302), .b(G26), .O(gate66inter2));
  inv1  gate2258(.a(s_244), .O(gate66inter3));
  inv1  gate2259(.a(s_245), .O(gate66inter4));
  nand2 gate2260(.a(gate66inter4), .b(gate66inter3), .O(gate66inter5));
  nor2  gate2261(.a(gate66inter5), .b(gate66inter2), .O(gate66inter6));
  inv1  gate2262(.a(G26), .O(gate66inter7));
  inv1  gate2263(.a(G302), .O(gate66inter8));
  nand2 gate2264(.a(gate66inter8), .b(gate66inter7), .O(gate66inter9));
  nand2 gate2265(.a(s_245), .b(gate66inter3), .O(gate66inter10));
  nor2  gate2266(.a(gate66inter10), .b(gate66inter9), .O(gate66inter11));
  nor2  gate2267(.a(gate66inter11), .b(gate66inter6), .O(gate66inter12));
  nand2 gate2268(.a(gate66inter12), .b(gate66inter1), .O(G387));
nand2 gate67( .a(G27), .b(G305), .O(G388) );
nand2 gate68( .a(G28), .b(G305), .O(G389) );
nand2 gate69( .a(G29), .b(G308), .O(G390) );
nand2 gate70( .a(G30), .b(G308), .O(G391) );
nand2 gate71( .a(G31), .b(G311), .O(G392) );
nand2 gate72( .a(G32), .b(G311), .O(G393) );
nand2 gate73( .a(G1), .b(G314), .O(G394) );
nand2 gate74( .a(G5), .b(G314), .O(G395) );
nand2 gate75( .a(G9), .b(G317), .O(G396) );
nand2 gate76( .a(G13), .b(G317), .O(G397) );

  xor2  gate687(.a(G320), .b(G2), .O(gate77inter0));
  nand2 gate688(.a(gate77inter0), .b(s_20), .O(gate77inter1));
  and2  gate689(.a(G320), .b(G2), .O(gate77inter2));
  inv1  gate690(.a(s_20), .O(gate77inter3));
  inv1  gate691(.a(s_21), .O(gate77inter4));
  nand2 gate692(.a(gate77inter4), .b(gate77inter3), .O(gate77inter5));
  nor2  gate693(.a(gate77inter5), .b(gate77inter2), .O(gate77inter6));
  inv1  gate694(.a(G2), .O(gate77inter7));
  inv1  gate695(.a(G320), .O(gate77inter8));
  nand2 gate696(.a(gate77inter8), .b(gate77inter7), .O(gate77inter9));
  nand2 gate697(.a(s_21), .b(gate77inter3), .O(gate77inter10));
  nor2  gate698(.a(gate77inter10), .b(gate77inter9), .O(gate77inter11));
  nor2  gate699(.a(gate77inter11), .b(gate77inter6), .O(gate77inter12));
  nand2 gate700(.a(gate77inter12), .b(gate77inter1), .O(G398));

  xor2  gate575(.a(G320), .b(G6), .O(gate78inter0));
  nand2 gate576(.a(gate78inter0), .b(s_4), .O(gate78inter1));
  and2  gate577(.a(G320), .b(G6), .O(gate78inter2));
  inv1  gate578(.a(s_4), .O(gate78inter3));
  inv1  gate579(.a(s_5), .O(gate78inter4));
  nand2 gate580(.a(gate78inter4), .b(gate78inter3), .O(gate78inter5));
  nor2  gate581(.a(gate78inter5), .b(gate78inter2), .O(gate78inter6));
  inv1  gate582(.a(G6), .O(gate78inter7));
  inv1  gate583(.a(G320), .O(gate78inter8));
  nand2 gate584(.a(gate78inter8), .b(gate78inter7), .O(gate78inter9));
  nand2 gate585(.a(s_5), .b(gate78inter3), .O(gate78inter10));
  nor2  gate586(.a(gate78inter10), .b(gate78inter9), .O(gate78inter11));
  nor2  gate587(.a(gate78inter11), .b(gate78inter6), .O(gate78inter12));
  nand2 gate588(.a(gate78inter12), .b(gate78inter1), .O(G399));

  xor2  gate1317(.a(G323), .b(G10), .O(gate79inter0));
  nand2 gate1318(.a(gate79inter0), .b(s_110), .O(gate79inter1));
  and2  gate1319(.a(G323), .b(G10), .O(gate79inter2));
  inv1  gate1320(.a(s_110), .O(gate79inter3));
  inv1  gate1321(.a(s_111), .O(gate79inter4));
  nand2 gate1322(.a(gate79inter4), .b(gate79inter3), .O(gate79inter5));
  nor2  gate1323(.a(gate79inter5), .b(gate79inter2), .O(gate79inter6));
  inv1  gate1324(.a(G10), .O(gate79inter7));
  inv1  gate1325(.a(G323), .O(gate79inter8));
  nand2 gate1326(.a(gate79inter8), .b(gate79inter7), .O(gate79inter9));
  nand2 gate1327(.a(s_111), .b(gate79inter3), .O(gate79inter10));
  nor2  gate1328(.a(gate79inter10), .b(gate79inter9), .O(gate79inter11));
  nor2  gate1329(.a(gate79inter11), .b(gate79inter6), .O(gate79inter12));
  nand2 gate1330(.a(gate79inter12), .b(gate79inter1), .O(G400));
nand2 gate80( .a(G14), .b(G323), .O(G401) );

  xor2  gate1401(.a(G326), .b(G3), .O(gate81inter0));
  nand2 gate1402(.a(gate81inter0), .b(s_122), .O(gate81inter1));
  and2  gate1403(.a(G326), .b(G3), .O(gate81inter2));
  inv1  gate1404(.a(s_122), .O(gate81inter3));
  inv1  gate1405(.a(s_123), .O(gate81inter4));
  nand2 gate1406(.a(gate81inter4), .b(gate81inter3), .O(gate81inter5));
  nor2  gate1407(.a(gate81inter5), .b(gate81inter2), .O(gate81inter6));
  inv1  gate1408(.a(G3), .O(gate81inter7));
  inv1  gate1409(.a(G326), .O(gate81inter8));
  nand2 gate1410(.a(gate81inter8), .b(gate81inter7), .O(gate81inter9));
  nand2 gate1411(.a(s_123), .b(gate81inter3), .O(gate81inter10));
  nor2  gate1412(.a(gate81inter10), .b(gate81inter9), .O(gate81inter11));
  nor2  gate1413(.a(gate81inter11), .b(gate81inter6), .O(gate81inter12));
  nand2 gate1414(.a(gate81inter12), .b(gate81inter1), .O(G402));

  xor2  gate1191(.a(G326), .b(G7), .O(gate82inter0));
  nand2 gate1192(.a(gate82inter0), .b(s_92), .O(gate82inter1));
  and2  gate1193(.a(G326), .b(G7), .O(gate82inter2));
  inv1  gate1194(.a(s_92), .O(gate82inter3));
  inv1  gate1195(.a(s_93), .O(gate82inter4));
  nand2 gate1196(.a(gate82inter4), .b(gate82inter3), .O(gate82inter5));
  nor2  gate1197(.a(gate82inter5), .b(gate82inter2), .O(gate82inter6));
  inv1  gate1198(.a(G7), .O(gate82inter7));
  inv1  gate1199(.a(G326), .O(gate82inter8));
  nand2 gate1200(.a(gate82inter8), .b(gate82inter7), .O(gate82inter9));
  nand2 gate1201(.a(s_93), .b(gate82inter3), .O(gate82inter10));
  nor2  gate1202(.a(gate82inter10), .b(gate82inter9), .O(gate82inter11));
  nor2  gate1203(.a(gate82inter11), .b(gate82inter6), .O(gate82inter12));
  nand2 gate1204(.a(gate82inter12), .b(gate82inter1), .O(G403));

  xor2  gate1835(.a(G329), .b(G11), .O(gate83inter0));
  nand2 gate1836(.a(gate83inter0), .b(s_184), .O(gate83inter1));
  and2  gate1837(.a(G329), .b(G11), .O(gate83inter2));
  inv1  gate1838(.a(s_184), .O(gate83inter3));
  inv1  gate1839(.a(s_185), .O(gate83inter4));
  nand2 gate1840(.a(gate83inter4), .b(gate83inter3), .O(gate83inter5));
  nor2  gate1841(.a(gate83inter5), .b(gate83inter2), .O(gate83inter6));
  inv1  gate1842(.a(G11), .O(gate83inter7));
  inv1  gate1843(.a(G329), .O(gate83inter8));
  nand2 gate1844(.a(gate83inter8), .b(gate83inter7), .O(gate83inter9));
  nand2 gate1845(.a(s_185), .b(gate83inter3), .O(gate83inter10));
  nor2  gate1846(.a(gate83inter10), .b(gate83inter9), .O(gate83inter11));
  nor2  gate1847(.a(gate83inter11), .b(gate83inter6), .O(gate83inter12));
  nand2 gate1848(.a(gate83inter12), .b(gate83inter1), .O(G404));

  xor2  gate1695(.a(G329), .b(G15), .O(gate84inter0));
  nand2 gate1696(.a(gate84inter0), .b(s_164), .O(gate84inter1));
  and2  gate1697(.a(G329), .b(G15), .O(gate84inter2));
  inv1  gate1698(.a(s_164), .O(gate84inter3));
  inv1  gate1699(.a(s_165), .O(gate84inter4));
  nand2 gate1700(.a(gate84inter4), .b(gate84inter3), .O(gate84inter5));
  nor2  gate1701(.a(gate84inter5), .b(gate84inter2), .O(gate84inter6));
  inv1  gate1702(.a(G15), .O(gate84inter7));
  inv1  gate1703(.a(G329), .O(gate84inter8));
  nand2 gate1704(.a(gate84inter8), .b(gate84inter7), .O(gate84inter9));
  nand2 gate1705(.a(s_165), .b(gate84inter3), .O(gate84inter10));
  nor2  gate1706(.a(gate84inter10), .b(gate84inter9), .O(gate84inter11));
  nor2  gate1707(.a(gate84inter11), .b(gate84inter6), .O(gate84inter12));
  nand2 gate1708(.a(gate84inter12), .b(gate84inter1), .O(G405));
nand2 gate85( .a(G4), .b(G332), .O(G406) );

  xor2  gate1429(.a(G332), .b(G8), .O(gate86inter0));
  nand2 gate1430(.a(gate86inter0), .b(s_126), .O(gate86inter1));
  and2  gate1431(.a(G332), .b(G8), .O(gate86inter2));
  inv1  gate1432(.a(s_126), .O(gate86inter3));
  inv1  gate1433(.a(s_127), .O(gate86inter4));
  nand2 gate1434(.a(gate86inter4), .b(gate86inter3), .O(gate86inter5));
  nor2  gate1435(.a(gate86inter5), .b(gate86inter2), .O(gate86inter6));
  inv1  gate1436(.a(G8), .O(gate86inter7));
  inv1  gate1437(.a(G332), .O(gate86inter8));
  nand2 gate1438(.a(gate86inter8), .b(gate86inter7), .O(gate86inter9));
  nand2 gate1439(.a(s_127), .b(gate86inter3), .O(gate86inter10));
  nor2  gate1440(.a(gate86inter10), .b(gate86inter9), .O(gate86inter11));
  nor2  gate1441(.a(gate86inter11), .b(gate86inter6), .O(gate86inter12));
  nand2 gate1442(.a(gate86inter12), .b(gate86inter1), .O(G407));

  xor2  gate2185(.a(G335), .b(G12), .O(gate87inter0));
  nand2 gate2186(.a(gate87inter0), .b(s_234), .O(gate87inter1));
  and2  gate2187(.a(G335), .b(G12), .O(gate87inter2));
  inv1  gate2188(.a(s_234), .O(gate87inter3));
  inv1  gate2189(.a(s_235), .O(gate87inter4));
  nand2 gate2190(.a(gate87inter4), .b(gate87inter3), .O(gate87inter5));
  nor2  gate2191(.a(gate87inter5), .b(gate87inter2), .O(gate87inter6));
  inv1  gate2192(.a(G12), .O(gate87inter7));
  inv1  gate2193(.a(G335), .O(gate87inter8));
  nand2 gate2194(.a(gate87inter8), .b(gate87inter7), .O(gate87inter9));
  nand2 gate2195(.a(s_235), .b(gate87inter3), .O(gate87inter10));
  nor2  gate2196(.a(gate87inter10), .b(gate87inter9), .O(gate87inter11));
  nor2  gate2197(.a(gate87inter11), .b(gate87inter6), .O(gate87inter12));
  nand2 gate2198(.a(gate87inter12), .b(gate87inter1), .O(G408));
nand2 gate88( .a(G16), .b(G335), .O(G409) );

  xor2  gate799(.a(G338), .b(G17), .O(gate89inter0));
  nand2 gate800(.a(gate89inter0), .b(s_36), .O(gate89inter1));
  and2  gate801(.a(G338), .b(G17), .O(gate89inter2));
  inv1  gate802(.a(s_36), .O(gate89inter3));
  inv1  gate803(.a(s_37), .O(gate89inter4));
  nand2 gate804(.a(gate89inter4), .b(gate89inter3), .O(gate89inter5));
  nor2  gate805(.a(gate89inter5), .b(gate89inter2), .O(gate89inter6));
  inv1  gate806(.a(G17), .O(gate89inter7));
  inv1  gate807(.a(G338), .O(gate89inter8));
  nand2 gate808(.a(gate89inter8), .b(gate89inter7), .O(gate89inter9));
  nand2 gate809(.a(s_37), .b(gate89inter3), .O(gate89inter10));
  nor2  gate810(.a(gate89inter10), .b(gate89inter9), .O(gate89inter11));
  nor2  gate811(.a(gate89inter11), .b(gate89inter6), .O(gate89inter12));
  nand2 gate812(.a(gate89inter12), .b(gate89inter1), .O(G410));
nand2 gate90( .a(G21), .b(G338), .O(G411) );

  xor2  gate2311(.a(G341), .b(G25), .O(gate91inter0));
  nand2 gate2312(.a(gate91inter0), .b(s_252), .O(gate91inter1));
  and2  gate2313(.a(G341), .b(G25), .O(gate91inter2));
  inv1  gate2314(.a(s_252), .O(gate91inter3));
  inv1  gate2315(.a(s_253), .O(gate91inter4));
  nand2 gate2316(.a(gate91inter4), .b(gate91inter3), .O(gate91inter5));
  nor2  gate2317(.a(gate91inter5), .b(gate91inter2), .O(gate91inter6));
  inv1  gate2318(.a(G25), .O(gate91inter7));
  inv1  gate2319(.a(G341), .O(gate91inter8));
  nand2 gate2320(.a(gate91inter8), .b(gate91inter7), .O(gate91inter9));
  nand2 gate2321(.a(s_253), .b(gate91inter3), .O(gate91inter10));
  nor2  gate2322(.a(gate91inter10), .b(gate91inter9), .O(gate91inter11));
  nor2  gate2323(.a(gate91inter11), .b(gate91inter6), .O(gate91inter12));
  nand2 gate2324(.a(gate91inter12), .b(gate91inter1), .O(G412));

  xor2  gate1289(.a(G341), .b(G29), .O(gate92inter0));
  nand2 gate1290(.a(gate92inter0), .b(s_106), .O(gate92inter1));
  and2  gate1291(.a(G341), .b(G29), .O(gate92inter2));
  inv1  gate1292(.a(s_106), .O(gate92inter3));
  inv1  gate1293(.a(s_107), .O(gate92inter4));
  nand2 gate1294(.a(gate92inter4), .b(gate92inter3), .O(gate92inter5));
  nor2  gate1295(.a(gate92inter5), .b(gate92inter2), .O(gate92inter6));
  inv1  gate1296(.a(G29), .O(gate92inter7));
  inv1  gate1297(.a(G341), .O(gate92inter8));
  nand2 gate1298(.a(gate92inter8), .b(gate92inter7), .O(gate92inter9));
  nand2 gate1299(.a(s_107), .b(gate92inter3), .O(gate92inter10));
  nor2  gate1300(.a(gate92inter10), .b(gate92inter9), .O(gate92inter11));
  nor2  gate1301(.a(gate92inter11), .b(gate92inter6), .O(gate92inter12));
  nand2 gate1302(.a(gate92inter12), .b(gate92inter1), .O(G413));
nand2 gate93( .a(G18), .b(G344), .O(G414) );
nand2 gate94( .a(G22), .b(G344), .O(G415) );

  xor2  gate2157(.a(G347), .b(G26), .O(gate95inter0));
  nand2 gate2158(.a(gate95inter0), .b(s_230), .O(gate95inter1));
  and2  gate2159(.a(G347), .b(G26), .O(gate95inter2));
  inv1  gate2160(.a(s_230), .O(gate95inter3));
  inv1  gate2161(.a(s_231), .O(gate95inter4));
  nand2 gate2162(.a(gate95inter4), .b(gate95inter3), .O(gate95inter5));
  nor2  gate2163(.a(gate95inter5), .b(gate95inter2), .O(gate95inter6));
  inv1  gate2164(.a(G26), .O(gate95inter7));
  inv1  gate2165(.a(G347), .O(gate95inter8));
  nand2 gate2166(.a(gate95inter8), .b(gate95inter7), .O(gate95inter9));
  nand2 gate2167(.a(s_231), .b(gate95inter3), .O(gate95inter10));
  nor2  gate2168(.a(gate95inter10), .b(gate95inter9), .O(gate95inter11));
  nor2  gate2169(.a(gate95inter11), .b(gate95inter6), .O(gate95inter12));
  nand2 gate2170(.a(gate95inter12), .b(gate95inter1), .O(G416));
nand2 gate96( .a(G30), .b(G347), .O(G417) );
nand2 gate97( .a(G19), .b(G350), .O(G418) );

  xor2  gate1163(.a(G350), .b(G23), .O(gate98inter0));
  nand2 gate1164(.a(gate98inter0), .b(s_88), .O(gate98inter1));
  and2  gate1165(.a(G350), .b(G23), .O(gate98inter2));
  inv1  gate1166(.a(s_88), .O(gate98inter3));
  inv1  gate1167(.a(s_89), .O(gate98inter4));
  nand2 gate1168(.a(gate98inter4), .b(gate98inter3), .O(gate98inter5));
  nor2  gate1169(.a(gate98inter5), .b(gate98inter2), .O(gate98inter6));
  inv1  gate1170(.a(G23), .O(gate98inter7));
  inv1  gate1171(.a(G350), .O(gate98inter8));
  nand2 gate1172(.a(gate98inter8), .b(gate98inter7), .O(gate98inter9));
  nand2 gate1173(.a(s_89), .b(gate98inter3), .O(gate98inter10));
  nor2  gate1174(.a(gate98inter10), .b(gate98inter9), .O(gate98inter11));
  nor2  gate1175(.a(gate98inter11), .b(gate98inter6), .O(gate98inter12));
  nand2 gate1176(.a(gate98inter12), .b(gate98inter1), .O(G419));
nand2 gate99( .a(G27), .b(G353), .O(G420) );
nand2 gate100( .a(G31), .b(G353), .O(G421) );

  xor2  gate883(.a(G356), .b(G20), .O(gate101inter0));
  nand2 gate884(.a(gate101inter0), .b(s_48), .O(gate101inter1));
  and2  gate885(.a(G356), .b(G20), .O(gate101inter2));
  inv1  gate886(.a(s_48), .O(gate101inter3));
  inv1  gate887(.a(s_49), .O(gate101inter4));
  nand2 gate888(.a(gate101inter4), .b(gate101inter3), .O(gate101inter5));
  nor2  gate889(.a(gate101inter5), .b(gate101inter2), .O(gate101inter6));
  inv1  gate890(.a(G20), .O(gate101inter7));
  inv1  gate891(.a(G356), .O(gate101inter8));
  nand2 gate892(.a(gate101inter8), .b(gate101inter7), .O(gate101inter9));
  nand2 gate893(.a(s_49), .b(gate101inter3), .O(gate101inter10));
  nor2  gate894(.a(gate101inter10), .b(gate101inter9), .O(gate101inter11));
  nor2  gate895(.a(gate101inter11), .b(gate101inter6), .O(gate101inter12));
  nand2 gate896(.a(gate101inter12), .b(gate101inter1), .O(G422));

  xor2  gate1513(.a(G356), .b(G24), .O(gate102inter0));
  nand2 gate1514(.a(gate102inter0), .b(s_138), .O(gate102inter1));
  and2  gate1515(.a(G356), .b(G24), .O(gate102inter2));
  inv1  gate1516(.a(s_138), .O(gate102inter3));
  inv1  gate1517(.a(s_139), .O(gate102inter4));
  nand2 gate1518(.a(gate102inter4), .b(gate102inter3), .O(gate102inter5));
  nor2  gate1519(.a(gate102inter5), .b(gate102inter2), .O(gate102inter6));
  inv1  gate1520(.a(G24), .O(gate102inter7));
  inv1  gate1521(.a(G356), .O(gate102inter8));
  nand2 gate1522(.a(gate102inter8), .b(gate102inter7), .O(gate102inter9));
  nand2 gate1523(.a(s_139), .b(gate102inter3), .O(gate102inter10));
  nor2  gate1524(.a(gate102inter10), .b(gate102inter9), .O(gate102inter11));
  nor2  gate1525(.a(gate102inter11), .b(gate102inter6), .O(gate102inter12));
  nand2 gate1526(.a(gate102inter12), .b(gate102inter1), .O(G423));

  xor2  gate1219(.a(G359), .b(G28), .O(gate103inter0));
  nand2 gate1220(.a(gate103inter0), .b(s_96), .O(gate103inter1));
  and2  gate1221(.a(G359), .b(G28), .O(gate103inter2));
  inv1  gate1222(.a(s_96), .O(gate103inter3));
  inv1  gate1223(.a(s_97), .O(gate103inter4));
  nand2 gate1224(.a(gate103inter4), .b(gate103inter3), .O(gate103inter5));
  nor2  gate1225(.a(gate103inter5), .b(gate103inter2), .O(gate103inter6));
  inv1  gate1226(.a(G28), .O(gate103inter7));
  inv1  gate1227(.a(G359), .O(gate103inter8));
  nand2 gate1228(.a(gate103inter8), .b(gate103inter7), .O(gate103inter9));
  nand2 gate1229(.a(s_97), .b(gate103inter3), .O(gate103inter10));
  nor2  gate1230(.a(gate103inter10), .b(gate103inter9), .O(gate103inter11));
  nor2  gate1231(.a(gate103inter11), .b(gate103inter6), .O(gate103inter12));
  nand2 gate1232(.a(gate103inter12), .b(gate103inter1), .O(G424));
nand2 gate104( .a(G32), .b(G359), .O(G425) );
nand2 gate105( .a(G362), .b(G363), .O(G426) );
nand2 gate106( .a(G364), .b(G365), .O(G429) );

  xor2  gate1611(.a(G367), .b(G366), .O(gate107inter0));
  nand2 gate1612(.a(gate107inter0), .b(s_152), .O(gate107inter1));
  and2  gate1613(.a(G367), .b(G366), .O(gate107inter2));
  inv1  gate1614(.a(s_152), .O(gate107inter3));
  inv1  gate1615(.a(s_153), .O(gate107inter4));
  nand2 gate1616(.a(gate107inter4), .b(gate107inter3), .O(gate107inter5));
  nor2  gate1617(.a(gate107inter5), .b(gate107inter2), .O(gate107inter6));
  inv1  gate1618(.a(G366), .O(gate107inter7));
  inv1  gate1619(.a(G367), .O(gate107inter8));
  nand2 gate1620(.a(gate107inter8), .b(gate107inter7), .O(gate107inter9));
  nand2 gate1621(.a(s_153), .b(gate107inter3), .O(gate107inter10));
  nor2  gate1622(.a(gate107inter10), .b(gate107inter9), .O(gate107inter11));
  nor2  gate1623(.a(gate107inter11), .b(gate107inter6), .O(gate107inter12));
  nand2 gate1624(.a(gate107inter12), .b(gate107inter1), .O(G432));
nand2 gate108( .a(G368), .b(G369), .O(G435) );
nand2 gate109( .a(G370), .b(G371), .O(G438) );

  xor2  gate1205(.a(G373), .b(G372), .O(gate110inter0));
  nand2 gate1206(.a(gate110inter0), .b(s_94), .O(gate110inter1));
  and2  gate1207(.a(G373), .b(G372), .O(gate110inter2));
  inv1  gate1208(.a(s_94), .O(gate110inter3));
  inv1  gate1209(.a(s_95), .O(gate110inter4));
  nand2 gate1210(.a(gate110inter4), .b(gate110inter3), .O(gate110inter5));
  nor2  gate1211(.a(gate110inter5), .b(gate110inter2), .O(gate110inter6));
  inv1  gate1212(.a(G372), .O(gate110inter7));
  inv1  gate1213(.a(G373), .O(gate110inter8));
  nand2 gate1214(.a(gate110inter8), .b(gate110inter7), .O(gate110inter9));
  nand2 gate1215(.a(s_95), .b(gate110inter3), .O(gate110inter10));
  nor2  gate1216(.a(gate110inter10), .b(gate110inter9), .O(gate110inter11));
  nor2  gate1217(.a(gate110inter11), .b(gate110inter6), .O(gate110inter12));
  nand2 gate1218(.a(gate110inter12), .b(gate110inter1), .O(G441));
nand2 gate111( .a(G374), .b(G375), .O(G444) );

  xor2  gate743(.a(G377), .b(G376), .O(gate112inter0));
  nand2 gate744(.a(gate112inter0), .b(s_28), .O(gate112inter1));
  and2  gate745(.a(G377), .b(G376), .O(gate112inter2));
  inv1  gate746(.a(s_28), .O(gate112inter3));
  inv1  gate747(.a(s_29), .O(gate112inter4));
  nand2 gate748(.a(gate112inter4), .b(gate112inter3), .O(gate112inter5));
  nor2  gate749(.a(gate112inter5), .b(gate112inter2), .O(gate112inter6));
  inv1  gate750(.a(G376), .O(gate112inter7));
  inv1  gate751(.a(G377), .O(gate112inter8));
  nand2 gate752(.a(gate112inter8), .b(gate112inter7), .O(gate112inter9));
  nand2 gate753(.a(s_29), .b(gate112inter3), .O(gate112inter10));
  nor2  gate754(.a(gate112inter10), .b(gate112inter9), .O(gate112inter11));
  nor2  gate755(.a(gate112inter11), .b(gate112inter6), .O(gate112inter12));
  nand2 gate756(.a(gate112inter12), .b(gate112inter1), .O(G447));

  xor2  gate1443(.a(G379), .b(G378), .O(gate113inter0));
  nand2 gate1444(.a(gate113inter0), .b(s_128), .O(gate113inter1));
  and2  gate1445(.a(G379), .b(G378), .O(gate113inter2));
  inv1  gate1446(.a(s_128), .O(gate113inter3));
  inv1  gate1447(.a(s_129), .O(gate113inter4));
  nand2 gate1448(.a(gate113inter4), .b(gate113inter3), .O(gate113inter5));
  nor2  gate1449(.a(gate113inter5), .b(gate113inter2), .O(gate113inter6));
  inv1  gate1450(.a(G378), .O(gate113inter7));
  inv1  gate1451(.a(G379), .O(gate113inter8));
  nand2 gate1452(.a(gate113inter8), .b(gate113inter7), .O(gate113inter9));
  nand2 gate1453(.a(s_129), .b(gate113inter3), .O(gate113inter10));
  nor2  gate1454(.a(gate113inter10), .b(gate113inter9), .O(gate113inter11));
  nor2  gate1455(.a(gate113inter11), .b(gate113inter6), .O(gate113inter12));
  nand2 gate1456(.a(gate113inter12), .b(gate113inter1), .O(G450));
nand2 gate114( .a(G380), .b(G381), .O(G453) );
nand2 gate115( .a(G382), .b(G383), .O(G456) );
nand2 gate116( .a(G384), .b(G385), .O(G459) );
nand2 gate117( .a(G386), .b(G387), .O(G462) );
nand2 gate118( .a(G388), .b(G389), .O(G465) );

  xor2  gate2241(.a(G391), .b(G390), .O(gate119inter0));
  nand2 gate2242(.a(gate119inter0), .b(s_242), .O(gate119inter1));
  and2  gate2243(.a(G391), .b(G390), .O(gate119inter2));
  inv1  gate2244(.a(s_242), .O(gate119inter3));
  inv1  gate2245(.a(s_243), .O(gate119inter4));
  nand2 gate2246(.a(gate119inter4), .b(gate119inter3), .O(gate119inter5));
  nor2  gate2247(.a(gate119inter5), .b(gate119inter2), .O(gate119inter6));
  inv1  gate2248(.a(G390), .O(gate119inter7));
  inv1  gate2249(.a(G391), .O(gate119inter8));
  nand2 gate2250(.a(gate119inter8), .b(gate119inter7), .O(gate119inter9));
  nand2 gate2251(.a(s_243), .b(gate119inter3), .O(gate119inter10));
  nor2  gate2252(.a(gate119inter10), .b(gate119inter9), .O(gate119inter11));
  nor2  gate2253(.a(gate119inter11), .b(gate119inter6), .O(gate119inter12));
  nand2 gate2254(.a(gate119inter12), .b(gate119inter1), .O(G468));

  xor2  gate2213(.a(G393), .b(G392), .O(gate120inter0));
  nand2 gate2214(.a(gate120inter0), .b(s_238), .O(gate120inter1));
  and2  gate2215(.a(G393), .b(G392), .O(gate120inter2));
  inv1  gate2216(.a(s_238), .O(gate120inter3));
  inv1  gate2217(.a(s_239), .O(gate120inter4));
  nand2 gate2218(.a(gate120inter4), .b(gate120inter3), .O(gate120inter5));
  nor2  gate2219(.a(gate120inter5), .b(gate120inter2), .O(gate120inter6));
  inv1  gate2220(.a(G392), .O(gate120inter7));
  inv1  gate2221(.a(G393), .O(gate120inter8));
  nand2 gate2222(.a(gate120inter8), .b(gate120inter7), .O(gate120inter9));
  nand2 gate2223(.a(s_239), .b(gate120inter3), .O(gate120inter10));
  nor2  gate2224(.a(gate120inter10), .b(gate120inter9), .O(gate120inter11));
  nor2  gate2225(.a(gate120inter11), .b(gate120inter6), .O(gate120inter12));
  nand2 gate2226(.a(gate120inter12), .b(gate120inter1), .O(G471));
nand2 gate121( .a(G394), .b(G395), .O(G474) );

  xor2  gate1723(.a(G397), .b(G396), .O(gate122inter0));
  nand2 gate1724(.a(gate122inter0), .b(s_168), .O(gate122inter1));
  and2  gate1725(.a(G397), .b(G396), .O(gate122inter2));
  inv1  gate1726(.a(s_168), .O(gate122inter3));
  inv1  gate1727(.a(s_169), .O(gate122inter4));
  nand2 gate1728(.a(gate122inter4), .b(gate122inter3), .O(gate122inter5));
  nor2  gate1729(.a(gate122inter5), .b(gate122inter2), .O(gate122inter6));
  inv1  gate1730(.a(G396), .O(gate122inter7));
  inv1  gate1731(.a(G397), .O(gate122inter8));
  nand2 gate1732(.a(gate122inter8), .b(gate122inter7), .O(gate122inter9));
  nand2 gate1733(.a(s_169), .b(gate122inter3), .O(gate122inter10));
  nor2  gate1734(.a(gate122inter10), .b(gate122inter9), .O(gate122inter11));
  nor2  gate1735(.a(gate122inter11), .b(gate122inter6), .O(gate122inter12));
  nand2 gate1736(.a(gate122inter12), .b(gate122inter1), .O(G477));
nand2 gate123( .a(G398), .b(G399), .O(G480) );
nand2 gate124( .a(G400), .b(G401), .O(G483) );

  xor2  gate1821(.a(G403), .b(G402), .O(gate125inter0));
  nand2 gate1822(.a(gate125inter0), .b(s_182), .O(gate125inter1));
  and2  gate1823(.a(G403), .b(G402), .O(gate125inter2));
  inv1  gate1824(.a(s_182), .O(gate125inter3));
  inv1  gate1825(.a(s_183), .O(gate125inter4));
  nand2 gate1826(.a(gate125inter4), .b(gate125inter3), .O(gate125inter5));
  nor2  gate1827(.a(gate125inter5), .b(gate125inter2), .O(gate125inter6));
  inv1  gate1828(.a(G402), .O(gate125inter7));
  inv1  gate1829(.a(G403), .O(gate125inter8));
  nand2 gate1830(.a(gate125inter8), .b(gate125inter7), .O(gate125inter9));
  nand2 gate1831(.a(s_183), .b(gate125inter3), .O(gate125inter10));
  nor2  gate1832(.a(gate125inter10), .b(gate125inter9), .O(gate125inter11));
  nor2  gate1833(.a(gate125inter11), .b(gate125inter6), .O(gate125inter12));
  nand2 gate1834(.a(gate125inter12), .b(gate125inter1), .O(G486));
nand2 gate126( .a(G404), .b(G405), .O(G489) );
nand2 gate127( .a(G406), .b(G407), .O(G492) );
nand2 gate128( .a(G408), .b(G409), .O(G495) );
nand2 gate129( .a(G410), .b(G411), .O(G498) );
nand2 gate130( .a(G412), .b(G413), .O(G501) );
nand2 gate131( .a(G414), .b(G415), .O(G504) );

  xor2  gate1639(.a(G417), .b(G416), .O(gate132inter0));
  nand2 gate1640(.a(gate132inter0), .b(s_156), .O(gate132inter1));
  and2  gate1641(.a(G417), .b(G416), .O(gate132inter2));
  inv1  gate1642(.a(s_156), .O(gate132inter3));
  inv1  gate1643(.a(s_157), .O(gate132inter4));
  nand2 gate1644(.a(gate132inter4), .b(gate132inter3), .O(gate132inter5));
  nor2  gate1645(.a(gate132inter5), .b(gate132inter2), .O(gate132inter6));
  inv1  gate1646(.a(G416), .O(gate132inter7));
  inv1  gate1647(.a(G417), .O(gate132inter8));
  nand2 gate1648(.a(gate132inter8), .b(gate132inter7), .O(gate132inter9));
  nand2 gate1649(.a(s_157), .b(gate132inter3), .O(gate132inter10));
  nor2  gate1650(.a(gate132inter10), .b(gate132inter9), .O(gate132inter11));
  nor2  gate1651(.a(gate132inter11), .b(gate132inter6), .O(gate132inter12));
  nand2 gate1652(.a(gate132inter12), .b(gate132inter1), .O(G507));

  xor2  gate2059(.a(G419), .b(G418), .O(gate133inter0));
  nand2 gate2060(.a(gate133inter0), .b(s_216), .O(gate133inter1));
  and2  gate2061(.a(G419), .b(G418), .O(gate133inter2));
  inv1  gate2062(.a(s_216), .O(gate133inter3));
  inv1  gate2063(.a(s_217), .O(gate133inter4));
  nand2 gate2064(.a(gate133inter4), .b(gate133inter3), .O(gate133inter5));
  nor2  gate2065(.a(gate133inter5), .b(gate133inter2), .O(gate133inter6));
  inv1  gate2066(.a(G418), .O(gate133inter7));
  inv1  gate2067(.a(G419), .O(gate133inter8));
  nand2 gate2068(.a(gate133inter8), .b(gate133inter7), .O(gate133inter9));
  nand2 gate2069(.a(s_217), .b(gate133inter3), .O(gate133inter10));
  nor2  gate2070(.a(gate133inter10), .b(gate133inter9), .O(gate133inter11));
  nor2  gate2071(.a(gate133inter11), .b(gate133inter6), .O(gate133inter12));
  nand2 gate2072(.a(gate133inter12), .b(gate133inter1), .O(G510));
nand2 gate134( .a(G420), .b(G421), .O(G513) );

  xor2  gate771(.a(G423), .b(G422), .O(gate135inter0));
  nand2 gate772(.a(gate135inter0), .b(s_32), .O(gate135inter1));
  and2  gate773(.a(G423), .b(G422), .O(gate135inter2));
  inv1  gate774(.a(s_32), .O(gate135inter3));
  inv1  gate775(.a(s_33), .O(gate135inter4));
  nand2 gate776(.a(gate135inter4), .b(gate135inter3), .O(gate135inter5));
  nor2  gate777(.a(gate135inter5), .b(gate135inter2), .O(gate135inter6));
  inv1  gate778(.a(G422), .O(gate135inter7));
  inv1  gate779(.a(G423), .O(gate135inter8));
  nand2 gate780(.a(gate135inter8), .b(gate135inter7), .O(gate135inter9));
  nand2 gate781(.a(s_33), .b(gate135inter3), .O(gate135inter10));
  nor2  gate782(.a(gate135inter10), .b(gate135inter9), .O(gate135inter11));
  nor2  gate783(.a(gate135inter11), .b(gate135inter6), .O(gate135inter12));
  nand2 gate784(.a(gate135inter12), .b(gate135inter1), .O(G516));
nand2 gate136( .a(G424), .b(G425), .O(G519) );
nand2 gate137( .a(G426), .b(G429), .O(G522) );

  xor2  gate2283(.a(G435), .b(G432), .O(gate138inter0));
  nand2 gate2284(.a(gate138inter0), .b(s_248), .O(gate138inter1));
  and2  gate2285(.a(G435), .b(G432), .O(gate138inter2));
  inv1  gate2286(.a(s_248), .O(gate138inter3));
  inv1  gate2287(.a(s_249), .O(gate138inter4));
  nand2 gate2288(.a(gate138inter4), .b(gate138inter3), .O(gate138inter5));
  nor2  gate2289(.a(gate138inter5), .b(gate138inter2), .O(gate138inter6));
  inv1  gate2290(.a(G432), .O(gate138inter7));
  inv1  gate2291(.a(G435), .O(gate138inter8));
  nand2 gate2292(.a(gate138inter8), .b(gate138inter7), .O(gate138inter9));
  nand2 gate2293(.a(s_249), .b(gate138inter3), .O(gate138inter10));
  nor2  gate2294(.a(gate138inter10), .b(gate138inter9), .O(gate138inter11));
  nor2  gate2295(.a(gate138inter11), .b(gate138inter6), .O(gate138inter12));
  nand2 gate2296(.a(gate138inter12), .b(gate138inter1), .O(G525));
nand2 gate139( .a(G438), .b(G441), .O(G528) );
nand2 gate140( .a(G444), .b(G447), .O(G531) );
nand2 gate141( .a(G450), .b(G453), .O(G534) );
nand2 gate142( .a(G456), .b(G459), .O(G537) );
nand2 gate143( .a(G462), .b(G465), .O(G540) );

  xor2  gate2087(.a(G471), .b(G468), .O(gate144inter0));
  nand2 gate2088(.a(gate144inter0), .b(s_220), .O(gate144inter1));
  and2  gate2089(.a(G471), .b(G468), .O(gate144inter2));
  inv1  gate2090(.a(s_220), .O(gate144inter3));
  inv1  gate2091(.a(s_221), .O(gate144inter4));
  nand2 gate2092(.a(gate144inter4), .b(gate144inter3), .O(gate144inter5));
  nor2  gate2093(.a(gate144inter5), .b(gate144inter2), .O(gate144inter6));
  inv1  gate2094(.a(G468), .O(gate144inter7));
  inv1  gate2095(.a(G471), .O(gate144inter8));
  nand2 gate2096(.a(gate144inter8), .b(gate144inter7), .O(gate144inter9));
  nand2 gate2097(.a(s_221), .b(gate144inter3), .O(gate144inter10));
  nor2  gate2098(.a(gate144inter10), .b(gate144inter9), .O(gate144inter11));
  nor2  gate2099(.a(gate144inter11), .b(gate144inter6), .O(gate144inter12));
  nand2 gate2100(.a(gate144inter12), .b(gate144inter1), .O(G543));
nand2 gate145( .a(G474), .b(G477), .O(G546) );
nand2 gate146( .a(G480), .b(G483), .O(G549) );

  xor2  gate631(.a(G489), .b(G486), .O(gate147inter0));
  nand2 gate632(.a(gate147inter0), .b(s_12), .O(gate147inter1));
  and2  gate633(.a(G489), .b(G486), .O(gate147inter2));
  inv1  gate634(.a(s_12), .O(gate147inter3));
  inv1  gate635(.a(s_13), .O(gate147inter4));
  nand2 gate636(.a(gate147inter4), .b(gate147inter3), .O(gate147inter5));
  nor2  gate637(.a(gate147inter5), .b(gate147inter2), .O(gate147inter6));
  inv1  gate638(.a(G486), .O(gate147inter7));
  inv1  gate639(.a(G489), .O(gate147inter8));
  nand2 gate640(.a(gate147inter8), .b(gate147inter7), .O(gate147inter9));
  nand2 gate641(.a(s_13), .b(gate147inter3), .O(gate147inter10));
  nor2  gate642(.a(gate147inter10), .b(gate147inter9), .O(gate147inter11));
  nor2  gate643(.a(gate147inter11), .b(gate147inter6), .O(gate147inter12));
  nand2 gate644(.a(gate147inter12), .b(gate147inter1), .O(G552));
nand2 gate148( .a(G492), .b(G495), .O(G555) );
nand2 gate149( .a(G498), .b(G501), .O(G558) );
nand2 gate150( .a(G504), .b(G507), .O(G561) );

  xor2  gate1989(.a(G513), .b(G510), .O(gate151inter0));
  nand2 gate1990(.a(gate151inter0), .b(s_206), .O(gate151inter1));
  and2  gate1991(.a(G513), .b(G510), .O(gate151inter2));
  inv1  gate1992(.a(s_206), .O(gate151inter3));
  inv1  gate1993(.a(s_207), .O(gate151inter4));
  nand2 gate1994(.a(gate151inter4), .b(gate151inter3), .O(gate151inter5));
  nor2  gate1995(.a(gate151inter5), .b(gate151inter2), .O(gate151inter6));
  inv1  gate1996(.a(G510), .O(gate151inter7));
  inv1  gate1997(.a(G513), .O(gate151inter8));
  nand2 gate1998(.a(gate151inter8), .b(gate151inter7), .O(gate151inter9));
  nand2 gate1999(.a(s_207), .b(gate151inter3), .O(gate151inter10));
  nor2  gate2000(.a(gate151inter10), .b(gate151inter9), .O(gate151inter11));
  nor2  gate2001(.a(gate151inter11), .b(gate151inter6), .O(gate151inter12));
  nand2 gate2002(.a(gate151inter12), .b(gate151inter1), .O(G564));

  xor2  gate2339(.a(G519), .b(G516), .O(gate152inter0));
  nand2 gate2340(.a(gate152inter0), .b(s_256), .O(gate152inter1));
  and2  gate2341(.a(G519), .b(G516), .O(gate152inter2));
  inv1  gate2342(.a(s_256), .O(gate152inter3));
  inv1  gate2343(.a(s_257), .O(gate152inter4));
  nand2 gate2344(.a(gate152inter4), .b(gate152inter3), .O(gate152inter5));
  nor2  gate2345(.a(gate152inter5), .b(gate152inter2), .O(gate152inter6));
  inv1  gate2346(.a(G516), .O(gate152inter7));
  inv1  gate2347(.a(G519), .O(gate152inter8));
  nand2 gate2348(.a(gate152inter8), .b(gate152inter7), .O(gate152inter9));
  nand2 gate2349(.a(s_257), .b(gate152inter3), .O(gate152inter10));
  nor2  gate2350(.a(gate152inter10), .b(gate152inter9), .O(gate152inter11));
  nor2  gate2351(.a(gate152inter11), .b(gate152inter6), .O(gate152inter12));
  nand2 gate2352(.a(gate152inter12), .b(gate152inter1), .O(G567));
nand2 gate153( .a(G426), .b(G522), .O(G570) );
nand2 gate154( .a(G429), .b(G522), .O(G571) );

  xor2  gate2409(.a(G525), .b(G432), .O(gate155inter0));
  nand2 gate2410(.a(gate155inter0), .b(s_266), .O(gate155inter1));
  and2  gate2411(.a(G525), .b(G432), .O(gate155inter2));
  inv1  gate2412(.a(s_266), .O(gate155inter3));
  inv1  gate2413(.a(s_267), .O(gate155inter4));
  nand2 gate2414(.a(gate155inter4), .b(gate155inter3), .O(gate155inter5));
  nor2  gate2415(.a(gate155inter5), .b(gate155inter2), .O(gate155inter6));
  inv1  gate2416(.a(G432), .O(gate155inter7));
  inv1  gate2417(.a(G525), .O(gate155inter8));
  nand2 gate2418(.a(gate155inter8), .b(gate155inter7), .O(gate155inter9));
  nand2 gate2419(.a(s_267), .b(gate155inter3), .O(gate155inter10));
  nor2  gate2420(.a(gate155inter10), .b(gate155inter9), .O(gate155inter11));
  nor2  gate2421(.a(gate155inter11), .b(gate155inter6), .O(gate155inter12));
  nand2 gate2422(.a(gate155inter12), .b(gate155inter1), .O(G572));

  xor2  gate1149(.a(G525), .b(G435), .O(gate156inter0));
  nand2 gate1150(.a(gate156inter0), .b(s_86), .O(gate156inter1));
  and2  gate1151(.a(G525), .b(G435), .O(gate156inter2));
  inv1  gate1152(.a(s_86), .O(gate156inter3));
  inv1  gate1153(.a(s_87), .O(gate156inter4));
  nand2 gate1154(.a(gate156inter4), .b(gate156inter3), .O(gate156inter5));
  nor2  gate1155(.a(gate156inter5), .b(gate156inter2), .O(gate156inter6));
  inv1  gate1156(.a(G435), .O(gate156inter7));
  inv1  gate1157(.a(G525), .O(gate156inter8));
  nand2 gate1158(.a(gate156inter8), .b(gate156inter7), .O(gate156inter9));
  nand2 gate1159(.a(s_87), .b(gate156inter3), .O(gate156inter10));
  nor2  gate1160(.a(gate156inter10), .b(gate156inter9), .O(gate156inter11));
  nor2  gate1161(.a(gate156inter11), .b(gate156inter6), .O(gate156inter12));
  nand2 gate1162(.a(gate156inter12), .b(gate156inter1), .O(G573));

  xor2  gate2297(.a(G528), .b(G438), .O(gate157inter0));
  nand2 gate2298(.a(gate157inter0), .b(s_250), .O(gate157inter1));
  and2  gate2299(.a(G528), .b(G438), .O(gate157inter2));
  inv1  gate2300(.a(s_250), .O(gate157inter3));
  inv1  gate2301(.a(s_251), .O(gate157inter4));
  nand2 gate2302(.a(gate157inter4), .b(gate157inter3), .O(gate157inter5));
  nor2  gate2303(.a(gate157inter5), .b(gate157inter2), .O(gate157inter6));
  inv1  gate2304(.a(G438), .O(gate157inter7));
  inv1  gate2305(.a(G528), .O(gate157inter8));
  nand2 gate2306(.a(gate157inter8), .b(gate157inter7), .O(gate157inter9));
  nand2 gate2307(.a(s_251), .b(gate157inter3), .O(gate157inter10));
  nor2  gate2308(.a(gate157inter10), .b(gate157inter9), .O(gate157inter11));
  nor2  gate2309(.a(gate157inter11), .b(gate157inter6), .O(gate157inter12));
  nand2 gate2310(.a(gate157inter12), .b(gate157inter1), .O(G574));
nand2 gate158( .a(G441), .b(G528), .O(G575) );
nand2 gate159( .a(G444), .b(G531), .O(G576) );
nand2 gate160( .a(G447), .b(G531), .O(G577) );
nand2 gate161( .a(G450), .b(G534), .O(G578) );

  xor2  gate981(.a(G534), .b(G453), .O(gate162inter0));
  nand2 gate982(.a(gate162inter0), .b(s_62), .O(gate162inter1));
  and2  gate983(.a(G534), .b(G453), .O(gate162inter2));
  inv1  gate984(.a(s_62), .O(gate162inter3));
  inv1  gate985(.a(s_63), .O(gate162inter4));
  nand2 gate986(.a(gate162inter4), .b(gate162inter3), .O(gate162inter5));
  nor2  gate987(.a(gate162inter5), .b(gate162inter2), .O(gate162inter6));
  inv1  gate988(.a(G453), .O(gate162inter7));
  inv1  gate989(.a(G534), .O(gate162inter8));
  nand2 gate990(.a(gate162inter8), .b(gate162inter7), .O(gate162inter9));
  nand2 gate991(.a(s_63), .b(gate162inter3), .O(gate162inter10));
  nor2  gate992(.a(gate162inter10), .b(gate162inter9), .O(gate162inter11));
  nor2  gate993(.a(gate162inter11), .b(gate162inter6), .O(gate162inter12));
  nand2 gate994(.a(gate162inter12), .b(gate162inter1), .O(G579));

  xor2  gate2353(.a(G537), .b(G456), .O(gate163inter0));
  nand2 gate2354(.a(gate163inter0), .b(s_258), .O(gate163inter1));
  and2  gate2355(.a(G537), .b(G456), .O(gate163inter2));
  inv1  gate2356(.a(s_258), .O(gate163inter3));
  inv1  gate2357(.a(s_259), .O(gate163inter4));
  nand2 gate2358(.a(gate163inter4), .b(gate163inter3), .O(gate163inter5));
  nor2  gate2359(.a(gate163inter5), .b(gate163inter2), .O(gate163inter6));
  inv1  gate2360(.a(G456), .O(gate163inter7));
  inv1  gate2361(.a(G537), .O(gate163inter8));
  nand2 gate2362(.a(gate163inter8), .b(gate163inter7), .O(gate163inter9));
  nand2 gate2363(.a(s_259), .b(gate163inter3), .O(gate163inter10));
  nor2  gate2364(.a(gate163inter10), .b(gate163inter9), .O(gate163inter11));
  nor2  gate2365(.a(gate163inter11), .b(gate163inter6), .O(gate163inter12));
  nand2 gate2366(.a(gate163inter12), .b(gate163inter1), .O(G580));
nand2 gate164( .a(G459), .b(G537), .O(G581) );
nand2 gate165( .a(G462), .b(G540), .O(G582) );

  xor2  gate1681(.a(G540), .b(G465), .O(gate166inter0));
  nand2 gate1682(.a(gate166inter0), .b(s_162), .O(gate166inter1));
  and2  gate1683(.a(G540), .b(G465), .O(gate166inter2));
  inv1  gate1684(.a(s_162), .O(gate166inter3));
  inv1  gate1685(.a(s_163), .O(gate166inter4));
  nand2 gate1686(.a(gate166inter4), .b(gate166inter3), .O(gate166inter5));
  nor2  gate1687(.a(gate166inter5), .b(gate166inter2), .O(gate166inter6));
  inv1  gate1688(.a(G465), .O(gate166inter7));
  inv1  gate1689(.a(G540), .O(gate166inter8));
  nand2 gate1690(.a(gate166inter8), .b(gate166inter7), .O(gate166inter9));
  nand2 gate1691(.a(s_163), .b(gate166inter3), .O(gate166inter10));
  nor2  gate1692(.a(gate166inter10), .b(gate166inter9), .O(gate166inter11));
  nor2  gate1693(.a(gate166inter11), .b(gate166inter6), .O(gate166inter12));
  nand2 gate1694(.a(gate166inter12), .b(gate166inter1), .O(G583));

  xor2  gate2171(.a(G543), .b(G468), .O(gate167inter0));
  nand2 gate2172(.a(gate167inter0), .b(s_232), .O(gate167inter1));
  and2  gate2173(.a(G543), .b(G468), .O(gate167inter2));
  inv1  gate2174(.a(s_232), .O(gate167inter3));
  inv1  gate2175(.a(s_233), .O(gate167inter4));
  nand2 gate2176(.a(gate167inter4), .b(gate167inter3), .O(gate167inter5));
  nor2  gate2177(.a(gate167inter5), .b(gate167inter2), .O(gate167inter6));
  inv1  gate2178(.a(G468), .O(gate167inter7));
  inv1  gate2179(.a(G543), .O(gate167inter8));
  nand2 gate2180(.a(gate167inter8), .b(gate167inter7), .O(gate167inter9));
  nand2 gate2181(.a(s_233), .b(gate167inter3), .O(gate167inter10));
  nor2  gate2182(.a(gate167inter10), .b(gate167inter9), .O(gate167inter11));
  nor2  gate2183(.a(gate167inter11), .b(gate167inter6), .O(gate167inter12));
  nand2 gate2184(.a(gate167inter12), .b(gate167inter1), .O(G584));
nand2 gate168( .a(G471), .b(G543), .O(G585) );
nand2 gate169( .a(G474), .b(G546), .O(G586) );
nand2 gate170( .a(G477), .b(G546), .O(G587) );

  xor2  gate1415(.a(G549), .b(G480), .O(gate171inter0));
  nand2 gate1416(.a(gate171inter0), .b(s_124), .O(gate171inter1));
  and2  gate1417(.a(G549), .b(G480), .O(gate171inter2));
  inv1  gate1418(.a(s_124), .O(gate171inter3));
  inv1  gate1419(.a(s_125), .O(gate171inter4));
  nand2 gate1420(.a(gate171inter4), .b(gate171inter3), .O(gate171inter5));
  nor2  gate1421(.a(gate171inter5), .b(gate171inter2), .O(gate171inter6));
  inv1  gate1422(.a(G480), .O(gate171inter7));
  inv1  gate1423(.a(G549), .O(gate171inter8));
  nand2 gate1424(.a(gate171inter8), .b(gate171inter7), .O(gate171inter9));
  nand2 gate1425(.a(s_125), .b(gate171inter3), .O(gate171inter10));
  nor2  gate1426(.a(gate171inter10), .b(gate171inter9), .O(gate171inter11));
  nor2  gate1427(.a(gate171inter11), .b(gate171inter6), .O(gate171inter12));
  nand2 gate1428(.a(gate171inter12), .b(gate171inter1), .O(G588));

  xor2  gate1737(.a(G549), .b(G483), .O(gate172inter0));
  nand2 gate1738(.a(gate172inter0), .b(s_170), .O(gate172inter1));
  and2  gate1739(.a(G549), .b(G483), .O(gate172inter2));
  inv1  gate1740(.a(s_170), .O(gate172inter3));
  inv1  gate1741(.a(s_171), .O(gate172inter4));
  nand2 gate1742(.a(gate172inter4), .b(gate172inter3), .O(gate172inter5));
  nor2  gate1743(.a(gate172inter5), .b(gate172inter2), .O(gate172inter6));
  inv1  gate1744(.a(G483), .O(gate172inter7));
  inv1  gate1745(.a(G549), .O(gate172inter8));
  nand2 gate1746(.a(gate172inter8), .b(gate172inter7), .O(gate172inter9));
  nand2 gate1747(.a(s_171), .b(gate172inter3), .O(gate172inter10));
  nor2  gate1748(.a(gate172inter10), .b(gate172inter9), .O(gate172inter11));
  nor2  gate1749(.a(gate172inter11), .b(gate172inter6), .O(gate172inter12));
  nand2 gate1750(.a(gate172inter12), .b(gate172inter1), .O(G589));
nand2 gate173( .a(G486), .b(G552), .O(G590) );
nand2 gate174( .a(G489), .b(G552), .O(G591) );
nand2 gate175( .a(G492), .b(G555), .O(G592) );
nand2 gate176( .a(G495), .b(G555), .O(G593) );
nand2 gate177( .a(G498), .b(G558), .O(G594) );
nand2 gate178( .a(G501), .b(G558), .O(G595) );
nand2 gate179( .a(G504), .b(G561), .O(G596) );

  xor2  gate1793(.a(G561), .b(G507), .O(gate180inter0));
  nand2 gate1794(.a(gate180inter0), .b(s_178), .O(gate180inter1));
  and2  gate1795(.a(G561), .b(G507), .O(gate180inter2));
  inv1  gate1796(.a(s_178), .O(gate180inter3));
  inv1  gate1797(.a(s_179), .O(gate180inter4));
  nand2 gate1798(.a(gate180inter4), .b(gate180inter3), .O(gate180inter5));
  nor2  gate1799(.a(gate180inter5), .b(gate180inter2), .O(gate180inter6));
  inv1  gate1800(.a(G507), .O(gate180inter7));
  inv1  gate1801(.a(G561), .O(gate180inter8));
  nand2 gate1802(.a(gate180inter8), .b(gate180inter7), .O(gate180inter9));
  nand2 gate1803(.a(s_179), .b(gate180inter3), .O(gate180inter10));
  nor2  gate1804(.a(gate180inter10), .b(gate180inter9), .O(gate180inter11));
  nor2  gate1805(.a(gate180inter11), .b(gate180inter6), .O(gate180inter12));
  nand2 gate1806(.a(gate180inter12), .b(gate180inter1), .O(G597));

  xor2  gate841(.a(G564), .b(G510), .O(gate181inter0));
  nand2 gate842(.a(gate181inter0), .b(s_42), .O(gate181inter1));
  and2  gate843(.a(G564), .b(G510), .O(gate181inter2));
  inv1  gate844(.a(s_42), .O(gate181inter3));
  inv1  gate845(.a(s_43), .O(gate181inter4));
  nand2 gate846(.a(gate181inter4), .b(gate181inter3), .O(gate181inter5));
  nor2  gate847(.a(gate181inter5), .b(gate181inter2), .O(gate181inter6));
  inv1  gate848(.a(G510), .O(gate181inter7));
  inv1  gate849(.a(G564), .O(gate181inter8));
  nand2 gate850(.a(gate181inter8), .b(gate181inter7), .O(gate181inter9));
  nand2 gate851(.a(s_43), .b(gate181inter3), .O(gate181inter10));
  nor2  gate852(.a(gate181inter10), .b(gate181inter9), .O(gate181inter11));
  nor2  gate853(.a(gate181inter11), .b(gate181inter6), .O(gate181inter12));
  nand2 gate854(.a(gate181inter12), .b(gate181inter1), .O(G598));
nand2 gate182( .a(G513), .b(G564), .O(G599) );
nand2 gate183( .a(G516), .b(G567), .O(G600) );

  xor2  gate673(.a(G567), .b(G519), .O(gate184inter0));
  nand2 gate674(.a(gate184inter0), .b(s_18), .O(gate184inter1));
  and2  gate675(.a(G567), .b(G519), .O(gate184inter2));
  inv1  gate676(.a(s_18), .O(gate184inter3));
  inv1  gate677(.a(s_19), .O(gate184inter4));
  nand2 gate678(.a(gate184inter4), .b(gate184inter3), .O(gate184inter5));
  nor2  gate679(.a(gate184inter5), .b(gate184inter2), .O(gate184inter6));
  inv1  gate680(.a(G519), .O(gate184inter7));
  inv1  gate681(.a(G567), .O(gate184inter8));
  nand2 gate682(.a(gate184inter8), .b(gate184inter7), .O(gate184inter9));
  nand2 gate683(.a(s_19), .b(gate184inter3), .O(gate184inter10));
  nor2  gate684(.a(gate184inter10), .b(gate184inter9), .O(gate184inter11));
  nor2  gate685(.a(gate184inter11), .b(gate184inter6), .O(gate184inter12));
  nand2 gate686(.a(gate184inter12), .b(gate184inter1), .O(G601));

  xor2  gate1891(.a(G571), .b(G570), .O(gate185inter0));
  nand2 gate1892(.a(gate185inter0), .b(s_192), .O(gate185inter1));
  and2  gate1893(.a(G571), .b(G570), .O(gate185inter2));
  inv1  gate1894(.a(s_192), .O(gate185inter3));
  inv1  gate1895(.a(s_193), .O(gate185inter4));
  nand2 gate1896(.a(gate185inter4), .b(gate185inter3), .O(gate185inter5));
  nor2  gate1897(.a(gate185inter5), .b(gate185inter2), .O(gate185inter6));
  inv1  gate1898(.a(G570), .O(gate185inter7));
  inv1  gate1899(.a(G571), .O(gate185inter8));
  nand2 gate1900(.a(gate185inter8), .b(gate185inter7), .O(gate185inter9));
  nand2 gate1901(.a(s_193), .b(gate185inter3), .O(gate185inter10));
  nor2  gate1902(.a(gate185inter10), .b(gate185inter9), .O(gate185inter11));
  nor2  gate1903(.a(gate185inter11), .b(gate185inter6), .O(gate185inter12));
  nand2 gate1904(.a(gate185inter12), .b(gate185inter1), .O(G602));

  xor2  gate1499(.a(G573), .b(G572), .O(gate186inter0));
  nand2 gate1500(.a(gate186inter0), .b(s_136), .O(gate186inter1));
  and2  gate1501(.a(G573), .b(G572), .O(gate186inter2));
  inv1  gate1502(.a(s_136), .O(gate186inter3));
  inv1  gate1503(.a(s_137), .O(gate186inter4));
  nand2 gate1504(.a(gate186inter4), .b(gate186inter3), .O(gate186inter5));
  nor2  gate1505(.a(gate186inter5), .b(gate186inter2), .O(gate186inter6));
  inv1  gate1506(.a(G572), .O(gate186inter7));
  inv1  gate1507(.a(G573), .O(gate186inter8));
  nand2 gate1508(.a(gate186inter8), .b(gate186inter7), .O(gate186inter9));
  nand2 gate1509(.a(s_137), .b(gate186inter3), .O(gate186inter10));
  nor2  gate1510(.a(gate186inter10), .b(gate186inter9), .O(gate186inter11));
  nor2  gate1511(.a(gate186inter11), .b(gate186inter6), .O(gate186inter12));
  nand2 gate1512(.a(gate186inter12), .b(gate186inter1), .O(G607));
nand2 gate187( .a(G574), .b(G575), .O(G612) );
nand2 gate188( .a(G576), .b(G577), .O(G617) );
nand2 gate189( .a(G578), .b(G579), .O(G622) );
nand2 gate190( .a(G580), .b(G581), .O(G627) );
nand2 gate191( .a(G582), .b(G583), .O(G632) );

  xor2  gate2199(.a(G585), .b(G584), .O(gate192inter0));
  nand2 gate2200(.a(gate192inter0), .b(s_236), .O(gate192inter1));
  and2  gate2201(.a(G585), .b(G584), .O(gate192inter2));
  inv1  gate2202(.a(s_236), .O(gate192inter3));
  inv1  gate2203(.a(s_237), .O(gate192inter4));
  nand2 gate2204(.a(gate192inter4), .b(gate192inter3), .O(gate192inter5));
  nor2  gate2205(.a(gate192inter5), .b(gate192inter2), .O(gate192inter6));
  inv1  gate2206(.a(G584), .O(gate192inter7));
  inv1  gate2207(.a(G585), .O(gate192inter8));
  nand2 gate2208(.a(gate192inter8), .b(gate192inter7), .O(gate192inter9));
  nand2 gate2209(.a(s_237), .b(gate192inter3), .O(gate192inter10));
  nor2  gate2210(.a(gate192inter10), .b(gate192inter9), .O(gate192inter11));
  nor2  gate2211(.a(gate192inter11), .b(gate192inter6), .O(gate192inter12));
  nand2 gate2212(.a(gate192inter12), .b(gate192inter1), .O(G637));
nand2 gate193( .a(G586), .b(G587), .O(G642) );
nand2 gate194( .a(G588), .b(G589), .O(G645) );
nand2 gate195( .a(G590), .b(G591), .O(G648) );
nand2 gate196( .a(G592), .b(G593), .O(G651) );
nand2 gate197( .a(G594), .b(G595), .O(G654) );
nand2 gate198( .a(G596), .b(G597), .O(G657) );
nand2 gate199( .a(G598), .b(G599), .O(G660) );

  xor2  gate1093(.a(G601), .b(G600), .O(gate200inter0));
  nand2 gate1094(.a(gate200inter0), .b(s_78), .O(gate200inter1));
  and2  gate1095(.a(G601), .b(G600), .O(gate200inter2));
  inv1  gate1096(.a(s_78), .O(gate200inter3));
  inv1  gate1097(.a(s_79), .O(gate200inter4));
  nand2 gate1098(.a(gate200inter4), .b(gate200inter3), .O(gate200inter5));
  nor2  gate1099(.a(gate200inter5), .b(gate200inter2), .O(gate200inter6));
  inv1  gate1100(.a(G600), .O(gate200inter7));
  inv1  gate1101(.a(G601), .O(gate200inter8));
  nand2 gate1102(.a(gate200inter8), .b(gate200inter7), .O(gate200inter9));
  nand2 gate1103(.a(s_79), .b(gate200inter3), .O(gate200inter10));
  nor2  gate1104(.a(gate200inter10), .b(gate200inter9), .O(gate200inter11));
  nor2  gate1105(.a(gate200inter11), .b(gate200inter6), .O(gate200inter12));
  nand2 gate1106(.a(gate200inter12), .b(gate200inter1), .O(G663));
nand2 gate201( .a(G602), .b(G607), .O(G666) );
nand2 gate202( .a(G612), .b(G617), .O(G669) );

  xor2  gate953(.a(G612), .b(G602), .O(gate203inter0));
  nand2 gate954(.a(gate203inter0), .b(s_58), .O(gate203inter1));
  and2  gate955(.a(G612), .b(G602), .O(gate203inter2));
  inv1  gate956(.a(s_58), .O(gate203inter3));
  inv1  gate957(.a(s_59), .O(gate203inter4));
  nand2 gate958(.a(gate203inter4), .b(gate203inter3), .O(gate203inter5));
  nor2  gate959(.a(gate203inter5), .b(gate203inter2), .O(gate203inter6));
  inv1  gate960(.a(G602), .O(gate203inter7));
  inv1  gate961(.a(G612), .O(gate203inter8));
  nand2 gate962(.a(gate203inter8), .b(gate203inter7), .O(gate203inter9));
  nand2 gate963(.a(s_59), .b(gate203inter3), .O(gate203inter10));
  nor2  gate964(.a(gate203inter10), .b(gate203inter9), .O(gate203inter11));
  nor2  gate965(.a(gate203inter11), .b(gate203inter6), .O(gate203inter12));
  nand2 gate966(.a(gate203inter12), .b(gate203inter1), .O(G672));
nand2 gate204( .a(G607), .b(G617), .O(G675) );
nand2 gate205( .a(G622), .b(G627), .O(G678) );

  xor2  gate1331(.a(G637), .b(G632), .O(gate206inter0));
  nand2 gate1332(.a(gate206inter0), .b(s_112), .O(gate206inter1));
  and2  gate1333(.a(G637), .b(G632), .O(gate206inter2));
  inv1  gate1334(.a(s_112), .O(gate206inter3));
  inv1  gate1335(.a(s_113), .O(gate206inter4));
  nand2 gate1336(.a(gate206inter4), .b(gate206inter3), .O(gate206inter5));
  nor2  gate1337(.a(gate206inter5), .b(gate206inter2), .O(gate206inter6));
  inv1  gate1338(.a(G632), .O(gate206inter7));
  inv1  gate1339(.a(G637), .O(gate206inter8));
  nand2 gate1340(.a(gate206inter8), .b(gate206inter7), .O(gate206inter9));
  nand2 gate1341(.a(s_113), .b(gate206inter3), .O(gate206inter10));
  nor2  gate1342(.a(gate206inter10), .b(gate206inter9), .O(gate206inter11));
  nor2  gate1343(.a(gate206inter11), .b(gate206inter6), .O(gate206inter12));
  nand2 gate1344(.a(gate206inter12), .b(gate206inter1), .O(G681));
nand2 gate207( .a(G622), .b(G632), .O(G684) );
nand2 gate208( .a(G627), .b(G637), .O(G687) );
nand2 gate209( .a(G602), .b(G666), .O(G690) );
nand2 gate210( .a(G607), .b(G666), .O(G691) );
nand2 gate211( .a(G612), .b(G669), .O(G692) );
nand2 gate212( .a(G617), .b(G669), .O(G693) );
nand2 gate213( .a(G602), .b(G672), .O(G694) );
nand2 gate214( .a(G612), .b(G672), .O(G695) );

  xor2  gate869(.a(G675), .b(G607), .O(gate215inter0));
  nand2 gate870(.a(gate215inter0), .b(s_46), .O(gate215inter1));
  and2  gate871(.a(G675), .b(G607), .O(gate215inter2));
  inv1  gate872(.a(s_46), .O(gate215inter3));
  inv1  gate873(.a(s_47), .O(gate215inter4));
  nand2 gate874(.a(gate215inter4), .b(gate215inter3), .O(gate215inter5));
  nor2  gate875(.a(gate215inter5), .b(gate215inter2), .O(gate215inter6));
  inv1  gate876(.a(G607), .O(gate215inter7));
  inv1  gate877(.a(G675), .O(gate215inter8));
  nand2 gate878(.a(gate215inter8), .b(gate215inter7), .O(gate215inter9));
  nand2 gate879(.a(s_47), .b(gate215inter3), .O(gate215inter10));
  nor2  gate880(.a(gate215inter10), .b(gate215inter9), .O(gate215inter11));
  nor2  gate881(.a(gate215inter11), .b(gate215inter6), .O(gate215inter12));
  nand2 gate882(.a(gate215inter12), .b(gate215inter1), .O(G696));
nand2 gate216( .a(G617), .b(G675), .O(G697) );
nand2 gate217( .a(G622), .b(G678), .O(G698) );
nand2 gate218( .a(G627), .b(G678), .O(G699) );

  xor2  gate1373(.a(G681), .b(G632), .O(gate219inter0));
  nand2 gate1374(.a(gate219inter0), .b(s_118), .O(gate219inter1));
  and2  gate1375(.a(G681), .b(G632), .O(gate219inter2));
  inv1  gate1376(.a(s_118), .O(gate219inter3));
  inv1  gate1377(.a(s_119), .O(gate219inter4));
  nand2 gate1378(.a(gate219inter4), .b(gate219inter3), .O(gate219inter5));
  nor2  gate1379(.a(gate219inter5), .b(gate219inter2), .O(gate219inter6));
  inv1  gate1380(.a(G632), .O(gate219inter7));
  inv1  gate1381(.a(G681), .O(gate219inter8));
  nand2 gate1382(.a(gate219inter8), .b(gate219inter7), .O(gate219inter9));
  nand2 gate1383(.a(s_119), .b(gate219inter3), .O(gate219inter10));
  nor2  gate1384(.a(gate219inter10), .b(gate219inter9), .O(gate219inter11));
  nor2  gate1385(.a(gate219inter11), .b(gate219inter6), .O(gate219inter12));
  nand2 gate1386(.a(gate219inter12), .b(gate219inter1), .O(G700));
nand2 gate220( .a(G637), .b(G681), .O(G701) );
nand2 gate221( .a(G622), .b(G684), .O(G702) );
nand2 gate222( .a(G632), .b(G684), .O(G703) );

  xor2  gate1807(.a(G687), .b(G627), .O(gate223inter0));
  nand2 gate1808(.a(gate223inter0), .b(s_180), .O(gate223inter1));
  and2  gate1809(.a(G687), .b(G627), .O(gate223inter2));
  inv1  gate1810(.a(s_180), .O(gate223inter3));
  inv1  gate1811(.a(s_181), .O(gate223inter4));
  nand2 gate1812(.a(gate223inter4), .b(gate223inter3), .O(gate223inter5));
  nor2  gate1813(.a(gate223inter5), .b(gate223inter2), .O(gate223inter6));
  inv1  gate1814(.a(G627), .O(gate223inter7));
  inv1  gate1815(.a(G687), .O(gate223inter8));
  nand2 gate1816(.a(gate223inter8), .b(gate223inter7), .O(gate223inter9));
  nand2 gate1817(.a(s_181), .b(gate223inter3), .O(gate223inter10));
  nor2  gate1818(.a(gate223inter10), .b(gate223inter9), .O(gate223inter11));
  nor2  gate1819(.a(gate223inter11), .b(gate223inter6), .O(gate223inter12));
  nand2 gate1820(.a(gate223inter12), .b(gate223inter1), .O(G704));
nand2 gate224( .a(G637), .b(G687), .O(G705) );
nand2 gate225( .a(G690), .b(G691), .O(G706) );
nand2 gate226( .a(G692), .b(G693), .O(G709) );
nand2 gate227( .a(G694), .b(G695), .O(G712) );

  xor2  gate603(.a(G697), .b(G696), .O(gate228inter0));
  nand2 gate604(.a(gate228inter0), .b(s_8), .O(gate228inter1));
  and2  gate605(.a(G697), .b(G696), .O(gate228inter2));
  inv1  gate606(.a(s_8), .O(gate228inter3));
  inv1  gate607(.a(s_9), .O(gate228inter4));
  nand2 gate608(.a(gate228inter4), .b(gate228inter3), .O(gate228inter5));
  nor2  gate609(.a(gate228inter5), .b(gate228inter2), .O(gate228inter6));
  inv1  gate610(.a(G696), .O(gate228inter7));
  inv1  gate611(.a(G697), .O(gate228inter8));
  nand2 gate612(.a(gate228inter8), .b(gate228inter7), .O(gate228inter9));
  nand2 gate613(.a(s_9), .b(gate228inter3), .O(gate228inter10));
  nor2  gate614(.a(gate228inter10), .b(gate228inter9), .O(gate228inter11));
  nor2  gate615(.a(gate228inter11), .b(gate228inter6), .O(gate228inter12));
  nand2 gate616(.a(gate228inter12), .b(gate228inter1), .O(G715));

  xor2  gate2143(.a(G699), .b(G698), .O(gate229inter0));
  nand2 gate2144(.a(gate229inter0), .b(s_228), .O(gate229inter1));
  and2  gate2145(.a(G699), .b(G698), .O(gate229inter2));
  inv1  gate2146(.a(s_228), .O(gate229inter3));
  inv1  gate2147(.a(s_229), .O(gate229inter4));
  nand2 gate2148(.a(gate229inter4), .b(gate229inter3), .O(gate229inter5));
  nor2  gate2149(.a(gate229inter5), .b(gate229inter2), .O(gate229inter6));
  inv1  gate2150(.a(G698), .O(gate229inter7));
  inv1  gate2151(.a(G699), .O(gate229inter8));
  nand2 gate2152(.a(gate229inter8), .b(gate229inter7), .O(gate229inter9));
  nand2 gate2153(.a(s_229), .b(gate229inter3), .O(gate229inter10));
  nor2  gate2154(.a(gate229inter10), .b(gate229inter9), .O(gate229inter11));
  nor2  gate2155(.a(gate229inter11), .b(gate229inter6), .O(gate229inter12));
  nand2 gate2156(.a(gate229inter12), .b(gate229inter1), .O(G718));

  xor2  gate2325(.a(G701), .b(G700), .O(gate230inter0));
  nand2 gate2326(.a(gate230inter0), .b(s_254), .O(gate230inter1));
  and2  gate2327(.a(G701), .b(G700), .O(gate230inter2));
  inv1  gate2328(.a(s_254), .O(gate230inter3));
  inv1  gate2329(.a(s_255), .O(gate230inter4));
  nand2 gate2330(.a(gate230inter4), .b(gate230inter3), .O(gate230inter5));
  nor2  gate2331(.a(gate230inter5), .b(gate230inter2), .O(gate230inter6));
  inv1  gate2332(.a(G700), .O(gate230inter7));
  inv1  gate2333(.a(G701), .O(gate230inter8));
  nand2 gate2334(.a(gate230inter8), .b(gate230inter7), .O(gate230inter9));
  nand2 gate2335(.a(s_255), .b(gate230inter3), .O(gate230inter10));
  nor2  gate2336(.a(gate230inter10), .b(gate230inter9), .O(gate230inter11));
  nor2  gate2337(.a(gate230inter11), .b(gate230inter6), .O(gate230inter12));
  nand2 gate2338(.a(gate230inter12), .b(gate230inter1), .O(G721));
nand2 gate231( .a(G702), .b(G703), .O(G724) );
nand2 gate232( .a(G704), .b(G705), .O(G727) );

  xor2  gate1485(.a(G718), .b(G242), .O(gate233inter0));
  nand2 gate1486(.a(gate233inter0), .b(s_134), .O(gate233inter1));
  and2  gate1487(.a(G718), .b(G242), .O(gate233inter2));
  inv1  gate1488(.a(s_134), .O(gate233inter3));
  inv1  gate1489(.a(s_135), .O(gate233inter4));
  nand2 gate1490(.a(gate233inter4), .b(gate233inter3), .O(gate233inter5));
  nor2  gate1491(.a(gate233inter5), .b(gate233inter2), .O(gate233inter6));
  inv1  gate1492(.a(G242), .O(gate233inter7));
  inv1  gate1493(.a(G718), .O(gate233inter8));
  nand2 gate1494(.a(gate233inter8), .b(gate233inter7), .O(gate233inter9));
  nand2 gate1495(.a(s_135), .b(gate233inter3), .O(gate233inter10));
  nor2  gate1496(.a(gate233inter10), .b(gate233inter9), .O(gate233inter11));
  nor2  gate1497(.a(gate233inter11), .b(gate233inter6), .O(gate233inter12));
  nand2 gate1498(.a(gate233inter12), .b(gate233inter1), .O(G730));

  xor2  gate1779(.a(G721), .b(G245), .O(gate234inter0));
  nand2 gate1780(.a(gate234inter0), .b(s_176), .O(gate234inter1));
  and2  gate1781(.a(G721), .b(G245), .O(gate234inter2));
  inv1  gate1782(.a(s_176), .O(gate234inter3));
  inv1  gate1783(.a(s_177), .O(gate234inter4));
  nand2 gate1784(.a(gate234inter4), .b(gate234inter3), .O(gate234inter5));
  nor2  gate1785(.a(gate234inter5), .b(gate234inter2), .O(gate234inter6));
  inv1  gate1786(.a(G245), .O(gate234inter7));
  inv1  gate1787(.a(G721), .O(gate234inter8));
  nand2 gate1788(.a(gate234inter8), .b(gate234inter7), .O(gate234inter9));
  nand2 gate1789(.a(s_177), .b(gate234inter3), .O(gate234inter10));
  nor2  gate1790(.a(gate234inter10), .b(gate234inter9), .O(gate234inter11));
  nor2  gate1791(.a(gate234inter11), .b(gate234inter6), .O(gate234inter12));
  nand2 gate1792(.a(gate234inter12), .b(gate234inter1), .O(G733));
nand2 gate235( .a(G248), .b(G724), .O(G736) );
nand2 gate236( .a(G251), .b(G727), .O(G739) );

  xor2  gate1023(.a(G706), .b(G254), .O(gate237inter0));
  nand2 gate1024(.a(gate237inter0), .b(s_68), .O(gate237inter1));
  and2  gate1025(.a(G706), .b(G254), .O(gate237inter2));
  inv1  gate1026(.a(s_68), .O(gate237inter3));
  inv1  gate1027(.a(s_69), .O(gate237inter4));
  nand2 gate1028(.a(gate237inter4), .b(gate237inter3), .O(gate237inter5));
  nor2  gate1029(.a(gate237inter5), .b(gate237inter2), .O(gate237inter6));
  inv1  gate1030(.a(G254), .O(gate237inter7));
  inv1  gate1031(.a(G706), .O(gate237inter8));
  nand2 gate1032(.a(gate237inter8), .b(gate237inter7), .O(gate237inter9));
  nand2 gate1033(.a(s_69), .b(gate237inter3), .O(gate237inter10));
  nor2  gate1034(.a(gate237inter10), .b(gate237inter9), .O(gate237inter11));
  nor2  gate1035(.a(gate237inter11), .b(gate237inter6), .O(gate237inter12));
  nand2 gate1036(.a(gate237inter12), .b(gate237inter1), .O(G742));
nand2 gate238( .a(G257), .b(G709), .O(G745) );

  xor2  gate1471(.a(G712), .b(G260), .O(gate239inter0));
  nand2 gate1472(.a(gate239inter0), .b(s_132), .O(gate239inter1));
  and2  gate1473(.a(G712), .b(G260), .O(gate239inter2));
  inv1  gate1474(.a(s_132), .O(gate239inter3));
  inv1  gate1475(.a(s_133), .O(gate239inter4));
  nand2 gate1476(.a(gate239inter4), .b(gate239inter3), .O(gate239inter5));
  nor2  gate1477(.a(gate239inter5), .b(gate239inter2), .O(gate239inter6));
  inv1  gate1478(.a(G260), .O(gate239inter7));
  inv1  gate1479(.a(G712), .O(gate239inter8));
  nand2 gate1480(.a(gate239inter8), .b(gate239inter7), .O(gate239inter9));
  nand2 gate1481(.a(s_133), .b(gate239inter3), .O(gate239inter10));
  nor2  gate1482(.a(gate239inter10), .b(gate239inter9), .O(gate239inter11));
  nor2  gate1483(.a(gate239inter11), .b(gate239inter6), .O(gate239inter12));
  nand2 gate1484(.a(gate239inter12), .b(gate239inter1), .O(G748));
nand2 gate240( .a(G263), .b(G715), .O(G751) );
nand2 gate241( .a(G242), .b(G730), .O(G754) );
nand2 gate242( .a(G718), .b(G730), .O(G755) );
nand2 gate243( .a(G245), .b(G733), .O(G756) );

  xor2  gate1555(.a(G733), .b(G721), .O(gate244inter0));
  nand2 gate1556(.a(gate244inter0), .b(s_144), .O(gate244inter1));
  and2  gate1557(.a(G733), .b(G721), .O(gate244inter2));
  inv1  gate1558(.a(s_144), .O(gate244inter3));
  inv1  gate1559(.a(s_145), .O(gate244inter4));
  nand2 gate1560(.a(gate244inter4), .b(gate244inter3), .O(gate244inter5));
  nor2  gate1561(.a(gate244inter5), .b(gate244inter2), .O(gate244inter6));
  inv1  gate1562(.a(G721), .O(gate244inter7));
  inv1  gate1563(.a(G733), .O(gate244inter8));
  nand2 gate1564(.a(gate244inter8), .b(gate244inter7), .O(gate244inter9));
  nand2 gate1565(.a(s_145), .b(gate244inter3), .O(gate244inter10));
  nor2  gate1566(.a(gate244inter10), .b(gate244inter9), .O(gate244inter11));
  nor2  gate1567(.a(gate244inter11), .b(gate244inter6), .O(gate244inter12));
  nand2 gate1568(.a(gate244inter12), .b(gate244inter1), .O(G757));
nand2 gate245( .a(G248), .b(G736), .O(G758) );
nand2 gate246( .a(G724), .b(G736), .O(G759) );
nand2 gate247( .a(G251), .b(G739), .O(G760) );
nand2 gate248( .a(G727), .b(G739), .O(G761) );

  xor2  gate2395(.a(G742), .b(G254), .O(gate249inter0));
  nand2 gate2396(.a(gate249inter0), .b(s_264), .O(gate249inter1));
  and2  gate2397(.a(G742), .b(G254), .O(gate249inter2));
  inv1  gate2398(.a(s_264), .O(gate249inter3));
  inv1  gate2399(.a(s_265), .O(gate249inter4));
  nand2 gate2400(.a(gate249inter4), .b(gate249inter3), .O(gate249inter5));
  nor2  gate2401(.a(gate249inter5), .b(gate249inter2), .O(gate249inter6));
  inv1  gate2402(.a(G254), .O(gate249inter7));
  inv1  gate2403(.a(G742), .O(gate249inter8));
  nand2 gate2404(.a(gate249inter8), .b(gate249inter7), .O(gate249inter9));
  nand2 gate2405(.a(s_265), .b(gate249inter3), .O(gate249inter10));
  nor2  gate2406(.a(gate249inter10), .b(gate249inter9), .O(gate249inter11));
  nor2  gate2407(.a(gate249inter11), .b(gate249inter6), .O(gate249inter12));
  nand2 gate2408(.a(gate249inter12), .b(gate249inter1), .O(G762));
nand2 gate250( .a(G706), .b(G742), .O(G763) );

  xor2  gate2003(.a(G745), .b(G257), .O(gate251inter0));
  nand2 gate2004(.a(gate251inter0), .b(s_208), .O(gate251inter1));
  and2  gate2005(.a(G745), .b(G257), .O(gate251inter2));
  inv1  gate2006(.a(s_208), .O(gate251inter3));
  inv1  gate2007(.a(s_209), .O(gate251inter4));
  nand2 gate2008(.a(gate251inter4), .b(gate251inter3), .O(gate251inter5));
  nor2  gate2009(.a(gate251inter5), .b(gate251inter2), .O(gate251inter6));
  inv1  gate2010(.a(G257), .O(gate251inter7));
  inv1  gate2011(.a(G745), .O(gate251inter8));
  nand2 gate2012(.a(gate251inter8), .b(gate251inter7), .O(gate251inter9));
  nand2 gate2013(.a(s_209), .b(gate251inter3), .O(gate251inter10));
  nor2  gate2014(.a(gate251inter10), .b(gate251inter9), .O(gate251inter11));
  nor2  gate2015(.a(gate251inter11), .b(gate251inter6), .O(gate251inter12));
  nand2 gate2016(.a(gate251inter12), .b(gate251inter1), .O(G764));

  xor2  gate1905(.a(G745), .b(G709), .O(gate252inter0));
  nand2 gate1906(.a(gate252inter0), .b(s_194), .O(gate252inter1));
  and2  gate1907(.a(G745), .b(G709), .O(gate252inter2));
  inv1  gate1908(.a(s_194), .O(gate252inter3));
  inv1  gate1909(.a(s_195), .O(gate252inter4));
  nand2 gate1910(.a(gate252inter4), .b(gate252inter3), .O(gate252inter5));
  nor2  gate1911(.a(gate252inter5), .b(gate252inter2), .O(gate252inter6));
  inv1  gate1912(.a(G709), .O(gate252inter7));
  inv1  gate1913(.a(G745), .O(gate252inter8));
  nand2 gate1914(.a(gate252inter8), .b(gate252inter7), .O(gate252inter9));
  nand2 gate1915(.a(s_195), .b(gate252inter3), .O(gate252inter10));
  nor2  gate1916(.a(gate252inter10), .b(gate252inter9), .O(gate252inter11));
  nor2  gate1917(.a(gate252inter11), .b(gate252inter6), .O(gate252inter12));
  nand2 gate1918(.a(gate252inter12), .b(gate252inter1), .O(G765));
nand2 gate253( .a(G260), .b(G748), .O(G766) );
nand2 gate254( .a(G712), .b(G748), .O(G767) );
nand2 gate255( .a(G263), .b(G751), .O(G768) );
nand2 gate256( .a(G715), .b(G751), .O(G769) );

  xor2  gate645(.a(G755), .b(G754), .O(gate257inter0));
  nand2 gate646(.a(gate257inter0), .b(s_14), .O(gate257inter1));
  and2  gate647(.a(G755), .b(G754), .O(gate257inter2));
  inv1  gate648(.a(s_14), .O(gate257inter3));
  inv1  gate649(.a(s_15), .O(gate257inter4));
  nand2 gate650(.a(gate257inter4), .b(gate257inter3), .O(gate257inter5));
  nor2  gate651(.a(gate257inter5), .b(gate257inter2), .O(gate257inter6));
  inv1  gate652(.a(G754), .O(gate257inter7));
  inv1  gate653(.a(G755), .O(gate257inter8));
  nand2 gate654(.a(gate257inter8), .b(gate257inter7), .O(gate257inter9));
  nand2 gate655(.a(s_15), .b(gate257inter3), .O(gate257inter10));
  nor2  gate656(.a(gate257inter10), .b(gate257inter9), .O(gate257inter11));
  nor2  gate657(.a(gate257inter11), .b(gate257inter6), .O(gate257inter12));
  nand2 gate658(.a(gate257inter12), .b(gate257inter1), .O(G770));

  xor2  gate967(.a(G757), .b(G756), .O(gate258inter0));
  nand2 gate968(.a(gate258inter0), .b(s_60), .O(gate258inter1));
  and2  gate969(.a(G757), .b(G756), .O(gate258inter2));
  inv1  gate970(.a(s_60), .O(gate258inter3));
  inv1  gate971(.a(s_61), .O(gate258inter4));
  nand2 gate972(.a(gate258inter4), .b(gate258inter3), .O(gate258inter5));
  nor2  gate973(.a(gate258inter5), .b(gate258inter2), .O(gate258inter6));
  inv1  gate974(.a(G756), .O(gate258inter7));
  inv1  gate975(.a(G757), .O(gate258inter8));
  nand2 gate976(.a(gate258inter8), .b(gate258inter7), .O(gate258inter9));
  nand2 gate977(.a(s_61), .b(gate258inter3), .O(gate258inter10));
  nor2  gate978(.a(gate258inter10), .b(gate258inter9), .O(gate258inter11));
  nor2  gate979(.a(gate258inter11), .b(gate258inter6), .O(gate258inter12));
  nand2 gate980(.a(gate258inter12), .b(gate258inter1), .O(G773));

  xor2  gate1233(.a(G759), .b(G758), .O(gate259inter0));
  nand2 gate1234(.a(gate259inter0), .b(s_98), .O(gate259inter1));
  and2  gate1235(.a(G759), .b(G758), .O(gate259inter2));
  inv1  gate1236(.a(s_98), .O(gate259inter3));
  inv1  gate1237(.a(s_99), .O(gate259inter4));
  nand2 gate1238(.a(gate259inter4), .b(gate259inter3), .O(gate259inter5));
  nor2  gate1239(.a(gate259inter5), .b(gate259inter2), .O(gate259inter6));
  inv1  gate1240(.a(G758), .O(gate259inter7));
  inv1  gate1241(.a(G759), .O(gate259inter8));
  nand2 gate1242(.a(gate259inter8), .b(gate259inter7), .O(gate259inter9));
  nand2 gate1243(.a(s_99), .b(gate259inter3), .O(gate259inter10));
  nor2  gate1244(.a(gate259inter10), .b(gate259inter9), .O(gate259inter11));
  nor2  gate1245(.a(gate259inter11), .b(gate259inter6), .O(gate259inter12));
  nand2 gate1246(.a(gate259inter12), .b(gate259inter1), .O(G776));
nand2 gate260( .a(G760), .b(G761), .O(G779) );
nand2 gate261( .a(G762), .b(G763), .O(G782) );
nand2 gate262( .a(G764), .b(G765), .O(G785) );
nand2 gate263( .a(G766), .b(G767), .O(G788) );

  xor2  gate617(.a(G769), .b(G768), .O(gate264inter0));
  nand2 gate618(.a(gate264inter0), .b(s_10), .O(gate264inter1));
  and2  gate619(.a(G769), .b(G768), .O(gate264inter2));
  inv1  gate620(.a(s_10), .O(gate264inter3));
  inv1  gate621(.a(s_11), .O(gate264inter4));
  nand2 gate622(.a(gate264inter4), .b(gate264inter3), .O(gate264inter5));
  nor2  gate623(.a(gate264inter5), .b(gate264inter2), .O(gate264inter6));
  inv1  gate624(.a(G768), .O(gate264inter7));
  inv1  gate625(.a(G769), .O(gate264inter8));
  nand2 gate626(.a(gate264inter8), .b(gate264inter7), .O(gate264inter9));
  nand2 gate627(.a(s_11), .b(gate264inter3), .O(gate264inter10));
  nor2  gate628(.a(gate264inter10), .b(gate264inter9), .O(gate264inter11));
  nor2  gate629(.a(gate264inter11), .b(gate264inter6), .O(gate264inter12));
  nand2 gate630(.a(gate264inter12), .b(gate264inter1), .O(G791));
nand2 gate265( .a(G642), .b(G770), .O(G794) );
nand2 gate266( .a(G645), .b(G773), .O(G797) );
nand2 gate267( .a(G648), .b(G776), .O(G800) );
nand2 gate268( .a(G651), .b(G779), .O(G803) );
nand2 gate269( .a(G654), .b(G782), .O(G806) );
nand2 gate270( .a(G657), .b(G785), .O(G809) );
nand2 gate271( .a(G660), .b(G788), .O(G812) );
nand2 gate272( .a(G663), .b(G791), .O(G815) );
nand2 gate273( .a(G642), .b(G794), .O(G818) );
nand2 gate274( .a(G770), .b(G794), .O(G819) );
nand2 gate275( .a(G645), .b(G797), .O(G820) );

  xor2  gate1079(.a(G797), .b(G773), .O(gate276inter0));
  nand2 gate1080(.a(gate276inter0), .b(s_76), .O(gate276inter1));
  and2  gate1081(.a(G797), .b(G773), .O(gate276inter2));
  inv1  gate1082(.a(s_76), .O(gate276inter3));
  inv1  gate1083(.a(s_77), .O(gate276inter4));
  nand2 gate1084(.a(gate276inter4), .b(gate276inter3), .O(gate276inter5));
  nor2  gate1085(.a(gate276inter5), .b(gate276inter2), .O(gate276inter6));
  inv1  gate1086(.a(G773), .O(gate276inter7));
  inv1  gate1087(.a(G797), .O(gate276inter8));
  nand2 gate1088(.a(gate276inter8), .b(gate276inter7), .O(gate276inter9));
  nand2 gate1089(.a(s_77), .b(gate276inter3), .O(gate276inter10));
  nor2  gate1090(.a(gate276inter10), .b(gate276inter9), .O(gate276inter11));
  nor2  gate1091(.a(gate276inter11), .b(gate276inter6), .O(gate276inter12));
  nand2 gate1092(.a(gate276inter12), .b(gate276inter1), .O(G821));

  xor2  gate1177(.a(G800), .b(G648), .O(gate277inter0));
  nand2 gate1178(.a(gate277inter0), .b(s_90), .O(gate277inter1));
  and2  gate1179(.a(G800), .b(G648), .O(gate277inter2));
  inv1  gate1180(.a(s_90), .O(gate277inter3));
  inv1  gate1181(.a(s_91), .O(gate277inter4));
  nand2 gate1182(.a(gate277inter4), .b(gate277inter3), .O(gate277inter5));
  nor2  gate1183(.a(gate277inter5), .b(gate277inter2), .O(gate277inter6));
  inv1  gate1184(.a(G648), .O(gate277inter7));
  inv1  gate1185(.a(G800), .O(gate277inter8));
  nand2 gate1186(.a(gate277inter8), .b(gate277inter7), .O(gate277inter9));
  nand2 gate1187(.a(s_91), .b(gate277inter3), .O(gate277inter10));
  nor2  gate1188(.a(gate277inter10), .b(gate277inter9), .O(gate277inter11));
  nor2  gate1189(.a(gate277inter11), .b(gate277inter6), .O(gate277inter12));
  nand2 gate1190(.a(gate277inter12), .b(gate277inter1), .O(G822));

  xor2  gate715(.a(G800), .b(G776), .O(gate278inter0));
  nand2 gate716(.a(gate278inter0), .b(s_24), .O(gate278inter1));
  and2  gate717(.a(G800), .b(G776), .O(gate278inter2));
  inv1  gate718(.a(s_24), .O(gate278inter3));
  inv1  gate719(.a(s_25), .O(gate278inter4));
  nand2 gate720(.a(gate278inter4), .b(gate278inter3), .O(gate278inter5));
  nor2  gate721(.a(gate278inter5), .b(gate278inter2), .O(gate278inter6));
  inv1  gate722(.a(G776), .O(gate278inter7));
  inv1  gate723(.a(G800), .O(gate278inter8));
  nand2 gate724(.a(gate278inter8), .b(gate278inter7), .O(gate278inter9));
  nand2 gate725(.a(s_25), .b(gate278inter3), .O(gate278inter10));
  nor2  gate726(.a(gate278inter10), .b(gate278inter9), .O(gate278inter11));
  nor2  gate727(.a(gate278inter11), .b(gate278inter6), .O(gate278inter12));
  nand2 gate728(.a(gate278inter12), .b(gate278inter1), .O(G823));
nand2 gate279( .a(G651), .b(G803), .O(G824) );
nand2 gate280( .a(G779), .b(G803), .O(G825) );
nand2 gate281( .a(G654), .b(G806), .O(G826) );
nand2 gate282( .a(G782), .b(G806), .O(G827) );
nand2 gate283( .a(G657), .b(G809), .O(G828) );
nand2 gate284( .a(G785), .b(G809), .O(G829) );
nand2 gate285( .a(G660), .b(G812), .O(G830) );

  xor2  gate701(.a(G812), .b(G788), .O(gate286inter0));
  nand2 gate702(.a(gate286inter0), .b(s_22), .O(gate286inter1));
  and2  gate703(.a(G812), .b(G788), .O(gate286inter2));
  inv1  gate704(.a(s_22), .O(gate286inter3));
  inv1  gate705(.a(s_23), .O(gate286inter4));
  nand2 gate706(.a(gate286inter4), .b(gate286inter3), .O(gate286inter5));
  nor2  gate707(.a(gate286inter5), .b(gate286inter2), .O(gate286inter6));
  inv1  gate708(.a(G788), .O(gate286inter7));
  inv1  gate709(.a(G812), .O(gate286inter8));
  nand2 gate710(.a(gate286inter8), .b(gate286inter7), .O(gate286inter9));
  nand2 gate711(.a(s_23), .b(gate286inter3), .O(gate286inter10));
  nor2  gate712(.a(gate286inter10), .b(gate286inter9), .O(gate286inter11));
  nor2  gate713(.a(gate286inter11), .b(gate286inter6), .O(gate286inter12));
  nand2 gate714(.a(gate286inter12), .b(gate286inter1), .O(G831));
nand2 gate287( .a(G663), .b(G815), .O(G832) );

  xor2  gate1009(.a(G815), .b(G791), .O(gate288inter0));
  nand2 gate1010(.a(gate288inter0), .b(s_66), .O(gate288inter1));
  and2  gate1011(.a(G815), .b(G791), .O(gate288inter2));
  inv1  gate1012(.a(s_66), .O(gate288inter3));
  inv1  gate1013(.a(s_67), .O(gate288inter4));
  nand2 gate1014(.a(gate288inter4), .b(gate288inter3), .O(gate288inter5));
  nor2  gate1015(.a(gate288inter5), .b(gate288inter2), .O(gate288inter6));
  inv1  gate1016(.a(G791), .O(gate288inter7));
  inv1  gate1017(.a(G815), .O(gate288inter8));
  nand2 gate1018(.a(gate288inter8), .b(gate288inter7), .O(gate288inter9));
  nand2 gate1019(.a(s_67), .b(gate288inter3), .O(gate288inter10));
  nor2  gate1020(.a(gate288inter10), .b(gate288inter9), .O(gate288inter11));
  nor2  gate1021(.a(gate288inter11), .b(gate288inter6), .O(gate288inter12));
  nand2 gate1022(.a(gate288inter12), .b(gate288inter1), .O(G833));
nand2 gate289( .a(G818), .b(G819), .O(G834) );

  xor2  gate2367(.a(G821), .b(G820), .O(gate290inter0));
  nand2 gate2368(.a(gate290inter0), .b(s_260), .O(gate290inter1));
  and2  gate2369(.a(G821), .b(G820), .O(gate290inter2));
  inv1  gate2370(.a(s_260), .O(gate290inter3));
  inv1  gate2371(.a(s_261), .O(gate290inter4));
  nand2 gate2372(.a(gate290inter4), .b(gate290inter3), .O(gate290inter5));
  nor2  gate2373(.a(gate290inter5), .b(gate290inter2), .O(gate290inter6));
  inv1  gate2374(.a(G820), .O(gate290inter7));
  inv1  gate2375(.a(G821), .O(gate290inter8));
  nand2 gate2376(.a(gate290inter8), .b(gate290inter7), .O(gate290inter9));
  nand2 gate2377(.a(s_261), .b(gate290inter3), .O(gate290inter10));
  nor2  gate2378(.a(gate290inter10), .b(gate290inter9), .O(gate290inter11));
  nor2  gate2379(.a(gate290inter11), .b(gate290inter6), .O(gate290inter12));
  nand2 gate2380(.a(gate290inter12), .b(gate290inter1), .O(G847));
nand2 gate291( .a(G822), .b(G823), .O(G860) );
nand2 gate292( .a(G824), .b(G825), .O(G873) );
nand2 gate293( .a(G828), .b(G829), .O(G886) );

  xor2  gate995(.a(G833), .b(G832), .O(gate294inter0));
  nand2 gate996(.a(gate294inter0), .b(s_64), .O(gate294inter1));
  and2  gate997(.a(G833), .b(G832), .O(gate294inter2));
  inv1  gate998(.a(s_64), .O(gate294inter3));
  inv1  gate999(.a(s_65), .O(gate294inter4));
  nand2 gate1000(.a(gate294inter4), .b(gate294inter3), .O(gate294inter5));
  nor2  gate1001(.a(gate294inter5), .b(gate294inter2), .O(gate294inter6));
  inv1  gate1002(.a(G832), .O(gate294inter7));
  inv1  gate1003(.a(G833), .O(gate294inter8));
  nand2 gate1004(.a(gate294inter8), .b(gate294inter7), .O(gate294inter9));
  nand2 gate1005(.a(s_65), .b(gate294inter3), .O(gate294inter10));
  nor2  gate1006(.a(gate294inter10), .b(gate294inter9), .O(gate294inter11));
  nor2  gate1007(.a(gate294inter11), .b(gate294inter6), .O(gate294inter12));
  nand2 gate1008(.a(gate294inter12), .b(gate294inter1), .O(G899));
nand2 gate295( .a(G830), .b(G831), .O(G912) );
nand2 gate296( .a(G826), .b(G827), .O(G925) );
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );

  xor2  gate2269(.a(G1036), .b(G1), .O(gate387inter0));
  nand2 gate2270(.a(gate387inter0), .b(s_246), .O(gate387inter1));
  and2  gate2271(.a(G1036), .b(G1), .O(gate387inter2));
  inv1  gate2272(.a(s_246), .O(gate387inter3));
  inv1  gate2273(.a(s_247), .O(gate387inter4));
  nand2 gate2274(.a(gate387inter4), .b(gate387inter3), .O(gate387inter5));
  nor2  gate2275(.a(gate387inter5), .b(gate387inter2), .O(gate387inter6));
  inv1  gate2276(.a(G1), .O(gate387inter7));
  inv1  gate2277(.a(G1036), .O(gate387inter8));
  nand2 gate2278(.a(gate387inter8), .b(gate387inter7), .O(gate387inter9));
  nand2 gate2279(.a(s_247), .b(gate387inter3), .O(gate387inter10));
  nor2  gate2280(.a(gate387inter10), .b(gate387inter9), .O(gate387inter11));
  nor2  gate2281(.a(gate387inter11), .b(gate387inter6), .O(gate387inter12));
  nand2 gate2282(.a(gate387inter12), .b(gate387inter1), .O(G1132));

  xor2  gate1541(.a(G1039), .b(G2), .O(gate388inter0));
  nand2 gate1542(.a(gate388inter0), .b(s_142), .O(gate388inter1));
  and2  gate1543(.a(G1039), .b(G2), .O(gate388inter2));
  inv1  gate1544(.a(s_142), .O(gate388inter3));
  inv1  gate1545(.a(s_143), .O(gate388inter4));
  nand2 gate1546(.a(gate388inter4), .b(gate388inter3), .O(gate388inter5));
  nor2  gate1547(.a(gate388inter5), .b(gate388inter2), .O(gate388inter6));
  inv1  gate1548(.a(G2), .O(gate388inter7));
  inv1  gate1549(.a(G1039), .O(gate388inter8));
  nand2 gate1550(.a(gate388inter8), .b(gate388inter7), .O(gate388inter9));
  nand2 gate1551(.a(s_143), .b(gate388inter3), .O(gate388inter10));
  nor2  gate1552(.a(gate388inter10), .b(gate388inter9), .O(gate388inter11));
  nor2  gate1553(.a(gate388inter11), .b(gate388inter6), .O(gate388inter12));
  nand2 gate1554(.a(gate388inter12), .b(gate388inter1), .O(G1135));

  xor2  gate729(.a(G1042), .b(G3), .O(gate389inter0));
  nand2 gate730(.a(gate389inter0), .b(s_26), .O(gate389inter1));
  and2  gate731(.a(G1042), .b(G3), .O(gate389inter2));
  inv1  gate732(.a(s_26), .O(gate389inter3));
  inv1  gate733(.a(s_27), .O(gate389inter4));
  nand2 gate734(.a(gate389inter4), .b(gate389inter3), .O(gate389inter5));
  nor2  gate735(.a(gate389inter5), .b(gate389inter2), .O(gate389inter6));
  inv1  gate736(.a(G3), .O(gate389inter7));
  inv1  gate737(.a(G1042), .O(gate389inter8));
  nand2 gate738(.a(gate389inter8), .b(gate389inter7), .O(gate389inter9));
  nand2 gate739(.a(s_27), .b(gate389inter3), .O(gate389inter10));
  nor2  gate740(.a(gate389inter10), .b(gate389inter9), .O(gate389inter11));
  nor2  gate741(.a(gate389inter11), .b(gate389inter6), .O(gate389inter12));
  nand2 gate742(.a(gate389inter12), .b(gate389inter1), .O(G1138));
nand2 gate390( .a(G4), .b(G1045), .O(G1141) );
nand2 gate391( .a(G5), .b(G1048), .O(G1144) );
nand2 gate392( .a(G6), .b(G1051), .O(G1147) );
nand2 gate393( .a(G7), .b(G1054), .O(G1150) );

  xor2  gate1849(.a(G1057), .b(G8), .O(gate394inter0));
  nand2 gate1850(.a(gate394inter0), .b(s_186), .O(gate394inter1));
  and2  gate1851(.a(G1057), .b(G8), .O(gate394inter2));
  inv1  gate1852(.a(s_186), .O(gate394inter3));
  inv1  gate1853(.a(s_187), .O(gate394inter4));
  nand2 gate1854(.a(gate394inter4), .b(gate394inter3), .O(gate394inter5));
  nor2  gate1855(.a(gate394inter5), .b(gate394inter2), .O(gate394inter6));
  inv1  gate1856(.a(G8), .O(gate394inter7));
  inv1  gate1857(.a(G1057), .O(gate394inter8));
  nand2 gate1858(.a(gate394inter8), .b(gate394inter7), .O(gate394inter9));
  nand2 gate1859(.a(s_187), .b(gate394inter3), .O(gate394inter10));
  nor2  gate1860(.a(gate394inter10), .b(gate394inter9), .O(gate394inter11));
  nor2  gate1861(.a(gate394inter11), .b(gate394inter6), .O(gate394inter12));
  nand2 gate1862(.a(gate394inter12), .b(gate394inter1), .O(G1153));
nand2 gate395( .a(G9), .b(G1060), .O(G1156) );
nand2 gate396( .a(G10), .b(G1063), .O(G1159) );

  xor2  gate855(.a(G1066), .b(G11), .O(gate397inter0));
  nand2 gate856(.a(gate397inter0), .b(s_44), .O(gate397inter1));
  and2  gate857(.a(G1066), .b(G11), .O(gate397inter2));
  inv1  gate858(.a(s_44), .O(gate397inter3));
  inv1  gate859(.a(s_45), .O(gate397inter4));
  nand2 gate860(.a(gate397inter4), .b(gate397inter3), .O(gate397inter5));
  nor2  gate861(.a(gate397inter5), .b(gate397inter2), .O(gate397inter6));
  inv1  gate862(.a(G11), .O(gate397inter7));
  inv1  gate863(.a(G1066), .O(gate397inter8));
  nand2 gate864(.a(gate397inter8), .b(gate397inter7), .O(gate397inter9));
  nand2 gate865(.a(s_45), .b(gate397inter3), .O(gate397inter10));
  nor2  gate866(.a(gate397inter10), .b(gate397inter9), .O(gate397inter11));
  nor2  gate867(.a(gate397inter11), .b(gate397inter6), .O(gate397inter12));
  nand2 gate868(.a(gate397inter12), .b(gate397inter1), .O(G1162));
nand2 gate398( .a(G12), .b(G1069), .O(G1165) );

  xor2  gate1121(.a(G1072), .b(G13), .O(gate399inter0));
  nand2 gate1122(.a(gate399inter0), .b(s_82), .O(gate399inter1));
  and2  gate1123(.a(G1072), .b(G13), .O(gate399inter2));
  inv1  gate1124(.a(s_82), .O(gate399inter3));
  inv1  gate1125(.a(s_83), .O(gate399inter4));
  nand2 gate1126(.a(gate399inter4), .b(gate399inter3), .O(gate399inter5));
  nor2  gate1127(.a(gate399inter5), .b(gate399inter2), .O(gate399inter6));
  inv1  gate1128(.a(G13), .O(gate399inter7));
  inv1  gate1129(.a(G1072), .O(gate399inter8));
  nand2 gate1130(.a(gate399inter8), .b(gate399inter7), .O(gate399inter9));
  nand2 gate1131(.a(s_83), .b(gate399inter3), .O(gate399inter10));
  nor2  gate1132(.a(gate399inter10), .b(gate399inter9), .O(gate399inter11));
  nor2  gate1133(.a(gate399inter11), .b(gate399inter6), .O(gate399inter12));
  nand2 gate1134(.a(gate399inter12), .b(gate399inter1), .O(G1168));
nand2 gate400( .a(G14), .b(G1075), .O(G1171) );
nand2 gate401( .a(G15), .b(G1078), .O(G1174) );
nand2 gate402( .a(G16), .b(G1081), .O(G1177) );
nand2 gate403( .a(G17), .b(G1084), .O(G1180) );

  xor2  gate1667(.a(G1087), .b(G18), .O(gate404inter0));
  nand2 gate1668(.a(gate404inter0), .b(s_160), .O(gate404inter1));
  and2  gate1669(.a(G1087), .b(G18), .O(gate404inter2));
  inv1  gate1670(.a(s_160), .O(gate404inter3));
  inv1  gate1671(.a(s_161), .O(gate404inter4));
  nand2 gate1672(.a(gate404inter4), .b(gate404inter3), .O(gate404inter5));
  nor2  gate1673(.a(gate404inter5), .b(gate404inter2), .O(gate404inter6));
  inv1  gate1674(.a(G18), .O(gate404inter7));
  inv1  gate1675(.a(G1087), .O(gate404inter8));
  nand2 gate1676(.a(gate404inter8), .b(gate404inter7), .O(gate404inter9));
  nand2 gate1677(.a(s_161), .b(gate404inter3), .O(gate404inter10));
  nor2  gate1678(.a(gate404inter10), .b(gate404inter9), .O(gate404inter11));
  nor2  gate1679(.a(gate404inter11), .b(gate404inter6), .O(gate404inter12));
  nand2 gate1680(.a(gate404inter12), .b(gate404inter1), .O(G1183));
nand2 gate405( .a(G19), .b(G1090), .O(G1186) );
nand2 gate406( .a(G20), .b(G1093), .O(G1189) );
nand2 gate407( .a(G21), .b(G1096), .O(G1192) );
nand2 gate408( .a(G22), .b(G1099), .O(G1195) );
nand2 gate409( .a(G23), .b(G1102), .O(G1198) );
nand2 gate410( .a(G24), .b(G1105), .O(G1201) );
nand2 gate411( .a(G25), .b(G1108), .O(G1204) );
nand2 gate412( .a(G26), .b(G1111), .O(G1207) );
nand2 gate413( .a(G27), .b(G1114), .O(G1210) );

  xor2  gate2423(.a(G1117), .b(G28), .O(gate414inter0));
  nand2 gate2424(.a(gate414inter0), .b(s_268), .O(gate414inter1));
  and2  gate2425(.a(G1117), .b(G28), .O(gate414inter2));
  inv1  gate2426(.a(s_268), .O(gate414inter3));
  inv1  gate2427(.a(s_269), .O(gate414inter4));
  nand2 gate2428(.a(gate414inter4), .b(gate414inter3), .O(gate414inter5));
  nor2  gate2429(.a(gate414inter5), .b(gate414inter2), .O(gate414inter6));
  inv1  gate2430(.a(G28), .O(gate414inter7));
  inv1  gate2431(.a(G1117), .O(gate414inter8));
  nand2 gate2432(.a(gate414inter8), .b(gate414inter7), .O(gate414inter9));
  nand2 gate2433(.a(s_269), .b(gate414inter3), .O(gate414inter10));
  nor2  gate2434(.a(gate414inter10), .b(gate414inter9), .O(gate414inter11));
  nor2  gate2435(.a(gate414inter11), .b(gate414inter6), .O(gate414inter12));
  nand2 gate2436(.a(gate414inter12), .b(gate414inter1), .O(G1213));
nand2 gate415( .a(G29), .b(G1120), .O(G1216) );

  xor2  gate827(.a(G1123), .b(G30), .O(gate416inter0));
  nand2 gate828(.a(gate416inter0), .b(s_40), .O(gate416inter1));
  and2  gate829(.a(G1123), .b(G30), .O(gate416inter2));
  inv1  gate830(.a(s_40), .O(gate416inter3));
  inv1  gate831(.a(s_41), .O(gate416inter4));
  nand2 gate832(.a(gate416inter4), .b(gate416inter3), .O(gate416inter5));
  nor2  gate833(.a(gate416inter5), .b(gate416inter2), .O(gate416inter6));
  inv1  gate834(.a(G30), .O(gate416inter7));
  inv1  gate835(.a(G1123), .O(gate416inter8));
  nand2 gate836(.a(gate416inter8), .b(gate416inter7), .O(gate416inter9));
  nand2 gate837(.a(s_41), .b(gate416inter3), .O(gate416inter10));
  nor2  gate838(.a(gate416inter10), .b(gate416inter9), .O(gate416inter11));
  nor2  gate839(.a(gate416inter11), .b(gate416inter6), .O(gate416inter12));
  nand2 gate840(.a(gate416inter12), .b(gate416inter1), .O(G1219));

  xor2  gate2129(.a(G1126), .b(G31), .O(gate417inter0));
  nand2 gate2130(.a(gate417inter0), .b(s_226), .O(gate417inter1));
  and2  gate2131(.a(G1126), .b(G31), .O(gate417inter2));
  inv1  gate2132(.a(s_226), .O(gate417inter3));
  inv1  gate2133(.a(s_227), .O(gate417inter4));
  nand2 gate2134(.a(gate417inter4), .b(gate417inter3), .O(gate417inter5));
  nor2  gate2135(.a(gate417inter5), .b(gate417inter2), .O(gate417inter6));
  inv1  gate2136(.a(G31), .O(gate417inter7));
  inv1  gate2137(.a(G1126), .O(gate417inter8));
  nand2 gate2138(.a(gate417inter8), .b(gate417inter7), .O(gate417inter9));
  nand2 gate2139(.a(s_227), .b(gate417inter3), .O(gate417inter10));
  nor2  gate2140(.a(gate417inter10), .b(gate417inter9), .O(gate417inter11));
  nor2  gate2141(.a(gate417inter11), .b(gate417inter6), .O(gate417inter12));
  nand2 gate2142(.a(gate417inter12), .b(gate417inter1), .O(G1222));

  xor2  gate2017(.a(G1129), .b(G32), .O(gate418inter0));
  nand2 gate2018(.a(gate418inter0), .b(s_210), .O(gate418inter1));
  and2  gate2019(.a(G1129), .b(G32), .O(gate418inter2));
  inv1  gate2020(.a(s_210), .O(gate418inter3));
  inv1  gate2021(.a(s_211), .O(gate418inter4));
  nand2 gate2022(.a(gate418inter4), .b(gate418inter3), .O(gate418inter5));
  nor2  gate2023(.a(gate418inter5), .b(gate418inter2), .O(gate418inter6));
  inv1  gate2024(.a(G32), .O(gate418inter7));
  inv1  gate2025(.a(G1129), .O(gate418inter8));
  nand2 gate2026(.a(gate418inter8), .b(gate418inter7), .O(gate418inter9));
  nand2 gate2027(.a(s_211), .b(gate418inter3), .O(gate418inter10));
  nor2  gate2028(.a(gate418inter10), .b(gate418inter9), .O(gate418inter11));
  nor2  gate2029(.a(gate418inter11), .b(gate418inter6), .O(gate418inter12));
  nand2 gate2030(.a(gate418inter12), .b(gate418inter1), .O(G1225));
nand2 gate419( .a(G1), .b(G1132), .O(G1228) );
nand2 gate420( .a(G1036), .b(G1132), .O(G1229) );
nand2 gate421( .a(G2), .b(G1135), .O(G1230) );

  xor2  gate1387(.a(G1135), .b(G1039), .O(gate422inter0));
  nand2 gate1388(.a(gate422inter0), .b(s_120), .O(gate422inter1));
  and2  gate1389(.a(G1135), .b(G1039), .O(gate422inter2));
  inv1  gate1390(.a(s_120), .O(gate422inter3));
  inv1  gate1391(.a(s_121), .O(gate422inter4));
  nand2 gate1392(.a(gate422inter4), .b(gate422inter3), .O(gate422inter5));
  nor2  gate1393(.a(gate422inter5), .b(gate422inter2), .O(gate422inter6));
  inv1  gate1394(.a(G1039), .O(gate422inter7));
  inv1  gate1395(.a(G1135), .O(gate422inter8));
  nand2 gate1396(.a(gate422inter8), .b(gate422inter7), .O(gate422inter9));
  nand2 gate1397(.a(s_121), .b(gate422inter3), .O(gate422inter10));
  nor2  gate1398(.a(gate422inter10), .b(gate422inter9), .O(gate422inter11));
  nor2  gate1399(.a(gate422inter11), .b(gate422inter6), .O(gate422inter12));
  nand2 gate1400(.a(gate422inter12), .b(gate422inter1), .O(G1231));
nand2 gate423( .a(G3), .b(G1138), .O(G1232) );
nand2 gate424( .a(G1042), .b(G1138), .O(G1233) );

  xor2  gate1933(.a(G1141), .b(G4), .O(gate425inter0));
  nand2 gate1934(.a(gate425inter0), .b(s_198), .O(gate425inter1));
  and2  gate1935(.a(G1141), .b(G4), .O(gate425inter2));
  inv1  gate1936(.a(s_198), .O(gate425inter3));
  inv1  gate1937(.a(s_199), .O(gate425inter4));
  nand2 gate1938(.a(gate425inter4), .b(gate425inter3), .O(gate425inter5));
  nor2  gate1939(.a(gate425inter5), .b(gate425inter2), .O(gate425inter6));
  inv1  gate1940(.a(G4), .O(gate425inter7));
  inv1  gate1941(.a(G1141), .O(gate425inter8));
  nand2 gate1942(.a(gate425inter8), .b(gate425inter7), .O(gate425inter9));
  nand2 gate1943(.a(s_199), .b(gate425inter3), .O(gate425inter10));
  nor2  gate1944(.a(gate425inter10), .b(gate425inter9), .O(gate425inter11));
  nor2  gate1945(.a(gate425inter11), .b(gate425inter6), .O(gate425inter12));
  nand2 gate1946(.a(gate425inter12), .b(gate425inter1), .O(G1234));
nand2 gate426( .a(G1045), .b(G1141), .O(G1235) );

  xor2  gate1597(.a(G1144), .b(G5), .O(gate427inter0));
  nand2 gate1598(.a(gate427inter0), .b(s_150), .O(gate427inter1));
  and2  gate1599(.a(G1144), .b(G5), .O(gate427inter2));
  inv1  gate1600(.a(s_150), .O(gate427inter3));
  inv1  gate1601(.a(s_151), .O(gate427inter4));
  nand2 gate1602(.a(gate427inter4), .b(gate427inter3), .O(gate427inter5));
  nor2  gate1603(.a(gate427inter5), .b(gate427inter2), .O(gate427inter6));
  inv1  gate1604(.a(G5), .O(gate427inter7));
  inv1  gate1605(.a(G1144), .O(gate427inter8));
  nand2 gate1606(.a(gate427inter8), .b(gate427inter7), .O(gate427inter9));
  nand2 gate1607(.a(s_151), .b(gate427inter3), .O(gate427inter10));
  nor2  gate1608(.a(gate427inter10), .b(gate427inter9), .O(gate427inter11));
  nor2  gate1609(.a(gate427inter11), .b(gate427inter6), .O(gate427inter12));
  nand2 gate1610(.a(gate427inter12), .b(gate427inter1), .O(G1236));
nand2 gate428( .a(G1048), .b(G1144), .O(G1237) );
nand2 gate429( .a(G6), .b(G1147), .O(G1238) );
nand2 gate430( .a(G1051), .b(G1147), .O(G1239) );
nand2 gate431( .a(G7), .b(G1150), .O(G1240) );
nand2 gate432( .a(G1054), .b(G1150), .O(G1241) );
nand2 gate433( .a(G8), .b(G1153), .O(G1242) );
nand2 gate434( .a(G1057), .b(G1153), .O(G1243) );
nand2 gate435( .a(G9), .b(G1156), .O(G1244) );
nand2 gate436( .a(G1060), .b(G1156), .O(G1245) );
nand2 gate437( .a(G10), .b(G1159), .O(G1246) );
nand2 gate438( .a(G1063), .b(G1159), .O(G1247) );

  xor2  gate813(.a(G1162), .b(G11), .O(gate439inter0));
  nand2 gate814(.a(gate439inter0), .b(s_38), .O(gate439inter1));
  and2  gate815(.a(G1162), .b(G11), .O(gate439inter2));
  inv1  gate816(.a(s_38), .O(gate439inter3));
  inv1  gate817(.a(s_39), .O(gate439inter4));
  nand2 gate818(.a(gate439inter4), .b(gate439inter3), .O(gate439inter5));
  nor2  gate819(.a(gate439inter5), .b(gate439inter2), .O(gate439inter6));
  inv1  gate820(.a(G11), .O(gate439inter7));
  inv1  gate821(.a(G1162), .O(gate439inter8));
  nand2 gate822(.a(gate439inter8), .b(gate439inter7), .O(gate439inter9));
  nand2 gate823(.a(s_39), .b(gate439inter3), .O(gate439inter10));
  nor2  gate824(.a(gate439inter10), .b(gate439inter9), .O(gate439inter11));
  nor2  gate825(.a(gate439inter11), .b(gate439inter6), .O(gate439inter12));
  nand2 gate826(.a(gate439inter12), .b(gate439inter1), .O(G1248));

  xor2  gate939(.a(G1162), .b(G1066), .O(gate440inter0));
  nand2 gate940(.a(gate440inter0), .b(s_56), .O(gate440inter1));
  and2  gate941(.a(G1162), .b(G1066), .O(gate440inter2));
  inv1  gate942(.a(s_56), .O(gate440inter3));
  inv1  gate943(.a(s_57), .O(gate440inter4));
  nand2 gate944(.a(gate440inter4), .b(gate440inter3), .O(gate440inter5));
  nor2  gate945(.a(gate440inter5), .b(gate440inter2), .O(gate440inter6));
  inv1  gate946(.a(G1066), .O(gate440inter7));
  inv1  gate947(.a(G1162), .O(gate440inter8));
  nand2 gate948(.a(gate440inter8), .b(gate440inter7), .O(gate440inter9));
  nand2 gate949(.a(s_57), .b(gate440inter3), .O(gate440inter10));
  nor2  gate950(.a(gate440inter10), .b(gate440inter9), .O(gate440inter11));
  nor2  gate951(.a(gate440inter11), .b(gate440inter6), .O(gate440inter12));
  nand2 gate952(.a(gate440inter12), .b(gate440inter1), .O(G1249));

  xor2  gate2437(.a(G1165), .b(G12), .O(gate441inter0));
  nand2 gate2438(.a(gate441inter0), .b(s_270), .O(gate441inter1));
  and2  gate2439(.a(G1165), .b(G12), .O(gate441inter2));
  inv1  gate2440(.a(s_270), .O(gate441inter3));
  inv1  gate2441(.a(s_271), .O(gate441inter4));
  nand2 gate2442(.a(gate441inter4), .b(gate441inter3), .O(gate441inter5));
  nor2  gate2443(.a(gate441inter5), .b(gate441inter2), .O(gate441inter6));
  inv1  gate2444(.a(G12), .O(gate441inter7));
  inv1  gate2445(.a(G1165), .O(gate441inter8));
  nand2 gate2446(.a(gate441inter8), .b(gate441inter7), .O(gate441inter9));
  nand2 gate2447(.a(s_271), .b(gate441inter3), .O(gate441inter10));
  nor2  gate2448(.a(gate441inter10), .b(gate441inter9), .O(gate441inter11));
  nor2  gate2449(.a(gate441inter11), .b(gate441inter6), .O(gate441inter12));
  nand2 gate2450(.a(gate441inter12), .b(gate441inter1), .O(G1250));
nand2 gate442( .a(G1069), .b(G1165), .O(G1251) );

  xor2  gate2115(.a(G1168), .b(G13), .O(gate443inter0));
  nand2 gate2116(.a(gate443inter0), .b(s_224), .O(gate443inter1));
  and2  gate2117(.a(G1168), .b(G13), .O(gate443inter2));
  inv1  gate2118(.a(s_224), .O(gate443inter3));
  inv1  gate2119(.a(s_225), .O(gate443inter4));
  nand2 gate2120(.a(gate443inter4), .b(gate443inter3), .O(gate443inter5));
  nor2  gate2121(.a(gate443inter5), .b(gate443inter2), .O(gate443inter6));
  inv1  gate2122(.a(G13), .O(gate443inter7));
  inv1  gate2123(.a(G1168), .O(gate443inter8));
  nand2 gate2124(.a(gate443inter8), .b(gate443inter7), .O(gate443inter9));
  nand2 gate2125(.a(s_225), .b(gate443inter3), .O(gate443inter10));
  nor2  gate2126(.a(gate443inter10), .b(gate443inter9), .O(gate443inter11));
  nor2  gate2127(.a(gate443inter11), .b(gate443inter6), .O(gate443inter12));
  nand2 gate2128(.a(gate443inter12), .b(gate443inter1), .O(G1252));

  xor2  gate1975(.a(G1168), .b(G1072), .O(gate444inter0));
  nand2 gate1976(.a(gate444inter0), .b(s_204), .O(gate444inter1));
  and2  gate1977(.a(G1168), .b(G1072), .O(gate444inter2));
  inv1  gate1978(.a(s_204), .O(gate444inter3));
  inv1  gate1979(.a(s_205), .O(gate444inter4));
  nand2 gate1980(.a(gate444inter4), .b(gate444inter3), .O(gate444inter5));
  nor2  gate1981(.a(gate444inter5), .b(gate444inter2), .O(gate444inter6));
  inv1  gate1982(.a(G1072), .O(gate444inter7));
  inv1  gate1983(.a(G1168), .O(gate444inter8));
  nand2 gate1984(.a(gate444inter8), .b(gate444inter7), .O(gate444inter9));
  nand2 gate1985(.a(s_205), .b(gate444inter3), .O(gate444inter10));
  nor2  gate1986(.a(gate444inter10), .b(gate444inter9), .O(gate444inter11));
  nor2  gate1987(.a(gate444inter11), .b(gate444inter6), .O(gate444inter12));
  nand2 gate1988(.a(gate444inter12), .b(gate444inter1), .O(G1253));

  xor2  gate1947(.a(G1171), .b(G14), .O(gate445inter0));
  nand2 gate1948(.a(gate445inter0), .b(s_200), .O(gate445inter1));
  and2  gate1949(.a(G1171), .b(G14), .O(gate445inter2));
  inv1  gate1950(.a(s_200), .O(gate445inter3));
  inv1  gate1951(.a(s_201), .O(gate445inter4));
  nand2 gate1952(.a(gate445inter4), .b(gate445inter3), .O(gate445inter5));
  nor2  gate1953(.a(gate445inter5), .b(gate445inter2), .O(gate445inter6));
  inv1  gate1954(.a(G14), .O(gate445inter7));
  inv1  gate1955(.a(G1171), .O(gate445inter8));
  nand2 gate1956(.a(gate445inter8), .b(gate445inter7), .O(gate445inter9));
  nand2 gate1957(.a(s_201), .b(gate445inter3), .O(gate445inter10));
  nor2  gate1958(.a(gate445inter10), .b(gate445inter9), .O(gate445inter11));
  nor2  gate1959(.a(gate445inter11), .b(gate445inter6), .O(gate445inter12));
  nand2 gate1960(.a(gate445inter12), .b(gate445inter1), .O(G1254));
nand2 gate446( .a(G1075), .b(G1171), .O(G1255) );

  xor2  gate1653(.a(G1174), .b(G15), .O(gate447inter0));
  nand2 gate1654(.a(gate447inter0), .b(s_158), .O(gate447inter1));
  and2  gate1655(.a(G1174), .b(G15), .O(gate447inter2));
  inv1  gate1656(.a(s_158), .O(gate447inter3));
  inv1  gate1657(.a(s_159), .O(gate447inter4));
  nand2 gate1658(.a(gate447inter4), .b(gate447inter3), .O(gate447inter5));
  nor2  gate1659(.a(gate447inter5), .b(gate447inter2), .O(gate447inter6));
  inv1  gate1660(.a(G15), .O(gate447inter7));
  inv1  gate1661(.a(G1174), .O(gate447inter8));
  nand2 gate1662(.a(gate447inter8), .b(gate447inter7), .O(gate447inter9));
  nand2 gate1663(.a(s_159), .b(gate447inter3), .O(gate447inter10));
  nor2  gate1664(.a(gate447inter10), .b(gate447inter9), .O(gate447inter11));
  nor2  gate1665(.a(gate447inter11), .b(gate447inter6), .O(gate447inter12));
  nand2 gate1666(.a(gate447inter12), .b(gate447inter1), .O(G1256));
nand2 gate448( .a(G1078), .b(G1174), .O(G1257) );
nand2 gate449( .a(G16), .b(G1177), .O(G1258) );
nand2 gate450( .a(G1081), .b(G1177), .O(G1259) );
nand2 gate451( .a(G17), .b(G1180), .O(G1260) );
nand2 gate452( .a(G1084), .b(G1180), .O(G1261) );

  xor2  gate547(.a(G1183), .b(G18), .O(gate453inter0));
  nand2 gate548(.a(gate453inter0), .b(s_0), .O(gate453inter1));
  and2  gate549(.a(G1183), .b(G18), .O(gate453inter2));
  inv1  gate550(.a(s_0), .O(gate453inter3));
  inv1  gate551(.a(s_1), .O(gate453inter4));
  nand2 gate552(.a(gate453inter4), .b(gate453inter3), .O(gate453inter5));
  nor2  gate553(.a(gate453inter5), .b(gate453inter2), .O(gate453inter6));
  inv1  gate554(.a(G18), .O(gate453inter7));
  inv1  gate555(.a(G1183), .O(gate453inter8));
  nand2 gate556(.a(gate453inter8), .b(gate453inter7), .O(gate453inter9));
  nand2 gate557(.a(s_1), .b(gate453inter3), .O(gate453inter10));
  nor2  gate558(.a(gate453inter10), .b(gate453inter9), .O(gate453inter11));
  nor2  gate559(.a(gate453inter11), .b(gate453inter6), .O(gate453inter12));
  nand2 gate560(.a(gate453inter12), .b(gate453inter1), .O(G1262));
nand2 gate454( .a(G1087), .b(G1183), .O(G1263) );
nand2 gate455( .a(G19), .b(G1186), .O(G1264) );
nand2 gate456( .a(G1090), .b(G1186), .O(G1265) );
nand2 gate457( .a(G20), .b(G1189), .O(G1266) );

  xor2  gate911(.a(G1189), .b(G1093), .O(gate458inter0));
  nand2 gate912(.a(gate458inter0), .b(s_52), .O(gate458inter1));
  and2  gate913(.a(G1189), .b(G1093), .O(gate458inter2));
  inv1  gate914(.a(s_52), .O(gate458inter3));
  inv1  gate915(.a(s_53), .O(gate458inter4));
  nand2 gate916(.a(gate458inter4), .b(gate458inter3), .O(gate458inter5));
  nor2  gate917(.a(gate458inter5), .b(gate458inter2), .O(gate458inter6));
  inv1  gate918(.a(G1093), .O(gate458inter7));
  inv1  gate919(.a(G1189), .O(gate458inter8));
  nand2 gate920(.a(gate458inter8), .b(gate458inter7), .O(gate458inter9));
  nand2 gate921(.a(s_53), .b(gate458inter3), .O(gate458inter10));
  nor2  gate922(.a(gate458inter10), .b(gate458inter9), .O(gate458inter11));
  nor2  gate923(.a(gate458inter11), .b(gate458inter6), .O(gate458inter12));
  nand2 gate924(.a(gate458inter12), .b(gate458inter1), .O(G1267));

  xor2  gate1261(.a(G1192), .b(G21), .O(gate459inter0));
  nand2 gate1262(.a(gate459inter0), .b(s_102), .O(gate459inter1));
  and2  gate1263(.a(G1192), .b(G21), .O(gate459inter2));
  inv1  gate1264(.a(s_102), .O(gate459inter3));
  inv1  gate1265(.a(s_103), .O(gate459inter4));
  nand2 gate1266(.a(gate459inter4), .b(gate459inter3), .O(gate459inter5));
  nor2  gate1267(.a(gate459inter5), .b(gate459inter2), .O(gate459inter6));
  inv1  gate1268(.a(G21), .O(gate459inter7));
  inv1  gate1269(.a(G1192), .O(gate459inter8));
  nand2 gate1270(.a(gate459inter8), .b(gate459inter7), .O(gate459inter9));
  nand2 gate1271(.a(s_103), .b(gate459inter3), .O(gate459inter10));
  nor2  gate1272(.a(gate459inter10), .b(gate459inter9), .O(gate459inter11));
  nor2  gate1273(.a(gate459inter11), .b(gate459inter6), .O(gate459inter12));
  nand2 gate1274(.a(gate459inter12), .b(gate459inter1), .O(G1268));

  xor2  gate1709(.a(G1192), .b(G1096), .O(gate460inter0));
  nand2 gate1710(.a(gate460inter0), .b(s_166), .O(gate460inter1));
  and2  gate1711(.a(G1192), .b(G1096), .O(gate460inter2));
  inv1  gate1712(.a(s_166), .O(gate460inter3));
  inv1  gate1713(.a(s_167), .O(gate460inter4));
  nand2 gate1714(.a(gate460inter4), .b(gate460inter3), .O(gate460inter5));
  nor2  gate1715(.a(gate460inter5), .b(gate460inter2), .O(gate460inter6));
  inv1  gate1716(.a(G1096), .O(gate460inter7));
  inv1  gate1717(.a(G1192), .O(gate460inter8));
  nand2 gate1718(.a(gate460inter8), .b(gate460inter7), .O(gate460inter9));
  nand2 gate1719(.a(s_167), .b(gate460inter3), .O(gate460inter10));
  nor2  gate1720(.a(gate460inter10), .b(gate460inter9), .O(gate460inter11));
  nor2  gate1721(.a(gate460inter11), .b(gate460inter6), .O(gate460inter12));
  nand2 gate1722(.a(gate460inter12), .b(gate460inter1), .O(G1269));
nand2 gate461( .a(G22), .b(G1195), .O(G1270) );
nand2 gate462( .a(G1099), .b(G1195), .O(G1271) );
nand2 gate463( .a(G23), .b(G1198), .O(G1272) );
nand2 gate464( .a(G1102), .b(G1198), .O(G1273) );
nand2 gate465( .a(G24), .b(G1201), .O(G1274) );
nand2 gate466( .a(G1105), .b(G1201), .O(G1275) );

  xor2  gate1527(.a(G1204), .b(G25), .O(gate467inter0));
  nand2 gate1528(.a(gate467inter0), .b(s_140), .O(gate467inter1));
  and2  gate1529(.a(G1204), .b(G25), .O(gate467inter2));
  inv1  gate1530(.a(s_140), .O(gate467inter3));
  inv1  gate1531(.a(s_141), .O(gate467inter4));
  nand2 gate1532(.a(gate467inter4), .b(gate467inter3), .O(gate467inter5));
  nor2  gate1533(.a(gate467inter5), .b(gate467inter2), .O(gate467inter6));
  inv1  gate1534(.a(G25), .O(gate467inter7));
  inv1  gate1535(.a(G1204), .O(gate467inter8));
  nand2 gate1536(.a(gate467inter8), .b(gate467inter7), .O(gate467inter9));
  nand2 gate1537(.a(s_141), .b(gate467inter3), .O(gate467inter10));
  nor2  gate1538(.a(gate467inter10), .b(gate467inter9), .O(gate467inter11));
  nor2  gate1539(.a(gate467inter11), .b(gate467inter6), .O(gate467inter12));
  nand2 gate1540(.a(gate467inter12), .b(gate467inter1), .O(G1276));
nand2 gate468( .a(G1108), .b(G1204), .O(G1277) );
nand2 gate469( .a(G26), .b(G1207), .O(G1278) );
nand2 gate470( .a(G1111), .b(G1207), .O(G1279) );

  xor2  gate1765(.a(G1210), .b(G27), .O(gate471inter0));
  nand2 gate1766(.a(gate471inter0), .b(s_174), .O(gate471inter1));
  and2  gate1767(.a(G1210), .b(G27), .O(gate471inter2));
  inv1  gate1768(.a(s_174), .O(gate471inter3));
  inv1  gate1769(.a(s_175), .O(gate471inter4));
  nand2 gate1770(.a(gate471inter4), .b(gate471inter3), .O(gate471inter5));
  nor2  gate1771(.a(gate471inter5), .b(gate471inter2), .O(gate471inter6));
  inv1  gate1772(.a(G27), .O(gate471inter7));
  inv1  gate1773(.a(G1210), .O(gate471inter8));
  nand2 gate1774(.a(gate471inter8), .b(gate471inter7), .O(gate471inter9));
  nand2 gate1775(.a(s_175), .b(gate471inter3), .O(gate471inter10));
  nor2  gate1776(.a(gate471inter10), .b(gate471inter9), .O(gate471inter11));
  nor2  gate1777(.a(gate471inter11), .b(gate471inter6), .O(gate471inter12));
  nand2 gate1778(.a(gate471inter12), .b(gate471inter1), .O(G1280));

  xor2  gate1051(.a(G1210), .b(G1114), .O(gate472inter0));
  nand2 gate1052(.a(gate472inter0), .b(s_72), .O(gate472inter1));
  and2  gate1053(.a(G1210), .b(G1114), .O(gate472inter2));
  inv1  gate1054(.a(s_72), .O(gate472inter3));
  inv1  gate1055(.a(s_73), .O(gate472inter4));
  nand2 gate1056(.a(gate472inter4), .b(gate472inter3), .O(gate472inter5));
  nor2  gate1057(.a(gate472inter5), .b(gate472inter2), .O(gate472inter6));
  inv1  gate1058(.a(G1114), .O(gate472inter7));
  inv1  gate1059(.a(G1210), .O(gate472inter8));
  nand2 gate1060(.a(gate472inter8), .b(gate472inter7), .O(gate472inter9));
  nand2 gate1061(.a(s_73), .b(gate472inter3), .O(gate472inter10));
  nor2  gate1062(.a(gate472inter10), .b(gate472inter9), .O(gate472inter11));
  nor2  gate1063(.a(gate472inter11), .b(gate472inter6), .O(gate472inter12));
  nand2 gate1064(.a(gate472inter12), .b(gate472inter1), .O(G1281));

  xor2  gate925(.a(G1213), .b(G28), .O(gate473inter0));
  nand2 gate926(.a(gate473inter0), .b(s_54), .O(gate473inter1));
  and2  gate927(.a(G1213), .b(G28), .O(gate473inter2));
  inv1  gate928(.a(s_54), .O(gate473inter3));
  inv1  gate929(.a(s_55), .O(gate473inter4));
  nand2 gate930(.a(gate473inter4), .b(gate473inter3), .O(gate473inter5));
  nor2  gate931(.a(gate473inter5), .b(gate473inter2), .O(gate473inter6));
  inv1  gate932(.a(G28), .O(gate473inter7));
  inv1  gate933(.a(G1213), .O(gate473inter8));
  nand2 gate934(.a(gate473inter8), .b(gate473inter7), .O(gate473inter9));
  nand2 gate935(.a(s_55), .b(gate473inter3), .O(gate473inter10));
  nor2  gate936(.a(gate473inter10), .b(gate473inter9), .O(gate473inter11));
  nor2  gate937(.a(gate473inter11), .b(gate473inter6), .O(gate473inter12));
  nand2 gate938(.a(gate473inter12), .b(gate473inter1), .O(G1282));
nand2 gate474( .a(G1117), .b(G1213), .O(G1283) );
nand2 gate475( .a(G29), .b(G1216), .O(G1284) );
nand2 gate476( .a(G1120), .b(G1216), .O(G1285) );

  xor2  gate785(.a(G1219), .b(G30), .O(gate477inter0));
  nand2 gate786(.a(gate477inter0), .b(s_34), .O(gate477inter1));
  and2  gate787(.a(G1219), .b(G30), .O(gate477inter2));
  inv1  gate788(.a(s_34), .O(gate477inter3));
  inv1  gate789(.a(s_35), .O(gate477inter4));
  nand2 gate790(.a(gate477inter4), .b(gate477inter3), .O(gate477inter5));
  nor2  gate791(.a(gate477inter5), .b(gate477inter2), .O(gate477inter6));
  inv1  gate792(.a(G30), .O(gate477inter7));
  inv1  gate793(.a(G1219), .O(gate477inter8));
  nand2 gate794(.a(gate477inter8), .b(gate477inter7), .O(gate477inter9));
  nand2 gate795(.a(s_35), .b(gate477inter3), .O(gate477inter10));
  nor2  gate796(.a(gate477inter10), .b(gate477inter9), .O(gate477inter11));
  nor2  gate797(.a(gate477inter11), .b(gate477inter6), .O(gate477inter12));
  nand2 gate798(.a(gate477inter12), .b(gate477inter1), .O(G1286));

  xor2  gate1359(.a(G1219), .b(G1123), .O(gate478inter0));
  nand2 gate1360(.a(gate478inter0), .b(s_116), .O(gate478inter1));
  and2  gate1361(.a(G1219), .b(G1123), .O(gate478inter2));
  inv1  gate1362(.a(s_116), .O(gate478inter3));
  inv1  gate1363(.a(s_117), .O(gate478inter4));
  nand2 gate1364(.a(gate478inter4), .b(gate478inter3), .O(gate478inter5));
  nor2  gate1365(.a(gate478inter5), .b(gate478inter2), .O(gate478inter6));
  inv1  gate1366(.a(G1123), .O(gate478inter7));
  inv1  gate1367(.a(G1219), .O(gate478inter8));
  nand2 gate1368(.a(gate478inter8), .b(gate478inter7), .O(gate478inter9));
  nand2 gate1369(.a(s_117), .b(gate478inter3), .O(gate478inter10));
  nor2  gate1370(.a(gate478inter10), .b(gate478inter9), .O(gate478inter11));
  nor2  gate1371(.a(gate478inter11), .b(gate478inter6), .O(gate478inter12));
  nand2 gate1372(.a(gate478inter12), .b(gate478inter1), .O(G1287));
nand2 gate479( .a(G31), .b(G1222), .O(G1288) );

  xor2  gate1247(.a(G1222), .b(G1126), .O(gate480inter0));
  nand2 gate1248(.a(gate480inter0), .b(s_100), .O(gate480inter1));
  and2  gate1249(.a(G1222), .b(G1126), .O(gate480inter2));
  inv1  gate1250(.a(s_100), .O(gate480inter3));
  inv1  gate1251(.a(s_101), .O(gate480inter4));
  nand2 gate1252(.a(gate480inter4), .b(gate480inter3), .O(gate480inter5));
  nor2  gate1253(.a(gate480inter5), .b(gate480inter2), .O(gate480inter6));
  inv1  gate1254(.a(G1126), .O(gate480inter7));
  inv1  gate1255(.a(G1222), .O(gate480inter8));
  nand2 gate1256(.a(gate480inter8), .b(gate480inter7), .O(gate480inter9));
  nand2 gate1257(.a(s_101), .b(gate480inter3), .O(gate480inter10));
  nor2  gate1258(.a(gate480inter10), .b(gate480inter9), .O(gate480inter11));
  nor2  gate1259(.a(gate480inter11), .b(gate480inter6), .O(gate480inter12));
  nand2 gate1260(.a(gate480inter12), .b(gate480inter1), .O(G1289));
nand2 gate481( .a(G32), .b(G1225), .O(G1290) );

  xor2  gate1303(.a(G1225), .b(G1129), .O(gate482inter0));
  nand2 gate1304(.a(gate482inter0), .b(s_108), .O(gate482inter1));
  and2  gate1305(.a(G1225), .b(G1129), .O(gate482inter2));
  inv1  gate1306(.a(s_108), .O(gate482inter3));
  inv1  gate1307(.a(s_109), .O(gate482inter4));
  nand2 gate1308(.a(gate482inter4), .b(gate482inter3), .O(gate482inter5));
  nor2  gate1309(.a(gate482inter5), .b(gate482inter2), .O(gate482inter6));
  inv1  gate1310(.a(G1129), .O(gate482inter7));
  inv1  gate1311(.a(G1225), .O(gate482inter8));
  nand2 gate1312(.a(gate482inter8), .b(gate482inter7), .O(gate482inter9));
  nand2 gate1313(.a(s_109), .b(gate482inter3), .O(gate482inter10));
  nor2  gate1314(.a(gate482inter10), .b(gate482inter9), .O(gate482inter11));
  nor2  gate1315(.a(gate482inter11), .b(gate482inter6), .O(gate482inter12));
  nand2 gate1316(.a(gate482inter12), .b(gate482inter1), .O(G1291));
nand2 gate483( .a(G1228), .b(G1229), .O(G1292) );
nand2 gate484( .a(G1230), .b(G1231), .O(G1293) );

  xor2  gate2227(.a(G1233), .b(G1232), .O(gate485inter0));
  nand2 gate2228(.a(gate485inter0), .b(s_240), .O(gate485inter1));
  and2  gate2229(.a(G1233), .b(G1232), .O(gate485inter2));
  inv1  gate2230(.a(s_240), .O(gate485inter3));
  inv1  gate2231(.a(s_241), .O(gate485inter4));
  nand2 gate2232(.a(gate485inter4), .b(gate485inter3), .O(gate485inter5));
  nor2  gate2233(.a(gate485inter5), .b(gate485inter2), .O(gate485inter6));
  inv1  gate2234(.a(G1232), .O(gate485inter7));
  inv1  gate2235(.a(G1233), .O(gate485inter8));
  nand2 gate2236(.a(gate485inter8), .b(gate485inter7), .O(gate485inter9));
  nand2 gate2237(.a(s_241), .b(gate485inter3), .O(gate485inter10));
  nor2  gate2238(.a(gate485inter10), .b(gate485inter9), .O(gate485inter11));
  nor2  gate2239(.a(gate485inter11), .b(gate485inter6), .O(gate485inter12));
  nand2 gate2240(.a(gate485inter12), .b(gate485inter1), .O(G1294));
nand2 gate486( .a(G1234), .b(G1235), .O(G1295) );
nand2 gate487( .a(G1236), .b(G1237), .O(G1296) );
nand2 gate488( .a(G1238), .b(G1239), .O(G1297) );
nand2 gate489( .a(G1240), .b(G1241), .O(G1298) );

  xor2  gate659(.a(G1243), .b(G1242), .O(gate490inter0));
  nand2 gate660(.a(gate490inter0), .b(s_16), .O(gate490inter1));
  and2  gate661(.a(G1243), .b(G1242), .O(gate490inter2));
  inv1  gate662(.a(s_16), .O(gate490inter3));
  inv1  gate663(.a(s_17), .O(gate490inter4));
  nand2 gate664(.a(gate490inter4), .b(gate490inter3), .O(gate490inter5));
  nor2  gate665(.a(gate490inter5), .b(gate490inter2), .O(gate490inter6));
  inv1  gate666(.a(G1242), .O(gate490inter7));
  inv1  gate667(.a(G1243), .O(gate490inter8));
  nand2 gate668(.a(gate490inter8), .b(gate490inter7), .O(gate490inter9));
  nand2 gate669(.a(s_17), .b(gate490inter3), .O(gate490inter10));
  nor2  gate670(.a(gate490inter10), .b(gate490inter9), .O(gate490inter11));
  nor2  gate671(.a(gate490inter11), .b(gate490inter6), .O(gate490inter12));
  nand2 gate672(.a(gate490inter12), .b(gate490inter1), .O(G1299));
nand2 gate491( .a(G1244), .b(G1245), .O(G1300) );
nand2 gate492( .a(G1246), .b(G1247), .O(G1301) );
nand2 gate493( .a(G1248), .b(G1249), .O(G1302) );
nand2 gate494( .a(G1250), .b(G1251), .O(G1303) );

  xor2  gate1457(.a(G1253), .b(G1252), .O(gate495inter0));
  nand2 gate1458(.a(gate495inter0), .b(s_130), .O(gate495inter1));
  and2  gate1459(.a(G1253), .b(G1252), .O(gate495inter2));
  inv1  gate1460(.a(s_130), .O(gate495inter3));
  inv1  gate1461(.a(s_131), .O(gate495inter4));
  nand2 gate1462(.a(gate495inter4), .b(gate495inter3), .O(gate495inter5));
  nor2  gate1463(.a(gate495inter5), .b(gate495inter2), .O(gate495inter6));
  inv1  gate1464(.a(G1252), .O(gate495inter7));
  inv1  gate1465(.a(G1253), .O(gate495inter8));
  nand2 gate1466(.a(gate495inter8), .b(gate495inter7), .O(gate495inter9));
  nand2 gate1467(.a(s_131), .b(gate495inter3), .O(gate495inter10));
  nor2  gate1468(.a(gate495inter10), .b(gate495inter9), .O(gate495inter11));
  nor2  gate1469(.a(gate495inter11), .b(gate495inter6), .O(gate495inter12));
  nand2 gate1470(.a(gate495inter12), .b(gate495inter1), .O(G1304));
nand2 gate496( .a(G1254), .b(G1255), .O(G1305) );

  xor2  gate1961(.a(G1257), .b(G1256), .O(gate497inter0));
  nand2 gate1962(.a(gate497inter0), .b(s_202), .O(gate497inter1));
  and2  gate1963(.a(G1257), .b(G1256), .O(gate497inter2));
  inv1  gate1964(.a(s_202), .O(gate497inter3));
  inv1  gate1965(.a(s_203), .O(gate497inter4));
  nand2 gate1966(.a(gate497inter4), .b(gate497inter3), .O(gate497inter5));
  nor2  gate1967(.a(gate497inter5), .b(gate497inter2), .O(gate497inter6));
  inv1  gate1968(.a(G1256), .O(gate497inter7));
  inv1  gate1969(.a(G1257), .O(gate497inter8));
  nand2 gate1970(.a(gate497inter8), .b(gate497inter7), .O(gate497inter9));
  nand2 gate1971(.a(s_203), .b(gate497inter3), .O(gate497inter10));
  nor2  gate1972(.a(gate497inter10), .b(gate497inter9), .O(gate497inter11));
  nor2  gate1973(.a(gate497inter11), .b(gate497inter6), .O(gate497inter12));
  nand2 gate1974(.a(gate497inter12), .b(gate497inter1), .O(G1306));

  xor2  gate1065(.a(G1259), .b(G1258), .O(gate498inter0));
  nand2 gate1066(.a(gate498inter0), .b(s_74), .O(gate498inter1));
  and2  gate1067(.a(G1259), .b(G1258), .O(gate498inter2));
  inv1  gate1068(.a(s_74), .O(gate498inter3));
  inv1  gate1069(.a(s_75), .O(gate498inter4));
  nand2 gate1070(.a(gate498inter4), .b(gate498inter3), .O(gate498inter5));
  nor2  gate1071(.a(gate498inter5), .b(gate498inter2), .O(gate498inter6));
  inv1  gate1072(.a(G1258), .O(gate498inter7));
  inv1  gate1073(.a(G1259), .O(gate498inter8));
  nand2 gate1074(.a(gate498inter8), .b(gate498inter7), .O(gate498inter9));
  nand2 gate1075(.a(s_75), .b(gate498inter3), .O(gate498inter10));
  nor2  gate1076(.a(gate498inter10), .b(gate498inter9), .O(gate498inter11));
  nor2  gate1077(.a(gate498inter11), .b(gate498inter6), .O(gate498inter12));
  nand2 gate1078(.a(gate498inter12), .b(gate498inter1), .O(G1307));
nand2 gate499( .a(G1260), .b(G1261), .O(G1308) );

  xor2  gate1863(.a(G1263), .b(G1262), .O(gate500inter0));
  nand2 gate1864(.a(gate500inter0), .b(s_188), .O(gate500inter1));
  and2  gate1865(.a(G1263), .b(G1262), .O(gate500inter2));
  inv1  gate1866(.a(s_188), .O(gate500inter3));
  inv1  gate1867(.a(s_189), .O(gate500inter4));
  nand2 gate1868(.a(gate500inter4), .b(gate500inter3), .O(gate500inter5));
  nor2  gate1869(.a(gate500inter5), .b(gate500inter2), .O(gate500inter6));
  inv1  gate1870(.a(G1262), .O(gate500inter7));
  inv1  gate1871(.a(G1263), .O(gate500inter8));
  nand2 gate1872(.a(gate500inter8), .b(gate500inter7), .O(gate500inter9));
  nand2 gate1873(.a(s_189), .b(gate500inter3), .O(gate500inter10));
  nor2  gate1874(.a(gate500inter10), .b(gate500inter9), .O(gate500inter11));
  nor2  gate1875(.a(gate500inter11), .b(gate500inter6), .O(gate500inter12));
  nand2 gate1876(.a(gate500inter12), .b(gate500inter1), .O(G1309));
nand2 gate501( .a(G1264), .b(G1265), .O(G1310) );
nand2 gate502( .a(G1266), .b(G1267), .O(G1311) );

  xor2  gate1877(.a(G1269), .b(G1268), .O(gate503inter0));
  nand2 gate1878(.a(gate503inter0), .b(s_190), .O(gate503inter1));
  and2  gate1879(.a(G1269), .b(G1268), .O(gate503inter2));
  inv1  gate1880(.a(s_190), .O(gate503inter3));
  inv1  gate1881(.a(s_191), .O(gate503inter4));
  nand2 gate1882(.a(gate503inter4), .b(gate503inter3), .O(gate503inter5));
  nor2  gate1883(.a(gate503inter5), .b(gate503inter2), .O(gate503inter6));
  inv1  gate1884(.a(G1268), .O(gate503inter7));
  inv1  gate1885(.a(G1269), .O(gate503inter8));
  nand2 gate1886(.a(gate503inter8), .b(gate503inter7), .O(gate503inter9));
  nand2 gate1887(.a(s_191), .b(gate503inter3), .O(gate503inter10));
  nor2  gate1888(.a(gate503inter10), .b(gate503inter9), .O(gate503inter11));
  nor2  gate1889(.a(gate503inter11), .b(gate503inter6), .O(gate503inter12));
  nand2 gate1890(.a(gate503inter12), .b(gate503inter1), .O(G1312));
nand2 gate504( .a(G1270), .b(G1271), .O(G1313) );
nand2 gate505( .a(G1272), .b(G1273), .O(G1314) );
nand2 gate506( .a(G1274), .b(G1275), .O(G1315) );

  xor2  gate1135(.a(G1277), .b(G1276), .O(gate507inter0));
  nand2 gate1136(.a(gate507inter0), .b(s_84), .O(gate507inter1));
  and2  gate1137(.a(G1277), .b(G1276), .O(gate507inter2));
  inv1  gate1138(.a(s_84), .O(gate507inter3));
  inv1  gate1139(.a(s_85), .O(gate507inter4));
  nand2 gate1140(.a(gate507inter4), .b(gate507inter3), .O(gate507inter5));
  nor2  gate1141(.a(gate507inter5), .b(gate507inter2), .O(gate507inter6));
  inv1  gate1142(.a(G1276), .O(gate507inter7));
  inv1  gate1143(.a(G1277), .O(gate507inter8));
  nand2 gate1144(.a(gate507inter8), .b(gate507inter7), .O(gate507inter9));
  nand2 gate1145(.a(s_85), .b(gate507inter3), .O(gate507inter10));
  nor2  gate1146(.a(gate507inter10), .b(gate507inter9), .O(gate507inter11));
  nor2  gate1147(.a(gate507inter11), .b(gate507inter6), .O(gate507inter12));
  nand2 gate1148(.a(gate507inter12), .b(gate507inter1), .O(G1316));
nand2 gate508( .a(G1278), .b(G1279), .O(G1317) );
nand2 gate509( .a(G1280), .b(G1281), .O(G1318) );

  xor2  gate1107(.a(G1283), .b(G1282), .O(gate510inter0));
  nand2 gate1108(.a(gate510inter0), .b(s_80), .O(gate510inter1));
  and2  gate1109(.a(G1283), .b(G1282), .O(gate510inter2));
  inv1  gate1110(.a(s_80), .O(gate510inter3));
  inv1  gate1111(.a(s_81), .O(gate510inter4));
  nand2 gate1112(.a(gate510inter4), .b(gate510inter3), .O(gate510inter5));
  nor2  gate1113(.a(gate510inter5), .b(gate510inter2), .O(gate510inter6));
  inv1  gate1114(.a(G1282), .O(gate510inter7));
  inv1  gate1115(.a(G1283), .O(gate510inter8));
  nand2 gate1116(.a(gate510inter8), .b(gate510inter7), .O(gate510inter9));
  nand2 gate1117(.a(s_81), .b(gate510inter3), .O(gate510inter10));
  nor2  gate1118(.a(gate510inter10), .b(gate510inter9), .O(gate510inter11));
  nor2  gate1119(.a(gate510inter11), .b(gate510inter6), .O(gate510inter12));
  nand2 gate1120(.a(gate510inter12), .b(gate510inter1), .O(G1319));
nand2 gate511( .a(G1284), .b(G1285), .O(G1320) );
nand2 gate512( .a(G1286), .b(G1287), .O(G1321) );

  xor2  gate2381(.a(G1289), .b(G1288), .O(gate513inter0));
  nand2 gate2382(.a(gate513inter0), .b(s_262), .O(gate513inter1));
  and2  gate2383(.a(G1289), .b(G1288), .O(gate513inter2));
  inv1  gate2384(.a(s_262), .O(gate513inter3));
  inv1  gate2385(.a(s_263), .O(gate513inter4));
  nand2 gate2386(.a(gate513inter4), .b(gate513inter3), .O(gate513inter5));
  nor2  gate2387(.a(gate513inter5), .b(gate513inter2), .O(gate513inter6));
  inv1  gate2388(.a(G1288), .O(gate513inter7));
  inv1  gate2389(.a(G1289), .O(gate513inter8));
  nand2 gate2390(.a(gate513inter8), .b(gate513inter7), .O(gate513inter9));
  nand2 gate2391(.a(s_263), .b(gate513inter3), .O(gate513inter10));
  nor2  gate2392(.a(gate513inter10), .b(gate513inter9), .O(gate513inter11));
  nor2  gate2393(.a(gate513inter11), .b(gate513inter6), .O(gate513inter12));
  nand2 gate2394(.a(gate513inter12), .b(gate513inter1), .O(G1322));

  xor2  gate1625(.a(G1291), .b(G1290), .O(gate514inter0));
  nand2 gate1626(.a(gate514inter0), .b(s_154), .O(gate514inter1));
  and2  gate1627(.a(G1291), .b(G1290), .O(gate514inter2));
  inv1  gate1628(.a(s_154), .O(gate514inter3));
  inv1  gate1629(.a(s_155), .O(gate514inter4));
  nand2 gate1630(.a(gate514inter4), .b(gate514inter3), .O(gate514inter5));
  nor2  gate1631(.a(gate514inter5), .b(gate514inter2), .O(gate514inter6));
  inv1  gate1632(.a(G1290), .O(gate514inter7));
  inv1  gate1633(.a(G1291), .O(gate514inter8));
  nand2 gate1634(.a(gate514inter8), .b(gate514inter7), .O(gate514inter9));
  nand2 gate1635(.a(s_155), .b(gate514inter3), .O(gate514inter10));
  nor2  gate1636(.a(gate514inter10), .b(gate514inter9), .O(gate514inter11));
  nor2  gate1637(.a(gate514inter11), .b(gate514inter6), .O(gate514inter12));
  nand2 gate1638(.a(gate514inter12), .b(gate514inter1), .O(G1323));
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule