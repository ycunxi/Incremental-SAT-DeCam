module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);

input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;//RE__PI;

input s_0,s_1;//RE__ALLOW(00,01,10,11);
input s_2,s_3;//RE__ALLOW(00,01,10,11);
input s_4,s_5;//RE__ALLOW(00,01,10,11);
input s_6,s_7;//RE__ALLOW(00,01,10,11);
input s_8,s_9;//RE__ALLOW(00,01,10,11);
input s_10,s_11;//RE__ALLOW(00,01,10,11);
input s_12,s_13;//RE__ALLOW(00,01,10,11);
input s_14,s_15;//RE__ALLOW(00,01,10,11);
input s_16,s_17;//RE__ALLOW(00,01,10,11);
input s_18,s_19;//RE__ALLOW(00,01,10,11);
input s_20,s_21;//RE__ALLOW(00,01,10,11);
input s_22,s_23;//RE__ALLOW(00,01,10,11);
input s_24,s_25;//RE__ALLOW(00,01,10,11);
input s_26,s_27;//RE__ALLOW(00,01,10,11);
input s_28,s_29;//RE__ALLOW(00,01,10,11);
input s_30,s_31;//RE__ALLOW(00,01,10,11);
input s_32,s_33;//RE__ALLOW(00,01,10,11);
input s_34,s_35;//RE__ALLOW(00,01,10,11);
input s_36,s_37;//RE__ALLOW(00,01,10,11);
input s_38,s_39;//RE__ALLOW(00,01,10,11);
input s_40,s_41;//RE__ALLOW(00,01,10,11);
input s_42,s_43;//RE__ALLOW(00,01,10,11);
input s_44,s_45;//RE__ALLOW(00,01,10,11);
input s_46,s_47;//RE__ALLOW(00,01,10,11);
input s_48,s_49;//RE__ALLOW(00,01,10,11);
input s_50,s_51;//RE__ALLOW(00,01,10,11);
input s_52,s_53;//RE__ALLOW(00,01,10,11);
input s_54,s_55;//RE__ALLOW(00,01,10,11);
input s_56,s_57;//RE__ALLOW(00,01,10,11);
input s_58,s_59;//RE__ALLOW(00,01,10,11);
input s_60,s_61;//RE__ALLOW(00,01,10,11);
input s_62,s_63;//RE__ALLOW(00,01,10,11);
input s_64,s_65;//RE__ALLOW(00,01,10,11);
input s_66,s_67;//RE__ALLOW(00,01,10,11);
input s_68,s_69;//RE__ALLOW(00,01,10,11);
input s_70,s_71;//RE__ALLOW(00,01,10,11);
input s_72,s_73;//RE__ALLOW(00,01,10,11);
input s_74,s_75;//RE__ALLOW(00,01,10,11);
input s_76,s_77;//RE__ALLOW(00,01,10,11);
input s_78,s_79;//RE__ALLOW(00,01,10,11);
input s_80,s_81;//RE__ALLOW(00,01,10,11);
input s_82,s_83;//RE__ALLOW(00,01,10,11);
input s_84,s_85;//RE__ALLOW(00,01,10,11);
input s_86,s_87;//RE__ALLOW(00,01,10,11);
input s_88,s_89;//RE__ALLOW(00,01,10,11);
input s_90,s_91;//RE__ALLOW(00,01,10,11);
input s_92,s_93;//RE__ALLOW(00,01,10,11);
input s_94,s_95;//RE__ALLOW(00,01,10,11);
input s_96,s_97;//RE__ALLOW(00,01,10,11);
input s_98,s_99;//RE__ALLOW(00,01,10,11);
input s_100,s_101;//RE__ALLOW(00,01,10,11);
input s_102,s_103;//RE__ALLOW(00,01,10,11);
input s_104,s_105;//RE__ALLOW(00,01,10,11);
input s_106,s_107;//RE__ALLOW(00,01,10,11);
input s_108,s_109;//RE__ALLOW(00,01,10,11);
input s_110,s_111;//RE__ALLOW(00,01,10,11);
input s_112,s_113;//RE__ALLOW(00,01,10,11);
input s_114,s_115;//RE__ALLOW(00,01,10,11);
input s_116,s_117;//RE__ALLOW(00,01,10,11);
input s_118,s_119;//RE__ALLOW(00,01,10,11);
input s_120,s_121;//RE__ALLOW(00,01,10,11);
input s_122,s_123;//RE__ALLOW(00,01,10,11);
input s_124,s_125;//RE__ALLOW(00,01,10,11);
input s_126,s_127;//RE__ALLOW(00,01,10,11);
input s_128,s_129;//RE__ALLOW(00,01,10,11);
input s_130,s_131;//RE__ALLOW(00,01,10,11);
input s_132,s_133;//RE__ALLOW(00,01,10,11);
input s_134,s_135;//RE__ALLOW(00,01,10,11);
input s_136,s_137;//RE__ALLOW(00,01,10,11);
input s_138,s_139;//RE__ALLOW(00,01,10,11);
input s_140,s_141;//RE__ALLOW(00,01,10,11);
input s_142,s_143;//RE__ALLOW(00,01,10,11);
input s_144,s_145;//RE__ALLOW(00,01,10,11);
input s_146,s_147;//RE__ALLOW(00,01,10,11);
input s_148,s_149;//RE__ALLOW(00,01,10,11);
input s_150,s_151;//RE__ALLOW(00,01,10,11);
input s_152,s_153;//RE__ALLOW(00,01,10,11);
input s_154,s_155;//RE__ALLOW(00,01,10,11);
input s_156,s_157;//RE__ALLOW(00,01,10,11);
input s_158,s_159;//RE__ALLOW(00,01,10,11);
input s_160,s_161;//RE__ALLOW(00,01,10,11);
input s_162,s_163;//RE__ALLOW(00,01,10,11);
input s_164,s_165;//RE__ALLOW(00,01,10,11);
input s_166,s_167;//RE__ALLOW(00,01,10,11);
input s_168,s_169;//RE__ALLOW(00,01,10,11);
input s_170,s_171;//RE__ALLOW(00,01,10,11);
input s_172,s_173;//RE__ALLOW(00,01,10,11);
input s_174,s_175;//RE__ALLOW(00,01,10,11);
input s_176,s_177;//RE__ALLOW(00,01,10,11);
input s_178,s_179;//RE__ALLOW(00,01,10,11);
input s_180,s_181;//RE__ALLOW(00,01,10,11);
input s_182,s_183;//RE__ALLOW(00,01,10,11);
input s_184,s_185;//RE__ALLOW(00,01,10,11);
input s_186,s_187;//RE__ALLOW(00,01,10,11);
input s_188,s_189;//RE__ALLOW(00,01,10,11);
input s_190,s_191;//RE__ALLOW(00,01,10,11);
input s_192,s_193;//RE__ALLOW(00,01,10,11);
input s_194,s_195;//RE__ALLOW(00,01,10,11);
input s_196,s_197;//RE__ALLOW(00,01,10,11);
input s_198,s_199;//RE__ALLOW(00,01,10,11);
input s_200,s_201;//RE__ALLOW(00,01,10,11);
input s_202,s_203;//RE__ALLOW(00,01,10,11);
input s_204,s_205;//RE__ALLOW(00,01,10,11);
input s_206,s_207;//RE__ALLOW(00,01,10,11);
input s_208,s_209;//RE__ALLOW(00,01,10,11);
input s_210,s_211;//RE__ALLOW(00,01,10,11);
input s_212,s_213;//RE__ALLOW(00,01,10,11);
input s_214,s_215;//RE__ALLOW(00,01,10,11);
input s_216,s_217;//RE__ALLOW(00,01,10,11);
input s_218,s_219;//RE__ALLOW(00,01,10,11);
input s_220,s_221;//RE__ALLOW(00,01,10,11);
input s_222,s_223;//RE__ALLOW(00,01,10,11);
input s_224,s_225;//RE__ALLOW(00,01,10,11);
input s_226,s_227;//RE__ALLOW(00,01,10,11);
input s_228,s_229;//RE__ALLOW(00,01,10,11);
input s_230,s_231;//RE__ALLOW(00,01,10,11);
input s_232,s_233;//RE__ALLOW(00,01,10,11);
input s_234,s_235;//RE__ALLOW(00,01,10,11);
input s_236,s_237;//RE__ALLOW(00,01,10,11);
input s_238,s_239;//RE__ALLOW(00,01,10,11);
input s_240,s_241;//RE__ALLOW(00,01,10,11);
input s_242,s_243;//RE__ALLOW(00,01,10,11);
input s_244,s_245;//RE__ALLOW(00,01,10,11);
input s_246,s_247;//RE__ALLOW(00,01,10,11);
input s_248,s_249;//RE__ALLOW(00,01,10,11);
input s_250,s_251;//RE__ALLOW(00,01,10,11);
input s_252,s_253;//RE__ALLOW(00,01,10,11);
input s_254,s_255;//RE__ALLOW(00,01,10,11);
input s_256,s_257;//RE__ALLOW(00,01,10,11);
input s_258,s_259;//RE__ALLOW(00,01,10,11);
input s_260,s_261;//RE__ALLOW(00,01,10,11);
input s_262,s_263;//RE__ALLOW(00,01,10,11);
input s_264,s_265;//RE__ALLOW(00,01,10,11);
input s_266,s_267;//RE__ALLOW(00,01,10,11);
input s_268,s_269;//RE__ALLOW(00,01,10,11);
input s_270,s_271;//RE__ALLOW(00,01,10,11);
input s_272,s_273;//RE__ALLOW(00,01,10,11);
input s_274,s_275;//RE__ALLOW(00,01,10,11);
input s_276,s_277;//RE__ALLOW(00,01,10,11);
input s_278,s_279;//RE__ALLOW(00,01,10,11);
input s_280,s_281;//RE__ALLOW(00,01,10,11);
input s_282,s_283;//RE__ALLOW(00,01,10,11);
input s_284,s_285;//RE__ALLOW(00,01,10,11);
input s_286,s_287;//RE__ALLOW(00,01,10,11);
input s_288,s_289;//RE__ALLOW(00,01,10,11);
input s_290,s_291;//RE__ALLOW(00,01,10,11);
input s_292,s_293;//RE__ALLOW(00,01,10,11);
input s_294,s_295;//RE__ALLOW(00,01,10,11);
input s_296,s_297;//RE__ALLOW(00,01,10,11);
input s_298,s_299;//RE__ALLOW(00,01,10,11);
input s_300,s_301;//RE__ALLOW(00,01,10,11);
input s_302,s_303;//RE__ALLOW(00,01,10,11);
input s_304,s_305;//RE__ALLOW(00,01,10,11);
input s_306,s_307;//RE__ALLOW(00,01,10,11);
input s_308,s_309;//RE__ALLOW(00,01,10,11);
input s_310,s_311;//RE__ALLOW(00,01,10,11);
input s_312,s_313;//RE__ALLOW(00,01,10,11);
input s_314,s_315;//RE__ALLOW(00,01,10,11);
input s_316,s_317;//RE__ALLOW(00,01,10,11);
input s_318,s_319;//RE__ALLOW(00,01,10,11);
input s_320,s_321;//RE__ALLOW(00,01,10,11);
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;

  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate19inter0, gate19inter1, gate19inter2, gate19inter3, gate19inter4, gate19inter5, gate19inter6, gate19inter7, gate19inter8, gate19inter9, gate19inter10, gate19inter11, gate19inter12, gate216inter0, gate216inter1, gate216inter2, gate216inter3, gate216inter4, gate216inter5, gate216inter6, gate216inter7, gate216inter8, gate216inter9, gate216inter10, gate216inter11, gate216inter12, gate74inter0, gate74inter1, gate74inter2, gate74inter3, gate74inter4, gate74inter5, gate74inter6, gate74inter7, gate74inter8, gate74inter9, gate74inter10, gate74inter11, gate74inter12, gate35inter0, gate35inter1, gate35inter2, gate35inter3, gate35inter4, gate35inter5, gate35inter6, gate35inter7, gate35inter8, gate35inter9, gate35inter10, gate35inter11, gate35inter12, gate399inter0, gate399inter1, gate399inter2, gate399inter3, gate399inter4, gate399inter5, gate399inter6, gate399inter7, gate399inter8, gate399inter9, gate399inter10, gate399inter11, gate399inter12, gate124inter0, gate124inter1, gate124inter2, gate124inter3, gate124inter4, gate124inter5, gate124inter6, gate124inter7, gate124inter8, gate124inter9, gate124inter10, gate124inter11, gate124inter12, gate496inter0, gate496inter1, gate496inter2, gate496inter3, gate496inter4, gate496inter5, gate496inter6, gate496inter7, gate496inter8, gate496inter9, gate496inter10, gate496inter11, gate496inter12, gate274inter0, gate274inter1, gate274inter2, gate274inter3, gate274inter4, gate274inter5, gate274inter6, gate274inter7, gate274inter8, gate274inter9, gate274inter10, gate274inter11, gate274inter12, gate471inter0, gate471inter1, gate471inter2, gate471inter3, gate471inter4, gate471inter5, gate471inter6, gate471inter7, gate471inter8, gate471inter9, gate471inter10, gate471inter11, gate471inter12, gate497inter0, gate497inter1, gate497inter2, gate497inter3, gate497inter4, gate497inter5, gate497inter6, gate497inter7, gate497inter8, gate497inter9, gate497inter10, gate497inter11, gate497inter12, gate195inter0, gate195inter1, gate195inter2, gate195inter3, gate195inter4, gate195inter5, gate195inter6, gate195inter7, gate195inter8, gate195inter9, gate195inter10, gate195inter11, gate195inter12, gate256inter0, gate256inter1, gate256inter2, gate256inter3, gate256inter4, gate256inter5, gate256inter6, gate256inter7, gate256inter8, gate256inter9, gate256inter10, gate256inter11, gate256inter12, gate101inter0, gate101inter1, gate101inter2, gate101inter3, gate101inter4, gate101inter5, gate101inter6, gate101inter7, gate101inter8, gate101inter9, gate101inter10, gate101inter11, gate101inter12, gate198inter0, gate198inter1, gate198inter2, gate198inter3, gate198inter4, gate198inter5, gate198inter6, gate198inter7, gate198inter8, gate198inter9, gate198inter10, gate198inter11, gate198inter12, gate231inter0, gate231inter1, gate231inter2, gate231inter3, gate231inter4, gate231inter5, gate231inter6, gate231inter7, gate231inter8, gate231inter9, gate231inter10, gate231inter11, gate231inter12, gate272inter0, gate272inter1, gate272inter2, gate272inter3, gate272inter4, gate272inter5, gate272inter6, gate272inter7, gate272inter8, gate272inter9, gate272inter10, gate272inter11, gate272inter12, gate47inter0, gate47inter1, gate47inter2, gate47inter3, gate47inter4, gate47inter5, gate47inter6, gate47inter7, gate47inter8, gate47inter9, gate47inter10, gate47inter11, gate47inter12, gate423inter0, gate423inter1, gate423inter2, gate423inter3, gate423inter4, gate423inter5, gate423inter6, gate423inter7, gate423inter8, gate423inter9, gate423inter10, gate423inter11, gate423inter12, gate71inter0, gate71inter1, gate71inter2, gate71inter3, gate71inter4, gate71inter5, gate71inter6, gate71inter7, gate71inter8, gate71inter9, gate71inter10, gate71inter11, gate71inter12, gate16inter0, gate16inter1, gate16inter2, gate16inter3, gate16inter4, gate16inter5, gate16inter6, gate16inter7, gate16inter8, gate16inter9, gate16inter10, gate16inter11, gate16inter12, gate174inter0, gate174inter1, gate174inter2, gate174inter3, gate174inter4, gate174inter5, gate174inter6, gate174inter7, gate174inter8, gate174inter9, gate174inter10, gate174inter11, gate174inter12, gate139inter0, gate139inter1, gate139inter2, gate139inter3, gate139inter4, gate139inter5, gate139inter6, gate139inter7, gate139inter8, gate139inter9, gate139inter10, gate139inter11, gate139inter12, gate454inter0, gate454inter1, gate454inter2, gate454inter3, gate454inter4, gate454inter5, gate454inter6, gate454inter7, gate454inter8, gate454inter9, gate454inter10, gate454inter11, gate454inter12, gate514inter0, gate514inter1, gate514inter2, gate514inter3, gate514inter4, gate514inter5, gate514inter6, gate514inter7, gate514inter8, gate514inter9, gate514inter10, gate514inter11, gate514inter12, gate128inter0, gate128inter1, gate128inter2, gate128inter3, gate128inter4, gate128inter5, gate128inter6, gate128inter7, gate128inter8, gate128inter9, gate128inter10, gate128inter11, gate128inter12, gate212inter0, gate212inter1, gate212inter2, gate212inter3, gate212inter4, gate212inter5, gate212inter6, gate212inter7, gate212inter8, gate212inter9, gate212inter10, gate212inter11, gate212inter12, gate455inter0, gate455inter1, gate455inter2, gate455inter3, gate455inter4, gate455inter5, gate455inter6, gate455inter7, gate455inter8, gate455inter9, gate455inter10, gate455inter11, gate455inter12, gate49inter0, gate49inter1, gate49inter2, gate49inter3, gate49inter4, gate49inter5, gate49inter6, gate49inter7, gate49inter8, gate49inter9, gate49inter10, gate49inter11, gate49inter12, gate193inter0, gate193inter1, gate193inter2, gate193inter3, gate193inter4, gate193inter5, gate193inter6, gate193inter7, gate193inter8, gate193inter9, gate193inter10, gate193inter11, gate193inter12, gate482inter0, gate482inter1, gate482inter2, gate482inter3, gate482inter4, gate482inter5, gate482inter6, gate482inter7, gate482inter8, gate482inter9, gate482inter10, gate482inter11, gate482inter12, gate20inter0, gate20inter1, gate20inter2, gate20inter3, gate20inter4, gate20inter5, gate20inter6, gate20inter7, gate20inter8, gate20inter9, gate20inter10, gate20inter11, gate20inter12, gate83inter0, gate83inter1, gate83inter2, gate83inter3, gate83inter4, gate83inter5, gate83inter6, gate83inter7, gate83inter8, gate83inter9, gate83inter10, gate83inter11, gate83inter12, gate110inter0, gate110inter1, gate110inter2, gate110inter3, gate110inter4, gate110inter5, gate110inter6, gate110inter7, gate110inter8, gate110inter9, gate110inter10, gate110inter11, gate110inter12, gate64inter0, gate64inter1, gate64inter2, gate64inter3, gate64inter4, gate64inter5, gate64inter6, gate64inter7, gate64inter8, gate64inter9, gate64inter10, gate64inter11, gate64inter12, gate389inter0, gate389inter1, gate389inter2, gate389inter3, gate389inter4, gate389inter5, gate389inter6, gate389inter7, gate389inter8, gate389inter9, gate389inter10, gate389inter11, gate389inter12, gate257inter0, gate257inter1, gate257inter2, gate257inter3, gate257inter4, gate257inter5, gate257inter6, gate257inter7, gate257inter8, gate257inter9, gate257inter10, gate257inter11, gate257inter12, gate136inter0, gate136inter1, gate136inter2, gate136inter3, gate136inter4, gate136inter5, gate136inter6, gate136inter7, gate136inter8, gate136inter9, gate136inter10, gate136inter11, gate136inter12, gate485inter0, gate485inter1, gate485inter2, gate485inter3, gate485inter4, gate485inter5, gate485inter6, gate485inter7, gate485inter8, gate485inter9, gate485inter10, gate485inter11, gate485inter12, gate73inter0, gate73inter1, gate73inter2, gate73inter3, gate73inter4, gate73inter5, gate73inter6, gate73inter7, gate73inter8, gate73inter9, gate73inter10, gate73inter11, gate73inter12, gate293inter0, gate293inter1, gate293inter2, gate293inter3, gate293inter4, gate293inter5, gate293inter6, gate293inter7, gate293inter8, gate293inter9, gate293inter10, gate293inter11, gate293inter12, gate211inter0, gate211inter1, gate211inter2, gate211inter3, gate211inter4, gate211inter5, gate211inter6, gate211inter7, gate211inter8, gate211inter9, gate211inter10, gate211inter11, gate211inter12, gate145inter0, gate145inter1, gate145inter2, gate145inter3, gate145inter4, gate145inter5, gate145inter6, gate145inter7, gate145inter8, gate145inter9, gate145inter10, gate145inter11, gate145inter12, gate236inter0, gate236inter1, gate236inter2, gate236inter3, gate236inter4, gate236inter5, gate236inter6, gate236inter7, gate236inter8, gate236inter9, gate236inter10, gate236inter11, gate236inter12, gate26inter0, gate26inter1, gate26inter2, gate26inter3, gate26inter4, gate26inter5, gate26inter6, gate26inter7, gate26inter8, gate26inter9, gate26inter10, gate26inter11, gate26inter12, gate480inter0, gate480inter1, gate480inter2, gate480inter3, gate480inter4, gate480inter5, gate480inter6, gate480inter7, gate480inter8, gate480inter9, gate480inter10, gate480inter11, gate480inter12, gate222inter0, gate222inter1, gate222inter2, gate222inter3, gate222inter4, gate222inter5, gate222inter6, gate222inter7, gate222inter8, gate222inter9, gate222inter10, gate222inter11, gate222inter12, gate196inter0, gate196inter1, gate196inter2, gate196inter3, gate196inter4, gate196inter5, gate196inter6, gate196inter7, gate196inter8, gate196inter9, gate196inter10, gate196inter11, gate196inter12, gate152inter0, gate152inter1, gate152inter2, gate152inter3, gate152inter4, gate152inter5, gate152inter6, gate152inter7, gate152inter8, gate152inter9, gate152inter10, gate152inter11, gate152inter12, gate457inter0, gate457inter1, gate457inter2, gate457inter3, gate457inter4, gate457inter5, gate457inter6, gate457inter7, gate457inter8, gate457inter9, gate457inter10, gate457inter11, gate457inter12, gate226inter0, gate226inter1, gate226inter2, gate226inter3, gate226inter4, gate226inter5, gate226inter6, gate226inter7, gate226inter8, gate226inter9, gate226inter10, gate226inter11, gate226inter12, gate170inter0, gate170inter1, gate170inter2, gate170inter3, gate170inter4, gate170inter5, gate170inter6, gate170inter7, gate170inter8, gate170inter9, gate170inter10, gate170inter11, gate170inter12, gate171inter0, gate171inter1, gate171inter2, gate171inter3, gate171inter4, gate171inter5, gate171inter6, gate171inter7, gate171inter8, gate171inter9, gate171inter10, gate171inter11, gate171inter12, gate17inter0, gate17inter1, gate17inter2, gate17inter3, gate17inter4, gate17inter5, gate17inter6, gate17inter7, gate17inter8, gate17inter9, gate17inter10, gate17inter11, gate17inter12, gate48inter0, gate48inter1, gate48inter2, gate48inter3, gate48inter4, gate48inter5, gate48inter6, gate48inter7, gate48inter8, gate48inter9, gate48inter10, gate48inter11, gate48inter12, gate443inter0, gate443inter1, gate443inter2, gate443inter3, gate443inter4, gate443inter5, gate443inter6, gate443inter7, gate443inter8, gate443inter9, gate443inter10, gate443inter11, gate443inter12, gate205inter0, gate205inter1, gate205inter2, gate205inter3, gate205inter4, gate205inter5, gate205inter6, gate205inter7, gate205inter8, gate205inter9, gate205inter10, gate205inter11, gate205inter12, gate255inter0, gate255inter1, gate255inter2, gate255inter3, gate255inter4, gate255inter5, gate255inter6, gate255inter7, gate255inter8, gate255inter9, gate255inter10, gate255inter11, gate255inter12, gate467inter0, gate467inter1, gate467inter2, gate467inter3, gate467inter4, gate467inter5, gate467inter6, gate467inter7, gate467inter8, gate467inter9, gate467inter10, gate467inter11, gate467inter12, gate194inter0, gate194inter1, gate194inter2, gate194inter3, gate194inter4, gate194inter5, gate194inter6, gate194inter7, gate194inter8, gate194inter9, gate194inter10, gate194inter11, gate194inter12, gate510inter0, gate510inter1, gate510inter2, gate510inter3, gate510inter4, gate510inter5, gate510inter6, gate510inter7, gate510inter8, gate510inter9, gate510inter10, gate510inter11, gate510inter12, gate232inter0, gate232inter1, gate232inter2, gate232inter3, gate232inter4, gate232inter5, gate232inter6, gate232inter7, gate232inter8, gate232inter9, gate232inter10, gate232inter11, gate232inter12, gate148inter0, gate148inter1, gate148inter2, gate148inter3, gate148inter4, gate148inter5, gate148inter6, gate148inter7, gate148inter8, gate148inter9, gate148inter10, gate148inter11, gate148inter12, gate104inter0, gate104inter1, gate104inter2, gate104inter3, gate104inter4, gate104inter5, gate104inter6, gate104inter7, gate104inter8, gate104inter9, gate104inter10, gate104inter11, gate104inter12, gate153inter0, gate153inter1, gate153inter2, gate153inter3, gate153inter4, gate153inter5, gate153inter6, gate153inter7, gate153inter8, gate153inter9, gate153inter10, gate153inter11, gate153inter12, gate448inter0, gate448inter1, gate448inter2, gate448inter3, gate448inter4, gate448inter5, gate448inter6, gate448inter7, gate448inter8, gate448inter9, gate448inter10, gate448inter11, gate448inter12, gate131inter0, gate131inter1, gate131inter2, gate131inter3, gate131inter4, gate131inter5, gate131inter6, gate131inter7, gate131inter8, gate131inter9, gate131inter10, gate131inter11, gate131inter12, gate204inter0, gate204inter1, gate204inter2, gate204inter3, gate204inter4, gate204inter5, gate204inter6, gate204inter7, gate204inter8, gate204inter9, gate204inter10, gate204inter11, gate204inter12, gate281inter0, gate281inter1, gate281inter2, gate281inter3, gate281inter4, gate281inter5, gate281inter6, gate281inter7, gate281inter8, gate281inter9, gate281inter10, gate281inter11, gate281inter12, gate119inter0, gate119inter1, gate119inter2, gate119inter3, gate119inter4, gate119inter5, gate119inter6, gate119inter7, gate119inter8, gate119inter9, gate119inter10, gate119inter11, gate119inter12, gate266inter0, gate266inter1, gate266inter2, gate266inter3, gate266inter4, gate266inter5, gate266inter6, gate266inter7, gate266inter8, gate266inter9, gate266inter10, gate266inter11, gate266inter12, gate436inter0, gate436inter1, gate436inter2, gate436inter3, gate436inter4, gate436inter5, gate436inter6, gate436inter7, gate436inter8, gate436inter9, gate436inter10, gate436inter11, gate436inter12, gate403inter0, gate403inter1, gate403inter2, gate403inter3, gate403inter4, gate403inter5, gate403inter6, gate403inter7, gate403inter8, gate403inter9, gate403inter10, gate403inter11, gate403inter12, gate494inter0, gate494inter1, gate494inter2, gate494inter3, gate494inter4, gate494inter5, gate494inter6, gate494inter7, gate494inter8, gate494inter9, gate494inter10, gate494inter11, gate494inter12, gate161inter0, gate161inter1, gate161inter2, gate161inter3, gate161inter4, gate161inter5, gate161inter6, gate161inter7, gate161inter8, gate161inter9, gate161inter10, gate161inter11, gate161inter12, gate506inter0, gate506inter1, gate506inter2, gate506inter3, gate506inter4, gate506inter5, gate506inter6, gate506inter7, gate506inter8, gate506inter9, gate506inter10, gate506inter11, gate506inter12, gate238inter0, gate238inter1, gate238inter2, gate238inter3, gate238inter4, gate238inter5, gate238inter6, gate238inter7, gate238inter8, gate238inter9, gate238inter10, gate238inter11, gate238inter12, gate229inter0, gate229inter1, gate229inter2, gate229inter3, gate229inter4, gate229inter5, gate229inter6, gate229inter7, gate229inter8, gate229inter9, gate229inter10, gate229inter11, gate229inter12, gate203inter0, gate203inter1, gate203inter2, gate203inter3, gate203inter4, gate203inter5, gate203inter6, gate203inter7, gate203inter8, gate203inter9, gate203inter10, gate203inter11, gate203inter12, gate115inter0, gate115inter1, gate115inter2, gate115inter3, gate115inter4, gate115inter5, gate115inter6, gate115inter7, gate115inter8, gate115inter9, gate115inter10, gate115inter11, gate115inter12, gate450inter0, gate450inter1, gate450inter2, gate450inter3, gate450inter4, gate450inter5, gate450inter6, gate450inter7, gate450inter8, gate450inter9, gate450inter10, gate450inter11, gate450inter12, gate237inter0, gate237inter1, gate237inter2, gate237inter3, gate237inter4, gate237inter5, gate237inter6, gate237inter7, gate237inter8, gate237inter9, gate237inter10, gate237inter11, gate237inter12, gate451inter0, gate451inter1, gate451inter2, gate451inter3, gate451inter4, gate451inter5, gate451inter6, gate451inter7, gate451inter8, gate451inter9, gate451inter10, gate451inter11, gate451inter12, gate10inter0, gate10inter1, gate10inter2, gate10inter3, gate10inter4, gate10inter5, gate10inter6, gate10inter7, gate10inter8, gate10inter9, gate10inter10, gate10inter11, gate10inter12, gate483inter0, gate483inter1, gate483inter2, gate483inter3, gate483inter4, gate483inter5, gate483inter6, gate483inter7, gate483inter8, gate483inter9, gate483inter10, gate483inter11, gate483inter12, gate286inter0, gate286inter1, gate286inter2, gate286inter3, gate286inter4, gate286inter5, gate286inter6, gate286inter7, gate286inter8, gate286inter9, gate286inter10, gate286inter11, gate286inter12, gate164inter0, gate164inter1, gate164inter2, gate164inter3, gate164inter4, gate164inter5, gate164inter6, gate164inter7, gate164inter8, gate164inter9, gate164inter10, gate164inter11, gate164inter12, gate411inter0, gate411inter1, gate411inter2, gate411inter3, gate411inter4, gate411inter5, gate411inter6, gate411inter7, gate411inter8, gate411inter9, gate411inter10, gate411inter11, gate411inter12, gate245inter0, gate245inter1, gate245inter2, gate245inter3, gate245inter4, gate245inter5, gate245inter6, gate245inter7, gate245inter8, gate245inter9, gate245inter10, gate245inter11, gate245inter12, gate405inter0, gate405inter1, gate405inter2, gate405inter3, gate405inter4, gate405inter5, gate405inter6, gate405inter7, gate405inter8, gate405inter9, gate405inter10, gate405inter11, gate405inter12, gate260inter0, gate260inter1, gate260inter2, gate260inter3, gate260inter4, gate260inter5, gate260inter6, gate260inter7, gate260inter8, gate260inter9, gate260inter10, gate260inter11, gate260inter12, gate57inter0, gate57inter1, gate57inter2, gate57inter3, gate57inter4, gate57inter5, gate57inter6, gate57inter7, gate57inter8, gate57inter9, gate57inter10, gate57inter11, gate57inter12, gate184inter0, gate184inter1, gate184inter2, gate184inter3, gate184inter4, gate184inter5, gate184inter6, gate184inter7, gate184inter8, gate184inter9, gate184inter10, gate184inter11, gate184inter12, gate501inter0, gate501inter1, gate501inter2, gate501inter3, gate501inter4, gate501inter5, gate501inter6, gate501inter7, gate501inter8, gate501inter9, gate501inter10, gate501inter11, gate501inter12, gate140inter0, gate140inter1, gate140inter2, gate140inter3, gate140inter4, gate140inter5, gate140inter6, gate140inter7, gate140inter8, gate140inter9, gate140inter10, gate140inter11, gate140inter12, gate42inter0, gate42inter1, gate42inter2, gate42inter3, gate42inter4, gate42inter5, gate42inter6, gate42inter7, gate42inter8, gate42inter9, gate42inter10, gate42inter11, gate42inter12, gate191inter0, gate191inter1, gate191inter2, gate191inter3, gate191inter4, gate191inter5, gate191inter6, gate191inter7, gate191inter8, gate191inter9, gate191inter10, gate191inter11, gate191inter12, gate122inter0, gate122inter1, gate122inter2, gate122inter3, gate122inter4, gate122inter5, gate122inter6, gate122inter7, gate122inter8, gate122inter9, gate122inter10, gate122inter11, gate122inter12, gate417inter0, gate417inter1, gate417inter2, gate417inter3, gate417inter4, gate417inter5, gate417inter6, gate417inter7, gate417inter8, gate417inter9, gate417inter10, gate417inter11, gate417inter12, gate440inter0, gate440inter1, gate440inter2, gate440inter3, gate440inter4, gate440inter5, gate440inter6, gate440inter7, gate440inter8, gate440inter9, gate440inter10, gate440inter11, gate440inter12, gate460inter0, gate460inter1, gate460inter2, gate460inter3, gate460inter4, gate460inter5, gate460inter6, gate460inter7, gate460inter8, gate460inter9, gate460inter10, gate460inter11, gate460inter12, gate113inter0, gate113inter1, gate113inter2, gate113inter3, gate113inter4, gate113inter5, gate113inter6, gate113inter7, gate113inter8, gate113inter9, gate113inter10, gate113inter11, gate113inter12, gate414inter0, gate414inter1, gate414inter2, gate414inter3, gate414inter4, gate414inter5, gate414inter6, gate414inter7, gate414inter8, gate414inter9, gate414inter10, gate414inter11, gate414inter12, gate291inter0, gate291inter1, gate291inter2, gate291inter3, gate291inter4, gate291inter5, gate291inter6, gate291inter7, gate291inter8, gate291inter9, gate291inter10, gate291inter11, gate291inter12, gate12inter0, gate12inter1, gate12inter2, gate12inter3, gate12inter4, gate12inter5, gate12inter6, gate12inter7, gate12inter8, gate12inter9, gate12inter10, gate12inter11, gate12inter12, gate265inter0, gate265inter1, gate265inter2, gate265inter3, gate265inter4, gate265inter5, gate265inter6, gate265inter7, gate265inter8, gate265inter9, gate265inter10, gate265inter11, gate265inter12, gate188inter0, gate188inter1, gate188inter2, gate188inter3, gate188inter4, gate188inter5, gate188inter6, gate188inter7, gate188inter8, gate188inter9, gate188inter10, gate188inter11, gate188inter12, gate96inter0, gate96inter1, gate96inter2, gate96inter3, gate96inter4, gate96inter5, gate96inter6, gate96inter7, gate96inter8, gate96inter9, gate96inter10, gate96inter11, gate96inter12, gate408inter0, gate408inter1, gate408inter2, gate408inter3, gate408inter4, gate408inter5, gate408inter6, gate408inter7, gate408inter8, gate408inter9, gate408inter10, gate408inter11, gate408inter12, gate166inter0, gate166inter1, gate166inter2, gate166inter3, gate166inter4, gate166inter5, gate166inter6, gate166inter7, gate166inter8, gate166inter9, gate166inter10, gate166inter11, gate166inter12, gate219inter0, gate219inter1, gate219inter2, gate219inter3, gate219inter4, gate219inter5, gate219inter6, gate219inter7, gate219inter8, gate219inter9, gate219inter10, gate219inter11, gate219inter12, gate218inter0, gate218inter1, gate218inter2, gate218inter3, gate218inter4, gate218inter5, gate218inter6, gate218inter7, gate218inter8, gate218inter9, gate218inter10, gate218inter11, gate218inter12, gate91inter0, gate91inter1, gate91inter2, gate91inter3, gate91inter4, gate91inter5, gate91inter6, gate91inter7, gate91inter8, gate91inter9, gate91inter10, gate91inter11, gate91inter12, gate412inter0, gate412inter1, gate412inter2, gate412inter3, gate412inter4, gate412inter5, gate412inter6, gate412inter7, gate412inter8, gate412inter9, gate412inter10, gate412inter11, gate412inter12, gate275inter0, gate275inter1, gate275inter2, gate275inter3, gate275inter4, gate275inter5, gate275inter6, gate275inter7, gate275inter8, gate275inter9, gate275inter10, gate275inter11, gate275inter12, gate100inter0, gate100inter1, gate100inter2, gate100inter3, gate100inter4, gate100inter5, gate100inter6, gate100inter7, gate100inter8, gate100inter9, gate100inter10, gate100inter11, gate100inter12, gate199inter0, gate199inter1, gate199inter2, gate199inter3, gate199inter4, gate199inter5, gate199inter6, gate199inter7, gate199inter8, gate199inter9, gate199inter10, gate199inter11, gate199inter12, gate89inter0, gate89inter1, gate89inter2, gate89inter3, gate89inter4, gate89inter5, gate89inter6, gate89inter7, gate89inter8, gate89inter9, gate89inter10, gate89inter11, gate89inter12, gate430inter0, gate430inter1, gate430inter2, gate430inter3, gate430inter4, gate430inter5, gate430inter6, gate430inter7, gate430inter8, gate430inter9, gate430inter10, gate430inter11, gate430inter12, gate263inter0, gate263inter1, gate263inter2, gate263inter3, gate263inter4, gate263inter5, gate263inter6, gate263inter7, gate263inter8, gate263inter9, gate263inter10, gate263inter11, gate263inter12, gate428inter0, gate428inter1, gate428inter2, gate428inter3, gate428inter4, gate428inter5, gate428inter6, gate428inter7, gate428inter8, gate428inter9, gate428inter10, gate428inter11, gate428inter12, gate154inter0, gate154inter1, gate154inter2, gate154inter3, gate154inter4, gate154inter5, gate154inter6, gate154inter7, gate154inter8, gate154inter9, gate154inter10, gate154inter11, gate154inter12, gate246inter0, gate246inter1, gate246inter2, gate246inter3, gate246inter4, gate246inter5, gate246inter6, gate246inter7, gate246inter8, gate246inter9, gate246inter10, gate246inter11, gate246inter12, gate24inter0, gate24inter1, gate24inter2, gate24inter3, gate24inter4, gate24inter5, gate24inter6, gate24inter7, gate24inter8, gate24inter9, gate24inter10, gate24inter11, gate24inter12, gate418inter0, gate418inter1, gate418inter2, gate418inter3, gate418inter4, gate418inter5, gate418inter6, gate418inter7, gate418inter8, gate418inter9, gate418inter10, gate418inter11, gate418inter12, gate81inter0, gate81inter1, gate81inter2, gate81inter3, gate81inter4, gate81inter5, gate81inter6, gate81inter7, gate81inter8, gate81inter9, gate81inter10, gate81inter11, gate81inter12, gate468inter0, gate468inter1, gate468inter2, gate468inter3, gate468inter4, gate468inter5, gate468inter6, gate468inter7, gate468inter8, gate468inter9, gate468inter10, gate468inter11, gate468inter12, gate464inter0, gate464inter1, gate464inter2, gate464inter3, gate464inter4, gate464inter5, gate464inter6, gate464inter7, gate464inter8, gate464inter9, gate464inter10, gate464inter11, gate464inter12, gate395inter0, gate395inter1, gate395inter2, gate395inter3, gate395inter4, gate395inter5, gate395inter6, gate395inter7, gate395inter8, gate395inter9, gate395inter10, gate395inter11, gate395inter12, gate44inter0, gate44inter1, gate44inter2, gate44inter3, gate44inter4, gate44inter5, gate44inter6, gate44inter7, gate44inter8, gate44inter9, gate44inter10, gate44inter11, gate44inter12, gate419inter0, gate419inter1, gate419inter2, gate419inter3, gate419inter4, gate419inter5, gate419inter6, gate419inter7, gate419inter8, gate419inter9, gate419inter10, gate419inter11, gate419inter12, gate69inter0, gate69inter1, gate69inter2, gate69inter3, gate69inter4, gate69inter5, gate69inter6, gate69inter7, gate69inter8, gate69inter9, gate69inter10, gate69inter11, gate69inter12, gate43inter0, gate43inter1, gate43inter2, gate43inter3, gate43inter4, gate43inter5, gate43inter6, gate43inter7, gate43inter8, gate43inter9, gate43inter10, gate43inter11, gate43inter12, gate155inter0, gate155inter1, gate155inter2, gate155inter3, gate155inter4, gate155inter5, gate155inter6, gate155inter7, gate155inter8, gate155inter9, gate155inter10, gate155inter11, gate155inter12, gate137inter0, gate137inter1, gate137inter2, gate137inter3, gate137inter4, gate137inter5, gate137inter6, gate137inter7, gate137inter8, gate137inter9, gate137inter10, gate137inter11, gate137inter12, gate144inter0, gate144inter1, gate144inter2, gate144inter3, gate144inter4, gate144inter5, gate144inter6, gate144inter7, gate144inter8, gate144inter9, gate144inter10, gate144inter11, gate144inter12, gate227inter0, gate227inter1, gate227inter2, gate227inter3, gate227inter4, gate227inter5, gate227inter6, gate227inter7, gate227inter8, gate227inter9, gate227inter10, gate227inter11, gate227inter12, gate79inter0, gate79inter1, gate79inter2, gate79inter3, gate79inter4, gate79inter5, gate79inter6, gate79inter7, gate79inter8, gate79inter9, gate79inter10, gate79inter11, gate79inter12, gate151inter0, gate151inter1, gate151inter2, gate151inter3, gate151inter4, gate151inter5, gate151inter6, gate151inter7, gate151inter8, gate151inter9, gate151inter10, gate151inter11, gate151inter12, gate36inter0, gate36inter1, gate36inter2, gate36inter3, gate36inter4, gate36inter5, gate36inter6, gate36inter7, gate36inter8, gate36inter9, gate36inter10, gate36inter11, gate36inter12, gate129inter0, gate129inter1, gate129inter2, gate129inter3, gate129inter4, gate129inter5, gate129inter6, gate129inter7, gate129inter8, gate129inter9, gate129inter10, gate129inter11, gate129inter12, gate207inter0, gate207inter1, gate207inter2, gate207inter3, gate207inter4, gate207inter5, gate207inter6, gate207inter7, gate207inter8, gate207inter9, gate207inter10, gate207inter11, gate207inter12, gate268inter0, gate268inter1, gate268inter2, gate268inter3, gate268inter4, gate268inter5, gate268inter6, gate268inter7, gate268inter8, gate268inter9, gate268inter10, gate268inter11, gate268inter12, gate250inter0, gate250inter1, gate250inter2, gate250inter3, gate250inter4, gate250inter5, gate250inter6, gate250inter7, gate250inter8, gate250inter9, gate250inter10, gate250inter11, gate250inter12, gate470inter0, gate470inter1, gate470inter2, gate470inter3, gate470inter4, gate470inter5, gate470inter6, gate470inter7, gate470inter8, gate470inter9, gate470inter10, gate470inter11, gate470inter12, gate27inter0, gate27inter1, gate27inter2, gate27inter3, gate27inter4, gate27inter5, gate27inter6, gate27inter7, gate27inter8, gate27inter9, gate27inter10, gate27inter11, gate27inter12, gate130inter0, gate130inter1, gate130inter2, gate130inter3, gate130inter4, gate130inter5, gate130inter6, gate130inter7, gate130inter8, gate130inter9, gate130inter10, gate130inter11, gate130inter12, gate240inter0, gate240inter1, gate240inter2, gate240inter3, gate240inter4, gate240inter5, gate240inter6, gate240inter7, gate240inter8, gate240inter9, gate240inter10, gate240inter11, gate240inter12, gate25inter0, gate25inter1, gate25inter2, gate25inter3, gate25inter4, gate25inter5, gate25inter6, gate25inter7, gate25inter8, gate25inter9, gate25inter10, gate25inter11, gate25inter12, gate490inter0, gate490inter1, gate490inter2, gate490inter3, gate490inter4, gate490inter5, gate490inter6, gate490inter7, gate490inter8, gate490inter9, gate490inter10, gate490inter11, gate490inter12, gate267inter0, gate267inter1, gate267inter2, gate267inter3, gate267inter4, gate267inter5, gate267inter6, gate267inter7, gate267inter8, gate267inter9, gate267inter10, gate267inter11, gate267inter12, gate135inter0, gate135inter1, gate135inter2, gate135inter3, gate135inter4, gate135inter5, gate135inter6, gate135inter7, gate135inter8, gate135inter9, gate135inter10, gate135inter11, gate135inter12, gate437inter0, gate437inter1, gate437inter2, gate437inter3, gate437inter4, gate437inter5, gate437inter6, gate437inter7, gate437inter8, gate437inter9, gate437inter10, gate437inter11, gate437inter12, gate202inter0, gate202inter1, gate202inter2, gate202inter3, gate202inter4, gate202inter5, gate202inter6, gate202inter7, gate202inter8, gate202inter9, gate202inter10, gate202inter11, gate202inter12, gate499inter0, gate499inter1, gate499inter2, gate499inter3, gate499inter4, gate499inter5, gate499inter6, gate499inter7, gate499inter8, gate499inter9, gate499inter10, gate499inter11, gate499inter12, gate103inter0, gate103inter1, gate103inter2, gate103inter3, gate103inter4, gate103inter5, gate103inter6, gate103inter7, gate103inter8, gate103inter9, gate103inter10, gate103inter11, gate103inter12, gate221inter0, gate221inter1, gate221inter2, gate221inter3, gate221inter4, gate221inter5, gate221inter6, gate221inter7, gate221inter8, gate221inter9, gate221inter10, gate221inter11, gate221inter12, gate427inter0, gate427inter1, gate427inter2, gate427inter3, gate427inter4, gate427inter5, gate427inter6, gate427inter7, gate427inter8, gate427inter9, gate427inter10, gate427inter11, gate427inter12, gate492inter0, gate492inter1, gate492inter2, gate492inter3, gate492inter4, gate492inter5, gate492inter6, gate492inter7, gate492inter8, gate492inter9, gate492inter10, gate492inter11, gate492inter12, gate296inter0, gate296inter1, gate296inter2, gate296inter3, gate296inter4, gate296inter5, gate296inter6, gate296inter7, gate296inter8, gate296inter9, gate296inter10, gate296inter11, gate296inter12, gate175inter0, gate175inter1, gate175inter2, gate175inter3, gate175inter4, gate175inter5, gate175inter6, gate175inter7, gate175inter8, gate175inter9, gate175inter10, gate175inter11, gate175inter12, gate230inter0, gate230inter1, gate230inter2, gate230inter3, gate230inter4, gate230inter5, gate230inter6, gate230inter7, gate230inter8, gate230inter9, gate230inter10, gate230inter11, gate230inter12;



and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );
nand2 gate9( .a(G1), .b(G2), .O(G266) );

  xor2  gate1695(.a(G4), .b(G3), .O(gate10inter0));
  nand2 gate1696(.a(gate10inter0), .b(s_164), .O(gate10inter1));
  and2  gate1697(.a(G4), .b(G3), .O(gate10inter2));
  inv1  gate1698(.a(s_164), .O(gate10inter3));
  inv1  gate1699(.a(s_165), .O(gate10inter4));
  nand2 gate1700(.a(gate10inter4), .b(gate10inter3), .O(gate10inter5));
  nor2  gate1701(.a(gate10inter5), .b(gate10inter2), .O(gate10inter6));
  inv1  gate1702(.a(G3), .O(gate10inter7));
  inv1  gate1703(.a(G4), .O(gate10inter8));
  nand2 gate1704(.a(gate10inter8), .b(gate10inter7), .O(gate10inter9));
  nand2 gate1705(.a(s_165), .b(gate10inter3), .O(gate10inter10));
  nor2  gate1706(.a(gate10inter10), .b(gate10inter9), .O(gate10inter11));
  nor2  gate1707(.a(gate10inter11), .b(gate10inter6), .O(gate10inter12));
  nand2 gate1708(.a(gate10inter12), .b(gate10inter1), .O(G269));
nand2 gate11( .a(G5), .b(G6), .O(G272) );

  xor2  gate1989(.a(G8), .b(G7), .O(gate12inter0));
  nand2 gate1990(.a(gate12inter0), .b(s_206), .O(gate12inter1));
  and2  gate1991(.a(G8), .b(G7), .O(gate12inter2));
  inv1  gate1992(.a(s_206), .O(gate12inter3));
  inv1  gate1993(.a(s_207), .O(gate12inter4));
  nand2 gate1994(.a(gate12inter4), .b(gate12inter3), .O(gate12inter5));
  nor2  gate1995(.a(gate12inter5), .b(gate12inter2), .O(gate12inter6));
  inv1  gate1996(.a(G7), .O(gate12inter7));
  inv1  gate1997(.a(G8), .O(gate12inter8));
  nand2 gate1998(.a(gate12inter8), .b(gate12inter7), .O(gate12inter9));
  nand2 gate1999(.a(s_207), .b(gate12inter3), .O(gate12inter10));
  nor2  gate2000(.a(gate12inter10), .b(gate12inter9), .O(gate12inter11));
  nor2  gate2001(.a(gate12inter11), .b(gate12inter6), .O(gate12inter12));
  nand2 gate2002(.a(gate12inter12), .b(gate12inter1), .O(G275));
nand2 gate13( .a(G9), .b(G10), .O(G278) );
nand2 gate14( .a(G11), .b(G12), .O(G281) );
nand2 gate15( .a(G13), .b(G14), .O(G284) );

  xor2  gate813(.a(G16), .b(G15), .O(gate16inter0));
  nand2 gate814(.a(gate16inter0), .b(s_38), .O(gate16inter1));
  and2  gate815(.a(G16), .b(G15), .O(gate16inter2));
  inv1  gate816(.a(s_38), .O(gate16inter3));
  inv1  gate817(.a(s_39), .O(gate16inter4));
  nand2 gate818(.a(gate16inter4), .b(gate16inter3), .O(gate16inter5));
  nor2  gate819(.a(gate16inter5), .b(gate16inter2), .O(gate16inter6));
  inv1  gate820(.a(G15), .O(gate16inter7));
  inv1  gate821(.a(G16), .O(gate16inter8));
  nand2 gate822(.a(gate16inter8), .b(gate16inter7), .O(gate16inter9));
  nand2 gate823(.a(s_39), .b(gate16inter3), .O(gate16inter10));
  nor2  gate824(.a(gate16inter10), .b(gate16inter9), .O(gate16inter11));
  nor2  gate825(.a(gate16inter11), .b(gate16inter6), .O(gate16inter12));
  nand2 gate826(.a(gate16inter12), .b(gate16inter1), .O(G287));

  xor2  gate1275(.a(G18), .b(G17), .O(gate17inter0));
  nand2 gate1276(.a(gate17inter0), .b(s_104), .O(gate17inter1));
  and2  gate1277(.a(G18), .b(G17), .O(gate17inter2));
  inv1  gate1278(.a(s_104), .O(gate17inter3));
  inv1  gate1279(.a(s_105), .O(gate17inter4));
  nand2 gate1280(.a(gate17inter4), .b(gate17inter3), .O(gate17inter5));
  nor2  gate1281(.a(gate17inter5), .b(gate17inter2), .O(gate17inter6));
  inv1  gate1282(.a(G17), .O(gate17inter7));
  inv1  gate1283(.a(G18), .O(gate17inter8));
  nand2 gate1284(.a(gate17inter8), .b(gate17inter7), .O(gate17inter9));
  nand2 gate1285(.a(s_105), .b(gate17inter3), .O(gate17inter10));
  nor2  gate1286(.a(gate17inter10), .b(gate17inter9), .O(gate17inter11));
  nor2  gate1287(.a(gate17inter11), .b(gate17inter6), .O(gate17inter12));
  nand2 gate1288(.a(gate17inter12), .b(gate17inter1), .O(G290));
nand2 gate18( .a(G19), .b(G20), .O(G293) );

  xor2  gate547(.a(G22), .b(G21), .O(gate19inter0));
  nand2 gate548(.a(gate19inter0), .b(s_0), .O(gate19inter1));
  and2  gate549(.a(G22), .b(G21), .O(gate19inter2));
  inv1  gate550(.a(s_0), .O(gate19inter3));
  inv1  gate551(.a(s_1), .O(gate19inter4));
  nand2 gate552(.a(gate19inter4), .b(gate19inter3), .O(gate19inter5));
  nor2  gate553(.a(gate19inter5), .b(gate19inter2), .O(gate19inter6));
  inv1  gate554(.a(G21), .O(gate19inter7));
  inv1  gate555(.a(G22), .O(gate19inter8));
  nand2 gate556(.a(gate19inter8), .b(gate19inter7), .O(gate19inter9));
  nand2 gate557(.a(s_1), .b(gate19inter3), .O(gate19inter10));
  nor2  gate558(.a(gate19inter10), .b(gate19inter9), .O(gate19inter11));
  nor2  gate559(.a(gate19inter11), .b(gate19inter6), .O(gate19inter12));
  nand2 gate560(.a(gate19inter12), .b(gate19inter1), .O(G296));

  xor2  gate967(.a(G24), .b(G23), .O(gate20inter0));
  nand2 gate968(.a(gate20inter0), .b(s_60), .O(gate20inter1));
  and2  gate969(.a(G24), .b(G23), .O(gate20inter2));
  inv1  gate970(.a(s_60), .O(gate20inter3));
  inv1  gate971(.a(s_61), .O(gate20inter4));
  nand2 gate972(.a(gate20inter4), .b(gate20inter3), .O(gate20inter5));
  nor2  gate973(.a(gate20inter5), .b(gate20inter2), .O(gate20inter6));
  inv1  gate974(.a(G23), .O(gate20inter7));
  inv1  gate975(.a(G24), .O(gate20inter8));
  nand2 gate976(.a(gate20inter8), .b(gate20inter7), .O(gate20inter9));
  nand2 gate977(.a(s_61), .b(gate20inter3), .O(gate20inter10));
  nor2  gate978(.a(gate20inter10), .b(gate20inter9), .O(gate20inter11));
  nor2  gate979(.a(gate20inter11), .b(gate20inter6), .O(gate20inter12));
  nand2 gate980(.a(gate20inter12), .b(gate20inter1), .O(G299));
nand2 gate21( .a(G25), .b(G26), .O(G302) );
nand2 gate22( .a(G27), .b(G28), .O(G305) );
nand2 gate23( .a(G29), .b(G30), .O(G308) );

  xor2  gate2255(.a(G32), .b(G31), .O(gate24inter0));
  nand2 gate2256(.a(gate24inter0), .b(s_244), .O(gate24inter1));
  and2  gate2257(.a(G32), .b(G31), .O(gate24inter2));
  inv1  gate2258(.a(s_244), .O(gate24inter3));
  inv1  gate2259(.a(s_245), .O(gate24inter4));
  nand2 gate2260(.a(gate24inter4), .b(gate24inter3), .O(gate24inter5));
  nor2  gate2261(.a(gate24inter5), .b(gate24inter2), .O(gate24inter6));
  inv1  gate2262(.a(G31), .O(gate24inter7));
  inv1  gate2263(.a(G32), .O(gate24inter8));
  nand2 gate2264(.a(gate24inter8), .b(gate24inter7), .O(gate24inter9));
  nand2 gate2265(.a(s_245), .b(gate24inter3), .O(gate24inter10));
  nor2  gate2266(.a(gate24inter10), .b(gate24inter9), .O(gate24inter11));
  nor2  gate2267(.a(gate24inter11), .b(gate24inter6), .O(gate24inter12));
  nand2 gate2268(.a(gate24inter12), .b(gate24inter1), .O(G311));

  xor2  gate2605(.a(G5), .b(G1), .O(gate25inter0));
  nand2 gate2606(.a(gate25inter0), .b(s_294), .O(gate25inter1));
  and2  gate2607(.a(G5), .b(G1), .O(gate25inter2));
  inv1  gate2608(.a(s_294), .O(gate25inter3));
  inv1  gate2609(.a(s_295), .O(gate25inter4));
  nand2 gate2610(.a(gate25inter4), .b(gate25inter3), .O(gate25inter5));
  nor2  gate2611(.a(gate25inter5), .b(gate25inter2), .O(gate25inter6));
  inv1  gate2612(.a(G1), .O(gate25inter7));
  inv1  gate2613(.a(G5), .O(gate25inter8));
  nand2 gate2614(.a(gate25inter8), .b(gate25inter7), .O(gate25inter9));
  nand2 gate2615(.a(s_295), .b(gate25inter3), .O(gate25inter10));
  nor2  gate2616(.a(gate25inter10), .b(gate25inter9), .O(gate25inter11));
  nor2  gate2617(.a(gate25inter11), .b(gate25inter6), .O(gate25inter12));
  nand2 gate2618(.a(gate25inter12), .b(gate25inter1), .O(G314));

  xor2  gate1149(.a(G13), .b(G9), .O(gate26inter0));
  nand2 gate1150(.a(gate26inter0), .b(s_86), .O(gate26inter1));
  and2  gate1151(.a(G13), .b(G9), .O(gate26inter2));
  inv1  gate1152(.a(s_86), .O(gate26inter3));
  inv1  gate1153(.a(s_87), .O(gate26inter4));
  nand2 gate1154(.a(gate26inter4), .b(gate26inter3), .O(gate26inter5));
  nor2  gate1155(.a(gate26inter5), .b(gate26inter2), .O(gate26inter6));
  inv1  gate1156(.a(G9), .O(gate26inter7));
  inv1  gate1157(.a(G13), .O(gate26inter8));
  nand2 gate1158(.a(gate26inter8), .b(gate26inter7), .O(gate26inter9));
  nand2 gate1159(.a(s_87), .b(gate26inter3), .O(gate26inter10));
  nor2  gate1160(.a(gate26inter10), .b(gate26inter9), .O(gate26inter11));
  nor2  gate1161(.a(gate26inter11), .b(gate26inter6), .O(gate26inter12));
  nand2 gate1162(.a(gate26inter12), .b(gate26inter1), .O(G317));

  xor2  gate2563(.a(G6), .b(G2), .O(gate27inter0));
  nand2 gate2564(.a(gate27inter0), .b(s_288), .O(gate27inter1));
  and2  gate2565(.a(G6), .b(G2), .O(gate27inter2));
  inv1  gate2566(.a(s_288), .O(gate27inter3));
  inv1  gate2567(.a(s_289), .O(gate27inter4));
  nand2 gate2568(.a(gate27inter4), .b(gate27inter3), .O(gate27inter5));
  nor2  gate2569(.a(gate27inter5), .b(gate27inter2), .O(gate27inter6));
  inv1  gate2570(.a(G2), .O(gate27inter7));
  inv1  gate2571(.a(G6), .O(gate27inter8));
  nand2 gate2572(.a(gate27inter8), .b(gate27inter7), .O(gate27inter9));
  nand2 gate2573(.a(s_289), .b(gate27inter3), .O(gate27inter10));
  nor2  gate2574(.a(gate27inter10), .b(gate27inter9), .O(gate27inter11));
  nor2  gate2575(.a(gate27inter11), .b(gate27inter6), .O(gate27inter12));
  nand2 gate2576(.a(gate27inter12), .b(gate27inter1), .O(G320));
nand2 gate28( .a(G10), .b(G14), .O(G323) );
nand2 gate29( .a(G3), .b(G7), .O(G326) );
nand2 gate30( .a(G11), .b(G15), .O(G329) );
nand2 gate31( .a(G4), .b(G8), .O(G332) );
nand2 gate32( .a(G12), .b(G16), .O(G335) );
nand2 gate33( .a(G17), .b(G21), .O(G338) );
nand2 gate34( .a(G25), .b(G29), .O(G341) );

  xor2  gate589(.a(G22), .b(G18), .O(gate35inter0));
  nand2 gate590(.a(gate35inter0), .b(s_6), .O(gate35inter1));
  and2  gate591(.a(G22), .b(G18), .O(gate35inter2));
  inv1  gate592(.a(s_6), .O(gate35inter3));
  inv1  gate593(.a(s_7), .O(gate35inter4));
  nand2 gate594(.a(gate35inter4), .b(gate35inter3), .O(gate35inter5));
  nor2  gate595(.a(gate35inter5), .b(gate35inter2), .O(gate35inter6));
  inv1  gate596(.a(G18), .O(gate35inter7));
  inv1  gate597(.a(G22), .O(gate35inter8));
  nand2 gate598(.a(gate35inter8), .b(gate35inter7), .O(gate35inter9));
  nand2 gate599(.a(s_7), .b(gate35inter3), .O(gate35inter10));
  nor2  gate600(.a(gate35inter10), .b(gate35inter9), .O(gate35inter11));
  nor2  gate601(.a(gate35inter11), .b(gate35inter6), .O(gate35inter12));
  nand2 gate602(.a(gate35inter12), .b(gate35inter1), .O(G344));

  xor2  gate2479(.a(G30), .b(G26), .O(gate36inter0));
  nand2 gate2480(.a(gate36inter0), .b(s_276), .O(gate36inter1));
  and2  gate2481(.a(G30), .b(G26), .O(gate36inter2));
  inv1  gate2482(.a(s_276), .O(gate36inter3));
  inv1  gate2483(.a(s_277), .O(gate36inter4));
  nand2 gate2484(.a(gate36inter4), .b(gate36inter3), .O(gate36inter5));
  nor2  gate2485(.a(gate36inter5), .b(gate36inter2), .O(gate36inter6));
  inv1  gate2486(.a(G26), .O(gate36inter7));
  inv1  gate2487(.a(G30), .O(gate36inter8));
  nand2 gate2488(.a(gate36inter8), .b(gate36inter7), .O(gate36inter9));
  nand2 gate2489(.a(s_277), .b(gate36inter3), .O(gate36inter10));
  nor2  gate2490(.a(gate36inter10), .b(gate36inter9), .O(gate36inter11));
  nor2  gate2491(.a(gate36inter11), .b(gate36inter6), .O(gate36inter12));
  nand2 gate2492(.a(gate36inter12), .b(gate36inter1), .O(G347));
nand2 gate37( .a(G19), .b(G23), .O(G350) );
nand2 gate38( .a(G27), .b(G31), .O(G353) );
nand2 gate39( .a(G20), .b(G24), .O(G356) );
nand2 gate40( .a(G28), .b(G32), .O(G359) );
nand2 gate41( .a(G1), .b(G266), .O(G362) );

  xor2  gate1863(.a(G266), .b(G2), .O(gate42inter0));
  nand2 gate1864(.a(gate42inter0), .b(s_188), .O(gate42inter1));
  and2  gate1865(.a(G266), .b(G2), .O(gate42inter2));
  inv1  gate1866(.a(s_188), .O(gate42inter3));
  inv1  gate1867(.a(s_189), .O(gate42inter4));
  nand2 gate1868(.a(gate42inter4), .b(gate42inter3), .O(gate42inter5));
  nor2  gate1869(.a(gate42inter5), .b(gate42inter2), .O(gate42inter6));
  inv1  gate1870(.a(G2), .O(gate42inter7));
  inv1  gate1871(.a(G266), .O(gate42inter8));
  nand2 gate1872(.a(gate42inter8), .b(gate42inter7), .O(gate42inter9));
  nand2 gate1873(.a(s_189), .b(gate42inter3), .O(gate42inter10));
  nor2  gate1874(.a(gate42inter10), .b(gate42inter9), .O(gate42inter11));
  nor2  gate1875(.a(gate42inter11), .b(gate42inter6), .O(gate42inter12));
  nand2 gate1876(.a(gate42inter12), .b(gate42inter1), .O(G363));

  xor2  gate2381(.a(G269), .b(G3), .O(gate43inter0));
  nand2 gate2382(.a(gate43inter0), .b(s_262), .O(gate43inter1));
  and2  gate2383(.a(G269), .b(G3), .O(gate43inter2));
  inv1  gate2384(.a(s_262), .O(gate43inter3));
  inv1  gate2385(.a(s_263), .O(gate43inter4));
  nand2 gate2386(.a(gate43inter4), .b(gate43inter3), .O(gate43inter5));
  nor2  gate2387(.a(gate43inter5), .b(gate43inter2), .O(gate43inter6));
  inv1  gate2388(.a(G3), .O(gate43inter7));
  inv1  gate2389(.a(G269), .O(gate43inter8));
  nand2 gate2390(.a(gate43inter8), .b(gate43inter7), .O(gate43inter9));
  nand2 gate2391(.a(s_263), .b(gate43inter3), .O(gate43inter10));
  nor2  gate2392(.a(gate43inter10), .b(gate43inter9), .O(gate43inter11));
  nor2  gate2393(.a(gate43inter11), .b(gate43inter6), .O(gate43inter12));
  nand2 gate2394(.a(gate43inter12), .b(gate43inter1), .O(G364));

  xor2  gate2339(.a(G269), .b(G4), .O(gate44inter0));
  nand2 gate2340(.a(gate44inter0), .b(s_256), .O(gate44inter1));
  and2  gate2341(.a(G269), .b(G4), .O(gate44inter2));
  inv1  gate2342(.a(s_256), .O(gate44inter3));
  inv1  gate2343(.a(s_257), .O(gate44inter4));
  nand2 gate2344(.a(gate44inter4), .b(gate44inter3), .O(gate44inter5));
  nor2  gate2345(.a(gate44inter5), .b(gate44inter2), .O(gate44inter6));
  inv1  gate2346(.a(G4), .O(gate44inter7));
  inv1  gate2347(.a(G269), .O(gate44inter8));
  nand2 gate2348(.a(gate44inter8), .b(gate44inter7), .O(gate44inter9));
  nand2 gate2349(.a(s_257), .b(gate44inter3), .O(gate44inter10));
  nor2  gate2350(.a(gate44inter10), .b(gate44inter9), .O(gate44inter11));
  nor2  gate2351(.a(gate44inter11), .b(gate44inter6), .O(gate44inter12));
  nand2 gate2352(.a(gate44inter12), .b(gate44inter1), .O(G365));
nand2 gate45( .a(G5), .b(G272), .O(G366) );
nand2 gate46( .a(G6), .b(G272), .O(G367) );

  xor2  gate771(.a(G275), .b(G7), .O(gate47inter0));
  nand2 gate772(.a(gate47inter0), .b(s_32), .O(gate47inter1));
  and2  gate773(.a(G275), .b(G7), .O(gate47inter2));
  inv1  gate774(.a(s_32), .O(gate47inter3));
  inv1  gate775(.a(s_33), .O(gate47inter4));
  nand2 gate776(.a(gate47inter4), .b(gate47inter3), .O(gate47inter5));
  nor2  gate777(.a(gate47inter5), .b(gate47inter2), .O(gate47inter6));
  inv1  gate778(.a(G7), .O(gate47inter7));
  inv1  gate779(.a(G275), .O(gate47inter8));
  nand2 gate780(.a(gate47inter8), .b(gate47inter7), .O(gate47inter9));
  nand2 gate781(.a(s_33), .b(gate47inter3), .O(gate47inter10));
  nor2  gate782(.a(gate47inter10), .b(gate47inter9), .O(gate47inter11));
  nor2  gate783(.a(gate47inter11), .b(gate47inter6), .O(gate47inter12));
  nand2 gate784(.a(gate47inter12), .b(gate47inter1), .O(G368));

  xor2  gate1289(.a(G275), .b(G8), .O(gate48inter0));
  nand2 gate1290(.a(gate48inter0), .b(s_106), .O(gate48inter1));
  and2  gate1291(.a(G275), .b(G8), .O(gate48inter2));
  inv1  gate1292(.a(s_106), .O(gate48inter3));
  inv1  gate1293(.a(s_107), .O(gate48inter4));
  nand2 gate1294(.a(gate48inter4), .b(gate48inter3), .O(gate48inter5));
  nor2  gate1295(.a(gate48inter5), .b(gate48inter2), .O(gate48inter6));
  inv1  gate1296(.a(G8), .O(gate48inter7));
  inv1  gate1297(.a(G275), .O(gate48inter8));
  nand2 gate1298(.a(gate48inter8), .b(gate48inter7), .O(gate48inter9));
  nand2 gate1299(.a(s_107), .b(gate48inter3), .O(gate48inter10));
  nor2  gate1300(.a(gate48inter10), .b(gate48inter9), .O(gate48inter11));
  nor2  gate1301(.a(gate48inter11), .b(gate48inter6), .O(gate48inter12));
  nand2 gate1302(.a(gate48inter12), .b(gate48inter1), .O(G369));

  xor2  gate925(.a(G278), .b(G9), .O(gate49inter0));
  nand2 gate926(.a(gate49inter0), .b(s_54), .O(gate49inter1));
  and2  gate927(.a(G278), .b(G9), .O(gate49inter2));
  inv1  gate928(.a(s_54), .O(gate49inter3));
  inv1  gate929(.a(s_55), .O(gate49inter4));
  nand2 gate930(.a(gate49inter4), .b(gate49inter3), .O(gate49inter5));
  nor2  gate931(.a(gate49inter5), .b(gate49inter2), .O(gate49inter6));
  inv1  gate932(.a(G9), .O(gate49inter7));
  inv1  gate933(.a(G278), .O(gate49inter8));
  nand2 gate934(.a(gate49inter8), .b(gate49inter7), .O(gate49inter9));
  nand2 gate935(.a(s_55), .b(gate49inter3), .O(gate49inter10));
  nor2  gate936(.a(gate49inter10), .b(gate49inter9), .O(gate49inter11));
  nor2  gate937(.a(gate49inter11), .b(gate49inter6), .O(gate49inter12));
  nand2 gate938(.a(gate49inter12), .b(gate49inter1), .O(G370));
nand2 gate50( .a(G10), .b(G278), .O(G371) );
nand2 gate51( .a(G11), .b(G281), .O(G372) );
nand2 gate52( .a(G12), .b(G281), .O(G373) );
nand2 gate53( .a(G13), .b(G284), .O(G374) );
nand2 gate54( .a(G14), .b(G284), .O(G375) );
nand2 gate55( .a(G15), .b(G287), .O(G376) );
nand2 gate56( .a(G16), .b(G287), .O(G377) );

  xor2  gate1807(.a(G290), .b(G17), .O(gate57inter0));
  nand2 gate1808(.a(gate57inter0), .b(s_180), .O(gate57inter1));
  and2  gate1809(.a(G290), .b(G17), .O(gate57inter2));
  inv1  gate1810(.a(s_180), .O(gate57inter3));
  inv1  gate1811(.a(s_181), .O(gate57inter4));
  nand2 gate1812(.a(gate57inter4), .b(gate57inter3), .O(gate57inter5));
  nor2  gate1813(.a(gate57inter5), .b(gate57inter2), .O(gate57inter6));
  inv1  gate1814(.a(G17), .O(gate57inter7));
  inv1  gate1815(.a(G290), .O(gate57inter8));
  nand2 gate1816(.a(gate57inter8), .b(gate57inter7), .O(gate57inter9));
  nand2 gate1817(.a(s_181), .b(gate57inter3), .O(gate57inter10));
  nor2  gate1818(.a(gate57inter10), .b(gate57inter9), .O(gate57inter11));
  nor2  gate1819(.a(gate57inter11), .b(gate57inter6), .O(gate57inter12));
  nand2 gate1820(.a(gate57inter12), .b(gate57inter1), .O(G378));
nand2 gate58( .a(G18), .b(G290), .O(G379) );
nand2 gate59( .a(G19), .b(G293), .O(G380) );
nand2 gate60( .a(G20), .b(G293), .O(G381) );
nand2 gate61( .a(G21), .b(G296), .O(G382) );
nand2 gate62( .a(G22), .b(G296), .O(G383) );
nand2 gate63( .a(G23), .b(G299), .O(G384) );

  xor2  gate1009(.a(G299), .b(G24), .O(gate64inter0));
  nand2 gate1010(.a(gate64inter0), .b(s_66), .O(gate64inter1));
  and2  gate1011(.a(G299), .b(G24), .O(gate64inter2));
  inv1  gate1012(.a(s_66), .O(gate64inter3));
  inv1  gate1013(.a(s_67), .O(gate64inter4));
  nand2 gate1014(.a(gate64inter4), .b(gate64inter3), .O(gate64inter5));
  nor2  gate1015(.a(gate64inter5), .b(gate64inter2), .O(gate64inter6));
  inv1  gate1016(.a(G24), .O(gate64inter7));
  inv1  gate1017(.a(G299), .O(gate64inter8));
  nand2 gate1018(.a(gate64inter8), .b(gate64inter7), .O(gate64inter9));
  nand2 gate1019(.a(s_67), .b(gate64inter3), .O(gate64inter10));
  nor2  gate1020(.a(gate64inter10), .b(gate64inter9), .O(gate64inter11));
  nor2  gate1021(.a(gate64inter11), .b(gate64inter6), .O(gate64inter12));
  nand2 gate1022(.a(gate64inter12), .b(gate64inter1), .O(G385));
nand2 gate65( .a(G25), .b(G302), .O(G386) );
nand2 gate66( .a(G26), .b(G302), .O(G387) );
nand2 gate67( .a(G27), .b(G305), .O(G388) );
nand2 gate68( .a(G28), .b(G305), .O(G389) );

  xor2  gate2367(.a(G308), .b(G29), .O(gate69inter0));
  nand2 gate2368(.a(gate69inter0), .b(s_260), .O(gate69inter1));
  and2  gate2369(.a(G308), .b(G29), .O(gate69inter2));
  inv1  gate2370(.a(s_260), .O(gate69inter3));
  inv1  gate2371(.a(s_261), .O(gate69inter4));
  nand2 gate2372(.a(gate69inter4), .b(gate69inter3), .O(gate69inter5));
  nor2  gate2373(.a(gate69inter5), .b(gate69inter2), .O(gate69inter6));
  inv1  gate2374(.a(G29), .O(gate69inter7));
  inv1  gate2375(.a(G308), .O(gate69inter8));
  nand2 gate2376(.a(gate69inter8), .b(gate69inter7), .O(gate69inter9));
  nand2 gate2377(.a(s_261), .b(gate69inter3), .O(gate69inter10));
  nor2  gate2378(.a(gate69inter10), .b(gate69inter9), .O(gate69inter11));
  nor2  gate2379(.a(gate69inter11), .b(gate69inter6), .O(gate69inter12));
  nand2 gate2380(.a(gate69inter12), .b(gate69inter1), .O(G390));
nand2 gate70( .a(G30), .b(G308), .O(G391) );

  xor2  gate799(.a(G311), .b(G31), .O(gate71inter0));
  nand2 gate800(.a(gate71inter0), .b(s_36), .O(gate71inter1));
  and2  gate801(.a(G311), .b(G31), .O(gate71inter2));
  inv1  gate802(.a(s_36), .O(gate71inter3));
  inv1  gate803(.a(s_37), .O(gate71inter4));
  nand2 gate804(.a(gate71inter4), .b(gate71inter3), .O(gate71inter5));
  nor2  gate805(.a(gate71inter5), .b(gate71inter2), .O(gate71inter6));
  inv1  gate806(.a(G31), .O(gate71inter7));
  inv1  gate807(.a(G311), .O(gate71inter8));
  nand2 gate808(.a(gate71inter8), .b(gate71inter7), .O(gate71inter9));
  nand2 gate809(.a(s_37), .b(gate71inter3), .O(gate71inter10));
  nor2  gate810(.a(gate71inter10), .b(gate71inter9), .O(gate71inter11));
  nor2  gate811(.a(gate71inter11), .b(gate71inter6), .O(gate71inter12));
  nand2 gate812(.a(gate71inter12), .b(gate71inter1), .O(G392));
nand2 gate72( .a(G32), .b(G311), .O(G393) );

  xor2  gate1079(.a(G314), .b(G1), .O(gate73inter0));
  nand2 gate1080(.a(gate73inter0), .b(s_76), .O(gate73inter1));
  and2  gate1081(.a(G314), .b(G1), .O(gate73inter2));
  inv1  gate1082(.a(s_76), .O(gate73inter3));
  inv1  gate1083(.a(s_77), .O(gate73inter4));
  nand2 gate1084(.a(gate73inter4), .b(gate73inter3), .O(gate73inter5));
  nor2  gate1085(.a(gate73inter5), .b(gate73inter2), .O(gate73inter6));
  inv1  gate1086(.a(G1), .O(gate73inter7));
  inv1  gate1087(.a(G314), .O(gate73inter8));
  nand2 gate1088(.a(gate73inter8), .b(gate73inter7), .O(gate73inter9));
  nand2 gate1089(.a(s_77), .b(gate73inter3), .O(gate73inter10));
  nor2  gate1090(.a(gate73inter10), .b(gate73inter9), .O(gate73inter11));
  nor2  gate1091(.a(gate73inter11), .b(gate73inter6), .O(gate73inter12));
  nand2 gate1092(.a(gate73inter12), .b(gate73inter1), .O(G394));

  xor2  gate575(.a(G314), .b(G5), .O(gate74inter0));
  nand2 gate576(.a(gate74inter0), .b(s_4), .O(gate74inter1));
  and2  gate577(.a(G314), .b(G5), .O(gate74inter2));
  inv1  gate578(.a(s_4), .O(gate74inter3));
  inv1  gate579(.a(s_5), .O(gate74inter4));
  nand2 gate580(.a(gate74inter4), .b(gate74inter3), .O(gate74inter5));
  nor2  gate581(.a(gate74inter5), .b(gate74inter2), .O(gate74inter6));
  inv1  gate582(.a(G5), .O(gate74inter7));
  inv1  gate583(.a(G314), .O(gate74inter8));
  nand2 gate584(.a(gate74inter8), .b(gate74inter7), .O(gate74inter9));
  nand2 gate585(.a(s_5), .b(gate74inter3), .O(gate74inter10));
  nor2  gate586(.a(gate74inter10), .b(gate74inter9), .O(gate74inter11));
  nor2  gate587(.a(gate74inter11), .b(gate74inter6), .O(gate74inter12));
  nand2 gate588(.a(gate74inter12), .b(gate74inter1), .O(G395));
nand2 gate75( .a(G9), .b(G317), .O(G396) );
nand2 gate76( .a(G13), .b(G317), .O(G397) );
nand2 gate77( .a(G2), .b(G320), .O(G398) );
nand2 gate78( .a(G6), .b(G320), .O(G399) );

  xor2  gate2451(.a(G323), .b(G10), .O(gate79inter0));
  nand2 gate2452(.a(gate79inter0), .b(s_272), .O(gate79inter1));
  and2  gate2453(.a(G323), .b(G10), .O(gate79inter2));
  inv1  gate2454(.a(s_272), .O(gate79inter3));
  inv1  gate2455(.a(s_273), .O(gate79inter4));
  nand2 gate2456(.a(gate79inter4), .b(gate79inter3), .O(gate79inter5));
  nor2  gate2457(.a(gate79inter5), .b(gate79inter2), .O(gate79inter6));
  inv1  gate2458(.a(G10), .O(gate79inter7));
  inv1  gate2459(.a(G323), .O(gate79inter8));
  nand2 gate2460(.a(gate79inter8), .b(gate79inter7), .O(gate79inter9));
  nand2 gate2461(.a(s_273), .b(gate79inter3), .O(gate79inter10));
  nor2  gate2462(.a(gate79inter10), .b(gate79inter9), .O(gate79inter11));
  nor2  gate2463(.a(gate79inter11), .b(gate79inter6), .O(gate79inter12));
  nand2 gate2464(.a(gate79inter12), .b(gate79inter1), .O(G400));
nand2 gate80( .a(G14), .b(G323), .O(G401) );

  xor2  gate2283(.a(G326), .b(G3), .O(gate81inter0));
  nand2 gate2284(.a(gate81inter0), .b(s_248), .O(gate81inter1));
  and2  gate2285(.a(G326), .b(G3), .O(gate81inter2));
  inv1  gate2286(.a(s_248), .O(gate81inter3));
  inv1  gate2287(.a(s_249), .O(gate81inter4));
  nand2 gate2288(.a(gate81inter4), .b(gate81inter3), .O(gate81inter5));
  nor2  gate2289(.a(gate81inter5), .b(gate81inter2), .O(gate81inter6));
  inv1  gate2290(.a(G3), .O(gate81inter7));
  inv1  gate2291(.a(G326), .O(gate81inter8));
  nand2 gate2292(.a(gate81inter8), .b(gate81inter7), .O(gate81inter9));
  nand2 gate2293(.a(s_249), .b(gate81inter3), .O(gate81inter10));
  nor2  gate2294(.a(gate81inter10), .b(gate81inter9), .O(gate81inter11));
  nor2  gate2295(.a(gate81inter11), .b(gate81inter6), .O(gate81inter12));
  nand2 gate2296(.a(gate81inter12), .b(gate81inter1), .O(G402));
nand2 gate82( .a(G7), .b(G326), .O(G403) );

  xor2  gate981(.a(G329), .b(G11), .O(gate83inter0));
  nand2 gate982(.a(gate83inter0), .b(s_62), .O(gate83inter1));
  and2  gate983(.a(G329), .b(G11), .O(gate83inter2));
  inv1  gate984(.a(s_62), .O(gate83inter3));
  inv1  gate985(.a(s_63), .O(gate83inter4));
  nand2 gate986(.a(gate83inter4), .b(gate83inter3), .O(gate83inter5));
  nor2  gate987(.a(gate83inter5), .b(gate83inter2), .O(gate83inter6));
  inv1  gate988(.a(G11), .O(gate83inter7));
  inv1  gate989(.a(G329), .O(gate83inter8));
  nand2 gate990(.a(gate83inter8), .b(gate83inter7), .O(gate83inter9));
  nand2 gate991(.a(s_63), .b(gate83inter3), .O(gate83inter10));
  nor2  gate992(.a(gate83inter10), .b(gate83inter9), .O(gate83inter11));
  nor2  gate993(.a(gate83inter11), .b(gate83inter6), .O(gate83inter12));
  nand2 gate994(.a(gate83inter12), .b(gate83inter1), .O(G404));
nand2 gate84( .a(G15), .b(G329), .O(G405) );
nand2 gate85( .a(G4), .b(G332), .O(G406) );
nand2 gate86( .a(G8), .b(G332), .O(G407) );
nand2 gate87( .a(G12), .b(G335), .O(G408) );
nand2 gate88( .a(G16), .b(G335), .O(G409) );

  xor2  gate2171(.a(G338), .b(G17), .O(gate89inter0));
  nand2 gate2172(.a(gate89inter0), .b(s_232), .O(gate89inter1));
  and2  gate2173(.a(G338), .b(G17), .O(gate89inter2));
  inv1  gate2174(.a(s_232), .O(gate89inter3));
  inv1  gate2175(.a(s_233), .O(gate89inter4));
  nand2 gate2176(.a(gate89inter4), .b(gate89inter3), .O(gate89inter5));
  nor2  gate2177(.a(gate89inter5), .b(gate89inter2), .O(gate89inter6));
  inv1  gate2178(.a(G17), .O(gate89inter7));
  inv1  gate2179(.a(G338), .O(gate89inter8));
  nand2 gate2180(.a(gate89inter8), .b(gate89inter7), .O(gate89inter9));
  nand2 gate2181(.a(s_233), .b(gate89inter3), .O(gate89inter10));
  nor2  gate2182(.a(gate89inter10), .b(gate89inter9), .O(gate89inter11));
  nor2  gate2183(.a(gate89inter11), .b(gate89inter6), .O(gate89inter12));
  nand2 gate2184(.a(gate89inter12), .b(gate89inter1), .O(G410));
nand2 gate90( .a(G21), .b(G338), .O(G411) );

  xor2  gate2101(.a(G341), .b(G25), .O(gate91inter0));
  nand2 gate2102(.a(gate91inter0), .b(s_222), .O(gate91inter1));
  and2  gate2103(.a(G341), .b(G25), .O(gate91inter2));
  inv1  gate2104(.a(s_222), .O(gate91inter3));
  inv1  gate2105(.a(s_223), .O(gate91inter4));
  nand2 gate2106(.a(gate91inter4), .b(gate91inter3), .O(gate91inter5));
  nor2  gate2107(.a(gate91inter5), .b(gate91inter2), .O(gate91inter6));
  inv1  gate2108(.a(G25), .O(gate91inter7));
  inv1  gate2109(.a(G341), .O(gate91inter8));
  nand2 gate2110(.a(gate91inter8), .b(gate91inter7), .O(gate91inter9));
  nand2 gate2111(.a(s_223), .b(gate91inter3), .O(gate91inter10));
  nor2  gate2112(.a(gate91inter10), .b(gate91inter9), .O(gate91inter11));
  nor2  gate2113(.a(gate91inter11), .b(gate91inter6), .O(gate91inter12));
  nand2 gate2114(.a(gate91inter12), .b(gate91inter1), .O(G412));
nand2 gate92( .a(G29), .b(G341), .O(G413) );
nand2 gate93( .a(G18), .b(G344), .O(G414) );
nand2 gate94( .a(G22), .b(G344), .O(G415) );
nand2 gate95( .a(G26), .b(G347), .O(G416) );

  xor2  gate2031(.a(G347), .b(G30), .O(gate96inter0));
  nand2 gate2032(.a(gate96inter0), .b(s_212), .O(gate96inter1));
  and2  gate2033(.a(G347), .b(G30), .O(gate96inter2));
  inv1  gate2034(.a(s_212), .O(gate96inter3));
  inv1  gate2035(.a(s_213), .O(gate96inter4));
  nand2 gate2036(.a(gate96inter4), .b(gate96inter3), .O(gate96inter5));
  nor2  gate2037(.a(gate96inter5), .b(gate96inter2), .O(gate96inter6));
  inv1  gate2038(.a(G30), .O(gate96inter7));
  inv1  gate2039(.a(G347), .O(gate96inter8));
  nand2 gate2040(.a(gate96inter8), .b(gate96inter7), .O(gate96inter9));
  nand2 gate2041(.a(s_213), .b(gate96inter3), .O(gate96inter10));
  nor2  gate2042(.a(gate96inter10), .b(gate96inter9), .O(gate96inter11));
  nor2  gate2043(.a(gate96inter11), .b(gate96inter6), .O(gate96inter12));
  nand2 gate2044(.a(gate96inter12), .b(gate96inter1), .O(G417));
nand2 gate97( .a(G19), .b(G350), .O(G418) );
nand2 gate98( .a(G23), .b(G350), .O(G419) );
nand2 gate99( .a(G27), .b(G353), .O(G420) );

  xor2  gate2143(.a(G353), .b(G31), .O(gate100inter0));
  nand2 gate2144(.a(gate100inter0), .b(s_228), .O(gate100inter1));
  and2  gate2145(.a(G353), .b(G31), .O(gate100inter2));
  inv1  gate2146(.a(s_228), .O(gate100inter3));
  inv1  gate2147(.a(s_229), .O(gate100inter4));
  nand2 gate2148(.a(gate100inter4), .b(gate100inter3), .O(gate100inter5));
  nor2  gate2149(.a(gate100inter5), .b(gate100inter2), .O(gate100inter6));
  inv1  gate2150(.a(G31), .O(gate100inter7));
  inv1  gate2151(.a(G353), .O(gate100inter8));
  nand2 gate2152(.a(gate100inter8), .b(gate100inter7), .O(gate100inter9));
  nand2 gate2153(.a(s_229), .b(gate100inter3), .O(gate100inter10));
  nor2  gate2154(.a(gate100inter10), .b(gate100inter9), .O(gate100inter11));
  nor2  gate2155(.a(gate100inter11), .b(gate100inter6), .O(gate100inter12));
  nand2 gate2156(.a(gate100inter12), .b(gate100inter1), .O(G421));

  xor2  gate715(.a(G356), .b(G20), .O(gate101inter0));
  nand2 gate716(.a(gate101inter0), .b(s_24), .O(gate101inter1));
  and2  gate717(.a(G356), .b(G20), .O(gate101inter2));
  inv1  gate718(.a(s_24), .O(gate101inter3));
  inv1  gate719(.a(s_25), .O(gate101inter4));
  nand2 gate720(.a(gate101inter4), .b(gate101inter3), .O(gate101inter5));
  nor2  gate721(.a(gate101inter5), .b(gate101inter2), .O(gate101inter6));
  inv1  gate722(.a(G20), .O(gate101inter7));
  inv1  gate723(.a(G356), .O(gate101inter8));
  nand2 gate724(.a(gate101inter8), .b(gate101inter7), .O(gate101inter9));
  nand2 gate725(.a(s_25), .b(gate101inter3), .O(gate101inter10));
  nor2  gate726(.a(gate101inter10), .b(gate101inter9), .O(gate101inter11));
  nor2  gate727(.a(gate101inter11), .b(gate101inter6), .O(gate101inter12));
  nand2 gate728(.a(gate101inter12), .b(gate101inter1), .O(G422));
nand2 gate102( .a(G24), .b(G356), .O(G423) );

  xor2  gate2703(.a(G359), .b(G28), .O(gate103inter0));
  nand2 gate2704(.a(gate103inter0), .b(s_308), .O(gate103inter1));
  and2  gate2705(.a(G359), .b(G28), .O(gate103inter2));
  inv1  gate2706(.a(s_308), .O(gate103inter3));
  inv1  gate2707(.a(s_309), .O(gate103inter4));
  nand2 gate2708(.a(gate103inter4), .b(gate103inter3), .O(gate103inter5));
  nor2  gate2709(.a(gate103inter5), .b(gate103inter2), .O(gate103inter6));
  inv1  gate2710(.a(G28), .O(gate103inter7));
  inv1  gate2711(.a(G359), .O(gate103inter8));
  nand2 gate2712(.a(gate103inter8), .b(gate103inter7), .O(gate103inter9));
  nand2 gate2713(.a(s_309), .b(gate103inter3), .O(gate103inter10));
  nor2  gate2714(.a(gate103inter10), .b(gate103inter9), .O(gate103inter11));
  nor2  gate2715(.a(gate103inter11), .b(gate103inter6), .O(gate103inter12));
  nand2 gate2716(.a(gate103inter12), .b(gate103inter1), .O(G424));

  xor2  gate1415(.a(G359), .b(G32), .O(gate104inter0));
  nand2 gate1416(.a(gate104inter0), .b(s_124), .O(gate104inter1));
  and2  gate1417(.a(G359), .b(G32), .O(gate104inter2));
  inv1  gate1418(.a(s_124), .O(gate104inter3));
  inv1  gate1419(.a(s_125), .O(gate104inter4));
  nand2 gate1420(.a(gate104inter4), .b(gate104inter3), .O(gate104inter5));
  nor2  gate1421(.a(gate104inter5), .b(gate104inter2), .O(gate104inter6));
  inv1  gate1422(.a(G32), .O(gate104inter7));
  inv1  gate1423(.a(G359), .O(gate104inter8));
  nand2 gate1424(.a(gate104inter8), .b(gate104inter7), .O(gate104inter9));
  nand2 gate1425(.a(s_125), .b(gate104inter3), .O(gate104inter10));
  nor2  gate1426(.a(gate104inter10), .b(gate104inter9), .O(gate104inter11));
  nor2  gate1427(.a(gate104inter11), .b(gate104inter6), .O(gate104inter12));
  nand2 gate1428(.a(gate104inter12), .b(gate104inter1), .O(G425));
nand2 gate105( .a(G362), .b(G363), .O(G426) );
nand2 gate106( .a(G364), .b(G365), .O(G429) );
nand2 gate107( .a(G366), .b(G367), .O(G432) );
nand2 gate108( .a(G368), .b(G369), .O(G435) );
nand2 gate109( .a(G370), .b(G371), .O(G438) );

  xor2  gate995(.a(G373), .b(G372), .O(gate110inter0));
  nand2 gate996(.a(gate110inter0), .b(s_64), .O(gate110inter1));
  and2  gate997(.a(G373), .b(G372), .O(gate110inter2));
  inv1  gate998(.a(s_64), .O(gate110inter3));
  inv1  gate999(.a(s_65), .O(gate110inter4));
  nand2 gate1000(.a(gate110inter4), .b(gate110inter3), .O(gate110inter5));
  nor2  gate1001(.a(gate110inter5), .b(gate110inter2), .O(gate110inter6));
  inv1  gate1002(.a(G372), .O(gate110inter7));
  inv1  gate1003(.a(G373), .O(gate110inter8));
  nand2 gate1004(.a(gate110inter8), .b(gate110inter7), .O(gate110inter9));
  nand2 gate1005(.a(s_65), .b(gate110inter3), .O(gate110inter10));
  nor2  gate1006(.a(gate110inter10), .b(gate110inter9), .O(gate110inter11));
  nor2  gate1007(.a(gate110inter11), .b(gate110inter6), .O(gate110inter12));
  nand2 gate1008(.a(gate110inter12), .b(gate110inter1), .O(G441));
nand2 gate111( .a(G374), .b(G375), .O(G444) );
nand2 gate112( .a(G376), .b(G377), .O(G447) );

  xor2  gate1947(.a(G379), .b(G378), .O(gate113inter0));
  nand2 gate1948(.a(gate113inter0), .b(s_200), .O(gate113inter1));
  and2  gate1949(.a(G379), .b(G378), .O(gate113inter2));
  inv1  gate1950(.a(s_200), .O(gate113inter3));
  inv1  gate1951(.a(s_201), .O(gate113inter4));
  nand2 gate1952(.a(gate113inter4), .b(gate113inter3), .O(gate113inter5));
  nor2  gate1953(.a(gate113inter5), .b(gate113inter2), .O(gate113inter6));
  inv1  gate1954(.a(G378), .O(gate113inter7));
  inv1  gate1955(.a(G379), .O(gate113inter8));
  nand2 gate1956(.a(gate113inter8), .b(gate113inter7), .O(gate113inter9));
  nand2 gate1957(.a(s_201), .b(gate113inter3), .O(gate113inter10));
  nor2  gate1958(.a(gate113inter10), .b(gate113inter9), .O(gate113inter11));
  nor2  gate1959(.a(gate113inter11), .b(gate113inter6), .O(gate113inter12));
  nand2 gate1960(.a(gate113inter12), .b(gate113inter1), .O(G450));
nand2 gate114( .a(G380), .b(G381), .O(G453) );

  xor2  gate1639(.a(G383), .b(G382), .O(gate115inter0));
  nand2 gate1640(.a(gate115inter0), .b(s_156), .O(gate115inter1));
  and2  gate1641(.a(G383), .b(G382), .O(gate115inter2));
  inv1  gate1642(.a(s_156), .O(gate115inter3));
  inv1  gate1643(.a(s_157), .O(gate115inter4));
  nand2 gate1644(.a(gate115inter4), .b(gate115inter3), .O(gate115inter5));
  nor2  gate1645(.a(gate115inter5), .b(gate115inter2), .O(gate115inter6));
  inv1  gate1646(.a(G382), .O(gate115inter7));
  inv1  gate1647(.a(G383), .O(gate115inter8));
  nand2 gate1648(.a(gate115inter8), .b(gate115inter7), .O(gate115inter9));
  nand2 gate1649(.a(s_157), .b(gate115inter3), .O(gate115inter10));
  nor2  gate1650(.a(gate115inter10), .b(gate115inter9), .O(gate115inter11));
  nor2  gate1651(.a(gate115inter11), .b(gate115inter6), .O(gate115inter12));
  nand2 gate1652(.a(gate115inter12), .b(gate115inter1), .O(G456));
nand2 gate116( .a(G384), .b(G385), .O(G459) );
nand2 gate117( .a(G386), .b(G387), .O(G462) );
nand2 gate118( .a(G388), .b(G389), .O(G465) );

  xor2  gate1499(.a(G391), .b(G390), .O(gate119inter0));
  nand2 gate1500(.a(gate119inter0), .b(s_136), .O(gate119inter1));
  and2  gate1501(.a(G391), .b(G390), .O(gate119inter2));
  inv1  gate1502(.a(s_136), .O(gate119inter3));
  inv1  gate1503(.a(s_137), .O(gate119inter4));
  nand2 gate1504(.a(gate119inter4), .b(gate119inter3), .O(gate119inter5));
  nor2  gate1505(.a(gate119inter5), .b(gate119inter2), .O(gate119inter6));
  inv1  gate1506(.a(G390), .O(gate119inter7));
  inv1  gate1507(.a(G391), .O(gate119inter8));
  nand2 gate1508(.a(gate119inter8), .b(gate119inter7), .O(gate119inter9));
  nand2 gate1509(.a(s_137), .b(gate119inter3), .O(gate119inter10));
  nor2  gate1510(.a(gate119inter10), .b(gate119inter9), .O(gate119inter11));
  nor2  gate1511(.a(gate119inter11), .b(gate119inter6), .O(gate119inter12));
  nand2 gate1512(.a(gate119inter12), .b(gate119inter1), .O(G468));
nand2 gate120( .a(G392), .b(G393), .O(G471) );
nand2 gate121( .a(G394), .b(G395), .O(G474) );

  xor2  gate1891(.a(G397), .b(G396), .O(gate122inter0));
  nand2 gate1892(.a(gate122inter0), .b(s_192), .O(gate122inter1));
  and2  gate1893(.a(G397), .b(G396), .O(gate122inter2));
  inv1  gate1894(.a(s_192), .O(gate122inter3));
  inv1  gate1895(.a(s_193), .O(gate122inter4));
  nand2 gate1896(.a(gate122inter4), .b(gate122inter3), .O(gate122inter5));
  nor2  gate1897(.a(gate122inter5), .b(gate122inter2), .O(gate122inter6));
  inv1  gate1898(.a(G396), .O(gate122inter7));
  inv1  gate1899(.a(G397), .O(gate122inter8));
  nand2 gate1900(.a(gate122inter8), .b(gate122inter7), .O(gate122inter9));
  nand2 gate1901(.a(s_193), .b(gate122inter3), .O(gate122inter10));
  nor2  gate1902(.a(gate122inter10), .b(gate122inter9), .O(gate122inter11));
  nor2  gate1903(.a(gate122inter11), .b(gate122inter6), .O(gate122inter12));
  nand2 gate1904(.a(gate122inter12), .b(gate122inter1), .O(G477));
nand2 gate123( .a(G398), .b(G399), .O(G480) );

  xor2  gate617(.a(G401), .b(G400), .O(gate124inter0));
  nand2 gate618(.a(gate124inter0), .b(s_10), .O(gate124inter1));
  and2  gate619(.a(G401), .b(G400), .O(gate124inter2));
  inv1  gate620(.a(s_10), .O(gate124inter3));
  inv1  gate621(.a(s_11), .O(gate124inter4));
  nand2 gate622(.a(gate124inter4), .b(gate124inter3), .O(gate124inter5));
  nor2  gate623(.a(gate124inter5), .b(gate124inter2), .O(gate124inter6));
  inv1  gate624(.a(G400), .O(gate124inter7));
  inv1  gate625(.a(G401), .O(gate124inter8));
  nand2 gate626(.a(gate124inter8), .b(gate124inter7), .O(gate124inter9));
  nand2 gate627(.a(s_11), .b(gate124inter3), .O(gate124inter10));
  nor2  gate628(.a(gate124inter10), .b(gate124inter9), .O(gate124inter11));
  nor2  gate629(.a(gate124inter11), .b(gate124inter6), .O(gate124inter12));
  nand2 gate630(.a(gate124inter12), .b(gate124inter1), .O(G483));
nand2 gate125( .a(G402), .b(G403), .O(G486) );
nand2 gate126( .a(G404), .b(G405), .O(G489) );
nand2 gate127( .a(G406), .b(G407), .O(G492) );

  xor2  gate883(.a(G409), .b(G408), .O(gate128inter0));
  nand2 gate884(.a(gate128inter0), .b(s_48), .O(gate128inter1));
  and2  gate885(.a(G409), .b(G408), .O(gate128inter2));
  inv1  gate886(.a(s_48), .O(gate128inter3));
  inv1  gate887(.a(s_49), .O(gate128inter4));
  nand2 gate888(.a(gate128inter4), .b(gate128inter3), .O(gate128inter5));
  nor2  gate889(.a(gate128inter5), .b(gate128inter2), .O(gate128inter6));
  inv1  gate890(.a(G408), .O(gate128inter7));
  inv1  gate891(.a(G409), .O(gate128inter8));
  nand2 gate892(.a(gate128inter8), .b(gate128inter7), .O(gate128inter9));
  nand2 gate893(.a(s_49), .b(gate128inter3), .O(gate128inter10));
  nor2  gate894(.a(gate128inter10), .b(gate128inter9), .O(gate128inter11));
  nor2  gate895(.a(gate128inter11), .b(gate128inter6), .O(gate128inter12));
  nand2 gate896(.a(gate128inter12), .b(gate128inter1), .O(G495));

  xor2  gate2493(.a(G411), .b(G410), .O(gate129inter0));
  nand2 gate2494(.a(gate129inter0), .b(s_278), .O(gate129inter1));
  and2  gate2495(.a(G411), .b(G410), .O(gate129inter2));
  inv1  gate2496(.a(s_278), .O(gate129inter3));
  inv1  gate2497(.a(s_279), .O(gate129inter4));
  nand2 gate2498(.a(gate129inter4), .b(gate129inter3), .O(gate129inter5));
  nor2  gate2499(.a(gate129inter5), .b(gate129inter2), .O(gate129inter6));
  inv1  gate2500(.a(G410), .O(gate129inter7));
  inv1  gate2501(.a(G411), .O(gate129inter8));
  nand2 gate2502(.a(gate129inter8), .b(gate129inter7), .O(gate129inter9));
  nand2 gate2503(.a(s_279), .b(gate129inter3), .O(gate129inter10));
  nor2  gate2504(.a(gate129inter10), .b(gate129inter9), .O(gate129inter11));
  nor2  gate2505(.a(gate129inter11), .b(gate129inter6), .O(gate129inter12));
  nand2 gate2506(.a(gate129inter12), .b(gate129inter1), .O(G498));

  xor2  gate2577(.a(G413), .b(G412), .O(gate130inter0));
  nand2 gate2578(.a(gate130inter0), .b(s_290), .O(gate130inter1));
  and2  gate2579(.a(G413), .b(G412), .O(gate130inter2));
  inv1  gate2580(.a(s_290), .O(gate130inter3));
  inv1  gate2581(.a(s_291), .O(gate130inter4));
  nand2 gate2582(.a(gate130inter4), .b(gate130inter3), .O(gate130inter5));
  nor2  gate2583(.a(gate130inter5), .b(gate130inter2), .O(gate130inter6));
  inv1  gate2584(.a(G412), .O(gate130inter7));
  inv1  gate2585(.a(G413), .O(gate130inter8));
  nand2 gate2586(.a(gate130inter8), .b(gate130inter7), .O(gate130inter9));
  nand2 gate2587(.a(s_291), .b(gate130inter3), .O(gate130inter10));
  nor2  gate2588(.a(gate130inter10), .b(gate130inter9), .O(gate130inter11));
  nor2  gate2589(.a(gate130inter11), .b(gate130inter6), .O(gate130inter12));
  nand2 gate2590(.a(gate130inter12), .b(gate130inter1), .O(G501));

  xor2  gate1457(.a(G415), .b(G414), .O(gate131inter0));
  nand2 gate1458(.a(gate131inter0), .b(s_130), .O(gate131inter1));
  and2  gate1459(.a(G415), .b(G414), .O(gate131inter2));
  inv1  gate1460(.a(s_130), .O(gate131inter3));
  inv1  gate1461(.a(s_131), .O(gate131inter4));
  nand2 gate1462(.a(gate131inter4), .b(gate131inter3), .O(gate131inter5));
  nor2  gate1463(.a(gate131inter5), .b(gate131inter2), .O(gate131inter6));
  inv1  gate1464(.a(G414), .O(gate131inter7));
  inv1  gate1465(.a(G415), .O(gate131inter8));
  nand2 gate1466(.a(gate131inter8), .b(gate131inter7), .O(gate131inter9));
  nand2 gate1467(.a(s_131), .b(gate131inter3), .O(gate131inter10));
  nor2  gate1468(.a(gate131inter10), .b(gate131inter9), .O(gate131inter11));
  nor2  gate1469(.a(gate131inter11), .b(gate131inter6), .O(gate131inter12));
  nand2 gate1470(.a(gate131inter12), .b(gate131inter1), .O(G504));
nand2 gate132( .a(G416), .b(G417), .O(G507) );
nand2 gate133( .a(G418), .b(G419), .O(G510) );
nand2 gate134( .a(G420), .b(G421), .O(G513) );

  xor2  gate2647(.a(G423), .b(G422), .O(gate135inter0));
  nand2 gate2648(.a(gate135inter0), .b(s_300), .O(gate135inter1));
  and2  gate2649(.a(G423), .b(G422), .O(gate135inter2));
  inv1  gate2650(.a(s_300), .O(gate135inter3));
  inv1  gate2651(.a(s_301), .O(gate135inter4));
  nand2 gate2652(.a(gate135inter4), .b(gate135inter3), .O(gate135inter5));
  nor2  gate2653(.a(gate135inter5), .b(gate135inter2), .O(gate135inter6));
  inv1  gate2654(.a(G422), .O(gate135inter7));
  inv1  gate2655(.a(G423), .O(gate135inter8));
  nand2 gate2656(.a(gate135inter8), .b(gate135inter7), .O(gate135inter9));
  nand2 gate2657(.a(s_301), .b(gate135inter3), .O(gate135inter10));
  nor2  gate2658(.a(gate135inter10), .b(gate135inter9), .O(gate135inter11));
  nor2  gate2659(.a(gate135inter11), .b(gate135inter6), .O(gate135inter12));
  nand2 gate2660(.a(gate135inter12), .b(gate135inter1), .O(G516));

  xor2  gate1051(.a(G425), .b(G424), .O(gate136inter0));
  nand2 gate1052(.a(gate136inter0), .b(s_72), .O(gate136inter1));
  and2  gate1053(.a(G425), .b(G424), .O(gate136inter2));
  inv1  gate1054(.a(s_72), .O(gate136inter3));
  inv1  gate1055(.a(s_73), .O(gate136inter4));
  nand2 gate1056(.a(gate136inter4), .b(gate136inter3), .O(gate136inter5));
  nor2  gate1057(.a(gate136inter5), .b(gate136inter2), .O(gate136inter6));
  inv1  gate1058(.a(G424), .O(gate136inter7));
  inv1  gate1059(.a(G425), .O(gate136inter8));
  nand2 gate1060(.a(gate136inter8), .b(gate136inter7), .O(gate136inter9));
  nand2 gate1061(.a(s_73), .b(gate136inter3), .O(gate136inter10));
  nor2  gate1062(.a(gate136inter10), .b(gate136inter9), .O(gate136inter11));
  nor2  gate1063(.a(gate136inter11), .b(gate136inter6), .O(gate136inter12));
  nand2 gate1064(.a(gate136inter12), .b(gate136inter1), .O(G519));

  xor2  gate2409(.a(G429), .b(G426), .O(gate137inter0));
  nand2 gate2410(.a(gate137inter0), .b(s_266), .O(gate137inter1));
  and2  gate2411(.a(G429), .b(G426), .O(gate137inter2));
  inv1  gate2412(.a(s_266), .O(gate137inter3));
  inv1  gate2413(.a(s_267), .O(gate137inter4));
  nand2 gate2414(.a(gate137inter4), .b(gate137inter3), .O(gate137inter5));
  nor2  gate2415(.a(gate137inter5), .b(gate137inter2), .O(gate137inter6));
  inv1  gate2416(.a(G426), .O(gate137inter7));
  inv1  gate2417(.a(G429), .O(gate137inter8));
  nand2 gate2418(.a(gate137inter8), .b(gate137inter7), .O(gate137inter9));
  nand2 gate2419(.a(s_267), .b(gate137inter3), .O(gate137inter10));
  nor2  gate2420(.a(gate137inter10), .b(gate137inter9), .O(gate137inter11));
  nor2  gate2421(.a(gate137inter11), .b(gate137inter6), .O(gate137inter12));
  nand2 gate2422(.a(gate137inter12), .b(gate137inter1), .O(G522));
nand2 gate138( .a(G432), .b(G435), .O(G525) );

  xor2  gate841(.a(G441), .b(G438), .O(gate139inter0));
  nand2 gate842(.a(gate139inter0), .b(s_42), .O(gate139inter1));
  and2  gate843(.a(G441), .b(G438), .O(gate139inter2));
  inv1  gate844(.a(s_42), .O(gate139inter3));
  inv1  gate845(.a(s_43), .O(gate139inter4));
  nand2 gate846(.a(gate139inter4), .b(gate139inter3), .O(gate139inter5));
  nor2  gate847(.a(gate139inter5), .b(gate139inter2), .O(gate139inter6));
  inv1  gate848(.a(G438), .O(gate139inter7));
  inv1  gate849(.a(G441), .O(gate139inter8));
  nand2 gate850(.a(gate139inter8), .b(gate139inter7), .O(gate139inter9));
  nand2 gate851(.a(s_43), .b(gate139inter3), .O(gate139inter10));
  nor2  gate852(.a(gate139inter10), .b(gate139inter9), .O(gate139inter11));
  nor2  gate853(.a(gate139inter11), .b(gate139inter6), .O(gate139inter12));
  nand2 gate854(.a(gate139inter12), .b(gate139inter1), .O(G528));

  xor2  gate1849(.a(G447), .b(G444), .O(gate140inter0));
  nand2 gate1850(.a(gate140inter0), .b(s_186), .O(gate140inter1));
  and2  gate1851(.a(G447), .b(G444), .O(gate140inter2));
  inv1  gate1852(.a(s_186), .O(gate140inter3));
  inv1  gate1853(.a(s_187), .O(gate140inter4));
  nand2 gate1854(.a(gate140inter4), .b(gate140inter3), .O(gate140inter5));
  nor2  gate1855(.a(gate140inter5), .b(gate140inter2), .O(gate140inter6));
  inv1  gate1856(.a(G444), .O(gate140inter7));
  inv1  gate1857(.a(G447), .O(gate140inter8));
  nand2 gate1858(.a(gate140inter8), .b(gate140inter7), .O(gate140inter9));
  nand2 gate1859(.a(s_187), .b(gate140inter3), .O(gate140inter10));
  nor2  gate1860(.a(gate140inter10), .b(gate140inter9), .O(gate140inter11));
  nor2  gate1861(.a(gate140inter11), .b(gate140inter6), .O(gate140inter12));
  nand2 gate1862(.a(gate140inter12), .b(gate140inter1), .O(G531));
nand2 gate141( .a(G450), .b(G453), .O(G534) );
nand2 gate142( .a(G456), .b(G459), .O(G537) );
nand2 gate143( .a(G462), .b(G465), .O(G540) );

  xor2  gate2423(.a(G471), .b(G468), .O(gate144inter0));
  nand2 gate2424(.a(gate144inter0), .b(s_268), .O(gate144inter1));
  and2  gate2425(.a(G471), .b(G468), .O(gate144inter2));
  inv1  gate2426(.a(s_268), .O(gate144inter3));
  inv1  gate2427(.a(s_269), .O(gate144inter4));
  nand2 gate2428(.a(gate144inter4), .b(gate144inter3), .O(gate144inter5));
  nor2  gate2429(.a(gate144inter5), .b(gate144inter2), .O(gate144inter6));
  inv1  gate2430(.a(G468), .O(gate144inter7));
  inv1  gate2431(.a(G471), .O(gate144inter8));
  nand2 gate2432(.a(gate144inter8), .b(gate144inter7), .O(gate144inter9));
  nand2 gate2433(.a(s_269), .b(gate144inter3), .O(gate144inter10));
  nor2  gate2434(.a(gate144inter10), .b(gate144inter9), .O(gate144inter11));
  nor2  gate2435(.a(gate144inter11), .b(gate144inter6), .O(gate144inter12));
  nand2 gate2436(.a(gate144inter12), .b(gate144inter1), .O(G543));

  xor2  gate1121(.a(G477), .b(G474), .O(gate145inter0));
  nand2 gate1122(.a(gate145inter0), .b(s_82), .O(gate145inter1));
  and2  gate1123(.a(G477), .b(G474), .O(gate145inter2));
  inv1  gate1124(.a(s_82), .O(gate145inter3));
  inv1  gate1125(.a(s_83), .O(gate145inter4));
  nand2 gate1126(.a(gate145inter4), .b(gate145inter3), .O(gate145inter5));
  nor2  gate1127(.a(gate145inter5), .b(gate145inter2), .O(gate145inter6));
  inv1  gate1128(.a(G474), .O(gate145inter7));
  inv1  gate1129(.a(G477), .O(gate145inter8));
  nand2 gate1130(.a(gate145inter8), .b(gate145inter7), .O(gate145inter9));
  nand2 gate1131(.a(s_83), .b(gate145inter3), .O(gate145inter10));
  nor2  gate1132(.a(gate145inter10), .b(gate145inter9), .O(gate145inter11));
  nor2  gate1133(.a(gate145inter11), .b(gate145inter6), .O(gate145inter12));
  nand2 gate1134(.a(gate145inter12), .b(gate145inter1), .O(G546));
nand2 gate146( .a(G480), .b(G483), .O(G549) );
nand2 gate147( .a(G486), .b(G489), .O(G552) );

  xor2  gate1401(.a(G495), .b(G492), .O(gate148inter0));
  nand2 gate1402(.a(gate148inter0), .b(s_122), .O(gate148inter1));
  and2  gate1403(.a(G495), .b(G492), .O(gate148inter2));
  inv1  gate1404(.a(s_122), .O(gate148inter3));
  inv1  gate1405(.a(s_123), .O(gate148inter4));
  nand2 gate1406(.a(gate148inter4), .b(gate148inter3), .O(gate148inter5));
  nor2  gate1407(.a(gate148inter5), .b(gate148inter2), .O(gate148inter6));
  inv1  gate1408(.a(G492), .O(gate148inter7));
  inv1  gate1409(.a(G495), .O(gate148inter8));
  nand2 gate1410(.a(gate148inter8), .b(gate148inter7), .O(gate148inter9));
  nand2 gate1411(.a(s_123), .b(gate148inter3), .O(gate148inter10));
  nor2  gate1412(.a(gate148inter10), .b(gate148inter9), .O(gate148inter11));
  nor2  gate1413(.a(gate148inter11), .b(gate148inter6), .O(gate148inter12));
  nand2 gate1414(.a(gate148inter12), .b(gate148inter1), .O(G555));
nand2 gate149( .a(G498), .b(G501), .O(G558) );
nand2 gate150( .a(G504), .b(G507), .O(G561) );

  xor2  gate2465(.a(G513), .b(G510), .O(gate151inter0));
  nand2 gate2466(.a(gate151inter0), .b(s_274), .O(gate151inter1));
  and2  gate2467(.a(G513), .b(G510), .O(gate151inter2));
  inv1  gate2468(.a(s_274), .O(gate151inter3));
  inv1  gate2469(.a(s_275), .O(gate151inter4));
  nand2 gate2470(.a(gate151inter4), .b(gate151inter3), .O(gate151inter5));
  nor2  gate2471(.a(gate151inter5), .b(gate151inter2), .O(gate151inter6));
  inv1  gate2472(.a(G510), .O(gate151inter7));
  inv1  gate2473(.a(G513), .O(gate151inter8));
  nand2 gate2474(.a(gate151inter8), .b(gate151inter7), .O(gate151inter9));
  nand2 gate2475(.a(s_275), .b(gate151inter3), .O(gate151inter10));
  nor2  gate2476(.a(gate151inter10), .b(gate151inter9), .O(gate151inter11));
  nor2  gate2477(.a(gate151inter11), .b(gate151inter6), .O(gate151inter12));
  nand2 gate2478(.a(gate151inter12), .b(gate151inter1), .O(G564));

  xor2  gate1205(.a(G519), .b(G516), .O(gate152inter0));
  nand2 gate1206(.a(gate152inter0), .b(s_94), .O(gate152inter1));
  and2  gate1207(.a(G519), .b(G516), .O(gate152inter2));
  inv1  gate1208(.a(s_94), .O(gate152inter3));
  inv1  gate1209(.a(s_95), .O(gate152inter4));
  nand2 gate1210(.a(gate152inter4), .b(gate152inter3), .O(gate152inter5));
  nor2  gate1211(.a(gate152inter5), .b(gate152inter2), .O(gate152inter6));
  inv1  gate1212(.a(G516), .O(gate152inter7));
  inv1  gate1213(.a(G519), .O(gate152inter8));
  nand2 gate1214(.a(gate152inter8), .b(gate152inter7), .O(gate152inter9));
  nand2 gate1215(.a(s_95), .b(gate152inter3), .O(gate152inter10));
  nor2  gate1216(.a(gate152inter10), .b(gate152inter9), .O(gate152inter11));
  nor2  gate1217(.a(gate152inter11), .b(gate152inter6), .O(gate152inter12));
  nand2 gate1218(.a(gate152inter12), .b(gate152inter1), .O(G567));

  xor2  gate1429(.a(G522), .b(G426), .O(gate153inter0));
  nand2 gate1430(.a(gate153inter0), .b(s_126), .O(gate153inter1));
  and2  gate1431(.a(G522), .b(G426), .O(gate153inter2));
  inv1  gate1432(.a(s_126), .O(gate153inter3));
  inv1  gate1433(.a(s_127), .O(gate153inter4));
  nand2 gate1434(.a(gate153inter4), .b(gate153inter3), .O(gate153inter5));
  nor2  gate1435(.a(gate153inter5), .b(gate153inter2), .O(gate153inter6));
  inv1  gate1436(.a(G426), .O(gate153inter7));
  inv1  gate1437(.a(G522), .O(gate153inter8));
  nand2 gate1438(.a(gate153inter8), .b(gate153inter7), .O(gate153inter9));
  nand2 gate1439(.a(s_127), .b(gate153inter3), .O(gate153inter10));
  nor2  gate1440(.a(gate153inter10), .b(gate153inter9), .O(gate153inter11));
  nor2  gate1441(.a(gate153inter11), .b(gate153inter6), .O(gate153inter12));
  nand2 gate1442(.a(gate153inter12), .b(gate153inter1), .O(G570));

  xor2  gate2227(.a(G522), .b(G429), .O(gate154inter0));
  nand2 gate2228(.a(gate154inter0), .b(s_240), .O(gate154inter1));
  and2  gate2229(.a(G522), .b(G429), .O(gate154inter2));
  inv1  gate2230(.a(s_240), .O(gate154inter3));
  inv1  gate2231(.a(s_241), .O(gate154inter4));
  nand2 gate2232(.a(gate154inter4), .b(gate154inter3), .O(gate154inter5));
  nor2  gate2233(.a(gate154inter5), .b(gate154inter2), .O(gate154inter6));
  inv1  gate2234(.a(G429), .O(gate154inter7));
  inv1  gate2235(.a(G522), .O(gate154inter8));
  nand2 gate2236(.a(gate154inter8), .b(gate154inter7), .O(gate154inter9));
  nand2 gate2237(.a(s_241), .b(gate154inter3), .O(gate154inter10));
  nor2  gate2238(.a(gate154inter10), .b(gate154inter9), .O(gate154inter11));
  nor2  gate2239(.a(gate154inter11), .b(gate154inter6), .O(gate154inter12));
  nand2 gate2240(.a(gate154inter12), .b(gate154inter1), .O(G571));

  xor2  gate2395(.a(G525), .b(G432), .O(gate155inter0));
  nand2 gate2396(.a(gate155inter0), .b(s_264), .O(gate155inter1));
  and2  gate2397(.a(G525), .b(G432), .O(gate155inter2));
  inv1  gate2398(.a(s_264), .O(gate155inter3));
  inv1  gate2399(.a(s_265), .O(gate155inter4));
  nand2 gate2400(.a(gate155inter4), .b(gate155inter3), .O(gate155inter5));
  nor2  gate2401(.a(gate155inter5), .b(gate155inter2), .O(gate155inter6));
  inv1  gate2402(.a(G432), .O(gate155inter7));
  inv1  gate2403(.a(G525), .O(gate155inter8));
  nand2 gate2404(.a(gate155inter8), .b(gate155inter7), .O(gate155inter9));
  nand2 gate2405(.a(s_265), .b(gate155inter3), .O(gate155inter10));
  nor2  gate2406(.a(gate155inter10), .b(gate155inter9), .O(gate155inter11));
  nor2  gate2407(.a(gate155inter11), .b(gate155inter6), .O(gate155inter12));
  nand2 gate2408(.a(gate155inter12), .b(gate155inter1), .O(G572));
nand2 gate156( .a(G435), .b(G525), .O(G573) );
nand2 gate157( .a(G438), .b(G528), .O(G574) );
nand2 gate158( .a(G441), .b(G528), .O(G575) );
nand2 gate159( .a(G444), .b(G531), .O(G576) );
nand2 gate160( .a(G447), .b(G531), .O(G577) );

  xor2  gate1569(.a(G534), .b(G450), .O(gate161inter0));
  nand2 gate1570(.a(gate161inter0), .b(s_146), .O(gate161inter1));
  and2  gate1571(.a(G534), .b(G450), .O(gate161inter2));
  inv1  gate1572(.a(s_146), .O(gate161inter3));
  inv1  gate1573(.a(s_147), .O(gate161inter4));
  nand2 gate1574(.a(gate161inter4), .b(gate161inter3), .O(gate161inter5));
  nor2  gate1575(.a(gate161inter5), .b(gate161inter2), .O(gate161inter6));
  inv1  gate1576(.a(G450), .O(gate161inter7));
  inv1  gate1577(.a(G534), .O(gate161inter8));
  nand2 gate1578(.a(gate161inter8), .b(gate161inter7), .O(gate161inter9));
  nand2 gate1579(.a(s_147), .b(gate161inter3), .O(gate161inter10));
  nor2  gate1580(.a(gate161inter10), .b(gate161inter9), .O(gate161inter11));
  nor2  gate1581(.a(gate161inter11), .b(gate161inter6), .O(gate161inter12));
  nand2 gate1582(.a(gate161inter12), .b(gate161inter1), .O(G578));
nand2 gate162( .a(G453), .b(G534), .O(G579) );
nand2 gate163( .a(G456), .b(G537), .O(G580) );

  xor2  gate1737(.a(G537), .b(G459), .O(gate164inter0));
  nand2 gate1738(.a(gate164inter0), .b(s_170), .O(gate164inter1));
  and2  gate1739(.a(G537), .b(G459), .O(gate164inter2));
  inv1  gate1740(.a(s_170), .O(gate164inter3));
  inv1  gate1741(.a(s_171), .O(gate164inter4));
  nand2 gate1742(.a(gate164inter4), .b(gate164inter3), .O(gate164inter5));
  nor2  gate1743(.a(gate164inter5), .b(gate164inter2), .O(gate164inter6));
  inv1  gate1744(.a(G459), .O(gate164inter7));
  inv1  gate1745(.a(G537), .O(gate164inter8));
  nand2 gate1746(.a(gate164inter8), .b(gate164inter7), .O(gate164inter9));
  nand2 gate1747(.a(s_171), .b(gate164inter3), .O(gate164inter10));
  nor2  gate1748(.a(gate164inter10), .b(gate164inter9), .O(gate164inter11));
  nor2  gate1749(.a(gate164inter11), .b(gate164inter6), .O(gate164inter12));
  nand2 gate1750(.a(gate164inter12), .b(gate164inter1), .O(G581));
nand2 gate165( .a(G462), .b(G540), .O(G582) );

  xor2  gate2059(.a(G540), .b(G465), .O(gate166inter0));
  nand2 gate2060(.a(gate166inter0), .b(s_216), .O(gate166inter1));
  and2  gate2061(.a(G540), .b(G465), .O(gate166inter2));
  inv1  gate2062(.a(s_216), .O(gate166inter3));
  inv1  gate2063(.a(s_217), .O(gate166inter4));
  nand2 gate2064(.a(gate166inter4), .b(gate166inter3), .O(gate166inter5));
  nor2  gate2065(.a(gate166inter5), .b(gate166inter2), .O(gate166inter6));
  inv1  gate2066(.a(G465), .O(gate166inter7));
  inv1  gate2067(.a(G540), .O(gate166inter8));
  nand2 gate2068(.a(gate166inter8), .b(gate166inter7), .O(gate166inter9));
  nand2 gate2069(.a(s_217), .b(gate166inter3), .O(gate166inter10));
  nor2  gate2070(.a(gate166inter10), .b(gate166inter9), .O(gate166inter11));
  nor2  gate2071(.a(gate166inter11), .b(gate166inter6), .O(gate166inter12));
  nand2 gate2072(.a(gate166inter12), .b(gate166inter1), .O(G583));
nand2 gate167( .a(G468), .b(G543), .O(G584) );
nand2 gate168( .a(G471), .b(G543), .O(G585) );
nand2 gate169( .a(G474), .b(G546), .O(G586) );

  xor2  gate1247(.a(G546), .b(G477), .O(gate170inter0));
  nand2 gate1248(.a(gate170inter0), .b(s_100), .O(gate170inter1));
  and2  gate1249(.a(G546), .b(G477), .O(gate170inter2));
  inv1  gate1250(.a(s_100), .O(gate170inter3));
  inv1  gate1251(.a(s_101), .O(gate170inter4));
  nand2 gate1252(.a(gate170inter4), .b(gate170inter3), .O(gate170inter5));
  nor2  gate1253(.a(gate170inter5), .b(gate170inter2), .O(gate170inter6));
  inv1  gate1254(.a(G477), .O(gate170inter7));
  inv1  gate1255(.a(G546), .O(gate170inter8));
  nand2 gate1256(.a(gate170inter8), .b(gate170inter7), .O(gate170inter9));
  nand2 gate1257(.a(s_101), .b(gate170inter3), .O(gate170inter10));
  nor2  gate1258(.a(gate170inter10), .b(gate170inter9), .O(gate170inter11));
  nor2  gate1259(.a(gate170inter11), .b(gate170inter6), .O(gate170inter12));
  nand2 gate1260(.a(gate170inter12), .b(gate170inter1), .O(G587));

  xor2  gate1261(.a(G549), .b(G480), .O(gate171inter0));
  nand2 gate1262(.a(gate171inter0), .b(s_102), .O(gate171inter1));
  and2  gate1263(.a(G549), .b(G480), .O(gate171inter2));
  inv1  gate1264(.a(s_102), .O(gate171inter3));
  inv1  gate1265(.a(s_103), .O(gate171inter4));
  nand2 gate1266(.a(gate171inter4), .b(gate171inter3), .O(gate171inter5));
  nor2  gate1267(.a(gate171inter5), .b(gate171inter2), .O(gate171inter6));
  inv1  gate1268(.a(G480), .O(gate171inter7));
  inv1  gate1269(.a(G549), .O(gate171inter8));
  nand2 gate1270(.a(gate171inter8), .b(gate171inter7), .O(gate171inter9));
  nand2 gate1271(.a(s_103), .b(gate171inter3), .O(gate171inter10));
  nor2  gate1272(.a(gate171inter10), .b(gate171inter9), .O(gate171inter11));
  nor2  gate1273(.a(gate171inter11), .b(gate171inter6), .O(gate171inter12));
  nand2 gate1274(.a(gate171inter12), .b(gate171inter1), .O(G588));
nand2 gate172( .a(G483), .b(G549), .O(G589) );
nand2 gate173( .a(G486), .b(G552), .O(G590) );

  xor2  gate827(.a(G552), .b(G489), .O(gate174inter0));
  nand2 gate828(.a(gate174inter0), .b(s_40), .O(gate174inter1));
  and2  gate829(.a(G552), .b(G489), .O(gate174inter2));
  inv1  gate830(.a(s_40), .O(gate174inter3));
  inv1  gate831(.a(s_41), .O(gate174inter4));
  nand2 gate832(.a(gate174inter4), .b(gate174inter3), .O(gate174inter5));
  nor2  gate833(.a(gate174inter5), .b(gate174inter2), .O(gate174inter6));
  inv1  gate834(.a(G489), .O(gate174inter7));
  inv1  gate835(.a(G552), .O(gate174inter8));
  nand2 gate836(.a(gate174inter8), .b(gate174inter7), .O(gate174inter9));
  nand2 gate837(.a(s_41), .b(gate174inter3), .O(gate174inter10));
  nor2  gate838(.a(gate174inter10), .b(gate174inter9), .O(gate174inter11));
  nor2  gate839(.a(gate174inter11), .b(gate174inter6), .O(gate174inter12));
  nand2 gate840(.a(gate174inter12), .b(gate174inter1), .O(G591));

  xor2  gate2773(.a(G555), .b(G492), .O(gate175inter0));
  nand2 gate2774(.a(gate175inter0), .b(s_318), .O(gate175inter1));
  and2  gate2775(.a(G555), .b(G492), .O(gate175inter2));
  inv1  gate2776(.a(s_318), .O(gate175inter3));
  inv1  gate2777(.a(s_319), .O(gate175inter4));
  nand2 gate2778(.a(gate175inter4), .b(gate175inter3), .O(gate175inter5));
  nor2  gate2779(.a(gate175inter5), .b(gate175inter2), .O(gate175inter6));
  inv1  gate2780(.a(G492), .O(gate175inter7));
  inv1  gate2781(.a(G555), .O(gate175inter8));
  nand2 gate2782(.a(gate175inter8), .b(gate175inter7), .O(gate175inter9));
  nand2 gate2783(.a(s_319), .b(gate175inter3), .O(gate175inter10));
  nor2  gate2784(.a(gate175inter10), .b(gate175inter9), .O(gate175inter11));
  nor2  gate2785(.a(gate175inter11), .b(gate175inter6), .O(gate175inter12));
  nand2 gate2786(.a(gate175inter12), .b(gate175inter1), .O(G592));
nand2 gate176( .a(G495), .b(G555), .O(G593) );
nand2 gate177( .a(G498), .b(G558), .O(G594) );
nand2 gate178( .a(G501), .b(G558), .O(G595) );
nand2 gate179( .a(G504), .b(G561), .O(G596) );
nand2 gate180( .a(G507), .b(G561), .O(G597) );
nand2 gate181( .a(G510), .b(G564), .O(G598) );
nand2 gate182( .a(G513), .b(G564), .O(G599) );
nand2 gate183( .a(G516), .b(G567), .O(G600) );

  xor2  gate1821(.a(G567), .b(G519), .O(gate184inter0));
  nand2 gate1822(.a(gate184inter0), .b(s_182), .O(gate184inter1));
  and2  gate1823(.a(G567), .b(G519), .O(gate184inter2));
  inv1  gate1824(.a(s_182), .O(gate184inter3));
  inv1  gate1825(.a(s_183), .O(gate184inter4));
  nand2 gate1826(.a(gate184inter4), .b(gate184inter3), .O(gate184inter5));
  nor2  gate1827(.a(gate184inter5), .b(gate184inter2), .O(gate184inter6));
  inv1  gate1828(.a(G519), .O(gate184inter7));
  inv1  gate1829(.a(G567), .O(gate184inter8));
  nand2 gate1830(.a(gate184inter8), .b(gate184inter7), .O(gate184inter9));
  nand2 gate1831(.a(s_183), .b(gate184inter3), .O(gate184inter10));
  nor2  gate1832(.a(gate184inter10), .b(gate184inter9), .O(gate184inter11));
  nor2  gate1833(.a(gate184inter11), .b(gate184inter6), .O(gate184inter12));
  nand2 gate1834(.a(gate184inter12), .b(gate184inter1), .O(G601));
nand2 gate185( .a(G570), .b(G571), .O(G602) );
nand2 gate186( .a(G572), .b(G573), .O(G607) );
nand2 gate187( .a(G574), .b(G575), .O(G612) );

  xor2  gate2017(.a(G577), .b(G576), .O(gate188inter0));
  nand2 gate2018(.a(gate188inter0), .b(s_210), .O(gate188inter1));
  and2  gate2019(.a(G577), .b(G576), .O(gate188inter2));
  inv1  gate2020(.a(s_210), .O(gate188inter3));
  inv1  gate2021(.a(s_211), .O(gate188inter4));
  nand2 gate2022(.a(gate188inter4), .b(gate188inter3), .O(gate188inter5));
  nor2  gate2023(.a(gate188inter5), .b(gate188inter2), .O(gate188inter6));
  inv1  gate2024(.a(G576), .O(gate188inter7));
  inv1  gate2025(.a(G577), .O(gate188inter8));
  nand2 gate2026(.a(gate188inter8), .b(gate188inter7), .O(gate188inter9));
  nand2 gate2027(.a(s_211), .b(gate188inter3), .O(gate188inter10));
  nor2  gate2028(.a(gate188inter10), .b(gate188inter9), .O(gate188inter11));
  nor2  gate2029(.a(gate188inter11), .b(gate188inter6), .O(gate188inter12));
  nand2 gate2030(.a(gate188inter12), .b(gate188inter1), .O(G617));
nand2 gate189( .a(G578), .b(G579), .O(G622) );
nand2 gate190( .a(G580), .b(G581), .O(G627) );

  xor2  gate1877(.a(G583), .b(G582), .O(gate191inter0));
  nand2 gate1878(.a(gate191inter0), .b(s_190), .O(gate191inter1));
  and2  gate1879(.a(G583), .b(G582), .O(gate191inter2));
  inv1  gate1880(.a(s_190), .O(gate191inter3));
  inv1  gate1881(.a(s_191), .O(gate191inter4));
  nand2 gate1882(.a(gate191inter4), .b(gate191inter3), .O(gate191inter5));
  nor2  gate1883(.a(gate191inter5), .b(gate191inter2), .O(gate191inter6));
  inv1  gate1884(.a(G582), .O(gate191inter7));
  inv1  gate1885(.a(G583), .O(gate191inter8));
  nand2 gate1886(.a(gate191inter8), .b(gate191inter7), .O(gate191inter9));
  nand2 gate1887(.a(s_191), .b(gate191inter3), .O(gate191inter10));
  nor2  gate1888(.a(gate191inter10), .b(gate191inter9), .O(gate191inter11));
  nor2  gate1889(.a(gate191inter11), .b(gate191inter6), .O(gate191inter12));
  nand2 gate1890(.a(gate191inter12), .b(gate191inter1), .O(G632));
nand2 gate192( .a(G584), .b(G585), .O(G637) );

  xor2  gate939(.a(G587), .b(G586), .O(gate193inter0));
  nand2 gate940(.a(gate193inter0), .b(s_56), .O(gate193inter1));
  and2  gate941(.a(G587), .b(G586), .O(gate193inter2));
  inv1  gate942(.a(s_56), .O(gate193inter3));
  inv1  gate943(.a(s_57), .O(gate193inter4));
  nand2 gate944(.a(gate193inter4), .b(gate193inter3), .O(gate193inter5));
  nor2  gate945(.a(gate193inter5), .b(gate193inter2), .O(gate193inter6));
  inv1  gate946(.a(G586), .O(gate193inter7));
  inv1  gate947(.a(G587), .O(gate193inter8));
  nand2 gate948(.a(gate193inter8), .b(gate193inter7), .O(gate193inter9));
  nand2 gate949(.a(s_57), .b(gate193inter3), .O(gate193inter10));
  nor2  gate950(.a(gate193inter10), .b(gate193inter9), .O(gate193inter11));
  nor2  gate951(.a(gate193inter11), .b(gate193inter6), .O(gate193inter12));
  nand2 gate952(.a(gate193inter12), .b(gate193inter1), .O(G642));

  xor2  gate1359(.a(G589), .b(G588), .O(gate194inter0));
  nand2 gate1360(.a(gate194inter0), .b(s_116), .O(gate194inter1));
  and2  gate1361(.a(G589), .b(G588), .O(gate194inter2));
  inv1  gate1362(.a(s_116), .O(gate194inter3));
  inv1  gate1363(.a(s_117), .O(gate194inter4));
  nand2 gate1364(.a(gate194inter4), .b(gate194inter3), .O(gate194inter5));
  nor2  gate1365(.a(gate194inter5), .b(gate194inter2), .O(gate194inter6));
  inv1  gate1366(.a(G588), .O(gate194inter7));
  inv1  gate1367(.a(G589), .O(gate194inter8));
  nand2 gate1368(.a(gate194inter8), .b(gate194inter7), .O(gate194inter9));
  nand2 gate1369(.a(s_117), .b(gate194inter3), .O(gate194inter10));
  nor2  gate1370(.a(gate194inter10), .b(gate194inter9), .O(gate194inter11));
  nor2  gate1371(.a(gate194inter11), .b(gate194inter6), .O(gate194inter12));
  nand2 gate1372(.a(gate194inter12), .b(gate194inter1), .O(G645));

  xor2  gate687(.a(G591), .b(G590), .O(gate195inter0));
  nand2 gate688(.a(gate195inter0), .b(s_20), .O(gate195inter1));
  and2  gate689(.a(G591), .b(G590), .O(gate195inter2));
  inv1  gate690(.a(s_20), .O(gate195inter3));
  inv1  gate691(.a(s_21), .O(gate195inter4));
  nand2 gate692(.a(gate195inter4), .b(gate195inter3), .O(gate195inter5));
  nor2  gate693(.a(gate195inter5), .b(gate195inter2), .O(gate195inter6));
  inv1  gate694(.a(G590), .O(gate195inter7));
  inv1  gate695(.a(G591), .O(gate195inter8));
  nand2 gate696(.a(gate195inter8), .b(gate195inter7), .O(gate195inter9));
  nand2 gate697(.a(s_21), .b(gate195inter3), .O(gate195inter10));
  nor2  gate698(.a(gate195inter10), .b(gate195inter9), .O(gate195inter11));
  nor2  gate699(.a(gate195inter11), .b(gate195inter6), .O(gate195inter12));
  nand2 gate700(.a(gate195inter12), .b(gate195inter1), .O(G648));

  xor2  gate1191(.a(G593), .b(G592), .O(gate196inter0));
  nand2 gate1192(.a(gate196inter0), .b(s_92), .O(gate196inter1));
  and2  gate1193(.a(G593), .b(G592), .O(gate196inter2));
  inv1  gate1194(.a(s_92), .O(gate196inter3));
  inv1  gate1195(.a(s_93), .O(gate196inter4));
  nand2 gate1196(.a(gate196inter4), .b(gate196inter3), .O(gate196inter5));
  nor2  gate1197(.a(gate196inter5), .b(gate196inter2), .O(gate196inter6));
  inv1  gate1198(.a(G592), .O(gate196inter7));
  inv1  gate1199(.a(G593), .O(gate196inter8));
  nand2 gate1200(.a(gate196inter8), .b(gate196inter7), .O(gate196inter9));
  nand2 gate1201(.a(s_93), .b(gate196inter3), .O(gate196inter10));
  nor2  gate1202(.a(gate196inter10), .b(gate196inter9), .O(gate196inter11));
  nor2  gate1203(.a(gate196inter11), .b(gate196inter6), .O(gate196inter12));
  nand2 gate1204(.a(gate196inter12), .b(gate196inter1), .O(G651));
nand2 gate197( .a(G594), .b(G595), .O(G654) );

  xor2  gate729(.a(G597), .b(G596), .O(gate198inter0));
  nand2 gate730(.a(gate198inter0), .b(s_26), .O(gate198inter1));
  and2  gate731(.a(G597), .b(G596), .O(gate198inter2));
  inv1  gate732(.a(s_26), .O(gate198inter3));
  inv1  gate733(.a(s_27), .O(gate198inter4));
  nand2 gate734(.a(gate198inter4), .b(gate198inter3), .O(gate198inter5));
  nor2  gate735(.a(gate198inter5), .b(gate198inter2), .O(gate198inter6));
  inv1  gate736(.a(G596), .O(gate198inter7));
  inv1  gate737(.a(G597), .O(gate198inter8));
  nand2 gate738(.a(gate198inter8), .b(gate198inter7), .O(gate198inter9));
  nand2 gate739(.a(s_27), .b(gate198inter3), .O(gate198inter10));
  nor2  gate740(.a(gate198inter10), .b(gate198inter9), .O(gate198inter11));
  nor2  gate741(.a(gate198inter11), .b(gate198inter6), .O(gate198inter12));
  nand2 gate742(.a(gate198inter12), .b(gate198inter1), .O(G657));

  xor2  gate2157(.a(G599), .b(G598), .O(gate199inter0));
  nand2 gate2158(.a(gate199inter0), .b(s_230), .O(gate199inter1));
  and2  gate2159(.a(G599), .b(G598), .O(gate199inter2));
  inv1  gate2160(.a(s_230), .O(gate199inter3));
  inv1  gate2161(.a(s_231), .O(gate199inter4));
  nand2 gate2162(.a(gate199inter4), .b(gate199inter3), .O(gate199inter5));
  nor2  gate2163(.a(gate199inter5), .b(gate199inter2), .O(gate199inter6));
  inv1  gate2164(.a(G598), .O(gate199inter7));
  inv1  gate2165(.a(G599), .O(gate199inter8));
  nand2 gate2166(.a(gate199inter8), .b(gate199inter7), .O(gate199inter9));
  nand2 gate2167(.a(s_231), .b(gate199inter3), .O(gate199inter10));
  nor2  gate2168(.a(gate199inter10), .b(gate199inter9), .O(gate199inter11));
  nor2  gate2169(.a(gate199inter11), .b(gate199inter6), .O(gate199inter12));
  nand2 gate2170(.a(gate199inter12), .b(gate199inter1), .O(G660));
nand2 gate200( .a(G600), .b(G601), .O(G663) );
nand2 gate201( .a(G602), .b(G607), .O(G666) );

  xor2  gate2675(.a(G617), .b(G612), .O(gate202inter0));
  nand2 gate2676(.a(gate202inter0), .b(s_304), .O(gate202inter1));
  and2  gate2677(.a(G617), .b(G612), .O(gate202inter2));
  inv1  gate2678(.a(s_304), .O(gate202inter3));
  inv1  gate2679(.a(s_305), .O(gate202inter4));
  nand2 gate2680(.a(gate202inter4), .b(gate202inter3), .O(gate202inter5));
  nor2  gate2681(.a(gate202inter5), .b(gate202inter2), .O(gate202inter6));
  inv1  gate2682(.a(G612), .O(gate202inter7));
  inv1  gate2683(.a(G617), .O(gate202inter8));
  nand2 gate2684(.a(gate202inter8), .b(gate202inter7), .O(gate202inter9));
  nand2 gate2685(.a(s_305), .b(gate202inter3), .O(gate202inter10));
  nor2  gate2686(.a(gate202inter10), .b(gate202inter9), .O(gate202inter11));
  nor2  gate2687(.a(gate202inter11), .b(gate202inter6), .O(gate202inter12));
  nand2 gate2688(.a(gate202inter12), .b(gate202inter1), .O(G669));

  xor2  gate1625(.a(G612), .b(G602), .O(gate203inter0));
  nand2 gate1626(.a(gate203inter0), .b(s_154), .O(gate203inter1));
  and2  gate1627(.a(G612), .b(G602), .O(gate203inter2));
  inv1  gate1628(.a(s_154), .O(gate203inter3));
  inv1  gate1629(.a(s_155), .O(gate203inter4));
  nand2 gate1630(.a(gate203inter4), .b(gate203inter3), .O(gate203inter5));
  nor2  gate1631(.a(gate203inter5), .b(gate203inter2), .O(gate203inter6));
  inv1  gate1632(.a(G602), .O(gate203inter7));
  inv1  gate1633(.a(G612), .O(gate203inter8));
  nand2 gate1634(.a(gate203inter8), .b(gate203inter7), .O(gate203inter9));
  nand2 gate1635(.a(s_155), .b(gate203inter3), .O(gate203inter10));
  nor2  gate1636(.a(gate203inter10), .b(gate203inter9), .O(gate203inter11));
  nor2  gate1637(.a(gate203inter11), .b(gate203inter6), .O(gate203inter12));
  nand2 gate1638(.a(gate203inter12), .b(gate203inter1), .O(G672));

  xor2  gate1471(.a(G617), .b(G607), .O(gate204inter0));
  nand2 gate1472(.a(gate204inter0), .b(s_132), .O(gate204inter1));
  and2  gate1473(.a(G617), .b(G607), .O(gate204inter2));
  inv1  gate1474(.a(s_132), .O(gate204inter3));
  inv1  gate1475(.a(s_133), .O(gate204inter4));
  nand2 gate1476(.a(gate204inter4), .b(gate204inter3), .O(gate204inter5));
  nor2  gate1477(.a(gate204inter5), .b(gate204inter2), .O(gate204inter6));
  inv1  gate1478(.a(G607), .O(gate204inter7));
  inv1  gate1479(.a(G617), .O(gate204inter8));
  nand2 gate1480(.a(gate204inter8), .b(gate204inter7), .O(gate204inter9));
  nand2 gate1481(.a(s_133), .b(gate204inter3), .O(gate204inter10));
  nor2  gate1482(.a(gate204inter10), .b(gate204inter9), .O(gate204inter11));
  nor2  gate1483(.a(gate204inter11), .b(gate204inter6), .O(gate204inter12));
  nand2 gate1484(.a(gate204inter12), .b(gate204inter1), .O(G675));

  xor2  gate1317(.a(G627), .b(G622), .O(gate205inter0));
  nand2 gate1318(.a(gate205inter0), .b(s_110), .O(gate205inter1));
  and2  gate1319(.a(G627), .b(G622), .O(gate205inter2));
  inv1  gate1320(.a(s_110), .O(gate205inter3));
  inv1  gate1321(.a(s_111), .O(gate205inter4));
  nand2 gate1322(.a(gate205inter4), .b(gate205inter3), .O(gate205inter5));
  nor2  gate1323(.a(gate205inter5), .b(gate205inter2), .O(gate205inter6));
  inv1  gate1324(.a(G622), .O(gate205inter7));
  inv1  gate1325(.a(G627), .O(gate205inter8));
  nand2 gate1326(.a(gate205inter8), .b(gate205inter7), .O(gate205inter9));
  nand2 gate1327(.a(s_111), .b(gate205inter3), .O(gate205inter10));
  nor2  gate1328(.a(gate205inter10), .b(gate205inter9), .O(gate205inter11));
  nor2  gate1329(.a(gate205inter11), .b(gate205inter6), .O(gate205inter12));
  nand2 gate1330(.a(gate205inter12), .b(gate205inter1), .O(G678));
nand2 gate206( .a(G632), .b(G637), .O(G681) );

  xor2  gate2507(.a(G632), .b(G622), .O(gate207inter0));
  nand2 gate2508(.a(gate207inter0), .b(s_280), .O(gate207inter1));
  and2  gate2509(.a(G632), .b(G622), .O(gate207inter2));
  inv1  gate2510(.a(s_280), .O(gate207inter3));
  inv1  gate2511(.a(s_281), .O(gate207inter4));
  nand2 gate2512(.a(gate207inter4), .b(gate207inter3), .O(gate207inter5));
  nor2  gate2513(.a(gate207inter5), .b(gate207inter2), .O(gate207inter6));
  inv1  gate2514(.a(G622), .O(gate207inter7));
  inv1  gate2515(.a(G632), .O(gate207inter8));
  nand2 gate2516(.a(gate207inter8), .b(gate207inter7), .O(gate207inter9));
  nand2 gate2517(.a(s_281), .b(gate207inter3), .O(gate207inter10));
  nor2  gate2518(.a(gate207inter10), .b(gate207inter9), .O(gate207inter11));
  nor2  gate2519(.a(gate207inter11), .b(gate207inter6), .O(gate207inter12));
  nand2 gate2520(.a(gate207inter12), .b(gate207inter1), .O(G684));
nand2 gate208( .a(G627), .b(G637), .O(G687) );
nand2 gate209( .a(G602), .b(G666), .O(G690) );
nand2 gate210( .a(G607), .b(G666), .O(G691) );

  xor2  gate1107(.a(G669), .b(G612), .O(gate211inter0));
  nand2 gate1108(.a(gate211inter0), .b(s_80), .O(gate211inter1));
  and2  gate1109(.a(G669), .b(G612), .O(gate211inter2));
  inv1  gate1110(.a(s_80), .O(gate211inter3));
  inv1  gate1111(.a(s_81), .O(gate211inter4));
  nand2 gate1112(.a(gate211inter4), .b(gate211inter3), .O(gate211inter5));
  nor2  gate1113(.a(gate211inter5), .b(gate211inter2), .O(gate211inter6));
  inv1  gate1114(.a(G612), .O(gate211inter7));
  inv1  gate1115(.a(G669), .O(gate211inter8));
  nand2 gate1116(.a(gate211inter8), .b(gate211inter7), .O(gate211inter9));
  nand2 gate1117(.a(s_81), .b(gate211inter3), .O(gate211inter10));
  nor2  gate1118(.a(gate211inter10), .b(gate211inter9), .O(gate211inter11));
  nor2  gate1119(.a(gate211inter11), .b(gate211inter6), .O(gate211inter12));
  nand2 gate1120(.a(gate211inter12), .b(gate211inter1), .O(G692));

  xor2  gate897(.a(G669), .b(G617), .O(gate212inter0));
  nand2 gate898(.a(gate212inter0), .b(s_50), .O(gate212inter1));
  and2  gate899(.a(G669), .b(G617), .O(gate212inter2));
  inv1  gate900(.a(s_50), .O(gate212inter3));
  inv1  gate901(.a(s_51), .O(gate212inter4));
  nand2 gate902(.a(gate212inter4), .b(gate212inter3), .O(gate212inter5));
  nor2  gate903(.a(gate212inter5), .b(gate212inter2), .O(gate212inter6));
  inv1  gate904(.a(G617), .O(gate212inter7));
  inv1  gate905(.a(G669), .O(gate212inter8));
  nand2 gate906(.a(gate212inter8), .b(gate212inter7), .O(gate212inter9));
  nand2 gate907(.a(s_51), .b(gate212inter3), .O(gate212inter10));
  nor2  gate908(.a(gate212inter10), .b(gate212inter9), .O(gate212inter11));
  nor2  gate909(.a(gate212inter11), .b(gate212inter6), .O(gate212inter12));
  nand2 gate910(.a(gate212inter12), .b(gate212inter1), .O(G693));
nand2 gate213( .a(G602), .b(G672), .O(G694) );
nand2 gate214( .a(G612), .b(G672), .O(G695) );
nand2 gate215( .a(G607), .b(G675), .O(G696) );

  xor2  gate561(.a(G675), .b(G617), .O(gate216inter0));
  nand2 gate562(.a(gate216inter0), .b(s_2), .O(gate216inter1));
  and2  gate563(.a(G675), .b(G617), .O(gate216inter2));
  inv1  gate564(.a(s_2), .O(gate216inter3));
  inv1  gate565(.a(s_3), .O(gate216inter4));
  nand2 gate566(.a(gate216inter4), .b(gate216inter3), .O(gate216inter5));
  nor2  gate567(.a(gate216inter5), .b(gate216inter2), .O(gate216inter6));
  inv1  gate568(.a(G617), .O(gate216inter7));
  inv1  gate569(.a(G675), .O(gate216inter8));
  nand2 gate570(.a(gate216inter8), .b(gate216inter7), .O(gate216inter9));
  nand2 gate571(.a(s_3), .b(gate216inter3), .O(gate216inter10));
  nor2  gate572(.a(gate216inter10), .b(gate216inter9), .O(gate216inter11));
  nor2  gate573(.a(gate216inter11), .b(gate216inter6), .O(gate216inter12));
  nand2 gate574(.a(gate216inter12), .b(gate216inter1), .O(G697));
nand2 gate217( .a(G622), .b(G678), .O(G698) );

  xor2  gate2087(.a(G678), .b(G627), .O(gate218inter0));
  nand2 gate2088(.a(gate218inter0), .b(s_220), .O(gate218inter1));
  and2  gate2089(.a(G678), .b(G627), .O(gate218inter2));
  inv1  gate2090(.a(s_220), .O(gate218inter3));
  inv1  gate2091(.a(s_221), .O(gate218inter4));
  nand2 gate2092(.a(gate218inter4), .b(gate218inter3), .O(gate218inter5));
  nor2  gate2093(.a(gate218inter5), .b(gate218inter2), .O(gate218inter6));
  inv1  gate2094(.a(G627), .O(gate218inter7));
  inv1  gate2095(.a(G678), .O(gate218inter8));
  nand2 gate2096(.a(gate218inter8), .b(gate218inter7), .O(gate218inter9));
  nand2 gate2097(.a(s_221), .b(gate218inter3), .O(gate218inter10));
  nor2  gate2098(.a(gate218inter10), .b(gate218inter9), .O(gate218inter11));
  nor2  gate2099(.a(gate218inter11), .b(gate218inter6), .O(gate218inter12));
  nand2 gate2100(.a(gate218inter12), .b(gate218inter1), .O(G699));

  xor2  gate2073(.a(G681), .b(G632), .O(gate219inter0));
  nand2 gate2074(.a(gate219inter0), .b(s_218), .O(gate219inter1));
  and2  gate2075(.a(G681), .b(G632), .O(gate219inter2));
  inv1  gate2076(.a(s_218), .O(gate219inter3));
  inv1  gate2077(.a(s_219), .O(gate219inter4));
  nand2 gate2078(.a(gate219inter4), .b(gate219inter3), .O(gate219inter5));
  nor2  gate2079(.a(gate219inter5), .b(gate219inter2), .O(gate219inter6));
  inv1  gate2080(.a(G632), .O(gate219inter7));
  inv1  gate2081(.a(G681), .O(gate219inter8));
  nand2 gate2082(.a(gate219inter8), .b(gate219inter7), .O(gate219inter9));
  nand2 gate2083(.a(s_219), .b(gate219inter3), .O(gate219inter10));
  nor2  gate2084(.a(gate219inter10), .b(gate219inter9), .O(gate219inter11));
  nor2  gate2085(.a(gate219inter11), .b(gate219inter6), .O(gate219inter12));
  nand2 gate2086(.a(gate219inter12), .b(gate219inter1), .O(G700));
nand2 gate220( .a(G637), .b(G681), .O(G701) );

  xor2  gate2717(.a(G684), .b(G622), .O(gate221inter0));
  nand2 gate2718(.a(gate221inter0), .b(s_310), .O(gate221inter1));
  and2  gate2719(.a(G684), .b(G622), .O(gate221inter2));
  inv1  gate2720(.a(s_310), .O(gate221inter3));
  inv1  gate2721(.a(s_311), .O(gate221inter4));
  nand2 gate2722(.a(gate221inter4), .b(gate221inter3), .O(gate221inter5));
  nor2  gate2723(.a(gate221inter5), .b(gate221inter2), .O(gate221inter6));
  inv1  gate2724(.a(G622), .O(gate221inter7));
  inv1  gate2725(.a(G684), .O(gate221inter8));
  nand2 gate2726(.a(gate221inter8), .b(gate221inter7), .O(gate221inter9));
  nand2 gate2727(.a(s_311), .b(gate221inter3), .O(gate221inter10));
  nor2  gate2728(.a(gate221inter10), .b(gate221inter9), .O(gate221inter11));
  nor2  gate2729(.a(gate221inter11), .b(gate221inter6), .O(gate221inter12));
  nand2 gate2730(.a(gate221inter12), .b(gate221inter1), .O(G702));

  xor2  gate1177(.a(G684), .b(G632), .O(gate222inter0));
  nand2 gate1178(.a(gate222inter0), .b(s_90), .O(gate222inter1));
  and2  gate1179(.a(G684), .b(G632), .O(gate222inter2));
  inv1  gate1180(.a(s_90), .O(gate222inter3));
  inv1  gate1181(.a(s_91), .O(gate222inter4));
  nand2 gate1182(.a(gate222inter4), .b(gate222inter3), .O(gate222inter5));
  nor2  gate1183(.a(gate222inter5), .b(gate222inter2), .O(gate222inter6));
  inv1  gate1184(.a(G632), .O(gate222inter7));
  inv1  gate1185(.a(G684), .O(gate222inter8));
  nand2 gate1186(.a(gate222inter8), .b(gate222inter7), .O(gate222inter9));
  nand2 gate1187(.a(s_91), .b(gate222inter3), .O(gate222inter10));
  nor2  gate1188(.a(gate222inter10), .b(gate222inter9), .O(gate222inter11));
  nor2  gate1189(.a(gate222inter11), .b(gate222inter6), .O(gate222inter12));
  nand2 gate1190(.a(gate222inter12), .b(gate222inter1), .O(G703));
nand2 gate223( .a(G627), .b(G687), .O(G704) );
nand2 gate224( .a(G637), .b(G687), .O(G705) );
nand2 gate225( .a(G690), .b(G691), .O(G706) );

  xor2  gate1233(.a(G693), .b(G692), .O(gate226inter0));
  nand2 gate1234(.a(gate226inter0), .b(s_98), .O(gate226inter1));
  and2  gate1235(.a(G693), .b(G692), .O(gate226inter2));
  inv1  gate1236(.a(s_98), .O(gate226inter3));
  inv1  gate1237(.a(s_99), .O(gate226inter4));
  nand2 gate1238(.a(gate226inter4), .b(gate226inter3), .O(gate226inter5));
  nor2  gate1239(.a(gate226inter5), .b(gate226inter2), .O(gate226inter6));
  inv1  gate1240(.a(G692), .O(gate226inter7));
  inv1  gate1241(.a(G693), .O(gate226inter8));
  nand2 gate1242(.a(gate226inter8), .b(gate226inter7), .O(gate226inter9));
  nand2 gate1243(.a(s_99), .b(gate226inter3), .O(gate226inter10));
  nor2  gate1244(.a(gate226inter10), .b(gate226inter9), .O(gate226inter11));
  nor2  gate1245(.a(gate226inter11), .b(gate226inter6), .O(gate226inter12));
  nand2 gate1246(.a(gate226inter12), .b(gate226inter1), .O(G709));

  xor2  gate2437(.a(G695), .b(G694), .O(gate227inter0));
  nand2 gate2438(.a(gate227inter0), .b(s_270), .O(gate227inter1));
  and2  gate2439(.a(G695), .b(G694), .O(gate227inter2));
  inv1  gate2440(.a(s_270), .O(gate227inter3));
  inv1  gate2441(.a(s_271), .O(gate227inter4));
  nand2 gate2442(.a(gate227inter4), .b(gate227inter3), .O(gate227inter5));
  nor2  gate2443(.a(gate227inter5), .b(gate227inter2), .O(gate227inter6));
  inv1  gate2444(.a(G694), .O(gate227inter7));
  inv1  gate2445(.a(G695), .O(gate227inter8));
  nand2 gate2446(.a(gate227inter8), .b(gate227inter7), .O(gate227inter9));
  nand2 gate2447(.a(s_271), .b(gate227inter3), .O(gate227inter10));
  nor2  gate2448(.a(gate227inter10), .b(gate227inter9), .O(gate227inter11));
  nor2  gate2449(.a(gate227inter11), .b(gate227inter6), .O(gate227inter12));
  nand2 gate2450(.a(gate227inter12), .b(gate227inter1), .O(G712));
nand2 gate228( .a(G696), .b(G697), .O(G715) );

  xor2  gate1611(.a(G699), .b(G698), .O(gate229inter0));
  nand2 gate1612(.a(gate229inter0), .b(s_152), .O(gate229inter1));
  and2  gate1613(.a(G699), .b(G698), .O(gate229inter2));
  inv1  gate1614(.a(s_152), .O(gate229inter3));
  inv1  gate1615(.a(s_153), .O(gate229inter4));
  nand2 gate1616(.a(gate229inter4), .b(gate229inter3), .O(gate229inter5));
  nor2  gate1617(.a(gate229inter5), .b(gate229inter2), .O(gate229inter6));
  inv1  gate1618(.a(G698), .O(gate229inter7));
  inv1  gate1619(.a(G699), .O(gate229inter8));
  nand2 gate1620(.a(gate229inter8), .b(gate229inter7), .O(gate229inter9));
  nand2 gate1621(.a(s_153), .b(gate229inter3), .O(gate229inter10));
  nor2  gate1622(.a(gate229inter10), .b(gate229inter9), .O(gate229inter11));
  nor2  gate1623(.a(gate229inter11), .b(gate229inter6), .O(gate229inter12));
  nand2 gate1624(.a(gate229inter12), .b(gate229inter1), .O(G718));

  xor2  gate2787(.a(G701), .b(G700), .O(gate230inter0));
  nand2 gate2788(.a(gate230inter0), .b(s_320), .O(gate230inter1));
  and2  gate2789(.a(G701), .b(G700), .O(gate230inter2));
  inv1  gate2790(.a(s_320), .O(gate230inter3));
  inv1  gate2791(.a(s_321), .O(gate230inter4));
  nand2 gate2792(.a(gate230inter4), .b(gate230inter3), .O(gate230inter5));
  nor2  gate2793(.a(gate230inter5), .b(gate230inter2), .O(gate230inter6));
  inv1  gate2794(.a(G700), .O(gate230inter7));
  inv1  gate2795(.a(G701), .O(gate230inter8));
  nand2 gate2796(.a(gate230inter8), .b(gate230inter7), .O(gate230inter9));
  nand2 gate2797(.a(s_321), .b(gate230inter3), .O(gate230inter10));
  nor2  gate2798(.a(gate230inter10), .b(gate230inter9), .O(gate230inter11));
  nor2  gate2799(.a(gate230inter11), .b(gate230inter6), .O(gate230inter12));
  nand2 gate2800(.a(gate230inter12), .b(gate230inter1), .O(G721));

  xor2  gate743(.a(G703), .b(G702), .O(gate231inter0));
  nand2 gate744(.a(gate231inter0), .b(s_28), .O(gate231inter1));
  and2  gate745(.a(G703), .b(G702), .O(gate231inter2));
  inv1  gate746(.a(s_28), .O(gate231inter3));
  inv1  gate747(.a(s_29), .O(gate231inter4));
  nand2 gate748(.a(gate231inter4), .b(gate231inter3), .O(gate231inter5));
  nor2  gate749(.a(gate231inter5), .b(gate231inter2), .O(gate231inter6));
  inv1  gate750(.a(G702), .O(gate231inter7));
  inv1  gate751(.a(G703), .O(gate231inter8));
  nand2 gate752(.a(gate231inter8), .b(gate231inter7), .O(gate231inter9));
  nand2 gate753(.a(s_29), .b(gate231inter3), .O(gate231inter10));
  nor2  gate754(.a(gate231inter10), .b(gate231inter9), .O(gate231inter11));
  nor2  gate755(.a(gate231inter11), .b(gate231inter6), .O(gate231inter12));
  nand2 gate756(.a(gate231inter12), .b(gate231inter1), .O(G724));

  xor2  gate1387(.a(G705), .b(G704), .O(gate232inter0));
  nand2 gate1388(.a(gate232inter0), .b(s_120), .O(gate232inter1));
  and2  gate1389(.a(G705), .b(G704), .O(gate232inter2));
  inv1  gate1390(.a(s_120), .O(gate232inter3));
  inv1  gate1391(.a(s_121), .O(gate232inter4));
  nand2 gate1392(.a(gate232inter4), .b(gate232inter3), .O(gate232inter5));
  nor2  gate1393(.a(gate232inter5), .b(gate232inter2), .O(gate232inter6));
  inv1  gate1394(.a(G704), .O(gate232inter7));
  inv1  gate1395(.a(G705), .O(gate232inter8));
  nand2 gate1396(.a(gate232inter8), .b(gate232inter7), .O(gate232inter9));
  nand2 gate1397(.a(s_121), .b(gate232inter3), .O(gate232inter10));
  nor2  gate1398(.a(gate232inter10), .b(gate232inter9), .O(gate232inter11));
  nor2  gate1399(.a(gate232inter11), .b(gate232inter6), .O(gate232inter12));
  nand2 gate1400(.a(gate232inter12), .b(gate232inter1), .O(G727));
nand2 gate233( .a(G242), .b(G718), .O(G730) );
nand2 gate234( .a(G245), .b(G721), .O(G733) );
nand2 gate235( .a(G248), .b(G724), .O(G736) );

  xor2  gate1135(.a(G727), .b(G251), .O(gate236inter0));
  nand2 gate1136(.a(gate236inter0), .b(s_84), .O(gate236inter1));
  and2  gate1137(.a(G727), .b(G251), .O(gate236inter2));
  inv1  gate1138(.a(s_84), .O(gate236inter3));
  inv1  gate1139(.a(s_85), .O(gate236inter4));
  nand2 gate1140(.a(gate236inter4), .b(gate236inter3), .O(gate236inter5));
  nor2  gate1141(.a(gate236inter5), .b(gate236inter2), .O(gate236inter6));
  inv1  gate1142(.a(G251), .O(gate236inter7));
  inv1  gate1143(.a(G727), .O(gate236inter8));
  nand2 gate1144(.a(gate236inter8), .b(gate236inter7), .O(gate236inter9));
  nand2 gate1145(.a(s_85), .b(gate236inter3), .O(gate236inter10));
  nor2  gate1146(.a(gate236inter10), .b(gate236inter9), .O(gate236inter11));
  nor2  gate1147(.a(gate236inter11), .b(gate236inter6), .O(gate236inter12));
  nand2 gate1148(.a(gate236inter12), .b(gate236inter1), .O(G739));

  xor2  gate1667(.a(G706), .b(G254), .O(gate237inter0));
  nand2 gate1668(.a(gate237inter0), .b(s_160), .O(gate237inter1));
  and2  gate1669(.a(G706), .b(G254), .O(gate237inter2));
  inv1  gate1670(.a(s_160), .O(gate237inter3));
  inv1  gate1671(.a(s_161), .O(gate237inter4));
  nand2 gate1672(.a(gate237inter4), .b(gate237inter3), .O(gate237inter5));
  nor2  gate1673(.a(gate237inter5), .b(gate237inter2), .O(gate237inter6));
  inv1  gate1674(.a(G254), .O(gate237inter7));
  inv1  gate1675(.a(G706), .O(gate237inter8));
  nand2 gate1676(.a(gate237inter8), .b(gate237inter7), .O(gate237inter9));
  nand2 gate1677(.a(s_161), .b(gate237inter3), .O(gate237inter10));
  nor2  gate1678(.a(gate237inter10), .b(gate237inter9), .O(gate237inter11));
  nor2  gate1679(.a(gate237inter11), .b(gate237inter6), .O(gate237inter12));
  nand2 gate1680(.a(gate237inter12), .b(gate237inter1), .O(G742));

  xor2  gate1597(.a(G709), .b(G257), .O(gate238inter0));
  nand2 gate1598(.a(gate238inter0), .b(s_150), .O(gate238inter1));
  and2  gate1599(.a(G709), .b(G257), .O(gate238inter2));
  inv1  gate1600(.a(s_150), .O(gate238inter3));
  inv1  gate1601(.a(s_151), .O(gate238inter4));
  nand2 gate1602(.a(gate238inter4), .b(gate238inter3), .O(gate238inter5));
  nor2  gate1603(.a(gate238inter5), .b(gate238inter2), .O(gate238inter6));
  inv1  gate1604(.a(G257), .O(gate238inter7));
  inv1  gate1605(.a(G709), .O(gate238inter8));
  nand2 gate1606(.a(gate238inter8), .b(gate238inter7), .O(gate238inter9));
  nand2 gate1607(.a(s_151), .b(gate238inter3), .O(gate238inter10));
  nor2  gate1608(.a(gate238inter10), .b(gate238inter9), .O(gate238inter11));
  nor2  gate1609(.a(gate238inter11), .b(gate238inter6), .O(gate238inter12));
  nand2 gate1610(.a(gate238inter12), .b(gate238inter1), .O(G745));
nand2 gate239( .a(G260), .b(G712), .O(G748) );

  xor2  gate2591(.a(G715), .b(G263), .O(gate240inter0));
  nand2 gate2592(.a(gate240inter0), .b(s_292), .O(gate240inter1));
  and2  gate2593(.a(G715), .b(G263), .O(gate240inter2));
  inv1  gate2594(.a(s_292), .O(gate240inter3));
  inv1  gate2595(.a(s_293), .O(gate240inter4));
  nand2 gate2596(.a(gate240inter4), .b(gate240inter3), .O(gate240inter5));
  nor2  gate2597(.a(gate240inter5), .b(gate240inter2), .O(gate240inter6));
  inv1  gate2598(.a(G263), .O(gate240inter7));
  inv1  gate2599(.a(G715), .O(gate240inter8));
  nand2 gate2600(.a(gate240inter8), .b(gate240inter7), .O(gate240inter9));
  nand2 gate2601(.a(s_293), .b(gate240inter3), .O(gate240inter10));
  nor2  gate2602(.a(gate240inter10), .b(gate240inter9), .O(gate240inter11));
  nor2  gate2603(.a(gate240inter11), .b(gate240inter6), .O(gate240inter12));
  nand2 gate2604(.a(gate240inter12), .b(gate240inter1), .O(G751));
nand2 gate241( .a(G242), .b(G730), .O(G754) );
nand2 gate242( .a(G718), .b(G730), .O(G755) );
nand2 gate243( .a(G245), .b(G733), .O(G756) );
nand2 gate244( .a(G721), .b(G733), .O(G757) );

  xor2  gate1765(.a(G736), .b(G248), .O(gate245inter0));
  nand2 gate1766(.a(gate245inter0), .b(s_174), .O(gate245inter1));
  and2  gate1767(.a(G736), .b(G248), .O(gate245inter2));
  inv1  gate1768(.a(s_174), .O(gate245inter3));
  inv1  gate1769(.a(s_175), .O(gate245inter4));
  nand2 gate1770(.a(gate245inter4), .b(gate245inter3), .O(gate245inter5));
  nor2  gate1771(.a(gate245inter5), .b(gate245inter2), .O(gate245inter6));
  inv1  gate1772(.a(G248), .O(gate245inter7));
  inv1  gate1773(.a(G736), .O(gate245inter8));
  nand2 gate1774(.a(gate245inter8), .b(gate245inter7), .O(gate245inter9));
  nand2 gate1775(.a(s_175), .b(gate245inter3), .O(gate245inter10));
  nor2  gate1776(.a(gate245inter10), .b(gate245inter9), .O(gate245inter11));
  nor2  gate1777(.a(gate245inter11), .b(gate245inter6), .O(gate245inter12));
  nand2 gate1778(.a(gate245inter12), .b(gate245inter1), .O(G758));

  xor2  gate2241(.a(G736), .b(G724), .O(gate246inter0));
  nand2 gate2242(.a(gate246inter0), .b(s_242), .O(gate246inter1));
  and2  gate2243(.a(G736), .b(G724), .O(gate246inter2));
  inv1  gate2244(.a(s_242), .O(gate246inter3));
  inv1  gate2245(.a(s_243), .O(gate246inter4));
  nand2 gate2246(.a(gate246inter4), .b(gate246inter3), .O(gate246inter5));
  nor2  gate2247(.a(gate246inter5), .b(gate246inter2), .O(gate246inter6));
  inv1  gate2248(.a(G724), .O(gate246inter7));
  inv1  gate2249(.a(G736), .O(gate246inter8));
  nand2 gate2250(.a(gate246inter8), .b(gate246inter7), .O(gate246inter9));
  nand2 gate2251(.a(s_243), .b(gate246inter3), .O(gate246inter10));
  nor2  gate2252(.a(gate246inter10), .b(gate246inter9), .O(gate246inter11));
  nor2  gate2253(.a(gate246inter11), .b(gate246inter6), .O(gate246inter12));
  nand2 gate2254(.a(gate246inter12), .b(gate246inter1), .O(G759));
nand2 gate247( .a(G251), .b(G739), .O(G760) );
nand2 gate248( .a(G727), .b(G739), .O(G761) );
nand2 gate249( .a(G254), .b(G742), .O(G762) );

  xor2  gate2535(.a(G742), .b(G706), .O(gate250inter0));
  nand2 gate2536(.a(gate250inter0), .b(s_284), .O(gate250inter1));
  and2  gate2537(.a(G742), .b(G706), .O(gate250inter2));
  inv1  gate2538(.a(s_284), .O(gate250inter3));
  inv1  gate2539(.a(s_285), .O(gate250inter4));
  nand2 gate2540(.a(gate250inter4), .b(gate250inter3), .O(gate250inter5));
  nor2  gate2541(.a(gate250inter5), .b(gate250inter2), .O(gate250inter6));
  inv1  gate2542(.a(G706), .O(gate250inter7));
  inv1  gate2543(.a(G742), .O(gate250inter8));
  nand2 gate2544(.a(gate250inter8), .b(gate250inter7), .O(gate250inter9));
  nand2 gate2545(.a(s_285), .b(gate250inter3), .O(gate250inter10));
  nor2  gate2546(.a(gate250inter10), .b(gate250inter9), .O(gate250inter11));
  nor2  gate2547(.a(gate250inter11), .b(gate250inter6), .O(gate250inter12));
  nand2 gate2548(.a(gate250inter12), .b(gate250inter1), .O(G763));
nand2 gate251( .a(G257), .b(G745), .O(G764) );
nand2 gate252( .a(G709), .b(G745), .O(G765) );
nand2 gate253( .a(G260), .b(G748), .O(G766) );
nand2 gate254( .a(G712), .b(G748), .O(G767) );

  xor2  gate1331(.a(G751), .b(G263), .O(gate255inter0));
  nand2 gate1332(.a(gate255inter0), .b(s_112), .O(gate255inter1));
  and2  gate1333(.a(G751), .b(G263), .O(gate255inter2));
  inv1  gate1334(.a(s_112), .O(gate255inter3));
  inv1  gate1335(.a(s_113), .O(gate255inter4));
  nand2 gate1336(.a(gate255inter4), .b(gate255inter3), .O(gate255inter5));
  nor2  gate1337(.a(gate255inter5), .b(gate255inter2), .O(gate255inter6));
  inv1  gate1338(.a(G263), .O(gate255inter7));
  inv1  gate1339(.a(G751), .O(gate255inter8));
  nand2 gate1340(.a(gate255inter8), .b(gate255inter7), .O(gate255inter9));
  nand2 gate1341(.a(s_113), .b(gate255inter3), .O(gate255inter10));
  nor2  gate1342(.a(gate255inter10), .b(gate255inter9), .O(gate255inter11));
  nor2  gate1343(.a(gate255inter11), .b(gate255inter6), .O(gate255inter12));
  nand2 gate1344(.a(gate255inter12), .b(gate255inter1), .O(G768));

  xor2  gate701(.a(G751), .b(G715), .O(gate256inter0));
  nand2 gate702(.a(gate256inter0), .b(s_22), .O(gate256inter1));
  and2  gate703(.a(G751), .b(G715), .O(gate256inter2));
  inv1  gate704(.a(s_22), .O(gate256inter3));
  inv1  gate705(.a(s_23), .O(gate256inter4));
  nand2 gate706(.a(gate256inter4), .b(gate256inter3), .O(gate256inter5));
  nor2  gate707(.a(gate256inter5), .b(gate256inter2), .O(gate256inter6));
  inv1  gate708(.a(G715), .O(gate256inter7));
  inv1  gate709(.a(G751), .O(gate256inter8));
  nand2 gate710(.a(gate256inter8), .b(gate256inter7), .O(gate256inter9));
  nand2 gate711(.a(s_23), .b(gate256inter3), .O(gate256inter10));
  nor2  gate712(.a(gate256inter10), .b(gate256inter9), .O(gate256inter11));
  nor2  gate713(.a(gate256inter11), .b(gate256inter6), .O(gate256inter12));
  nand2 gate714(.a(gate256inter12), .b(gate256inter1), .O(G769));

  xor2  gate1037(.a(G755), .b(G754), .O(gate257inter0));
  nand2 gate1038(.a(gate257inter0), .b(s_70), .O(gate257inter1));
  and2  gate1039(.a(G755), .b(G754), .O(gate257inter2));
  inv1  gate1040(.a(s_70), .O(gate257inter3));
  inv1  gate1041(.a(s_71), .O(gate257inter4));
  nand2 gate1042(.a(gate257inter4), .b(gate257inter3), .O(gate257inter5));
  nor2  gate1043(.a(gate257inter5), .b(gate257inter2), .O(gate257inter6));
  inv1  gate1044(.a(G754), .O(gate257inter7));
  inv1  gate1045(.a(G755), .O(gate257inter8));
  nand2 gate1046(.a(gate257inter8), .b(gate257inter7), .O(gate257inter9));
  nand2 gate1047(.a(s_71), .b(gate257inter3), .O(gate257inter10));
  nor2  gate1048(.a(gate257inter10), .b(gate257inter9), .O(gate257inter11));
  nor2  gate1049(.a(gate257inter11), .b(gate257inter6), .O(gate257inter12));
  nand2 gate1050(.a(gate257inter12), .b(gate257inter1), .O(G770));
nand2 gate258( .a(G756), .b(G757), .O(G773) );
nand2 gate259( .a(G758), .b(G759), .O(G776) );

  xor2  gate1793(.a(G761), .b(G760), .O(gate260inter0));
  nand2 gate1794(.a(gate260inter0), .b(s_178), .O(gate260inter1));
  and2  gate1795(.a(G761), .b(G760), .O(gate260inter2));
  inv1  gate1796(.a(s_178), .O(gate260inter3));
  inv1  gate1797(.a(s_179), .O(gate260inter4));
  nand2 gate1798(.a(gate260inter4), .b(gate260inter3), .O(gate260inter5));
  nor2  gate1799(.a(gate260inter5), .b(gate260inter2), .O(gate260inter6));
  inv1  gate1800(.a(G760), .O(gate260inter7));
  inv1  gate1801(.a(G761), .O(gate260inter8));
  nand2 gate1802(.a(gate260inter8), .b(gate260inter7), .O(gate260inter9));
  nand2 gate1803(.a(s_179), .b(gate260inter3), .O(gate260inter10));
  nor2  gate1804(.a(gate260inter10), .b(gate260inter9), .O(gate260inter11));
  nor2  gate1805(.a(gate260inter11), .b(gate260inter6), .O(gate260inter12));
  nand2 gate1806(.a(gate260inter12), .b(gate260inter1), .O(G779));
nand2 gate261( .a(G762), .b(G763), .O(G782) );
nand2 gate262( .a(G764), .b(G765), .O(G785) );

  xor2  gate2199(.a(G767), .b(G766), .O(gate263inter0));
  nand2 gate2200(.a(gate263inter0), .b(s_236), .O(gate263inter1));
  and2  gate2201(.a(G767), .b(G766), .O(gate263inter2));
  inv1  gate2202(.a(s_236), .O(gate263inter3));
  inv1  gate2203(.a(s_237), .O(gate263inter4));
  nand2 gate2204(.a(gate263inter4), .b(gate263inter3), .O(gate263inter5));
  nor2  gate2205(.a(gate263inter5), .b(gate263inter2), .O(gate263inter6));
  inv1  gate2206(.a(G766), .O(gate263inter7));
  inv1  gate2207(.a(G767), .O(gate263inter8));
  nand2 gate2208(.a(gate263inter8), .b(gate263inter7), .O(gate263inter9));
  nand2 gate2209(.a(s_237), .b(gate263inter3), .O(gate263inter10));
  nor2  gate2210(.a(gate263inter10), .b(gate263inter9), .O(gate263inter11));
  nor2  gate2211(.a(gate263inter11), .b(gate263inter6), .O(gate263inter12));
  nand2 gate2212(.a(gate263inter12), .b(gate263inter1), .O(G788));
nand2 gate264( .a(G768), .b(G769), .O(G791) );

  xor2  gate2003(.a(G770), .b(G642), .O(gate265inter0));
  nand2 gate2004(.a(gate265inter0), .b(s_208), .O(gate265inter1));
  and2  gate2005(.a(G770), .b(G642), .O(gate265inter2));
  inv1  gate2006(.a(s_208), .O(gate265inter3));
  inv1  gate2007(.a(s_209), .O(gate265inter4));
  nand2 gate2008(.a(gate265inter4), .b(gate265inter3), .O(gate265inter5));
  nor2  gate2009(.a(gate265inter5), .b(gate265inter2), .O(gate265inter6));
  inv1  gate2010(.a(G642), .O(gate265inter7));
  inv1  gate2011(.a(G770), .O(gate265inter8));
  nand2 gate2012(.a(gate265inter8), .b(gate265inter7), .O(gate265inter9));
  nand2 gate2013(.a(s_209), .b(gate265inter3), .O(gate265inter10));
  nor2  gate2014(.a(gate265inter10), .b(gate265inter9), .O(gate265inter11));
  nor2  gate2015(.a(gate265inter11), .b(gate265inter6), .O(gate265inter12));
  nand2 gate2016(.a(gate265inter12), .b(gate265inter1), .O(G794));

  xor2  gate1513(.a(G773), .b(G645), .O(gate266inter0));
  nand2 gate1514(.a(gate266inter0), .b(s_138), .O(gate266inter1));
  and2  gate1515(.a(G773), .b(G645), .O(gate266inter2));
  inv1  gate1516(.a(s_138), .O(gate266inter3));
  inv1  gate1517(.a(s_139), .O(gate266inter4));
  nand2 gate1518(.a(gate266inter4), .b(gate266inter3), .O(gate266inter5));
  nor2  gate1519(.a(gate266inter5), .b(gate266inter2), .O(gate266inter6));
  inv1  gate1520(.a(G645), .O(gate266inter7));
  inv1  gate1521(.a(G773), .O(gate266inter8));
  nand2 gate1522(.a(gate266inter8), .b(gate266inter7), .O(gate266inter9));
  nand2 gate1523(.a(s_139), .b(gate266inter3), .O(gate266inter10));
  nor2  gate1524(.a(gate266inter10), .b(gate266inter9), .O(gate266inter11));
  nor2  gate1525(.a(gate266inter11), .b(gate266inter6), .O(gate266inter12));
  nand2 gate1526(.a(gate266inter12), .b(gate266inter1), .O(G797));

  xor2  gate2633(.a(G776), .b(G648), .O(gate267inter0));
  nand2 gate2634(.a(gate267inter0), .b(s_298), .O(gate267inter1));
  and2  gate2635(.a(G776), .b(G648), .O(gate267inter2));
  inv1  gate2636(.a(s_298), .O(gate267inter3));
  inv1  gate2637(.a(s_299), .O(gate267inter4));
  nand2 gate2638(.a(gate267inter4), .b(gate267inter3), .O(gate267inter5));
  nor2  gate2639(.a(gate267inter5), .b(gate267inter2), .O(gate267inter6));
  inv1  gate2640(.a(G648), .O(gate267inter7));
  inv1  gate2641(.a(G776), .O(gate267inter8));
  nand2 gate2642(.a(gate267inter8), .b(gate267inter7), .O(gate267inter9));
  nand2 gate2643(.a(s_299), .b(gate267inter3), .O(gate267inter10));
  nor2  gate2644(.a(gate267inter10), .b(gate267inter9), .O(gate267inter11));
  nor2  gate2645(.a(gate267inter11), .b(gate267inter6), .O(gate267inter12));
  nand2 gate2646(.a(gate267inter12), .b(gate267inter1), .O(G800));

  xor2  gate2521(.a(G779), .b(G651), .O(gate268inter0));
  nand2 gate2522(.a(gate268inter0), .b(s_282), .O(gate268inter1));
  and2  gate2523(.a(G779), .b(G651), .O(gate268inter2));
  inv1  gate2524(.a(s_282), .O(gate268inter3));
  inv1  gate2525(.a(s_283), .O(gate268inter4));
  nand2 gate2526(.a(gate268inter4), .b(gate268inter3), .O(gate268inter5));
  nor2  gate2527(.a(gate268inter5), .b(gate268inter2), .O(gate268inter6));
  inv1  gate2528(.a(G651), .O(gate268inter7));
  inv1  gate2529(.a(G779), .O(gate268inter8));
  nand2 gate2530(.a(gate268inter8), .b(gate268inter7), .O(gate268inter9));
  nand2 gate2531(.a(s_283), .b(gate268inter3), .O(gate268inter10));
  nor2  gate2532(.a(gate268inter10), .b(gate268inter9), .O(gate268inter11));
  nor2  gate2533(.a(gate268inter11), .b(gate268inter6), .O(gate268inter12));
  nand2 gate2534(.a(gate268inter12), .b(gate268inter1), .O(G803));
nand2 gate269( .a(G654), .b(G782), .O(G806) );
nand2 gate270( .a(G657), .b(G785), .O(G809) );
nand2 gate271( .a(G660), .b(G788), .O(G812) );

  xor2  gate757(.a(G791), .b(G663), .O(gate272inter0));
  nand2 gate758(.a(gate272inter0), .b(s_30), .O(gate272inter1));
  and2  gate759(.a(G791), .b(G663), .O(gate272inter2));
  inv1  gate760(.a(s_30), .O(gate272inter3));
  inv1  gate761(.a(s_31), .O(gate272inter4));
  nand2 gate762(.a(gate272inter4), .b(gate272inter3), .O(gate272inter5));
  nor2  gate763(.a(gate272inter5), .b(gate272inter2), .O(gate272inter6));
  inv1  gate764(.a(G663), .O(gate272inter7));
  inv1  gate765(.a(G791), .O(gate272inter8));
  nand2 gate766(.a(gate272inter8), .b(gate272inter7), .O(gate272inter9));
  nand2 gate767(.a(s_31), .b(gate272inter3), .O(gate272inter10));
  nor2  gate768(.a(gate272inter10), .b(gate272inter9), .O(gate272inter11));
  nor2  gate769(.a(gate272inter11), .b(gate272inter6), .O(gate272inter12));
  nand2 gate770(.a(gate272inter12), .b(gate272inter1), .O(G815));
nand2 gate273( .a(G642), .b(G794), .O(G818) );

  xor2  gate645(.a(G794), .b(G770), .O(gate274inter0));
  nand2 gate646(.a(gate274inter0), .b(s_14), .O(gate274inter1));
  and2  gate647(.a(G794), .b(G770), .O(gate274inter2));
  inv1  gate648(.a(s_14), .O(gate274inter3));
  inv1  gate649(.a(s_15), .O(gate274inter4));
  nand2 gate650(.a(gate274inter4), .b(gate274inter3), .O(gate274inter5));
  nor2  gate651(.a(gate274inter5), .b(gate274inter2), .O(gate274inter6));
  inv1  gate652(.a(G770), .O(gate274inter7));
  inv1  gate653(.a(G794), .O(gate274inter8));
  nand2 gate654(.a(gate274inter8), .b(gate274inter7), .O(gate274inter9));
  nand2 gate655(.a(s_15), .b(gate274inter3), .O(gate274inter10));
  nor2  gate656(.a(gate274inter10), .b(gate274inter9), .O(gate274inter11));
  nor2  gate657(.a(gate274inter11), .b(gate274inter6), .O(gate274inter12));
  nand2 gate658(.a(gate274inter12), .b(gate274inter1), .O(G819));

  xor2  gate2129(.a(G797), .b(G645), .O(gate275inter0));
  nand2 gate2130(.a(gate275inter0), .b(s_226), .O(gate275inter1));
  and2  gate2131(.a(G797), .b(G645), .O(gate275inter2));
  inv1  gate2132(.a(s_226), .O(gate275inter3));
  inv1  gate2133(.a(s_227), .O(gate275inter4));
  nand2 gate2134(.a(gate275inter4), .b(gate275inter3), .O(gate275inter5));
  nor2  gate2135(.a(gate275inter5), .b(gate275inter2), .O(gate275inter6));
  inv1  gate2136(.a(G645), .O(gate275inter7));
  inv1  gate2137(.a(G797), .O(gate275inter8));
  nand2 gate2138(.a(gate275inter8), .b(gate275inter7), .O(gate275inter9));
  nand2 gate2139(.a(s_227), .b(gate275inter3), .O(gate275inter10));
  nor2  gate2140(.a(gate275inter10), .b(gate275inter9), .O(gate275inter11));
  nor2  gate2141(.a(gate275inter11), .b(gate275inter6), .O(gate275inter12));
  nand2 gate2142(.a(gate275inter12), .b(gate275inter1), .O(G820));
nand2 gate276( .a(G773), .b(G797), .O(G821) );
nand2 gate277( .a(G648), .b(G800), .O(G822) );
nand2 gate278( .a(G776), .b(G800), .O(G823) );
nand2 gate279( .a(G651), .b(G803), .O(G824) );
nand2 gate280( .a(G779), .b(G803), .O(G825) );

  xor2  gate1485(.a(G806), .b(G654), .O(gate281inter0));
  nand2 gate1486(.a(gate281inter0), .b(s_134), .O(gate281inter1));
  and2  gate1487(.a(G806), .b(G654), .O(gate281inter2));
  inv1  gate1488(.a(s_134), .O(gate281inter3));
  inv1  gate1489(.a(s_135), .O(gate281inter4));
  nand2 gate1490(.a(gate281inter4), .b(gate281inter3), .O(gate281inter5));
  nor2  gate1491(.a(gate281inter5), .b(gate281inter2), .O(gate281inter6));
  inv1  gate1492(.a(G654), .O(gate281inter7));
  inv1  gate1493(.a(G806), .O(gate281inter8));
  nand2 gate1494(.a(gate281inter8), .b(gate281inter7), .O(gate281inter9));
  nand2 gate1495(.a(s_135), .b(gate281inter3), .O(gate281inter10));
  nor2  gate1496(.a(gate281inter10), .b(gate281inter9), .O(gate281inter11));
  nor2  gate1497(.a(gate281inter11), .b(gate281inter6), .O(gate281inter12));
  nand2 gate1498(.a(gate281inter12), .b(gate281inter1), .O(G826));
nand2 gate282( .a(G782), .b(G806), .O(G827) );
nand2 gate283( .a(G657), .b(G809), .O(G828) );
nand2 gate284( .a(G785), .b(G809), .O(G829) );
nand2 gate285( .a(G660), .b(G812), .O(G830) );

  xor2  gate1723(.a(G812), .b(G788), .O(gate286inter0));
  nand2 gate1724(.a(gate286inter0), .b(s_168), .O(gate286inter1));
  and2  gate1725(.a(G812), .b(G788), .O(gate286inter2));
  inv1  gate1726(.a(s_168), .O(gate286inter3));
  inv1  gate1727(.a(s_169), .O(gate286inter4));
  nand2 gate1728(.a(gate286inter4), .b(gate286inter3), .O(gate286inter5));
  nor2  gate1729(.a(gate286inter5), .b(gate286inter2), .O(gate286inter6));
  inv1  gate1730(.a(G788), .O(gate286inter7));
  inv1  gate1731(.a(G812), .O(gate286inter8));
  nand2 gate1732(.a(gate286inter8), .b(gate286inter7), .O(gate286inter9));
  nand2 gate1733(.a(s_169), .b(gate286inter3), .O(gate286inter10));
  nor2  gate1734(.a(gate286inter10), .b(gate286inter9), .O(gate286inter11));
  nor2  gate1735(.a(gate286inter11), .b(gate286inter6), .O(gate286inter12));
  nand2 gate1736(.a(gate286inter12), .b(gate286inter1), .O(G831));
nand2 gate287( .a(G663), .b(G815), .O(G832) );
nand2 gate288( .a(G791), .b(G815), .O(G833) );
nand2 gate289( .a(G818), .b(G819), .O(G834) );
nand2 gate290( .a(G820), .b(G821), .O(G847) );

  xor2  gate1975(.a(G823), .b(G822), .O(gate291inter0));
  nand2 gate1976(.a(gate291inter0), .b(s_204), .O(gate291inter1));
  and2  gate1977(.a(G823), .b(G822), .O(gate291inter2));
  inv1  gate1978(.a(s_204), .O(gate291inter3));
  inv1  gate1979(.a(s_205), .O(gate291inter4));
  nand2 gate1980(.a(gate291inter4), .b(gate291inter3), .O(gate291inter5));
  nor2  gate1981(.a(gate291inter5), .b(gate291inter2), .O(gate291inter6));
  inv1  gate1982(.a(G822), .O(gate291inter7));
  inv1  gate1983(.a(G823), .O(gate291inter8));
  nand2 gate1984(.a(gate291inter8), .b(gate291inter7), .O(gate291inter9));
  nand2 gate1985(.a(s_205), .b(gate291inter3), .O(gate291inter10));
  nor2  gate1986(.a(gate291inter10), .b(gate291inter9), .O(gate291inter11));
  nor2  gate1987(.a(gate291inter11), .b(gate291inter6), .O(gate291inter12));
  nand2 gate1988(.a(gate291inter12), .b(gate291inter1), .O(G860));
nand2 gate292( .a(G824), .b(G825), .O(G873) );

  xor2  gate1093(.a(G829), .b(G828), .O(gate293inter0));
  nand2 gate1094(.a(gate293inter0), .b(s_78), .O(gate293inter1));
  and2  gate1095(.a(G829), .b(G828), .O(gate293inter2));
  inv1  gate1096(.a(s_78), .O(gate293inter3));
  inv1  gate1097(.a(s_79), .O(gate293inter4));
  nand2 gate1098(.a(gate293inter4), .b(gate293inter3), .O(gate293inter5));
  nor2  gate1099(.a(gate293inter5), .b(gate293inter2), .O(gate293inter6));
  inv1  gate1100(.a(G828), .O(gate293inter7));
  inv1  gate1101(.a(G829), .O(gate293inter8));
  nand2 gate1102(.a(gate293inter8), .b(gate293inter7), .O(gate293inter9));
  nand2 gate1103(.a(s_79), .b(gate293inter3), .O(gate293inter10));
  nor2  gate1104(.a(gate293inter10), .b(gate293inter9), .O(gate293inter11));
  nor2  gate1105(.a(gate293inter11), .b(gate293inter6), .O(gate293inter12));
  nand2 gate1106(.a(gate293inter12), .b(gate293inter1), .O(G886));
nand2 gate294( .a(G832), .b(G833), .O(G899) );
nand2 gate295( .a(G830), .b(G831), .O(G912) );

  xor2  gate2759(.a(G827), .b(G826), .O(gate296inter0));
  nand2 gate2760(.a(gate296inter0), .b(s_316), .O(gate296inter1));
  and2  gate2761(.a(G827), .b(G826), .O(gate296inter2));
  inv1  gate2762(.a(s_316), .O(gate296inter3));
  inv1  gate2763(.a(s_317), .O(gate296inter4));
  nand2 gate2764(.a(gate296inter4), .b(gate296inter3), .O(gate296inter5));
  nor2  gate2765(.a(gate296inter5), .b(gate296inter2), .O(gate296inter6));
  inv1  gate2766(.a(G826), .O(gate296inter7));
  inv1  gate2767(.a(G827), .O(gate296inter8));
  nand2 gate2768(.a(gate296inter8), .b(gate296inter7), .O(gate296inter9));
  nand2 gate2769(.a(s_317), .b(gate296inter3), .O(gate296inter10));
  nor2  gate2770(.a(gate296inter10), .b(gate296inter9), .O(gate296inter11));
  nor2  gate2771(.a(gate296inter11), .b(gate296inter6), .O(gate296inter12));
  nand2 gate2772(.a(gate296inter12), .b(gate296inter1), .O(G925));
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );
nand2 gate387( .a(G1), .b(G1036), .O(G1132) );
nand2 gate388( .a(G2), .b(G1039), .O(G1135) );

  xor2  gate1023(.a(G1042), .b(G3), .O(gate389inter0));
  nand2 gate1024(.a(gate389inter0), .b(s_68), .O(gate389inter1));
  and2  gate1025(.a(G1042), .b(G3), .O(gate389inter2));
  inv1  gate1026(.a(s_68), .O(gate389inter3));
  inv1  gate1027(.a(s_69), .O(gate389inter4));
  nand2 gate1028(.a(gate389inter4), .b(gate389inter3), .O(gate389inter5));
  nor2  gate1029(.a(gate389inter5), .b(gate389inter2), .O(gate389inter6));
  inv1  gate1030(.a(G3), .O(gate389inter7));
  inv1  gate1031(.a(G1042), .O(gate389inter8));
  nand2 gate1032(.a(gate389inter8), .b(gate389inter7), .O(gate389inter9));
  nand2 gate1033(.a(s_69), .b(gate389inter3), .O(gate389inter10));
  nor2  gate1034(.a(gate389inter10), .b(gate389inter9), .O(gate389inter11));
  nor2  gate1035(.a(gate389inter11), .b(gate389inter6), .O(gate389inter12));
  nand2 gate1036(.a(gate389inter12), .b(gate389inter1), .O(G1138));
nand2 gate390( .a(G4), .b(G1045), .O(G1141) );
nand2 gate391( .a(G5), .b(G1048), .O(G1144) );
nand2 gate392( .a(G6), .b(G1051), .O(G1147) );
nand2 gate393( .a(G7), .b(G1054), .O(G1150) );
nand2 gate394( .a(G8), .b(G1057), .O(G1153) );

  xor2  gate2325(.a(G1060), .b(G9), .O(gate395inter0));
  nand2 gate2326(.a(gate395inter0), .b(s_254), .O(gate395inter1));
  and2  gate2327(.a(G1060), .b(G9), .O(gate395inter2));
  inv1  gate2328(.a(s_254), .O(gate395inter3));
  inv1  gate2329(.a(s_255), .O(gate395inter4));
  nand2 gate2330(.a(gate395inter4), .b(gate395inter3), .O(gate395inter5));
  nor2  gate2331(.a(gate395inter5), .b(gate395inter2), .O(gate395inter6));
  inv1  gate2332(.a(G9), .O(gate395inter7));
  inv1  gate2333(.a(G1060), .O(gate395inter8));
  nand2 gate2334(.a(gate395inter8), .b(gate395inter7), .O(gate395inter9));
  nand2 gate2335(.a(s_255), .b(gate395inter3), .O(gate395inter10));
  nor2  gate2336(.a(gate395inter10), .b(gate395inter9), .O(gate395inter11));
  nor2  gate2337(.a(gate395inter11), .b(gate395inter6), .O(gate395inter12));
  nand2 gate2338(.a(gate395inter12), .b(gate395inter1), .O(G1156));
nand2 gate396( .a(G10), .b(G1063), .O(G1159) );
nand2 gate397( .a(G11), .b(G1066), .O(G1162) );
nand2 gate398( .a(G12), .b(G1069), .O(G1165) );

  xor2  gate603(.a(G1072), .b(G13), .O(gate399inter0));
  nand2 gate604(.a(gate399inter0), .b(s_8), .O(gate399inter1));
  and2  gate605(.a(G1072), .b(G13), .O(gate399inter2));
  inv1  gate606(.a(s_8), .O(gate399inter3));
  inv1  gate607(.a(s_9), .O(gate399inter4));
  nand2 gate608(.a(gate399inter4), .b(gate399inter3), .O(gate399inter5));
  nor2  gate609(.a(gate399inter5), .b(gate399inter2), .O(gate399inter6));
  inv1  gate610(.a(G13), .O(gate399inter7));
  inv1  gate611(.a(G1072), .O(gate399inter8));
  nand2 gate612(.a(gate399inter8), .b(gate399inter7), .O(gate399inter9));
  nand2 gate613(.a(s_9), .b(gate399inter3), .O(gate399inter10));
  nor2  gate614(.a(gate399inter10), .b(gate399inter9), .O(gate399inter11));
  nor2  gate615(.a(gate399inter11), .b(gate399inter6), .O(gate399inter12));
  nand2 gate616(.a(gate399inter12), .b(gate399inter1), .O(G1168));
nand2 gate400( .a(G14), .b(G1075), .O(G1171) );
nand2 gate401( .a(G15), .b(G1078), .O(G1174) );
nand2 gate402( .a(G16), .b(G1081), .O(G1177) );

  xor2  gate1541(.a(G1084), .b(G17), .O(gate403inter0));
  nand2 gate1542(.a(gate403inter0), .b(s_142), .O(gate403inter1));
  and2  gate1543(.a(G1084), .b(G17), .O(gate403inter2));
  inv1  gate1544(.a(s_142), .O(gate403inter3));
  inv1  gate1545(.a(s_143), .O(gate403inter4));
  nand2 gate1546(.a(gate403inter4), .b(gate403inter3), .O(gate403inter5));
  nor2  gate1547(.a(gate403inter5), .b(gate403inter2), .O(gate403inter6));
  inv1  gate1548(.a(G17), .O(gate403inter7));
  inv1  gate1549(.a(G1084), .O(gate403inter8));
  nand2 gate1550(.a(gate403inter8), .b(gate403inter7), .O(gate403inter9));
  nand2 gate1551(.a(s_143), .b(gate403inter3), .O(gate403inter10));
  nor2  gate1552(.a(gate403inter10), .b(gate403inter9), .O(gate403inter11));
  nor2  gate1553(.a(gate403inter11), .b(gate403inter6), .O(gate403inter12));
  nand2 gate1554(.a(gate403inter12), .b(gate403inter1), .O(G1180));
nand2 gate404( .a(G18), .b(G1087), .O(G1183) );

  xor2  gate1779(.a(G1090), .b(G19), .O(gate405inter0));
  nand2 gate1780(.a(gate405inter0), .b(s_176), .O(gate405inter1));
  and2  gate1781(.a(G1090), .b(G19), .O(gate405inter2));
  inv1  gate1782(.a(s_176), .O(gate405inter3));
  inv1  gate1783(.a(s_177), .O(gate405inter4));
  nand2 gate1784(.a(gate405inter4), .b(gate405inter3), .O(gate405inter5));
  nor2  gate1785(.a(gate405inter5), .b(gate405inter2), .O(gate405inter6));
  inv1  gate1786(.a(G19), .O(gate405inter7));
  inv1  gate1787(.a(G1090), .O(gate405inter8));
  nand2 gate1788(.a(gate405inter8), .b(gate405inter7), .O(gate405inter9));
  nand2 gate1789(.a(s_177), .b(gate405inter3), .O(gate405inter10));
  nor2  gate1790(.a(gate405inter10), .b(gate405inter9), .O(gate405inter11));
  nor2  gate1791(.a(gate405inter11), .b(gate405inter6), .O(gate405inter12));
  nand2 gate1792(.a(gate405inter12), .b(gate405inter1), .O(G1186));
nand2 gate406( .a(G20), .b(G1093), .O(G1189) );
nand2 gate407( .a(G21), .b(G1096), .O(G1192) );

  xor2  gate2045(.a(G1099), .b(G22), .O(gate408inter0));
  nand2 gate2046(.a(gate408inter0), .b(s_214), .O(gate408inter1));
  and2  gate2047(.a(G1099), .b(G22), .O(gate408inter2));
  inv1  gate2048(.a(s_214), .O(gate408inter3));
  inv1  gate2049(.a(s_215), .O(gate408inter4));
  nand2 gate2050(.a(gate408inter4), .b(gate408inter3), .O(gate408inter5));
  nor2  gate2051(.a(gate408inter5), .b(gate408inter2), .O(gate408inter6));
  inv1  gate2052(.a(G22), .O(gate408inter7));
  inv1  gate2053(.a(G1099), .O(gate408inter8));
  nand2 gate2054(.a(gate408inter8), .b(gate408inter7), .O(gate408inter9));
  nand2 gate2055(.a(s_215), .b(gate408inter3), .O(gate408inter10));
  nor2  gate2056(.a(gate408inter10), .b(gate408inter9), .O(gate408inter11));
  nor2  gate2057(.a(gate408inter11), .b(gate408inter6), .O(gate408inter12));
  nand2 gate2058(.a(gate408inter12), .b(gate408inter1), .O(G1195));
nand2 gate409( .a(G23), .b(G1102), .O(G1198) );
nand2 gate410( .a(G24), .b(G1105), .O(G1201) );

  xor2  gate1751(.a(G1108), .b(G25), .O(gate411inter0));
  nand2 gate1752(.a(gate411inter0), .b(s_172), .O(gate411inter1));
  and2  gate1753(.a(G1108), .b(G25), .O(gate411inter2));
  inv1  gate1754(.a(s_172), .O(gate411inter3));
  inv1  gate1755(.a(s_173), .O(gate411inter4));
  nand2 gate1756(.a(gate411inter4), .b(gate411inter3), .O(gate411inter5));
  nor2  gate1757(.a(gate411inter5), .b(gate411inter2), .O(gate411inter6));
  inv1  gate1758(.a(G25), .O(gate411inter7));
  inv1  gate1759(.a(G1108), .O(gate411inter8));
  nand2 gate1760(.a(gate411inter8), .b(gate411inter7), .O(gate411inter9));
  nand2 gate1761(.a(s_173), .b(gate411inter3), .O(gate411inter10));
  nor2  gate1762(.a(gate411inter10), .b(gate411inter9), .O(gate411inter11));
  nor2  gate1763(.a(gate411inter11), .b(gate411inter6), .O(gate411inter12));
  nand2 gate1764(.a(gate411inter12), .b(gate411inter1), .O(G1204));

  xor2  gate2115(.a(G1111), .b(G26), .O(gate412inter0));
  nand2 gate2116(.a(gate412inter0), .b(s_224), .O(gate412inter1));
  and2  gate2117(.a(G1111), .b(G26), .O(gate412inter2));
  inv1  gate2118(.a(s_224), .O(gate412inter3));
  inv1  gate2119(.a(s_225), .O(gate412inter4));
  nand2 gate2120(.a(gate412inter4), .b(gate412inter3), .O(gate412inter5));
  nor2  gate2121(.a(gate412inter5), .b(gate412inter2), .O(gate412inter6));
  inv1  gate2122(.a(G26), .O(gate412inter7));
  inv1  gate2123(.a(G1111), .O(gate412inter8));
  nand2 gate2124(.a(gate412inter8), .b(gate412inter7), .O(gate412inter9));
  nand2 gate2125(.a(s_225), .b(gate412inter3), .O(gate412inter10));
  nor2  gate2126(.a(gate412inter10), .b(gate412inter9), .O(gate412inter11));
  nor2  gate2127(.a(gate412inter11), .b(gate412inter6), .O(gate412inter12));
  nand2 gate2128(.a(gate412inter12), .b(gate412inter1), .O(G1207));
nand2 gate413( .a(G27), .b(G1114), .O(G1210) );

  xor2  gate1961(.a(G1117), .b(G28), .O(gate414inter0));
  nand2 gate1962(.a(gate414inter0), .b(s_202), .O(gate414inter1));
  and2  gate1963(.a(G1117), .b(G28), .O(gate414inter2));
  inv1  gate1964(.a(s_202), .O(gate414inter3));
  inv1  gate1965(.a(s_203), .O(gate414inter4));
  nand2 gate1966(.a(gate414inter4), .b(gate414inter3), .O(gate414inter5));
  nor2  gate1967(.a(gate414inter5), .b(gate414inter2), .O(gate414inter6));
  inv1  gate1968(.a(G28), .O(gate414inter7));
  inv1  gate1969(.a(G1117), .O(gate414inter8));
  nand2 gate1970(.a(gate414inter8), .b(gate414inter7), .O(gate414inter9));
  nand2 gate1971(.a(s_203), .b(gate414inter3), .O(gate414inter10));
  nor2  gate1972(.a(gate414inter10), .b(gate414inter9), .O(gate414inter11));
  nor2  gate1973(.a(gate414inter11), .b(gate414inter6), .O(gate414inter12));
  nand2 gate1974(.a(gate414inter12), .b(gate414inter1), .O(G1213));
nand2 gate415( .a(G29), .b(G1120), .O(G1216) );
nand2 gate416( .a(G30), .b(G1123), .O(G1219) );

  xor2  gate1905(.a(G1126), .b(G31), .O(gate417inter0));
  nand2 gate1906(.a(gate417inter0), .b(s_194), .O(gate417inter1));
  and2  gate1907(.a(G1126), .b(G31), .O(gate417inter2));
  inv1  gate1908(.a(s_194), .O(gate417inter3));
  inv1  gate1909(.a(s_195), .O(gate417inter4));
  nand2 gate1910(.a(gate417inter4), .b(gate417inter3), .O(gate417inter5));
  nor2  gate1911(.a(gate417inter5), .b(gate417inter2), .O(gate417inter6));
  inv1  gate1912(.a(G31), .O(gate417inter7));
  inv1  gate1913(.a(G1126), .O(gate417inter8));
  nand2 gate1914(.a(gate417inter8), .b(gate417inter7), .O(gate417inter9));
  nand2 gate1915(.a(s_195), .b(gate417inter3), .O(gate417inter10));
  nor2  gate1916(.a(gate417inter10), .b(gate417inter9), .O(gate417inter11));
  nor2  gate1917(.a(gate417inter11), .b(gate417inter6), .O(gate417inter12));
  nand2 gate1918(.a(gate417inter12), .b(gate417inter1), .O(G1222));

  xor2  gate2269(.a(G1129), .b(G32), .O(gate418inter0));
  nand2 gate2270(.a(gate418inter0), .b(s_246), .O(gate418inter1));
  and2  gate2271(.a(G1129), .b(G32), .O(gate418inter2));
  inv1  gate2272(.a(s_246), .O(gate418inter3));
  inv1  gate2273(.a(s_247), .O(gate418inter4));
  nand2 gate2274(.a(gate418inter4), .b(gate418inter3), .O(gate418inter5));
  nor2  gate2275(.a(gate418inter5), .b(gate418inter2), .O(gate418inter6));
  inv1  gate2276(.a(G32), .O(gate418inter7));
  inv1  gate2277(.a(G1129), .O(gate418inter8));
  nand2 gate2278(.a(gate418inter8), .b(gate418inter7), .O(gate418inter9));
  nand2 gate2279(.a(s_247), .b(gate418inter3), .O(gate418inter10));
  nor2  gate2280(.a(gate418inter10), .b(gate418inter9), .O(gate418inter11));
  nor2  gate2281(.a(gate418inter11), .b(gate418inter6), .O(gate418inter12));
  nand2 gate2282(.a(gate418inter12), .b(gate418inter1), .O(G1225));

  xor2  gate2353(.a(G1132), .b(G1), .O(gate419inter0));
  nand2 gate2354(.a(gate419inter0), .b(s_258), .O(gate419inter1));
  and2  gate2355(.a(G1132), .b(G1), .O(gate419inter2));
  inv1  gate2356(.a(s_258), .O(gate419inter3));
  inv1  gate2357(.a(s_259), .O(gate419inter4));
  nand2 gate2358(.a(gate419inter4), .b(gate419inter3), .O(gate419inter5));
  nor2  gate2359(.a(gate419inter5), .b(gate419inter2), .O(gate419inter6));
  inv1  gate2360(.a(G1), .O(gate419inter7));
  inv1  gate2361(.a(G1132), .O(gate419inter8));
  nand2 gate2362(.a(gate419inter8), .b(gate419inter7), .O(gate419inter9));
  nand2 gate2363(.a(s_259), .b(gate419inter3), .O(gate419inter10));
  nor2  gate2364(.a(gate419inter10), .b(gate419inter9), .O(gate419inter11));
  nor2  gate2365(.a(gate419inter11), .b(gate419inter6), .O(gate419inter12));
  nand2 gate2366(.a(gate419inter12), .b(gate419inter1), .O(G1228));
nand2 gate420( .a(G1036), .b(G1132), .O(G1229) );
nand2 gate421( .a(G2), .b(G1135), .O(G1230) );
nand2 gate422( .a(G1039), .b(G1135), .O(G1231) );

  xor2  gate785(.a(G1138), .b(G3), .O(gate423inter0));
  nand2 gate786(.a(gate423inter0), .b(s_34), .O(gate423inter1));
  and2  gate787(.a(G1138), .b(G3), .O(gate423inter2));
  inv1  gate788(.a(s_34), .O(gate423inter3));
  inv1  gate789(.a(s_35), .O(gate423inter4));
  nand2 gate790(.a(gate423inter4), .b(gate423inter3), .O(gate423inter5));
  nor2  gate791(.a(gate423inter5), .b(gate423inter2), .O(gate423inter6));
  inv1  gate792(.a(G3), .O(gate423inter7));
  inv1  gate793(.a(G1138), .O(gate423inter8));
  nand2 gate794(.a(gate423inter8), .b(gate423inter7), .O(gate423inter9));
  nand2 gate795(.a(s_35), .b(gate423inter3), .O(gate423inter10));
  nor2  gate796(.a(gate423inter10), .b(gate423inter9), .O(gate423inter11));
  nor2  gate797(.a(gate423inter11), .b(gate423inter6), .O(gate423inter12));
  nand2 gate798(.a(gate423inter12), .b(gate423inter1), .O(G1232));
nand2 gate424( .a(G1042), .b(G1138), .O(G1233) );
nand2 gate425( .a(G4), .b(G1141), .O(G1234) );
nand2 gate426( .a(G1045), .b(G1141), .O(G1235) );

  xor2  gate2731(.a(G1144), .b(G5), .O(gate427inter0));
  nand2 gate2732(.a(gate427inter0), .b(s_312), .O(gate427inter1));
  and2  gate2733(.a(G1144), .b(G5), .O(gate427inter2));
  inv1  gate2734(.a(s_312), .O(gate427inter3));
  inv1  gate2735(.a(s_313), .O(gate427inter4));
  nand2 gate2736(.a(gate427inter4), .b(gate427inter3), .O(gate427inter5));
  nor2  gate2737(.a(gate427inter5), .b(gate427inter2), .O(gate427inter6));
  inv1  gate2738(.a(G5), .O(gate427inter7));
  inv1  gate2739(.a(G1144), .O(gate427inter8));
  nand2 gate2740(.a(gate427inter8), .b(gate427inter7), .O(gate427inter9));
  nand2 gate2741(.a(s_313), .b(gate427inter3), .O(gate427inter10));
  nor2  gate2742(.a(gate427inter10), .b(gate427inter9), .O(gate427inter11));
  nor2  gate2743(.a(gate427inter11), .b(gate427inter6), .O(gate427inter12));
  nand2 gate2744(.a(gate427inter12), .b(gate427inter1), .O(G1236));

  xor2  gate2213(.a(G1144), .b(G1048), .O(gate428inter0));
  nand2 gate2214(.a(gate428inter0), .b(s_238), .O(gate428inter1));
  and2  gate2215(.a(G1144), .b(G1048), .O(gate428inter2));
  inv1  gate2216(.a(s_238), .O(gate428inter3));
  inv1  gate2217(.a(s_239), .O(gate428inter4));
  nand2 gate2218(.a(gate428inter4), .b(gate428inter3), .O(gate428inter5));
  nor2  gate2219(.a(gate428inter5), .b(gate428inter2), .O(gate428inter6));
  inv1  gate2220(.a(G1048), .O(gate428inter7));
  inv1  gate2221(.a(G1144), .O(gate428inter8));
  nand2 gate2222(.a(gate428inter8), .b(gate428inter7), .O(gate428inter9));
  nand2 gate2223(.a(s_239), .b(gate428inter3), .O(gate428inter10));
  nor2  gate2224(.a(gate428inter10), .b(gate428inter9), .O(gate428inter11));
  nor2  gate2225(.a(gate428inter11), .b(gate428inter6), .O(gate428inter12));
  nand2 gate2226(.a(gate428inter12), .b(gate428inter1), .O(G1237));
nand2 gate429( .a(G6), .b(G1147), .O(G1238) );

  xor2  gate2185(.a(G1147), .b(G1051), .O(gate430inter0));
  nand2 gate2186(.a(gate430inter0), .b(s_234), .O(gate430inter1));
  and2  gate2187(.a(G1147), .b(G1051), .O(gate430inter2));
  inv1  gate2188(.a(s_234), .O(gate430inter3));
  inv1  gate2189(.a(s_235), .O(gate430inter4));
  nand2 gate2190(.a(gate430inter4), .b(gate430inter3), .O(gate430inter5));
  nor2  gate2191(.a(gate430inter5), .b(gate430inter2), .O(gate430inter6));
  inv1  gate2192(.a(G1051), .O(gate430inter7));
  inv1  gate2193(.a(G1147), .O(gate430inter8));
  nand2 gate2194(.a(gate430inter8), .b(gate430inter7), .O(gate430inter9));
  nand2 gate2195(.a(s_235), .b(gate430inter3), .O(gate430inter10));
  nor2  gate2196(.a(gate430inter10), .b(gate430inter9), .O(gate430inter11));
  nor2  gate2197(.a(gate430inter11), .b(gate430inter6), .O(gate430inter12));
  nand2 gate2198(.a(gate430inter12), .b(gate430inter1), .O(G1239));
nand2 gate431( .a(G7), .b(G1150), .O(G1240) );
nand2 gate432( .a(G1054), .b(G1150), .O(G1241) );
nand2 gate433( .a(G8), .b(G1153), .O(G1242) );
nand2 gate434( .a(G1057), .b(G1153), .O(G1243) );
nand2 gate435( .a(G9), .b(G1156), .O(G1244) );

  xor2  gate1527(.a(G1156), .b(G1060), .O(gate436inter0));
  nand2 gate1528(.a(gate436inter0), .b(s_140), .O(gate436inter1));
  and2  gate1529(.a(G1156), .b(G1060), .O(gate436inter2));
  inv1  gate1530(.a(s_140), .O(gate436inter3));
  inv1  gate1531(.a(s_141), .O(gate436inter4));
  nand2 gate1532(.a(gate436inter4), .b(gate436inter3), .O(gate436inter5));
  nor2  gate1533(.a(gate436inter5), .b(gate436inter2), .O(gate436inter6));
  inv1  gate1534(.a(G1060), .O(gate436inter7));
  inv1  gate1535(.a(G1156), .O(gate436inter8));
  nand2 gate1536(.a(gate436inter8), .b(gate436inter7), .O(gate436inter9));
  nand2 gate1537(.a(s_141), .b(gate436inter3), .O(gate436inter10));
  nor2  gate1538(.a(gate436inter10), .b(gate436inter9), .O(gate436inter11));
  nor2  gate1539(.a(gate436inter11), .b(gate436inter6), .O(gate436inter12));
  nand2 gate1540(.a(gate436inter12), .b(gate436inter1), .O(G1245));

  xor2  gate2661(.a(G1159), .b(G10), .O(gate437inter0));
  nand2 gate2662(.a(gate437inter0), .b(s_302), .O(gate437inter1));
  and2  gate2663(.a(G1159), .b(G10), .O(gate437inter2));
  inv1  gate2664(.a(s_302), .O(gate437inter3));
  inv1  gate2665(.a(s_303), .O(gate437inter4));
  nand2 gate2666(.a(gate437inter4), .b(gate437inter3), .O(gate437inter5));
  nor2  gate2667(.a(gate437inter5), .b(gate437inter2), .O(gate437inter6));
  inv1  gate2668(.a(G10), .O(gate437inter7));
  inv1  gate2669(.a(G1159), .O(gate437inter8));
  nand2 gate2670(.a(gate437inter8), .b(gate437inter7), .O(gate437inter9));
  nand2 gate2671(.a(s_303), .b(gate437inter3), .O(gate437inter10));
  nor2  gate2672(.a(gate437inter10), .b(gate437inter9), .O(gate437inter11));
  nor2  gate2673(.a(gate437inter11), .b(gate437inter6), .O(gate437inter12));
  nand2 gate2674(.a(gate437inter12), .b(gate437inter1), .O(G1246));
nand2 gate438( .a(G1063), .b(G1159), .O(G1247) );
nand2 gate439( .a(G11), .b(G1162), .O(G1248) );

  xor2  gate1919(.a(G1162), .b(G1066), .O(gate440inter0));
  nand2 gate1920(.a(gate440inter0), .b(s_196), .O(gate440inter1));
  and2  gate1921(.a(G1162), .b(G1066), .O(gate440inter2));
  inv1  gate1922(.a(s_196), .O(gate440inter3));
  inv1  gate1923(.a(s_197), .O(gate440inter4));
  nand2 gate1924(.a(gate440inter4), .b(gate440inter3), .O(gate440inter5));
  nor2  gate1925(.a(gate440inter5), .b(gate440inter2), .O(gate440inter6));
  inv1  gate1926(.a(G1066), .O(gate440inter7));
  inv1  gate1927(.a(G1162), .O(gate440inter8));
  nand2 gate1928(.a(gate440inter8), .b(gate440inter7), .O(gate440inter9));
  nand2 gate1929(.a(s_197), .b(gate440inter3), .O(gate440inter10));
  nor2  gate1930(.a(gate440inter10), .b(gate440inter9), .O(gate440inter11));
  nor2  gate1931(.a(gate440inter11), .b(gate440inter6), .O(gate440inter12));
  nand2 gate1932(.a(gate440inter12), .b(gate440inter1), .O(G1249));
nand2 gate441( .a(G12), .b(G1165), .O(G1250) );
nand2 gate442( .a(G1069), .b(G1165), .O(G1251) );

  xor2  gate1303(.a(G1168), .b(G13), .O(gate443inter0));
  nand2 gate1304(.a(gate443inter0), .b(s_108), .O(gate443inter1));
  and2  gate1305(.a(G1168), .b(G13), .O(gate443inter2));
  inv1  gate1306(.a(s_108), .O(gate443inter3));
  inv1  gate1307(.a(s_109), .O(gate443inter4));
  nand2 gate1308(.a(gate443inter4), .b(gate443inter3), .O(gate443inter5));
  nor2  gate1309(.a(gate443inter5), .b(gate443inter2), .O(gate443inter6));
  inv1  gate1310(.a(G13), .O(gate443inter7));
  inv1  gate1311(.a(G1168), .O(gate443inter8));
  nand2 gate1312(.a(gate443inter8), .b(gate443inter7), .O(gate443inter9));
  nand2 gate1313(.a(s_109), .b(gate443inter3), .O(gate443inter10));
  nor2  gate1314(.a(gate443inter10), .b(gate443inter9), .O(gate443inter11));
  nor2  gate1315(.a(gate443inter11), .b(gate443inter6), .O(gate443inter12));
  nand2 gate1316(.a(gate443inter12), .b(gate443inter1), .O(G1252));
nand2 gate444( .a(G1072), .b(G1168), .O(G1253) );
nand2 gate445( .a(G14), .b(G1171), .O(G1254) );
nand2 gate446( .a(G1075), .b(G1171), .O(G1255) );
nand2 gate447( .a(G15), .b(G1174), .O(G1256) );

  xor2  gate1443(.a(G1174), .b(G1078), .O(gate448inter0));
  nand2 gate1444(.a(gate448inter0), .b(s_128), .O(gate448inter1));
  and2  gate1445(.a(G1174), .b(G1078), .O(gate448inter2));
  inv1  gate1446(.a(s_128), .O(gate448inter3));
  inv1  gate1447(.a(s_129), .O(gate448inter4));
  nand2 gate1448(.a(gate448inter4), .b(gate448inter3), .O(gate448inter5));
  nor2  gate1449(.a(gate448inter5), .b(gate448inter2), .O(gate448inter6));
  inv1  gate1450(.a(G1078), .O(gate448inter7));
  inv1  gate1451(.a(G1174), .O(gate448inter8));
  nand2 gate1452(.a(gate448inter8), .b(gate448inter7), .O(gate448inter9));
  nand2 gate1453(.a(s_129), .b(gate448inter3), .O(gate448inter10));
  nor2  gate1454(.a(gate448inter10), .b(gate448inter9), .O(gate448inter11));
  nor2  gate1455(.a(gate448inter11), .b(gate448inter6), .O(gate448inter12));
  nand2 gate1456(.a(gate448inter12), .b(gate448inter1), .O(G1257));
nand2 gate449( .a(G16), .b(G1177), .O(G1258) );

  xor2  gate1653(.a(G1177), .b(G1081), .O(gate450inter0));
  nand2 gate1654(.a(gate450inter0), .b(s_158), .O(gate450inter1));
  and2  gate1655(.a(G1177), .b(G1081), .O(gate450inter2));
  inv1  gate1656(.a(s_158), .O(gate450inter3));
  inv1  gate1657(.a(s_159), .O(gate450inter4));
  nand2 gate1658(.a(gate450inter4), .b(gate450inter3), .O(gate450inter5));
  nor2  gate1659(.a(gate450inter5), .b(gate450inter2), .O(gate450inter6));
  inv1  gate1660(.a(G1081), .O(gate450inter7));
  inv1  gate1661(.a(G1177), .O(gate450inter8));
  nand2 gate1662(.a(gate450inter8), .b(gate450inter7), .O(gate450inter9));
  nand2 gate1663(.a(s_159), .b(gate450inter3), .O(gate450inter10));
  nor2  gate1664(.a(gate450inter10), .b(gate450inter9), .O(gate450inter11));
  nor2  gate1665(.a(gate450inter11), .b(gate450inter6), .O(gate450inter12));
  nand2 gate1666(.a(gate450inter12), .b(gate450inter1), .O(G1259));

  xor2  gate1681(.a(G1180), .b(G17), .O(gate451inter0));
  nand2 gate1682(.a(gate451inter0), .b(s_162), .O(gate451inter1));
  and2  gate1683(.a(G1180), .b(G17), .O(gate451inter2));
  inv1  gate1684(.a(s_162), .O(gate451inter3));
  inv1  gate1685(.a(s_163), .O(gate451inter4));
  nand2 gate1686(.a(gate451inter4), .b(gate451inter3), .O(gate451inter5));
  nor2  gate1687(.a(gate451inter5), .b(gate451inter2), .O(gate451inter6));
  inv1  gate1688(.a(G17), .O(gate451inter7));
  inv1  gate1689(.a(G1180), .O(gate451inter8));
  nand2 gate1690(.a(gate451inter8), .b(gate451inter7), .O(gate451inter9));
  nand2 gate1691(.a(s_163), .b(gate451inter3), .O(gate451inter10));
  nor2  gate1692(.a(gate451inter10), .b(gate451inter9), .O(gate451inter11));
  nor2  gate1693(.a(gate451inter11), .b(gate451inter6), .O(gate451inter12));
  nand2 gate1694(.a(gate451inter12), .b(gate451inter1), .O(G1260));
nand2 gate452( .a(G1084), .b(G1180), .O(G1261) );
nand2 gate453( .a(G18), .b(G1183), .O(G1262) );

  xor2  gate855(.a(G1183), .b(G1087), .O(gate454inter0));
  nand2 gate856(.a(gate454inter0), .b(s_44), .O(gate454inter1));
  and2  gate857(.a(G1183), .b(G1087), .O(gate454inter2));
  inv1  gate858(.a(s_44), .O(gate454inter3));
  inv1  gate859(.a(s_45), .O(gate454inter4));
  nand2 gate860(.a(gate454inter4), .b(gate454inter3), .O(gate454inter5));
  nor2  gate861(.a(gate454inter5), .b(gate454inter2), .O(gate454inter6));
  inv1  gate862(.a(G1087), .O(gate454inter7));
  inv1  gate863(.a(G1183), .O(gate454inter8));
  nand2 gate864(.a(gate454inter8), .b(gate454inter7), .O(gate454inter9));
  nand2 gate865(.a(s_45), .b(gate454inter3), .O(gate454inter10));
  nor2  gate866(.a(gate454inter10), .b(gate454inter9), .O(gate454inter11));
  nor2  gate867(.a(gate454inter11), .b(gate454inter6), .O(gate454inter12));
  nand2 gate868(.a(gate454inter12), .b(gate454inter1), .O(G1263));

  xor2  gate911(.a(G1186), .b(G19), .O(gate455inter0));
  nand2 gate912(.a(gate455inter0), .b(s_52), .O(gate455inter1));
  and2  gate913(.a(G1186), .b(G19), .O(gate455inter2));
  inv1  gate914(.a(s_52), .O(gate455inter3));
  inv1  gate915(.a(s_53), .O(gate455inter4));
  nand2 gate916(.a(gate455inter4), .b(gate455inter3), .O(gate455inter5));
  nor2  gate917(.a(gate455inter5), .b(gate455inter2), .O(gate455inter6));
  inv1  gate918(.a(G19), .O(gate455inter7));
  inv1  gate919(.a(G1186), .O(gate455inter8));
  nand2 gate920(.a(gate455inter8), .b(gate455inter7), .O(gate455inter9));
  nand2 gate921(.a(s_53), .b(gate455inter3), .O(gate455inter10));
  nor2  gate922(.a(gate455inter10), .b(gate455inter9), .O(gate455inter11));
  nor2  gate923(.a(gate455inter11), .b(gate455inter6), .O(gate455inter12));
  nand2 gate924(.a(gate455inter12), .b(gate455inter1), .O(G1264));
nand2 gate456( .a(G1090), .b(G1186), .O(G1265) );

  xor2  gate1219(.a(G1189), .b(G20), .O(gate457inter0));
  nand2 gate1220(.a(gate457inter0), .b(s_96), .O(gate457inter1));
  and2  gate1221(.a(G1189), .b(G20), .O(gate457inter2));
  inv1  gate1222(.a(s_96), .O(gate457inter3));
  inv1  gate1223(.a(s_97), .O(gate457inter4));
  nand2 gate1224(.a(gate457inter4), .b(gate457inter3), .O(gate457inter5));
  nor2  gate1225(.a(gate457inter5), .b(gate457inter2), .O(gate457inter6));
  inv1  gate1226(.a(G20), .O(gate457inter7));
  inv1  gate1227(.a(G1189), .O(gate457inter8));
  nand2 gate1228(.a(gate457inter8), .b(gate457inter7), .O(gate457inter9));
  nand2 gate1229(.a(s_97), .b(gate457inter3), .O(gate457inter10));
  nor2  gate1230(.a(gate457inter10), .b(gate457inter9), .O(gate457inter11));
  nor2  gate1231(.a(gate457inter11), .b(gate457inter6), .O(gate457inter12));
  nand2 gate1232(.a(gate457inter12), .b(gate457inter1), .O(G1266));
nand2 gate458( .a(G1093), .b(G1189), .O(G1267) );
nand2 gate459( .a(G21), .b(G1192), .O(G1268) );

  xor2  gate1933(.a(G1192), .b(G1096), .O(gate460inter0));
  nand2 gate1934(.a(gate460inter0), .b(s_198), .O(gate460inter1));
  and2  gate1935(.a(G1192), .b(G1096), .O(gate460inter2));
  inv1  gate1936(.a(s_198), .O(gate460inter3));
  inv1  gate1937(.a(s_199), .O(gate460inter4));
  nand2 gate1938(.a(gate460inter4), .b(gate460inter3), .O(gate460inter5));
  nor2  gate1939(.a(gate460inter5), .b(gate460inter2), .O(gate460inter6));
  inv1  gate1940(.a(G1096), .O(gate460inter7));
  inv1  gate1941(.a(G1192), .O(gate460inter8));
  nand2 gate1942(.a(gate460inter8), .b(gate460inter7), .O(gate460inter9));
  nand2 gate1943(.a(s_199), .b(gate460inter3), .O(gate460inter10));
  nor2  gate1944(.a(gate460inter10), .b(gate460inter9), .O(gate460inter11));
  nor2  gate1945(.a(gate460inter11), .b(gate460inter6), .O(gate460inter12));
  nand2 gate1946(.a(gate460inter12), .b(gate460inter1), .O(G1269));
nand2 gate461( .a(G22), .b(G1195), .O(G1270) );
nand2 gate462( .a(G1099), .b(G1195), .O(G1271) );
nand2 gate463( .a(G23), .b(G1198), .O(G1272) );

  xor2  gate2311(.a(G1198), .b(G1102), .O(gate464inter0));
  nand2 gate2312(.a(gate464inter0), .b(s_252), .O(gate464inter1));
  and2  gate2313(.a(G1198), .b(G1102), .O(gate464inter2));
  inv1  gate2314(.a(s_252), .O(gate464inter3));
  inv1  gate2315(.a(s_253), .O(gate464inter4));
  nand2 gate2316(.a(gate464inter4), .b(gate464inter3), .O(gate464inter5));
  nor2  gate2317(.a(gate464inter5), .b(gate464inter2), .O(gate464inter6));
  inv1  gate2318(.a(G1102), .O(gate464inter7));
  inv1  gate2319(.a(G1198), .O(gate464inter8));
  nand2 gate2320(.a(gate464inter8), .b(gate464inter7), .O(gate464inter9));
  nand2 gate2321(.a(s_253), .b(gate464inter3), .O(gate464inter10));
  nor2  gate2322(.a(gate464inter10), .b(gate464inter9), .O(gate464inter11));
  nor2  gate2323(.a(gate464inter11), .b(gate464inter6), .O(gate464inter12));
  nand2 gate2324(.a(gate464inter12), .b(gate464inter1), .O(G1273));
nand2 gate465( .a(G24), .b(G1201), .O(G1274) );
nand2 gate466( .a(G1105), .b(G1201), .O(G1275) );

  xor2  gate1345(.a(G1204), .b(G25), .O(gate467inter0));
  nand2 gate1346(.a(gate467inter0), .b(s_114), .O(gate467inter1));
  and2  gate1347(.a(G1204), .b(G25), .O(gate467inter2));
  inv1  gate1348(.a(s_114), .O(gate467inter3));
  inv1  gate1349(.a(s_115), .O(gate467inter4));
  nand2 gate1350(.a(gate467inter4), .b(gate467inter3), .O(gate467inter5));
  nor2  gate1351(.a(gate467inter5), .b(gate467inter2), .O(gate467inter6));
  inv1  gate1352(.a(G25), .O(gate467inter7));
  inv1  gate1353(.a(G1204), .O(gate467inter8));
  nand2 gate1354(.a(gate467inter8), .b(gate467inter7), .O(gate467inter9));
  nand2 gate1355(.a(s_115), .b(gate467inter3), .O(gate467inter10));
  nor2  gate1356(.a(gate467inter10), .b(gate467inter9), .O(gate467inter11));
  nor2  gate1357(.a(gate467inter11), .b(gate467inter6), .O(gate467inter12));
  nand2 gate1358(.a(gate467inter12), .b(gate467inter1), .O(G1276));

  xor2  gate2297(.a(G1204), .b(G1108), .O(gate468inter0));
  nand2 gate2298(.a(gate468inter0), .b(s_250), .O(gate468inter1));
  and2  gate2299(.a(G1204), .b(G1108), .O(gate468inter2));
  inv1  gate2300(.a(s_250), .O(gate468inter3));
  inv1  gate2301(.a(s_251), .O(gate468inter4));
  nand2 gate2302(.a(gate468inter4), .b(gate468inter3), .O(gate468inter5));
  nor2  gate2303(.a(gate468inter5), .b(gate468inter2), .O(gate468inter6));
  inv1  gate2304(.a(G1108), .O(gate468inter7));
  inv1  gate2305(.a(G1204), .O(gate468inter8));
  nand2 gate2306(.a(gate468inter8), .b(gate468inter7), .O(gate468inter9));
  nand2 gate2307(.a(s_251), .b(gate468inter3), .O(gate468inter10));
  nor2  gate2308(.a(gate468inter10), .b(gate468inter9), .O(gate468inter11));
  nor2  gate2309(.a(gate468inter11), .b(gate468inter6), .O(gate468inter12));
  nand2 gate2310(.a(gate468inter12), .b(gate468inter1), .O(G1277));
nand2 gate469( .a(G26), .b(G1207), .O(G1278) );

  xor2  gate2549(.a(G1207), .b(G1111), .O(gate470inter0));
  nand2 gate2550(.a(gate470inter0), .b(s_286), .O(gate470inter1));
  and2  gate2551(.a(G1207), .b(G1111), .O(gate470inter2));
  inv1  gate2552(.a(s_286), .O(gate470inter3));
  inv1  gate2553(.a(s_287), .O(gate470inter4));
  nand2 gate2554(.a(gate470inter4), .b(gate470inter3), .O(gate470inter5));
  nor2  gate2555(.a(gate470inter5), .b(gate470inter2), .O(gate470inter6));
  inv1  gate2556(.a(G1111), .O(gate470inter7));
  inv1  gate2557(.a(G1207), .O(gate470inter8));
  nand2 gate2558(.a(gate470inter8), .b(gate470inter7), .O(gate470inter9));
  nand2 gate2559(.a(s_287), .b(gate470inter3), .O(gate470inter10));
  nor2  gate2560(.a(gate470inter10), .b(gate470inter9), .O(gate470inter11));
  nor2  gate2561(.a(gate470inter11), .b(gate470inter6), .O(gate470inter12));
  nand2 gate2562(.a(gate470inter12), .b(gate470inter1), .O(G1279));

  xor2  gate659(.a(G1210), .b(G27), .O(gate471inter0));
  nand2 gate660(.a(gate471inter0), .b(s_16), .O(gate471inter1));
  and2  gate661(.a(G1210), .b(G27), .O(gate471inter2));
  inv1  gate662(.a(s_16), .O(gate471inter3));
  inv1  gate663(.a(s_17), .O(gate471inter4));
  nand2 gate664(.a(gate471inter4), .b(gate471inter3), .O(gate471inter5));
  nor2  gate665(.a(gate471inter5), .b(gate471inter2), .O(gate471inter6));
  inv1  gate666(.a(G27), .O(gate471inter7));
  inv1  gate667(.a(G1210), .O(gate471inter8));
  nand2 gate668(.a(gate471inter8), .b(gate471inter7), .O(gate471inter9));
  nand2 gate669(.a(s_17), .b(gate471inter3), .O(gate471inter10));
  nor2  gate670(.a(gate471inter10), .b(gate471inter9), .O(gate471inter11));
  nor2  gate671(.a(gate471inter11), .b(gate471inter6), .O(gate471inter12));
  nand2 gate672(.a(gate471inter12), .b(gate471inter1), .O(G1280));
nand2 gate472( .a(G1114), .b(G1210), .O(G1281) );
nand2 gate473( .a(G28), .b(G1213), .O(G1282) );
nand2 gate474( .a(G1117), .b(G1213), .O(G1283) );
nand2 gate475( .a(G29), .b(G1216), .O(G1284) );
nand2 gate476( .a(G1120), .b(G1216), .O(G1285) );
nand2 gate477( .a(G30), .b(G1219), .O(G1286) );
nand2 gate478( .a(G1123), .b(G1219), .O(G1287) );
nand2 gate479( .a(G31), .b(G1222), .O(G1288) );

  xor2  gate1163(.a(G1222), .b(G1126), .O(gate480inter0));
  nand2 gate1164(.a(gate480inter0), .b(s_88), .O(gate480inter1));
  and2  gate1165(.a(G1222), .b(G1126), .O(gate480inter2));
  inv1  gate1166(.a(s_88), .O(gate480inter3));
  inv1  gate1167(.a(s_89), .O(gate480inter4));
  nand2 gate1168(.a(gate480inter4), .b(gate480inter3), .O(gate480inter5));
  nor2  gate1169(.a(gate480inter5), .b(gate480inter2), .O(gate480inter6));
  inv1  gate1170(.a(G1126), .O(gate480inter7));
  inv1  gate1171(.a(G1222), .O(gate480inter8));
  nand2 gate1172(.a(gate480inter8), .b(gate480inter7), .O(gate480inter9));
  nand2 gate1173(.a(s_89), .b(gate480inter3), .O(gate480inter10));
  nor2  gate1174(.a(gate480inter10), .b(gate480inter9), .O(gate480inter11));
  nor2  gate1175(.a(gate480inter11), .b(gate480inter6), .O(gate480inter12));
  nand2 gate1176(.a(gate480inter12), .b(gate480inter1), .O(G1289));
nand2 gate481( .a(G32), .b(G1225), .O(G1290) );

  xor2  gate953(.a(G1225), .b(G1129), .O(gate482inter0));
  nand2 gate954(.a(gate482inter0), .b(s_58), .O(gate482inter1));
  and2  gate955(.a(G1225), .b(G1129), .O(gate482inter2));
  inv1  gate956(.a(s_58), .O(gate482inter3));
  inv1  gate957(.a(s_59), .O(gate482inter4));
  nand2 gate958(.a(gate482inter4), .b(gate482inter3), .O(gate482inter5));
  nor2  gate959(.a(gate482inter5), .b(gate482inter2), .O(gate482inter6));
  inv1  gate960(.a(G1129), .O(gate482inter7));
  inv1  gate961(.a(G1225), .O(gate482inter8));
  nand2 gate962(.a(gate482inter8), .b(gate482inter7), .O(gate482inter9));
  nand2 gate963(.a(s_59), .b(gate482inter3), .O(gate482inter10));
  nor2  gate964(.a(gate482inter10), .b(gate482inter9), .O(gate482inter11));
  nor2  gate965(.a(gate482inter11), .b(gate482inter6), .O(gate482inter12));
  nand2 gate966(.a(gate482inter12), .b(gate482inter1), .O(G1291));

  xor2  gate1709(.a(G1229), .b(G1228), .O(gate483inter0));
  nand2 gate1710(.a(gate483inter0), .b(s_166), .O(gate483inter1));
  and2  gate1711(.a(G1229), .b(G1228), .O(gate483inter2));
  inv1  gate1712(.a(s_166), .O(gate483inter3));
  inv1  gate1713(.a(s_167), .O(gate483inter4));
  nand2 gate1714(.a(gate483inter4), .b(gate483inter3), .O(gate483inter5));
  nor2  gate1715(.a(gate483inter5), .b(gate483inter2), .O(gate483inter6));
  inv1  gate1716(.a(G1228), .O(gate483inter7));
  inv1  gate1717(.a(G1229), .O(gate483inter8));
  nand2 gate1718(.a(gate483inter8), .b(gate483inter7), .O(gate483inter9));
  nand2 gate1719(.a(s_167), .b(gate483inter3), .O(gate483inter10));
  nor2  gate1720(.a(gate483inter10), .b(gate483inter9), .O(gate483inter11));
  nor2  gate1721(.a(gate483inter11), .b(gate483inter6), .O(gate483inter12));
  nand2 gate1722(.a(gate483inter12), .b(gate483inter1), .O(G1292));
nand2 gate484( .a(G1230), .b(G1231), .O(G1293) );

  xor2  gate1065(.a(G1233), .b(G1232), .O(gate485inter0));
  nand2 gate1066(.a(gate485inter0), .b(s_74), .O(gate485inter1));
  and2  gate1067(.a(G1233), .b(G1232), .O(gate485inter2));
  inv1  gate1068(.a(s_74), .O(gate485inter3));
  inv1  gate1069(.a(s_75), .O(gate485inter4));
  nand2 gate1070(.a(gate485inter4), .b(gate485inter3), .O(gate485inter5));
  nor2  gate1071(.a(gate485inter5), .b(gate485inter2), .O(gate485inter6));
  inv1  gate1072(.a(G1232), .O(gate485inter7));
  inv1  gate1073(.a(G1233), .O(gate485inter8));
  nand2 gate1074(.a(gate485inter8), .b(gate485inter7), .O(gate485inter9));
  nand2 gate1075(.a(s_75), .b(gate485inter3), .O(gate485inter10));
  nor2  gate1076(.a(gate485inter10), .b(gate485inter9), .O(gate485inter11));
  nor2  gate1077(.a(gate485inter11), .b(gate485inter6), .O(gate485inter12));
  nand2 gate1078(.a(gate485inter12), .b(gate485inter1), .O(G1294));
nand2 gate486( .a(G1234), .b(G1235), .O(G1295) );
nand2 gate487( .a(G1236), .b(G1237), .O(G1296) );
nand2 gate488( .a(G1238), .b(G1239), .O(G1297) );
nand2 gate489( .a(G1240), .b(G1241), .O(G1298) );

  xor2  gate2619(.a(G1243), .b(G1242), .O(gate490inter0));
  nand2 gate2620(.a(gate490inter0), .b(s_296), .O(gate490inter1));
  and2  gate2621(.a(G1243), .b(G1242), .O(gate490inter2));
  inv1  gate2622(.a(s_296), .O(gate490inter3));
  inv1  gate2623(.a(s_297), .O(gate490inter4));
  nand2 gate2624(.a(gate490inter4), .b(gate490inter3), .O(gate490inter5));
  nor2  gate2625(.a(gate490inter5), .b(gate490inter2), .O(gate490inter6));
  inv1  gate2626(.a(G1242), .O(gate490inter7));
  inv1  gate2627(.a(G1243), .O(gate490inter8));
  nand2 gate2628(.a(gate490inter8), .b(gate490inter7), .O(gate490inter9));
  nand2 gate2629(.a(s_297), .b(gate490inter3), .O(gate490inter10));
  nor2  gate2630(.a(gate490inter10), .b(gate490inter9), .O(gate490inter11));
  nor2  gate2631(.a(gate490inter11), .b(gate490inter6), .O(gate490inter12));
  nand2 gate2632(.a(gate490inter12), .b(gate490inter1), .O(G1299));
nand2 gate491( .a(G1244), .b(G1245), .O(G1300) );

  xor2  gate2745(.a(G1247), .b(G1246), .O(gate492inter0));
  nand2 gate2746(.a(gate492inter0), .b(s_314), .O(gate492inter1));
  and2  gate2747(.a(G1247), .b(G1246), .O(gate492inter2));
  inv1  gate2748(.a(s_314), .O(gate492inter3));
  inv1  gate2749(.a(s_315), .O(gate492inter4));
  nand2 gate2750(.a(gate492inter4), .b(gate492inter3), .O(gate492inter5));
  nor2  gate2751(.a(gate492inter5), .b(gate492inter2), .O(gate492inter6));
  inv1  gate2752(.a(G1246), .O(gate492inter7));
  inv1  gate2753(.a(G1247), .O(gate492inter8));
  nand2 gate2754(.a(gate492inter8), .b(gate492inter7), .O(gate492inter9));
  nand2 gate2755(.a(s_315), .b(gate492inter3), .O(gate492inter10));
  nor2  gate2756(.a(gate492inter10), .b(gate492inter9), .O(gate492inter11));
  nor2  gate2757(.a(gate492inter11), .b(gate492inter6), .O(gate492inter12));
  nand2 gate2758(.a(gate492inter12), .b(gate492inter1), .O(G1301));
nand2 gate493( .a(G1248), .b(G1249), .O(G1302) );

  xor2  gate1555(.a(G1251), .b(G1250), .O(gate494inter0));
  nand2 gate1556(.a(gate494inter0), .b(s_144), .O(gate494inter1));
  and2  gate1557(.a(G1251), .b(G1250), .O(gate494inter2));
  inv1  gate1558(.a(s_144), .O(gate494inter3));
  inv1  gate1559(.a(s_145), .O(gate494inter4));
  nand2 gate1560(.a(gate494inter4), .b(gate494inter3), .O(gate494inter5));
  nor2  gate1561(.a(gate494inter5), .b(gate494inter2), .O(gate494inter6));
  inv1  gate1562(.a(G1250), .O(gate494inter7));
  inv1  gate1563(.a(G1251), .O(gate494inter8));
  nand2 gate1564(.a(gate494inter8), .b(gate494inter7), .O(gate494inter9));
  nand2 gate1565(.a(s_145), .b(gate494inter3), .O(gate494inter10));
  nor2  gate1566(.a(gate494inter10), .b(gate494inter9), .O(gate494inter11));
  nor2  gate1567(.a(gate494inter11), .b(gate494inter6), .O(gate494inter12));
  nand2 gate1568(.a(gate494inter12), .b(gate494inter1), .O(G1303));
nand2 gate495( .a(G1252), .b(G1253), .O(G1304) );

  xor2  gate631(.a(G1255), .b(G1254), .O(gate496inter0));
  nand2 gate632(.a(gate496inter0), .b(s_12), .O(gate496inter1));
  and2  gate633(.a(G1255), .b(G1254), .O(gate496inter2));
  inv1  gate634(.a(s_12), .O(gate496inter3));
  inv1  gate635(.a(s_13), .O(gate496inter4));
  nand2 gate636(.a(gate496inter4), .b(gate496inter3), .O(gate496inter5));
  nor2  gate637(.a(gate496inter5), .b(gate496inter2), .O(gate496inter6));
  inv1  gate638(.a(G1254), .O(gate496inter7));
  inv1  gate639(.a(G1255), .O(gate496inter8));
  nand2 gate640(.a(gate496inter8), .b(gate496inter7), .O(gate496inter9));
  nand2 gate641(.a(s_13), .b(gate496inter3), .O(gate496inter10));
  nor2  gate642(.a(gate496inter10), .b(gate496inter9), .O(gate496inter11));
  nor2  gate643(.a(gate496inter11), .b(gate496inter6), .O(gate496inter12));
  nand2 gate644(.a(gate496inter12), .b(gate496inter1), .O(G1305));

  xor2  gate673(.a(G1257), .b(G1256), .O(gate497inter0));
  nand2 gate674(.a(gate497inter0), .b(s_18), .O(gate497inter1));
  and2  gate675(.a(G1257), .b(G1256), .O(gate497inter2));
  inv1  gate676(.a(s_18), .O(gate497inter3));
  inv1  gate677(.a(s_19), .O(gate497inter4));
  nand2 gate678(.a(gate497inter4), .b(gate497inter3), .O(gate497inter5));
  nor2  gate679(.a(gate497inter5), .b(gate497inter2), .O(gate497inter6));
  inv1  gate680(.a(G1256), .O(gate497inter7));
  inv1  gate681(.a(G1257), .O(gate497inter8));
  nand2 gate682(.a(gate497inter8), .b(gate497inter7), .O(gate497inter9));
  nand2 gate683(.a(s_19), .b(gate497inter3), .O(gate497inter10));
  nor2  gate684(.a(gate497inter10), .b(gate497inter9), .O(gate497inter11));
  nor2  gate685(.a(gate497inter11), .b(gate497inter6), .O(gate497inter12));
  nand2 gate686(.a(gate497inter12), .b(gate497inter1), .O(G1306));
nand2 gate498( .a(G1258), .b(G1259), .O(G1307) );

  xor2  gate2689(.a(G1261), .b(G1260), .O(gate499inter0));
  nand2 gate2690(.a(gate499inter0), .b(s_306), .O(gate499inter1));
  and2  gate2691(.a(G1261), .b(G1260), .O(gate499inter2));
  inv1  gate2692(.a(s_306), .O(gate499inter3));
  inv1  gate2693(.a(s_307), .O(gate499inter4));
  nand2 gate2694(.a(gate499inter4), .b(gate499inter3), .O(gate499inter5));
  nor2  gate2695(.a(gate499inter5), .b(gate499inter2), .O(gate499inter6));
  inv1  gate2696(.a(G1260), .O(gate499inter7));
  inv1  gate2697(.a(G1261), .O(gate499inter8));
  nand2 gate2698(.a(gate499inter8), .b(gate499inter7), .O(gate499inter9));
  nand2 gate2699(.a(s_307), .b(gate499inter3), .O(gate499inter10));
  nor2  gate2700(.a(gate499inter10), .b(gate499inter9), .O(gate499inter11));
  nor2  gate2701(.a(gate499inter11), .b(gate499inter6), .O(gate499inter12));
  nand2 gate2702(.a(gate499inter12), .b(gate499inter1), .O(G1308));
nand2 gate500( .a(G1262), .b(G1263), .O(G1309) );

  xor2  gate1835(.a(G1265), .b(G1264), .O(gate501inter0));
  nand2 gate1836(.a(gate501inter0), .b(s_184), .O(gate501inter1));
  and2  gate1837(.a(G1265), .b(G1264), .O(gate501inter2));
  inv1  gate1838(.a(s_184), .O(gate501inter3));
  inv1  gate1839(.a(s_185), .O(gate501inter4));
  nand2 gate1840(.a(gate501inter4), .b(gate501inter3), .O(gate501inter5));
  nor2  gate1841(.a(gate501inter5), .b(gate501inter2), .O(gate501inter6));
  inv1  gate1842(.a(G1264), .O(gate501inter7));
  inv1  gate1843(.a(G1265), .O(gate501inter8));
  nand2 gate1844(.a(gate501inter8), .b(gate501inter7), .O(gate501inter9));
  nand2 gate1845(.a(s_185), .b(gate501inter3), .O(gate501inter10));
  nor2  gate1846(.a(gate501inter10), .b(gate501inter9), .O(gate501inter11));
  nor2  gate1847(.a(gate501inter11), .b(gate501inter6), .O(gate501inter12));
  nand2 gate1848(.a(gate501inter12), .b(gate501inter1), .O(G1310));
nand2 gate502( .a(G1266), .b(G1267), .O(G1311) );
nand2 gate503( .a(G1268), .b(G1269), .O(G1312) );
nand2 gate504( .a(G1270), .b(G1271), .O(G1313) );
nand2 gate505( .a(G1272), .b(G1273), .O(G1314) );

  xor2  gate1583(.a(G1275), .b(G1274), .O(gate506inter0));
  nand2 gate1584(.a(gate506inter0), .b(s_148), .O(gate506inter1));
  and2  gate1585(.a(G1275), .b(G1274), .O(gate506inter2));
  inv1  gate1586(.a(s_148), .O(gate506inter3));
  inv1  gate1587(.a(s_149), .O(gate506inter4));
  nand2 gate1588(.a(gate506inter4), .b(gate506inter3), .O(gate506inter5));
  nor2  gate1589(.a(gate506inter5), .b(gate506inter2), .O(gate506inter6));
  inv1  gate1590(.a(G1274), .O(gate506inter7));
  inv1  gate1591(.a(G1275), .O(gate506inter8));
  nand2 gate1592(.a(gate506inter8), .b(gate506inter7), .O(gate506inter9));
  nand2 gate1593(.a(s_149), .b(gate506inter3), .O(gate506inter10));
  nor2  gate1594(.a(gate506inter10), .b(gate506inter9), .O(gate506inter11));
  nor2  gate1595(.a(gate506inter11), .b(gate506inter6), .O(gate506inter12));
  nand2 gate1596(.a(gate506inter12), .b(gate506inter1), .O(G1315));
nand2 gate507( .a(G1276), .b(G1277), .O(G1316) );
nand2 gate508( .a(G1278), .b(G1279), .O(G1317) );
nand2 gate509( .a(G1280), .b(G1281), .O(G1318) );

  xor2  gate1373(.a(G1283), .b(G1282), .O(gate510inter0));
  nand2 gate1374(.a(gate510inter0), .b(s_118), .O(gate510inter1));
  and2  gate1375(.a(G1283), .b(G1282), .O(gate510inter2));
  inv1  gate1376(.a(s_118), .O(gate510inter3));
  inv1  gate1377(.a(s_119), .O(gate510inter4));
  nand2 gate1378(.a(gate510inter4), .b(gate510inter3), .O(gate510inter5));
  nor2  gate1379(.a(gate510inter5), .b(gate510inter2), .O(gate510inter6));
  inv1  gate1380(.a(G1282), .O(gate510inter7));
  inv1  gate1381(.a(G1283), .O(gate510inter8));
  nand2 gate1382(.a(gate510inter8), .b(gate510inter7), .O(gate510inter9));
  nand2 gate1383(.a(s_119), .b(gate510inter3), .O(gate510inter10));
  nor2  gate1384(.a(gate510inter10), .b(gate510inter9), .O(gate510inter11));
  nor2  gate1385(.a(gate510inter11), .b(gate510inter6), .O(gate510inter12));
  nand2 gate1386(.a(gate510inter12), .b(gate510inter1), .O(G1319));
nand2 gate511( .a(G1284), .b(G1285), .O(G1320) );
nand2 gate512( .a(G1286), .b(G1287), .O(G1321) );
nand2 gate513( .a(G1288), .b(G1289), .O(G1322) );

  xor2  gate869(.a(G1291), .b(G1290), .O(gate514inter0));
  nand2 gate870(.a(gate514inter0), .b(s_46), .O(gate514inter1));
  and2  gate871(.a(G1291), .b(G1290), .O(gate514inter2));
  inv1  gate872(.a(s_46), .O(gate514inter3));
  inv1  gate873(.a(s_47), .O(gate514inter4));
  nand2 gate874(.a(gate514inter4), .b(gate514inter3), .O(gate514inter5));
  nor2  gate875(.a(gate514inter5), .b(gate514inter2), .O(gate514inter6));
  inv1  gate876(.a(G1290), .O(gate514inter7));
  inv1  gate877(.a(G1291), .O(gate514inter8));
  nand2 gate878(.a(gate514inter8), .b(gate514inter7), .O(gate514inter9));
  nand2 gate879(.a(s_47), .b(gate514inter3), .O(gate514inter10));
  nor2  gate880(.a(gate514inter10), .b(gate514inter9), .O(gate514inter11));
  nor2  gate881(.a(gate514inter11), .b(gate514inter6), .O(gate514inter12));
  nand2 gate882(.a(gate514inter12), .b(gate514inter1), .O(G1323));
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule