module c499 (N1,N5,N9,N13,N17,N21,N25,N29,N33,N37,
             N41,N45,N49,N53,N57,N61,N65,N69,N73,N77,
             N81,N85,N89,N93,N97,N101,N105,N109,N113,N117,
             N121,N125,N129,N130,N131,N132,N133,N134,N135,N136,
             N137,N724,N725,N726,N727,N728,N729,N730,N731,N732,
             N733,N734,N735,N736,N737,N738,N739,N740,N741,N742,
             N743,N744,N745,N746,N747,N748,N749,N750,N751,N752,
             N753,N754,N755);

input N1,N5,N9,N13,N17,N21,N25,N29,N33,N37,
      N41,N45,N49,N53,N57,N61,N65,N69,N73,N77,
      N81,N85,N89,N93,N97,N101,N105,N109,N113,N117,
      N121,N125,N129,N130,N131,N132,N133,N134,N135,N136,
      N137;//RE__PI;

input s_0,s_1;//RE__ALLOW(00,01,10,11);
input s_2,s_3;//RE__ALLOW(00,01,10,11);
input s_4,s_5;//RE__ALLOW(00,01,10,11);
input s_6,s_7;//RE__ALLOW(00,01,10,11);
input s_8,s_9;//RE__ALLOW(00,01,10,11);
input s_10,s_11;//RE__ALLOW(00,01,10,11);
input s_12,s_13;//RE__ALLOW(00,01,10,11);
input s_14,s_15;//RE__ALLOW(00,01,10,11);
input s_16,s_17;//RE__ALLOW(00,01,10,11);
input s_18,s_19;//RE__ALLOW(00,01,10,11);
input s_20,s_21;//RE__ALLOW(00,01,10,11);
output N724,N725,N726,N727,N728,N729,N730,N731,N732,N733,
       N734,N735,N736,N737,N738,N739,N740,N741,N742,N743,
       N744,N745,N746,N747,N748,N749,N750,N751,N752,N753,
       N754,N755;

wire N250,N251,N252,N253,N254,N255,N256,N257,N258,N259,
     N260,N261,N262,N263,N264,N265,N266,N267,N268,N269,
     N270,N271,N272,N273,N274,N275,N276,N277,N278,N279,
     N280,N281,N282,N283,N284,N285,N286,N287,N288,N289,
     N290,N293,N296,N299,N302,N305,N308,N311,N314,N315,
     N316,N317,N318,N319,N320,N321,N338,N339,N340,N341,
     N342,N343,N344,N345,N346,N347,N348,N349,N350,N351,
     N352,N353,N354,N367,N380,N393,N406,N419,N432,N445,
     N554,N555,N556,N557,N558,N559,N560,N561,N562,N563,
     N564,N565,N566,N567,N568,N569,N570,N571,N572,N573,
     N574,N575,N576,N577,N578,N579,N580,N581,N582,N583,
     N584,N585,N586,N587,N588,N589,N590,N591,N592,N593,
     N594,N595,N596,N597,N598,N599,N600,N601,N602,N607,
     N620,N625,N630,N635,N640,N645,N650,N655,N692,N693,
     N694,N695,N696,N697,N698,N699,N700,N701,N702,N703,
     N704,N705,N706,N707,N708,N709,N710,N711,N712,N713,
     N714,N715,N716,N717,N718,N719,N720,N721,N722,N723, gate185inter0, gate185inter1, gate185inter2, gate185inter3, gate185inter4, gate185inter5, gate185inter6, gate185inter7, gate185inter8, gate185inter9, gate185inter10, gate185inter11, gate185inter12, gate41inter0, gate41inter1, gate41inter2, gate41inter3, gate41inter4, gate41inter5, gate41inter6, gate41inter7, gate41inter8, gate41inter9, gate41inter10, gate41inter11, gate41inter12, gate55inter0, gate55inter1, gate55inter2, gate55inter3, gate55inter4, gate55inter5, gate55inter6, gate55inter7, gate55inter8, gate55inter9, gate55inter10, gate55inter11, gate55inter12, gate5inter0, gate5inter1, gate5inter2, gate5inter3, gate5inter4, gate5inter5, gate5inter6, gate5inter7, gate5inter8, gate5inter9, gate5inter10, gate5inter11, gate5inter12, gate65inter0, gate65inter1, gate65inter2, gate65inter3, gate65inter4, gate65inter5, gate65inter6, gate65inter7, gate65inter8, gate65inter9, gate65inter10, gate65inter11, gate65inter12, gate29inter0, gate29inter1, gate29inter2, gate29inter3, gate29inter4, gate29inter5, gate29inter6, gate29inter7, gate29inter8, gate29inter9, gate29inter10, gate29inter11, gate29inter12, gate173inter0, gate173inter1, gate173inter2, gate173inter3, gate173inter4, gate173inter5, gate173inter6, gate173inter7, gate173inter8, gate173inter9, gate173inter10, gate173inter11, gate173inter12, gate48inter0, gate48inter1, gate48inter2, gate48inter3, gate48inter4, gate48inter5, gate48inter6, gate48inter7, gate48inter8, gate48inter9, gate48inter10, gate48inter11, gate48inter12, gate177inter0, gate177inter1, gate177inter2, gate177inter3, gate177inter4, gate177inter5, gate177inter6, gate177inter7, gate177inter8, gate177inter9, gate177inter10, gate177inter11, gate177inter12, gate6inter0, gate6inter1, gate6inter2, gate6inter3, gate6inter4, gate6inter5, gate6inter6, gate6inter7, gate6inter8, gate6inter9, gate6inter10, gate6inter11, gate6inter12, gate3inter0, gate3inter1, gate3inter2, gate3inter3, gate3inter4, gate3inter5, gate3inter6, gate3inter7, gate3inter8, gate3inter9, gate3inter10, gate3inter11, gate3inter12;



xor2 gate1( .a(N1), .b(N5), .O(N250) );
xor2 gate2( .a(N9), .b(N13), .O(N251) );

  xor2  gate343(.a(N21), .b(N17), .O(gate3inter0));
  nand2 gate344(.a(gate3inter0), .b(s_20), .O(gate3inter1));
  and2  gate345(.a(N21), .b(N17), .O(gate3inter2));
  inv1  gate346(.a(s_20), .O(gate3inter3));
  inv1  gate347(.a(s_21), .O(gate3inter4));
  nand2 gate348(.a(gate3inter4), .b(gate3inter3), .O(gate3inter5));
  nor2  gate349(.a(gate3inter5), .b(gate3inter2), .O(gate3inter6));
  inv1  gate350(.a(N17), .O(gate3inter7));
  inv1  gate351(.a(N21), .O(gate3inter8));
  nand2 gate352(.a(gate3inter8), .b(gate3inter7), .O(gate3inter9));
  nand2 gate353(.a(s_21), .b(gate3inter3), .O(gate3inter10));
  nor2  gate354(.a(gate3inter10), .b(gate3inter9), .O(gate3inter11));
  nor2  gate355(.a(gate3inter11), .b(gate3inter6), .O(gate3inter12));
  nand2 gate356(.a(gate3inter12), .b(gate3inter1), .O(N252));
xor2 gate4( .a(N25), .b(N29), .O(N253) );

  xor2  gate245(.a(N37), .b(N33), .O(gate5inter0));
  nand2 gate246(.a(gate5inter0), .b(s_6), .O(gate5inter1));
  and2  gate247(.a(N37), .b(N33), .O(gate5inter2));
  inv1  gate248(.a(s_6), .O(gate5inter3));
  inv1  gate249(.a(s_7), .O(gate5inter4));
  nand2 gate250(.a(gate5inter4), .b(gate5inter3), .O(gate5inter5));
  nor2  gate251(.a(gate5inter5), .b(gate5inter2), .O(gate5inter6));
  inv1  gate252(.a(N33), .O(gate5inter7));
  inv1  gate253(.a(N37), .O(gate5inter8));
  nand2 gate254(.a(gate5inter8), .b(gate5inter7), .O(gate5inter9));
  nand2 gate255(.a(s_7), .b(gate5inter3), .O(gate5inter10));
  nor2  gate256(.a(gate5inter10), .b(gate5inter9), .O(gate5inter11));
  nor2  gate257(.a(gate5inter11), .b(gate5inter6), .O(gate5inter12));
  nand2 gate258(.a(gate5inter12), .b(gate5inter1), .O(N254));

  xor2  gate329(.a(N45), .b(N41), .O(gate6inter0));
  nand2 gate330(.a(gate6inter0), .b(s_18), .O(gate6inter1));
  and2  gate331(.a(N45), .b(N41), .O(gate6inter2));
  inv1  gate332(.a(s_18), .O(gate6inter3));
  inv1  gate333(.a(s_19), .O(gate6inter4));
  nand2 gate334(.a(gate6inter4), .b(gate6inter3), .O(gate6inter5));
  nor2  gate335(.a(gate6inter5), .b(gate6inter2), .O(gate6inter6));
  inv1  gate336(.a(N41), .O(gate6inter7));
  inv1  gate337(.a(N45), .O(gate6inter8));
  nand2 gate338(.a(gate6inter8), .b(gate6inter7), .O(gate6inter9));
  nand2 gate339(.a(s_19), .b(gate6inter3), .O(gate6inter10));
  nor2  gate340(.a(gate6inter10), .b(gate6inter9), .O(gate6inter11));
  nor2  gate341(.a(gate6inter11), .b(gate6inter6), .O(gate6inter12));
  nand2 gate342(.a(gate6inter12), .b(gate6inter1), .O(N255));
xor2 gate7( .a(N49), .b(N53), .O(N256) );
xor2 gate8( .a(N57), .b(N61), .O(N257) );
xor2 gate9( .a(N65), .b(N69), .O(N258) );
xor2 gate10( .a(N73), .b(N77), .O(N259) );
xor2 gate11( .a(N81), .b(N85), .O(N260) );
xor2 gate12( .a(N89), .b(N93), .O(N261) );
xor2 gate13( .a(N97), .b(N101), .O(N262) );
xor2 gate14( .a(N105), .b(N109), .O(N263) );
xor2 gate15( .a(N113), .b(N117), .O(N264) );
xor2 gate16( .a(N121), .b(N125), .O(N265) );
and2 gate17( .a(N129), .b(N137), .O(N266) );
and2 gate18( .a(N130), .b(N137), .O(N267) );
and2 gate19( .a(N131), .b(N137), .O(N268) );
and2 gate20( .a(N132), .b(N137), .O(N269) );
and2 gate21( .a(N133), .b(N137), .O(N270) );
and2 gate22( .a(N134), .b(N137), .O(N271) );
and2 gate23( .a(N135), .b(N137), .O(N272) );
and2 gate24( .a(N136), .b(N137), .O(N273) );
xor2 gate25( .a(N1), .b(N17), .O(N274) );
xor2 gate26( .a(N33), .b(N49), .O(N275) );
xor2 gate27( .a(N5), .b(N21), .O(N276) );
xor2 gate28( .a(N37), .b(N53), .O(N277) );

  xor2  gate273(.a(N25), .b(N9), .O(gate29inter0));
  nand2 gate274(.a(gate29inter0), .b(s_10), .O(gate29inter1));
  and2  gate275(.a(N25), .b(N9), .O(gate29inter2));
  inv1  gate276(.a(s_10), .O(gate29inter3));
  inv1  gate277(.a(s_11), .O(gate29inter4));
  nand2 gate278(.a(gate29inter4), .b(gate29inter3), .O(gate29inter5));
  nor2  gate279(.a(gate29inter5), .b(gate29inter2), .O(gate29inter6));
  inv1  gate280(.a(N9), .O(gate29inter7));
  inv1  gate281(.a(N25), .O(gate29inter8));
  nand2 gate282(.a(gate29inter8), .b(gate29inter7), .O(gate29inter9));
  nand2 gate283(.a(s_11), .b(gate29inter3), .O(gate29inter10));
  nor2  gate284(.a(gate29inter10), .b(gate29inter9), .O(gate29inter11));
  nor2  gate285(.a(gate29inter11), .b(gate29inter6), .O(gate29inter12));
  nand2 gate286(.a(gate29inter12), .b(gate29inter1), .O(N278));
xor2 gate30( .a(N41), .b(N57), .O(N279) );
xor2 gate31( .a(N13), .b(N29), .O(N280) );
xor2 gate32( .a(N45), .b(N61), .O(N281) );
xor2 gate33( .a(N65), .b(N81), .O(N282) );
xor2 gate34( .a(N97), .b(N113), .O(N283) );
xor2 gate35( .a(N69), .b(N85), .O(N284) );
xor2 gate36( .a(N101), .b(N117), .O(N285) );
xor2 gate37( .a(N73), .b(N89), .O(N286) );
xor2 gate38( .a(N105), .b(N121), .O(N287) );
xor2 gate39( .a(N77), .b(N93), .O(N288) );
xor2 gate40( .a(N109), .b(N125), .O(N289) );

  xor2  gate217(.a(N251), .b(N250), .O(gate41inter0));
  nand2 gate218(.a(gate41inter0), .b(s_2), .O(gate41inter1));
  and2  gate219(.a(N251), .b(N250), .O(gate41inter2));
  inv1  gate220(.a(s_2), .O(gate41inter3));
  inv1  gate221(.a(s_3), .O(gate41inter4));
  nand2 gate222(.a(gate41inter4), .b(gate41inter3), .O(gate41inter5));
  nor2  gate223(.a(gate41inter5), .b(gate41inter2), .O(gate41inter6));
  inv1  gate224(.a(N250), .O(gate41inter7));
  inv1  gate225(.a(N251), .O(gate41inter8));
  nand2 gate226(.a(gate41inter8), .b(gate41inter7), .O(gate41inter9));
  nand2 gate227(.a(s_3), .b(gate41inter3), .O(gate41inter10));
  nor2  gate228(.a(gate41inter10), .b(gate41inter9), .O(gate41inter11));
  nor2  gate229(.a(gate41inter11), .b(gate41inter6), .O(gate41inter12));
  nand2 gate230(.a(gate41inter12), .b(gate41inter1), .O(N290));
xor2 gate42( .a(N252), .b(N253), .O(N293) );
xor2 gate43( .a(N254), .b(N255), .O(N296) );
xor2 gate44( .a(N256), .b(N257), .O(N299) );
xor2 gate45( .a(N258), .b(N259), .O(N302) );
xor2 gate46( .a(N260), .b(N261), .O(N305) );
xor2 gate47( .a(N262), .b(N263), .O(N308) );

  xor2  gate301(.a(N265), .b(N264), .O(gate48inter0));
  nand2 gate302(.a(gate48inter0), .b(s_14), .O(gate48inter1));
  and2  gate303(.a(N265), .b(N264), .O(gate48inter2));
  inv1  gate304(.a(s_14), .O(gate48inter3));
  inv1  gate305(.a(s_15), .O(gate48inter4));
  nand2 gate306(.a(gate48inter4), .b(gate48inter3), .O(gate48inter5));
  nor2  gate307(.a(gate48inter5), .b(gate48inter2), .O(gate48inter6));
  inv1  gate308(.a(N264), .O(gate48inter7));
  inv1  gate309(.a(N265), .O(gate48inter8));
  nand2 gate310(.a(gate48inter8), .b(gate48inter7), .O(gate48inter9));
  nand2 gate311(.a(s_15), .b(gate48inter3), .O(gate48inter10));
  nor2  gate312(.a(gate48inter10), .b(gate48inter9), .O(gate48inter11));
  nor2  gate313(.a(gate48inter11), .b(gate48inter6), .O(gate48inter12));
  nand2 gate314(.a(gate48inter12), .b(gate48inter1), .O(N311));
xor2 gate49( .a(N274), .b(N275), .O(N314) );
xor2 gate50( .a(N276), .b(N277), .O(N315) );
xor2 gate51( .a(N278), .b(N279), .O(N316) );
xor2 gate52( .a(N280), .b(N281), .O(N317) );
xor2 gate53( .a(N282), .b(N283), .O(N318) );
xor2 gate54( .a(N284), .b(N285), .O(N319) );

  xor2  gate231(.a(N287), .b(N286), .O(gate55inter0));
  nand2 gate232(.a(gate55inter0), .b(s_4), .O(gate55inter1));
  and2  gate233(.a(N287), .b(N286), .O(gate55inter2));
  inv1  gate234(.a(s_4), .O(gate55inter3));
  inv1  gate235(.a(s_5), .O(gate55inter4));
  nand2 gate236(.a(gate55inter4), .b(gate55inter3), .O(gate55inter5));
  nor2  gate237(.a(gate55inter5), .b(gate55inter2), .O(gate55inter6));
  inv1  gate238(.a(N286), .O(gate55inter7));
  inv1  gate239(.a(N287), .O(gate55inter8));
  nand2 gate240(.a(gate55inter8), .b(gate55inter7), .O(gate55inter9));
  nand2 gate241(.a(s_5), .b(gate55inter3), .O(gate55inter10));
  nor2  gate242(.a(gate55inter10), .b(gate55inter9), .O(gate55inter11));
  nor2  gate243(.a(gate55inter11), .b(gate55inter6), .O(gate55inter12));
  nand2 gate244(.a(gate55inter12), .b(gate55inter1), .O(N320));
xor2 gate56( .a(N288), .b(N289), .O(N321) );
xor2 gate57( .a(N290), .b(N293), .O(N338) );
xor2 gate58( .a(N296), .b(N299), .O(N339) );
xor2 gate59( .a(N290), .b(N296), .O(N340) );
xor2 gate60( .a(N293), .b(N299), .O(N341) );
xor2 gate61( .a(N302), .b(N305), .O(N342) );
xor2 gate62( .a(N308), .b(N311), .O(N343) );
xor2 gate63( .a(N302), .b(N308), .O(N344) );
xor2 gate64( .a(N305), .b(N311), .O(N345) );

  xor2  gate259(.a(N342), .b(N266), .O(gate65inter0));
  nand2 gate260(.a(gate65inter0), .b(s_8), .O(gate65inter1));
  and2  gate261(.a(N342), .b(N266), .O(gate65inter2));
  inv1  gate262(.a(s_8), .O(gate65inter3));
  inv1  gate263(.a(s_9), .O(gate65inter4));
  nand2 gate264(.a(gate65inter4), .b(gate65inter3), .O(gate65inter5));
  nor2  gate265(.a(gate65inter5), .b(gate65inter2), .O(gate65inter6));
  inv1  gate266(.a(N266), .O(gate65inter7));
  inv1  gate267(.a(N342), .O(gate65inter8));
  nand2 gate268(.a(gate65inter8), .b(gate65inter7), .O(gate65inter9));
  nand2 gate269(.a(s_9), .b(gate65inter3), .O(gate65inter10));
  nor2  gate270(.a(gate65inter10), .b(gate65inter9), .O(gate65inter11));
  nor2  gate271(.a(gate65inter11), .b(gate65inter6), .O(gate65inter12));
  nand2 gate272(.a(gate65inter12), .b(gate65inter1), .O(N346));
xor2 gate66( .a(N267), .b(N343), .O(N347) );
xor2 gate67( .a(N268), .b(N344), .O(N348) );
xor2 gate68( .a(N269), .b(N345), .O(N349) );
xor2 gate69( .a(N270), .b(N338), .O(N350) );
xor2 gate70( .a(N271), .b(N339), .O(N351) );
xor2 gate71( .a(N272), .b(N340), .O(N352) );
xor2 gate72( .a(N273), .b(N341), .O(N353) );
xor2 gate73( .a(N314), .b(N346), .O(N354) );
xor2 gate74( .a(N315), .b(N347), .O(N367) );
xor2 gate75( .a(N316), .b(N348), .O(N380) );
xor2 gate76( .a(N317), .b(N349), .O(N393) );
xor2 gate77( .a(N318), .b(N350), .O(N406) );
xor2 gate78( .a(N319), .b(N351), .O(N419) );
xor2 gate79( .a(N320), .b(N352), .O(N432) );
xor2 gate80( .a(N321), .b(N353), .O(N445) );
inv1 gate81( .a(N354), .O(N554) );
inv1 gate82( .a(N367), .O(N555) );
inv1 gate83( .a(N380), .O(N556) );
inv1 gate84( .a(N354), .O(N557) );
inv1 gate85( .a(N367), .O(N558) );
inv1 gate86( .a(N393), .O(N559) );
inv1 gate87( .a(N354), .O(N560) );
inv1 gate88( .a(N380), .O(N561) );
inv1 gate89( .a(N393), .O(N562) );
inv1 gate90( .a(N367), .O(N563) );
inv1 gate91( .a(N380), .O(N564) );
inv1 gate92( .a(N393), .O(N565) );
inv1 gate93( .a(N419), .O(N566) );
inv1 gate94( .a(N445), .O(N567) );
inv1 gate95( .a(N419), .O(N568) );
inv1 gate96( .a(N432), .O(N569) );
inv1 gate97( .a(N406), .O(N570) );
inv1 gate98( .a(N445), .O(N571) );
inv1 gate99( .a(N406), .O(N572) );
inv1 gate100( .a(N432), .O(N573) );
inv1 gate101( .a(N406), .O(N574) );
inv1 gate102( .a(N419), .O(N575) );
inv1 gate103( .a(N432), .O(N576) );
inv1 gate104( .a(N406), .O(N577) );
inv1 gate105( .a(N419), .O(N578) );
inv1 gate106( .a(N445), .O(N579) );
inv1 gate107( .a(N406), .O(N580) );
inv1 gate108( .a(N432), .O(N581) );
inv1 gate109( .a(N445), .O(N582) );
inv1 gate110( .a(N419), .O(N583) );
inv1 gate111( .a(N432), .O(N584) );
inv1 gate112( .a(N445), .O(N585) );
inv1 gate113( .a(N367), .O(N586) );
inv1 gate114( .a(N393), .O(N587) );
inv1 gate115( .a(N367), .O(N588) );
inv1 gate116( .a(N380), .O(N589) );
inv1 gate117( .a(N354), .O(N590) );
inv1 gate118( .a(N393), .O(N591) );
inv1 gate119( .a(N354), .O(N592) );
inv1 gate120( .a(N380), .O(N593) );
and4 gate121( .a(N554), .b(N555), .c(N556), .d(N393), .O(N594) );
and4 gate122( .a(N557), .b(N558), .c(N380), .d(N559), .O(N595) );
and4 gate123( .a(N560), .b(N367), .c(N561), .d(N562), .O(N596) );
and4 gate124( .a(N354), .b(N563), .c(N564), .d(N565), .O(N597) );
and4 gate125( .a(N574), .b(N575), .c(N576), .d(N445), .O(N598) );
and4 gate126( .a(N577), .b(N578), .c(N432), .d(N579), .O(N599) );
and4 gate127( .a(N580), .b(N419), .c(N581), .d(N582), .O(N600) );
and4 gate128( .a(N406), .b(N583), .c(N584), .d(N585), .O(N601) );
or4 gate129( .a(N594), .b(N595), .c(N596), .d(N597), .O(N602) );
or4 gate130( .a(N598), .b(N599), .c(N600), .d(N601), .O(N607) );
and5 gate131( .a(N406), .b(N566), .c(N432), .d(N567), .e(N602), .O(N620) );
and5 gate132( .a(N406), .b(N568), .c(N569), .d(N445), .e(N602), .O(N625) );
and5 gate133( .a(N570), .b(N419), .c(N432), .d(N571), .e(N602), .O(N630) );
and5 gate134( .a(N572), .b(N419), .c(N573), .d(N445), .e(N602), .O(N635) );
and5 gate135( .a(N354), .b(N586), .c(N380), .d(N587), .e(N607), .O(N640) );
and5 gate136( .a(N354), .b(N588), .c(N589), .d(N393), .e(N607), .O(N645) );
and5 gate137( .a(N590), .b(N367), .c(N380), .d(N591), .e(N607), .O(N650) );
and5 gate138( .a(N592), .b(N367), .c(N593), .d(N393), .e(N607), .O(N655) );
and2 gate139( .a(N354), .b(N620), .O(N692) );
and2 gate140( .a(N367), .b(N620), .O(N693) );
and2 gate141( .a(N380), .b(N620), .O(N694) );
and2 gate142( .a(N393), .b(N620), .O(N695) );
and2 gate143( .a(N354), .b(N625), .O(N696) );
and2 gate144( .a(N367), .b(N625), .O(N697) );
and2 gate145( .a(N380), .b(N625), .O(N698) );
and2 gate146( .a(N393), .b(N625), .O(N699) );
and2 gate147( .a(N354), .b(N630), .O(N700) );
and2 gate148( .a(N367), .b(N630), .O(N701) );
and2 gate149( .a(N380), .b(N630), .O(N702) );
and2 gate150( .a(N393), .b(N630), .O(N703) );
and2 gate151( .a(N354), .b(N635), .O(N704) );
and2 gate152( .a(N367), .b(N635), .O(N705) );
and2 gate153( .a(N380), .b(N635), .O(N706) );
and2 gate154( .a(N393), .b(N635), .O(N707) );
and2 gate155( .a(N406), .b(N640), .O(N708) );
and2 gate156( .a(N419), .b(N640), .O(N709) );
and2 gate157( .a(N432), .b(N640), .O(N710) );
and2 gate158( .a(N445), .b(N640), .O(N711) );
and2 gate159( .a(N406), .b(N645), .O(N712) );
and2 gate160( .a(N419), .b(N645), .O(N713) );
and2 gate161( .a(N432), .b(N645), .O(N714) );
and2 gate162( .a(N445), .b(N645), .O(N715) );
and2 gate163( .a(N406), .b(N650), .O(N716) );
and2 gate164( .a(N419), .b(N650), .O(N717) );
and2 gate165( .a(N432), .b(N650), .O(N718) );
and2 gate166( .a(N445), .b(N650), .O(N719) );
and2 gate167( .a(N406), .b(N655), .O(N720) );
and2 gate168( .a(N419), .b(N655), .O(N721) );
and2 gate169( .a(N432), .b(N655), .O(N722) );
and2 gate170( .a(N445), .b(N655), .O(N723) );
xor2 gate171( .a(N1), .b(N692), .O(N724) );
xor2 gate172( .a(N5), .b(N693), .O(N725) );

  xor2  gate287(.a(N694), .b(N9), .O(gate173inter0));
  nand2 gate288(.a(gate173inter0), .b(s_12), .O(gate173inter1));
  and2  gate289(.a(N694), .b(N9), .O(gate173inter2));
  inv1  gate290(.a(s_12), .O(gate173inter3));
  inv1  gate291(.a(s_13), .O(gate173inter4));
  nand2 gate292(.a(gate173inter4), .b(gate173inter3), .O(gate173inter5));
  nor2  gate293(.a(gate173inter5), .b(gate173inter2), .O(gate173inter6));
  inv1  gate294(.a(N9), .O(gate173inter7));
  inv1  gate295(.a(N694), .O(gate173inter8));
  nand2 gate296(.a(gate173inter8), .b(gate173inter7), .O(gate173inter9));
  nand2 gate297(.a(s_13), .b(gate173inter3), .O(gate173inter10));
  nor2  gate298(.a(gate173inter10), .b(gate173inter9), .O(gate173inter11));
  nor2  gate299(.a(gate173inter11), .b(gate173inter6), .O(gate173inter12));
  nand2 gate300(.a(gate173inter12), .b(gate173inter1), .O(N726));
xor2 gate174( .a(N13), .b(N695), .O(N727) );
xor2 gate175( .a(N17), .b(N696), .O(N728) );
xor2 gate176( .a(N21), .b(N697), .O(N729) );

  xor2  gate315(.a(N698), .b(N25), .O(gate177inter0));
  nand2 gate316(.a(gate177inter0), .b(s_16), .O(gate177inter1));
  and2  gate317(.a(N698), .b(N25), .O(gate177inter2));
  inv1  gate318(.a(s_16), .O(gate177inter3));
  inv1  gate319(.a(s_17), .O(gate177inter4));
  nand2 gate320(.a(gate177inter4), .b(gate177inter3), .O(gate177inter5));
  nor2  gate321(.a(gate177inter5), .b(gate177inter2), .O(gate177inter6));
  inv1  gate322(.a(N25), .O(gate177inter7));
  inv1  gate323(.a(N698), .O(gate177inter8));
  nand2 gate324(.a(gate177inter8), .b(gate177inter7), .O(gate177inter9));
  nand2 gate325(.a(s_17), .b(gate177inter3), .O(gate177inter10));
  nor2  gate326(.a(gate177inter10), .b(gate177inter9), .O(gate177inter11));
  nor2  gate327(.a(gate177inter11), .b(gate177inter6), .O(gate177inter12));
  nand2 gate328(.a(gate177inter12), .b(gate177inter1), .O(N730));
xor2 gate178( .a(N29), .b(N699), .O(N731) );
xor2 gate179( .a(N33), .b(N700), .O(N732) );
xor2 gate180( .a(N37), .b(N701), .O(N733) );
xor2 gate181( .a(N41), .b(N702), .O(N734) );
xor2 gate182( .a(N45), .b(N703), .O(N735) );
xor2 gate183( .a(N49), .b(N704), .O(N736) );
xor2 gate184( .a(N53), .b(N705), .O(N737) );

  xor2  gate203(.a(N706), .b(N57), .O(gate185inter0));
  nand2 gate204(.a(gate185inter0), .b(s_0), .O(gate185inter1));
  and2  gate205(.a(N706), .b(N57), .O(gate185inter2));
  inv1  gate206(.a(s_0), .O(gate185inter3));
  inv1  gate207(.a(s_1), .O(gate185inter4));
  nand2 gate208(.a(gate185inter4), .b(gate185inter3), .O(gate185inter5));
  nor2  gate209(.a(gate185inter5), .b(gate185inter2), .O(gate185inter6));
  inv1  gate210(.a(N57), .O(gate185inter7));
  inv1  gate211(.a(N706), .O(gate185inter8));
  nand2 gate212(.a(gate185inter8), .b(gate185inter7), .O(gate185inter9));
  nand2 gate213(.a(s_1), .b(gate185inter3), .O(gate185inter10));
  nor2  gate214(.a(gate185inter10), .b(gate185inter9), .O(gate185inter11));
  nor2  gate215(.a(gate185inter11), .b(gate185inter6), .O(gate185inter12));
  nand2 gate216(.a(gate185inter12), .b(gate185inter1), .O(N738));
xor2 gate186( .a(N61), .b(N707), .O(N739) );
xor2 gate187( .a(N65), .b(N708), .O(N740) );
xor2 gate188( .a(N69), .b(N709), .O(N741) );
xor2 gate189( .a(N73), .b(N710), .O(N742) );
xor2 gate190( .a(N77), .b(N711), .O(N743) );
xor2 gate191( .a(N81), .b(N712), .O(N744) );
xor2 gate192( .a(N85), .b(N713), .O(N745) );
xor2 gate193( .a(N89), .b(N714), .O(N746) );
xor2 gate194( .a(N93), .b(N715), .O(N747) );
xor2 gate195( .a(N97), .b(N716), .O(N748) );
xor2 gate196( .a(N101), .b(N717), .O(N749) );
xor2 gate197( .a(N105), .b(N718), .O(N750) );
xor2 gate198( .a(N109), .b(N719), .O(N751) );
xor2 gate199( .a(N113), .b(N720), .O(N752) );
xor2 gate200( .a(N117), .b(N721), .O(N753) );
xor2 gate201( .a(N121), .b(N722), .O(N754) );
xor2 gate202( .a(N125), .b(N723), .O(N755) );

endmodule