module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);

input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;//RE__PI;

input s_0,s_1;//RE__ALLOW(00,01,10,11);
input s_2,s_3;//RE__ALLOW(00,01,10,11);
input s_4,s_5;//RE__ALLOW(00,01,10,11);
input s_6,s_7;//RE__ALLOW(00,01,10,11);
input s_8,s_9;//RE__ALLOW(00,01,10,11);
input s_10,s_11;//RE__ALLOW(00,01,10,11);
input s_12,s_13;//RE__ALLOW(00,01,10,11);
input s_14,s_15;//RE__ALLOW(00,01,10,11);
input s_16,s_17;//RE__ALLOW(00,01,10,11);
input s_18,s_19;//RE__ALLOW(00,01,10,11);
input s_20,s_21;//RE__ALLOW(00,01,10,11);
input s_22,s_23;//RE__ALLOW(00,01,10,11);
input s_24,s_25;//RE__ALLOW(00,01,10,11);
input s_26,s_27;//RE__ALLOW(00,01,10,11);
input s_28,s_29;//RE__ALLOW(00,01,10,11);
input s_30,s_31;//RE__ALLOW(00,01,10,11);
input s_32,s_33;//RE__ALLOW(00,01,10,11);
input s_34,s_35;//RE__ALLOW(00,01,10,11);
input s_36,s_37;//RE__ALLOW(00,01,10,11);
input s_38,s_39;//RE__ALLOW(00,01,10,11);
input s_40,s_41;//RE__ALLOW(00,01,10,11);
input s_42,s_43;//RE__ALLOW(00,01,10,11);
input s_44,s_45;//RE__ALLOW(00,01,10,11);
input s_46,s_47;//RE__ALLOW(00,01,10,11);
input s_48,s_49;//RE__ALLOW(00,01,10,11);
input s_50,s_51;//RE__ALLOW(00,01,10,11);
input s_52,s_53;//RE__ALLOW(00,01,10,11);
input s_54,s_55;//RE__ALLOW(00,01,10,11);
input s_56,s_57;//RE__ALLOW(00,01,10,11);
input s_58,s_59;//RE__ALLOW(00,01,10,11);
input s_60,s_61;//RE__ALLOW(00,01,10,11);
input s_62,s_63;//RE__ALLOW(00,01,10,11);
input s_64,s_65;//RE__ALLOW(00,01,10,11);
input s_66,s_67;//RE__ALLOW(00,01,10,11);
input s_68,s_69;//RE__ALLOW(00,01,10,11);
input s_70,s_71;//RE__ALLOW(00,01,10,11);
input s_72,s_73;//RE__ALLOW(00,01,10,11);
input s_74,s_75;//RE__ALLOW(00,01,10,11);
input s_76,s_77;//RE__ALLOW(00,01,10,11);
input s_78,s_79;//RE__ALLOW(00,01,10,11);
input s_80,s_81;//RE__ALLOW(00,01,10,11);
input s_82,s_83;//RE__ALLOW(00,01,10,11);
input s_84,s_85;//RE__ALLOW(00,01,10,11);
input s_86,s_87;//RE__ALLOW(00,01,10,11);
input s_88,s_89;//RE__ALLOW(00,01,10,11);
input s_90,s_91;//RE__ALLOW(00,01,10,11);
input s_92,s_93;//RE__ALLOW(00,01,10,11);
input s_94,s_95;//RE__ALLOW(00,01,10,11);
input s_96,s_97;//RE__ALLOW(00,01,10,11);
input s_98,s_99;//RE__ALLOW(00,01,10,11);
input s_100,s_101;//RE__ALLOW(00,01,10,11);
input s_102,s_103;//RE__ALLOW(00,01,10,11);
input s_104,s_105;//RE__ALLOW(00,01,10,11);
input s_106,s_107;//RE__ALLOW(00,01,10,11);
input s_108,s_109;//RE__ALLOW(00,01,10,11);
input s_110,s_111;//RE__ALLOW(00,01,10,11);
input s_112,s_113;//RE__ALLOW(00,01,10,11);
input s_114,s_115;//RE__ALLOW(00,01,10,11);
input s_116,s_117;//RE__ALLOW(00,01,10,11);
input s_118,s_119;//RE__ALLOW(00,01,10,11);
input s_120,s_121;//RE__ALLOW(00,01,10,11);
input s_122,s_123;//RE__ALLOW(00,01,10,11);
input s_124,s_125;//RE__ALLOW(00,01,10,11);
input s_126,s_127;//RE__ALLOW(00,01,10,11);
input s_128,s_129;//RE__ALLOW(00,01,10,11);
input s_130,s_131;//RE__ALLOW(00,01,10,11);
input s_132,s_133;//RE__ALLOW(00,01,10,11);
input s_134,s_135;//RE__ALLOW(00,01,10,11);
input s_136,s_137;//RE__ALLOW(00,01,10,11);
input s_138,s_139;//RE__ALLOW(00,01,10,11);
input s_140,s_141;//RE__ALLOW(00,01,10,11);
input s_142,s_143;//RE__ALLOW(00,01,10,11);
input s_144,s_145;//RE__ALLOW(00,01,10,11);
input s_146,s_147;//RE__ALLOW(00,01,10,11);
input s_148,s_149;//RE__ALLOW(00,01,10,11);
input s_150,s_151;//RE__ALLOW(00,01,10,11);
input s_152,s_153;//RE__ALLOW(00,01,10,11);
input s_154,s_155;//RE__ALLOW(00,01,10,11);
input s_156,s_157;//RE__ALLOW(00,01,10,11);
input s_158,s_159;//RE__ALLOW(00,01,10,11);
input s_160,s_161;//RE__ALLOW(00,01,10,11);
input s_162,s_163;//RE__ALLOW(00,01,10,11);
input s_164,s_165;//RE__ALLOW(00,01,10,11);
input s_166,s_167;//RE__ALLOW(00,01,10,11);
input s_168,s_169;//RE__ALLOW(00,01,10,11);
input s_170,s_171;//RE__ALLOW(00,01,10,11);
input s_172,s_173;//RE__ALLOW(00,01,10,11);
input s_174,s_175;//RE__ALLOW(00,01,10,11);
input s_176,s_177;//RE__ALLOW(00,01,10,11);
input s_178,s_179;//RE__ALLOW(00,01,10,11);
input s_180,s_181;//RE__ALLOW(00,01,10,11);
input s_182,s_183;//RE__ALLOW(00,01,10,11);
input s_184,s_185;//RE__ALLOW(00,01,10,11);
input s_186,s_187;//RE__ALLOW(00,01,10,11);
input s_188,s_189;//RE__ALLOW(00,01,10,11);
input s_190,s_191;//RE__ALLOW(00,01,10,11);
input s_192,s_193;//RE__ALLOW(00,01,10,11);
input s_194,s_195;//RE__ALLOW(00,01,10,11);
input s_196,s_197;//RE__ALLOW(00,01,10,11);
input s_198,s_199;//RE__ALLOW(00,01,10,11);
input s_200,s_201;//RE__ALLOW(00,01,10,11);
input s_202,s_203;//RE__ALLOW(00,01,10,11);
input s_204,s_205;//RE__ALLOW(00,01,10,11);
input s_206,s_207;//RE__ALLOW(00,01,10,11);
input s_208,s_209;//RE__ALLOW(00,01,10,11);
input s_210,s_211;//RE__ALLOW(00,01,10,11);
input s_212,s_213;//RE__ALLOW(00,01,10,11);
input s_214,s_215;//RE__ALLOW(00,01,10,11);
input s_216,s_217;//RE__ALLOW(00,01,10,11);
input s_218,s_219;//RE__ALLOW(00,01,10,11);
input s_220,s_221;//RE__ALLOW(00,01,10,11);
input s_222,s_223;//RE__ALLOW(00,01,10,11);
input s_224,s_225;//RE__ALLOW(00,01,10,11);
input s_226,s_227;//RE__ALLOW(00,01,10,11);
input s_228,s_229;//RE__ALLOW(00,01,10,11);
input s_230,s_231;//RE__ALLOW(00,01,10,11);
input s_232,s_233;//RE__ALLOW(00,01,10,11);
input s_234,s_235;//RE__ALLOW(00,01,10,11);
input s_236,s_237;//RE__ALLOW(00,01,10,11);
input s_238,s_239;//RE__ALLOW(00,01,10,11);
input s_240,s_241;//RE__ALLOW(00,01,10,11);
input s_242,s_243;//RE__ALLOW(00,01,10,11);
input s_244,s_245;//RE__ALLOW(00,01,10,11);
input s_246,s_247;//RE__ALLOW(00,01,10,11);
input s_248,s_249;//RE__ALLOW(00,01,10,11);
input s_250,s_251;//RE__ALLOW(00,01,10,11);
input s_252,s_253;//RE__ALLOW(00,01,10,11);
input s_254,s_255;//RE__ALLOW(00,01,10,11);
input s_256,s_257;//RE__ALLOW(00,01,10,11);
input s_258,s_259;//RE__ALLOW(00,01,10,11);
input s_260,s_261;//RE__ALLOW(00,01,10,11);
input s_262,s_263;//RE__ALLOW(00,01,10,11);
input s_264,s_265;//RE__ALLOW(00,01,10,11);
input s_266,s_267;//RE__ALLOW(00,01,10,11);
input s_268,s_269;//RE__ALLOW(00,01,10,11);
input s_270,s_271;//RE__ALLOW(00,01,10,11);
input s_272,s_273;//RE__ALLOW(00,01,10,11);
input s_274,s_275;//RE__ALLOW(00,01,10,11);
input s_276,s_277;//RE__ALLOW(00,01,10,11);
input s_278,s_279;//RE__ALLOW(00,01,10,11);
input s_280,s_281;//RE__ALLOW(00,01,10,11);
input s_282,s_283;//RE__ALLOW(00,01,10,11);
input s_284,s_285;//RE__ALLOW(00,01,10,11);
input s_286,s_287;//RE__ALLOW(00,01,10,11);
input s_288,s_289;//RE__ALLOW(00,01,10,11);
input s_290,s_291;//RE__ALLOW(00,01,10,11);
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;

  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate195inter0, gate195inter1, gate195inter2, gate195inter3, gate195inter4, gate195inter5, gate195inter6, gate195inter7, gate195inter8, gate195inter9, gate195inter10, gate195inter11, gate195inter12, gate84inter0, gate84inter1, gate84inter2, gate84inter3, gate84inter4, gate84inter5, gate84inter6, gate84inter7, gate84inter8, gate84inter9, gate84inter10, gate84inter11, gate84inter12, gate176inter0, gate176inter1, gate176inter2, gate176inter3, gate176inter4, gate176inter5, gate176inter6, gate176inter7, gate176inter8, gate176inter9, gate176inter10, gate176inter11, gate176inter12, gate242inter0, gate242inter1, gate242inter2, gate242inter3, gate242inter4, gate242inter5, gate242inter6, gate242inter7, gate242inter8, gate242inter9, gate242inter10, gate242inter11, gate242inter12, gate103inter0, gate103inter1, gate103inter2, gate103inter3, gate103inter4, gate103inter5, gate103inter6, gate103inter7, gate103inter8, gate103inter9, gate103inter10, gate103inter11, gate103inter12, gate197inter0, gate197inter1, gate197inter2, gate197inter3, gate197inter4, gate197inter5, gate197inter6, gate197inter7, gate197inter8, gate197inter9, gate197inter10, gate197inter11, gate197inter12, gate70inter0, gate70inter1, gate70inter2, gate70inter3, gate70inter4, gate70inter5, gate70inter6, gate70inter7, gate70inter8, gate70inter9, gate70inter10, gate70inter11, gate70inter12, gate144inter0, gate144inter1, gate144inter2, gate144inter3, gate144inter4, gate144inter5, gate144inter6, gate144inter7, gate144inter8, gate144inter9, gate144inter10, gate144inter11, gate144inter12, gate492inter0, gate492inter1, gate492inter2, gate492inter3, gate492inter4, gate492inter5, gate492inter6, gate492inter7, gate492inter8, gate492inter9, gate492inter10, gate492inter11, gate492inter12, gate173inter0, gate173inter1, gate173inter2, gate173inter3, gate173inter4, gate173inter5, gate173inter6, gate173inter7, gate173inter8, gate173inter9, gate173inter10, gate173inter11, gate173inter12, gate495inter0, gate495inter1, gate495inter2, gate495inter3, gate495inter4, gate495inter5, gate495inter6, gate495inter7, gate495inter8, gate495inter9, gate495inter10, gate495inter11, gate495inter12, gate291inter0, gate291inter1, gate291inter2, gate291inter3, gate291inter4, gate291inter5, gate291inter6, gate291inter7, gate291inter8, gate291inter9, gate291inter10, gate291inter11, gate291inter12, gate429inter0, gate429inter1, gate429inter2, gate429inter3, gate429inter4, gate429inter5, gate429inter6, gate429inter7, gate429inter8, gate429inter9, gate429inter10, gate429inter11, gate429inter12, gate292inter0, gate292inter1, gate292inter2, gate292inter3, gate292inter4, gate292inter5, gate292inter6, gate292inter7, gate292inter8, gate292inter9, gate292inter10, gate292inter11, gate292inter12, gate463inter0, gate463inter1, gate463inter2, gate463inter3, gate463inter4, gate463inter5, gate463inter6, gate463inter7, gate463inter8, gate463inter9, gate463inter10, gate463inter11, gate463inter12, gate267inter0, gate267inter1, gate267inter2, gate267inter3, gate267inter4, gate267inter5, gate267inter6, gate267inter7, gate267inter8, gate267inter9, gate267inter10, gate267inter11, gate267inter12, gate182inter0, gate182inter1, gate182inter2, gate182inter3, gate182inter4, gate182inter5, gate182inter6, gate182inter7, gate182inter8, gate182inter9, gate182inter10, gate182inter11, gate182inter12, gate127inter0, gate127inter1, gate127inter2, gate127inter3, gate127inter4, gate127inter5, gate127inter6, gate127inter7, gate127inter8, gate127inter9, gate127inter10, gate127inter11, gate127inter12, gate269inter0, gate269inter1, gate269inter2, gate269inter3, gate269inter4, gate269inter5, gate269inter6, gate269inter7, gate269inter8, gate269inter9, gate269inter10, gate269inter11, gate269inter12, gate110inter0, gate110inter1, gate110inter2, gate110inter3, gate110inter4, gate110inter5, gate110inter6, gate110inter7, gate110inter8, gate110inter9, gate110inter10, gate110inter11, gate110inter12, gate504inter0, gate504inter1, gate504inter2, gate504inter3, gate504inter4, gate504inter5, gate504inter6, gate504inter7, gate504inter8, gate504inter9, gate504inter10, gate504inter11, gate504inter12, gate172inter0, gate172inter1, gate172inter2, gate172inter3, gate172inter4, gate172inter5, gate172inter6, gate172inter7, gate172inter8, gate172inter9, gate172inter10, gate172inter11, gate172inter12, gate499inter0, gate499inter1, gate499inter2, gate499inter3, gate499inter4, gate499inter5, gate499inter6, gate499inter7, gate499inter8, gate499inter9, gate499inter10, gate499inter11, gate499inter12, gate177inter0, gate177inter1, gate177inter2, gate177inter3, gate177inter4, gate177inter5, gate177inter6, gate177inter7, gate177inter8, gate177inter9, gate177inter10, gate177inter11, gate177inter12, gate214inter0, gate214inter1, gate214inter2, gate214inter3, gate214inter4, gate214inter5, gate214inter6, gate214inter7, gate214inter8, gate214inter9, gate214inter10, gate214inter11, gate214inter12, gate198inter0, gate198inter1, gate198inter2, gate198inter3, gate198inter4, gate198inter5, gate198inter6, gate198inter7, gate198inter8, gate198inter9, gate198inter10, gate198inter11, gate198inter12, gate290inter0, gate290inter1, gate290inter2, gate290inter3, gate290inter4, gate290inter5, gate290inter6, gate290inter7, gate290inter8, gate290inter9, gate290inter10, gate290inter11, gate290inter12, gate53inter0, gate53inter1, gate53inter2, gate53inter3, gate53inter4, gate53inter5, gate53inter6, gate53inter7, gate53inter8, gate53inter9, gate53inter10, gate53inter11, gate53inter12, gate10inter0, gate10inter1, gate10inter2, gate10inter3, gate10inter4, gate10inter5, gate10inter6, gate10inter7, gate10inter8, gate10inter9, gate10inter10, gate10inter11, gate10inter12, gate67inter0, gate67inter1, gate67inter2, gate67inter3, gate67inter4, gate67inter5, gate67inter6, gate67inter7, gate67inter8, gate67inter9, gate67inter10, gate67inter11, gate67inter12, gate391inter0, gate391inter1, gate391inter2, gate391inter3, gate391inter4, gate391inter5, gate391inter6, gate391inter7, gate391inter8, gate391inter9, gate391inter10, gate391inter11, gate391inter12, gate410inter0, gate410inter1, gate410inter2, gate410inter3, gate410inter4, gate410inter5, gate410inter6, gate410inter7, gate410inter8, gate410inter9, gate410inter10, gate410inter11, gate410inter12, gate166inter0, gate166inter1, gate166inter2, gate166inter3, gate166inter4, gate166inter5, gate166inter6, gate166inter7, gate166inter8, gate166inter9, gate166inter10, gate166inter11, gate166inter12, gate258inter0, gate258inter1, gate258inter2, gate258inter3, gate258inter4, gate258inter5, gate258inter6, gate258inter7, gate258inter8, gate258inter9, gate258inter10, gate258inter11, gate258inter12, gate14inter0, gate14inter1, gate14inter2, gate14inter3, gate14inter4, gate14inter5, gate14inter6, gate14inter7, gate14inter8, gate14inter9, gate14inter10, gate14inter11, gate14inter12, gate238inter0, gate238inter1, gate238inter2, gate238inter3, gate238inter4, gate238inter5, gate238inter6, gate238inter7, gate238inter8, gate238inter9, gate238inter10, gate238inter11, gate238inter12, gate60inter0, gate60inter1, gate60inter2, gate60inter3, gate60inter4, gate60inter5, gate60inter6, gate60inter7, gate60inter8, gate60inter9, gate60inter10, gate60inter11, gate60inter12, gate206inter0, gate206inter1, gate206inter2, gate206inter3, gate206inter4, gate206inter5, gate206inter6, gate206inter7, gate206inter8, gate206inter9, gate206inter10, gate206inter11, gate206inter12, gate43inter0, gate43inter1, gate43inter2, gate43inter3, gate43inter4, gate43inter5, gate43inter6, gate43inter7, gate43inter8, gate43inter9, gate43inter10, gate43inter11, gate43inter12, gate396inter0, gate396inter1, gate396inter2, gate396inter3, gate396inter4, gate396inter5, gate396inter6, gate396inter7, gate396inter8, gate396inter9, gate396inter10, gate396inter11, gate396inter12, gate94inter0, gate94inter1, gate94inter2, gate94inter3, gate94inter4, gate94inter5, gate94inter6, gate94inter7, gate94inter8, gate94inter9, gate94inter10, gate94inter11, gate94inter12, gate237inter0, gate237inter1, gate237inter2, gate237inter3, gate237inter4, gate237inter5, gate237inter6, gate237inter7, gate237inter8, gate237inter9, gate237inter10, gate237inter11, gate237inter12, gate159inter0, gate159inter1, gate159inter2, gate159inter3, gate159inter4, gate159inter5, gate159inter6, gate159inter7, gate159inter8, gate159inter9, gate159inter10, gate159inter11, gate159inter12, gate403inter0, gate403inter1, gate403inter2, gate403inter3, gate403inter4, gate403inter5, gate403inter6, gate403inter7, gate403inter8, gate403inter9, gate403inter10, gate403inter11, gate403inter12, gate31inter0, gate31inter1, gate31inter2, gate31inter3, gate31inter4, gate31inter5, gate31inter6, gate31inter7, gate31inter8, gate31inter9, gate31inter10, gate31inter11, gate31inter12, gate249inter0, gate249inter1, gate249inter2, gate249inter3, gate249inter4, gate249inter5, gate249inter6, gate249inter7, gate249inter8, gate249inter9, gate249inter10, gate249inter11, gate249inter12, gate13inter0, gate13inter1, gate13inter2, gate13inter3, gate13inter4, gate13inter5, gate13inter6, gate13inter7, gate13inter8, gate13inter9, gate13inter10, gate13inter11, gate13inter12, gate419inter0, gate419inter1, gate419inter2, gate419inter3, gate419inter4, gate419inter5, gate419inter6, gate419inter7, gate419inter8, gate419inter9, gate419inter10, gate419inter11, gate419inter12, gate38inter0, gate38inter1, gate38inter2, gate38inter3, gate38inter4, gate38inter5, gate38inter6, gate38inter7, gate38inter8, gate38inter9, gate38inter10, gate38inter11, gate38inter12, gate41inter0, gate41inter1, gate41inter2, gate41inter3, gate41inter4, gate41inter5, gate41inter6, gate41inter7, gate41inter8, gate41inter9, gate41inter10, gate41inter11, gate41inter12, gate494inter0, gate494inter1, gate494inter2, gate494inter3, gate494inter4, gate494inter5, gate494inter6, gate494inter7, gate494inter8, gate494inter9, gate494inter10, gate494inter11, gate494inter12, gate295inter0, gate295inter1, gate295inter2, gate295inter3, gate295inter4, gate295inter5, gate295inter6, gate295inter7, gate295inter8, gate295inter9, gate295inter10, gate295inter11, gate295inter12, gate509inter0, gate509inter1, gate509inter2, gate509inter3, gate509inter4, gate509inter5, gate509inter6, gate509inter7, gate509inter8, gate509inter9, gate509inter10, gate509inter11, gate509inter12, gate404inter0, gate404inter1, gate404inter2, gate404inter3, gate404inter4, gate404inter5, gate404inter6, gate404inter7, gate404inter8, gate404inter9, gate404inter10, gate404inter11, gate404inter12, gate513inter0, gate513inter1, gate513inter2, gate513inter3, gate513inter4, gate513inter5, gate513inter6, gate513inter7, gate513inter8, gate513inter9, gate513inter10, gate513inter11, gate513inter12, gate293inter0, gate293inter1, gate293inter2, gate293inter3, gate293inter4, gate293inter5, gate293inter6, gate293inter7, gate293inter8, gate293inter9, gate293inter10, gate293inter11, gate293inter12, gate113inter0, gate113inter1, gate113inter2, gate113inter3, gate113inter4, gate113inter5, gate113inter6, gate113inter7, gate113inter8, gate113inter9, gate113inter10, gate113inter11, gate113inter12, gate274inter0, gate274inter1, gate274inter2, gate274inter3, gate274inter4, gate274inter5, gate274inter6, gate274inter7, gate274inter8, gate274inter9, gate274inter10, gate274inter11, gate274inter12, gate395inter0, gate395inter1, gate395inter2, gate395inter3, gate395inter4, gate395inter5, gate395inter6, gate395inter7, gate395inter8, gate395inter9, gate395inter10, gate395inter11, gate395inter12, gate392inter0, gate392inter1, gate392inter2, gate392inter3, gate392inter4, gate392inter5, gate392inter6, gate392inter7, gate392inter8, gate392inter9, gate392inter10, gate392inter11, gate392inter12, gate99inter0, gate99inter1, gate99inter2, gate99inter3, gate99inter4, gate99inter5, gate99inter6, gate99inter7, gate99inter8, gate99inter9, gate99inter10, gate99inter11, gate99inter12, gate55inter0, gate55inter1, gate55inter2, gate55inter3, gate55inter4, gate55inter5, gate55inter6, gate55inter7, gate55inter8, gate55inter9, gate55inter10, gate55inter11, gate55inter12, gate125inter0, gate125inter1, gate125inter2, gate125inter3, gate125inter4, gate125inter5, gate125inter6, gate125inter7, gate125inter8, gate125inter9, gate125inter10, gate125inter11, gate125inter12, gate133inter0, gate133inter1, gate133inter2, gate133inter3, gate133inter4, gate133inter5, gate133inter6, gate133inter7, gate133inter8, gate133inter9, gate133inter10, gate133inter11, gate133inter12, gate121inter0, gate121inter1, gate121inter2, gate121inter3, gate121inter4, gate121inter5, gate121inter6, gate121inter7, gate121inter8, gate121inter9, gate121inter10, gate121inter11, gate121inter12, gate417inter0, gate417inter1, gate417inter2, gate417inter3, gate417inter4, gate417inter5, gate417inter6, gate417inter7, gate417inter8, gate417inter9, gate417inter10, gate417inter11, gate417inter12, gate448inter0, gate448inter1, gate448inter2, gate448inter3, gate448inter4, gate448inter5, gate448inter6, gate448inter7, gate448inter8, gate448inter9, gate448inter10, gate448inter11, gate448inter12, gate439inter0, gate439inter1, gate439inter2, gate439inter3, gate439inter4, gate439inter5, gate439inter6, gate439inter7, gate439inter8, gate439inter9, gate439inter10, gate439inter11, gate439inter12, gate61inter0, gate61inter1, gate61inter2, gate61inter3, gate61inter4, gate61inter5, gate61inter6, gate61inter7, gate61inter8, gate61inter9, gate61inter10, gate61inter11, gate61inter12, gate151inter0, gate151inter1, gate151inter2, gate151inter3, gate151inter4, gate151inter5, gate151inter6, gate151inter7, gate151inter8, gate151inter9, gate151inter10, gate151inter11, gate151inter12, gate22inter0, gate22inter1, gate22inter2, gate22inter3, gate22inter4, gate22inter5, gate22inter6, gate22inter7, gate22inter8, gate22inter9, gate22inter10, gate22inter11, gate22inter12, gate476inter0, gate476inter1, gate476inter2, gate476inter3, gate476inter4, gate476inter5, gate476inter6, gate476inter7, gate476inter8, gate476inter9, gate476inter10, gate476inter11, gate476inter12, gate19inter0, gate19inter1, gate19inter2, gate19inter3, gate19inter4, gate19inter5, gate19inter6, gate19inter7, gate19inter8, gate19inter9, gate19inter10, gate19inter11, gate19inter12, gate15inter0, gate15inter1, gate15inter2, gate15inter3, gate15inter4, gate15inter5, gate15inter6, gate15inter7, gate15inter8, gate15inter9, gate15inter10, gate15inter11, gate15inter12, gate388inter0, gate388inter1, gate388inter2, gate388inter3, gate388inter4, gate388inter5, gate388inter6, gate388inter7, gate388inter8, gate388inter9, gate388inter10, gate388inter11, gate388inter12, gate89inter0, gate89inter1, gate89inter2, gate89inter3, gate89inter4, gate89inter5, gate89inter6, gate89inter7, gate89inter8, gate89inter9, gate89inter10, gate89inter11, gate89inter12, gate134inter0, gate134inter1, gate134inter2, gate134inter3, gate134inter4, gate134inter5, gate134inter6, gate134inter7, gate134inter8, gate134inter9, gate134inter10, gate134inter11, gate134inter12, gate181inter0, gate181inter1, gate181inter2, gate181inter3, gate181inter4, gate181inter5, gate181inter6, gate181inter7, gate181inter8, gate181inter9, gate181inter10, gate181inter11, gate181inter12, gate225inter0, gate225inter1, gate225inter2, gate225inter3, gate225inter4, gate225inter5, gate225inter6, gate225inter7, gate225inter8, gate225inter9, gate225inter10, gate225inter11, gate225inter12, gate387inter0, gate387inter1, gate387inter2, gate387inter3, gate387inter4, gate387inter5, gate387inter6, gate387inter7, gate387inter8, gate387inter9, gate387inter10, gate387inter11, gate387inter12, gate162inter0, gate162inter1, gate162inter2, gate162inter3, gate162inter4, gate162inter5, gate162inter6, gate162inter7, gate162inter8, gate162inter9, gate162inter10, gate162inter11, gate162inter12, gate497inter0, gate497inter1, gate497inter2, gate497inter3, gate497inter4, gate497inter5, gate497inter6, gate497inter7, gate497inter8, gate497inter9, gate497inter10, gate497inter11, gate497inter12, gate487inter0, gate487inter1, gate487inter2, gate487inter3, gate487inter4, gate487inter5, gate487inter6, gate487inter7, gate487inter8, gate487inter9, gate487inter10, gate487inter11, gate487inter12, gate54inter0, gate54inter1, gate54inter2, gate54inter3, gate54inter4, gate54inter5, gate54inter6, gate54inter7, gate54inter8, gate54inter9, gate54inter10, gate54inter11, gate54inter12, gate221inter0, gate221inter1, gate221inter2, gate221inter3, gate221inter4, gate221inter5, gate221inter6, gate221inter7, gate221inter8, gate221inter9, gate221inter10, gate221inter11, gate221inter12, gate212inter0, gate212inter1, gate212inter2, gate212inter3, gate212inter4, gate212inter5, gate212inter6, gate212inter7, gate212inter8, gate212inter9, gate212inter10, gate212inter11, gate212inter12, gate466inter0, gate466inter1, gate466inter2, gate466inter3, gate466inter4, gate466inter5, gate466inter6, gate466inter7, gate466inter8, gate466inter9, gate466inter10, gate466inter11, gate466inter12, gate130inter0, gate130inter1, gate130inter2, gate130inter3, gate130inter4, gate130inter5, gate130inter6, gate130inter7, gate130inter8, gate130inter9, gate130inter10, gate130inter11, gate130inter12, gate409inter0, gate409inter1, gate409inter2, gate409inter3, gate409inter4, gate409inter5, gate409inter6, gate409inter7, gate409inter8, gate409inter9, gate409inter10, gate409inter11, gate409inter12, gate507inter0, gate507inter1, gate507inter2, gate507inter3, gate507inter4, gate507inter5, gate507inter6, gate507inter7, gate507inter8, gate507inter9, gate507inter10, gate507inter11, gate507inter12, gate283inter0, gate283inter1, gate283inter2, gate283inter3, gate283inter4, gate283inter5, gate283inter6, gate283inter7, gate283inter8, gate283inter9, gate283inter10, gate283inter11, gate283inter12, gate482inter0, gate482inter1, gate482inter2, gate482inter3, gate482inter4, gate482inter5, gate482inter6, gate482inter7, gate482inter8, gate482inter9, gate482inter10, gate482inter11, gate482inter12, gate411inter0, gate411inter1, gate411inter2, gate411inter3, gate411inter4, gate411inter5, gate411inter6, gate411inter7, gate411inter8, gate411inter9, gate411inter10, gate411inter11, gate411inter12, gate243inter0, gate243inter1, gate243inter2, gate243inter3, gate243inter4, gate243inter5, gate243inter6, gate243inter7, gate243inter8, gate243inter9, gate243inter10, gate243inter11, gate243inter12, gate119inter0, gate119inter1, gate119inter2, gate119inter3, gate119inter4, gate119inter5, gate119inter6, gate119inter7, gate119inter8, gate119inter9, gate119inter10, gate119inter11, gate119inter12, gate124inter0, gate124inter1, gate124inter2, gate124inter3, gate124inter4, gate124inter5, gate124inter6, gate124inter7, gate124inter8, gate124inter9, gate124inter10, gate124inter11, gate124inter12, gate143inter0, gate143inter1, gate143inter2, gate143inter3, gate143inter4, gate143inter5, gate143inter6, gate143inter7, gate143inter8, gate143inter9, gate143inter10, gate143inter11, gate143inter12, gate471inter0, gate471inter1, gate471inter2, gate471inter3, gate471inter4, gate471inter5, gate471inter6, gate471inter7, gate471inter8, gate471inter9, gate471inter10, gate471inter11, gate471inter12, gate194inter0, gate194inter1, gate194inter2, gate194inter3, gate194inter4, gate194inter5, gate194inter6, gate194inter7, gate194inter8, gate194inter9, gate194inter10, gate194inter11, gate194inter12, gate486inter0, gate486inter1, gate486inter2, gate486inter3, gate486inter4, gate486inter5, gate486inter6, gate486inter7, gate486inter8, gate486inter9, gate486inter10, gate486inter11, gate486inter12, gate48inter0, gate48inter1, gate48inter2, gate48inter3, gate48inter4, gate48inter5, gate48inter6, gate48inter7, gate48inter8, gate48inter9, gate48inter10, gate48inter11, gate48inter12, gate474inter0, gate474inter1, gate474inter2, gate474inter3, gate474inter4, gate474inter5, gate474inter6, gate474inter7, gate474inter8, gate474inter9, gate474inter10, gate474inter11, gate474inter12, gate461inter0, gate461inter1, gate461inter2, gate461inter3, gate461inter4, gate461inter5, gate461inter6, gate461inter7, gate461inter8, gate461inter9, gate461inter10, gate461inter11, gate461inter12, gate481inter0, gate481inter1, gate481inter2, gate481inter3, gate481inter4, gate481inter5, gate481inter6, gate481inter7, gate481inter8, gate481inter9, gate481inter10, gate481inter11, gate481inter12, gate288inter0, gate288inter1, gate288inter2, gate288inter3, gate288inter4, gate288inter5, gate288inter6, gate288inter7, gate288inter8, gate288inter9, gate288inter10, gate288inter11, gate288inter12, gate398inter0, gate398inter1, gate398inter2, gate398inter3, gate398inter4, gate398inter5, gate398inter6, gate398inter7, gate398inter8, gate398inter9, gate398inter10, gate398inter11, gate398inter12, gate294inter0, gate294inter1, gate294inter2, gate294inter3, gate294inter4, gate294inter5, gate294inter6, gate294inter7, gate294inter8, gate294inter9, gate294inter10, gate294inter11, gate294inter12, gate236inter0, gate236inter1, gate236inter2, gate236inter3, gate236inter4, gate236inter5, gate236inter6, gate236inter7, gate236inter8, gate236inter9, gate236inter10, gate236inter11, gate236inter12, gate97inter0, gate97inter1, gate97inter2, gate97inter3, gate97inter4, gate97inter5, gate97inter6, gate97inter7, gate97inter8, gate97inter9, gate97inter10, gate97inter11, gate97inter12, gate66inter0, gate66inter1, gate66inter2, gate66inter3, gate66inter4, gate66inter5, gate66inter6, gate66inter7, gate66inter8, gate66inter9, gate66inter10, gate66inter11, gate66inter12, gate72inter0, gate72inter1, gate72inter2, gate72inter3, gate72inter4, gate72inter5, gate72inter6, gate72inter7, gate72inter8, gate72inter9, gate72inter10, gate72inter11, gate72inter12, gate420inter0, gate420inter1, gate420inter2, gate420inter3, gate420inter4, gate420inter5, gate420inter6, gate420inter7, gate420inter8, gate420inter9, gate420inter10, gate420inter11, gate420inter12, gate271inter0, gate271inter1, gate271inter2, gate271inter3, gate271inter4, gate271inter5, gate271inter6, gate271inter7, gate271inter8, gate271inter9, gate271inter10, gate271inter11, gate271inter12, gate27inter0, gate27inter1, gate27inter2, gate27inter3, gate27inter4, gate27inter5, gate27inter6, gate27inter7, gate27inter8, gate27inter9, gate27inter10, gate27inter11, gate27inter12, gate241inter0, gate241inter1, gate241inter2, gate241inter3, gate241inter4, gate241inter5, gate241inter6, gate241inter7, gate241inter8, gate241inter9, gate241inter10, gate241inter11, gate241inter12, gate93inter0, gate93inter1, gate93inter2, gate93inter3, gate93inter4, gate93inter5, gate93inter6, gate93inter7, gate93inter8, gate93inter9, gate93inter10, gate93inter11, gate93inter12, gate454inter0, gate454inter1, gate454inter2, gate454inter3, gate454inter4, gate454inter5, gate454inter6, gate454inter7, gate454inter8, gate454inter9, gate454inter10, gate454inter11, gate454inter12, gate140inter0, gate140inter1, gate140inter2, gate140inter3, gate140inter4, gate140inter5, gate140inter6, gate140inter7, gate140inter8, gate140inter9, gate140inter10, gate140inter11, gate140inter12, gate502inter0, gate502inter1, gate502inter2, gate502inter3, gate502inter4, gate502inter5, gate502inter6, gate502inter7, gate502inter8, gate502inter9, gate502inter10, gate502inter11, gate502inter12, gate402inter0, gate402inter1, gate402inter2, gate402inter3, gate402inter4, gate402inter5, gate402inter6, gate402inter7, gate402inter8, gate402inter9, gate402inter10, gate402inter11, gate402inter12, gate235inter0, gate235inter1, gate235inter2, gate235inter3, gate235inter4, gate235inter5, gate235inter6, gate235inter7, gate235inter8, gate235inter9, gate235inter10, gate235inter11, gate235inter12, gate145inter0, gate145inter1, gate145inter2, gate145inter3, gate145inter4, gate145inter5, gate145inter6, gate145inter7, gate145inter8, gate145inter9, gate145inter10, gate145inter11, gate145inter12, gate449inter0, gate449inter1, gate449inter2, gate449inter3, gate449inter4, gate449inter5, gate449inter6, gate449inter7, gate449inter8, gate449inter9, gate449inter10, gate449inter11, gate449inter12, gate281inter0, gate281inter1, gate281inter2, gate281inter3, gate281inter4, gate281inter5, gate281inter6, gate281inter7, gate281inter8, gate281inter9, gate281inter10, gate281inter11, gate281inter12, gate76inter0, gate76inter1, gate76inter2, gate76inter3, gate76inter4, gate76inter5, gate76inter6, gate76inter7, gate76inter8, gate76inter9, gate76inter10, gate76inter11, gate76inter12, gate155inter0, gate155inter1, gate155inter2, gate155inter3, gate155inter4, gate155inter5, gate155inter6, gate155inter7, gate155inter8, gate155inter9, gate155inter10, gate155inter11, gate155inter12, gate137inter0, gate137inter1, gate137inter2, gate137inter3, gate137inter4, gate137inter5, gate137inter6, gate137inter7, gate137inter8, gate137inter9, gate137inter10, gate137inter11, gate137inter12, gate200inter0, gate200inter1, gate200inter2, gate200inter3, gate200inter4, gate200inter5, gate200inter6, gate200inter7, gate200inter8, gate200inter9, gate200inter10, gate200inter11, gate200inter12, gate158inter0, gate158inter1, gate158inter2, gate158inter3, gate158inter4, gate158inter5, gate158inter6, gate158inter7, gate158inter8, gate158inter9, gate158inter10, gate158inter11, gate158inter12, gate468inter0, gate468inter1, gate468inter2, gate468inter3, gate468inter4, gate468inter5, gate468inter6, gate468inter7, gate468inter8, gate468inter9, gate468inter10, gate468inter11, gate468inter12, gate219inter0, gate219inter1, gate219inter2, gate219inter3, gate219inter4, gate219inter5, gate219inter6, gate219inter7, gate219inter8, gate219inter9, gate219inter10, gate219inter11, gate219inter12, gate101inter0, gate101inter1, gate101inter2, gate101inter3, gate101inter4, gate101inter5, gate101inter6, gate101inter7, gate101inter8, gate101inter9, gate101inter10, gate101inter11, gate101inter12, gate456inter0, gate456inter1, gate456inter2, gate456inter3, gate456inter4, gate456inter5, gate456inter6, gate456inter7, gate456inter8, gate456inter9, gate456inter10, gate456inter11, gate456inter12, gate289inter0, gate289inter1, gate289inter2, gate289inter3, gate289inter4, gate289inter5, gate289inter6, gate289inter7, gate289inter8, gate289inter9, gate289inter10, gate289inter11, gate289inter12, gate211inter0, gate211inter1, gate211inter2, gate211inter3, gate211inter4, gate211inter5, gate211inter6, gate211inter7, gate211inter8, gate211inter9, gate211inter10, gate211inter11, gate211inter12, gate462inter0, gate462inter1, gate462inter2, gate462inter3, gate462inter4, gate462inter5, gate462inter6, gate462inter7, gate462inter8, gate462inter9, gate462inter10, gate462inter11, gate462inter12, gate205inter0, gate205inter1, gate205inter2, gate205inter3, gate205inter4, gate205inter5, gate205inter6, gate205inter7, gate205inter8, gate205inter9, gate205inter10, gate205inter11, gate205inter12, gate120inter0, gate120inter1, gate120inter2, gate120inter3, gate120inter4, gate120inter5, gate120inter6, gate120inter7, gate120inter8, gate120inter9, gate120inter10, gate120inter11, gate120inter12, gate16inter0, gate16inter1, gate16inter2, gate16inter3, gate16inter4, gate16inter5, gate16inter6, gate16inter7, gate16inter8, gate16inter9, gate16inter10, gate16inter11, gate16inter12, gate56inter0, gate56inter1, gate56inter2, gate56inter3, gate56inter4, gate56inter5, gate56inter6, gate56inter7, gate56inter8, gate56inter9, gate56inter10, gate56inter11, gate56inter12, gate282inter0, gate282inter1, gate282inter2, gate282inter3, gate282inter4, gate282inter5, gate282inter6, gate282inter7, gate282inter8, gate282inter9, gate282inter10, gate282inter11, gate282inter12, gate488inter0, gate488inter1, gate488inter2, gate488inter3, gate488inter4, gate488inter5, gate488inter6, gate488inter7, gate488inter8, gate488inter9, gate488inter10, gate488inter11, gate488inter12, gate514inter0, gate514inter1, gate514inter2, gate514inter3, gate514inter4, gate514inter5, gate514inter6, gate514inter7, gate514inter8, gate514inter9, gate514inter10, gate514inter11, gate514inter12, gate434inter0, gate434inter1, gate434inter2, gate434inter3, gate434inter4, gate434inter5, gate434inter6, gate434inter7, gate434inter8, gate434inter9, gate434inter10, gate434inter11, gate434inter12, gate156inter0, gate156inter1, gate156inter2, gate156inter3, gate156inter4, gate156inter5, gate156inter6, gate156inter7, gate156inter8, gate156inter9, gate156inter10, gate156inter11, gate156inter12, gate139inter0, gate139inter1, gate139inter2, gate139inter3, gate139inter4, gate139inter5, gate139inter6, gate139inter7, gate139inter8, gate139inter9, gate139inter10, gate139inter11, gate139inter12;



and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );
nand2 gate9( .a(G1), .b(G2), .O(G266) );

  xor2  gate939(.a(G4), .b(G3), .O(gate10inter0));
  nand2 gate940(.a(gate10inter0), .b(s_56), .O(gate10inter1));
  and2  gate941(.a(G4), .b(G3), .O(gate10inter2));
  inv1  gate942(.a(s_56), .O(gate10inter3));
  inv1  gate943(.a(s_57), .O(gate10inter4));
  nand2 gate944(.a(gate10inter4), .b(gate10inter3), .O(gate10inter5));
  nor2  gate945(.a(gate10inter5), .b(gate10inter2), .O(gate10inter6));
  inv1  gate946(.a(G3), .O(gate10inter7));
  inv1  gate947(.a(G4), .O(gate10inter8));
  nand2 gate948(.a(gate10inter8), .b(gate10inter7), .O(gate10inter9));
  nand2 gate949(.a(s_57), .b(gate10inter3), .O(gate10inter10));
  nor2  gate950(.a(gate10inter10), .b(gate10inter9), .O(gate10inter11));
  nor2  gate951(.a(gate10inter11), .b(gate10inter6), .O(gate10inter12));
  nand2 gate952(.a(gate10inter12), .b(gate10inter1), .O(G269));
nand2 gate11( .a(G5), .b(G6), .O(G272) );
nand2 gate12( .a(G7), .b(G8), .O(G275) );

  xor2  gate1191(.a(G10), .b(G9), .O(gate13inter0));
  nand2 gate1192(.a(gate13inter0), .b(s_92), .O(gate13inter1));
  and2  gate1193(.a(G10), .b(G9), .O(gate13inter2));
  inv1  gate1194(.a(s_92), .O(gate13inter3));
  inv1  gate1195(.a(s_93), .O(gate13inter4));
  nand2 gate1196(.a(gate13inter4), .b(gate13inter3), .O(gate13inter5));
  nor2  gate1197(.a(gate13inter5), .b(gate13inter2), .O(gate13inter6));
  inv1  gate1198(.a(G9), .O(gate13inter7));
  inv1  gate1199(.a(G10), .O(gate13inter8));
  nand2 gate1200(.a(gate13inter8), .b(gate13inter7), .O(gate13inter9));
  nand2 gate1201(.a(s_93), .b(gate13inter3), .O(gate13inter10));
  nor2  gate1202(.a(gate13inter10), .b(gate13inter9), .O(gate13inter11));
  nor2  gate1203(.a(gate13inter11), .b(gate13inter6), .O(gate13inter12));
  nand2 gate1204(.a(gate13inter12), .b(gate13inter1), .O(G278));

  xor2  gate1023(.a(G12), .b(G11), .O(gate14inter0));
  nand2 gate1024(.a(gate14inter0), .b(s_68), .O(gate14inter1));
  and2  gate1025(.a(G12), .b(G11), .O(gate14inter2));
  inv1  gate1026(.a(s_68), .O(gate14inter3));
  inv1  gate1027(.a(s_69), .O(gate14inter4));
  nand2 gate1028(.a(gate14inter4), .b(gate14inter3), .O(gate14inter5));
  nor2  gate1029(.a(gate14inter5), .b(gate14inter2), .O(gate14inter6));
  inv1  gate1030(.a(G11), .O(gate14inter7));
  inv1  gate1031(.a(G12), .O(gate14inter8));
  nand2 gate1032(.a(gate14inter8), .b(gate14inter7), .O(gate14inter9));
  nand2 gate1033(.a(s_69), .b(gate14inter3), .O(gate14inter10));
  nor2  gate1034(.a(gate14inter10), .b(gate14inter9), .O(gate14inter11));
  nor2  gate1035(.a(gate14inter11), .b(gate14inter6), .O(gate14inter12));
  nand2 gate1036(.a(gate14inter12), .b(gate14inter1), .O(G281));

  xor2  gate1569(.a(G14), .b(G13), .O(gate15inter0));
  nand2 gate1570(.a(gate15inter0), .b(s_146), .O(gate15inter1));
  and2  gate1571(.a(G14), .b(G13), .O(gate15inter2));
  inv1  gate1572(.a(s_146), .O(gate15inter3));
  inv1  gate1573(.a(s_147), .O(gate15inter4));
  nand2 gate1574(.a(gate15inter4), .b(gate15inter3), .O(gate15inter5));
  nor2  gate1575(.a(gate15inter5), .b(gate15inter2), .O(gate15inter6));
  inv1  gate1576(.a(G13), .O(gate15inter7));
  inv1  gate1577(.a(G14), .O(gate15inter8));
  nand2 gate1578(.a(gate15inter8), .b(gate15inter7), .O(gate15inter9));
  nand2 gate1579(.a(s_147), .b(gate15inter3), .O(gate15inter10));
  nor2  gate1580(.a(gate15inter10), .b(gate15inter9), .O(gate15inter11));
  nor2  gate1581(.a(gate15inter11), .b(gate15inter6), .O(gate15inter12));
  nand2 gate1582(.a(gate15inter12), .b(gate15inter1), .O(G284));

  xor2  gate2479(.a(G16), .b(G15), .O(gate16inter0));
  nand2 gate2480(.a(gate16inter0), .b(s_276), .O(gate16inter1));
  and2  gate2481(.a(G16), .b(G15), .O(gate16inter2));
  inv1  gate2482(.a(s_276), .O(gate16inter3));
  inv1  gate2483(.a(s_277), .O(gate16inter4));
  nand2 gate2484(.a(gate16inter4), .b(gate16inter3), .O(gate16inter5));
  nor2  gate2485(.a(gate16inter5), .b(gate16inter2), .O(gate16inter6));
  inv1  gate2486(.a(G15), .O(gate16inter7));
  inv1  gate2487(.a(G16), .O(gate16inter8));
  nand2 gate2488(.a(gate16inter8), .b(gate16inter7), .O(gate16inter9));
  nand2 gate2489(.a(s_277), .b(gate16inter3), .O(gate16inter10));
  nor2  gate2490(.a(gate16inter10), .b(gate16inter9), .O(gate16inter11));
  nor2  gate2491(.a(gate16inter11), .b(gate16inter6), .O(gate16inter12));
  nand2 gate2492(.a(gate16inter12), .b(gate16inter1), .O(G287));
nand2 gate17( .a(G17), .b(G18), .O(G290) );
nand2 gate18( .a(G19), .b(G20), .O(G293) );

  xor2  gate1555(.a(G22), .b(G21), .O(gate19inter0));
  nand2 gate1556(.a(gate19inter0), .b(s_144), .O(gate19inter1));
  and2  gate1557(.a(G22), .b(G21), .O(gate19inter2));
  inv1  gate1558(.a(s_144), .O(gate19inter3));
  inv1  gate1559(.a(s_145), .O(gate19inter4));
  nand2 gate1560(.a(gate19inter4), .b(gate19inter3), .O(gate19inter5));
  nor2  gate1561(.a(gate19inter5), .b(gate19inter2), .O(gate19inter6));
  inv1  gate1562(.a(G21), .O(gate19inter7));
  inv1  gate1563(.a(G22), .O(gate19inter8));
  nand2 gate1564(.a(gate19inter8), .b(gate19inter7), .O(gate19inter9));
  nand2 gate1565(.a(s_145), .b(gate19inter3), .O(gate19inter10));
  nor2  gate1566(.a(gate19inter10), .b(gate19inter9), .O(gate19inter11));
  nor2  gate1567(.a(gate19inter11), .b(gate19inter6), .O(gate19inter12));
  nand2 gate1568(.a(gate19inter12), .b(gate19inter1), .O(G296));
nand2 gate20( .a(G23), .b(G24), .O(G299) );
nand2 gate21( .a(G25), .b(G26), .O(G302) );

  xor2  gate1527(.a(G28), .b(G27), .O(gate22inter0));
  nand2 gate1528(.a(gate22inter0), .b(s_140), .O(gate22inter1));
  and2  gate1529(.a(G28), .b(G27), .O(gate22inter2));
  inv1  gate1530(.a(s_140), .O(gate22inter3));
  inv1  gate1531(.a(s_141), .O(gate22inter4));
  nand2 gate1532(.a(gate22inter4), .b(gate22inter3), .O(gate22inter5));
  nor2  gate1533(.a(gate22inter5), .b(gate22inter2), .O(gate22inter6));
  inv1  gate1534(.a(G27), .O(gate22inter7));
  inv1  gate1535(.a(G28), .O(gate22inter8));
  nand2 gate1536(.a(gate22inter8), .b(gate22inter7), .O(gate22inter9));
  nand2 gate1537(.a(s_141), .b(gate22inter3), .O(gate22inter10));
  nor2  gate1538(.a(gate22inter10), .b(gate22inter9), .O(gate22inter11));
  nor2  gate1539(.a(gate22inter11), .b(gate22inter6), .O(gate22inter12));
  nand2 gate1540(.a(gate22inter12), .b(gate22inter1), .O(G305));
nand2 gate23( .a(G29), .b(G30), .O(G308) );
nand2 gate24( .a(G31), .b(G32), .O(G311) );
nand2 gate25( .a(G1), .b(G5), .O(G314) );
nand2 gate26( .a(G9), .b(G13), .O(G317) );

  xor2  gate2129(.a(G6), .b(G2), .O(gate27inter0));
  nand2 gate2130(.a(gate27inter0), .b(s_226), .O(gate27inter1));
  and2  gate2131(.a(G6), .b(G2), .O(gate27inter2));
  inv1  gate2132(.a(s_226), .O(gate27inter3));
  inv1  gate2133(.a(s_227), .O(gate27inter4));
  nand2 gate2134(.a(gate27inter4), .b(gate27inter3), .O(gate27inter5));
  nor2  gate2135(.a(gate27inter5), .b(gate27inter2), .O(gate27inter6));
  inv1  gate2136(.a(G2), .O(gate27inter7));
  inv1  gate2137(.a(G6), .O(gate27inter8));
  nand2 gate2138(.a(gate27inter8), .b(gate27inter7), .O(gate27inter9));
  nand2 gate2139(.a(s_227), .b(gate27inter3), .O(gate27inter10));
  nor2  gate2140(.a(gate27inter10), .b(gate27inter9), .O(gate27inter11));
  nor2  gate2141(.a(gate27inter11), .b(gate27inter6), .O(gate27inter12));
  nand2 gate2142(.a(gate27inter12), .b(gate27inter1), .O(G320));
nand2 gate28( .a(G10), .b(G14), .O(G323) );
nand2 gate29( .a(G3), .b(G7), .O(G326) );
nand2 gate30( .a(G11), .b(G15), .O(G329) );

  xor2  gate1163(.a(G8), .b(G4), .O(gate31inter0));
  nand2 gate1164(.a(gate31inter0), .b(s_88), .O(gate31inter1));
  and2  gate1165(.a(G8), .b(G4), .O(gate31inter2));
  inv1  gate1166(.a(s_88), .O(gate31inter3));
  inv1  gate1167(.a(s_89), .O(gate31inter4));
  nand2 gate1168(.a(gate31inter4), .b(gate31inter3), .O(gate31inter5));
  nor2  gate1169(.a(gate31inter5), .b(gate31inter2), .O(gate31inter6));
  inv1  gate1170(.a(G4), .O(gate31inter7));
  inv1  gate1171(.a(G8), .O(gate31inter8));
  nand2 gate1172(.a(gate31inter8), .b(gate31inter7), .O(gate31inter9));
  nand2 gate1173(.a(s_89), .b(gate31inter3), .O(gate31inter10));
  nor2  gate1174(.a(gate31inter10), .b(gate31inter9), .O(gate31inter11));
  nor2  gate1175(.a(gate31inter11), .b(gate31inter6), .O(gate31inter12));
  nand2 gate1176(.a(gate31inter12), .b(gate31inter1), .O(G332));
nand2 gate32( .a(G12), .b(G16), .O(G335) );
nand2 gate33( .a(G17), .b(G21), .O(G338) );
nand2 gate34( .a(G25), .b(G29), .O(G341) );
nand2 gate35( .a(G18), .b(G22), .O(G344) );
nand2 gate36( .a(G26), .b(G30), .O(G347) );
nand2 gate37( .a(G19), .b(G23), .O(G350) );

  xor2  gate1219(.a(G31), .b(G27), .O(gate38inter0));
  nand2 gate1220(.a(gate38inter0), .b(s_96), .O(gate38inter1));
  and2  gate1221(.a(G31), .b(G27), .O(gate38inter2));
  inv1  gate1222(.a(s_96), .O(gate38inter3));
  inv1  gate1223(.a(s_97), .O(gate38inter4));
  nand2 gate1224(.a(gate38inter4), .b(gate38inter3), .O(gate38inter5));
  nor2  gate1225(.a(gate38inter5), .b(gate38inter2), .O(gate38inter6));
  inv1  gate1226(.a(G27), .O(gate38inter7));
  inv1  gate1227(.a(G31), .O(gate38inter8));
  nand2 gate1228(.a(gate38inter8), .b(gate38inter7), .O(gate38inter9));
  nand2 gate1229(.a(s_97), .b(gate38inter3), .O(gate38inter10));
  nor2  gate1230(.a(gate38inter10), .b(gate38inter9), .O(gate38inter11));
  nor2  gate1231(.a(gate38inter11), .b(gate38inter6), .O(gate38inter12));
  nand2 gate1232(.a(gate38inter12), .b(gate38inter1), .O(G353));
nand2 gate39( .a(G20), .b(G24), .O(G356) );
nand2 gate40( .a(G28), .b(G32), .O(G359) );

  xor2  gate1233(.a(G266), .b(G1), .O(gate41inter0));
  nand2 gate1234(.a(gate41inter0), .b(s_98), .O(gate41inter1));
  and2  gate1235(.a(G266), .b(G1), .O(gate41inter2));
  inv1  gate1236(.a(s_98), .O(gate41inter3));
  inv1  gate1237(.a(s_99), .O(gate41inter4));
  nand2 gate1238(.a(gate41inter4), .b(gate41inter3), .O(gate41inter5));
  nor2  gate1239(.a(gate41inter5), .b(gate41inter2), .O(gate41inter6));
  inv1  gate1240(.a(G1), .O(gate41inter7));
  inv1  gate1241(.a(G266), .O(gate41inter8));
  nand2 gate1242(.a(gate41inter8), .b(gate41inter7), .O(gate41inter9));
  nand2 gate1243(.a(s_99), .b(gate41inter3), .O(gate41inter10));
  nor2  gate1244(.a(gate41inter10), .b(gate41inter9), .O(gate41inter11));
  nor2  gate1245(.a(gate41inter11), .b(gate41inter6), .O(gate41inter12));
  nand2 gate1246(.a(gate41inter12), .b(gate41inter1), .O(G362));
nand2 gate42( .a(G2), .b(G266), .O(G363) );

  xor2  gate1079(.a(G269), .b(G3), .O(gate43inter0));
  nand2 gate1080(.a(gate43inter0), .b(s_76), .O(gate43inter1));
  and2  gate1081(.a(G269), .b(G3), .O(gate43inter2));
  inv1  gate1082(.a(s_76), .O(gate43inter3));
  inv1  gate1083(.a(s_77), .O(gate43inter4));
  nand2 gate1084(.a(gate43inter4), .b(gate43inter3), .O(gate43inter5));
  nor2  gate1085(.a(gate43inter5), .b(gate43inter2), .O(gate43inter6));
  inv1  gate1086(.a(G3), .O(gate43inter7));
  inv1  gate1087(.a(G269), .O(gate43inter8));
  nand2 gate1088(.a(gate43inter8), .b(gate43inter7), .O(gate43inter9));
  nand2 gate1089(.a(s_77), .b(gate43inter3), .O(gate43inter10));
  nor2  gate1090(.a(gate43inter10), .b(gate43inter9), .O(gate43inter11));
  nor2  gate1091(.a(gate43inter11), .b(gate43inter6), .O(gate43inter12));
  nand2 gate1092(.a(gate43inter12), .b(gate43inter1), .O(G364));
nand2 gate44( .a(G4), .b(G269), .O(G365) );
nand2 gate45( .a(G5), .b(G272), .O(G366) );
nand2 gate46( .a(G6), .b(G272), .O(G367) );
nand2 gate47( .a(G7), .b(G275), .O(G368) );

  xor2  gate1947(.a(G275), .b(G8), .O(gate48inter0));
  nand2 gate1948(.a(gate48inter0), .b(s_200), .O(gate48inter1));
  and2  gate1949(.a(G275), .b(G8), .O(gate48inter2));
  inv1  gate1950(.a(s_200), .O(gate48inter3));
  inv1  gate1951(.a(s_201), .O(gate48inter4));
  nand2 gate1952(.a(gate48inter4), .b(gate48inter3), .O(gate48inter5));
  nor2  gate1953(.a(gate48inter5), .b(gate48inter2), .O(gate48inter6));
  inv1  gate1954(.a(G8), .O(gate48inter7));
  inv1  gate1955(.a(G275), .O(gate48inter8));
  nand2 gate1956(.a(gate48inter8), .b(gate48inter7), .O(gate48inter9));
  nand2 gate1957(.a(s_201), .b(gate48inter3), .O(gate48inter10));
  nor2  gate1958(.a(gate48inter10), .b(gate48inter9), .O(gate48inter11));
  nor2  gate1959(.a(gate48inter11), .b(gate48inter6), .O(gate48inter12));
  nand2 gate1960(.a(gate48inter12), .b(gate48inter1), .O(G369));
nand2 gate49( .a(G9), .b(G278), .O(G370) );
nand2 gate50( .a(G10), .b(G278), .O(G371) );
nand2 gate51( .a(G11), .b(G281), .O(G372) );
nand2 gate52( .a(G12), .b(G281), .O(G373) );

  xor2  gate925(.a(G284), .b(G13), .O(gate53inter0));
  nand2 gate926(.a(gate53inter0), .b(s_54), .O(gate53inter1));
  and2  gate927(.a(G284), .b(G13), .O(gate53inter2));
  inv1  gate928(.a(s_54), .O(gate53inter3));
  inv1  gate929(.a(s_55), .O(gate53inter4));
  nand2 gate930(.a(gate53inter4), .b(gate53inter3), .O(gate53inter5));
  nor2  gate931(.a(gate53inter5), .b(gate53inter2), .O(gate53inter6));
  inv1  gate932(.a(G13), .O(gate53inter7));
  inv1  gate933(.a(G284), .O(gate53inter8));
  nand2 gate934(.a(gate53inter8), .b(gate53inter7), .O(gate53inter9));
  nand2 gate935(.a(s_55), .b(gate53inter3), .O(gate53inter10));
  nor2  gate936(.a(gate53inter10), .b(gate53inter9), .O(gate53inter11));
  nor2  gate937(.a(gate53inter11), .b(gate53inter6), .O(gate53inter12));
  nand2 gate938(.a(gate53inter12), .b(gate53inter1), .O(G374));

  xor2  gate1709(.a(G284), .b(G14), .O(gate54inter0));
  nand2 gate1710(.a(gate54inter0), .b(s_166), .O(gate54inter1));
  and2  gate1711(.a(G284), .b(G14), .O(gate54inter2));
  inv1  gate1712(.a(s_166), .O(gate54inter3));
  inv1  gate1713(.a(s_167), .O(gate54inter4));
  nand2 gate1714(.a(gate54inter4), .b(gate54inter3), .O(gate54inter5));
  nor2  gate1715(.a(gate54inter5), .b(gate54inter2), .O(gate54inter6));
  inv1  gate1716(.a(G14), .O(gate54inter7));
  inv1  gate1717(.a(G284), .O(gate54inter8));
  nand2 gate1718(.a(gate54inter8), .b(gate54inter7), .O(gate54inter9));
  nand2 gate1719(.a(s_167), .b(gate54inter3), .O(gate54inter10));
  nor2  gate1720(.a(gate54inter10), .b(gate54inter9), .O(gate54inter11));
  nor2  gate1721(.a(gate54inter11), .b(gate54inter6), .O(gate54inter12));
  nand2 gate1722(.a(gate54inter12), .b(gate54inter1), .O(G375));

  xor2  gate1401(.a(G287), .b(G15), .O(gate55inter0));
  nand2 gate1402(.a(gate55inter0), .b(s_122), .O(gate55inter1));
  and2  gate1403(.a(G287), .b(G15), .O(gate55inter2));
  inv1  gate1404(.a(s_122), .O(gate55inter3));
  inv1  gate1405(.a(s_123), .O(gate55inter4));
  nand2 gate1406(.a(gate55inter4), .b(gate55inter3), .O(gate55inter5));
  nor2  gate1407(.a(gate55inter5), .b(gate55inter2), .O(gate55inter6));
  inv1  gate1408(.a(G15), .O(gate55inter7));
  inv1  gate1409(.a(G287), .O(gate55inter8));
  nand2 gate1410(.a(gate55inter8), .b(gate55inter7), .O(gate55inter9));
  nand2 gate1411(.a(s_123), .b(gate55inter3), .O(gate55inter10));
  nor2  gate1412(.a(gate55inter10), .b(gate55inter9), .O(gate55inter11));
  nor2  gate1413(.a(gate55inter11), .b(gate55inter6), .O(gate55inter12));
  nand2 gate1414(.a(gate55inter12), .b(gate55inter1), .O(G376));

  xor2  gate2493(.a(G287), .b(G16), .O(gate56inter0));
  nand2 gate2494(.a(gate56inter0), .b(s_278), .O(gate56inter1));
  and2  gate2495(.a(G287), .b(G16), .O(gate56inter2));
  inv1  gate2496(.a(s_278), .O(gate56inter3));
  inv1  gate2497(.a(s_279), .O(gate56inter4));
  nand2 gate2498(.a(gate56inter4), .b(gate56inter3), .O(gate56inter5));
  nor2  gate2499(.a(gate56inter5), .b(gate56inter2), .O(gate56inter6));
  inv1  gate2500(.a(G16), .O(gate56inter7));
  inv1  gate2501(.a(G287), .O(gate56inter8));
  nand2 gate2502(.a(gate56inter8), .b(gate56inter7), .O(gate56inter9));
  nand2 gate2503(.a(s_279), .b(gate56inter3), .O(gate56inter10));
  nor2  gate2504(.a(gate56inter10), .b(gate56inter9), .O(gate56inter11));
  nor2  gate2505(.a(gate56inter11), .b(gate56inter6), .O(gate56inter12));
  nand2 gate2506(.a(gate56inter12), .b(gate56inter1), .O(G377));
nand2 gate57( .a(G17), .b(G290), .O(G378) );
nand2 gate58( .a(G18), .b(G290), .O(G379) );
nand2 gate59( .a(G19), .b(G293), .O(G380) );

  xor2  gate1051(.a(G293), .b(G20), .O(gate60inter0));
  nand2 gate1052(.a(gate60inter0), .b(s_72), .O(gate60inter1));
  and2  gate1053(.a(G293), .b(G20), .O(gate60inter2));
  inv1  gate1054(.a(s_72), .O(gate60inter3));
  inv1  gate1055(.a(s_73), .O(gate60inter4));
  nand2 gate1056(.a(gate60inter4), .b(gate60inter3), .O(gate60inter5));
  nor2  gate1057(.a(gate60inter5), .b(gate60inter2), .O(gate60inter6));
  inv1  gate1058(.a(G20), .O(gate60inter7));
  inv1  gate1059(.a(G293), .O(gate60inter8));
  nand2 gate1060(.a(gate60inter8), .b(gate60inter7), .O(gate60inter9));
  nand2 gate1061(.a(s_73), .b(gate60inter3), .O(gate60inter10));
  nor2  gate1062(.a(gate60inter10), .b(gate60inter9), .O(gate60inter11));
  nor2  gate1063(.a(gate60inter11), .b(gate60inter6), .O(gate60inter12));
  nand2 gate1064(.a(gate60inter12), .b(gate60inter1), .O(G381));

  xor2  gate1499(.a(G296), .b(G21), .O(gate61inter0));
  nand2 gate1500(.a(gate61inter0), .b(s_136), .O(gate61inter1));
  and2  gate1501(.a(G296), .b(G21), .O(gate61inter2));
  inv1  gate1502(.a(s_136), .O(gate61inter3));
  inv1  gate1503(.a(s_137), .O(gate61inter4));
  nand2 gate1504(.a(gate61inter4), .b(gate61inter3), .O(gate61inter5));
  nor2  gate1505(.a(gate61inter5), .b(gate61inter2), .O(gate61inter6));
  inv1  gate1506(.a(G21), .O(gate61inter7));
  inv1  gate1507(.a(G296), .O(gate61inter8));
  nand2 gate1508(.a(gate61inter8), .b(gate61inter7), .O(gate61inter9));
  nand2 gate1509(.a(s_137), .b(gate61inter3), .O(gate61inter10));
  nor2  gate1510(.a(gate61inter10), .b(gate61inter9), .O(gate61inter11));
  nor2  gate1511(.a(gate61inter11), .b(gate61inter6), .O(gate61inter12));
  nand2 gate1512(.a(gate61inter12), .b(gate61inter1), .O(G382));
nand2 gate62( .a(G22), .b(G296), .O(G383) );
nand2 gate63( .a(G23), .b(G299), .O(G384) );
nand2 gate64( .a(G24), .b(G299), .O(G385) );
nand2 gate65( .a(G25), .b(G302), .O(G386) );

  xor2  gate2073(.a(G302), .b(G26), .O(gate66inter0));
  nand2 gate2074(.a(gate66inter0), .b(s_218), .O(gate66inter1));
  and2  gate2075(.a(G302), .b(G26), .O(gate66inter2));
  inv1  gate2076(.a(s_218), .O(gate66inter3));
  inv1  gate2077(.a(s_219), .O(gate66inter4));
  nand2 gate2078(.a(gate66inter4), .b(gate66inter3), .O(gate66inter5));
  nor2  gate2079(.a(gate66inter5), .b(gate66inter2), .O(gate66inter6));
  inv1  gate2080(.a(G26), .O(gate66inter7));
  inv1  gate2081(.a(G302), .O(gate66inter8));
  nand2 gate2082(.a(gate66inter8), .b(gate66inter7), .O(gate66inter9));
  nand2 gate2083(.a(s_219), .b(gate66inter3), .O(gate66inter10));
  nor2  gate2084(.a(gate66inter10), .b(gate66inter9), .O(gate66inter11));
  nor2  gate2085(.a(gate66inter11), .b(gate66inter6), .O(gate66inter12));
  nand2 gate2086(.a(gate66inter12), .b(gate66inter1), .O(G387));

  xor2  gate953(.a(G305), .b(G27), .O(gate67inter0));
  nand2 gate954(.a(gate67inter0), .b(s_58), .O(gate67inter1));
  and2  gate955(.a(G305), .b(G27), .O(gate67inter2));
  inv1  gate956(.a(s_58), .O(gate67inter3));
  inv1  gate957(.a(s_59), .O(gate67inter4));
  nand2 gate958(.a(gate67inter4), .b(gate67inter3), .O(gate67inter5));
  nor2  gate959(.a(gate67inter5), .b(gate67inter2), .O(gate67inter6));
  inv1  gate960(.a(G27), .O(gate67inter7));
  inv1  gate961(.a(G305), .O(gate67inter8));
  nand2 gate962(.a(gate67inter8), .b(gate67inter7), .O(gate67inter9));
  nand2 gate963(.a(s_59), .b(gate67inter3), .O(gate67inter10));
  nor2  gate964(.a(gate67inter10), .b(gate67inter9), .O(gate67inter11));
  nor2  gate965(.a(gate67inter11), .b(gate67inter6), .O(gate67inter12));
  nand2 gate966(.a(gate67inter12), .b(gate67inter1), .O(G388));
nand2 gate68( .a(G28), .b(G305), .O(G389) );
nand2 gate69( .a(G29), .b(G308), .O(G390) );

  xor2  gate631(.a(G308), .b(G30), .O(gate70inter0));
  nand2 gate632(.a(gate70inter0), .b(s_12), .O(gate70inter1));
  and2  gate633(.a(G308), .b(G30), .O(gate70inter2));
  inv1  gate634(.a(s_12), .O(gate70inter3));
  inv1  gate635(.a(s_13), .O(gate70inter4));
  nand2 gate636(.a(gate70inter4), .b(gate70inter3), .O(gate70inter5));
  nor2  gate637(.a(gate70inter5), .b(gate70inter2), .O(gate70inter6));
  inv1  gate638(.a(G30), .O(gate70inter7));
  inv1  gate639(.a(G308), .O(gate70inter8));
  nand2 gate640(.a(gate70inter8), .b(gate70inter7), .O(gate70inter9));
  nand2 gate641(.a(s_13), .b(gate70inter3), .O(gate70inter10));
  nor2  gate642(.a(gate70inter10), .b(gate70inter9), .O(gate70inter11));
  nor2  gate643(.a(gate70inter11), .b(gate70inter6), .O(gate70inter12));
  nand2 gate644(.a(gate70inter12), .b(gate70inter1), .O(G391));
nand2 gate71( .a(G31), .b(G311), .O(G392) );

  xor2  gate2087(.a(G311), .b(G32), .O(gate72inter0));
  nand2 gate2088(.a(gate72inter0), .b(s_220), .O(gate72inter1));
  and2  gate2089(.a(G311), .b(G32), .O(gate72inter2));
  inv1  gate2090(.a(s_220), .O(gate72inter3));
  inv1  gate2091(.a(s_221), .O(gate72inter4));
  nand2 gate2092(.a(gate72inter4), .b(gate72inter3), .O(gate72inter5));
  nor2  gate2093(.a(gate72inter5), .b(gate72inter2), .O(gate72inter6));
  inv1  gate2094(.a(G32), .O(gate72inter7));
  inv1  gate2095(.a(G311), .O(gate72inter8));
  nand2 gate2096(.a(gate72inter8), .b(gate72inter7), .O(gate72inter9));
  nand2 gate2097(.a(s_221), .b(gate72inter3), .O(gate72inter10));
  nor2  gate2098(.a(gate72inter10), .b(gate72inter9), .O(gate72inter11));
  nor2  gate2099(.a(gate72inter11), .b(gate72inter6), .O(gate72inter12));
  nand2 gate2100(.a(gate72inter12), .b(gate72inter1), .O(G393));
nand2 gate73( .a(G1), .b(G314), .O(G394) );
nand2 gate74( .a(G5), .b(G314), .O(G395) );
nand2 gate75( .a(G9), .b(G317), .O(G396) );

  xor2  gate2283(.a(G317), .b(G13), .O(gate76inter0));
  nand2 gate2284(.a(gate76inter0), .b(s_248), .O(gate76inter1));
  and2  gate2285(.a(G317), .b(G13), .O(gate76inter2));
  inv1  gate2286(.a(s_248), .O(gate76inter3));
  inv1  gate2287(.a(s_249), .O(gate76inter4));
  nand2 gate2288(.a(gate76inter4), .b(gate76inter3), .O(gate76inter5));
  nor2  gate2289(.a(gate76inter5), .b(gate76inter2), .O(gate76inter6));
  inv1  gate2290(.a(G13), .O(gate76inter7));
  inv1  gate2291(.a(G317), .O(gate76inter8));
  nand2 gate2292(.a(gate76inter8), .b(gate76inter7), .O(gate76inter9));
  nand2 gate2293(.a(s_249), .b(gate76inter3), .O(gate76inter10));
  nor2  gate2294(.a(gate76inter10), .b(gate76inter9), .O(gate76inter11));
  nor2  gate2295(.a(gate76inter11), .b(gate76inter6), .O(gate76inter12));
  nand2 gate2296(.a(gate76inter12), .b(gate76inter1), .O(G397));
nand2 gate77( .a(G2), .b(G320), .O(G398) );
nand2 gate78( .a(G6), .b(G320), .O(G399) );
nand2 gate79( .a(G10), .b(G323), .O(G400) );
nand2 gate80( .a(G14), .b(G323), .O(G401) );
nand2 gate81( .a(G3), .b(G326), .O(G402) );
nand2 gate82( .a(G7), .b(G326), .O(G403) );
nand2 gate83( .a(G11), .b(G329), .O(G404) );

  xor2  gate561(.a(G329), .b(G15), .O(gate84inter0));
  nand2 gate562(.a(gate84inter0), .b(s_2), .O(gate84inter1));
  and2  gate563(.a(G329), .b(G15), .O(gate84inter2));
  inv1  gate564(.a(s_2), .O(gate84inter3));
  inv1  gate565(.a(s_3), .O(gate84inter4));
  nand2 gate566(.a(gate84inter4), .b(gate84inter3), .O(gate84inter5));
  nor2  gate567(.a(gate84inter5), .b(gate84inter2), .O(gate84inter6));
  inv1  gate568(.a(G15), .O(gate84inter7));
  inv1  gate569(.a(G329), .O(gate84inter8));
  nand2 gate570(.a(gate84inter8), .b(gate84inter7), .O(gate84inter9));
  nand2 gate571(.a(s_3), .b(gate84inter3), .O(gate84inter10));
  nor2  gate572(.a(gate84inter10), .b(gate84inter9), .O(gate84inter11));
  nor2  gate573(.a(gate84inter11), .b(gate84inter6), .O(gate84inter12));
  nand2 gate574(.a(gate84inter12), .b(gate84inter1), .O(G405));
nand2 gate85( .a(G4), .b(G332), .O(G406) );
nand2 gate86( .a(G8), .b(G332), .O(G407) );
nand2 gate87( .a(G12), .b(G335), .O(G408) );
nand2 gate88( .a(G16), .b(G335), .O(G409) );

  xor2  gate1597(.a(G338), .b(G17), .O(gate89inter0));
  nand2 gate1598(.a(gate89inter0), .b(s_150), .O(gate89inter1));
  and2  gate1599(.a(G338), .b(G17), .O(gate89inter2));
  inv1  gate1600(.a(s_150), .O(gate89inter3));
  inv1  gate1601(.a(s_151), .O(gate89inter4));
  nand2 gate1602(.a(gate89inter4), .b(gate89inter3), .O(gate89inter5));
  nor2  gate1603(.a(gate89inter5), .b(gate89inter2), .O(gate89inter6));
  inv1  gate1604(.a(G17), .O(gate89inter7));
  inv1  gate1605(.a(G338), .O(gate89inter8));
  nand2 gate1606(.a(gate89inter8), .b(gate89inter7), .O(gate89inter9));
  nand2 gate1607(.a(s_151), .b(gate89inter3), .O(gate89inter10));
  nor2  gate1608(.a(gate89inter10), .b(gate89inter9), .O(gate89inter11));
  nor2  gate1609(.a(gate89inter11), .b(gate89inter6), .O(gate89inter12));
  nand2 gate1610(.a(gate89inter12), .b(gate89inter1), .O(G410));
nand2 gate90( .a(G21), .b(G338), .O(G411) );
nand2 gate91( .a(G25), .b(G341), .O(G412) );
nand2 gate92( .a(G29), .b(G341), .O(G413) );

  xor2  gate2157(.a(G344), .b(G18), .O(gate93inter0));
  nand2 gate2158(.a(gate93inter0), .b(s_230), .O(gate93inter1));
  and2  gate2159(.a(G344), .b(G18), .O(gate93inter2));
  inv1  gate2160(.a(s_230), .O(gate93inter3));
  inv1  gate2161(.a(s_231), .O(gate93inter4));
  nand2 gate2162(.a(gate93inter4), .b(gate93inter3), .O(gate93inter5));
  nor2  gate2163(.a(gate93inter5), .b(gate93inter2), .O(gate93inter6));
  inv1  gate2164(.a(G18), .O(gate93inter7));
  inv1  gate2165(.a(G344), .O(gate93inter8));
  nand2 gate2166(.a(gate93inter8), .b(gate93inter7), .O(gate93inter9));
  nand2 gate2167(.a(s_231), .b(gate93inter3), .O(gate93inter10));
  nor2  gate2168(.a(gate93inter10), .b(gate93inter9), .O(gate93inter11));
  nor2  gate2169(.a(gate93inter11), .b(gate93inter6), .O(gate93inter12));
  nand2 gate2170(.a(gate93inter12), .b(gate93inter1), .O(G414));

  xor2  gate1107(.a(G344), .b(G22), .O(gate94inter0));
  nand2 gate1108(.a(gate94inter0), .b(s_80), .O(gate94inter1));
  and2  gate1109(.a(G344), .b(G22), .O(gate94inter2));
  inv1  gate1110(.a(s_80), .O(gate94inter3));
  inv1  gate1111(.a(s_81), .O(gate94inter4));
  nand2 gate1112(.a(gate94inter4), .b(gate94inter3), .O(gate94inter5));
  nor2  gate1113(.a(gate94inter5), .b(gate94inter2), .O(gate94inter6));
  inv1  gate1114(.a(G22), .O(gate94inter7));
  inv1  gate1115(.a(G344), .O(gate94inter8));
  nand2 gate1116(.a(gate94inter8), .b(gate94inter7), .O(gate94inter9));
  nand2 gate1117(.a(s_81), .b(gate94inter3), .O(gate94inter10));
  nor2  gate1118(.a(gate94inter10), .b(gate94inter9), .O(gate94inter11));
  nor2  gate1119(.a(gate94inter11), .b(gate94inter6), .O(gate94inter12));
  nand2 gate1120(.a(gate94inter12), .b(gate94inter1), .O(G415));
nand2 gate95( .a(G26), .b(G347), .O(G416) );
nand2 gate96( .a(G30), .b(G347), .O(G417) );

  xor2  gate2059(.a(G350), .b(G19), .O(gate97inter0));
  nand2 gate2060(.a(gate97inter0), .b(s_216), .O(gate97inter1));
  and2  gate2061(.a(G350), .b(G19), .O(gate97inter2));
  inv1  gate2062(.a(s_216), .O(gate97inter3));
  inv1  gate2063(.a(s_217), .O(gate97inter4));
  nand2 gate2064(.a(gate97inter4), .b(gate97inter3), .O(gate97inter5));
  nor2  gate2065(.a(gate97inter5), .b(gate97inter2), .O(gate97inter6));
  inv1  gate2066(.a(G19), .O(gate97inter7));
  inv1  gate2067(.a(G350), .O(gate97inter8));
  nand2 gate2068(.a(gate97inter8), .b(gate97inter7), .O(gate97inter9));
  nand2 gate2069(.a(s_217), .b(gate97inter3), .O(gate97inter10));
  nor2  gate2070(.a(gate97inter10), .b(gate97inter9), .O(gate97inter11));
  nor2  gate2071(.a(gate97inter11), .b(gate97inter6), .O(gate97inter12));
  nand2 gate2072(.a(gate97inter12), .b(gate97inter1), .O(G418));
nand2 gate98( .a(G23), .b(G350), .O(G419) );

  xor2  gate1387(.a(G353), .b(G27), .O(gate99inter0));
  nand2 gate1388(.a(gate99inter0), .b(s_120), .O(gate99inter1));
  and2  gate1389(.a(G353), .b(G27), .O(gate99inter2));
  inv1  gate1390(.a(s_120), .O(gate99inter3));
  inv1  gate1391(.a(s_121), .O(gate99inter4));
  nand2 gate1392(.a(gate99inter4), .b(gate99inter3), .O(gate99inter5));
  nor2  gate1393(.a(gate99inter5), .b(gate99inter2), .O(gate99inter6));
  inv1  gate1394(.a(G27), .O(gate99inter7));
  inv1  gate1395(.a(G353), .O(gate99inter8));
  nand2 gate1396(.a(gate99inter8), .b(gate99inter7), .O(gate99inter9));
  nand2 gate1397(.a(s_121), .b(gate99inter3), .O(gate99inter10));
  nor2  gate1398(.a(gate99inter10), .b(gate99inter9), .O(gate99inter11));
  nor2  gate1399(.a(gate99inter11), .b(gate99inter6), .O(gate99inter12));
  nand2 gate1400(.a(gate99inter12), .b(gate99inter1), .O(G420));
nand2 gate100( .a(G31), .b(G353), .O(G421) );

  xor2  gate2381(.a(G356), .b(G20), .O(gate101inter0));
  nand2 gate2382(.a(gate101inter0), .b(s_262), .O(gate101inter1));
  and2  gate2383(.a(G356), .b(G20), .O(gate101inter2));
  inv1  gate2384(.a(s_262), .O(gate101inter3));
  inv1  gate2385(.a(s_263), .O(gate101inter4));
  nand2 gate2386(.a(gate101inter4), .b(gate101inter3), .O(gate101inter5));
  nor2  gate2387(.a(gate101inter5), .b(gate101inter2), .O(gate101inter6));
  inv1  gate2388(.a(G20), .O(gate101inter7));
  inv1  gate2389(.a(G356), .O(gate101inter8));
  nand2 gate2390(.a(gate101inter8), .b(gate101inter7), .O(gate101inter9));
  nand2 gate2391(.a(s_263), .b(gate101inter3), .O(gate101inter10));
  nor2  gate2392(.a(gate101inter10), .b(gate101inter9), .O(gate101inter11));
  nor2  gate2393(.a(gate101inter11), .b(gate101inter6), .O(gate101inter12));
  nand2 gate2394(.a(gate101inter12), .b(gate101inter1), .O(G422));
nand2 gate102( .a(G24), .b(G356), .O(G423) );

  xor2  gate603(.a(G359), .b(G28), .O(gate103inter0));
  nand2 gate604(.a(gate103inter0), .b(s_8), .O(gate103inter1));
  and2  gate605(.a(G359), .b(G28), .O(gate103inter2));
  inv1  gate606(.a(s_8), .O(gate103inter3));
  inv1  gate607(.a(s_9), .O(gate103inter4));
  nand2 gate608(.a(gate103inter4), .b(gate103inter3), .O(gate103inter5));
  nor2  gate609(.a(gate103inter5), .b(gate103inter2), .O(gate103inter6));
  inv1  gate610(.a(G28), .O(gate103inter7));
  inv1  gate611(.a(G359), .O(gate103inter8));
  nand2 gate612(.a(gate103inter8), .b(gate103inter7), .O(gate103inter9));
  nand2 gate613(.a(s_9), .b(gate103inter3), .O(gate103inter10));
  nor2  gate614(.a(gate103inter10), .b(gate103inter9), .O(gate103inter11));
  nor2  gate615(.a(gate103inter11), .b(gate103inter6), .O(gate103inter12));
  nand2 gate616(.a(gate103inter12), .b(gate103inter1), .O(G424));
nand2 gate104( .a(G32), .b(G359), .O(G425) );
nand2 gate105( .a(G362), .b(G363), .O(G426) );
nand2 gate106( .a(G364), .b(G365), .O(G429) );
nand2 gate107( .a(G366), .b(G367), .O(G432) );
nand2 gate108( .a(G368), .b(G369), .O(G435) );
nand2 gate109( .a(G370), .b(G371), .O(G438) );

  xor2  gate813(.a(G373), .b(G372), .O(gate110inter0));
  nand2 gate814(.a(gate110inter0), .b(s_38), .O(gate110inter1));
  and2  gate815(.a(G373), .b(G372), .O(gate110inter2));
  inv1  gate816(.a(s_38), .O(gate110inter3));
  inv1  gate817(.a(s_39), .O(gate110inter4));
  nand2 gate818(.a(gate110inter4), .b(gate110inter3), .O(gate110inter5));
  nor2  gate819(.a(gate110inter5), .b(gate110inter2), .O(gate110inter6));
  inv1  gate820(.a(G372), .O(gate110inter7));
  inv1  gate821(.a(G373), .O(gate110inter8));
  nand2 gate822(.a(gate110inter8), .b(gate110inter7), .O(gate110inter9));
  nand2 gate823(.a(s_39), .b(gate110inter3), .O(gate110inter10));
  nor2  gate824(.a(gate110inter10), .b(gate110inter9), .O(gate110inter11));
  nor2  gate825(.a(gate110inter11), .b(gate110inter6), .O(gate110inter12));
  nand2 gate826(.a(gate110inter12), .b(gate110inter1), .O(G441));
nand2 gate111( .a(G374), .b(G375), .O(G444) );
nand2 gate112( .a(G376), .b(G377), .O(G447) );

  xor2  gate1331(.a(G379), .b(G378), .O(gate113inter0));
  nand2 gate1332(.a(gate113inter0), .b(s_112), .O(gate113inter1));
  and2  gate1333(.a(G379), .b(G378), .O(gate113inter2));
  inv1  gate1334(.a(s_112), .O(gate113inter3));
  inv1  gate1335(.a(s_113), .O(gate113inter4));
  nand2 gate1336(.a(gate113inter4), .b(gate113inter3), .O(gate113inter5));
  nor2  gate1337(.a(gate113inter5), .b(gate113inter2), .O(gate113inter6));
  inv1  gate1338(.a(G378), .O(gate113inter7));
  inv1  gate1339(.a(G379), .O(gate113inter8));
  nand2 gate1340(.a(gate113inter8), .b(gate113inter7), .O(gate113inter9));
  nand2 gate1341(.a(s_113), .b(gate113inter3), .O(gate113inter10));
  nor2  gate1342(.a(gate113inter10), .b(gate113inter9), .O(gate113inter11));
  nor2  gate1343(.a(gate113inter11), .b(gate113inter6), .O(gate113inter12));
  nand2 gate1344(.a(gate113inter12), .b(gate113inter1), .O(G450));
nand2 gate114( .a(G380), .b(G381), .O(G453) );
nand2 gate115( .a(G382), .b(G383), .O(G456) );
nand2 gate116( .a(G384), .b(G385), .O(G459) );
nand2 gate117( .a(G386), .b(G387), .O(G462) );
nand2 gate118( .a(G388), .b(G389), .O(G465) );

  xor2  gate1863(.a(G391), .b(G390), .O(gate119inter0));
  nand2 gate1864(.a(gate119inter0), .b(s_188), .O(gate119inter1));
  and2  gate1865(.a(G391), .b(G390), .O(gate119inter2));
  inv1  gate1866(.a(s_188), .O(gate119inter3));
  inv1  gate1867(.a(s_189), .O(gate119inter4));
  nand2 gate1868(.a(gate119inter4), .b(gate119inter3), .O(gate119inter5));
  nor2  gate1869(.a(gate119inter5), .b(gate119inter2), .O(gate119inter6));
  inv1  gate1870(.a(G390), .O(gate119inter7));
  inv1  gate1871(.a(G391), .O(gate119inter8));
  nand2 gate1872(.a(gate119inter8), .b(gate119inter7), .O(gate119inter9));
  nand2 gate1873(.a(s_189), .b(gate119inter3), .O(gate119inter10));
  nor2  gate1874(.a(gate119inter10), .b(gate119inter9), .O(gate119inter11));
  nor2  gate1875(.a(gate119inter11), .b(gate119inter6), .O(gate119inter12));
  nand2 gate1876(.a(gate119inter12), .b(gate119inter1), .O(G468));

  xor2  gate2465(.a(G393), .b(G392), .O(gate120inter0));
  nand2 gate2466(.a(gate120inter0), .b(s_274), .O(gate120inter1));
  and2  gate2467(.a(G393), .b(G392), .O(gate120inter2));
  inv1  gate2468(.a(s_274), .O(gate120inter3));
  inv1  gate2469(.a(s_275), .O(gate120inter4));
  nand2 gate2470(.a(gate120inter4), .b(gate120inter3), .O(gate120inter5));
  nor2  gate2471(.a(gate120inter5), .b(gate120inter2), .O(gate120inter6));
  inv1  gate2472(.a(G392), .O(gate120inter7));
  inv1  gate2473(.a(G393), .O(gate120inter8));
  nand2 gate2474(.a(gate120inter8), .b(gate120inter7), .O(gate120inter9));
  nand2 gate2475(.a(s_275), .b(gate120inter3), .O(gate120inter10));
  nor2  gate2476(.a(gate120inter10), .b(gate120inter9), .O(gate120inter11));
  nor2  gate2477(.a(gate120inter11), .b(gate120inter6), .O(gate120inter12));
  nand2 gate2478(.a(gate120inter12), .b(gate120inter1), .O(G471));

  xor2  gate1443(.a(G395), .b(G394), .O(gate121inter0));
  nand2 gate1444(.a(gate121inter0), .b(s_128), .O(gate121inter1));
  and2  gate1445(.a(G395), .b(G394), .O(gate121inter2));
  inv1  gate1446(.a(s_128), .O(gate121inter3));
  inv1  gate1447(.a(s_129), .O(gate121inter4));
  nand2 gate1448(.a(gate121inter4), .b(gate121inter3), .O(gate121inter5));
  nor2  gate1449(.a(gate121inter5), .b(gate121inter2), .O(gate121inter6));
  inv1  gate1450(.a(G394), .O(gate121inter7));
  inv1  gate1451(.a(G395), .O(gate121inter8));
  nand2 gate1452(.a(gate121inter8), .b(gate121inter7), .O(gate121inter9));
  nand2 gate1453(.a(s_129), .b(gate121inter3), .O(gate121inter10));
  nor2  gate1454(.a(gate121inter10), .b(gate121inter9), .O(gate121inter11));
  nor2  gate1455(.a(gate121inter11), .b(gate121inter6), .O(gate121inter12));
  nand2 gate1456(.a(gate121inter12), .b(gate121inter1), .O(G474));
nand2 gate122( .a(G396), .b(G397), .O(G477) );
nand2 gate123( .a(G398), .b(G399), .O(G480) );

  xor2  gate1877(.a(G401), .b(G400), .O(gate124inter0));
  nand2 gate1878(.a(gate124inter0), .b(s_190), .O(gate124inter1));
  and2  gate1879(.a(G401), .b(G400), .O(gate124inter2));
  inv1  gate1880(.a(s_190), .O(gate124inter3));
  inv1  gate1881(.a(s_191), .O(gate124inter4));
  nand2 gate1882(.a(gate124inter4), .b(gate124inter3), .O(gate124inter5));
  nor2  gate1883(.a(gate124inter5), .b(gate124inter2), .O(gate124inter6));
  inv1  gate1884(.a(G400), .O(gate124inter7));
  inv1  gate1885(.a(G401), .O(gate124inter8));
  nand2 gate1886(.a(gate124inter8), .b(gate124inter7), .O(gate124inter9));
  nand2 gate1887(.a(s_191), .b(gate124inter3), .O(gate124inter10));
  nor2  gate1888(.a(gate124inter10), .b(gate124inter9), .O(gate124inter11));
  nor2  gate1889(.a(gate124inter11), .b(gate124inter6), .O(gate124inter12));
  nand2 gate1890(.a(gate124inter12), .b(gate124inter1), .O(G483));

  xor2  gate1415(.a(G403), .b(G402), .O(gate125inter0));
  nand2 gate1416(.a(gate125inter0), .b(s_124), .O(gate125inter1));
  and2  gate1417(.a(G403), .b(G402), .O(gate125inter2));
  inv1  gate1418(.a(s_124), .O(gate125inter3));
  inv1  gate1419(.a(s_125), .O(gate125inter4));
  nand2 gate1420(.a(gate125inter4), .b(gate125inter3), .O(gate125inter5));
  nor2  gate1421(.a(gate125inter5), .b(gate125inter2), .O(gate125inter6));
  inv1  gate1422(.a(G402), .O(gate125inter7));
  inv1  gate1423(.a(G403), .O(gate125inter8));
  nand2 gate1424(.a(gate125inter8), .b(gate125inter7), .O(gate125inter9));
  nand2 gate1425(.a(s_125), .b(gate125inter3), .O(gate125inter10));
  nor2  gate1426(.a(gate125inter10), .b(gate125inter9), .O(gate125inter11));
  nor2  gate1427(.a(gate125inter11), .b(gate125inter6), .O(gate125inter12));
  nand2 gate1428(.a(gate125inter12), .b(gate125inter1), .O(G486));
nand2 gate126( .a(G404), .b(G405), .O(G489) );

  xor2  gate785(.a(G407), .b(G406), .O(gate127inter0));
  nand2 gate786(.a(gate127inter0), .b(s_34), .O(gate127inter1));
  and2  gate787(.a(G407), .b(G406), .O(gate127inter2));
  inv1  gate788(.a(s_34), .O(gate127inter3));
  inv1  gate789(.a(s_35), .O(gate127inter4));
  nand2 gate790(.a(gate127inter4), .b(gate127inter3), .O(gate127inter5));
  nor2  gate791(.a(gate127inter5), .b(gate127inter2), .O(gate127inter6));
  inv1  gate792(.a(G406), .O(gate127inter7));
  inv1  gate793(.a(G407), .O(gate127inter8));
  nand2 gate794(.a(gate127inter8), .b(gate127inter7), .O(gate127inter9));
  nand2 gate795(.a(s_35), .b(gate127inter3), .O(gate127inter10));
  nor2  gate796(.a(gate127inter10), .b(gate127inter9), .O(gate127inter11));
  nor2  gate797(.a(gate127inter11), .b(gate127inter6), .O(gate127inter12));
  nand2 gate798(.a(gate127inter12), .b(gate127inter1), .O(G492));
nand2 gate128( .a(G408), .b(G409), .O(G495) );
nand2 gate129( .a(G410), .b(G411), .O(G498) );

  xor2  gate1765(.a(G413), .b(G412), .O(gate130inter0));
  nand2 gate1766(.a(gate130inter0), .b(s_174), .O(gate130inter1));
  and2  gate1767(.a(G413), .b(G412), .O(gate130inter2));
  inv1  gate1768(.a(s_174), .O(gate130inter3));
  inv1  gate1769(.a(s_175), .O(gate130inter4));
  nand2 gate1770(.a(gate130inter4), .b(gate130inter3), .O(gate130inter5));
  nor2  gate1771(.a(gate130inter5), .b(gate130inter2), .O(gate130inter6));
  inv1  gate1772(.a(G412), .O(gate130inter7));
  inv1  gate1773(.a(G413), .O(gate130inter8));
  nand2 gate1774(.a(gate130inter8), .b(gate130inter7), .O(gate130inter9));
  nand2 gate1775(.a(s_175), .b(gate130inter3), .O(gate130inter10));
  nor2  gate1776(.a(gate130inter10), .b(gate130inter9), .O(gate130inter11));
  nor2  gate1777(.a(gate130inter11), .b(gate130inter6), .O(gate130inter12));
  nand2 gate1778(.a(gate130inter12), .b(gate130inter1), .O(G501));
nand2 gate131( .a(G414), .b(G415), .O(G504) );
nand2 gate132( .a(G416), .b(G417), .O(G507) );

  xor2  gate1429(.a(G419), .b(G418), .O(gate133inter0));
  nand2 gate1430(.a(gate133inter0), .b(s_126), .O(gate133inter1));
  and2  gate1431(.a(G419), .b(G418), .O(gate133inter2));
  inv1  gate1432(.a(s_126), .O(gate133inter3));
  inv1  gate1433(.a(s_127), .O(gate133inter4));
  nand2 gate1434(.a(gate133inter4), .b(gate133inter3), .O(gate133inter5));
  nor2  gate1435(.a(gate133inter5), .b(gate133inter2), .O(gate133inter6));
  inv1  gate1436(.a(G418), .O(gate133inter7));
  inv1  gate1437(.a(G419), .O(gate133inter8));
  nand2 gate1438(.a(gate133inter8), .b(gate133inter7), .O(gate133inter9));
  nand2 gate1439(.a(s_127), .b(gate133inter3), .O(gate133inter10));
  nor2  gate1440(.a(gate133inter10), .b(gate133inter9), .O(gate133inter11));
  nor2  gate1441(.a(gate133inter11), .b(gate133inter6), .O(gate133inter12));
  nand2 gate1442(.a(gate133inter12), .b(gate133inter1), .O(G510));

  xor2  gate1611(.a(G421), .b(G420), .O(gate134inter0));
  nand2 gate1612(.a(gate134inter0), .b(s_152), .O(gate134inter1));
  and2  gate1613(.a(G421), .b(G420), .O(gate134inter2));
  inv1  gate1614(.a(s_152), .O(gate134inter3));
  inv1  gate1615(.a(s_153), .O(gate134inter4));
  nand2 gate1616(.a(gate134inter4), .b(gate134inter3), .O(gate134inter5));
  nor2  gate1617(.a(gate134inter5), .b(gate134inter2), .O(gate134inter6));
  inv1  gate1618(.a(G420), .O(gate134inter7));
  inv1  gate1619(.a(G421), .O(gate134inter8));
  nand2 gate1620(.a(gate134inter8), .b(gate134inter7), .O(gate134inter9));
  nand2 gate1621(.a(s_153), .b(gate134inter3), .O(gate134inter10));
  nor2  gate1622(.a(gate134inter10), .b(gate134inter9), .O(gate134inter11));
  nor2  gate1623(.a(gate134inter11), .b(gate134inter6), .O(gate134inter12));
  nand2 gate1624(.a(gate134inter12), .b(gate134inter1), .O(G513));
nand2 gate135( .a(G422), .b(G423), .O(G516) );
nand2 gate136( .a(G424), .b(G425), .O(G519) );

  xor2  gate2311(.a(G429), .b(G426), .O(gate137inter0));
  nand2 gate2312(.a(gate137inter0), .b(s_252), .O(gate137inter1));
  and2  gate2313(.a(G429), .b(G426), .O(gate137inter2));
  inv1  gate2314(.a(s_252), .O(gate137inter3));
  inv1  gate2315(.a(s_253), .O(gate137inter4));
  nand2 gate2316(.a(gate137inter4), .b(gate137inter3), .O(gate137inter5));
  nor2  gate2317(.a(gate137inter5), .b(gate137inter2), .O(gate137inter6));
  inv1  gate2318(.a(G426), .O(gate137inter7));
  inv1  gate2319(.a(G429), .O(gate137inter8));
  nand2 gate2320(.a(gate137inter8), .b(gate137inter7), .O(gate137inter9));
  nand2 gate2321(.a(s_253), .b(gate137inter3), .O(gate137inter10));
  nor2  gate2322(.a(gate137inter10), .b(gate137inter9), .O(gate137inter11));
  nor2  gate2323(.a(gate137inter11), .b(gate137inter6), .O(gate137inter12));
  nand2 gate2324(.a(gate137inter12), .b(gate137inter1), .O(G522));
nand2 gate138( .a(G432), .b(G435), .O(G525) );

  xor2  gate2577(.a(G441), .b(G438), .O(gate139inter0));
  nand2 gate2578(.a(gate139inter0), .b(s_290), .O(gate139inter1));
  and2  gate2579(.a(G441), .b(G438), .O(gate139inter2));
  inv1  gate2580(.a(s_290), .O(gate139inter3));
  inv1  gate2581(.a(s_291), .O(gate139inter4));
  nand2 gate2582(.a(gate139inter4), .b(gate139inter3), .O(gate139inter5));
  nor2  gate2583(.a(gate139inter5), .b(gate139inter2), .O(gate139inter6));
  inv1  gate2584(.a(G438), .O(gate139inter7));
  inv1  gate2585(.a(G441), .O(gate139inter8));
  nand2 gate2586(.a(gate139inter8), .b(gate139inter7), .O(gate139inter9));
  nand2 gate2587(.a(s_291), .b(gate139inter3), .O(gate139inter10));
  nor2  gate2588(.a(gate139inter10), .b(gate139inter9), .O(gate139inter11));
  nor2  gate2589(.a(gate139inter11), .b(gate139inter6), .O(gate139inter12));
  nand2 gate2590(.a(gate139inter12), .b(gate139inter1), .O(G528));

  xor2  gate2185(.a(G447), .b(G444), .O(gate140inter0));
  nand2 gate2186(.a(gate140inter0), .b(s_234), .O(gate140inter1));
  and2  gate2187(.a(G447), .b(G444), .O(gate140inter2));
  inv1  gate2188(.a(s_234), .O(gate140inter3));
  inv1  gate2189(.a(s_235), .O(gate140inter4));
  nand2 gate2190(.a(gate140inter4), .b(gate140inter3), .O(gate140inter5));
  nor2  gate2191(.a(gate140inter5), .b(gate140inter2), .O(gate140inter6));
  inv1  gate2192(.a(G444), .O(gate140inter7));
  inv1  gate2193(.a(G447), .O(gate140inter8));
  nand2 gate2194(.a(gate140inter8), .b(gate140inter7), .O(gate140inter9));
  nand2 gate2195(.a(s_235), .b(gate140inter3), .O(gate140inter10));
  nor2  gate2196(.a(gate140inter10), .b(gate140inter9), .O(gate140inter11));
  nor2  gate2197(.a(gate140inter11), .b(gate140inter6), .O(gate140inter12));
  nand2 gate2198(.a(gate140inter12), .b(gate140inter1), .O(G531));
nand2 gate141( .a(G450), .b(G453), .O(G534) );
nand2 gate142( .a(G456), .b(G459), .O(G537) );

  xor2  gate1891(.a(G465), .b(G462), .O(gate143inter0));
  nand2 gate1892(.a(gate143inter0), .b(s_192), .O(gate143inter1));
  and2  gate1893(.a(G465), .b(G462), .O(gate143inter2));
  inv1  gate1894(.a(s_192), .O(gate143inter3));
  inv1  gate1895(.a(s_193), .O(gate143inter4));
  nand2 gate1896(.a(gate143inter4), .b(gate143inter3), .O(gate143inter5));
  nor2  gate1897(.a(gate143inter5), .b(gate143inter2), .O(gate143inter6));
  inv1  gate1898(.a(G462), .O(gate143inter7));
  inv1  gate1899(.a(G465), .O(gate143inter8));
  nand2 gate1900(.a(gate143inter8), .b(gate143inter7), .O(gate143inter9));
  nand2 gate1901(.a(s_193), .b(gate143inter3), .O(gate143inter10));
  nor2  gate1902(.a(gate143inter10), .b(gate143inter9), .O(gate143inter11));
  nor2  gate1903(.a(gate143inter11), .b(gate143inter6), .O(gate143inter12));
  nand2 gate1904(.a(gate143inter12), .b(gate143inter1), .O(G540));

  xor2  gate645(.a(G471), .b(G468), .O(gate144inter0));
  nand2 gate646(.a(gate144inter0), .b(s_14), .O(gate144inter1));
  and2  gate647(.a(G471), .b(G468), .O(gate144inter2));
  inv1  gate648(.a(s_14), .O(gate144inter3));
  inv1  gate649(.a(s_15), .O(gate144inter4));
  nand2 gate650(.a(gate144inter4), .b(gate144inter3), .O(gate144inter5));
  nor2  gate651(.a(gate144inter5), .b(gate144inter2), .O(gate144inter6));
  inv1  gate652(.a(G468), .O(gate144inter7));
  inv1  gate653(.a(G471), .O(gate144inter8));
  nand2 gate654(.a(gate144inter8), .b(gate144inter7), .O(gate144inter9));
  nand2 gate655(.a(s_15), .b(gate144inter3), .O(gate144inter10));
  nor2  gate656(.a(gate144inter10), .b(gate144inter9), .O(gate144inter11));
  nor2  gate657(.a(gate144inter11), .b(gate144inter6), .O(gate144inter12));
  nand2 gate658(.a(gate144inter12), .b(gate144inter1), .O(G543));

  xor2  gate2241(.a(G477), .b(G474), .O(gate145inter0));
  nand2 gate2242(.a(gate145inter0), .b(s_242), .O(gate145inter1));
  and2  gate2243(.a(G477), .b(G474), .O(gate145inter2));
  inv1  gate2244(.a(s_242), .O(gate145inter3));
  inv1  gate2245(.a(s_243), .O(gate145inter4));
  nand2 gate2246(.a(gate145inter4), .b(gate145inter3), .O(gate145inter5));
  nor2  gate2247(.a(gate145inter5), .b(gate145inter2), .O(gate145inter6));
  inv1  gate2248(.a(G474), .O(gate145inter7));
  inv1  gate2249(.a(G477), .O(gate145inter8));
  nand2 gate2250(.a(gate145inter8), .b(gate145inter7), .O(gate145inter9));
  nand2 gate2251(.a(s_243), .b(gate145inter3), .O(gate145inter10));
  nor2  gate2252(.a(gate145inter10), .b(gate145inter9), .O(gate145inter11));
  nor2  gate2253(.a(gate145inter11), .b(gate145inter6), .O(gate145inter12));
  nand2 gate2254(.a(gate145inter12), .b(gate145inter1), .O(G546));
nand2 gate146( .a(G480), .b(G483), .O(G549) );
nand2 gate147( .a(G486), .b(G489), .O(G552) );
nand2 gate148( .a(G492), .b(G495), .O(G555) );
nand2 gate149( .a(G498), .b(G501), .O(G558) );
nand2 gate150( .a(G504), .b(G507), .O(G561) );

  xor2  gate1513(.a(G513), .b(G510), .O(gate151inter0));
  nand2 gate1514(.a(gate151inter0), .b(s_138), .O(gate151inter1));
  and2  gate1515(.a(G513), .b(G510), .O(gate151inter2));
  inv1  gate1516(.a(s_138), .O(gate151inter3));
  inv1  gate1517(.a(s_139), .O(gate151inter4));
  nand2 gate1518(.a(gate151inter4), .b(gate151inter3), .O(gate151inter5));
  nor2  gate1519(.a(gate151inter5), .b(gate151inter2), .O(gate151inter6));
  inv1  gate1520(.a(G510), .O(gate151inter7));
  inv1  gate1521(.a(G513), .O(gate151inter8));
  nand2 gate1522(.a(gate151inter8), .b(gate151inter7), .O(gate151inter9));
  nand2 gate1523(.a(s_139), .b(gate151inter3), .O(gate151inter10));
  nor2  gate1524(.a(gate151inter10), .b(gate151inter9), .O(gate151inter11));
  nor2  gate1525(.a(gate151inter11), .b(gate151inter6), .O(gate151inter12));
  nand2 gate1526(.a(gate151inter12), .b(gate151inter1), .O(G564));
nand2 gate152( .a(G516), .b(G519), .O(G567) );
nand2 gate153( .a(G426), .b(G522), .O(G570) );
nand2 gate154( .a(G429), .b(G522), .O(G571) );

  xor2  gate2297(.a(G525), .b(G432), .O(gate155inter0));
  nand2 gate2298(.a(gate155inter0), .b(s_250), .O(gate155inter1));
  and2  gate2299(.a(G525), .b(G432), .O(gate155inter2));
  inv1  gate2300(.a(s_250), .O(gate155inter3));
  inv1  gate2301(.a(s_251), .O(gate155inter4));
  nand2 gate2302(.a(gate155inter4), .b(gate155inter3), .O(gate155inter5));
  nor2  gate2303(.a(gate155inter5), .b(gate155inter2), .O(gate155inter6));
  inv1  gate2304(.a(G432), .O(gate155inter7));
  inv1  gate2305(.a(G525), .O(gate155inter8));
  nand2 gate2306(.a(gate155inter8), .b(gate155inter7), .O(gate155inter9));
  nand2 gate2307(.a(s_251), .b(gate155inter3), .O(gate155inter10));
  nor2  gate2308(.a(gate155inter10), .b(gate155inter9), .O(gate155inter11));
  nor2  gate2309(.a(gate155inter11), .b(gate155inter6), .O(gate155inter12));
  nand2 gate2310(.a(gate155inter12), .b(gate155inter1), .O(G572));

  xor2  gate2563(.a(G525), .b(G435), .O(gate156inter0));
  nand2 gate2564(.a(gate156inter0), .b(s_288), .O(gate156inter1));
  and2  gate2565(.a(G525), .b(G435), .O(gate156inter2));
  inv1  gate2566(.a(s_288), .O(gate156inter3));
  inv1  gate2567(.a(s_289), .O(gate156inter4));
  nand2 gate2568(.a(gate156inter4), .b(gate156inter3), .O(gate156inter5));
  nor2  gate2569(.a(gate156inter5), .b(gate156inter2), .O(gate156inter6));
  inv1  gate2570(.a(G435), .O(gate156inter7));
  inv1  gate2571(.a(G525), .O(gate156inter8));
  nand2 gate2572(.a(gate156inter8), .b(gate156inter7), .O(gate156inter9));
  nand2 gate2573(.a(s_289), .b(gate156inter3), .O(gate156inter10));
  nor2  gate2574(.a(gate156inter10), .b(gate156inter9), .O(gate156inter11));
  nor2  gate2575(.a(gate156inter11), .b(gate156inter6), .O(gate156inter12));
  nand2 gate2576(.a(gate156inter12), .b(gate156inter1), .O(G573));
nand2 gate157( .a(G438), .b(G528), .O(G574) );

  xor2  gate2339(.a(G528), .b(G441), .O(gate158inter0));
  nand2 gate2340(.a(gate158inter0), .b(s_256), .O(gate158inter1));
  and2  gate2341(.a(G528), .b(G441), .O(gate158inter2));
  inv1  gate2342(.a(s_256), .O(gate158inter3));
  inv1  gate2343(.a(s_257), .O(gate158inter4));
  nand2 gate2344(.a(gate158inter4), .b(gate158inter3), .O(gate158inter5));
  nor2  gate2345(.a(gate158inter5), .b(gate158inter2), .O(gate158inter6));
  inv1  gate2346(.a(G441), .O(gate158inter7));
  inv1  gate2347(.a(G528), .O(gate158inter8));
  nand2 gate2348(.a(gate158inter8), .b(gate158inter7), .O(gate158inter9));
  nand2 gate2349(.a(s_257), .b(gate158inter3), .O(gate158inter10));
  nor2  gate2350(.a(gate158inter10), .b(gate158inter9), .O(gate158inter11));
  nor2  gate2351(.a(gate158inter11), .b(gate158inter6), .O(gate158inter12));
  nand2 gate2352(.a(gate158inter12), .b(gate158inter1), .O(G575));

  xor2  gate1135(.a(G531), .b(G444), .O(gate159inter0));
  nand2 gate1136(.a(gate159inter0), .b(s_84), .O(gate159inter1));
  and2  gate1137(.a(G531), .b(G444), .O(gate159inter2));
  inv1  gate1138(.a(s_84), .O(gate159inter3));
  inv1  gate1139(.a(s_85), .O(gate159inter4));
  nand2 gate1140(.a(gate159inter4), .b(gate159inter3), .O(gate159inter5));
  nor2  gate1141(.a(gate159inter5), .b(gate159inter2), .O(gate159inter6));
  inv1  gate1142(.a(G444), .O(gate159inter7));
  inv1  gate1143(.a(G531), .O(gate159inter8));
  nand2 gate1144(.a(gate159inter8), .b(gate159inter7), .O(gate159inter9));
  nand2 gate1145(.a(s_85), .b(gate159inter3), .O(gate159inter10));
  nor2  gate1146(.a(gate159inter10), .b(gate159inter9), .O(gate159inter11));
  nor2  gate1147(.a(gate159inter11), .b(gate159inter6), .O(gate159inter12));
  nand2 gate1148(.a(gate159inter12), .b(gate159inter1), .O(G576));
nand2 gate160( .a(G447), .b(G531), .O(G577) );
nand2 gate161( .a(G450), .b(G534), .O(G578) );

  xor2  gate1667(.a(G534), .b(G453), .O(gate162inter0));
  nand2 gate1668(.a(gate162inter0), .b(s_160), .O(gate162inter1));
  and2  gate1669(.a(G534), .b(G453), .O(gate162inter2));
  inv1  gate1670(.a(s_160), .O(gate162inter3));
  inv1  gate1671(.a(s_161), .O(gate162inter4));
  nand2 gate1672(.a(gate162inter4), .b(gate162inter3), .O(gate162inter5));
  nor2  gate1673(.a(gate162inter5), .b(gate162inter2), .O(gate162inter6));
  inv1  gate1674(.a(G453), .O(gate162inter7));
  inv1  gate1675(.a(G534), .O(gate162inter8));
  nand2 gate1676(.a(gate162inter8), .b(gate162inter7), .O(gate162inter9));
  nand2 gate1677(.a(s_161), .b(gate162inter3), .O(gate162inter10));
  nor2  gate1678(.a(gate162inter10), .b(gate162inter9), .O(gate162inter11));
  nor2  gate1679(.a(gate162inter11), .b(gate162inter6), .O(gate162inter12));
  nand2 gate1680(.a(gate162inter12), .b(gate162inter1), .O(G579));
nand2 gate163( .a(G456), .b(G537), .O(G580) );
nand2 gate164( .a(G459), .b(G537), .O(G581) );
nand2 gate165( .a(G462), .b(G540), .O(G582) );

  xor2  gate995(.a(G540), .b(G465), .O(gate166inter0));
  nand2 gate996(.a(gate166inter0), .b(s_64), .O(gate166inter1));
  and2  gate997(.a(G540), .b(G465), .O(gate166inter2));
  inv1  gate998(.a(s_64), .O(gate166inter3));
  inv1  gate999(.a(s_65), .O(gate166inter4));
  nand2 gate1000(.a(gate166inter4), .b(gate166inter3), .O(gate166inter5));
  nor2  gate1001(.a(gate166inter5), .b(gate166inter2), .O(gate166inter6));
  inv1  gate1002(.a(G465), .O(gate166inter7));
  inv1  gate1003(.a(G540), .O(gate166inter8));
  nand2 gate1004(.a(gate166inter8), .b(gate166inter7), .O(gate166inter9));
  nand2 gate1005(.a(s_65), .b(gate166inter3), .O(gate166inter10));
  nor2  gate1006(.a(gate166inter10), .b(gate166inter9), .O(gate166inter11));
  nor2  gate1007(.a(gate166inter11), .b(gate166inter6), .O(gate166inter12));
  nand2 gate1008(.a(gate166inter12), .b(gate166inter1), .O(G583));
nand2 gate167( .a(G468), .b(G543), .O(G584) );
nand2 gate168( .a(G471), .b(G543), .O(G585) );
nand2 gate169( .a(G474), .b(G546), .O(G586) );
nand2 gate170( .a(G477), .b(G546), .O(G587) );
nand2 gate171( .a(G480), .b(G549), .O(G588) );

  xor2  gate841(.a(G549), .b(G483), .O(gate172inter0));
  nand2 gate842(.a(gate172inter0), .b(s_42), .O(gate172inter1));
  and2  gate843(.a(G549), .b(G483), .O(gate172inter2));
  inv1  gate844(.a(s_42), .O(gate172inter3));
  inv1  gate845(.a(s_43), .O(gate172inter4));
  nand2 gate846(.a(gate172inter4), .b(gate172inter3), .O(gate172inter5));
  nor2  gate847(.a(gate172inter5), .b(gate172inter2), .O(gate172inter6));
  inv1  gate848(.a(G483), .O(gate172inter7));
  inv1  gate849(.a(G549), .O(gate172inter8));
  nand2 gate850(.a(gate172inter8), .b(gate172inter7), .O(gate172inter9));
  nand2 gate851(.a(s_43), .b(gate172inter3), .O(gate172inter10));
  nor2  gate852(.a(gate172inter10), .b(gate172inter9), .O(gate172inter11));
  nor2  gate853(.a(gate172inter11), .b(gate172inter6), .O(gate172inter12));
  nand2 gate854(.a(gate172inter12), .b(gate172inter1), .O(G589));

  xor2  gate673(.a(G552), .b(G486), .O(gate173inter0));
  nand2 gate674(.a(gate173inter0), .b(s_18), .O(gate173inter1));
  and2  gate675(.a(G552), .b(G486), .O(gate173inter2));
  inv1  gate676(.a(s_18), .O(gate173inter3));
  inv1  gate677(.a(s_19), .O(gate173inter4));
  nand2 gate678(.a(gate173inter4), .b(gate173inter3), .O(gate173inter5));
  nor2  gate679(.a(gate173inter5), .b(gate173inter2), .O(gate173inter6));
  inv1  gate680(.a(G486), .O(gate173inter7));
  inv1  gate681(.a(G552), .O(gate173inter8));
  nand2 gate682(.a(gate173inter8), .b(gate173inter7), .O(gate173inter9));
  nand2 gate683(.a(s_19), .b(gate173inter3), .O(gate173inter10));
  nor2  gate684(.a(gate173inter10), .b(gate173inter9), .O(gate173inter11));
  nor2  gate685(.a(gate173inter11), .b(gate173inter6), .O(gate173inter12));
  nand2 gate686(.a(gate173inter12), .b(gate173inter1), .O(G590));
nand2 gate174( .a(G489), .b(G552), .O(G591) );
nand2 gate175( .a(G492), .b(G555), .O(G592) );

  xor2  gate575(.a(G555), .b(G495), .O(gate176inter0));
  nand2 gate576(.a(gate176inter0), .b(s_4), .O(gate176inter1));
  and2  gate577(.a(G555), .b(G495), .O(gate176inter2));
  inv1  gate578(.a(s_4), .O(gate176inter3));
  inv1  gate579(.a(s_5), .O(gate176inter4));
  nand2 gate580(.a(gate176inter4), .b(gate176inter3), .O(gate176inter5));
  nor2  gate581(.a(gate176inter5), .b(gate176inter2), .O(gate176inter6));
  inv1  gate582(.a(G495), .O(gate176inter7));
  inv1  gate583(.a(G555), .O(gate176inter8));
  nand2 gate584(.a(gate176inter8), .b(gate176inter7), .O(gate176inter9));
  nand2 gate585(.a(s_5), .b(gate176inter3), .O(gate176inter10));
  nor2  gate586(.a(gate176inter10), .b(gate176inter9), .O(gate176inter11));
  nor2  gate587(.a(gate176inter11), .b(gate176inter6), .O(gate176inter12));
  nand2 gate588(.a(gate176inter12), .b(gate176inter1), .O(G593));

  xor2  gate869(.a(G558), .b(G498), .O(gate177inter0));
  nand2 gate870(.a(gate177inter0), .b(s_46), .O(gate177inter1));
  and2  gate871(.a(G558), .b(G498), .O(gate177inter2));
  inv1  gate872(.a(s_46), .O(gate177inter3));
  inv1  gate873(.a(s_47), .O(gate177inter4));
  nand2 gate874(.a(gate177inter4), .b(gate177inter3), .O(gate177inter5));
  nor2  gate875(.a(gate177inter5), .b(gate177inter2), .O(gate177inter6));
  inv1  gate876(.a(G498), .O(gate177inter7));
  inv1  gate877(.a(G558), .O(gate177inter8));
  nand2 gate878(.a(gate177inter8), .b(gate177inter7), .O(gate177inter9));
  nand2 gate879(.a(s_47), .b(gate177inter3), .O(gate177inter10));
  nor2  gate880(.a(gate177inter10), .b(gate177inter9), .O(gate177inter11));
  nor2  gate881(.a(gate177inter11), .b(gate177inter6), .O(gate177inter12));
  nand2 gate882(.a(gate177inter12), .b(gate177inter1), .O(G594));
nand2 gate178( .a(G501), .b(G558), .O(G595) );
nand2 gate179( .a(G504), .b(G561), .O(G596) );
nand2 gate180( .a(G507), .b(G561), .O(G597) );

  xor2  gate1625(.a(G564), .b(G510), .O(gate181inter0));
  nand2 gate1626(.a(gate181inter0), .b(s_154), .O(gate181inter1));
  and2  gate1627(.a(G564), .b(G510), .O(gate181inter2));
  inv1  gate1628(.a(s_154), .O(gate181inter3));
  inv1  gate1629(.a(s_155), .O(gate181inter4));
  nand2 gate1630(.a(gate181inter4), .b(gate181inter3), .O(gate181inter5));
  nor2  gate1631(.a(gate181inter5), .b(gate181inter2), .O(gate181inter6));
  inv1  gate1632(.a(G510), .O(gate181inter7));
  inv1  gate1633(.a(G564), .O(gate181inter8));
  nand2 gate1634(.a(gate181inter8), .b(gate181inter7), .O(gate181inter9));
  nand2 gate1635(.a(s_155), .b(gate181inter3), .O(gate181inter10));
  nor2  gate1636(.a(gate181inter10), .b(gate181inter9), .O(gate181inter11));
  nor2  gate1637(.a(gate181inter11), .b(gate181inter6), .O(gate181inter12));
  nand2 gate1638(.a(gate181inter12), .b(gate181inter1), .O(G598));

  xor2  gate771(.a(G564), .b(G513), .O(gate182inter0));
  nand2 gate772(.a(gate182inter0), .b(s_32), .O(gate182inter1));
  and2  gate773(.a(G564), .b(G513), .O(gate182inter2));
  inv1  gate774(.a(s_32), .O(gate182inter3));
  inv1  gate775(.a(s_33), .O(gate182inter4));
  nand2 gate776(.a(gate182inter4), .b(gate182inter3), .O(gate182inter5));
  nor2  gate777(.a(gate182inter5), .b(gate182inter2), .O(gate182inter6));
  inv1  gate778(.a(G513), .O(gate182inter7));
  inv1  gate779(.a(G564), .O(gate182inter8));
  nand2 gate780(.a(gate182inter8), .b(gate182inter7), .O(gate182inter9));
  nand2 gate781(.a(s_33), .b(gate182inter3), .O(gate182inter10));
  nor2  gate782(.a(gate182inter10), .b(gate182inter9), .O(gate182inter11));
  nor2  gate783(.a(gate182inter11), .b(gate182inter6), .O(gate182inter12));
  nand2 gate784(.a(gate182inter12), .b(gate182inter1), .O(G599));
nand2 gate183( .a(G516), .b(G567), .O(G600) );
nand2 gate184( .a(G519), .b(G567), .O(G601) );
nand2 gate185( .a(G570), .b(G571), .O(G602) );
nand2 gate186( .a(G572), .b(G573), .O(G607) );
nand2 gate187( .a(G574), .b(G575), .O(G612) );
nand2 gate188( .a(G576), .b(G577), .O(G617) );
nand2 gate189( .a(G578), .b(G579), .O(G622) );
nand2 gate190( .a(G580), .b(G581), .O(G627) );
nand2 gate191( .a(G582), .b(G583), .O(G632) );
nand2 gate192( .a(G584), .b(G585), .O(G637) );
nand2 gate193( .a(G586), .b(G587), .O(G642) );

  xor2  gate1919(.a(G589), .b(G588), .O(gate194inter0));
  nand2 gate1920(.a(gate194inter0), .b(s_196), .O(gate194inter1));
  and2  gate1921(.a(G589), .b(G588), .O(gate194inter2));
  inv1  gate1922(.a(s_196), .O(gate194inter3));
  inv1  gate1923(.a(s_197), .O(gate194inter4));
  nand2 gate1924(.a(gate194inter4), .b(gate194inter3), .O(gate194inter5));
  nor2  gate1925(.a(gate194inter5), .b(gate194inter2), .O(gate194inter6));
  inv1  gate1926(.a(G588), .O(gate194inter7));
  inv1  gate1927(.a(G589), .O(gate194inter8));
  nand2 gate1928(.a(gate194inter8), .b(gate194inter7), .O(gate194inter9));
  nand2 gate1929(.a(s_197), .b(gate194inter3), .O(gate194inter10));
  nor2  gate1930(.a(gate194inter10), .b(gate194inter9), .O(gate194inter11));
  nor2  gate1931(.a(gate194inter11), .b(gate194inter6), .O(gate194inter12));
  nand2 gate1932(.a(gate194inter12), .b(gate194inter1), .O(G645));

  xor2  gate547(.a(G591), .b(G590), .O(gate195inter0));
  nand2 gate548(.a(gate195inter0), .b(s_0), .O(gate195inter1));
  and2  gate549(.a(G591), .b(G590), .O(gate195inter2));
  inv1  gate550(.a(s_0), .O(gate195inter3));
  inv1  gate551(.a(s_1), .O(gate195inter4));
  nand2 gate552(.a(gate195inter4), .b(gate195inter3), .O(gate195inter5));
  nor2  gate553(.a(gate195inter5), .b(gate195inter2), .O(gate195inter6));
  inv1  gate554(.a(G590), .O(gate195inter7));
  inv1  gate555(.a(G591), .O(gate195inter8));
  nand2 gate556(.a(gate195inter8), .b(gate195inter7), .O(gate195inter9));
  nand2 gate557(.a(s_1), .b(gate195inter3), .O(gate195inter10));
  nor2  gate558(.a(gate195inter10), .b(gate195inter9), .O(gate195inter11));
  nor2  gate559(.a(gate195inter11), .b(gate195inter6), .O(gate195inter12));
  nand2 gate560(.a(gate195inter12), .b(gate195inter1), .O(G648));
nand2 gate196( .a(G592), .b(G593), .O(G651) );

  xor2  gate617(.a(G595), .b(G594), .O(gate197inter0));
  nand2 gate618(.a(gate197inter0), .b(s_10), .O(gate197inter1));
  and2  gate619(.a(G595), .b(G594), .O(gate197inter2));
  inv1  gate620(.a(s_10), .O(gate197inter3));
  inv1  gate621(.a(s_11), .O(gate197inter4));
  nand2 gate622(.a(gate197inter4), .b(gate197inter3), .O(gate197inter5));
  nor2  gate623(.a(gate197inter5), .b(gate197inter2), .O(gate197inter6));
  inv1  gate624(.a(G594), .O(gate197inter7));
  inv1  gate625(.a(G595), .O(gate197inter8));
  nand2 gate626(.a(gate197inter8), .b(gate197inter7), .O(gate197inter9));
  nand2 gate627(.a(s_11), .b(gate197inter3), .O(gate197inter10));
  nor2  gate628(.a(gate197inter10), .b(gate197inter9), .O(gate197inter11));
  nor2  gate629(.a(gate197inter11), .b(gate197inter6), .O(gate197inter12));
  nand2 gate630(.a(gate197inter12), .b(gate197inter1), .O(G654));

  xor2  gate897(.a(G597), .b(G596), .O(gate198inter0));
  nand2 gate898(.a(gate198inter0), .b(s_50), .O(gate198inter1));
  and2  gate899(.a(G597), .b(G596), .O(gate198inter2));
  inv1  gate900(.a(s_50), .O(gate198inter3));
  inv1  gate901(.a(s_51), .O(gate198inter4));
  nand2 gate902(.a(gate198inter4), .b(gate198inter3), .O(gate198inter5));
  nor2  gate903(.a(gate198inter5), .b(gate198inter2), .O(gate198inter6));
  inv1  gate904(.a(G596), .O(gate198inter7));
  inv1  gate905(.a(G597), .O(gate198inter8));
  nand2 gate906(.a(gate198inter8), .b(gate198inter7), .O(gate198inter9));
  nand2 gate907(.a(s_51), .b(gate198inter3), .O(gate198inter10));
  nor2  gate908(.a(gate198inter10), .b(gate198inter9), .O(gate198inter11));
  nor2  gate909(.a(gate198inter11), .b(gate198inter6), .O(gate198inter12));
  nand2 gate910(.a(gate198inter12), .b(gate198inter1), .O(G657));
nand2 gate199( .a(G598), .b(G599), .O(G660) );

  xor2  gate2325(.a(G601), .b(G600), .O(gate200inter0));
  nand2 gate2326(.a(gate200inter0), .b(s_254), .O(gate200inter1));
  and2  gate2327(.a(G601), .b(G600), .O(gate200inter2));
  inv1  gate2328(.a(s_254), .O(gate200inter3));
  inv1  gate2329(.a(s_255), .O(gate200inter4));
  nand2 gate2330(.a(gate200inter4), .b(gate200inter3), .O(gate200inter5));
  nor2  gate2331(.a(gate200inter5), .b(gate200inter2), .O(gate200inter6));
  inv1  gate2332(.a(G600), .O(gate200inter7));
  inv1  gate2333(.a(G601), .O(gate200inter8));
  nand2 gate2334(.a(gate200inter8), .b(gate200inter7), .O(gate200inter9));
  nand2 gate2335(.a(s_255), .b(gate200inter3), .O(gate200inter10));
  nor2  gate2336(.a(gate200inter10), .b(gate200inter9), .O(gate200inter11));
  nor2  gate2337(.a(gate200inter11), .b(gate200inter6), .O(gate200inter12));
  nand2 gate2338(.a(gate200inter12), .b(gate200inter1), .O(G663));
nand2 gate201( .a(G602), .b(G607), .O(G666) );
nand2 gate202( .a(G612), .b(G617), .O(G669) );
nand2 gate203( .a(G602), .b(G612), .O(G672) );
nand2 gate204( .a(G607), .b(G617), .O(G675) );

  xor2  gate2451(.a(G627), .b(G622), .O(gate205inter0));
  nand2 gate2452(.a(gate205inter0), .b(s_272), .O(gate205inter1));
  and2  gate2453(.a(G627), .b(G622), .O(gate205inter2));
  inv1  gate2454(.a(s_272), .O(gate205inter3));
  inv1  gate2455(.a(s_273), .O(gate205inter4));
  nand2 gate2456(.a(gate205inter4), .b(gate205inter3), .O(gate205inter5));
  nor2  gate2457(.a(gate205inter5), .b(gate205inter2), .O(gate205inter6));
  inv1  gate2458(.a(G622), .O(gate205inter7));
  inv1  gate2459(.a(G627), .O(gate205inter8));
  nand2 gate2460(.a(gate205inter8), .b(gate205inter7), .O(gate205inter9));
  nand2 gate2461(.a(s_273), .b(gate205inter3), .O(gate205inter10));
  nor2  gate2462(.a(gate205inter10), .b(gate205inter9), .O(gate205inter11));
  nor2  gate2463(.a(gate205inter11), .b(gate205inter6), .O(gate205inter12));
  nand2 gate2464(.a(gate205inter12), .b(gate205inter1), .O(G678));

  xor2  gate1065(.a(G637), .b(G632), .O(gate206inter0));
  nand2 gate1066(.a(gate206inter0), .b(s_74), .O(gate206inter1));
  and2  gate1067(.a(G637), .b(G632), .O(gate206inter2));
  inv1  gate1068(.a(s_74), .O(gate206inter3));
  inv1  gate1069(.a(s_75), .O(gate206inter4));
  nand2 gate1070(.a(gate206inter4), .b(gate206inter3), .O(gate206inter5));
  nor2  gate1071(.a(gate206inter5), .b(gate206inter2), .O(gate206inter6));
  inv1  gate1072(.a(G632), .O(gate206inter7));
  inv1  gate1073(.a(G637), .O(gate206inter8));
  nand2 gate1074(.a(gate206inter8), .b(gate206inter7), .O(gate206inter9));
  nand2 gate1075(.a(s_75), .b(gate206inter3), .O(gate206inter10));
  nor2  gate1076(.a(gate206inter10), .b(gate206inter9), .O(gate206inter11));
  nor2  gate1077(.a(gate206inter11), .b(gate206inter6), .O(gate206inter12));
  nand2 gate1078(.a(gate206inter12), .b(gate206inter1), .O(G681));
nand2 gate207( .a(G622), .b(G632), .O(G684) );
nand2 gate208( .a(G627), .b(G637), .O(G687) );
nand2 gate209( .a(G602), .b(G666), .O(G690) );
nand2 gate210( .a(G607), .b(G666), .O(G691) );

  xor2  gate2423(.a(G669), .b(G612), .O(gate211inter0));
  nand2 gate2424(.a(gate211inter0), .b(s_268), .O(gate211inter1));
  and2  gate2425(.a(G669), .b(G612), .O(gate211inter2));
  inv1  gate2426(.a(s_268), .O(gate211inter3));
  inv1  gate2427(.a(s_269), .O(gate211inter4));
  nand2 gate2428(.a(gate211inter4), .b(gate211inter3), .O(gate211inter5));
  nor2  gate2429(.a(gate211inter5), .b(gate211inter2), .O(gate211inter6));
  inv1  gate2430(.a(G612), .O(gate211inter7));
  inv1  gate2431(.a(G669), .O(gate211inter8));
  nand2 gate2432(.a(gate211inter8), .b(gate211inter7), .O(gate211inter9));
  nand2 gate2433(.a(s_269), .b(gate211inter3), .O(gate211inter10));
  nor2  gate2434(.a(gate211inter10), .b(gate211inter9), .O(gate211inter11));
  nor2  gate2435(.a(gate211inter11), .b(gate211inter6), .O(gate211inter12));
  nand2 gate2436(.a(gate211inter12), .b(gate211inter1), .O(G692));

  xor2  gate1737(.a(G669), .b(G617), .O(gate212inter0));
  nand2 gate1738(.a(gate212inter0), .b(s_170), .O(gate212inter1));
  and2  gate1739(.a(G669), .b(G617), .O(gate212inter2));
  inv1  gate1740(.a(s_170), .O(gate212inter3));
  inv1  gate1741(.a(s_171), .O(gate212inter4));
  nand2 gate1742(.a(gate212inter4), .b(gate212inter3), .O(gate212inter5));
  nor2  gate1743(.a(gate212inter5), .b(gate212inter2), .O(gate212inter6));
  inv1  gate1744(.a(G617), .O(gate212inter7));
  inv1  gate1745(.a(G669), .O(gate212inter8));
  nand2 gate1746(.a(gate212inter8), .b(gate212inter7), .O(gate212inter9));
  nand2 gate1747(.a(s_171), .b(gate212inter3), .O(gate212inter10));
  nor2  gate1748(.a(gate212inter10), .b(gate212inter9), .O(gate212inter11));
  nor2  gate1749(.a(gate212inter11), .b(gate212inter6), .O(gate212inter12));
  nand2 gate1750(.a(gate212inter12), .b(gate212inter1), .O(G693));
nand2 gate213( .a(G602), .b(G672), .O(G694) );

  xor2  gate883(.a(G672), .b(G612), .O(gate214inter0));
  nand2 gate884(.a(gate214inter0), .b(s_48), .O(gate214inter1));
  and2  gate885(.a(G672), .b(G612), .O(gate214inter2));
  inv1  gate886(.a(s_48), .O(gate214inter3));
  inv1  gate887(.a(s_49), .O(gate214inter4));
  nand2 gate888(.a(gate214inter4), .b(gate214inter3), .O(gate214inter5));
  nor2  gate889(.a(gate214inter5), .b(gate214inter2), .O(gate214inter6));
  inv1  gate890(.a(G612), .O(gate214inter7));
  inv1  gate891(.a(G672), .O(gate214inter8));
  nand2 gate892(.a(gate214inter8), .b(gate214inter7), .O(gate214inter9));
  nand2 gate893(.a(s_49), .b(gate214inter3), .O(gate214inter10));
  nor2  gate894(.a(gate214inter10), .b(gate214inter9), .O(gate214inter11));
  nor2  gate895(.a(gate214inter11), .b(gate214inter6), .O(gate214inter12));
  nand2 gate896(.a(gate214inter12), .b(gate214inter1), .O(G695));
nand2 gate215( .a(G607), .b(G675), .O(G696) );
nand2 gate216( .a(G617), .b(G675), .O(G697) );
nand2 gate217( .a(G622), .b(G678), .O(G698) );
nand2 gate218( .a(G627), .b(G678), .O(G699) );

  xor2  gate2367(.a(G681), .b(G632), .O(gate219inter0));
  nand2 gate2368(.a(gate219inter0), .b(s_260), .O(gate219inter1));
  and2  gate2369(.a(G681), .b(G632), .O(gate219inter2));
  inv1  gate2370(.a(s_260), .O(gate219inter3));
  inv1  gate2371(.a(s_261), .O(gate219inter4));
  nand2 gate2372(.a(gate219inter4), .b(gate219inter3), .O(gate219inter5));
  nor2  gate2373(.a(gate219inter5), .b(gate219inter2), .O(gate219inter6));
  inv1  gate2374(.a(G632), .O(gate219inter7));
  inv1  gate2375(.a(G681), .O(gate219inter8));
  nand2 gate2376(.a(gate219inter8), .b(gate219inter7), .O(gate219inter9));
  nand2 gate2377(.a(s_261), .b(gate219inter3), .O(gate219inter10));
  nor2  gate2378(.a(gate219inter10), .b(gate219inter9), .O(gate219inter11));
  nor2  gate2379(.a(gate219inter11), .b(gate219inter6), .O(gate219inter12));
  nand2 gate2380(.a(gate219inter12), .b(gate219inter1), .O(G700));
nand2 gate220( .a(G637), .b(G681), .O(G701) );

  xor2  gate1723(.a(G684), .b(G622), .O(gate221inter0));
  nand2 gate1724(.a(gate221inter0), .b(s_168), .O(gate221inter1));
  and2  gate1725(.a(G684), .b(G622), .O(gate221inter2));
  inv1  gate1726(.a(s_168), .O(gate221inter3));
  inv1  gate1727(.a(s_169), .O(gate221inter4));
  nand2 gate1728(.a(gate221inter4), .b(gate221inter3), .O(gate221inter5));
  nor2  gate1729(.a(gate221inter5), .b(gate221inter2), .O(gate221inter6));
  inv1  gate1730(.a(G622), .O(gate221inter7));
  inv1  gate1731(.a(G684), .O(gate221inter8));
  nand2 gate1732(.a(gate221inter8), .b(gate221inter7), .O(gate221inter9));
  nand2 gate1733(.a(s_169), .b(gate221inter3), .O(gate221inter10));
  nor2  gate1734(.a(gate221inter10), .b(gate221inter9), .O(gate221inter11));
  nor2  gate1735(.a(gate221inter11), .b(gate221inter6), .O(gate221inter12));
  nand2 gate1736(.a(gate221inter12), .b(gate221inter1), .O(G702));
nand2 gate222( .a(G632), .b(G684), .O(G703) );
nand2 gate223( .a(G627), .b(G687), .O(G704) );
nand2 gate224( .a(G637), .b(G687), .O(G705) );

  xor2  gate1639(.a(G691), .b(G690), .O(gate225inter0));
  nand2 gate1640(.a(gate225inter0), .b(s_156), .O(gate225inter1));
  and2  gate1641(.a(G691), .b(G690), .O(gate225inter2));
  inv1  gate1642(.a(s_156), .O(gate225inter3));
  inv1  gate1643(.a(s_157), .O(gate225inter4));
  nand2 gate1644(.a(gate225inter4), .b(gate225inter3), .O(gate225inter5));
  nor2  gate1645(.a(gate225inter5), .b(gate225inter2), .O(gate225inter6));
  inv1  gate1646(.a(G690), .O(gate225inter7));
  inv1  gate1647(.a(G691), .O(gate225inter8));
  nand2 gate1648(.a(gate225inter8), .b(gate225inter7), .O(gate225inter9));
  nand2 gate1649(.a(s_157), .b(gate225inter3), .O(gate225inter10));
  nor2  gate1650(.a(gate225inter10), .b(gate225inter9), .O(gate225inter11));
  nor2  gate1651(.a(gate225inter11), .b(gate225inter6), .O(gate225inter12));
  nand2 gate1652(.a(gate225inter12), .b(gate225inter1), .O(G706));
nand2 gate226( .a(G692), .b(G693), .O(G709) );
nand2 gate227( .a(G694), .b(G695), .O(G712) );
nand2 gate228( .a(G696), .b(G697), .O(G715) );
nand2 gate229( .a(G698), .b(G699), .O(G718) );
nand2 gate230( .a(G700), .b(G701), .O(G721) );
nand2 gate231( .a(G702), .b(G703), .O(G724) );
nand2 gate232( .a(G704), .b(G705), .O(G727) );
nand2 gate233( .a(G242), .b(G718), .O(G730) );
nand2 gate234( .a(G245), .b(G721), .O(G733) );

  xor2  gate2227(.a(G724), .b(G248), .O(gate235inter0));
  nand2 gate2228(.a(gate235inter0), .b(s_240), .O(gate235inter1));
  and2  gate2229(.a(G724), .b(G248), .O(gate235inter2));
  inv1  gate2230(.a(s_240), .O(gate235inter3));
  inv1  gate2231(.a(s_241), .O(gate235inter4));
  nand2 gate2232(.a(gate235inter4), .b(gate235inter3), .O(gate235inter5));
  nor2  gate2233(.a(gate235inter5), .b(gate235inter2), .O(gate235inter6));
  inv1  gate2234(.a(G248), .O(gate235inter7));
  inv1  gate2235(.a(G724), .O(gate235inter8));
  nand2 gate2236(.a(gate235inter8), .b(gate235inter7), .O(gate235inter9));
  nand2 gate2237(.a(s_241), .b(gate235inter3), .O(gate235inter10));
  nor2  gate2238(.a(gate235inter10), .b(gate235inter9), .O(gate235inter11));
  nor2  gate2239(.a(gate235inter11), .b(gate235inter6), .O(gate235inter12));
  nand2 gate2240(.a(gate235inter12), .b(gate235inter1), .O(G736));

  xor2  gate2045(.a(G727), .b(G251), .O(gate236inter0));
  nand2 gate2046(.a(gate236inter0), .b(s_214), .O(gate236inter1));
  and2  gate2047(.a(G727), .b(G251), .O(gate236inter2));
  inv1  gate2048(.a(s_214), .O(gate236inter3));
  inv1  gate2049(.a(s_215), .O(gate236inter4));
  nand2 gate2050(.a(gate236inter4), .b(gate236inter3), .O(gate236inter5));
  nor2  gate2051(.a(gate236inter5), .b(gate236inter2), .O(gate236inter6));
  inv1  gate2052(.a(G251), .O(gate236inter7));
  inv1  gate2053(.a(G727), .O(gate236inter8));
  nand2 gate2054(.a(gate236inter8), .b(gate236inter7), .O(gate236inter9));
  nand2 gate2055(.a(s_215), .b(gate236inter3), .O(gate236inter10));
  nor2  gate2056(.a(gate236inter10), .b(gate236inter9), .O(gate236inter11));
  nor2  gate2057(.a(gate236inter11), .b(gate236inter6), .O(gate236inter12));
  nand2 gate2058(.a(gate236inter12), .b(gate236inter1), .O(G739));

  xor2  gate1121(.a(G706), .b(G254), .O(gate237inter0));
  nand2 gate1122(.a(gate237inter0), .b(s_82), .O(gate237inter1));
  and2  gate1123(.a(G706), .b(G254), .O(gate237inter2));
  inv1  gate1124(.a(s_82), .O(gate237inter3));
  inv1  gate1125(.a(s_83), .O(gate237inter4));
  nand2 gate1126(.a(gate237inter4), .b(gate237inter3), .O(gate237inter5));
  nor2  gate1127(.a(gate237inter5), .b(gate237inter2), .O(gate237inter6));
  inv1  gate1128(.a(G254), .O(gate237inter7));
  inv1  gate1129(.a(G706), .O(gate237inter8));
  nand2 gate1130(.a(gate237inter8), .b(gate237inter7), .O(gate237inter9));
  nand2 gate1131(.a(s_83), .b(gate237inter3), .O(gate237inter10));
  nor2  gate1132(.a(gate237inter10), .b(gate237inter9), .O(gate237inter11));
  nor2  gate1133(.a(gate237inter11), .b(gate237inter6), .O(gate237inter12));
  nand2 gate1134(.a(gate237inter12), .b(gate237inter1), .O(G742));

  xor2  gate1037(.a(G709), .b(G257), .O(gate238inter0));
  nand2 gate1038(.a(gate238inter0), .b(s_70), .O(gate238inter1));
  and2  gate1039(.a(G709), .b(G257), .O(gate238inter2));
  inv1  gate1040(.a(s_70), .O(gate238inter3));
  inv1  gate1041(.a(s_71), .O(gate238inter4));
  nand2 gate1042(.a(gate238inter4), .b(gate238inter3), .O(gate238inter5));
  nor2  gate1043(.a(gate238inter5), .b(gate238inter2), .O(gate238inter6));
  inv1  gate1044(.a(G257), .O(gate238inter7));
  inv1  gate1045(.a(G709), .O(gate238inter8));
  nand2 gate1046(.a(gate238inter8), .b(gate238inter7), .O(gate238inter9));
  nand2 gate1047(.a(s_71), .b(gate238inter3), .O(gate238inter10));
  nor2  gate1048(.a(gate238inter10), .b(gate238inter9), .O(gate238inter11));
  nor2  gate1049(.a(gate238inter11), .b(gate238inter6), .O(gate238inter12));
  nand2 gate1050(.a(gate238inter12), .b(gate238inter1), .O(G745));
nand2 gate239( .a(G260), .b(G712), .O(G748) );
nand2 gate240( .a(G263), .b(G715), .O(G751) );

  xor2  gate2143(.a(G730), .b(G242), .O(gate241inter0));
  nand2 gate2144(.a(gate241inter0), .b(s_228), .O(gate241inter1));
  and2  gate2145(.a(G730), .b(G242), .O(gate241inter2));
  inv1  gate2146(.a(s_228), .O(gate241inter3));
  inv1  gate2147(.a(s_229), .O(gate241inter4));
  nand2 gate2148(.a(gate241inter4), .b(gate241inter3), .O(gate241inter5));
  nor2  gate2149(.a(gate241inter5), .b(gate241inter2), .O(gate241inter6));
  inv1  gate2150(.a(G242), .O(gate241inter7));
  inv1  gate2151(.a(G730), .O(gate241inter8));
  nand2 gate2152(.a(gate241inter8), .b(gate241inter7), .O(gate241inter9));
  nand2 gate2153(.a(s_229), .b(gate241inter3), .O(gate241inter10));
  nor2  gate2154(.a(gate241inter10), .b(gate241inter9), .O(gate241inter11));
  nor2  gate2155(.a(gate241inter11), .b(gate241inter6), .O(gate241inter12));
  nand2 gate2156(.a(gate241inter12), .b(gate241inter1), .O(G754));

  xor2  gate589(.a(G730), .b(G718), .O(gate242inter0));
  nand2 gate590(.a(gate242inter0), .b(s_6), .O(gate242inter1));
  and2  gate591(.a(G730), .b(G718), .O(gate242inter2));
  inv1  gate592(.a(s_6), .O(gate242inter3));
  inv1  gate593(.a(s_7), .O(gate242inter4));
  nand2 gate594(.a(gate242inter4), .b(gate242inter3), .O(gate242inter5));
  nor2  gate595(.a(gate242inter5), .b(gate242inter2), .O(gate242inter6));
  inv1  gate596(.a(G718), .O(gate242inter7));
  inv1  gate597(.a(G730), .O(gate242inter8));
  nand2 gate598(.a(gate242inter8), .b(gate242inter7), .O(gate242inter9));
  nand2 gate599(.a(s_7), .b(gate242inter3), .O(gate242inter10));
  nor2  gate600(.a(gate242inter10), .b(gate242inter9), .O(gate242inter11));
  nor2  gate601(.a(gate242inter11), .b(gate242inter6), .O(gate242inter12));
  nand2 gate602(.a(gate242inter12), .b(gate242inter1), .O(G755));

  xor2  gate1849(.a(G733), .b(G245), .O(gate243inter0));
  nand2 gate1850(.a(gate243inter0), .b(s_186), .O(gate243inter1));
  and2  gate1851(.a(G733), .b(G245), .O(gate243inter2));
  inv1  gate1852(.a(s_186), .O(gate243inter3));
  inv1  gate1853(.a(s_187), .O(gate243inter4));
  nand2 gate1854(.a(gate243inter4), .b(gate243inter3), .O(gate243inter5));
  nor2  gate1855(.a(gate243inter5), .b(gate243inter2), .O(gate243inter6));
  inv1  gate1856(.a(G245), .O(gate243inter7));
  inv1  gate1857(.a(G733), .O(gate243inter8));
  nand2 gate1858(.a(gate243inter8), .b(gate243inter7), .O(gate243inter9));
  nand2 gate1859(.a(s_187), .b(gate243inter3), .O(gate243inter10));
  nor2  gate1860(.a(gate243inter10), .b(gate243inter9), .O(gate243inter11));
  nor2  gate1861(.a(gate243inter11), .b(gate243inter6), .O(gate243inter12));
  nand2 gate1862(.a(gate243inter12), .b(gate243inter1), .O(G756));
nand2 gate244( .a(G721), .b(G733), .O(G757) );
nand2 gate245( .a(G248), .b(G736), .O(G758) );
nand2 gate246( .a(G724), .b(G736), .O(G759) );
nand2 gate247( .a(G251), .b(G739), .O(G760) );
nand2 gate248( .a(G727), .b(G739), .O(G761) );

  xor2  gate1177(.a(G742), .b(G254), .O(gate249inter0));
  nand2 gate1178(.a(gate249inter0), .b(s_90), .O(gate249inter1));
  and2  gate1179(.a(G742), .b(G254), .O(gate249inter2));
  inv1  gate1180(.a(s_90), .O(gate249inter3));
  inv1  gate1181(.a(s_91), .O(gate249inter4));
  nand2 gate1182(.a(gate249inter4), .b(gate249inter3), .O(gate249inter5));
  nor2  gate1183(.a(gate249inter5), .b(gate249inter2), .O(gate249inter6));
  inv1  gate1184(.a(G254), .O(gate249inter7));
  inv1  gate1185(.a(G742), .O(gate249inter8));
  nand2 gate1186(.a(gate249inter8), .b(gate249inter7), .O(gate249inter9));
  nand2 gate1187(.a(s_91), .b(gate249inter3), .O(gate249inter10));
  nor2  gate1188(.a(gate249inter10), .b(gate249inter9), .O(gate249inter11));
  nor2  gate1189(.a(gate249inter11), .b(gate249inter6), .O(gate249inter12));
  nand2 gate1190(.a(gate249inter12), .b(gate249inter1), .O(G762));
nand2 gate250( .a(G706), .b(G742), .O(G763) );
nand2 gate251( .a(G257), .b(G745), .O(G764) );
nand2 gate252( .a(G709), .b(G745), .O(G765) );
nand2 gate253( .a(G260), .b(G748), .O(G766) );
nand2 gate254( .a(G712), .b(G748), .O(G767) );
nand2 gate255( .a(G263), .b(G751), .O(G768) );
nand2 gate256( .a(G715), .b(G751), .O(G769) );
nand2 gate257( .a(G754), .b(G755), .O(G770) );

  xor2  gate1009(.a(G757), .b(G756), .O(gate258inter0));
  nand2 gate1010(.a(gate258inter0), .b(s_66), .O(gate258inter1));
  and2  gate1011(.a(G757), .b(G756), .O(gate258inter2));
  inv1  gate1012(.a(s_66), .O(gate258inter3));
  inv1  gate1013(.a(s_67), .O(gate258inter4));
  nand2 gate1014(.a(gate258inter4), .b(gate258inter3), .O(gate258inter5));
  nor2  gate1015(.a(gate258inter5), .b(gate258inter2), .O(gate258inter6));
  inv1  gate1016(.a(G756), .O(gate258inter7));
  inv1  gate1017(.a(G757), .O(gate258inter8));
  nand2 gate1018(.a(gate258inter8), .b(gate258inter7), .O(gate258inter9));
  nand2 gate1019(.a(s_67), .b(gate258inter3), .O(gate258inter10));
  nor2  gate1020(.a(gate258inter10), .b(gate258inter9), .O(gate258inter11));
  nor2  gate1021(.a(gate258inter11), .b(gate258inter6), .O(gate258inter12));
  nand2 gate1022(.a(gate258inter12), .b(gate258inter1), .O(G773));
nand2 gate259( .a(G758), .b(G759), .O(G776) );
nand2 gate260( .a(G760), .b(G761), .O(G779) );
nand2 gate261( .a(G762), .b(G763), .O(G782) );
nand2 gate262( .a(G764), .b(G765), .O(G785) );
nand2 gate263( .a(G766), .b(G767), .O(G788) );
nand2 gate264( .a(G768), .b(G769), .O(G791) );
nand2 gate265( .a(G642), .b(G770), .O(G794) );
nand2 gate266( .a(G645), .b(G773), .O(G797) );

  xor2  gate757(.a(G776), .b(G648), .O(gate267inter0));
  nand2 gate758(.a(gate267inter0), .b(s_30), .O(gate267inter1));
  and2  gate759(.a(G776), .b(G648), .O(gate267inter2));
  inv1  gate760(.a(s_30), .O(gate267inter3));
  inv1  gate761(.a(s_31), .O(gate267inter4));
  nand2 gate762(.a(gate267inter4), .b(gate267inter3), .O(gate267inter5));
  nor2  gate763(.a(gate267inter5), .b(gate267inter2), .O(gate267inter6));
  inv1  gate764(.a(G648), .O(gate267inter7));
  inv1  gate765(.a(G776), .O(gate267inter8));
  nand2 gate766(.a(gate267inter8), .b(gate267inter7), .O(gate267inter9));
  nand2 gate767(.a(s_31), .b(gate267inter3), .O(gate267inter10));
  nor2  gate768(.a(gate267inter10), .b(gate267inter9), .O(gate267inter11));
  nor2  gate769(.a(gate267inter11), .b(gate267inter6), .O(gate267inter12));
  nand2 gate770(.a(gate267inter12), .b(gate267inter1), .O(G800));
nand2 gate268( .a(G651), .b(G779), .O(G803) );

  xor2  gate799(.a(G782), .b(G654), .O(gate269inter0));
  nand2 gate800(.a(gate269inter0), .b(s_36), .O(gate269inter1));
  and2  gate801(.a(G782), .b(G654), .O(gate269inter2));
  inv1  gate802(.a(s_36), .O(gate269inter3));
  inv1  gate803(.a(s_37), .O(gate269inter4));
  nand2 gate804(.a(gate269inter4), .b(gate269inter3), .O(gate269inter5));
  nor2  gate805(.a(gate269inter5), .b(gate269inter2), .O(gate269inter6));
  inv1  gate806(.a(G654), .O(gate269inter7));
  inv1  gate807(.a(G782), .O(gate269inter8));
  nand2 gate808(.a(gate269inter8), .b(gate269inter7), .O(gate269inter9));
  nand2 gate809(.a(s_37), .b(gate269inter3), .O(gate269inter10));
  nor2  gate810(.a(gate269inter10), .b(gate269inter9), .O(gate269inter11));
  nor2  gate811(.a(gate269inter11), .b(gate269inter6), .O(gate269inter12));
  nand2 gate812(.a(gate269inter12), .b(gate269inter1), .O(G806));
nand2 gate270( .a(G657), .b(G785), .O(G809) );

  xor2  gate2115(.a(G788), .b(G660), .O(gate271inter0));
  nand2 gate2116(.a(gate271inter0), .b(s_224), .O(gate271inter1));
  and2  gate2117(.a(G788), .b(G660), .O(gate271inter2));
  inv1  gate2118(.a(s_224), .O(gate271inter3));
  inv1  gate2119(.a(s_225), .O(gate271inter4));
  nand2 gate2120(.a(gate271inter4), .b(gate271inter3), .O(gate271inter5));
  nor2  gate2121(.a(gate271inter5), .b(gate271inter2), .O(gate271inter6));
  inv1  gate2122(.a(G660), .O(gate271inter7));
  inv1  gate2123(.a(G788), .O(gate271inter8));
  nand2 gate2124(.a(gate271inter8), .b(gate271inter7), .O(gate271inter9));
  nand2 gate2125(.a(s_225), .b(gate271inter3), .O(gate271inter10));
  nor2  gate2126(.a(gate271inter10), .b(gate271inter9), .O(gate271inter11));
  nor2  gate2127(.a(gate271inter11), .b(gate271inter6), .O(gate271inter12));
  nand2 gate2128(.a(gate271inter12), .b(gate271inter1), .O(G812));
nand2 gate272( .a(G663), .b(G791), .O(G815) );
nand2 gate273( .a(G642), .b(G794), .O(G818) );

  xor2  gate1345(.a(G794), .b(G770), .O(gate274inter0));
  nand2 gate1346(.a(gate274inter0), .b(s_114), .O(gate274inter1));
  and2  gate1347(.a(G794), .b(G770), .O(gate274inter2));
  inv1  gate1348(.a(s_114), .O(gate274inter3));
  inv1  gate1349(.a(s_115), .O(gate274inter4));
  nand2 gate1350(.a(gate274inter4), .b(gate274inter3), .O(gate274inter5));
  nor2  gate1351(.a(gate274inter5), .b(gate274inter2), .O(gate274inter6));
  inv1  gate1352(.a(G770), .O(gate274inter7));
  inv1  gate1353(.a(G794), .O(gate274inter8));
  nand2 gate1354(.a(gate274inter8), .b(gate274inter7), .O(gate274inter9));
  nand2 gate1355(.a(s_115), .b(gate274inter3), .O(gate274inter10));
  nor2  gate1356(.a(gate274inter10), .b(gate274inter9), .O(gate274inter11));
  nor2  gate1357(.a(gate274inter11), .b(gate274inter6), .O(gate274inter12));
  nand2 gate1358(.a(gate274inter12), .b(gate274inter1), .O(G819));
nand2 gate275( .a(G645), .b(G797), .O(G820) );
nand2 gate276( .a(G773), .b(G797), .O(G821) );
nand2 gate277( .a(G648), .b(G800), .O(G822) );
nand2 gate278( .a(G776), .b(G800), .O(G823) );
nand2 gate279( .a(G651), .b(G803), .O(G824) );
nand2 gate280( .a(G779), .b(G803), .O(G825) );

  xor2  gate2269(.a(G806), .b(G654), .O(gate281inter0));
  nand2 gate2270(.a(gate281inter0), .b(s_246), .O(gate281inter1));
  and2  gate2271(.a(G806), .b(G654), .O(gate281inter2));
  inv1  gate2272(.a(s_246), .O(gate281inter3));
  inv1  gate2273(.a(s_247), .O(gate281inter4));
  nand2 gate2274(.a(gate281inter4), .b(gate281inter3), .O(gate281inter5));
  nor2  gate2275(.a(gate281inter5), .b(gate281inter2), .O(gate281inter6));
  inv1  gate2276(.a(G654), .O(gate281inter7));
  inv1  gate2277(.a(G806), .O(gate281inter8));
  nand2 gate2278(.a(gate281inter8), .b(gate281inter7), .O(gate281inter9));
  nand2 gate2279(.a(s_247), .b(gate281inter3), .O(gate281inter10));
  nor2  gate2280(.a(gate281inter10), .b(gate281inter9), .O(gate281inter11));
  nor2  gate2281(.a(gate281inter11), .b(gate281inter6), .O(gate281inter12));
  nand2 gate2282(.a(gate281inter12), .b(gate281inter1), .O(G826));

  xor2  gate2507(.a(G806), .b(G782), .O(gate282inter0));
  nand2 gate2508(.a(gate282inter0), .b(s_280), .O(gate282inter1));
  and2  gate2509(.a(G806), .b(G782), .O(gate282inter2));
  inv1  gate2510(.a(s_280), .O(gate282inter3));
  inv1  gate2511(.a(s_281), .O(gate282inter4));
  nand2 gate2512(.a(gate282inter4), .b(gate282inter3), .O(gate282inter5));
  nor2  gate2513(.a(gate282inter5), .b(gate282inter2), .O(gate282inter6));
  inv1  gate2514(.a(G782), .O(gate282inter7));
  inv1  gate2515(.a(G806), .O(gate282inter8));
  nand2 gate2516(.a(gate282inter8), .b(gate282inter7), .O(gate282inter9));
  nand2 gate2517(.a(s_281), .b(gate282inter3), .O(gate282inter10));
  nor2  gate2518(.a(gate282inter10), .b(gate282inter9), .O(gate282inter11));
  nor2  gate2519(.a(gate282inter11), .b(gate282inter6), .O(gate282inter12));
  nand2 gate2520(.a(gate282inter12), .b(gate282inter1), .O(G827));

  xor2  gate1807(.a(G809), .b(G657), .O(gate283inter0));
  nand2 gate1808(.a(gate283inter0), .b(s_180), .O(gate283inter1));
  and2  gate1809(.a(G809), .b(G657), .O(gate283inter2));
  inv1  gate1810(.a(s_180), .O(gate283inter3));
  inv1  gate1811(.a(s_181), .O(gate283inter4));
  nand2 gate1812(.a(gate283inter4), .b(gate283inter3), .O(gate283inter5));
  nor2  gate1813(.a(gate283inter5), .b(gate283inter2), .O(gate283inter6));
  inv1  gate1814(.a(G657), .O(gate283inter7));
  inv1  gate1815(.a(G809), .O(gate283inter8));
  nand2 gate1816(.a(gate283inter8), .b(gate283inter7), .O(gate283inter9));
  nand2 gate1817(.a(s_181), .b(gate283inter3), .O(gate283inter10));
  nor2  gate1818(.a(gate283inter10), .b(gate283inter9), .O(gate283inter11));
  nor2  gate1819(.a(gate283inter11), .b(gate283inter6), .O(gate283inter12));
  nand2 gate1820(.a(gate283inter12), .b(gate283inter1), .O(G828));
nand2 gate284( .a(G785), .b(G809), .O(G829) );
nand2 gate285( .a(G660), .b(G812), .O(G830) );
nand2 gate286( .a(G788), .b(G812), .O(G831) );
nand2 gate287( .a(G663), .b(G815), .O(G832) );

  xor2  gate2003(.a(G815), .b(G791), .O(gate288inter0));
  nand2 gate2004(.a(gate288inter0), .b(s_208), .O(gate288inter1));
  and2  gate2005(.a(G815), .b(G791), .O(gate288inter2));
  inv1  gate2006(.a(s_208), .O(gate288inter3));
  inv1  gate2007(.a(s_209), .O(gate288inter4));
  nand2 gate2008(.a(gate288inter4), .b(gate288inter3), .O(gate288inter5));
  nor2  gate2009(.a(gate288inter5), .b(gate288inter2), .O(gate288inter6));
  inv1  gate2010(.a(G791), .O(gate288inter7));
  inv1  gate2011(.a(G815), .O(gate288inter8));
  nand2 gate2012(.a(gate288inter8), .b(gate288inter7), .O(gate288inter9));
  nand2 gate2013(.a(s_209), .b(gate288inter3), .O(gate288inter10));
  nor2  gate2014(.a(gate288inter10), .b(gate288inter9), .O(gate288inter11));
  nor2  gate2015(.a(gate288inter11), .b(gate288inter6), .O(gate288inter12));
  nand2 gate2016(.a(gate288inter12), .b(gate288inter1), .O(G833));

  xor2  gate2409(.a(G819), .b(G818), .O(gate289inter0));
  nand2 gate2410(.a(gate289inter0), .b(s_266), .O(gate289inter1));
  and2  gate2411(.a(G819), .b(G818), .O(gate289inter2));
  inv1  gate2412(.a(s_266), .O(gate289inter3));
  inv1  gate2413(.a(s_267), .O(gate289inter4));
  nand2 gate2414(.a(gate289inter4), .b(gate289inter3), .O(gate289inter5));
  nor2  gate2415(.a(gate289inter5), .b(gate289inter2), .O(gate289inter6));
  inv1  gate2416(.a(G818), .O(gate289inter7));
  inv1  gate2417(.a(G819), .O(gate289inter8));
  nand2 gate2418(.a(gate289inter8), .b(gate289inter7), .O(gate289inter9));
  nand2 gate2419(.a(s_267), .b(gate289inter3), .O(gate289inter10));
  nor2  gate2420(.a(gate289inter10), .b(gate289inter9), .O(gate289inter11));
  nor2  gate2421(.a(gate289inter11), .b(gate289inter6), .O(gate289inter12));
  nand2 gate2422(.a(gate289inter12), .b(gate289inter1), .O(G834));

  xor2  gate911(.a(G821), .b(G820), .O(gate290inter0));
  nand2 gate912(.a(gate290inter0), .b(s_52), .O(gate290inter1));
  and2  gate913(.a(G821), .b(G820), .O(gate290inter2));
  inv1  gate914(.a(s_52), .O(gate290inter3));
  inv1  gate915(.a(s_53), .O(gate290inter4));
  nand2 gate916(.a(gate290inter4), .b(gate290inter3), .O(gate290inter5));
  nor2  gate917(.a(gate290inter5), .b(gate290inter2), .O(gate290inter6));
  inv1  gate918(.a(G820), .O(gate290inter7));
  inv1  gate919(.a(G821), .O(gate290inter8));
  nand2 gate920(.a(gate290inter8), .b(gate290inter7), .O(gate290inter9));
  nand2 gate921(.a(s_53), .b(gate290inter3), .O(gate290inter10));
  nor2  gate922(.a(gate290inter10), .b(gate290inter9), .O(gate290inter11));
  nor2  gate923(.a(gate290inter11), .b(gate290inter6), .O(gate290inter12));
  nand2 gate924(.a(gate290inter12), .b(gate290inter1), .O(G847));

  xor2  gate701(.a(G823), .b(G822), .O(gate291inter0));
  nand2 gate702(.a(gate291inter0), .b(s_22), .O(gate291inter1));
  and2  gate703(.a(G823), .b(G822), .O(gate291inter2));
  inv1  gate704(.a(s_22), .O(gate291inter3));
  inv1  gate705(.a(s_23), .O(gate291inter4));
  nand2 gate706(.a(gate291inter4), .b(gate291inter3), .O(gate291inter5));
  nor2  gate707(.a(gate291inter5), .b(gate291inter2), .O(gate291inter6));
  inv1  gate708(.a(G822), .O(gate291inter7));
  inv1  gate709(.a(G823), .O(gate291inter8));
  nand2 gate710(.a(gate291inter8), .b(gate291inter7), .O(gate291inter9));
  nand2 gate711(.a(s_23), .b(gate291inter3), .O(gate291inter10));
  nor2  gate712(.a(gate291inter10), .b(gate291inter9), .O(gate291inter11));
  nor2  gate713(.a(gate291inter11), .b(gate291inter6), .O(gate291inter12));
  nand2 gate714(.a(gate291inter12), .b(gate291inter1), .O(G860));

  xor2  gate729(.a(G825), .b(G824), .O(gate292inter0));
  nand2 gate730(.a(gate292inter0), .b(s_26), .O(gate292inter1));
  and2  gate731(.a(G825), .b(G824), .O(gate292inter2));
  inv1  gate732(.a(s_26), .O(gate292inter3));
  inv1  gate733(.a(s_27), .O(gate292inter4));
  nand2 gate734(.a(gate292inter4), .b(gate292inter3), .O(gate292inter5));
  nor2  gate735(.a(gate292inter5), .b(gate292inter2), .O(gate292inter6));
  inv1  gate736(.a(G824), .O(gate292inter7));
  inv1  gate737(.a(G825), .O(gate292inter8));
  nand2 gate738(.a(gate292inter8), .b(gate292inter7), .O(gate292inter9));
  nand2 gate739(.a(s_27), .b(gate292inter3), .O(gate292inter10));
  nor2  gate740(.a(gate292inter10), .b(gate292inter9), .O(gate292inter11));
  nor2  gate741(.a(gate292inter11), .b(gate292inter6), .O(gate292inter12));
  nand2 gate742(.a(gate292inter12), .b(gate292inter1), .O(G873));

  xor2  gate1317(.a(G829), .b(G828), .O(gate293inter0));
  nand2 gate1318(.a(gate293inter0), .b(s_110), .O(gate293inter1));
  and2  gate1319(.a(G829), .b(G828), .O(gate293inter2));
  inv1  gate1320(.a(s_110), .O(gate293inter3));
  inv1  gate1321(.a(s_111), .O(gate293inter4));
  nand2 gate1322(.a(gate293inter4), .b(gate293inter3), .O(gate293inter5));
  nor2  gate1323(.a(gate293inter5), .b(gate293inter2), .O(gate293inter6));
  inv1  gate1324(.a(G828), .O(gate293inter7));
  inv1  gate1325(.a(G829), .O(gate293inter8));
  nand2 gate1326(.a(gate293inter8), .b(gate293inter7), .O(gate293inter9));
  nand2 gate1327(.a(s_111), .b(gate293inter3), .O(gate293inter10));
  nor2  gate1328(.a(gate293inter10), .b(gate293inter9), .O(gate293inter11));
  nor2  gate1329(.a(gate293inter11), .b(gate293inter6), .O(gate293inter12));
  nand2 gate1330(.a(gate293inter12), .b(gate293inter1), .O(G886));

  xor2  gate2031(.a(G833), .b(G832), .O(gate294inter0));
  nand2 gate2032(.a(gate294inter0), .b(s_212), .O(gate294inter1));
  and2  gate2033(.a(G833), .b(G832), .O(gate294inter2));
  inv1  gate2034(.a(s_212), .O(gate294inter3));
  inv1  gate2035(.a(s_213), .O(gate294inter4));
  nand2 gate2036(.a(gate294inter4), .b(gate294inter3), .O(gate294inter5));
  nor2  gate2037(.a(gate294inter5), .b(gate294inter2), .O(gate294inter6));
  inv1  gate2038(.a(G832), .O(gate294inter7));
  inv1  gate2039(.a(G833), .O(gate294inter8));
  nand2 gate2040(.a(gate294inter8), .b(gate294inter7), .O(gate294inter9));
  nand2 gate2041(.a(s_213), .b(gate294inter3), .O(gate294inter10));
  nor2  gate2042(.a(gate294inter10), .b(gate294inter9), .O(gate294inter11));
  nor2  gate2043(.a(gate294inter11), .b(gate294inter6), .O(gate294inter12));
  nand2 gate2044(.a(gate294inter12), .b(gate294inter1), .O(G899));

  xor2  gate1261(.a(G831), .b(G830), .O(gate295inter0));
  nand2 gate1262(.a(gate295inter0), .b(s_102), .O(gate295inter1));
  and2  gate1263(.a(G831), .b(G830), .O(gate295inter2));
  inv1  gate1264(.a(s_102), .O(gate295inter3));
  inv1  gate1265(.a(s_103), .O(gate295inter4));
  nand2 gate1266(.a(gate295inter4), .b(gate295inter3), .O(gate295inter5));
  nor2  gate1267(.a(gate295inter5), .b(gate295inter2), .O(gate295inter6));
  inv1  gate1268(.a(G830), .O(gate295inter7));
  inv1  gate1269(.a(G831), .O(gate295inter8));
  nand2 gate1270(.a(gate295inter8), .b(gate295inter7), .O(gate295inter9));
  nand2 gate1271(.a(s_103), .b(gate295inter3), .O(gate295inter10));
  nor2  gate1272(.a(gate295inter10), .b(gate295inter9), .O(gate295inter11));
  nor2  gate1273(.a(gate295inter11), .b(gate295inter6), .O(gate295inter12));
  nand2 gate1274(.a(gate295inter12), .b(gate295inter1), .O(G912));
nand2 gate296( .a(G826), .b(G827), .O(G925) );
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );

  xor2  gate1653(.a(G1036), .b(G1), .O(gate387inter0));
  nand2 gate1654(.a(gate387inter0), .b(s_158), .O(gate387inter1));
  and2  gate1655(.a(G1036), .b(G1), .O(gate387inter2));
  inv1  gate1656(.a(s_158), .O(gate387inter3));
  inv1  gate1657(.a(s_159), .O(gate387inter4));
  nand2 gate1658(.a(gate387inter4), .b(gate387inter3), .O(gate387inter5));
  nor2  gate1659(.a(gate387inter5), .b(gate387inter2), .O(gate387inter6));
  inv1  gate1660(.a(G1), .O(gate387inter7));
  inv1  gate1661(.a(G1036), .O(gate387inter8));
  nand2 gate1662(.a(gate387inter8), .b(gate387inter7), .O(gate387inter9));
  nand2 gate1663(.a(s_159), .b(gate387inter3), .O(gate387inter10));
  nor2  gate1664(.a(gate387inter10), .b(gate387inter9), .O(gate387inter11));
  nor2  gate1665(.a(gate387inter11), .b(gate387inter6), .O(gate387inter12));
  nand2 gate1666(.a(gate387inter12), .b(gate387inter1), .O(G1132));

  xor2  gate1583(.a(G1039), .b(G2), .O(gate388inter0));
  nand2 gate1584(.a(gate388inter0), .b(s_148), .O(gate388inter1));
  and2  gate1585(.a(G1039), .b(G2), .O(gate388inter2));
  inv1  gate1586(.a(s_148), .O(gate388inter3));
  inv1  gate1587(.a(s_149), .O(gate388inter4));
  nand2 gate1588(.a(gate388inter4), .b(gate388inter3), .O(gate388inter5));
  nor2  gate1589(.a(gate388inter5), .b(gate388inter2), .O(gate388inter6));
  inv1  gate1590(.a(G2), .O(gate388inter7));
  inv1  gate1591(.a(G1039), .O(gate388inter8));
  nand2 gate1592(.a(gate388inter8), .b(gate388inter7), .O(gate388inter9));
  nand2 gate1593(.a(s_149), .b(gate388inter3), .O(gate388inter10));
  nor2  gate1594(.a(gate388inter10), .b(gate388inter9), .O(gate388inter11));
  nor2  gate1595(.a(gate388inter11), .b(gate388inter6), .O(gate388inter12));
  nand2 gate1596(.a(gate388inter12), .b(gate388inter1), .O(G1135));
nand2 gate389( .a(G3), .b(G1042), .O(G1138) );
nand2 gate390( .a(G4), .b(G1045), .O(G1141) );

  xor2  gate967(.a(G1048), .b(G5), .O(gate391inter0));
  nand2 gate968(.a(gate391inter0), .b(s_60), .O(gate391inter1));
  and2  gate969(.a(G1048), .b(G5), .O(gate391inter2));
  inv1  gate970(.a(s_60), .O(gate391inter3));
  inv1  gate971(.a(s_61), .O(gate391inter4));
  nand2 gate972(.a(gate391inter4), .b(gate391inter3), .O(gate391inter5));
  nor2  gate973(.a(gate391inter5), .b(gate391inter2), .O(gate391inter6));
  inv1  gate974(.a(G5), .O(gate391inter7));
  inv1  gate975(.a(G1048), .O(gate391inter8));
  nand2 gate976(.a(gate391inter8), .b(gate391inter7), .O(gate391inter9));
  nand2 gate977(.a(s_61), .b(gate391inter3), .O(gate391inter10));
  nor2  gate978(.a(gate391inter10), .b(gate391inter9), .O(gate391inter11));
  nor2  gate979(.a(gate391inter11), .b(gate391inter6), .O(gate391inter12));
  nand2 gate980(.a(gate391inter12), .b(gate391inter1), .O(G1144));

  xor2  gate1373(.a(G1051), .b(G6), .O(gate392inter0));
  nand2 gate1374(.a(gate392inter0), .b(s_118), .O(gate392inter1));
  and2  gate1375(.a(G1051), .b(G6), .O(gate392inter2));
  inv1  gate1376(.a(s_118), .O(gate392inter3));
  inv1  gate1377(.a(s_119), .O(gate392inter4));
  nand2 gate1378(.a(gate392inter4), .b(gate392inter3), .O(gate392inter5));
  nor2  gate1379(.a(gate392inter5), .b(gate392inter2), .O(gate392inter6));
  inv1  gate1380(.a(G6), .O(gate392inter7));
  inv1  gate1381(.a(G1051), .O(gate392inter8));
  nand2 gate1382(.a(gate392inter8), .b(gate392inter7), .O(gate392inter9));
  nand2 gate1383(.a(s_119), .b(gate392inter3), .O(gate392inter10));
  nor2  gate1384(.a(gate392inter10), .b(gate392inter9), .O(gate392inter11));
  nor2  gate1385(.a(gate392inter11), .b(gate392inter6), .O(gate392inter12));
  nand2 gate1386(.a(gate392inter12), .b(gate392inter1), .O(G1147));
nand2 gate393( .a(G7), .b(G1054), .O(G1150) );
nand2 gate394( .a(G8), .b(G1057), .O(G1153) );

  xor2  gate1359(.a(G1060), .b(G9), .O(gate395inter0));
  nand2 gate1360(.a(gate395inter0), .b(s_116), .O(gate395inter1));
  and2  gate1361(.a(G1060), .b(G9), .O(gate395inter2));
  inv1  gate1362(.a(s_116), .O(gate395inter3));
  inv1  gate1363(.a(s_117), .O(gate395inter4));
  nand2 gate1364(.a(gate395inter4), .b(gate395inter3), .O(gate395inter5));
  nor2  gate1365(.a(gate395inter5), .b(gate395inter2), .O(gate395inter6));
  inv1  gate1366(.a(G9), .O(gate395inter7));
  inv1  gate1367(.a(G1060), .O(gate395inter8));
  nand2 gate1368(.a(gate395inter8), .b(gate395inter7), .O(gate395inter9));
  nand2 gate1369(.a(s_117), .b(gate395inter3), .O(gate395inter10));
  nor2  gate1370(.a(gate395inter10), .b(gate395inter9), .O(gate395inter11));
  nor2  gate1371(.a(gate395inter11), .b(gate395inter6), .O(gate395inter12));
  nand2 gate1372(.a(gate395inter12), .b(gate395inter1), .O(G1156));

  xor2  gate1093(.a(G1063), .b(G10), .O(gate396inter0));
  nand2 gate1094(.a(gate396inter0), .b(s_78), .O(gate396inter1));
  and2  gate1095(.a(G1063), .b(G10), .O(gate396inter2));
  inv1  gate1096(.a(s_78), .O(gate396inter3));
  inv1  gate1097(.a(s_79), .O(gate396inter4));
  nand2 gate1098(.a(gate396inter4), .b(gate396inter3), .O(gate396inter5));
  nor2  gate1099(.a(gate396inter5), .b(gate396inter2), .O(gate396inter6));
  inv1  gate1100(.a(G10), .O(gate396inter7));
  inv1  gate1101(.a(G1063), .O(gate396inter8));
  nand2 gate1102(.a(gate396inter8), .b(gate396inter7), .O(gate396inter9));
  nand2 gate1103(.a(s_79), .b(gate396inter3), .O(gate396inter10));
  nor2  gate1104(.a(gate396inter10), .b(gate396inter9), .O(gate396inter11));
  nor2  gate1105(.a(gate396inter11), .b(gate396inter6), .O(gate396inter12));
  nand2 gate1106(.a(gate396inter12), .b(gate396inter1), .O(G1159));
nand2 gate397( .a(G11), .b(G1066), .O(G1162) );

  xor2  gate2017(.a(G1069), .b(G12), .O(gate398inter0));
  nand2 gate2018(.a(gate398inter0), .b(s_210), .O(gate398inter1));
  and2  gate2019(.a(G1069), .b(G12), .O(gate398inter2));
  inv1  gate2020(.a(s_210), .O(gate398inter3));
  inv1  gate2021(.a(s_211), .O(gate398inter4));
  nand2 gate2022(.a(gate398inter4), .b(gate398inter3), .O(gate398inter5));
  nor2  gate2023(.a(gate398inter5), .b(gate398inter2), .O(gate398inter6));
  inv1  gate2024(.a(G12), .O(gate398inter7));
  inv1  gate2025(.a(G1069), .O(gate398inter8));
  nand2 gate2026(.a(gate398inter8), .b(gate398inter7), .O(gate398inter9));
  nand2 gate2027(.a(s_211), .b(gate398inter3), .O(gate398inter10));
  nor2  gate2028(.a(gate398inter10), .b(gate398inter9), .O(gate398inter11));
  nor2  gate2029(.a(gate398inter11), .b(gate398inter6), .O(gate398inter12));
  nand2 gate2030(.a(gate398inter12), .b(gate398inter1), .O(G1165));
nand2 gate399( .a(G13), .b(G1072), .O(G1168) );
nand2 gate400( .a(G14), .b(G1075), .O(G1171) );
nand2 gate401( .a(G15), .b(G1078), .O(G1174) );

  xor2  gate2213(.a(G1081), .b(G16), .O(gate402inter0));
  nand2 gate2214(.a(gate402inter0), .b(s_238), .O(gate402inter1));
  and2  gate2215(.a(G1081), .b(G16), .O(gate402inter2));
  inv1  gate2216(.a(s_238), .O(gate402inter3));
  inv1  gate2217(.a(s_239), .O(gate402inter4));
  nand2 gate2218(.a(gate402inter4), .b(gate402inter3), .O(gate402inter5));
  nor2  gate2219(.a(gate402inter5), .b(gate402inter2), .O(gate402inter6));
  inv1  gate2220(.a(G16), .O(gate402inter7));
  inv1  gate2221(.a(G1081), .O(gate402inter8));
  nand2 gate2222(.a(gate402inter8), .b(gate402inter7), .O(gate402inter9));
  nand2 gate2223(.a(s_239), .b(gate402inter3), .O(gate402inter10));
  nor2  gate2224(.a(gate402inter10), .b(gate402inter9), .O(gate402inter11));
  nor2  gate2225(.a(gate402inter11), .b(gate402inter6), .O(gate402inter12));
  nand2 gate2226(.a(gate402inter12), .b(gate402inter1), .O(G1177));

  xor2  gate1149(.a(G1084), .b(G17), .O(gate403inter0));
  nand2 gate1150(.a(gate403inter0), .b(s_86), .O(gate403inter1));
  and2  gate1151(.a(G1084), .b(G17), .O(gate403inter2));
  inv1  gate1152(.a(s_86), .O(gate403inter3));
  inv1  gate1153(.a(s_87), .O(gate403inter4));
  nand2 gate1154(.a(gate403inter4), .b(gate403inter3), .O(gate403inter5));
  nor2  gate1155(.a(gate403inter5), .b(gate403inter2), .O(gate403inter6));
  inv1  gate1156(.a(G17), .O(gate403inter7));
  inv1  gate1157(.a(G1084), .O(gate403inter8));
  nand2 gate1158(.a(gate403inter8), .b(gate403inter7), .O(gate403inter9));
  nand2 gate1159(.a(s_87), .b(gate403inter3), .O(gate403inter10));
  nor2  gate1160(.a(gate403inter10), .b(gate403inter9), .O(gate403inter11));
  nor2  gate1161(.a(gate403inter11), .b(gate403inter6), .O(gate403inter12));
  nand2 gate1162(.a(gate403inter12), .b(gate403inter1), .O(G1180));

  xor2  gate1289(.a(G1087), .b(G18), .O(gate404inter0));
  nand2 gate1290(.a(gate404inter0), .b(s_106), .O(gate404inter1));
  and2  gate1291(.a(G1087), .b(G18), .O(gate404inter2));
  inv1  gate1292(.a(s_106), .O(gate404inter3));
  inv1  gate1293(.a(s_107), .O(gate404inter4));
  nand2 gate1294(.a(gate404inter4), .b(gate404inter3), .O(gate404inter5));
  nor2  gate1295(.a(gate404inter5), .b(gate404inter2), .O(gate404inter6));
  inv1  gate1296(.a(G18), .O(gate404inter7));
  inv1  gate1297(.a(G1087), .O(gate404inter8));
  nand2 gate1298(.a(gate404inter8), .b(gate404inter7), .O(gate404inter9));
  nand2 gate1299(.a(s_107), .b(gate404inter3), .O(gate404inter10));
  nor2  gate1300(.a(gate404inter10), .b(gate404inter9), .O(gate404inter11));
  nor2  gate1301(.a(gate404inter11), .b(gate404inter6), .O(gate404inter12));
  nand2 gate1302(.a(gate404inter12), .b(gate404inter1), .O(G1183));
nand2 gate405( .a(G19), .b(G1090), .O(G1186) );
nand2 gate406( .a(G20), .b(G1093), .O(G1189) );
nand2 gate407( .a(G21), .b(G1096), .O(G1192) );
nand2 gate408( .a(G22), .b(G1099), .O(G1195) );

  xor2  gate1779(.a(G1102), .b(G23), .O(gate409inter0));
  nand2 gate1780(.a(gate409inter0), .b(s_176), .O(gate409inter1));
  and2  gate1781(.a(G1102), .b(G23), .O(gate409inter2));
  inv1  gate1782(.a(s_176), .O(gate409inter3));
  inv1  gate1783(.a(s_177), .O(gate409inter4));
  nand2 gate1784(.a(gate409inter4), .b(gate409inter3), .O(gate409inter5));
  nor2  gate1785(.a(gate409inter5), .b(gate409inter2), .O(gate409inter6));
  inv1  gate1786(.a(G23), .O(gate409inter7));
  inv1  gate1787(.a(G1102), .O(gate409inter8));
  nand2 gate1788(.a(gate409inter8), .b(gate409inter7), .O(gate409inter9));
  nand2 gate1789(.a(s_177), .b(gate409inter3), .O(gate409inter10));
  nor2  gate1790(.a(gate409inter10), .b(gate409inter9), .O(gate409inter11));
  nor2  gate1791(.a(gate409inter11), .b(gate409inter6), .O(gate409inter12));
  nand2 gate1792(.a(gate409inter12), .b(gate409inter1), .O(G1198));

  xor2  gate981(.a(G1105), .b(G24), .O(gate410inter0));
  nand2 gate982(.a(gate410inter0), .b(s_62), .O(gate410inter1));
  and2  gate983(.a(G1105), .b(G24), .O(gate410inter2));
  inv1  gate984(.a(s_62), .O(gate410inter3));
  inv1  gate985(.a(s_63), .O(gate410inter4));
  nand2 gate986(.a(gate410inter4), .b(gate410inter3), .O(gate410inter5));
  nor2  gate987(.a(gate410inter5), .b(gate410inter2), .O(gate410inter6));
  inv1  gate988(.a(G24), .O(gate410inter7));
  inv1  gate989(.a(G1105), .O(gate410inter8));
  nand2 gate990(.a(gate410inter8), .b(gate410inter7), .O(gate410inter9));
  nand2 gate991(.a(s_63), .b(gate410inter3), .O(gate410inter10));
  nor2  gate992(.a(gate410inter10), .b(gate410inter9), .O(gate410inter11));
  nor2  gate993(.a(gate410inter11), .b(gate410inter6), .O(gate410inter12));
  nand2 gate994(.a(gate410inter12), .b(gate410inter1), .O(G1201));

  xor2  gate1835(.a(G1108), .b(G25), .O(gate411inter0));
  nand2 gate1836(.a(gate411inter0), .b(s_184), .O(gate411inter1));
  and2  gate1837(.a(G1108), .b(G25), .O(gate411inter2));
  inv1  gate1838(.a(s_184), .O(gate411inter3));
  inv1  gate1839(.a(s_185), .O(gate411inter4));
  nand2 gate1840(.a(gate411inter4), .b(gate411inter3), .O(gate411inter5));
  nor2  gate1841(.a(gate411inter5), .b(gate411inter2), .O(gate411inter6));
  inv1  gate1842(.a(G25), .O(gate411inter7));
  inv1  gate1843(.a(G1108), .O(gate411inter8));
  nand2 gate1844(.a(gate411inter8), .b(gate411inter7), .O(gate411inter9));
  nand2 gate1845(.a(s_185), .b(gate411inter3), .O(gate411inter10));
  nor2  gate1846(.a(gate411inter10), .b(gate411inter9), .O(gate411inter11));
  nor2  gate1847(.a(gate411inter11), .b(gate411inter6), .O(gate411inter12));
  nand2 gate1848(.a(gate411inter12), .b(gate411inter1), .O(G1204));
nand2 gate412( .a(G26), .b(G1111), .O(G1207) );
nand2 gate413( .a(G27), .b(G1114), .O(G1210) );
nand2 gate414( .a(G28), .b(G1117), .O(G1213) );
nand2 gate415( .a(G29), .b(G1120), .O(G1216) );
nand2 gate416( .a(G30), .b(G1123), .O(G1219) );

  xor2  gate1457(.a(G1126), .b(G31), .O(gate417inter0));
  nand2 gate1458(.a(gate417inter0), .b(s_130), .O(gate417inter1));
  and2  gate1459(.a(G1126), .b(G31), .O(gate417inter2));
  inv1  gate1460(.a(s_130), .O(gate417inter3));
  inv1  gate1461(.a(s_131), .O(gate417inter4));
  nand2 gate1462(.a(gate417inter4), .b(gate417inter3), .O(gate417inter5));
  nor2  gate1463(.a(gate417inter5), .b(gate417inter2), .O(gate417inter6));
  inv1  gate1464(.a(G31), .O(gate417inter7));
  inv1  gate1465(.a(G1126), .O(gate417inter8));
  nand2 gate1466(.a(gate417inter8), .b(gate417inter7), .O(gate417inter9));
  nand2 gate1467(.a(s_131), .b(gate417inter3), .O(gate417inter10));
  nor2  gate1468(.a(gate417inter10), .b(gate417inter9), .O(gate417inter11));
  nor2  gate1469(.a(gate417inter11), .b(gate417inter6), .O(gate417inter12));
  nand2 gate1470(.a(gate417inter12), .b(gate417inter1), .O(G1222));
nand2 gate418( .a(G32), .b(G1129), .O(G1225) );

  xor2  gate1205(.a(G1132), .b(G1), .O(gate419inter0));
  nand2 gate1206(.a(gate419inter0), .b(s_94), .O(gate419inter1));
  and2  gate1207(.a(G1132), .b(G1), .O(gate419inter2));
  inv1  gate1208(.a(s_94), .O(gate419inter3));
  inv1  gate1209(.a(s_95), .O(gate419inter4));
  nand2 gate1210(.a(gate419inter4), .b(gate419inter3), .O(gate419inter5));
  nor2  gate1211(.a(gate419inter5), .b(gate419inter2), .O(gate419inter6));
  inv1  gate1212(.a(G1), .O(gate419inter7));
  inv1  gate1213(.a(G1132), .O(gate419inter8));
  nand2 gate1214(.a(gate419inter8), .b(gate419inter7), .O(gate419inter9));
  nand2 gate1215(.a(s_95), .b(gate419inter3), .O(gate419inter10));
  nor2  gate1216(.a(gate419inter10), .b(gate419inter9), .O(gate419inter11));
  nor2  gate1217(.a(gate419inter11), .b(gate419inter6), .O(gate419inter12));
  nand2 gate1218(.a(gate419inter12), .b(gate419inter1), .O(G1228));

  xor2  gate2101(.a(G1132), .b(G1036), .O(gate420inter0));
  nand2 gate2102(.a(gate420inter0), .b(s_222), .O(gate420inter1));
  and2  gate2103(.a(G1132), .b(G1036), .O(gate420inter2));
  inv1  gate2104(.a(s_222), .O(gate420inter3));
  inv1  gate2105(.a(s_223), .O(gate420inter4));
  nand2 gate2106(.a(gate420inter4), .b(gate420inter3), .O(gate420inter5));
  nor2  gate2107(.a(gate420inter5), .b(gate420inter2), .O(gate420inter6));
  inv1  gate2108(.a(G1036), .O(gate420inter7));
  inv1  gate2109(.a(G1132), .O(gate420inter8));
  nand2 gate2110(.a(gate420inter8), .b(gate420inter7), .O(gate420inter9));
  nand2 gate2111(.a(s_223), .b(gate420inter3), .O(gate420inter10));
  nor2  gate2112(.a(gate420inter10), .b(gate420inter9), .O(gate420inter11));
  nor2  gate2113(.a(gate420inter11), .b(gate420inter6), .O(gate420inter12));
  nand2 gate2114(.a(gate420inter12), .b(gate420inter1), .O(G1229));
nand2 gate421( .a(G2), .b(G1135), .O(G1230) );
nand2 gate422( .a(G1039), .b(G1135), .O(G1231) );
nand2 gate423( .a(G3), .b(G1138), .O(G1232) );
nand2 gate424( .a(G1042), .b(G1138), .O(G1233) );
nand2 gate425( .a(G4), .b(G1141), .O(G1234) );
nand2 gate426( .a(G1045), .b(G1141), .O(G1235) );
nand2 gate427( .a(G5), .b(G1144), .O(G1236) );
nand2 gate428( .a(G1048), .b(G1144), .O(G1237) );

  xor2  gate715(.a(G1147), .b(G6), .O(gate429inter0));
  nand2 gate716(.a(gate429inter0), .b(s_24), .O(gate429inter1));
  and2  gate717(.a(G1147), .b(G6), .O(gate429inter2));
  inv1  gate718(.a(s_24), .O(gate429inter3));
  inv1  gate719(.a(s_25), .O(gate429inter4));
  nand2 gate720(.a(gate429inter4), .b(gate429inter3), .O(gate429inter5));
  nor2  gate721(.a(gate429inter5), .b(gate429inter2), .O(gate429inter6));
  inv1  gate722(.a(G6), .O(gate429inter7));
  inv1  gate723(.a(G1147), .O(gate429inter8));
  nand2 gate724(.a(gate429inter8), .b(gate429inter7), .O(gate429inter9));
  nand2 gate725(.a(s_25), .b(gate429inter3), .O(gate429inter10));
  nor2  gate726(.a(gate429inter10), .b(gate429inter9), .O(gate429inter11));
  nor2  gate727(.a(gate429inter11), .b(gate429inter6), .O(gate429inter12));
  nand2 gate728(.a(gate429inter12), .b(gate429inter1), .O(G1238));
nand2 gate430( .a(G1051), .b(G1147), .O(G1239) );
nand2 gate431( .a(G7), .b(G1150), .O(G1240) );
nand2 gate432( .a(G1054), .b(G1150), .O(G1241) );
nand2 gate433( .a(G8), .b(G1153), .O(G1242) );

  xor2  gate2549(.a(G1153), .b(G1057), .O(gate434inter0));
  nand2 gate2550(.a(gate434inter0), .b(s_286), .O(gate434inter1));
  and2  gate2551(.a(G1153), .b(G1057), .O(gate434inter2));
  inv1  gate2552(.a(s_286), .O(gate434inter3));
  inv1  gate2553(.a(s_287), .O(gate434inter4));
  nand2 gate2554(.a(gate434inter4), .b(gate434inter3), .O(gate434inter5));
  nor2  gate2555(.a(gate434inter5), .b(gate434inter2), .O(gate434inter6));
  inv1  gate2556(.a(G1057), .O(gate434inter7));
  inv1  gate2557(.a(G1153), .O(gate434inter8));
  nand2 gate2558(.a(gate434inter8), .b(gate434inter7), .O(gate434inter9));
  nand2 gate2559(.a(s_287), .b(gate434inter3), .O(gate434inter10));
  nor2  gate2560(.a(gate434inter10), .b(gate434inter9), .O(gate434inter11));
  nor2  gate2561(.a(gate434inter11), .b(gate434inter6), .O(gate434inter12));
  nand2 gate2562(.a(gate434inter12), .b(gate434inter1), .O(G1243));
nand2 gate435( .a(G9), .b(G1156), .O(G1244) );
nand2 gate436( .a(G1060), .b(G1156), .O(G1245) );
nand2 gate437( .a(G10), .b(G1159), .O(G1246) );
nand2 gate438( .a(G1063), .b(G1159), .O(G1247) );

  xor2  gate1485(.a(G1162), .b(G11), .O(gate439inter0));
  nand2 gate1486(.a(gate439inter0), .b(s_134), .O(gate439inter1));
  and2  gate1487(.a(G1162), .b(G11), .O(gate439inter2));
  inv1  gate1488(.a(s_134), .O(gate439inter3));
  inv1  gate1489(.a(s_135), .O(gate439inter4));
  nand2 gate1490(.a(gate439inter4), .b(gate439inter3), .O(gate439inter5));
  nor2  gate1491(.a(gate439inter5), .b(gate439inter2), .O(gate439inter6));
  inv1  gate1492(.a(G11), .O(gate439inter7));
  inv1  gate1493(.a(G1162), .O(gate439inter8));
  nand2 gate1494(.a(gate439inter8), .b(gate439inter7), .O(gate439inter9));
  nand2 gate1495(.a(s_135), .b(gate439inter3), .O(gate439inter10));
  nor2  gate1496(.a(gate439inter10), .b(gate439inter9), .O(gate439inter11));
  nor2  gate1497(.a(gate439inter11), .b(gate439inter6), .O(gate439inter12));
  nand2 gate1498(.a(gate439inter12), .b(gate439inter1), .O(G1248));
nand2 gate440( .a(G1066), .b(G1162), .O(G1249) );
nand2 gate441( .a(G12), .b(G1165), .O(G1250) );
nand2 gate442( .a(G1069), .b(G1165), .O(G1251) );
nand2 gate443( .a(G13), .b(G1168), .O(G1252) );
nand2 gate444( .a(G1072), .b(G1168), .O(G1253) );
nand2 gate445( .a(G14), .b(G1171), .O(G1254) );
nand2 gate446( .a(G1075), .b(G1171), .O(G1255) );
nand2 gate447( .a(G15), .b(G1174), .O(G1256) );

  xor2  gate1471(.a(G1174), .b(G1078), .O(gate448inter0));
  nand2 gate1472(.a(gate448inter0), .b(s_132), .O(gate448inter1));
  and2  gate1473(.a(G1174), .b(G1078), .O(gate448inter2));
  inv1  gate1474(.a(s_132), .O(gate448inter3));
  inv1  gate1475(.a(s_133), .O(gate448inter4));
  nand2 gate1476(.a(gate448inter4), .b(gate448inter3), .O(gate448inter5));
  nor2  gate1477(.a(gate448inter5), .b(gate448inter2), .O(gate448inter6));
  inv1  gate1478(.a(G1078), .O(gate448inter7));
  inv1  gate1479(.a(G1174), .O(gate448inter8));
  nand2 gate1480(.a(gate448inter8), .b(gate448inter7), .O(gate448inter9));
  nand2 gate1481(.a(s_133), .b(gate448inter3), .O(gate448inter10));
  nor2  gate1482(.a(gate448inter10), .b(gate448inter9), .O(gate448inter11));
  nor2  gate1483(.a(gate448inter11), .b(gate448inter6), .O(gate448inter12));
  nand2 gate1484(.a(gate448inter12), .b(gate448inter1), .O(G1257));

  xor2  gate2255(.a(G1177), .b(G16), .O(gate449inter0));
  nand2 gate2256(.a(gate449inter0), .b(s_244), .O(gate449inter1));
  and2  gate2257(.a(G1177), .b(G16), .O(gate449inter2));
  inv1  gate2258(.a(s_244), .O(gate449inter3));
  inv1  gate2259(.a(s_245), .O(gate449inter4));
  nand2 gate2260(.a(gate449inter4), .b(gate449inter3), .O(gate449inter5));
  nor2  gate2261(.a(gate449inter5), .b(gate449inter2), .O(gate449inter6));
  inv1  gate2262(.a(G16), .O(gate449inter7));
  inv1  gate2263(.a(G1177), .O(gate449inter8));
  nand2 gate2264(.a(gate449inter8), .b(gate449inter7), .O(gate449inter9));
  nand2 gate2265(.a(s_245), .b(gate449inter3), .O(gate449inter10));
  nor2  gate2266(.a(gate449inter10), .b(gate449inter9), .O(gate449inter11));
  nor2  gate2267(.a(gate449inter11), .b(gate449inter6), .O(gate449inter12));
  nand2 gate2268(.a(gate449inter12), .b(gate449inter1), .O(G1258));
nand2 gate450( .a(G1081), .b(G1177), .O(G1259) );
nand2 gate451( .a(G17), .b(G1180), .O(G1260) );
nand2 gate452( .a(G1084), .b(G1180), .O(G1261) );
nand2 gate453( .a(G18), .b(G1183), .O(G1262) );

  xor2  gate2171(.a(G1183), .b(G1087), .O(gate454inter0));
  nand2 gate2172(.a(gate454inter0), .b(s_232), .O(gate454inter1));
  and2  gate2173(.a(G1183), .b(G1087), .O(gate454inter2));
  inv1  gate2174(.a(s_232), .O(gate454inter3));
  inv1  gate2175(.a(s_233), .O(gate454inter4));
  nand2 gate2176(.a(gate454inter4), .b(gate454inter3), .O(gate454inter5));
  nor2  gate2177(.a(gate454inter5), .b(gate454inter2), .O(gate454inter6));
  inv1  gate2178(.a(G1087), .O(gate454inter7));
  inv1  gate2179(.a(G1183), .O(gate454inter8));
  nand2 gate2180(.a(gate454inter8), .b(gate454inter7), .O(gate454inter9));
  nand2 gate2181(.a(s_233), .b(gate454inter3), .O(gate454inter10));
  nor2  gate2182(.a(gate454inter10), .b(gate454inter9), .O(gate454inter11));
  nor2  gate2183(.a(gate454inter11), .b(gate454inter6), .O(gate454inter12));
  nand2 gate2184(.a(gate454inter12), .b(gate454inter1), .O(G1263));
nand2 gate455( .a(G19), .b(G1186), .O(G1264) );

  xor2  gate2395(.a(G1186), .b(G1090), .O(gate456inter0));
  nand2 gate2396(.a(gate456inter0), .b(s_264), .O(gate456inter1));
  and2  gate2397(.a(G1186), .b(G1090), .O(gate456inter2));
  inv1  gate2398(.a(s_264), .O(gate456inter3));
  inv1  gate2399(.a(s_265), .O(gate456inter4));
  nand2 gate2400(.a(gate456inter4), .b(gate456inter3), .O(gate456inter5));
  nor2  gate2401(.a(gate456inter5), .b(gate456inter2), .O(gate456inter6));
  inv1  gate2402(.a(G1090), .O(gate456inter7));
  inv1  gate2403(.a(G1186), .O(gate456inter8));
  nand2 gate2404(.a(gate456inter8), .b(gate456inter7), .O(gate456inter9));
  nand2 gate2405(.a(s_265), .b(gate456inter3), .O(gate456inter10));
  nor2  gate2406(.a(gate456inter10), .b(gate456inter9), .O(gate456inter11));
  nor2  gate2407(.a(gate456inter11), .b(gate456inter6), .O(gate456inter12));
  nand2 gate2408(.a(gate456inter12), .b(gate456inter1), .O(G1265));
nand2 gate457( .a(G20), .b(G1189), .O(G1266) );
nand2 gate458( .a(G1093), .b(G1189), .O(G1267) );
nand2 gate459( .a(G21), .b(G1192), .O(G1268) );
nand2 gate460( .a(G1096), .b(G1192), .O(G1269) );

  xor2  gate1975(.a(G1195), .b(G22), .O(gate461inter0));
  nand2 gate1976(.a(gate461inter0), .b(s_204), .O(gate461inter1));
  and2  gate1977(.a(G1195), .b(G22), .O(gate461inter2));
  inv1  gate1978(.a(s_204), .O(gate461inter3));
  inv1  gate1979(.a(s_205), .O(gate461inter4));
  nand2 gate1980(.a(gate461inter4), .b(gate461inter3), .O(gate461inter5));
  nor2  gate1981(.a(gate461inter5), .b(gate461inter2), .O(gate461inter6));
  inv1  gate1982(.a(G22), .O(gate461inter7));
  inv1  gate1983(.a(G1195), .O(gate461inter8));
  nand2 gate1984(.a(gate461inter8), .b(gate461inter7), .O(gate461inter9));
  nand2 gate1985(.a(s_205), .b(gate461inter3), .O(gate461inter10));
  nor2  gate1986(.a(gate461inter10), .b(gate461inter9), .O(gate461inter11));
  nor2  gate1987(.a(gate461inter11), .b(gate461inter6), .O(gate461inter12));
  nand2 gate1988(.a(gate461inter12), .b(gate461inter1), .O(G1270));

  xor2  gate2437(.a(G1195), .b(G1099), .O(gate462inter0));
  nand2 gate2438(.a(gate462inter0), .b(s_270), .O(gate462inter1));
  and2  gate2439(.a(G1195), .b(G1099), .O(gate462inter2));
  inv1  gate2440(.a(s_270), .O(gate462inter3));
  inv1  gate2441(.a(s_271), .O(gate462inter4));
  nand2 gate2442(.a(gate462inter4), .b(gate462inter3), .O(gate462inter5));
  nor2  gate2443(.a(gate462inter5), .b(gate462inter2), .O(gate462inter6));
  inv1  gate2444(.a(G1099), .O(gate462inter7));
  inv1  gate2445(.a(G1195), .O(gate462inter8));
  nand2 gate2446(.a(gate462inter8), .b(gate462inter7), .O(gate462inter9));
  nand2 gate2447(.a(s_271), .b(gate462inter3), .O(gate462inter10));
  nor2  gate2448(.a(gate462inter10), .b(gate462inter9), .O(gate462inter11));
  nor2  gate2449(.a(gate462inter11), .b(gate462inter6), .O(gate462inter12));
  nand2 gate2450(.a(gate462inter12), .b(gate462inter1), .O(G1271));

  xor2  gate743(.a(G1198), .b(G23), .O(gate463inter0));
  nand2 gate744(.a(gate463inter0), .b(s_28), .O(gate463inter1));
  and2  gate745(.a(G1198), .b(G23), .O(gate463inter2));
  inv1  gate746(.a(s_28), .O(gate463inter3));
  inv1  gate747(.a(s_29), .O(gate463inter4));
  nand2 gate748(.a(gate463inter4), .b(gate463inter3), .O(gate463inter5));
  nor2  gate749(.a(gate463inter5), .b(gate463inter2), .O(gate463inter6));
  inv1  gate750(.a(G23), .O(gate463inter7));
  inv1  gate751(.a(G1198), .O(gate463inter8));
  nand2 gate752(.a(gate463inter8), .b(gate463inter7), .O(gate463inter9));
  nand2 gate753(.a(s_29), .b(gate463inter3), .O(gate463inter10));
  nor2  gate754(.a(gate463inter10), .b(gate463inter9), .O(gate463inter11));
  nor2  gate755(.a(gate463inter11), .b(gate463inter6), .O(gate463inter12));
  nand2 gate756(.a(gate463inter12), .b(gate463inter1), .O(G1272));
nand2 gate464( .a(G1102), .b(G1198), .O(G1273) );
nand2 gate465( .a(G24), .b(G1201), .O(G1274) );

  xor2  gate1751(.a(G1201), .b(G1105), .O(gate466inter0));
  nand2 gate1752(.a(gate466inter0), .b(s_172), .O(gate466inter1));
  and2  gate1753(.a(G1201), .b(G1105), .O(gate466inter2));
  inv1  gate1754(.a(s_172), .O(gate466inter3));
  inv1  gate1755(.a(s_173), .O(gate466inter4));
  nand2 gate1756(.a(gate466inter4), .b(gate466inter3), .O(gate466inter5));
  nor2  gate1757(.a(gate466inter5), .b(gate466inter2), .O(gate466inter6));
  inv1  gate1758(.a(G1105), .O(gate466inter7));
  inv1  gate1759(.a(G1201), .O(gate466inter8));
  nand2 gate1760(.a(gate466inter8), .b(gate466inter7), .O(gate466inter9));
  nand2 gate1761(.a(s_173), .b(gate466inter3), .O(gate466inter10));
  nor2  gate1762(.a(gate466inter10), .b(gate466inter9), .O(gate466inter11));
  nor2  gate1763(.a(gate466inter11), .b(gate466inter6), .O(gate466inter12));
  nand2 gate1764(.a(gate466inter12), .b(gate466inter1), .O(G1275));
nand2 gate467( .a(G25), .b(G1204), .O(G1276) );

  xor2  gate2353(.a(G1204), .b(G1108), .O(gate468inter0));
  nand2 gate2354(.a(gate468inter0), .b(s_258), .O(gate468inter1));
  and2  gate2355(.a(G1204), .b(G1108), .O(gate468inter2));
  inv1  gate2356(.a(s_258), .O(gate468inter3));
  inv1  gate2357(.a(s_259), .O(gate468inter4));
  nand2 gate2358(.a(gate468inter4), .b(gate468inter3), .O(gate468inter5));
  nor2  gate2359(.a(gate468inter5), .b(gate468inter2), .O(gate468inter6));
  inv1  gate2360(.a(G1108), .O(gate468inter7));
  inv1  gate2361(.a(G1204), .O(gate468inter8));
  nand2 gate2362(.a(gate468inter8), .b(gate468inter7), .O(gate468inter9));
  nand2 gate2363(.a(s_259), .b(gate468inter3), .O(gate468inter10));
  nor2  gate2364(.a(gate468inter10), .b(gate468inter9), .O(gate468inter11));
  nor2  gate2365(.a(gate468inter11), .b(gate468inter6), .O(gate468inter12));
  nand2 gate2366(.a(gate468inter12), .b(gate468inter1), .O(G1277));
nand2 gate469( .a(G26), .b(G1207), .O(G1278) );
nand2 gate470( .a(G1111), .b(G1207), .O(G1279) );

  xor2  gate1905(.a(G1210), .b(G27), .O(gate471inter0));
  nand2 gate1906(.a(gate471inter0), .b(s_194), .O(gate471inter1));
  and2  gate1907(.a(G1210), .b(G27), .O(gate471inter2));
  inv1  gate1908(.a(s_194), .O(gate471inter3));
  inv1  gate1909(.a(s_195), .O(gate471inter4));
  nand2 gate1910(.a(gate471inter4), .b(gate471inter3), .O(gate471inter5));
  nor2  gate1911(.a(gate471inter5), .b(gate471inter2), .O(gate471inter6));
  inv1  gate1912(.a(G27), .O(gate471inter7));
  inv1  gate1913(.a(G1210), .O(gate471inter8));
  nand2 gate1914(.a(gate471inter8), .b(gate471inter7), .O(gate471inter9));
  nand2 gate1915(.a(s_195), .b(gate471inter3), .O(gate471inter10));
  nor2  gate1916(.a(gate471inter10), .b(gate471inter9), .O(gate471inter11));
  nor2  gate1917(.a(gate471inter11), .b(gate471inter6), .O(gate471inter12));
  nand2 gate1918(.a(gate471inter12), .b(gate471inter1), .O(G1280));
nand2 gate472( .a(G1114), .b(G1210), .O(G1281) );
nand2 gate473( .a(G28), .b(G1213), .O(G1282) );

  xor2  gate1961(.a(G1213), .b(G1117), .O(gate474inter0));
  nand2 gate1962(.a(gate474inter0), .b(s_202), .O(gate474inter1));
  and2  gate1963(.a(G1213), .b(G1117), .O(gate474inter2));
  inv1  gate1964(.a(s_202), .O(gate474inter3));
  inv1  gate1965(.a(s_203), .O(gate474inter4));
  nand2 gate1966(.a(gate474inter4), .b(gate474inter3), .O(gate474inter5));
  nor2  gate1967(.a(gate474inter5), .b(gate474inter2), .O(gate474inter6));
  inv1  gate1968(.a(G1117), .O(gate474inter7));
  inv1  gate1969(.a(G1213), .O(gate474inter8));
  nand2 gate1970(.a(gate474inter8), .b(gate474inter7), .O(gate474inter9));
  nand2 gate1971(.a(s_203), .b(gate474inter3), .O(gate474inter10));
  nor2  gate1972(.a(gate474inter10), .b(gate474inter9), .O(gate474inter11));
  nor2  gate1973(.a(gate474inter11), .b(gate474inter6), .O(gate474inter12));
  nand2 gate1974(.a(gate474inter12), .b(gate474inter1), .O(G1283));
nand2 gate475( .a(G29), .b(G1216), .O(G1284) );

  xor2  gate1541(.a(G1216), .b(G1120), .O(gate476inter0));
  nand2 gate1542(.a(gate476inter0), .b(s_142), .O(gate476inter1));
  and2  gate1543(.a(G1216), .b(G1120), .O(gate476inter2));
  inv1  gate1544(.a(s_142), .O(gate476inter3));
  inv1  gate1545(.a(s_143), .O(gate476inter4));
  nand2 gate1546(.a(gate476inter4), .b(gate476inter3), .O(gate476inter5));
  nor2  gate1547(.a(gate476inter5), .b(gate476inter2), .O(gate476inter6));
  inv1  gate1548(.a(G1120), .O(gate476inter7));
  inv1  gate1549(.a(G1216), .O(gate476inter8));
  nand2 gate1550(.a(gate476inter8), .b(gate476inter7), .O(gate476inter9));
  nand2 gate1551(.a(s_143), .b(gate476inter3), .O(gate476inter10));
  nor2  gate1552(.a(gate476inter10), .b(gate476inter9), .O(gate476inter11));
  nor2  gate1553(.a(gate476inter11), .b(gate476inter6), .O(gate476inter12));
  nand2 gate1554(.a(gate476inter12), .b(gate476inter1), .O(G1285));
nand2 gate477( .a(G30), .b(G1219), .O(G1286) );
nand2 gate478( .a(G1123), .b(G1219), .O(G1287) );
nand2 gate479( .a(G31), .b(G1222), .O(G1288) );
nand2 gate480( .a(G1126), .b(G1222), .O(G1289) );

  xor2  gate1989(.a(G1225), .b(G32), .O(gate481inter0));
  nand2 gate1990(.a(gate481inter0), .b(s_206), .O(gate481inter1));
  and2  gate1991(.a(G1225), .b(G32), .O(gate481inter2));
  inv1  gate1992(.a(s_206), .O(gate481inter3));
  inv1  gate1993(.a(s_207), .O(gate481inter4));
  nand2 gate1994(.a(gate481inter4), .b(gate481inter3), .O(gate481inter5));
  nor2  gate1995(.a(gate481inter5), .b(gate481inter2), .O(gate481inter6));
  inv1  gate1996(.a(G32), .O(gate481inter7));
  inv1  gate1997(.a(G1225), .O(gate481inter8));
  nand2 gate1998(.a(gate481inter8), .b(gate481inter7), .O(gate481inter9));
  nand2 gate1999(.a(s_207), .b(gate481inter3), .O(gate481inter10));
  nor2  gate2000(.a(gate481inter10), .b(gate481inter9), .O(gate481inter11));
  nor2  gate2001(.a(gate481inter11), .b(gate481inter6), .O(gate481inter12));
  nand2 gate2002(.a(gate481inter12), .b(gate481inter1), .O(G1290));

  xor2  gate1821(.a(G1225), .b(G1129), .O(gate482inter0));
  nand2 gate1822(.a(gate482inter0), .b(s_182), .O(gate482inter1));
  and2  gate1823(.a(G1225), .b(G1129), .O(gate482inter2));
  inv1  gate1824(.a(s_182), .O(gate482inter3));
  inv1  gate1825(.a(s_183), .O(gate482inter4));
  nand2 gate1826(.a(gate482inter4), .b(gate482inter3), .O(gate482inter5));
  nor2  gate1827(.a(gate482inter5), .b(gate482inter2), .O(gate482inter6));
  inv1  gate1828(.a(G1129), .O(gate482inter7));
  inv1  gate1829(.a(G1225), .O(gate482inter8));
  nand2 gate1830(.a(gate482inter8), .b(gate482inter7), .O(gate482inter9));
  nand2 gate1831(.a(s_183), .b(gate482inter3), .O(gate482inter10));
  nor2  gate1832(.a(gate482inter10), .b(gate482inter9), .O(gate482inter11));
  nor2  gate1833(.a(gate482inter11), .b(gate482inter6), .O(gate482inter12));
  nand2 gate1834(.a(gate482inter12), .b(gate482inter1), .O(G1291));
nand2 gate483( .a(G1228), .b(G1229), .O(G1292) );
nand2 gate484( .a(G1230), .b(G1231), .O(G1293) );
nand2 gate485( .a(G1232), .b(G1233), .O(G1294) );

  xor2  gate1933(.a(G1235), .b(G1234), .O(gate486inter0));
  nand2 gate1934(.a(gate486inter0), .b(s_198), .O(gate486inter1));
  and2  gate1935(.a(G1235), .b(G1234), .O(gate486inter2));
  inv1  gate1936(.a(s_198), .O(gate486inter3));
  inv1  gate1937(.a(s_199), .O(gate486inter4));
  nand2 gate1938(.a(gate486inter4), .b(gate486inter3), .O(gate486inter5));
  nor2  gate1939(.a(gate486inter5), .b(gate486inter2), .O(gate486inter6));
  inv1  gate1940(.a(G1234), .O(gate486inter7));
  inv1  gate1941(.a(G1235), .O(gate486inter8));
  nand2 gate1942(.a(gate486inter8), .b(gate486inter7), .O(gate486inter9));
  nand2 gate1943(.a(s_199), .b(gate486inter3), .O(gate486inter10));
  nor2  gate1944(.a(gate486inter10), .b(gate486inter9), .O(gate486inter11));
  nor2  gate1945(.a(gate486inter11), .b(gate486inter6), .O(gate486inter12));
  nand2 gate1946(.a(gate486inter12), .b(gate486inter1), .O(G1295));

  xor2  gate1695(.a(G1237), .b(G1236), .O(gate487inter0));
  nand2 gate1696(.a(gate487inter0), .b(s_164), .O(gate487inter1));
  and2  gate1697(.a(G1237), .b(G1236), .O(gate487inter2));
  inv1  gate1698(.a(s_164), .O(gate487inter3));
  inv1  gate1699(.a(s_165), .O(gate487inter4));
  nand2 gate1700(.a(gate487inter4), .b(gate487inter3), .O(gate487inter5));
  nor2  gate1701(.a(gate487inter5), .b(gate487inter2), .O(gate487inter6));
  inv1  gate1702(.a(G1236), .O(gate487inter7));
  inv1  gate1703(.a(G1237), .O(gate487inter8));
  nand2 gate1704(.a(gate487inter8), .b(gate487inter7), .O(gate487inter9));
  nand2 gate1705(.a(s_165), .b(gate487inter3), .O(gate487inter10));
  nor2  gate1706(.a(gate487inter10), .b(gate487inter9), .O(gate487inter11));
  nor2  gate1707(.a(gate487inter11), .b(gate487inter6), .O(gate487inter12));
  nand2 gate1708(.a(gate487inter12), .b(gate487inter1), .O(G1296));

  xor2  gate2521(.a(G1239), .b(G1238), .O(gate488inter0));
  nand2 gate2522(.a(gate488inter0), .b(s_282), .O(gate488inter1));
  and2  gate2523(.a(G1239), .b(G1238), .O(gate488inter2));
  inv1  gate2524(.a(s_282), .O(gate488inter3));
  inv1  gate2525(.a(s_283), .O(gate488inter4));
  nand2 gate2526(.a(gate488inter4), .b(gate488inter3), .O(gate488inter5));
  nor2  gate2527(.a(gate488inter5), .b(gate488inter2), .O(gate488inter6));
  inv1  gate2528(.a(G1238), .O(gate488inter7));
  inv1  gate2529(.a(G1239), .O(gate488inter8));
  nand2 gate2530(.a(gate488inter8), .b(gate488inter7), .O(gate488inter9));
  nand2 gate2531(.a(s_283), .b(gate488inter3), .O(gate488inter10));
  nor2  gate2532(.a(gate488inter10), .b(gate488inter9), .O(gate488inter11));
  nor2  gate2533(.a(gate488inter11), .b(gate488inter6), .O(gate488inter12));
  nand2 gate2534(.a(gate488inter12), .b(gate488inter1), .O(G1297));
nand2 gate489( .a(G1240), .b(G1241), .O(G1298) );
nand2 gate490( .a(G1242), .b(G1243), .O(G1299) );
nand2 gate491( .a(G1244), .b(G1245), .O(G1300) );

  xor2  gate659(.a(G1247), .b(G1246), .O(gate492inter0));
  nand2 gate660(.a(gate492inter0), .b(s_16), .O(gate492inter1));
  and2  gate661(.a(G1247), .b(G1246), .O(gate492inter2));
  inv1  gate662(.a(s_16), .O(gate492inter3));
  inv1  gate663(.a(s_17), .O(gate492inter4));
  nand2 gate664(.a(gate492inter4), .b(gate492inter3), .O(gate492inter5));
  nor2  gate665(.a(gate492inter5), .b(gate492inter2), .O(gate492inter6));
  inv1  gate666(.a(G1246), .O(gate492inter7));
  inv1  gate667(.a(G1247), .O(gate492inter8));
  nand2 gate668(.a(gate492inter8), .b(gate492inter7), .O(gate492inter9));
  nand2 gate669(.a(s_17), .b(gate492inter3), .O(gate492inter10));
  nor2  gate670(.a(gate492inter10), .b(gate492inter9), .O(gate492inter11));
  nor2  gate671(.a(gate492inter11), .b(gate492inter6), .O(gate492inter12));
  nand2 gate672(.a(gate492inter12), .b(gate492inter1), .O(G1301));
nand2 gate493( .a(G1248), .b(G1249), .O(G1302) );

  xor2  gate1247(.a(G1251), .b(G1250), .O(gate494inter0));
  nand2 gate1248(.a(gate494inter0), .b(s_100), .O(gate494inter1));
  and2  gate1249(.a(G1251), .b(G1250), .O(gate494inter2));
  inv1  gate1250(.a(s_100), .O(gate494inter3));
  inv1  gate1251(.a(s_101), .O(gate494inter4));
  nand2 gate1252(.a(gate494inter4), .b(gate494inter3), .O(gate494inter5));
  nor2  gate1253(.a(gate494inter5), .b(gate494inter2), .O(gate494inter6));
  inv1  gate1254(.a(G1250), .O(gate494inter7));
  inv1  gate1255(.a(G1251), .O(gate494inter8));
  nand2 gate1256(.a(gate494inter8), .b(gate494inter7), .O(gate494inter9));
  nand2 gate1257(.a(s_101), .b(gate494inter3), .O(gate494inter10));
  nor2  gate1258(.a(gate494inter10), .b(gate494inter9), .O(gate494inter11));
  nor2  gate1259(.a(gate494inter11), .b(gate494inter6), .O(gate494inter12));
  nand2 gate1260(.a(gate494inter12), .b(gate494inter1), .O(G1303));

  xor2  gate687(.a(G1253), .b(G1252), .O(gate495inter0));
  nand2 gate688(.a(gate495inter0), .b(s_20), .O(gate495inter1));
  and2  gate689(.a(G1253), .b(G1252), .O(gate495inter2));
  inv1  gate690(.a(s_20), .O(gate495inter3));
  inv1  gate691(.a(s_21), .O(gate495inter4));
  nand2 gate692(.a(gate495inter4), .b(gate495inter3), .O(gate495inter5));
  nor2  gate693(.a(gate495inter5), .b(gate495inter2), .O(gate495inter6));
  inv1  gate694(.a(G1252), .O(gate495inter7));
  inv1  gate695(.a(G1253), .O(gate495inter8));
  nand2 gate696(.a(gate495inter8), .b(gate495inter7), .O(gate495inter9));
  nand2 gate697(.a(s_21), .b(gate495inter3), .O(gate495inter10));
  nor2  gate698(.a(gate495inter10), .b(gate495inter9), .O(gate495inter11));
  nor2  gate699(.a(gate495inter11), .b(gate495inter6), .O(gate495inter12));
  nand2 gate700(.a(gate495inter12), .b(gate495inter1), .O(G1304));
nand2 gate496( .a(G1254), .b(G1255), .O(G1305) );

  xor2  gate1681(.a(G1257), .b(G1256), .O(gate497inter0));
  nand2 gate1682(.a(gate497inter0), .b(s_162), .O(gate497inter1));
  and2  gate1683(.a(G1257), .b(G1256), .O(gate497inter2));
  inv1  gate1684(.a(s_162), .O(gate497inter3));
  inv1  gate1685(.a(s_163), .O(gate497inter4));
  nand2 gate1686(.a(gate497inter4), .b(gate497inter3), .O(gate497inter5));
  nor2  gate1687(.a(gate497inter5), .b(gate497inter2), .O(gate497inter6));
  inv1  gate1688(.a(G1256), .O(gate497inter7));
  inv1  gate1689(.a(G1257), .O(gate497inter8));
  nand2 gate1690(.a(gate497inter8), .b(gate497inter7), .O(gate497inter9));
  nand2 gate1691(.a(s_163), .b(gate497inter3), .O(gate497inter10));
  nor2  gate1692(.a(gate497inter10), .b(gate497inter9), .O(gate497inter11));
  nor2  gate1693(.a(gate497inter11), .b(gate497inter6), .O(gate497inter12));
  nand2 gate1694(.a(gate497inter12), .b(gate497inter1), .O(G1306));
nand2 gate498( .a(G1258), .b(G1259), .O(G1307) );

  xor2  gate855(.a(G1261), .b(G1260), .O(gate499inter0));
  nand2 gate856(.a(gate499inter0), .b(s_44), .O(gate499inter1));
  and2  gate857(.a(G1261), .b(G1260), .O(gate499inter2));
  inv1  gate858(.a(s_44), .O(gate499inter3));
  inv1  gate859(.a(s_45), .O(gate499inter4));
  nand2 gate860(.a(gate499inter4), .b(gate499inter3), .O(gate499inter5));
  nor2  gate861(.a(gate499inter5), .b(gate499inter2), .O(gate499inter6));
  inv1  gate862(.a(G1260), .O(gate499inter7));
  inv1  gate863(.a(G1261), .O(gate499inter8));
  nand2 gate864(.a(gate499inter8), .b(gate499inter7), .O(gate499inter9));
  nand2 gate865(.a(s_45), .b(gate499inter3), .O(gate499inter10));
  nor2  gate866(.a(gate499inter10), .b(gate499inter9), .O(gate499inter11));
  nor2  gate867(.a(gate499inter11), .b(gate499inter6), .O(gate499inter12));
  nand2 gate868(.a(gate499inter12), .b(gate499inter1), .O(G1308));
nand2 gate500( .a(G1262), .b(G1263), .O(G1309) );
nand2 gate501( .a(G1264), .b(G1265), .O(G1310) );

  xor2  gate2199(.a(G1267), .b(G1266), .O(gate502inter0));
  nand2 gate2200(.a(gate502inter0), .b(s_236), .O(gate502inter1));
  and2  gate2201(.a(G1267), .b(G1266), .O(gate502inter2));
  inv1  gate2202(.a(s_236), .O(gate502inter3));
  inv1  gate2203(.a(s_237), .O(gate502inter4));
  nand2 gate2204(.a(gate502inter4), .b(gate502inter3), .O(gate502inter5));
  nor2  gate2205(.a(gate502inter5), .b(gate502inter2), .O(gate502inter6));
  inv1  gate2206(.a(G1266), .O(gate502inter7));
  inv1  gate2207(.a(G1267), .O(gate502inter8));
  nand2 gate2208(.a(gate502inter8), .b(gate502inter7), .O(gate502inter9));
  nand2 gate2209(.a(s_237), .b(gate502inter3), .O(gate502inter10));
  nor2  gate2210(.a(gate502inter10), .b(gate502inter9), .O(gate502inter11));
  nor2  gate2211(.a(gate502inter11), .b(gate502inter6), .O(gate502inter12));
  nand2 gate2212(.a(gate502inter12), .b(gate502inter1), .O(G1311));
nand2 gate503( .a(G1268), .b(G1269), .O(G1312) );

  xor2  gate827(.a(G1271), .b(G1270), .O(gate504inter0));
  nand2 gate828(.a(gate504inter0), .b(s_40), .O(gate504inter1));
  and2  gate829(.a(G1271), .b(G1270), .O(gate504inter2));
  inv1  gate830(.a(s_40), .O(gate504inter3));
  inv1  gate831(.a(s_41), .O(gate504inter4));
  nand2 gate832(.a(gate504inter4), .b(gate504inter3), .O(gate504inter5));
  nor2  gate833(.a(gate504inter5), .b(gate504inter2), .O(gate504inter6));
  inv1  gate834(.a(G1270), .O(gate504inter7));
  inv1  gate835(.a(G1271), .O(gate504inter8));
  nand2 gate836(.a(gate504inter8), .b(gate504inter7), .O(gate504inter9));
  nand2 gate837(.a(s_41), .b(gate504inter3), .O(gate504inter10));
  nor2  gate838(.a(gate504inter10), .b(gate504inter9), .O(gate504inter11));
  nor2  gate839(.a(gate504inter11), .b(gate504inter6), .O(gate504inter12));
  nand2 gate840(.a(gate504inter12), .b(gate504inter1), .O(G1313));
nand2 gate505( .a(G1272), .b(G1273), .O(G1314) );
nand2 gate506( .a(G1274), .b(G1275), .O(G1315) );

  xor2  gate1793(.a(G1277), .b(G1276), .O(gate507inter0));
  nand2 gate1794(.a(gate507inter0), .b(s_178), .O(gate507inter1));
  and2  gate1795(.a(G1277), .b(G1276), .O(gate507inter2));
  inv1  gate1796(.a(s_178), .O(gate507inter3));
  inv1  gate1797(.a(s_179), .O(gate507inter4));
  nand2 gate1798(.a(gate507inter4), .b(gate507inter3), .O(gate507inter5));
  nor2  gate1799(.a(gate507inter5), .b(gate507inter2), .O(gate507inter6));
  inv1  gate1800(.a(G1276), .O(gate507inter7));
  inv1  gate1801(.a(G1277), .O(gate507inter8));
  nand2 gate1802(.a(gate507inter8), .b(gate507inter7), .O(gate507inter9));
  nand2 gate1803(.a(s_179), .b(gate507inter3), .O(gate507inter10));
  nor2  gate1804(.a(gate507inter10), .b(gate507inter9), .O(gate507inter11));
  nor2  gate1805(.a(gate507inter11), .b(gate507inter6), .O(gate507inter12));
  nand2 gate1806(.a(gate507inter12), .b(gate507inter1), .O(G1316));
nand2 gate508( .a(G1278), .b(G1279), .O(G1317) );

  xor2  gate1275(.a(G1281), .b(G1280), .O(gate509inter0));
  nand2 gate1276(.a(gate509inter0), .b(s_104), .O(gate509inter1));
  and2  gate1277(.a(G1281), .b(G1280), .O(gate509inter2));
  inv1  gate1278(.a(s_104), .O(gate509inter3));
  inv1  gate1279(.a(s_105), .O(gate509inter4));
  nand2 gate1280(.a(gate509inter4), .b(gate509inter3), .O(gate509inter5));
  nor2  gate1281(.a(gate509inter5), .b(gate509inter2), .O(gate509inter6));
  inv1  gate1282(.a(G1280), .O(gate509inter7));
  inv1  gate1283(.a(G1281), .O(gate509inter8));
  nand2 gate1284(.a(gate509inter8), .b(gate509inter7), .O(gate509inter9));
  nand2 gate1285(.a(s_105), .b(gate509inter3), .O(gate509inter10));
  nor2  gate1286(.a(gate509inter10), .b(gate509inter9), .O(gate509inter11));
  nor2  gate1287(.a(gate509inter11), .b(gate509inter6), .O(gate509inter12));
  nand2 gate1288(.a(gate509inter12), .b(gate509inter1), .O(G1318));
nand2 gate510( .a(G1282), .b(G1283), .O(G1319) );
nand2 gate511( .a(G1284), .b(G1285), .O(G1320) );
nand2 gate512( .a(G1286), .b(G1287), .O(G1321) );

  xor2  gate1303(.a(G1289), .b(G1288), .O(gate513inter0));
  nand2 gate1304(.a(gate513inter0), .b(s_108), .O(gate513inter1));
  and2  gate1305(.a(G1289), .b(G1288), .O(gate513inter2));
  inv1  gate1306(.a(s_108), .O(gate513inter3));
  inv1  gate1307(.a(s_109), .O(gate513inter4));
  nand2 gate1308(.a(gate513inter4), .b(gate513inter3), .O(gate513inter5));
  nor2  gate1309(.a(gate513inter5), .b(gate513inter2), .O(gate513inter6));
  inv1  gate1310(.a(G1288), .O(gate513inter7));
  inv1  gate1311(.a(G1289), .O(gate513inter8));
  nand2 gate1312(.a(gate513inter8), .b(gate513inter7), .O(gate513inter9));
  nand2 gate1313(.a(s_109), .b(gate513inter3), .O(gate513inter10));
  nor2  gate1314(.a(gate513inter10), .b(gate513inter9), .O(gate513inter11));
  nor2  gate1315(.a(gate513inter11), .b(gate513inter6), .O(gate513inter12));
  nand2 gate1316(.a(gate513inter12), .b(gate513inter1), .O(G1322));

  xor2  gate2535(.a(G1291), .b(G1290), .O(gate514inter0));
  nand2 gate2536(.a(gate514inter0), .b(s_284), .O(gate514inter1));
  and2  gate2537(.a(G1291), .b(G1290), .O(gate514inter2));
  inv1  gate2538(.a(s_284), .O(gate514inter3));
  inv1  gate2539(.a(s_285), .O(gate514inter4));
  nand2 gate2540(.a(gate514inter4), .b(gate514inter3), .O(gate514inter5));
  nor2  gate2541(.a(gate514inter5), .b(gate514inter2), .O(gate514inter6));
  inv1  gate2542(.a(G1290), .O(gate514inter7));
  inv1  gate2543(.a(G1291), .O(gate514inter8));
  nand2 gate2544(.a(gate514inter8), .b(gate514inter7), .O(gate514inter9));
  nand2 gate2545(.a(s_285), .b(gate514inter3), .O(gate514inter10));
  nor2  gate2546(.a(gate514inter10), .b(gate514inter9), .O(gate514inter11));
  nor2  gate2547(.a(gate514inter11), .b(gate514inter6), .O(gate514inter12));
  nand2 gate2548(.a(gate514inter12), .b(gate514inter1), .O(G1323));
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule