module c432 (N1,N4,N8,N11,N14,N17,N21,N24,N27,N30,
             N34,N37,N40,N43,N47,N50,N53,N56,N60,N63,
             N66,N69,N73,N76,N79,N82,N86,N89,N92,N95,
             N99,N102,N105,N108,N112,N115,N223,N329,N370,N421,
             N430,N431,N432);

input N1,N4,N8,N11,N14,N17,N21,N24,N27,N30,
      N34,N37,N40,N43,N47,N50,N53,N56,N60,N63,
      N66,N69,N73,N76,N79,N82,N86,N89,N92,N95,
      N99,N102,N105,N108,N112,N115;//RE__PI;

input s_0,s_1;//RE__ALLOW(00,01,10,11);
input s_2,s_3;//RE__ALLOW(00,01,10,11);
input s_4,s_5;//RE__ALLOW(00,01,10,11);
input s_6,s_7;//RE__ALLOW(00,01,10,11);
input s_8,s_9;//RE__ALLOW(00,01,10,11);
input s_10,s_11;//RE__ALLOW(00,01,10,11);
input s_12,s_13;//RE__ALLOW(00,01,10,11);
input s_14,s_15;//RE__ALLOW(00,01,10,11);
input s_16,s_17;//RE__ALLOW(00,01,10,11);
input s_18,s_19;//RE__ALLOW(00,01,10,11);
input s_20,s_21;//RE__ALLOW(00,01,10,11);
input s_22,s_23;//RE__ALLOW(00,01,10,11);
input s_24,s_25;//RE__ALLOW(00,01,10,11);
input s_26,s_27;//RE__ALLOW(00,01,10,11);
input s_28,s_29;//RE__ALLOW(00,01,10,11);
input s_30,s_31;//RE__ALLOW(00,01,10,11);
input s_32,s_33;//RE__ALLOW(00,01,10,11);
input s_34,s_35;//RE__ALLOW(00,01,10,11);
input s_36,s_37;//RE__ALLOW(00,01,10,11);
input s_38,s_39;//RE__ALLOW(00,01,10,11);
input s_40,s_41;//RE__ALLOW(00,01,10,11);
input s_42,s_43;//RE__ALLOW(00,01,10,11);
input s_44,s_45;//RE__ALLOW(00,01,10,11);
input s_46,s_47;//RE__ALLOW(00,01,10,11);
input s_48,s_49;//RE__ALLOW(00,01,10,11);
input s_50,s_51;//RE__ALLOW(00,01,10,11);
input s_52,s_53;//RE__ALLOW(00,01,10,11);
input s_54,s_55;//RE__ALLOW(00,01,10,11);
input s_56,s_57;//RE__ALLOW(00,01,10,11);
input s_58,s_59;//RE__ALLOW(00,01,10,11);
input s_60,s_61;//RE__ALLOW(00,01,10,11);
output N223,N329,N370,N421,N430,N431,N432;

wire N118,N119,N122,N123,N126,N127,N130,N131,N134,N135,
     N138,N139,N142,N143,N146,N147,N150,N151,N154,N157,
     N158,N159,N162,N165,N168,N171,N174,N177,N180,N183,
     N184,N185,N186,N187,N188,N189,N190,N191,N192,N193,
     N194,N195,N196,N197,N198,N199,N203,N213,N224,N227,
     N230,N233,N236,N239,N242,N243,N246,N247,N250,N251,
     N254,N255,N256,N257,N258,N259,N260,N263,N264,N267,
     N270,N273,N276,N279,N282,N285,N288,N289,N290,N291,
     N292,N293,N294,N295,N296,N300,N301,N302,N303,N304,
     N305,N306,N307,N308,N309,N319,N330,N331,N332,N333,
     N334,N335,N336,N337,N338,N339,N340,N341,N342,N343,
     N344,N345,N346,N347,N348,N349,N350,N351,N352,N353,
     N354,N355,N356,N357,N360,N371,N372,N373,N374,N375,
     N376,N377,N378,N379,N380,N381,N386,N393,N399,N404,
     N407,N411,N414,N415,N416,N417,N418,N419,N420,N422,
     N425,N428,N429, gate23inter0, gate23inter1, gate23inter2, gate23inter3, gate23inter4, gate23inter5, gate23inter6, gate23inter7, gate23inter8, gate23inter9, gate23inter10, gate23inter11, gate23inter12, gate83inter0, gate83inter1, gate83inter2, gate83inter3, gate83inter4, gate83inter5, gate83inter6, gate83inter7, gate83inter8, gate83inter9, gate83inter10, gate83inter11, gate83inter12, gate124inter0, gate124inter1, gate124inter2, gate124inter3, gate124inter4, gate124inter5, gate124inter6, gate124inter7, gate124inter8, gate124inter9, gate124inter10, gate124inter11, gate124inter12, gate57inter0, gate57inter1, gate57inter2, gate57inter3, gate57inter4, gate57inter5, gate57inter6, gate57inter7, gate57inter8, gate57inter9, gate57inter10, gate57inter11, gate57inter12, gate123inter0, gate123inter1, gate123inter2, gate123inter3, gate123inter4, gate123inter5, gate123inter6, gate123inter7, gate123inter8, gate123inter9, gate123inter10, gate123inter11, gate123inter12, gate43inter0, gate43inter1, gate43inter2, gate43inter3, gate43inter4, gate43inter5, gate43inter6, gate43inter7, gate43inter8, gate43inter9, gate43inter10, gate43inter11, gate43inter12, gate74inter0, gate74inter1, gate74inter2, gate74inter3, gate74inter4, gate74inter5, gate74inter6, gate74inter7, gate74inter8, gate74inter9, gate74inter10, gate74inter11, gate74inter12, gate69inter0, gate69inter1, gate69inter2, gate69inter3, gate69inter4, gate69inter5, gate69inter6, gate69inter7, gate69inter8, gate69inter9, gate69inter10, gate69inter11, gate69inter12, gate78inter0, gate78inter1, gate78inter2, gate78inter3, gate78inter4, gate78inter5, gate78inter6, gate78inter7, gate78inter8, gate78inter9, gate78inter10, gate78inter11, gate78inter12, gate34inter0, gate34inter1, gate34inter2, gate34inter3, gate34inter4, gate34inter5, gate34inter6, gate34inter7, gate34inter8, gate34inter9, gate34inter10, gate34inter11, gate34inter12, gate136inter0, gate136inter1, gate136inter2, gate136inter3, gate136inter4, gate136inter5, gate136inter6, gate136inter7, gate136inter8, gate136inter9, gate136inter10, gate136inter11, gate136inter12, gate117inter0, gate117inter1, gate117inter2, gate117inter3, gate117inter4, gate117inter5, gate117inter6, gate117inter7, gate117inter8, gate117inter9, gate117inter10, gate117inter11, gate117inter12, gate102inter0, gate102inter1, gate102inter2, gate102inter3, gate102inter4, gate102inter5, gate102inter6, gate102inter7, gate102inter8, gate102inter9, gate102inter10, gate102inter11, gate102inter12, gate132inter0, gate132inter1, gate132inter2, gate132inter3, gate132inter4, gate132inter5, gate132inter6, gate132inter7, gate132inter8, gate132inter9, gate132inter10, gate132inter11, gate132inter12, gate80inter0, gate80inter1, gate80inter2, gate80inter3, gate80inter4, gate80inter5, gate80inter6, gate80inter7, gate80inter8, gate80inter9, gate80inter10, gate80inter11, gate80inter12, gate116inter0, gate116inter1, gate116inter2, gate116inter3, gate116inter4, gate116inter5, gate116inter6, gate116inter7, gate116inter8, gate116inter9, gate116inter10, gate116inter11, gate116inter12, gate41inter0, gate41inter1, gate41inter2, gate41inter3, gate41inter4, gate41inter5, gate41inter6, gate41inter7, gate41inter8, gate41inter9, gate41inter10, gate41inter11, gate41inter12, gate53inter0, gate53inter1, gate53inter2, gate53inter3, gate53inter4, gate53inter5, gate53inter6, gate53inter7, gate53inter8, gate53inter9, gate53inter10, gate53inter11, gate53inter12, gate55inter0, gate55inter1, gate55inter2, gate55inter3, gate55inter4, gate55inter5, gate55inter6, gate55inter7, gate55inter8, gate55inter9, gate55inter10, gate55inter11, gate55inter12, gate64inter0, gate64inter1, gate64inter2, gate64inter3, gate64inter4, gate64inter5, gate64inter6, gate64inter7, gate64inter8, gate64inter9, gate64inter10, gate64inter11, gate64inter12, gate109inter0, gate109inter1, gate109inter2, gate109inter3, gate109inter4, gate109inter5, gate109inter6, gate109inter7, gate109inter8, gate109inter9, gate109inter10, gate109inter11, gate109inter12, gate111inter0, gate111inter1, gate111inter2, gate111inter3, gate111inter4, gate111inter5, gate111inter6, gate111inter7, gate111inter8, gate111inter9, gate111inter10, gate111inter11, gate111inter12, gate82inter0, gate82inter1, gate82inter2, gate82inter3, gate82inter4, gate82inter5, gate82inter6, gate82inter7, gate82inter8, gate82inter9, gate82inter10, gate82inter11, gate82inter12, gate107inter0, gate107inter1, gate107inter2, gate107inter3, gate107inter4, gate107inter5, gate107inter6, gate107inter7, gate107inter8, gate107inter9, gate107inter10, gate107inter11, gate107inter12, gate32inter0, gate32inter1, gate32inter2, gate32inter3, gate32inter4, gate32inter5, gate32inter6, gate32inter7, gate32inter8, gate32inter9, gate32inter10, gate32inter11, gate32inter12, gate72inter0, gate72inter1, gate72inter2, gate72inter3, gate72inter4, gate72inter5, gate72inter6, gate72inter7, gate72inter8, gate72inter9, gate72inter10, gate72inter11, gate72inter12, gate62inter0, gate62inter1, gate62inter2, gate62inter3, gate62inter4, gate62inter5, gate62inter6, gate62inter7, gate62inter8, gate62inter9, gate62inter10, gate62inter11, gate62inter12, gate76inter0, gate76inter1, gate76inter2, gate76inter3, gate76inter4, gate76inter5, gate76inter6, gate76inter7, gate76inter8, gate76inter9, gate76inter10, gate76inter11, gate76inter12, gate61inter0, gate61inter1, gate61inter2, gate61inter3, gate61inter4, gate61inter5, gate61inter6, gate61inter7, gate61inter8, gate61inter9, gate61inter10, gate61inter11, gate61inter12, gate119inter0, gate119inter1, gate119inter2, gate119inter3, gate119inter4, gate119inter5, gate119inter6, gate119inter7, gate119inter8, gate119inter9, gate119inter10, gate119inter11, gate119inter12, gate73inter0, gate73inter1, gate73inter2, gate73inter3, gate73inter4, gate73inter5, gate73inter6, gate73inter7, gate73inter8, gate73inter9, gate73inter10, gate73inter11, gate73inter12;



inv1 gate1( .a(N1), .O(N118) );
inv1 gate2( .a(N4), .O(N119) );
inv1 gate3( .a(N11), .O(N122) );
inv1 gate4( .a(N17), .O(N123) );
inv1 gate5( .a(N24), .O(N126) );
inv1 gate6( .a(N30), .O(N127) );
inv1 gate7( .a(N37), .O(N130) );
inv1 gate8( .a(N43), .O(N131) );
inv1 gate9( .a(N50), .O(N134) );
inv1 gate10( .a(N56), .O(N135) );
inv1 gate11( .a(N63), .O(N138) );
inv1 gate12( .a(N69), .O(N139) );
inv1 gate13( .a(N76), .O(N142) );
inv1 gate14( .a(N82), .O(N143) );
inv1 gate15( .a(N89), .O(N146) );
inv1 gate16( .a(N95), .O(N147) );
inv1 gate17( .a(N102), .O(N150) );
inv1 gate18( .a(N108), .O(N151) );
nand2 gate19( .a(N118), .b(N4), .O(N154) );
nor2 gate20( .a(N8), .b(N119), .O(N157) );
nor2 gate21( .a(N14), .b(N119), .O(N158) );
nand2 gate22( .a(N122), .b(N17), .O(N159) );

  xor2  gate161(.a(N30), .b(N126), .O(gate23inter0));
  nand2 gate162(.a(gate23inter0), .b(s_0), .O(gate23inter1));
  and2  gate163(.a(N30), .b(N126), .O(gate23inter2));
  inv1  gate164(.a(s_0), .O(gate23inter3));
  inv1  gate165(.a(s_1), .O(gate23inter4));
  nand2 gate166(.a(gate23inter4), .b(gate23inter3), .O(gate23inter5));
  nor2  gate167(.a(gate23inter5), .b(gate23inter2), .O(gate23inter6));
  inv1  gate168(.a(N126), .O(gate23inter7));
  inv1  gate169(.a(N30), .O(gate23inter8));
  nand2 gate170(.a(gate23inter8), .b(gate23inter7), .O(gate23inter9));
  nand2 gate171(.a(s_1), .b(gate23inter3), .O(gate23inter10));
  nor2  gate172(.a(gate23inter10), .b(gate23inter9), .O(gate23inter11));
  nor2  gate173(.a(gate23inter11), .b(gate23inter6), .O(gate23inter12));
  nand2 gate174(.a(gate23inter12), .b(gate23inter1), .O(N162));
nand2 gate24( .a(N130), .b(N43), .O(N165) );
nand2 gate25( .a(N134), .b(N56), .O(N168) );
nand2 gate26( .a(N138), .b(N69), .O(N171) );
nand2 gate27( .a(N142), .b(N82), .O(N174) );
nand2 gate28( .a(N146), .b(N95), .O(N177) );
nand2 gate29( .a(N150), .b(N108), .O(N180) );
nor2 gate30( .a(N21), .b(N123), .O(N183) );
nor2 gate31( .a(N27), .b(N123), .O(N184) );

  xor2  gate497(.a(N127), .b(N34), .O(gate32inter0));
  nand2 gate498(.a(gate32inter0), .b(s_48), .O(gate32inter1));
  and2  gate499(.a(N127), .b(N34), .O(gate32inter2));
  inv1  gate500(.a(s_48), .O(gate32inter3));
  inv1  gate501(.a(s_49), .O(gate32inter4));
  nand2 gate502(.a(gate32inter4), .b(gate32inter3), .O(gate32inter5));
  nor2  gate503(.a(gate32inter5), .b(gate32inter2), .O(gate32inter6));
  inv1  gate504(.a(N34), .O(gate32inter7));
  inv1  gate505(.a(N127), .O(gate32inter8));
  nand2 gate506(.a(gate32inter8), .b(gate32inter7), .O(gate32inter9));
  nand2 gate507(.a(s_49), .b(gate32inter3), .O(gate32inter10));
  nor2  gate508(.a(gate32inter10), .b(gate32inter9), .O(gate32inter11));
  nor2  gate509(.a(gate32inter11), .b(gate32inter6), .O(gate32inter12));
  nand2 gate510(.a(gate32inter12), .b(gate32inter1), .O(N185));
nor2 gate33( .a(N40), .b(N127), .O(N186) );

  xor2  gate287(.a(N131), .b(N47), .O(gate34inter0));
  nand2 gate288(.a(gate34inter0), .b(s_18), .O(gate34inter1));
  and2  gate289(.a(N131), .b(N47), .O(gate34inter2));
  inv1  gate290(.a(s_18), .O(gate34inter3));
  inv1  gate291(.a(s_19), .O(gate34inter4));
  nand2 gate292(.a(gate34inter4), .b(gate34inter3), .O(gate34inter5));
  nor2  gate293(.a(gate34inter5), .b(gate34inter2), .O(gate34inter6));
  inv1  gate294(.a(N47), .O(gate34inter7));
  inv1  gate295(.a(N131), .O(gate34inter8));
  nand2 gate296(.a(gate34inter8), .b(gate34inter7), .O(gate34inter9));
  nand2 gate297(.a(s_19), .b(gate34inter3), .O(gate34inter10));
  nor2  gate298(.a(gate34inter10), .b(gate34inter9), .O(gate34inter11));
  nor2  gate299(.a(gate34inter11), .b(gate34inter6), .O(gate34inter12));
  nand2 gate300(.a(gate34inter12), .b(gate34inter1), .O(N187));
nor2 gate35( .a(N53), .b(N131), .O(N188) );
nor2 gate36( .a(N60), .b(N135), .O(N189) );
nor2 gate37( .a(N66), .b(N135), .O(N190) );
nor2 gate38( .a(N73), .b(N139), .O(N191) );
nor2 gate39( .a(N79), .b(N139), .O(N192) );
nor2 gate40( .a(N86), .b(N143), .O(N193) );

  xor2  gate385(.a(N143), .b(N92), .O(gate41inter0));
  nand2 gate386(.a(gate41inter0), .b(s_32), .O(gate41inter1));
  and2  gate387(.a(N143), .b(N92), .O(gate41inter2));
  inv1  gate388(.a(s_32), .O(gate41inter3));
  inv1  gate389(.a(s_33), .O(gate41inter4));
  nand2 gate390(.a(gate41inter4), .b(gate41inter3), .O(gate41inter5));
  nor2  gate391(.a(gate41inter5), .b(gate41inter2), .O(gate41inter6));
  inv1  gate392(.a(N92), .O(gate41inter7));
  inv1  gate393(.a(N143), .O(gate41inter8));
  nand2 gate394(.a(gate41inter8), .b(gate41inter7), .O(gate41inter9));
  nand2 gate395(.a(s_33), .b(gate41inter3), .O(gate41inter10));
  nor2  gate396(.a(gate41inter10), .b(gate41inter9), .O(gate41inter11));
  nor2  gate397(.a(gate41inter11), .b(gate41inter6), .O(gate41inter12));
  nand2 gate398(.a(gate41inter12), .b(gate41inter1), .O(N194));
nor2 gate42( .a(N99), .b(N147), .O(N195) );

  xor2  gate231(.a(N147), .b(N105), .O(gate43inter0));
  nand2 gate232(.a(gate43inter0), .b(s_10), .O(gate43inter1));
  and2  gate233(.a(N147), .b(N105), .O(gate43inter2));
  inv1  gate234(.a(s_10), .O(gate43inter3));
  inv1  gate235(.a(s_11), .O(gate43inter4));
  nand2 gate236(.a(gate43inter4), .b(gate43inter3), .O(gate43inter5));
  nor2  gate237(.a(gate43inter5), .b(gate43inter2), .O(gate43inter6));
  inv1  gate238(.a(N105), .O(gate43inter7));
  inv1  gate239(.a(N147), .O(gate43inter8));
  nand2 gate240(.a(gate43inter8), .b(gate43inter7), .O(gate43inter9));
  nand2 gate241(.a(s_11), .b(gate43inter3), .O(gate43inter10));
  nor2  gate242(.a(gate43inter10), .b(gate43inter9), .O(gate43inter11));
  nor2  gate243(.a(gate43inter11), .b(gate43inter6), .O(gate43inter12));
  nand2 gate244(.a(gate43inter12), .b(gate43inter1), .O(N196));
nor2 gate44( .a(N112), .b(N151), .O(N197) );
nor2 gate45( .a(N115), .b(N151), .O(N198) );
and9 gate46( .a(N154), .b(N159), .c(N162), .d(N165), .e(N168), .f(N171), .g(N174), .h(N177), .i(N180), .O(N199) );
inv1 gate47( .a(N199), .O(N203) );
inv1 gate48( .a(N199), .O(N213) );
inv1 gate49( .a(N199), .O(N223) );
xor2 gate50( .a(N203), .b(N154), .O(N224) );
xor2 gate51( .a(N203), .b(N159), .O(N227) );
xor2 gate52( .a(N203), .b(N162), .O(N230) );

  xor2  gate399(.a(N165), .b(N203), .O(gate53inter0));
  nand2 gate400(.a(gate53inter0), .b(s_34), .O(gate53inter1));
  and2  gate401(.a(N165), .b(N203), .O(gate53inter2));
  inv1  gate402(.a(s_34), .O(gate53inter3));
  inv1  gate403(.a(s_35), .O(gate53inter4));
  nand2 gate404(.a(gate53inter4), .b(gate53inter3), .O(gate53inter5));
  nor2  gate405(.a(gate53inter5), .b(gate53inter2), .O(gate53inter6));
  inv1  gate406(.a(N203), .O(gate53inter7));
  inv1  gate407(.a(N165), .O(gate53inter8));
  nand2 gate408(.a(gate53inter8), .b(gate53inter7), .O(gate53inter9));
  nand2 gate409(.a(s_35), .b(gate53inter3), .O(gate53inter10));
  nor2  gate410(.a(gate53inter10), .b(gate53inter9), .O(gate53inter11));
  nor2  gate411(.a(gate53inter11), .b(gate53inter6), .O(gate53inter12));
  nand2 gate412(.a(gate53inter12), .b(gate53inter1), .O(N233));
xor2 gate54( .a(N203), .b(N168), .O(N236) );

  xor2  gate413(.a(N171), .b(N203), .O(gate55inter0));
  nand2 gate414(.a(gate55inter0), .b(s_36), .O(gate55inter1));
  and2  gate415(.a(N171), .b(N203), .O(gate55inter2));
  inv1  gate416(.a(s_36), .O(gate55inter3));
  inv1  gate417(.a(s_37), .O(gate55inter4));
  nand2 gate418(.a(gate55inter4), .b(gate55inter3), .O(gate55inter5));
  nor2  gate419(.a(gate55inter5), .b(gate55inter2), .O(gate55inter6));
  inv1  gate420(.a(N203), .O(gate55inter7));
  inv1  gate421(.a(N171), .O(gate55inter8));
  nand2 gate422(.a(gate55inter8), .b(gate55inter7), .O(gate55inter9));
  nand2 gate423(.a(s_37), .b(gate55inter3), .O(gate55inter10));
  nor2  gate424(.a(gate55inter10), .b(gate55inter9), .O(gate55inter11));
  nor2  gate425(.a(gate55inter11), .b(gate55inter6), .O(gate55inter12));
  nand2 gate426(.a(gate55inter12), .b(gate55inter1), .O(N239));
nand2 gate56( .a(N1), .b(N213), .O(N242) );

  xor2  gate203(.a(N174), .b(N203), .O(gate57inter0));
  nand2 gate204(.a(gate57inter0), .b(s_6), .O(gate57inter1));
  and2  gate205(.a(N174), .b(N203), .O(gate57inter2));
  inv1  gate206(.a(s_6), .O(gate57inter3));
  inv1  gate207(.a(s_7), .O(gate57inter4));
  nand2 gate208(.a(gate57inter4), .b(gate57inter3), .O(gate57inter5));
  nor2  gate209(.a(gate57inter5), .b(gate57inter2), .O(gate57inter6));
  inv1  gate210(.a(N203), .O(gate57inter7));
  inv1  gate211(.a(N174), .O(gate57inter8));
  nand2 gate212(.a(gate57inter8), .b(gate57inter7), .O(gate57inter9));
  nand2 gate213(.a(s_7), .b(gate57inter3), .O(gate57inter10));
  nor2  gate214(.a(gate57inter10), .b(gate57inter9), .O(gate57inter11));
  nor2  gate215(.a(gate57inter11), .b(gate57inter6), .O(gate57inter12));
  nand2 gate216(.a(gate57inter12), .b(gate57inter1), .O(N243));
nand2 gate58( .a(N213), .b(N11), .O(N246) );
xor2 gate59( .a(N203), .b(N177), .O(N247) );
nand2 gate60( .a(N213), .b(N24), .O(N250) );

  xor2  gate553(.a(N180), .b(N203), .O(gate61inter0));
  nand2 gate554(.a(gate61inter0), .b(s_56), .O(gate61inter1));
  and2  gate555(.a(N180), .b(N203), .O(gate61inter2));
  inv1  gate556(.a(s_56), .O(gate61inter3));
  inv1  gate557(.a(s_57), .O(gate61inter4));
  nand2 gate558(.a(gate61inter4), .b(gate61inter3), .O(gate61inter5));
  nor2  gate559(.a(gate61inter5), .b(gate61inter2), .O(gate61inter6));
  inv1  gate560(.a(N203), .O(gate61inter7));
  inv1  gate561(.a(N180), .O(gate61inter8));
  nand2 gate562(.a(gate61inter8), .b(gate61inter7), .O(gate61inter9));
  nand2 gate563(.a(s_57), .b(gate61inter3), .O(gate61inter10));
  nor2  gate564(.a(gate61inter10), .b(gate61inter9), .O(gate61inter11));
  nor2  gate565(.a(gate61inter11), .b(gate61inter6), .O(gate61inter12));
  nand2 gate566(.a(gate61inter12), .b(gate61inter1), .O(N251));

  xor2  gate525(.a(N37), .b(N213), .O(gate62inter0));
  nand2 gate526(.a(gate62inter0), .b(s_52), .O(gate62inter1));
  and2  gate527(.a(N37), .b(N213), .O(gate62inter2));
  inv1  gate528(.a(s_52), .O(gate62inter3));
  inv1  gate529(.a(s_53), .O(gate62inter4));
  nand2 gate530(.a(gate62inter4), .b(gate62inter3), .O(gate62inter5));
  nor2  gate531(.a(gate62inter5), .b(gate62inter2), .O(gate62inter6));
  inv1  gate532(.a(N213), .O(gate62inter7));
  inv1  gate533(.a(N37), .O(gate62inter8));
  nand2 gate534(.a(gate62inter8), .b(gate62inter7), .O(gate62inter9));
  nand2 gate535(.a(s_53), .b(gate62inter3), .O(gate62inter10));
  nor2  gate536(.a(gate62inter10), .b(gate62inter9), .O(gate62inter11));
  nor2  gate537(.a(gate62inter11), .b(gate62inter6), .O(gate62inter12));
  nand2 gate538(.a(gate62inter12), .b(gate62inter1), .O(N254));
nand2 gate63( .a(N213), .b(N50), .O(N255) );

  xor2  gate427(.a(N63), .b(N213), .O(gate64inter0));
  nand2 gate428(.a(gate64inter0), .b(s_38), .O(gate64inter1));
  and2  gate429(.a(N63), .b(N213), .O(gate64inter2));
  inv1  gate430(.a(s_38), .O(gate64inter3));
  inv1  gate431(.a(s_39), .O(gate64inter4));
  nand2 gate432(.a(gate64inter4), .b(gate64inter3), .O(gate64inter5));
  nor2  gate433(.a(gate64inter5), .b(gate64inter2), .O(gate64inter6));
  inv1  gate434(.a(N213), .O(gate64inter7));
  inv1  gate435(.a(N63), .O(gate64inter8));
  nand2 gate436(.a(gate64inter8), .b(gate64inter7), .O(gate64inter9));
  nand2 gate437(.a(s_39), .b(gate64inter3), .O(gate64inter10));
  nor2  gate438(.a(gate64inter10), .b(gate64inter9), .O(gate64inter11));
  nor2  gate439(.a(gate64inter11), .b(gate64inter6), .O(gate64inter12));
  nand2 gate440(.a(gate64inter12), .b(gate64inter1), .O(N256));
nand2 gate65( .a(N213), .b(N76), .O(N257) );
nand2 gate66( .a(N213), .b(N89), .O(N258) );
nand2 gate67( .a(N213), .b(N102), .O(N259) );
nand2 gate68( .a(N224), .b(N157), .O(N260) );

  xor2  gate259(.a(N158), .b(N224), .O(gate69inter0));
  nand2 gate260(.a(gate69inter0), .b(s_14), .O(gate69inter1));
  and2  gate261(.a(N158), .b(N224), .O(gate69inter2));
  inv1  gate262(.a(s_14), .O(gate69inter3));
  inv1  gate263(.a(s_15), .O(gate69inter4));
  nand2 gate264(.a(gate69inter4), .b(gate69inter3), .O(gate69inter5));
  nor2  gate265(.a(gate69inter5), .b(gate69inter2), .O(gate69inter6));
  inv1  gate266(.a(N224), .O(gate69inter7));
  inv1  gate267(.a(N158), .O(gate69inter8));
  nand2 gate268(.a(gate69inter8), .b(gate69inter7), .O(gate69inter9));
  nand2 gate269(.a(s_15), .b(gate69inter3), .O(gate69inter10));
  nor2  gate270(.a(gate69inter10), .b(gate69inter9), .O(gate69inter11));
  nor2  gate271(.a(gate69inter11), .b(gate69inter6), .O(gate69inter12));
  nand2 gate272(.a(gate69inter12), .b(gate69inter1), .O(N263));
nand2 gate70( .a(N227), .b(N183), .O(N264) );
nand2 gate71( .a(N230), .b(N185), .O(N267) );

  xor2  gate511(.a(N187), .b(N233), .O(gate72inter0));
  nand2 gate512(.a(gate72inter0), .b(s_50), .O(gate72inter1));
  and2  gate513(.a(N187), .b(N233), .O(gate72inter2));
  inv1  gate514(.a(s_50), .O(gate72inter3));
  inv1  gate515(.a(s_51), .O(gate72inter4));
  nand2 gate516(.a(gate72inter4), .b(gate72inter3), .O(gate72inter5));
  nor2  gate517(.a(gate72inter5), .b(gate72inter2), .O(gate72inter6));
  inv1  gate518(.a(N233), .O(gate72inter7));
  inv1  gate519(.a(N187), .O(gate72inter8));
  nand2 gate520(.a(gate72inter8), .b(gate72inter7), .O(gate72inter9));
  nand2 gate521(.a(s_51), .b(gate72inter3), .O(gate72inter10));
  nor2  gate522(.a(gate72inter10), .b(gate72inter9), .O(gate72inter11));
  nor2  gate523(.a(gate72inter11), .b(gate72inter6), .O(gate72inter12));
  nand2 gate524(.a(gate72inter12), .b(gate72inter1), .O(N270));

  xor2  gate581(.a(N189), .b(N236), .O(gate73inter0));
  nand2 gate582(.a(gate73inter0), .b(s_60), .O(gate73inter1));
  and2  gate583(.a(N189), .b(N236), .O(gate73inter2));
  inv1  gate584(.a(s_60), .O(gate73inter3));
  inv1  gate585(.a(s_61), .O(gate73inter4));
  nand2 gate586(.a(gate73inter4), .b(gate73inter3), .O(gate73inter5));
  nor2  gate587(.a(gate73inter5), .b(gate73inter2), .O(gate73inter6));
  inv1  gate588(.a(N236), .O(gate73inter7));
  inv1  gate589(.a(N189), .O(gate73inter8));
  nand2 gate590(.a(gate73inter8), .b(gate73inter7), .O(gate73inter9));
  nand2 gate591(.a(s_61), .b(gate73inter3), .O(gate73inter10));
  nor2  gate592(.a(gate73inter10), .b(gate73inter9), .O(gate73inter11));
  nor2  gate593(.a(gate73inter11), .b(gate73inter6), .O(gate73inter12));
  nand2 gate594(.a(gate73inter12), .b(gate73inter1), .O(N273));

  xor2  gate245(.a(N191), .b(N239), .O(gate74inter0));
  nand2 gate246(.a(gate74inter0), .b(s_12), .O(gate74inter1));
  and2  gate247(.a(N191), .b(N239), .O(gate74inter2));
  inv1  gate248(.a(s_12), .O(gate74inter3));
  inv1  gate249(.a(s_13), .O(gate74inter4));
  nand2 gate250(.a(gate74inter4), .b(gate74inter3), .O(gate74inter5));
  nor2  gate251(.a(gate74inter5), .b(gate74inter2), .O(gate74inter6));
  inv1  gate252(.a(N239), .O(gate74inter7));
  inv1  gate253(.a(N191), .O(gate74inter8));
  nand2 gate254(.a(gate74inter8), .b(gate74inter7), .O(gate74inter9));
  nand2 gate255(.a(s_13), .b(gate74inter3), .O(gate74inter10));
  nor2  gate256(.a(gate74inter10), .b(gate74inter9), .O(gate74inter11));
  nor2  gate257(.a(gate74inter11), .b(gate74inter6), .O(gate74inter12));
  nand2 gate258(.a(gate74inter12), .b(gate74inter1), .O(N276));
nand2 gate75( .a(N243), .b(N193), .O(N279) );

  xor2  gate539(.a(N195), .b(N247), .O(gate76inter0));
  nand2 gate540(.a(gate76inter0), .b(s_54), .O(gate76inter1));
  and2  gate541(.a(N195), .b(N247), .O(gate76inter2));
  inv1  gate542(.a(s_54), .O(gate76inter3));
  inv1  gate543(.a(s_55), .O(gate76inter4));
  nand2 gate544(.a(gate76inter4), .b(gate76inter3), .O(gate76inter5));
  nor2  gate545(.a(gate76inter5), .b(gate76inter2), .O(gate76inter6));
  inv1  gate546(.a(N247), .O(gate76inter7));
  inv1  gate547(.a(N195), .O(gate76inter8));
  nand2 gate548(.a(gate76inter8), .b(gate76inter7), .O(gate76inter9));
  nand2 gate549(.a(s_55), .b(gate76inter3), .O(gate76inter10));
  nor2  gate550(.a(gate76inter10), .b(gate76inter9), .O(gate76inter11));
  nor2  gate551(.a(gate76inter11), .b(gate76inter6), .O(gate76inter12));
  nand2 gate552(.a(gate76inter12), .b(gate76inter1), .O(N282));
nand2 gate77( .a(N251), .b(N197), .O(N285) );

  xor2  gate273(.a(N184), .b(N227), .O(gate78inter0));
  nand2 gate274(.a(gate78inter0), .b(s_16), .O(gate78inter1));
  and2  gate275(.a(N184), .b(N227), .O(gate78inter2));
  inv1  gate276(.a(s_16), .O(gate78inter3));
  inv1  gate277(.a(s_17), .O(gate78inter4));
  nand2 gate278(.a(gate78inter4), .b(gate78inter3), .O(gate78inter5));
  nor2  gate279(.a(gate78inter5), .b(gate78inter2), .O(gate78inter6));
  inv1  gate280(.a(N227), .O(gate78inter7));
  inv1  gate281(.a(N184), .O(gate78inter8));
  nand2 gate282(.a(gate78inter8), .b(gate78inter7), .O(gate78inter9));
  nand2 gate283(.a(s_17), .b(gate78inter3), .O(gate78inter10));
  nor2  gate284(.a(gate78inter10), .b(gate78inter9), .O(gate78inter11));
  nor2  gate285(.a(gate78inter11), .b(gate78inter6), .O(gate78inter12));
  nand2 gate286(.a(gate78inter12), .b(gate78inter1), .O(N288));
nand2 gate79( .a(N230), .b(N186), .O(N289) );

  xor2  gate357(.a(N188), .b(N233), .O(gate80inter0));
  nand2 gate358(.a(gate80inter0), .b(s_28), .O(gate80inter1));
  and2  gate359(.a(N188), .b(N233), .O(gate80inter2));
  inv1  gate360(.a(s_28), .O(gate80inter3));
  inv1  gate361(.a(s_29), .O(gate80inter4));
  nand2 gate362(.a(gate80inter4), .b(gate80inter3), .O(gate80inter5));
  nor2  gate363(.a(gate80inter5), .b(gate80inter2), .O(gate80inter6));
  inv1  gate364(.a(N233), .O(gate80inter7));
  inv1  gate365(.a(N188), .O(gate80inter8));
  nand2 gate366(.a(gate80inter8), .b(gate80inter7), .O(gate80inter9));
  nand2 gate367(.a(s_29), .b(gate80inter3), .O(gate80inter10));
  nor2  gate368(.a(gate80inter10), .b(gate80inter9), .O(gate80inter11));
  nor2  gate369(.a(gate80inter11), .b(gate80inter6), .O(gate80inter12));
  nand2 gate370(.a(gate80inter12), .b(gate80inter1), .O(N290));
nand2 gate81( .a(N236), .b(N190), .O(N291) );

  xor2  gate469(.a(N192), .b(N239), .O(gate82inter0));
  nand2 gate470(.a(gate82inter0), .b(s_44), .O(gate82inter1));
  and2  gate471(.a(N192), .b(N239), .O(gate82inter2));
  inv1  gate472(.a(s_44), .O(gate82inter3));
  inv1  gate473(.a(s_45), .O(gate82inter4));
  nand2 gate474(.a(gate82inter4), .b(gate82inter3), .O(gate82inter5));
  nor2  gate475(.a(gate82inter5), .b(gate82inter2), .O(gate82inter6));
  inv1  gate476(.a(N239), .O(gate82inter7));
  inv1  gate477(.a(N192), .O(gate82inter8));
  nand2 gate478(.a(gate82inter8), .b(gate82inter7), .O(gate82inter9));
  nand2 gate479(.a(s_45), .b(gate82inter3), .O(gate82inter10));
  nor2  gate480(.a(gate82inter10), .b(gate82inter9), .O(gate82inter11));
  nor2  gate481(.a(gate82inter11), .b(gate82inter6), .O(gate82inter12));
  nand2 gate482(.a(gate82inter12), .b(gate82inter1), .O(N292));

  xor2  gate175(.a(N194), .b(N243), .O(gate83inter0));
  nand2 gate176(.a(gate83inter0), .b(s_2), .O(gate83inter1));
  and2  gate177(.a(N194), .b(N243), .O(gate83inter2));
  inv1  gate178(.a(s_2), .O(gate83inter3));
  inv1  gate179(.a(s_3), .O(gate83inter4));
  nand2 gate180(.a(gate83inter4), .b(gate83inter3), .O(gate83inter5));
  nor2  gate181(.a(gate83inter5), .b(gate83inter2), .O(gate83inter6));
  inv1  gate182(.a(N243), .O(gate83inter7));
  inv1  gate183(.a(N194), .O(gate83inter8));
  nand2 gate184(.a(gate83inter8), .b(gate83inter7), .O(gate83inter9));
  nand2 gate185(.a(s_3), .b(gate83inter3), .O(gate83inter10));
  nor2  gate186(.a(gate83inter10), .b(gate83inter9), .O(gate83inter11));
  nor2  gate187(.a(gate83inter11), .b(gate83inter6), .O(gate83inter12));
  nand2 gate188(.a(gate83inter12), .b(gate83inter1), .O(N293));
nand2 gate84( .a(N247), .b(N196), .O(N294) );
nand2 gate85( .a(N251), .b(N198), .O(N295) );
and9 gate86( .a(N260), .b(N264), .c(N267), .d(N270), .e(N273), .f(N276), .g(N279), .h(N282), .i(N285), .O(N296) );
inv1 gate87( .a(N263), .O(N300) );
inv1 gate88( .a(N288), .O(N301) );
inv1 gate89( .a(N289), .O(N302) );
inv1 gate90( .a(N290), .O(N303) );
inv1 gate91( .a(N291), .O(N304) );
inv1 gate92( .a(N292), .O(N305) );
inv1 gate93( .a(N293), .O(N306) );
inv1 gate94( .a(N294), .O(N307) );
inv1 gate95( .a(N295), .O(N308) );
inv1 gate96( .a(N296), .O(N309) );
inv1 gate97( .a(N296), .O(N319) );
inv1 gate98( .a(N296), .O(N329) );
xor2 gate99( .a(N309), .b(N260), .O(N330) );
xor2 gate100( .a(N309), .b(N264), .O(N331) );
xor2 gate101( .a(N309), .b(N267), .O(N332) );

  xor2  gate329(.a(N270), .b(N309), .O(gate102inter0));
  nand2 gate330(.a(gate102inter0), .b(s_24), .O(gate102inter1));
  and2  gate331(.a(N270), .b(N309), .O(gate102inter2));
  inv1  gate332(.a(s_24), .O(gate102inter3));
  inv1  gate333(.a(s_25), .O(gate102inter4));
  nand2 gate334(.a(gate102inter4), .b(gate102inter3), .O(gate102inter5));
  nor2  gate335(.a(gate102inter5), .b(gate102inter2), .O(gate102inter6));
  inv1  gate336(.a(N309), .O(gate102inter7));
  inv1  gate337(.a(N270), .O(gate102inter8));
  nand2 gate338(.a(gate102inter8), .b(gate102inter7), .O(gate102inter9));
  nand2 gate339(.a(s_25), .b(gate102inter3), .O(gate102inter10));
  nor2  gate340(.a(gate102inter10), .b(gate102inter9), .O(gate102inter11));
  nor2  gate341(.a(gate102inter11), .b(gate102inter6), .O(gate102inter12));
  nand2 gate342(.a(gate102inter12), .b(gate102inter1), .O(N333));
nand2 gate103( .a(N8), .b(N319), .O(N334) );
xor2 gate104( .a(N309), .b(N273), .O(N335) );
nand2 gate105( .a(N319), .b(N21), .O(N336) );
xor2 gate106( .a(N309), .b(N276), .O(N337) );

  xor2  gate483(.a(N34), .b(N319), .O(gate107inter0));
  nand2 gate484(.a(gate107inter0), .b(s_46), .O(gate107inter1));
  and2  gate485(.a(N34), .b(N319), .O(gate107inter2));
  inv1  gate486(.a(s_46), .O(gate107inter3));
  inv1  gate487(.a(s_47), .O(gate107inter4));
  nand2 gate488(.a(gate107inter4), .b(gate107inter3), .O(gate107inter5));
  nor2  gate489(.a(gate107inter5), .b(gate107inter2), .O(gate107inter6));
  inv1  gate490(.a(N319), .O(gate107inter7));
  inv1  gate491(.a(N34), .O(gate107inter8));
  nand2 gate492(.a(gate107inter8), .b(gate107inter7), .O(gate107inter9));
  nand2 gate493(.a(s_47), .b(gate107inter3), .O(gate107inter10));
  nor2  gate494(.a(gate107inter10), .b(gate107inter9), .O(gate107inter11));
  nor2  gate495(.a(gate107inter11), .b(gate107inter6), .O(gate107inter12));
  nand2 gate496(.a(gate107inter12), .b(gate107inter1), .O(N338));
xor2 gate108( .a(N309), .b(N279), .O(N339) );

  xor2  gate441(.a(N47), .b(N319), .O(gate109inter0));
  nand2 gate442(.a(gate109inter0), .b(s_40), .O(gate109inter1));
  and2  gate443(.a(N47), .b(N319), .O(gate109inter2));
  inv1  gate444(.a(s_40), .O(gate109inter3));
  inv1  gate445(.a(s_41), .O(gate109inter4));
  nand2 gate446(.a(gate109inter4), .b(gate109inter3), .O(gate109inter5));
  nor2  gate447(.a(gate109inter5), .b(gate109inter2), .O(gate109inter6));
  inv1  gate448(.a(N319), .O(gate109inter7));
  inv1  gate449(.a(N47), .O(gate109inter8));
  nand2 gate450(.a(gate109inter8), .b(gate109inter7), .O(gate109inter9));
  nand2 gate451(.a(s_41), .b(gate109inter3), .O(gate109inter10));
  nor2  gate452(.a(gate109inter10), .b(gate109inter9), .O(gate109inter11));
  nor2  gate453(.a(gate109inter11), .b(gate109inter6), .O(gate109inter12));
  nand2 gate454(.a(gate109inter12), .b(gate109inter1), .O(N340));
xor2 gate110( .a(N309), .b(N282), .O(N341) );

  xor2  gate455(.a(N60), .b(N319), .O(gate111inter0));
  nand2 gate456(.a(gate111inter0), .b(s_42), .O(gate111inter1));
  and2  gate457(.a(N60), .b(N319), .O(gate111inter2));
  inv1  gate458(.a(s_42), .O(gate111inter3));
  inv1  gate459(.a(s_43), .O(gate111inter4));
  nand2 gate460(.a(gate111inter4), .b(gate111inter3), .O(gate111inter5));
  nor2  gate461(.a(gate111inter5), .b(gate111inter2), .O(gate111inter6));
  inv1  gate462(.a(N319), .O(gate111inter7));
  inv1  gate463(.a(N60), .O(gate111inter8));
  nand2 gate464(.a(gate111inter8), .b(gate111inter7), .O(gate111inter9));
  nand2 gate465(.a(s_43), .b(gate111inter3), .O(gate111inter10));
  nor2  gate466(.a(gate111inter10), .b(gate111inter9), .O(gate111inter11));
  nor2  gate467(.a(gate111inter11), .b(gate111inter6), .O(gate111inter12));
  nand2 gate468(.a(gate111inter12), .b(gate111inter1), .O(N342));
xor2 gate112( .a(N309), .b(N285), .O(N343) );
nand2 gate113( .a(N319), .b(N73), .O(N344) );
nand2 gate114( .a(N319), .b(N86), .O(N345) );
nand2 gate115( .a(N319), .b(N99), .O(N346) );

  xor2  gate371(.a(N112), .b(N319), .O(gate116inter0));
  nand2 gate372(.a(gate116inter0), .b(s_30), .O(gate116inter1));
  and2  gate373(.a(N112), .b(N319), .O(gate116inter2));
  inv1  gate374(.a(s_30), .O(gate116inter3));
  inv1  gate375(.a(s_31), .O(gate116inter4));
  nand2 gate376(.a(gate116inter4), .b(gate116inter3), .O(gate116inter5));
  nor2  gate377(.a(gate116inter5), .b(gate116inter2), .O(gate116inter6));
  inv1  gate378(.a(N319), .O(gate116inter7));
  inv1  gate379(.a(N112), .O(gate116inter8));
  nand2 gate380(.a(gate116inter8), .b(gate116inter7), .O(gate116inter9));
  nand2 gate381(.a(s_31), .b(gate116inter3), .O(gate116inter10));
  nor2  gate382(.a(gate116inter10), .b(gate116inter9), .O(gate116inter11));
  nor2  gate383(.a(gate116inter11), .b(gate116inter6), .O(gate116inter12));
  nand2 gate384(.a(gate116inter12), .b(gate116inter1), .O(N347));

  xor2  gate315(.a(N300), .b(N330), .O(gate117inter0));
  nand2 gate316(.a(gate117inter0), .b(s_22), .O(gate117inter1));
  and2  gate317(.a(N300), .b(N330), .O(gate117inter2));
  inv1  gate318(.a(s_22), .O(gate117inter3));
  inv1  gate319(.a(s_23), .O(gate117inter4));
  nand2 gate320(.a(gate117inter4), .b(gate117inter3), .O(gate117inter5));
  nor2  gate321(.a(gate117inter5), .b(gate117inter2), .O(gate117inter6));
  inv1  gate322(.a(N330), .O(gate117inter7));
  inv1  gate323(.a(N300), .O(gate117inter8));
  nand2 gate324(.a(gate117inter8), .b(gate117inter7), .O(gate117inter9));
  nand2 gate325(.a(s_23), .b(gate117inter3), .O(gate117inter10));
  nor2  gate326(.a(gate117inter10), .b(gate117inter9), .O(gate117inter11));
  nor2  gate327(.a(gate117inter11), .b(gate117inter6), .O(gate117inter12));
  nand2 gate328(.a(gate117inter12), .b(gate117inter1), .O(N348));
nand2 gate118( .a(N331), .b(N301), .O(N349) );

  xor2  gate567(.a(N302), .b(N332), .O(gate119inter0));
  nand2 gate568(.a(gate119inter0), .b(s_58), .O(gate119inter1));
  and2  gate569(.a(N302), .b(N332), .O(gate119inter2));
  inv1  gate570(.a(s_58), .O(gate119inter3));
  inv1  gate571(.a(s_59), .O(gate119inter4));
  nand2 gate572(.a(gate119inter4), .b(gate119inter3), .O(gate119inter5));
  nor2  gate573(.a(gate119inter5), .b(gate119inter2), .O(gate119inter6));
  inv1  gate574(.a(N332), .O(gate119inter7));
  inv1  gate575(.a(N302), .O(gate119inter8));
  nand2 gate576(.a(gate119inter8), .b(gate119inter7), .O(gate119inter9));
  nand2 gate577(.a(s_59), .b(gate119inter3), .O(gate119inter10));
  nor2  gate578(.a(gate119inter10), .b(gate119inter9), .O(gate119inter11));
  nor2  gate579(.a(gate119inter11), .b(gate119inter6), .O(gate119inter12));
  nand2 gate580(.a(gate119inter12), .b(gate119inter1), .O(N350));
nand2 gate120( .a(N333), .b(N303), .O(N351) );
nand2 gate121( .a(N335), .b(N304), .O(N352) );
nand2 gate122( .a(N337), .b(N305), .O(N353) );

  xor2  gate217(.a(N306), .b(N339), .O(gate123inter0));
  nand2 gate218(.a(gate123inter0), .b(s_8), .O(gate123inter1));
  and2  gate219(.a(N306), .b(N339), .O(gate123inter2));
  inv1  gate220(.a(s_8), .O(gate123inter3));
  inv1  gate221(.a(s_9), .O(gate123inter4));
  nand2 gate222(.a(gate123inter4), .b(gate123inter3), .O(gate123inter5));
  nor2  gate223(.a(gate123inter5), .b(gate123inter2), .O(gate123inter6));
  inv1  gate224(.a(N339), .O(gate123inter7));
  inv1  gate225(.a(N306), .O(gate123inter8));
  nand2 gate226(.a(gate123inter8), .b(gate123inter7), .O(gate123inter9));
  nand2 gate227(.a(s_9), .b(gate123inter3), .O(gate123inter10));
  nor2  gate228(.a(gate123inter10), .b(gate123inter9), .O(gate123inter11));
  nor2  gate229(.a(gate123inter11), .b(gate123inter6), .O(gate123inter12));
  nand2 gate230(.a(gate123inter12), .b(gate123inter1), .O(N354));

  xor2  gate189(.a(N307), .b(N341), .O(gate124inter0));
  nand2 gate190(.a(gate124inter0), .b(s_4), .O(gate124inter1));
  and2  gate191(.a(N307), .b(N341), .O(gate124inter2));
  inv1  gate192(.a(s_4), .O(gate124inter3));
  inv1  gate193(.a(s_5), .O(gate124inter4));
  nand2 gate194(.a(gate124inter4), .b(gate124inter3), .O(gate124inter5));
  nor2  gate195(.a(gate124inter5), .b(gate124inter2), .O(gate124inter6));
  inv1  gate196(.a(N341), .O(gate124inter7));
  inv1  gate197(.a(N307), .O(gate124inter8));
  nand2 gate198(.a(gate124inter8), .b(gate124inter7), .O(gate124inter9));
  nand2 gate199(.a(s_5), .b(gate124inter3), .O(gate124inter10));
  nor2  gate200(.a(gate124inter10), .b(gate124inter9), .O(gate124inter11));
  nor2  gate201(.a(gate124inter11), .b(gate124inter6), .O(gate124inter12));
  nand2 gate202(.a(gate124inter12), .b(gate124inter1), .O(N355));
nand2 gate125( .a(N343), .b(N308), .O(N356) );
and9 gate126( .a(N348), .b(N349), .c(N350), .d(N351), .e(N352), .f(N353), .g(N354), .h(N355), .i(N356), .O(N357) );
inv1 gate127( .a(N357), .O(N360) );
inv1 gate128( .a(N357), .O(N370) );
nand2 gate129( .a(N14), .b(N360), .O(N371) );
nand2 gate130( .a(N360), .b(N27), .O(N372) );
nand2 gate131( .a(N360), .b(N40), .O(N373) );

  xor2  gate343(.a(N53), .b(N360), .O(gate132inter0));
  nand2 gate344(.a(gate132inter0), .b(s_26), .O(gate132inter1));
  and2  gate345(.a(N53), .b(N360), .O(gate132inter2));
  inv1  gate346(.a(s_26), .O(gate132inter3));
  inv1  gate347(.a(s_27), .O(gate132inter4));
  nand2 gate348(.a(gate132inter4), .b(gate132inter3), .O(gate132inter5));
  nor2  gate349(.a(gate132inter5), .b(gate132inter2), .O(gate132inter6));
  inv1  gate350(.a(N360), .O(gate132inter7));
  inv1  gate351(.a(N53), .O(gate132inter8));
  nand2 gate352(.a(gate132inter8), .b(gate132inter7), .O(gate132inter9));
  nand2 gate353(.a(s_27), .b(gate132inter3), .O(gate132inter10));
  nor2  gate354(.a(gate132inter10), .b(gate132inter9), .O(gate132inter11));
  nor2  gate355(.a(gate132inter11), .b(gate132inter6), .O(gate132inter12));
  nand2 gate356(.a(gate132inter12), .b(gate132inter1), .O(N374));
nand2 gate133( .a(N360), .b(N66), .O(N375) );
nand2 gate134( .a(N360), .b(N79), .O(N376) );
nand2 gate135( .a(N360), .b(N92), .O(N377) );

  xor2  gate301(.a(N105), .b(N360), .O(gate136inter0));
  nand2 gate302(.a(gate136inter0), .b(s_20), .O(gate136inter1));
  and2  gate303(.a(N105), .b(N360), .O(gate136inter2));
  inv1  gate304(.a(s_20), .O(gate136inter3));
  inv1  gate305(.a(s_21), .O(gate136inter4));
  nand2 gate306(.a(gate136inter4), .b(gate136inter3), .O(gate136inter5));
  nor2  gate307(.a(gate136inter5), .b(gate136inter2), .O(gate136inter6));
  inv1  gate308(.a(N360), .O(gate136inter7));
  inv1  gate309(.a(N105), .O(gate136inter8));
  nand2 gate310(.a(gate136inter8), .b(gate136inter7), .O(gate136inter9));
  nand2 gate311(.a(s_21), .b(gate136inter3), .O(gate136inter10));
  nor2  gate312(.a(gate136inter10), .b(gate136inter9), .O(gate136inter11));
  nor2  gate313(.a(gate136inter11), .b(gate136inter6), .O(gate136inter12));
  nand2 gate314(.a(gate136inter12), .b(gate136inter1), .O(N378));
nand2 gate137( .a(N360), .b(N115), .O(N379) );
nand4 gate138( .a(N4), .b(N242), .c(N334), .d(N371), .O(N380) );
nand4 gate139( .a(N246), .b(N336), .c(N372), .d(N17), .O(N381) );
nand4 gate140( .a(N250), .b(N338), .c(N373), .d(N30), .O(N386) );
nand4 gate141( .a(N254), .b(N340), .c(N374), .d(N43), .O(N393) );
nand4 gate142( .a(N255), .b(N342), .c(N375), .d(N56), .O(N399) );
nand4 gate143( .a(N256), .b(N344), .c(N376), .d(N69), .O(N404) );
nand4 gate144( .a(N257), .b(N345), .c(N377), .d(N82), .O(N407) );
nand4 gate145( .a(N258), .b(N346), .c(N378), .d(N95), .O(N411) );
nand4 gate146( .a(N259), .b(N347), .c(N379), .d(N108), .O(N414) );
inv1 gate147( .a(N380), .O(N415) );
and8 gate148( .a(N381), .b(N386), .c(N393), .d(N399), .e(N404), .f(N407), .g(N411), .h(N414), .O(N416) );
inv1 gate149( .a(N393), .O(N417) );
inv1 gate150( .a(N404), .O(N418) );
inv1 gate151( .a(N407), .O(N419) );
inv1 gate152( .a(N411), .O(N420) );
nor2 gate153( .a(N415), .b(N416), .O(N421) );
nand2 gate154( .a(N386), .b(N417), .O(N422) );
nand4 gate155( .a(N386), .b(N393), .c(N418), .d(N399), .O(N425) );
nand3 gate156( .a(N399), .b(N393), .c(N419), .O(N428) );
nand4 gate157( .a(N386), .b(N393), .c(N407), .d(N420), .O(N429) );
nand4 gate158( .a(N381), .b(N386), .c(N422), .d(N399), .O(N430) );
nand4 gate159( .a(N381), .b(N386), .c(N425), .d(N428), .O(N431) );
nand4 gate160( .a(N381), .b(N422), .c(N425), .d(N429), .O(N432) );

endmodule