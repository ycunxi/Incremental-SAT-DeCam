module c1908 (N1,N4,N7,N10,N13,N16,N19,N22,N25,N28,
              N31,N34,N37,N40,N43,N46,N49,N53,N56,N60,
              N63,N66,N69,N72,N76,N79,N82,N85,N88,N91,
              N94,N99,N104,N2753,N2754,N2755,N2756,N2762,N2767,N2768,
              N2779,N2780,N2781,N2782,N2783,N2784,N2785,N2786,N2787,N2811,
              N2886,N2887,N2888,N2889,N2890,N2891,N2892,N2899);
input N1,N4,N7,N10,N13,N16,N19,N22,N25,N28,
      N31,N34,N37,N40,N43,N46,N49,N53,N56,N60,
      N63,N66,N69,N72,N76,N79,N82,N85,N88,N91,
      N94,N99,N104;
  input s_0, s_1, s_2, s_3, s_4, s_5, s_6, s_7, s_8, s_9, s_10, s_11, s_12, s_13, s_14, s_15, s_16, s_17, s_18, s_19, s_20, s_21, s_22, s_23, s_24, s_25, s_26, s_27, s_28, s_29, s_30, s_31, s_32, s_33, s_34, s_35, s_36, s_37, s_38, s_39, s_40, s_41, s_42, s_43, s_44, s_45, s_46, s_47, s_48, s_49, s_50, s_51, s_52, s_53, s_54, s_55, s_56, s_57, s_58, s_59, s_60, s_61, s_62, s_63, s_64, s_65, s_66, s_67, s_68, s_69, s_70, s_71, s_72, s_73, s_74, s_75, s_76, s_77, s_78, s_79, s_80, s_81, s_82, s_83, s_84, s_85, s_86, s_87, s_88, s_89, s_90, s_91, s_92, s_93, s_94, s_95, s_96, s_97, s_98, s_99, s_100, s_101, s_102, s_103, s_104, s_105, s_106, s_107, s_108, s_109, s_110, s_111, s_112, s_113, s_114, s_115, s_116, s_117, s_118, s_119, s_120, s_121, s_122, s_123, s_124, s_125, s_126, s_127, s_128, s_129, s_130, s_131, s_132, s_133, s_134, s_135, s_136, s_137, s_138, s_139, s_140, s_141, s_142, s_143, s_144, s_145, s_146, s_147, s_148, s_149, s_150, s_151, s_152, s_153, s_154, s_155, s_156, s_157, s_158, s_159, s_160, s_161, s_162, s_163, s_164, s_165, s_166, s_167, s_168, s_169, s_170, s_171, s_172, s_173, s_174, s_175, s_176, s_177, s_178, s_179, s_180, s_181, s_182, s_183, s_184, s_185, s_186, s_187, s_188, s_189, s_190, s_191, s_192, s_193, s_194, s_195, s_196, s_197, s_198, s_199, s_200, s_201, s_202, s_203, s_204, s_205, s_206, s_207, s_208, s_209, s_210, s_211;
output N2753,N2754,N2755,N2756,N2762,N2767,N2768,N2779,N2780,N2781,
       N2782,N2783,N2784,N2785,N2786,N2787,N2811,N2886,N2887,N2888,
       N2889,N2890,N2891,N2892,N2899;
wire N190,N194,N197,N201,N206,N209,N212,N216,N220,N225,
     N229,N232,N235,N239,N243,N247,N251,N252,N253,N256,
     N257,N260,N263,N266,N269,N272,N275,N276,N277,N280,
     N283,N290,N297,N300,N303,N306,N313,N316,N319,N326,
     N331,N338,N343,N346,N349,N352,N355,N358,N361,N364,
     N367,N370,N373,N376,N379,N382,N385,N388,N534,N535,
     N536,N537,N538,N539,N540,N541,N542,N543,N544,N545,
     N546,N547,N548,N549,N550,N551,N552,N553,N554,N555,
     N556,N559,N562,N565,N568,N571,N574,N577,N580,N583,
     N586,N589,N592,N595,N598,N601,N602,N603,N608,N612,
     N616,N619,N622,N625,N628,N631,N634,N637,N640,N643,
     N646,N649,N652,N655,N658,N661,N664,N667,N670,N673,
     N676,N679,N682,N685,N688,N691,N694,N697,N700,N703,
     N706,N709,N712,N715,N718,N721,N724,N727,N730,N733,
     N736,N739,N742,N745,N748,N751,N886,N887,N888,N889,
     N890,N891,N892,N893,N894,N895,N896,N897,N898,N899,
     N903,N907,N910,N913,N914,N915,N916,N917,N918,N919,
     N920,N921,N922,N923,N926,N935,N938,N939,N942,N943,
     N946,N947,N950,N951,N954,N955,N958,N959,N962,N965,
     N968,N969,N972,N973,N976,N977,N980,N981,N984,N985,
     N988,N989,N990,N991,N992,N993,N994,N997,N998,N1001,
     N1002,N1003,N1004,N1005,N1006,N1007,N1008,N1009,N1010,N1013,
     N1016,N1019,N1022,N1025,N1028,N1031,N1034,N1037,N1040,N1043,
     N1046,N1049,N1054,N1055,N1063,N1064,N1067,N1068,N1119,N1120,
     N1121,N1122,N1128,N1129,N1130,N1131,N1132,N1133,N1148,N1149,
     N1150,N1151,N1152,N1153,N1154,N1155,N1156,N1157,N1158,N1159,
     N1160,N1161,N1162,N1163,N1164,N1167,N1168,N1171,N1188,N1205,
     N1206,N1207,N1208,N1209,N1210,N1211,N1212,N1213,N1214,N1215,
     N1216,N1217,N1218,N1219,N1220,N1221,N1222,N1223,N1224,N1225,
     N1226,N1227,N1228,N1229,N1230,N1231,N1232,N1235,N1238,N1239,
     N1240,N1241,N1242,N1243,N1246,N1249,N1252,N1255,N1258,N1261,
     N1264,N1267,N1309,N1310,N1311,N1312,N1313,N1314,N1315,N1316,
     N1317,N1318,N1319,N1322,N1327,N1328,N1334,N1344,N1345,N1346,
     N1348,N1349,N1350,N1351,N1352,N1355,N1358,N1361,N1364,N1367,
     N1370,N1373,N1376,N1379,N1383,N1386,N1387,N1388,N1389,N1390,
     N1393,N1396,N1397,N1398,N1399,N1409,N1412,N1413,N1416,N1419,
     N1433,N1434,N1438,N1439,N1440,N1443,N1444,N1445,N1446,N1447,
     N1448,N1451,N1452,N1453,N1454,N1455,N1456,N1457,N1458,N1459,
     N1460,N1461,N1462,N1463,N1464,N1468,N1469,N1470,N1471,N1472,
     N1475,N1476,N1478,N1481,N1484,N1487,N1488,N1489,N1490,N1491,
     N1492,N1493,N1494,N1495,N1496,N1498,N1499,N1500,N1501,N1504,
     N1510,N1513,N1514,N1517,N1520,N1521,N1522,N1526,N1527,N1528,
     N1529,N1530,N1531,N1532,N1534,N1537,N1540,N1546,N1554,N1557,
     N1561,N1567,N1568,N1569,N1571,N1576,N1588,N1591,N1593,N1594,
     N1595,N1596,N1600,N1603,N1606,N1609,N1612,N1615,N1620,N1623,
     N1635,N1636,N1638,N1639,N1640,N1643,N1647,N1651,N1658,N1661,
     N1664,N1671,N1672,N1675,N1677,N1678,N1679,N1680,N1681,N1682,
     N1683,N1685,N1688,N1697,N1701,N1706,N1707,N1708,N1709,N1710,
     N1711,N1712,N1713,N1714,N1717,N1720,N1721,N1723,N1727,N1728,
     N1730,N1731,N1734,N1740,N1741,N1742,N1746,N1747,N1748,N1751,
     N1759,N1761,N1762,N1763,N1764,N1768,N1769,N1772,N1773,N1774,
     N1777,N1783,N1784,N1785,N1786,N1787,N1788,N1791,N1792,N1795,
     N1796,N1798,N1801,N1802,N1807,N1808,N1809,N1810,N1812,N1815,
     N1818,N1821,N1822,N1823,N1824,N1825,N1826,N1827,N1830,N1837,
     N1838,N1841,N1848,N1849,N1850,N1852,N1855,N1856,N1857,N1858,
     N1864,N1865,N1866,N1869,N1872,N1875,N1878,N1879,N1882,N1883,
     N1884,N1885,N1889,N1895,N1896,N1897,N1898,N1902,N1910,N1911,
     N1912,N1913,N1915,N1919,N1920,N1921,N1922,N1923,N1924,N1927,
     N1930,N1933,N1936,N1937,N1938,N1941,N1942,N1944,N1947,N1950,
     N1953,N1958,N1961,N1965,N1968,N1975,N1976,N1977,N1978,N1979,
     N1980,N1985,N1987,N1999,N2000,N2002,N2003,N2004,N2005,N2006,
     N2007,N2008,N2009,N2012,N2013,N2014,N2015,N2016,N2018,N2019,
     N2020,N2021,N2022,N2023,N2024,N2025,N2026,N2027,N2030,N2033,
     N2036,N2037,N2038,N2039,N2040,N2041,N2042,N2047,N2052,N2055,
     N2060,N2061,N2062,N2067,N2068,N2071,N2076,N2077,N2078,N2081,
     N2086,N2089,N2104,N2119,N2129,N2143,N2148,N2151,N2196,N2199,
     N2202,N2205,N2214,N2215,N2216,N2217,N2222,N2223,N2224,N2225,
     N2226,N2227,N2228,N2229,N2230,N2231,N2232,N2233,N2234,N2235,
     N2236,N2237,N2240,N2241,N2244,N2245,N2250,N2253,N2256,N2257,
     N2260,N2263,N2266,N2269,N2272,N2279,N2286,N2297,N2315,N2326,
     N2340,N2353,N2361,N2375,N2384,N2385,N2386,N2426,N2427,N2537,
     N2540,N2543,N2546,N2549,N2552,N2555,N2558,N2561,N2564,N2567,
     N2570,N2573,N2576,N2594,N2597,N2600,N2603,N2606,N2611,N2614,
     N2617,N2620,N2627,N2628,N2629,N2630,N2631,N2632,N2633,N2634,
     N2639,N2642,N2645,N2648,N2651,N2655,N2658,N2661,N2664,N2669,
     N2670,N2671,N2672,N2673,N2674,N2675,N2676,N2682,N2683,N2688,
     N2689,N2690,N2691,N2710,N2720,N2721,N2722,N2723,N2724,N2725,
     N2726,N2727,N2728,N2729,N2730,N2731,N2732,N2733,N2734,N2735,
     N2736,N2737,N2738,N2739,N2740,N2741,N2742,N2743,N2744,N2745,
     N2746,N2747,N2750,N2757,N2758,N2759,N2760,N2761,N2763,N2764,
     N2765,N2766,N2773,N2776,N2788,N2789,N2800,N2807,N2808,N2809,
     N2810,N2812,N2815,N2818,N2821,N2824,N2827,N2828,N2829,N2843,
     N2846,N2850,N2851,N2852,N2853,N2854,N2857,N2858,N2859,N2860,
     N2861,N2862,N2863,N2866,N2867,N2868,N2869,N2870,N2871,N2872,
     N2873,N2874,N2875,N2876,N2877,N2878,N2879,N2880,N2881,N2882,
     N2883,N2895,N2896,N2897,N2898, gate300inter0, gate300inter1, gate300inter2, gate300inter3, gate300inter4, gate300inter5, gate300inter6, gate300inter7, gate300inter8, gate300inter9, gate300inter10, gate300inter11, gate300inter12, gate788inter0, gate788inter1, gate788inter2, gate788inter3, gate788inter4, gate788inter5, gate788inter6, gate788inter7, gate788inter8, gate788inter9, gate788inter10, gate788inter11, gate788inter12, gate540inter0, gate540inter1, gate540inter2, gate540inter3, gate540inter4, gate540inter5, gate540inter6, gate540inter7, gate540inter8, gate540inter9, gate540inter10, gate540inter11, gate540inter12, gate322inter0, gate322inter1, gate322inter2, gate322inter3, gate322inter4, gate322inter5, gate322inter6, gate322inter7, gate322inter8, gate322inter9, gate322inter10, gate322inter11, gate322inter12, gate425inter0, gate425inter1, gate425inter2, gate425inter3, gate425inter4, gate425inter5, gate425inter6, gate425inter7, gate425inter8, gate425inter9, gate425inter10, gate425inter11, gate425inter12, gate277inter0, gate277inter1, gate277inter2, gate277inter3, gate277inter4, gate277inter5, gate277inter6, gate277inter7, gate277inter8, gate277inter9, gate277inter10, gate277inter11, gate277inter12, gate161inter0, gate161inter1, gate161inter2, gate161inter3, gate161inter4, gate161inter5, gate161inter6, gate161inter7, gate161inter8, gate161inter9, gate161inter10, gate161inter11, gate161inter12, gate596inter0, gate596inter1, gate596inter2, gate596inter3, gate596inter4, gate596inter5, gate596inter6, gate596inter7, gate596inter8, gate596inter9, gate596inter10, gate596inter11, gate596inter12, gate251inter0, gate251inter1, gate251inter2, gate251inter3, gate251inter4, gate251inter5, gate251inter6, gate251inter7, gate251inter8, gate251inter9, gate251inter10, gate251inter11, gate251inter12, gate610inter0, gate610inter1, gate610inter2, gate610inter3, gate610inter4, gate610inter5, gate610inter6, gate610inter7, gate610inter8, gate610inter9, gate610inter10, gate610inter11, gate610inter12, gate248inter0, gate248inter1, gate248inter2, gate248inter3, gate248inter4, gate248inter5, gate248inter6, gate248inter7, gate248inter8, gate248inter9, gate248inter10, gate248inter11, gate248inter12, gate637inter0, gate637inter1, gate637inter2, gate637inter3, gate637inter4, gate637inter5, gate637inter6, gate637inter7, gate637inter8, gate637inter9, gate637inter10, gate637inter11, gate637inter12, gate314inter0, gate314inter1, gate314inter2, gate314inter3, gate314inter4, gate314inter5, gate314inter6, gate314inter7, gate314inter8, gate314inter9, gate314inter10, gate314inter11, gate314inter12, gate762inter0, gate762inter1, gate762inter2, gate762inter3, gate762inter4, gate762inter5, gate762inter6, gate762inter7, gate762inter8, gate762inter9, gate762inter10, gate762inter11, gate762inter12, gate663inter0, gate663inter1, gate663inter2, gate663inter3, gate663inter4, gate663inter5, gate663inter6, gate663inter7, gate663inter8, gate663inter9, gate663inter10, gate663inter11, gate663inter12, gate364inter0, gate364inter1, gate364inter2, gate364inter3, gate364inter4, gate364inter5, gate364inter6, gate364inter7, gate364inter8, gate364inter9, gate364inter10, gate364inter11, gate364inter12, gate799inter0, gate799inter1, gate799inter2, gate799inter3, gate799inter4, gate799inter5, gate799inter6, gate799inter7, gate799inter8, gate799inter9, gate799inter10, gate799inter11, gate799inter12, gate541inter0, gate541inter1, gate541inter2, gate541inter3, gate541inter4, gate541inter5, gate541inter6, gate541inter7, gate541inter8, gate541inter9, gate541inter10, gate541inter11, gate541inter12, gate862inter0, gate862inter1, gate862inter2, gate862inter3, gate862inter4, gate862inter5, gate862inter6, gate862inter7, gate862inter8, gate862inter9, gate862inter10, gate862inter11, gate862inter12, gate874inter0, gate874inter1, gate874inter2, gate874inter3, gate874inter4, gate874inter5, gate874inter6, gate874inter7, gate874inter8, gate874inter9, gate874inter10, gate874inter11, gate874inter12, gate843inter0, gate843inter1, gate843inter2, gate843inter3, gate843inter4, gate843inter5, gate843inter6, gate843inter7, gate843inter8, gate843inter9, gate843inter10, gate843inter11, gate843inter12, gate483inter0, gate483inter1, gate483inter2, gate483inter3, gate483inter4, gate483inter5, gate483inter6, gate483inter7, gate483inter8, gate483inter9, gate483inter10, gate483inter11, gate483inter12, gate684inter0, gate684inter1, gate684inter2, gate684inter3, gate684inter4, gate684inter5, gate684inter6, gate684inter7, gate684inter8, gate684inter9, gate684inter10, gate684inter11, gate684inter12, gate273inter0, gate273inter1, gate273inter2, gate273inter3, gate273inter4, gate273inter5, gate273inter6, gate273inter7, gate273inter8, gate273inter9, gate273inter10, gate273inter11, gate273inter12, gate345inter0, gate345inter1, gate345inter2, gate345inter3, gate345inter4, gate345inter5, gate345inter6, gate345inter7, gate345inter8, gate345inter9, gate345inter10, gate345inter11, gate345inter12, gate306inter0, gate306inter1, gate306inter2, gate306inter3, gate306inter4, gate306inter5, gate306inter6, gate306inter7, gate306inter8, gate306inter9, gate306inter10, gate306inter11, gate306inter12, gate643inter0, gate643inter1, gate643inter2, gate643inter3, gate643inter4, gate643inter5, gate643inter6, gate643inter7, gate643inter8, gate643inter9, gate643inter10, gate643inter11, gate643inter12, gate824inter0, gate824inter1, gate824inter2, gate824inter3, gate824inter4, gate824inter5, gate824inter6, gate824inter7, gate824inter8, gate824inter9, gate824inter10, gate824inter11, gate824inter12, gate466inter0, gate466inter1, gate466inter2, gate466inter3, gate466inter4, gate466inter5, gate466inter6, gate466inter7, gate466inter8, gate466inter9, gate466inter10, gate466inter11, gate466inter12, gate562inter0, gate562inter1, gate562inter2, gate562inter3, gate562inter4, gate562inter5, gate562inter6, gate562inter7, gate562inter8, gate562inter9, gate562inter10, gate562inter11, gate562inter12, gate819inter0, gate819inter1, gate819inter2, gate819inter3, gate819inter4, gate819inter5, gate819inter6, gate819inter7, gate819inter8, gate819inter9, gate819inter10, gate819inter11, gate819inter12, gate405inter0, gate405inter1, gate405inter2, gate405inter3, gate405inter4, gate405inter5, gate405inter6, gate405inter7, gate405inter8, gate405inter9, gate405inter10, gate405inter11, gate405inter12, gate853inter0, gate853inter1, gate853inter2, gate853inter3, gate853inter4, gate853inter5, gate853inter6, gate853inter7, gate853inter8, gate853inter9, gate853inter10, gate853inter11, gate853inter12, gate665inter0, gate665inter1, gate665inter2, gate665inter3, gate665inter4, gate665inter5, gate665inter6, gate665inter7, gate665inter8, gate665inter9, gate665inter10, gate665inter11, gate665inter12, gate508inter0, gate508inter1, gate508inter2, gate508inter3, gate508inter4, gate508inter5, gate508inter6, gate508inter7, gate508inter8, gate508inter9, gate508inter10, gate508inter11, gate508inter12, gate628inter0, gate628inter1, gate628inter2, gate628inter3, gate628inter4, gate628inter5, gate628inter6, gate628inter7, gate628inter8, gate628inter9, gate628inter10, gate628inter11, gate628inter12, gate632inter0, gate632inter1, gate632inter2, gate632inter3, gate632inter4, gate632inter5, gate632inter6, gate632inter7, gate632inter8, gate632inter9, gate632inter10, gate632inter11, gate632inter12, gate304inter0, gate304inter1, gate304inter2, gate304inter3, gate304inter4, gate304inter5, gate304inter6, gate304inter7, gate304inter8, gate304inter9, gate304inter10, gate304inter11, gate304inter12, gate234inter0, gate234inter1, gate234inter2, gate234inter3, gate234inter4, gate234inter5, gate234inter6, gate234inter7, gate234inter8, gate234inter9, gate234inter10, gate234inter11, gate234inter12, gate75inter0, gate75inter1, gate75inter2, gate75inter3, gate75inter4, gate75inter5, gate75inter6, gate75inter7, gate75inter8, gate75inter9, gate75inter10, gate75inter11, gate75inter12, gate816inter0, gate816inter1, gate816inter2, gate816inter3, gate816inter4, gate816inter5, gate816inter6, gate816inter7, gate816inter8, gate816inter9, gate816inter10, gate816inter11, gate816inter12, gate325inter0, gate325inter1, gate325inter2, gate325inter3, gate325inter4, gate325inter5, gate325inter6, gate325inter7, gate325inter8, gate325inter9, gate325inter10, gate325inter11, gate325inter12, gate79inter0, gate79inter1, gate79inter2, gate79inter3, gate79inter4, gate79inter5, gate79inter6, gate79inter7, gate79inter8, gate79inter9, gate79inter10, gate79inter11, gate79inter12, gate600inter0, gate600inter1, gate600inter2, gate600inter3, gate600inter4, gate600inter5, gate600inter6, gate600inter7, gate600inter8, gate600inter9, gate600inter10, gate600inter11, gate600inter12, gate809inter0, gate809inter1, gate809inter2, gate809inter3, gate809inter4, gate809inter5, gate809inter6, gate809inter7, gate809inter8, gate809inter9, gate809inter10, gate809inter11, gate809inter12, gate511inter0, gate511inter1, gate511inter2, gate511inter3, gate511inter4, gate511inter5, gate511inter6, gate511inter7, gate511inter8, gate511inter9, gate511inter10, gate511inter11, gate511inter12, gate259inter0, gate259inter1, gate259inter2, gate259inter3, gate259inter4, gate259inter5, gate259inter6, gate259inter7, gate259inter8, gate259inter9, gate259inter10, gate259inter11, gate259inter12, gate565inter0, gate565inter1, gate565inter2, gate565inter3, gate565inter4, gate565inter5, gate565inter6, gate565inter7, gate565inter8, gate565inter9, gate565inter10, gate565inter11, gate565inter12, gate559inter0, gate559inter1, gate559inter2, gate559inter3, gate559inter4, gate559inter5, gate559inter6, gate559inter7, gate559inter8, gate559inter9, gate559inter10, gate559inter11, gate559inter12, gate582inter0, gate582inter1, gate582inter2, gate582inter3, gate582inter4, gate582inter5, gate582inter6, gate582inter7, gate582inter8, gate582inter9, gate582inter10, gate582inter11, gate582inter12, gate269inter0, gate269inter1, gate269inter2, gate269inter3, gate269inter4, gate269inter5, gate269inter6, gate269inter7, gate269inter8, gate269inter9, gate269inter10, gate269inter11, gate269inter12, gate319inter0, gate319inter1, gate319inter2, gate319inter3, gate319inter4, gate319inter5, gate319inter6, gate319inter7, gate319inter8, gate319inter9, gate319inter10, gate319inter11, gate319inter12, gate782inter0, gate782inter1, gate782inter2, gate782inter3, gate782inter4, gate782inter5, gate782inter6, gate782inter7, gate782inter8, gate782inter9, gate782inter10, gate782inter11, gate782inter12, gate784inter0, gate784inter1, gate784inter2, gate784inter3, gate784inter4, gate784inter5, gate784inter6, gate784inter7, gate784inter8, gate784inter9, gate784inter10, gate784inter11, gate784inter12, gate812inter0, gate812inter1, gate812inter2, gate812inter3, gate812inter4, gate812inter5, gate812inter6, gate812inter7, gate812inter8, gate812inter9, gate812inter10, gate812inter11, gate812inter12, gate402inter0, gate402inter1, gate402inter2, gate402inter3, gate402inter4, gate402inter5, gate402inter6, gate402inter7, gate402inter8, gate402inter9, gate402inter10, gate402inter11, gate402inter12, gate501inter0, gate501inter1, gate501inter2, gate501inter3, gate501inter4, gate501inter5, gate501inter6, gate501inter7, gate501inter8, gate501inter9, gate501inter10, gate501inter11, gate501inter12, gate394inter0, gate394inter1, gate394inter2, gate394inter3, gate394inter4, gate394inter5, gate394inter6, gate394inter7, gate394inter8, gate394inter9, gate394inter10, gate394inter11, gate394inter12, gate316inter0, gate316inter1, gate316inter2, gate316inter3, gate316inter4, gate316inter5, gate316inter6, gate316inter7, gate316inter8, gate316inter9, gate316inter10, gate316inter11, gate316inter12, gate587inter0, gate587inter1, gate587inter2, gate587inter3, gate587inter4, gate587inter5, gate587inter6, gate587inter7, gate587inter8, gate587inter9, gate587inter10, gate587inter11, gate587inter12, gate510inter0, gate510inter1, gate510inter2, gate510inter3, gate510inter4, gate510inter5, gate510inter6, gate510inter7, gate510inter8, gate510inter9, gate510inter10, gate510inter11, gate510inter12, gate421inter0, gate421inter1, gate421inter2, gate421inter3, gate421inter4, gate421inter5, gate421inter6, gate421inter7, gate421inter8, gate421inter9, gate421inter10, gate421inter11, gate421inter12, gate344inter0, gate344inter1, gate344inter2, gate344inter3, gate344inter4, gate344inter5, gate344inter6, gate344inter7, gate344inter8, gate344inter9, gate344inter10, gate344inter11, gate344inter12, gate415inter0, gate415inter1, gate415inter2, gate415inter3, gate415inter4, gate415inter5, gate415inter6, gate415inter7, gate415inter8, gate415inter9, gate415inter10, gate415inter11, gate415inter12, gate840inter0, gate840inter1, gate840inter2, gate840inter3, gate840inter4, gate840inter5, gate840inter6, gate840inter7, gate840inter8, gate840inter9, gate840inter10, gate840inter11, gate840inter12, gate547inter0, gate547inter1, gate547inter2, gate547inter3, gate547inter4, gate547inter5, gate547inter6, gate547inter7, gate547inter8, gate547inter9, gate547inter10, gate547inter11, gate547inter12, gate552inter0, gate552inter1, gate552inter2, gate552inter3, gate552inter4, gate552inter5, gate552inter6, gate552inter7, gate552inter8, gate552inter9, gate552inter10, gate552inter11, gate552inter12, gate673inter0, gate673inter1, gate673inter2, gate673inter3, gate673inter4, gate673inter5, gate673inter6, gate673inter7, gate673inter8, gate673inter9, gate673inter10, gate673inter11, gate673inter12, gate77inter0, gate77inter1, gate77inter2, gate77inter3, gate77inter4, gate77inter5, gate77inter6, gate77inter7, gate77inter8, gate77inter9, gate77inter10, gate77inter11, gate77inter12, gate235inter0, gate235inter1, gate235inter2, gate235inter3, gate235inter4, gate235inter5, gate235inter6, gate235inter7, gate235inter8, gate235inter9, gate235inter10, gate235inter11, gate235inter12, gate826inter0, gate826inter1, gate826inter2, gate826inter3, gate826inter4, gate826inter5, gate826inter6, gate826inter7, gate826inter8, gate826inter9, gate826inter10, gate826inter11, gate826inter12, gate503inter0, gate503inter1, gate503inter2, gate503inter3, gate503inter4, gate503inter5, gate503inter6, gate503inter7, gate503inter8, gate503inter9, gate503inter10, gate503inter11, gate503inter12, gate336inter0, gate336inter1, gate336inter2, gate336inter3, gate336inter4, gate336inter5, gate336inter6, gate336inter7, gate336inter8, gate336inter9, gate336inter10, gate336inter11, gate336inter12, gate328inter0, gate328inter1, gate328inter2, gate328inter3, gate328inter4, gate328inter5, gate328inter6, gate328inter7, gate328inter8, gate328inter9, gate328inter10, gate328inter11, gate328inter12, gate245inter0, gate245inter1, gate245inter2, gate245inter3, gate245inter4, gate245inter5, gate245inter6, gate245inter7, gate245inter8, gate245inter9, gate245inter10, gate245inter11, gate245inter12, gate98inter0, gate98inter1, gate98inter2, gate98inter3, gate98inter4, gate98inter5, gate98inter6, gate98inter7, gate98inter8, gate98inter9, gate98inter10, gate98inter11, gate98inter12, gate303inter0, gate303inter1, gate303inter2, gate303inter3, gate303inter4, gate303inter5, gate303inter6, gate303inter7, gate303inter8, gate303inter9, gate303inter10, gate303inter11, gate303inter12, gate649inter0, gate649inter1, gate649inter2, gate649inter3, gate649inter4, gate649inter5, gate649inter6, gate649inter7, gate649inter8, gate649inter9, gate649inter10, gate649inter11, gate649inter12, gate856inter0, gate856inter1, gate856inter2, gate856inter3, gate856inter4, gate856inter5, gate856inter6, gate856inter7, gate856inter8, gate856inter9, gate856inter10, gate856inter11, gate856inter12, gate839inter0, gate839inter1, gate839inter2, gate839inter3, gate839inter4, gate839inter5, gate839inter6, gate839inter7, gate839inter8, gate839inter9, gate839inter10, gate839inter11, gate839inter12, gate635inter0, gate635inter1, gate635inter2, gate635inter3, gate635inter4, gate635inter5, gate635inter6, gate635inter7, gate635inter8, gate635inter9, gate635inter10, gate635inter11, gate635inter12, gate343inter0, gate343inter1, gate343inter2, gate343inter3, gate343inter4, gate343inter5, gate343inter6, gate343inter7, gate343inter8, gate343inter9, gate343inter10, gate343inter11, gate343inter12, gate835inter0, gate835inter1, gate835inter2, gate835inter3, gate835inter4, gate835inter5, gate835inter6, gate835inter7, gate835inter8, gate835inter9, gate835inter10, gate835inter11, gate835inter12, gate247inter0, gate247inter1, gate247inter2, gate247inter3, gate247inter4, gate247inter5, gate247inter6, gate247inter7, gate247inter8, gate247inter9, gate247inter10, gate247inter11, gate247inter12, gate558inter0, gate558inter1, gate558inter2, gate558inter3, gate558inter4, gate558inter5, gate558inter6, gate558inter7, gate558inter8, gate558inter9, gate558inter10, gate558inter11, gate558inter12, gate563inter0, gate563inter1, gate563inter2, gate563inter3, gate563inter4, gate563inter5, gate563inter6, gate563inter7, gate563inter8, gate563inter9, gate563inter10, gate563inter11, gate563inter12, gate876inter0, gate876inter1, gate876inter2, gate876inter3, gate876inter4, gate876inter5, gate876inter6, gate876inter7, gate876inter8, gate876inter9, gate876inter10, gate876inter11, gate876inter12, gate754inter0, gate754inter1, gate754inter2, gate754inter3, gate754inter4, gate754inter5, gate754inter6, gate754inter7, gate754inter8, gate754inter9, gate754inter10, gate754inter11, gate754inter12, gate162inter0, gate162inter1, gate162inter2, gate162inter3, gate162inter4, gate162inter5, gate162inter6, gate162inter7, gate162inter8, gate162inter9, gate162inter10, gate162inter11, gate162inter12, gate341inter0, gate341inter1, gate341inter2, gate341inter3, gate341inter4, gate341inter5, gate341inter6, gate341inter7, gate341inter8, gate341inter9, gate341inter10, gate341inter11, gate341inter12, gate675inter0, gate675inter1, gate675inter2, gate675inter3, gate675inter4, gate675inter5, gate675inter6, gate675inter7, gate675inter8, gate675inter9, gate675inter10, gate675inter11, gate675inter12, gate546inter0, gate546inter1, gate546inter2, gate546inter3, gate546inter4, gate546inter5, gate546inter6, gate546inter7, gate546inter8, gate546inter9, gate546inter10, gate546inter11, gate546inter12, gate486inter0, gate486inter1, gate486inter2, gate486inter3, gate486inter4, gate486inter5, gate486inter6, gate486inter7, gate486inter8, gate486inter9, gate486inter10, gate486inter11, gate486inter12, gate500inter0, gate500inter1, gate500inter2, gate500inter3, gate500inter4, gate500inter5, gate500inter6, gate500inter7, gate500inter8, gate500inter9, gate500inter10, gate500inter11, gate500inter12, gate822inter0, gate822inter1, gate822inter2, gate822inter3, gate822inter4, gate822inter5, gate822inter6, gate822inter7, gate822inter8, gate822inter9, gate822inter10, gate822inter11, gate822inter12, gate561inter0, gate561inter1, gate561inter2, gate561inter3, gate561inter4, gate561inter5, gate561inter6, gate561inter7, gate561inter8, gate561inter9, gate561inter10, gate561inter11, gate561inter12, gate326inter0, gate326inter1, gate326inter2, gate326inter3, gate326inter4, gate326inter5, gate326inter6, gate326inter7, gate326inter8, gate326inter9, gate326inter10, gate326inter11, gate326inter12, gate100inter0, gate100inter1, gate100inter2, gate100inter3, gate100inter4, gate100inter5, gate100inter6, gate100inter7, gate100inter8, gate100inter9, gate100inter10, gate100inter11, gate100inter12, gate368inter0, gate368inter1, gate368inter2, gate368inter3, gate368inter4, gate368inter5, gate368inter6, gate368inter7, gate368inter8, gate368inter9, gate368inter10, gate368inter11, gate368inter12, gate305inter0, gate305inter1, gate305inter2, gate305inter3, gate305inter4, gate305inter5, gate305inter6, gate305inter7, gate305inter8, gate305inter9, gate305inter10, gate305inter11, gate305inter12, gate624inter0, gate624inter1, gate624inter2, gate624inter3, gate624inter4, gate624inter5, gate624inter6, gate624inter7, gate624inter8, gate624inter9, gate624inter10, gate624inter11, gate624inter12, gate416inter0, gate416inter1, gate416inter2, gate416inter3, gate416inter4, gate416inter5, gate416inter6, gate416inter7, gate416inter8, gate416inter9, gate416inter10, gate416inter11, gate416inter12, gate865inter0, gate865inter1, gate865inter2, gate865inter3, gate865inter4, gate865inter5, gate865inter6, gate865inter7, gate865inter8, gate865inter9, gate865inter10, gate865inter11, gate865inter12, gate286inter0, gate286inter1, gate286inter2, gate286inter3, gate286inter4, gate286inter5, gate286inter6, gate286inter7, gate286inter8, gate286inter9, gate286inter10, gate286inter11, gate286inter12, gate281inter0, gate281inter1, gate281inter2, gate281inter3, gate281inter4, gate281inter5, gate281inter6, gate281inter7, gate281inter8, gate281inter9, gate281inter10, gate281inter11, gate281inter12, gate403inter0, gate403inter1, gate403inter2, gate403inter3, gate403inter4, gate403inter5, gate403inter6, gate403inter7, gate403inter8, gate403inter9, gate403inter10, gate403inter11, gate403inter12;


inv1 gate1( .a(N1), .O(N190) );
inv1 gate2( .a(N4), .O(N194) );
inv1 gate3( .a(N7), .O(N197) );
inv1 gate4( .a(N10), .O(N201) );
inv1 gate5( .a(N13), .O(N206) );
inv1 gate6( .a(N16), .O(N209) );
inv1 gate7( .a(N19), .O(N212) );
inv1 gate8( .a(N22), .O(N216) );
inv1 gate9( .a(N25), .O(N220) );
inv1 gate10( .a(N28), .O(N225) );
inv1 gate11( .a(N31), .O(N229) );
inv1 gate12( .a(N34), .O(N232) );
inv1 gate13( .a(N37), .O(N235) );
inv1 gate14( .a(N40), .O(N239) );
inv1 gate15( .a(N43), .O(N243) );
inv1 gate16( .a(N46), .O(N247) );
nand2 gate17( .a(N63), .b(N88), .O(N251) );
nand2 gate18( .a(N66), .b(N91), .O(N252) );
inv1 gate19( .a(N72), .O(N253) );
inv1 gate20( .a(N72), .O(N256) );
buf1 gate21( .a(N69), .O(N257) );
buf1 gate22( .a(N69), .O(N260) );
inv1 gate23( .a(N76), .O(N263) );
inv1 gate24( .a(N79), .O(N266) );
inv1 gate25( .a(N82), .O(N269) );
inv1 gate26( .a(N85), .O(N272) );
inv1 gate27( .a(N104), .O(N275) );
inv1 gate28( .a(N104), .O(N276) );
inv1 gate29( .a(N88), .O(N277) );
inv1 gate30( .a(N91), .O(N280) );
buf1 gate31( .a(N94), .O(N283) );
inv1 gate32( .a(N94), .O(N290) );
buf1 gate33( .a(N94), .O(N297) );
inv1 gate34( .a(N94), .O(N300) );
buf1 gate35( .a(N99), .O(N303) );
inv1 gate36( .a(N99), .O(N306) );
inv1 gate37( .a(N99), .O(N313) );
buf1 gate38( .a(N104), .O(N316) );
inv1 gate39( .a(N104), .O(N319) );
buf1 gate40( .a(N104), .O(N326) );
buf1 gate41( .a(N104), .O(N331) );
inv1 gate42( .a(N104), .O(N338) );
buf1 gate43( .a(N1), .O(N343) );
buf1 gate44( .a(N4), .O(N346) );
buf1 gate45( .a(N7), .O(N349) );
buf1 gate46( .a(N10), .O(N352) );
buf1 gate47( .a(N13), .O(N355) );
buf1 gate48( .a(N16), .O(N358) );
buf1 gate49( .a(N19), .O(N361) );
buf1 gate50( .a(N22), .O(N364) );
buf1 gate51( .a(N25), .O(N367) );
buf1 gate52( .a(N28), .O(N370) );
buf1 gate53( .a(N31), .O(N373) );
buf1 gate54( .a(N34), .O(N376) );
buf1 gate55( .a(N37), .O(N379) );
buf1 gate56( .a(N40), .O(N382) );
buf1 gate57( .a(N43), .O(N385) );
buf1 gate58( .a(N46), .O(N388) );
inv1 gate59( .a(N343), .O(N534) );
inv1 gate60( .a(N346), .O(N535) );
inv1 gate61( .a(N349), .O(N536) );
inv1 gate62( .a(N352), .O(N537) );
inv1 gate63( .a(N355), .O(N538) );
inv1 gate64( .a(N358), .O(N539) );
inv1 gate65( .a(N361), .O(N540) );
inv1 gate66( .a(N364), .O(N541) );
inv1 gate67( .a(N367), .O(N542) );
inv1 gate68( .a(N370), .O(N543) );
inv1 gate69( .a(N373), .O(N544) );
inv1 gate70( .a(N376), .O(N545) );
inv1 gate71( .a(N379), .O(N546) );
inv1 gate72( .a(N382), .O(N547) );
inv1 gate73( .a(N385), .O(N548) );
inv1 gate74( .a(N388), .O(N549) );

  xor2  gate1427(.a(N331), .b(N306), .O(gate75inter0));
  nand2 gate1428(.a(gate75inter0), .b(s_78), .O(gate75inter1));
  and2  gate1429(.a(N331), .b(N306), .O(gate75inter2));
  inv1  gate1430(.a(s_78), .O(gate75inter3));
  inv1  gate1431(.a(s_79), .O(gate75inter4));
  nand2 gate1432(.a(gate75inter4), .b(gate75inter3), .O(gate75inter5));
  nor2  gate1433(.a(gate75inter5), .b(gate75inter2), .O(gate75inter6));
  inv1  gate1434(.a(N306), .O(gate75inter7));
  inv1  gate1435(.a(N331), .O(gate75inter8));
  nand2 gate1436(.a(gate75inter8), .b(gate75inter7), .O(gate75inter9));
  nand2 gate1437(.a(s_79), .b(gate75inter3), .O(gate75inter10));
  nor2  gate1438(.a(gate75inter10), .b(gate75inter9), .O(gate75inter11));
  nor2  gate1439(.a(gate75inter11), .b(gate75inter6), .O(gate75inter12));
  nand2 gate1440(.a(gate75inter12), .b(gate75inter1), .O(N550));
nand2 gate76( .a(N306), .b(N331), .O(N551) );

  xor2  gate1833(.a(N331), .b(N306), .O(gate77inter0));
  nand2 gate1834(.a(gate77inter0), .b(s_136), .O(gate77inter1));
  and2  gate1835(.a(N331), .b(N306), .O(gate77inter2));
  inv1  gate1836(.a(s_136), .O(gate77inter3));
  inv1  gate1837(.a(s_137), .O(gate77inter4));
  nand2 gate1838(.a(gate77inter4), .b(gate77inter3), .O(gate77inter5));
  nor2  gate1839(.a(gate77inter5), .b(gate77inter2), .O(gate77inter6));
  inv1  gate1840(.a(N306), .O(gate77inter7));
  inv1  gate1841(.a(N331), .O(gate77inter8));
  nand2 gate1842(.a(gate77inter8), .b(gate77inter7), .O(gate77inter9));
  nand2 gate1843(.a(s_137), .b(gate77inter3), .O(gate77inter10));
  nor2  gate1844(.a(gate77inter10), .b(gate77inter9), .O(gate77inter11));
  nor2  gate1845(.a(gate77inter11), .b(gate77inter6), .O(gate77inter12));
  nand2 gate1846(.a(gate77inter12), .b(gate77inter1), .O(N552));
nand2 gate78( .a(N306), .b(N331), .O(N553) );

  xor2  gate1469(.a(N331), .b(N306), .O(gate79inter0));
  nand2 gate1470(.a(gate79inter0), .b(s_84), .O(gate79inter1));
  and2  gate1471(.a(N331), .b(N306), .O(gate79inter2));
  inv1  gate1472(.a(s_84), .O(gate79inter3));
  inv1  gate1473(.a(s_85), .O(gate79inter4));
  nand2 gate1474(.a(gate79inter4), .b(gate79inter3), .O(gate79inter5));
  nor2  gate1475(.a(gate79inter5), .b(gate79inter2), .O(gate79inter6));
  inv1  gate1476(.a(N306), .O(gate79inter7));
  inv1  gate1477(.a(N331), .O(gate79inter8));
  nand2 gate1478(.a(gate79inter8), .b(gate79inter7), .O(gate79inter9));
  nand2 gate1479(.a(s_85), .b(gate79inter3), .O(gate79inter10));
  nor2  gate1480(.a(gate79inter10), .b(gate79inter9), .O(gate79inter11));
  nor2  gate1481(.a(gate79inter11), .b(gate79inter6), .O(gate79inter12));
  nand2 gate1482(.a(gate79inter12), .b(gate79inter1), .O(N554));
nand2 gate80( .a(N306), .b(N331), .O(N555) );
buf1 gate81( .a(N190), .O(N556) );
buf1 gate82( .a(N194), .O(N559) );
buf1 gate83( .a(N206), .O(N562) );
buf1 gate84( .a(N209), .O(N565) );
buf1 gate85( .a(N225), .O(N568) );
buf1 gate86( .a(N243), .O(N571) );
and2 gate87( .a(N63), .b(N319), .O(N574) );
buf1 gate88( .a(N220), .O(N577) );
buf1 gate89( .a(N229), .O(N580) );
buf1 gate90( .a(N232), .O(N583) );
and2 gate91( .a(N66), .b(N319), .O(N586) );
buf1 gate92( .a(N239), .O(N589) );
and3 gate93( .a(N49), .b(N253), .c(N319), .O(N592) );
buf1 gate94( .a(N247), .O(N595) );
buf1 gate95( .a(N239), .O(N598) );
nand2 gate96( .a(N326), .b(N277), .O(N601) );
nand2 gate97( .a(N326), .b(N280), .O(N602) );

  xor2  gate1931(.a(N72), .b(N260), .O(gate98inter0));
  nand2 gate1932(.a(gate98inter0), .b(s_150), .O(gate98inter1));
  and2  gate1933(.a(N72), .b(N260), .O(gate98inter2));
  inv1  gate1934(.a(s_150), .O(gate98inter3));
  inv1  gate1935(.a(s_151), .O(gate98inter4));
  nand2 gate1936(.a(gate98inter4), .b(gate98inter3), .O(gate98inter5));
  nor2  gate1937(.a(gate98inter5), .b(gate98inter2), .O(gate98inter6));
  inv1  gate1938(.a(N260), .O(gate98inter7));
  inv1  gate1939(.a(N72), .O(gate98inter8));
  nand2 gate1940(.a(gate98inter8), .b(gate98inter7), .O(gate98inter9));
  nand2 gate1941(.a(s_151), .b(gate98inter3), .O(gate98inter10));
  nor2  gate1942(.a(gate98inter10), .b(gate98inter9), .O(gate98inter11));
  nor2  gate1943(.a(gate98inter11), .b(gate98inter6), .O(gate98inter12));
  nand2 gate1944(.a(gate98inter12), .b(gate98inter1), .O(N603));
nand2 gate99( .a(N260), .b(N300), .O(N608) );

  xor2  gate2239(.a(N300), .b(N256), .O(gate100inter0));
  nand2 gate2240(.a(gate100inter0), .b(s_194), .O(gate100inter1));
  and2  gate2241(.a(N300), .b(N256), .O(gate100inter2));
  inv1  gate2242(.a(s_194), .O(gate100inter3));
  inv1  gate2243(.a(s_195), .O(gate100inter4));
  nand2 gate2244(.a(gate100inter4), .b(gate100inter3), .O(gate100inter5));
  nor2  gate2245(.a(gate100inter5), .b(gate100inter2), .O(gate100inter6));
  inv1  gate2246(.a(N256), .O(gate100inter7));
  inv1  gate2247(.a(N300), .O(gate100inter8));
  nand2 gate2248(.a(gate100inter8), .b(gate100inter7), .O(gate100inter9));
  nand2 gate2249(.a(s_195), .b(gate100inter3), .O(gate100inter10));
  nor2  gate2250(.a(gate100inter10), .b(gate100inter9), .O(gate100inter11));
  nor2  gate2251(.a(gate100inter11), .b(gate100inter6), .O(gate100inter12));
  nand2 gate2252(.a(gate100inter12), .b(gate100inter1), .O(N612));
buf1 gate101( .a(N201), .O(N616) );
buf1 gate102( .a(N216), .O(N619) );
buf1 gate103( .a(N220), .O(N622) );
buf1 gate104( .a(N239), .O(N625) );
buf1 gate105( .a(N190), .O(N628) );
buf1 gate106( .a(N190), .O(N631) );
buf1 gate107( .a(N194), .O(N634) );
buf1 gate108( .a(N229), .O(N637) );
buf1 gate109( .a(N197), .O(N640) );
and3 gate110( .a(N56), .b(N257), .c(N319), .O(N643) );
buf1 gate111( .a(N232), .O(N646) );
buf1 gate112( .a(N201), .O(N649) );
buf1 gate113( .a(N235), .O(N652) );
and3 gate114( .a(N60), .b(N257), .c(N319), .O(N655) );
buf1 gate115( .a(N263), .O(N658) );
buf1 gate116( .a(N263), .O(N661) );
buf1 gate117( .a(N266), .O(N664) );
buf1 gate118( .a(N266), .O(N667) );
buf1 gate119( .a(N269), .O(N670) );
buf1 gate120( .a(N269), .O(N673) );
buf1 gate121( .a(N272), .O(N676) );
buf1 gate122( .a(N272), .O(N679) );
and2 gate123( .a(N251), .b(N316), .O(N682) );
and2 gate124( .a(N252), .b(N316), .O(N685) );
buf1 gate125( .a(N197), .O(N688) );
buf1 gate126( .a(N197), .O(N691) );
buf1 gate127( .a(N212), .O(N694) );
buf1 gate128( .a(N212), .O(N697) );
buf1 gate129( .a(N247), .O(N700) );
buf1 gate130( .a(N247), .O(N703) );
buf1 gate131( .a(N235), .O(N706) );
buf1 gate132( .a(N235), .O(N709) );
buf1 gate133( .a(N201), .O(N712) );
buf1 gate134( .a(N201), .O(N715) );
buf1 gate135( .a(N206), .O(N718) );
buf1 gate136( .a(N216), .O(N721) );
and3 gate137( .a(N53), .b(N253), .c(N319), .O(N724) );
buf1 gate138( .a(N243), .O(N727) );
buf1 gate139( .a(N220), .O(N730) );
buf1 gate140( .a(N220), .O(N733) );
buf1 gate141( .a(N209), .O(N736) );
buf1 gate142( .a(N216), .O(N739) );
buf1 gate143( .a(N225), .O(N742) );
buf1 gate144( .a(N243), .O(N745) );
buf1 gate145( .a(N212), .O(N748) );
buf1 gate146( .a(N225), .O(N751) );
inv1 gate147( .a(N682), .O(N886) );
inv1 gate148( .a(N685), .O(N887) );
inv1 gate149( .a(N616), .O(N888) );
inv1 gate150( .a(N619), .O(N889) );
inv1 gate151( .a(N622), .O(N890) );
inv1 gate152( .a(N625), .O(N891) );
inv1 gate153( .a(N631), .O(N892) );
inv1 gate154( .a(N643), .O(N893) );
inv1 gate155( .a(N649), .O(N894) );
inv1 gate156( .a(N652), .O(N895) );
inv1 gate157( .a(N655), .O(N896) );
and2 gate158( .a(N49), .b(N612), .O(N897) );
and2 gate159( .a(N56), .b(N608), .O(N898) );
nand2 gate160( .a(N53), .b(N612), .O(N899) );

  xor2  gate965(.a(N608), .b(N60), .O(gate161inter0));
  nand2 gate966(.a(gate161inter0), .b(s_12), .O(gate161inter1));
  and2  gate967(.a(N608), .b(N60), .O(gate161inter2));
  inv1  gate968(.a(s_12), .O(gate161inter3));
  inv1  gate969(.a(s_13), .O(gate161inter4));
  nand2 gate970(.a(gate161inter4), .b(gate161inter3), .O(gate161inter5));
  nor2  gate971(.a(gate161inter5), .b(gate161inter2), .O(gate161inter6));
  inv1  gate972(.a(N60), .O(gate161inter7));
  inv1  gate973(.a(N608), .O(gate161inter8));
  nand2 gate974(.a(gate161inter8), .b(gate161inter7), .O(gate161inter9));
  nand2 gate975(.a(s_13), .b(gate161inter3), .O(gate161inter10));
  nor2  gate976(.a(gate161inter10), .b(gate161inter9), .O(gate161inter11));
  nor2  gate977(.a(gate161inter11), .b(gate161inter6), .O(gate161inter12));
  nand2 gate978(.a(gate161inter12), .b(gate161inter1), .O(N903));

  xor2  gate2113(.a(N612), .b(N49), .O(gate162inter0));
  nand2 gate2114(.a(gate162inter0), .b(s_176), .O(gate162inter1));
  and2  gate2115(.a(N612), .b(N49), .O(gate162inter2));
  inv1  gate2116(.a(s_176), .O(gate162inter3));
  inv1  gate2117(.a(s_177), .O(gate162inter4));
  nand2 gate2118(.a(gate162inter4), .b(gate162inter3), .O(gate162inter5));
  nor2  gate2119(.a(gate162inter5), .b(gate162inter2), .O(gate162inter6));
  inv1  gate2120(.a(N49), .O(gate162inter7));
  inv1  gate2121(.a(N612), .O(gate162inter8));
  nand2 gate2122(.a(gate162inter8), .b(gate162inter7), .O(gate162inter9));
  nand2 gate2123(.a(s_177), .b(gate162inter3), .O(gate162inter10));
  nor2  gate2124(.a(gate162inter10), .b(gate162inter9), .O(gate162inter11));
  nor2  gate2125(.a(gate162inter11), .b(gate162inter6), .O(gate162inter12));
  nand2 gate2126(.a(gate162inter12), .b(gate162inter1), .O(N907));
nand2 gate163( .a(N56), .b(N608), .O(N910) );
inv1 gate164( .a(N661), .O(N913) );
inv1 gate165( .a(N658), .O(N914) );
inv1 gate166( .a(N667), .O(N915) );
inv1 gate167( .a(N664), .O(N916) );
inv1 gate168( .a(N673), .O(N917) );
inv1 gate169( .a(N670), .O(N918) );
inv1 gate170( .a(N679), .O(N919) );
inv1 gate171( .a(N676), .O(N920) );
nand4 gate172( .a(N277), .b(N297), .c(N326), .d(N603), .O(N921) );
nand4 gate173( .a(N280), .b(N297), .c(N326), .d(N603), .O(N922) );
nand3 gate174( .a(N303), .b(N338), .c(N603), .O(N923) );
and3 gate175( .a(N303), .b(N338), .c(N603), .O(N926) );
buf1 gate176( .a(N556), .O(N935) );
inv1 gate177( .a(N688), .O(N938) );
buf1 gate178( .a(N556), .O(N939) );
inv1 gate179( .a(N691), .O(N942) );
buf1 gate180( .a(N562), .O(N943) );
inv1 gate181( .a(N694), .O(N946) );
buf1 gate182( .a(N562), .O(N947) );
inv1 gate183( .a(N697), .O(N950) );
buf1 gate184( .a(N568), .O(N951) );
inv1 gate185( .a(N700), .O(N954) );
buf1 gate186( .a(N568), .O(N955) );
inv1 gate187( .a(N703), .O(N958) );
buf1 gate188( .a(N574), .O(N959) );
buf1 gate189( .a(N574), .O(N962) );
buf1 gate190( .a(N580), .O(N965) );
inv1 gate191( .a(N706), .O(N968) );
buf1 gate192( .a(N580), .O(N969) );
inv1 gate193( .a(N709), .O(N972) );
buf1 gate194( .a(N586), .O(N973) );
inv1 gate195( .a(N712), .O(N976) );
buf1 gate196( .a(N586), .O(N977) );
inv1 gate197( .a(N715), .O(N980) );
buf1 gate198( .a(N592), .O(N981) );
inv1 gate199( .a(N628), .O(N984) );
buf1 gate200( .a(N592), .O(N985) );
inv1 gate201( .a(N718), .O(N988) );
inv1 gate202( .a(N721), .O(N989) );
inv1 gate203( .a(N634), .O(N990) );
inv1 gate204( .a(N724), .O(N991) );
inv1 gate205( .a(N727), .O(N992) );
inv1 gate206( .a(N637), .O(N993) );
buf1 gate207( .a(N595), .O(N994) );
inv1 gate208( .a(N730), .O(N997) );
buf1 gate209( .a(N595), .O(N998) );
inv1 gate210( .a(N733), .O(N1001) );
inv1 gate211( .a(N736), .O(N1002) );
inv1 gate212( .a(N739), .O(N1003) );
inv1 gate213( .a(N640), .O(N1004) );
inv1 gate214( .a(N742), .O(N1005) );
inv1 gate215( .a(N745), .O(N1006) );
inv1 gate216( .a(N646), .O(N1007) );
inv1 gate217( .a(N748), .O(N1008) );
inv1 gate218( .a(N751), .O(N1009) );
buf1 gate219( .a(N559), .O(N1010) );
buf1 gate220( .a(N559), .O(N1013) );
buf1 gate221( .a(N565), .O(N1016) );
buf1 gate222( .a(N565), .O(N1019) );
buf1 gate223( .a(N571), .O(N1022) );
buf1 gate224( .a(N571), .O(N1025) );
buf1 gate225( .a(N577), .O(N1028) );
buf1 gate226( .a(N577), .O(N1031) );
buf1 gate227( .a(N583), .O(N1034) );
buf1 gate228( .a(N583), .O(N1037) );
buf1 gate229( .a(N589), .O(N1040) );
buf1 gate230( .a(N589), .O(N1043) );
buf1 gate231( .a(N598), .O(N1046) );
buf1 gate232( .a(N598), .O(N1049) );
nand2 gate233( .a(N619), .b(N888), .O(N1054) );

  xor2  gate1413(.a(N889), .b(N616), .O(gate234inter0));
  nand2 gate1414(.a(gate234inter0), .b(s_76), .O(gate234inter1));
  and2  gate1415(.a(N889), .b(N616), .O(gate234inter2));
  inv1  gate1416(.a(s_76), .O(gate234inter3));
  inv1  gate1417(.a(s_77), .O(gate234inter4));
  nand2 gate1418(.a(gate234inter4), .b(gate234inter3), .O(gate234inter5));
  nor2  gate1419(.a(gate234inter5), .b(gate234inter2), .O(gate234inter6));
  inv1  gate1420(.a(N616), .O(gate234inter7));
  inv1  gate1421(.a(N889), .O(gate234inter8));
  nand2 gate1422(.a(gate234inter8), .b(gate234inter7), .O(gate234inter9));
  nand2 gate1423(.a(s_77), .b(gate234inter3), .O(gate234inter10));
  nor2  gate1424(.a(gate234inter10), .b(gate234inter9), .O(gate234inter11));
  nor2  gate1425(.a(gate234inter11), .b(gate234inter6), .O(gate234inter12));
  nand2 gate1426(.a(gate234inter12), .b(gate234inter1), .O(N1055));

  xor2  gate1847(.a(N890), .b(N625), .O(gate235inter0));
  nand2 gate1848(.a(gate235inter0), .b(s_138), .O(gate235inter1));
  and2  gate1849(.a(N890), .b(N625), .O(gate235inter2));
  inv1  gate1850(.a(s_138), .O(gate235inter3));
  inv1  gate1851(.a(s_139), .O(gate235inter4));
  nand2 gate1852(.a(gate235inter4), .b(gate235inter3), .O(gate235inter5));
  nor2  gate1853(.a(gate235inter5), .b(gate235inter2), .O(gate235inter6));
  inv1  gate1854(.a(N625), .O(gate235inter7));
  inv1  gate1855(.a(N890), .O(gate235inter8));
  nand2 gate1856(.a(gate235inter8), .b(gate235inter7), .O(gate235inter9));
  nand2 gate1857(.a(s_139), .b(gate235inter3), .O(gate235inter10));
  nor2  gate1858(.a(gate235inter10), .b(gate235inter9), .O(gate235inter11));
  nor2  gate1859(.a(gate235inter11), .b(gate235inter6), .O(gate235inter12));
  nand2 gate1860(.a(gate235inter12), .b(gate235inter1), .O(N1063));
nand2 gate236( .a(N622), .b(N891), .O(N1064) );
nand2 gate237( .a(N655), .b(N895), .O(N1067) );
nand2 gate238( .a(N652), .b(N896), .O(N1068) );
nand2 gate239( .a(N721), .b(N988), .O(N1119) );
nand2 gate240( .a(N718), .b(N989), .O(N1120) );
nand2 gate241( .a(N727), .b(N991), .O(N1121) );
nand2 gate242( .a(N724), .b(N992), .O(N1122) );
nand2 gate243( .a(N739), .b(N1002), .O(N1128) );
nand2 gate244( .a(N736), .b(N1003), .O(N1129) );

  xor2  gate1917(.a(N1005), .b(N745), .O(gate245inter0));
  nand2 gate1918(.a(gate245inter0), .b(s_148), .O(gate245inter1));
  and2  gate1919(.a(N1005), .b(N745), .O(gate245inter2));
  inv1  gate1920(.a(s_148), .O(gate245inter3));
  inv1  gate1921(.a(s_149), .O(gate245inter4));
  nand2 gate1922(.a(gate245inter4), .b(gate245inter3), .O(gate245inter5));
  nor2  gate1923(.a(gate245inter5), .b(gate245inter2), .O(gate245inter6));
  inv1  gate1924(.a(N745), .O(gate245inter7));
  inv1  gate1925(.a(N1005), .O(gate245inter8));
  nand2 gate1926(.a(gate245inter8), .b(gate245inter7), .O(gate245inter9));
  nand2 gate1927(.a(s_149), .b(gate245inter3), .O(gate245inter10));
  nor2  gate1928(.a(gate245inter10), .b(gate245inter9), .O(gate245inter11));
  nor2  gate1929(.a(gate245inter11), .b(gate245inter6), .O(gate245inter12));
  nand2 gate1930(.a(gate245inter12), .b(gate245inter1), .O(N1130));
nand2 gate246( .a(N742), .b(N1006), .O(N1131) );

  xor2  gate2043(.a(N1008), .b(N751), .O(gate247inter0));
  nand2 gate2044(.a(gate247inter0), .b(s_166), .O(gate247inter1));
  and2  gate2045(.a(N1008), .b(N751), .O(gate247inter2));
  inv1  gate2046(.a(s_166), .O(gate247inter3));
  inv1  gate2047(.a(s_167), .O(gate247inter4));
  nand2 gate2048(.a(gate247inter4), .b(gate247inter3), .O(gate247inter5));
  nor2  gate2049(.a(gate247inter5), .b(gate247inter2), .O(gate247inter6));
  inv1  gate2050(.a(N751), .O(gate247inter7));
  inv1  gate2051(.a(N1008), .O(gate247inter8));
  nand2 gate2052(.a(gate247inter8), .b(gate247inter7), .O(gate247inter9));
  nand2 gate2053(.a(s_167), .b(gate247inter3), .O(gate247inter10));
  nor2  gate2054(.a(gate247inter10), .b(gate247inter9), .O(gate247inter11));
  nor2  gate2055(.a(gate247inter11), .b(gate247inter6), .O(gate247inter12));
  nand2 gate2056(.a(gate247inter12), .b(gate247inter1), .O(N1132));

  xor2  gate1021(.a(N1009), .b(N748), .O(gate248inter0));
  nand2 gate1022(.a(gate248inter0), .b(s_20), .O(gate248inter1));
  and2  gate1023(.a(N1009), .b(N748), .O(gate248inter2));
  inv1  gate1024(.a(s_20), .O(gate248inter3));
  inv1  gate1025(.a(s_21), .O(gate248inter4));
  nand2 gate1026(.a(gate248inter4), .b(gate248inter3), .O(gate248inter5));
  nor2  gate1027(.a(gate248inter5), .b(gate248inter2), .O(gate248inter6));
  inv1  gate1028(.a(N748), .O(gate248inter7));
  inv1  gate1029(.a(N1009), .O(gate248inter8));
  nand2 gate1030(.a(gate248inter8), .b(gate248inter7), .O(gate248inter9));
  nand2 gate1031(.a(s_21), .b(gate248inter3), .O(gate248inter10));
  nor2  gate1032(.a(gate248inter10), .b(gate248inter9), .O(gate248inter11));
  nor2  gate1033(.a(gate248inter11), .b(gate248inter6), .O(gate248inter12));
  nand2 gate1034(.a(gate248inter12), .b(gate248inter1), .O(N1133));
inv1 gate249( .a(N939), .O(N1148) );
inv1 gate250( .a(N935), .O(N1149) );

  xor2  gate993(.a(N1055), .b(N1054), .O(gate251inter0));
  nand2 gate994(.a(gate251inter0), .b(s_16), .O(gate251inter1));
  and2  gate995(.a(N1055), .b(N1054), .O(gate251inter2));
  inv1  gate996(.a(s_16), .O(gate251inter3));
  inv1  gate997(.a(s_17), .O(gate251inter4));
  nand2 gate998(.a(gate251inter4), .b(gate251inter3), .O(gate251inter5));
  nor2  gate999(.a(gate251inter5), .b(gate251inter2), .O(gate251inter6));
  inv1  gate1000(.a(N1054), .O(gate251inter7));
  inv1  gate1001(.a(N1055), .O(gate251inter8));
  nand2 gate1002(.a(gate251inter8), .b(gate251inter7), .O(gate251inter9));
  nand2 gate1003(.a(s_17), .b(gate251inter3), .O(gate251inter10));
  nor2  gate1004(.a(gate251inter10), .b(gate251inter9), .O(gate251inter11));
  nor2  gate1005(.a(gate251inter11), .b(gate251inter6), .O(gate251inter12));
  nand2 gate1006(.a(gate251inter12), .b(gate251inter1), .O(N1150));
inv1 gate252( .a(N943), .O(N1151) );
inv1 gate253( .a(N947), .O(N1152) );
inv1 gate254( .a(N955), .O(N1153) );
inv1 gate255( .a(N951), .O(N1154) );
inv1 gate256( .a(N962), .O(N1155) );
inv1 gate257( .a(N969), .O(N1156) );
inv1 gate258( .a(N977), .O(N1157) );

  xor2  gate1525(.a(N1064), .b(N1063), .O(gate259inter0));
  nand2 gate1526(.a(gate259inter0), .b(s_92), .O(gate259inter1));
  and2  gate1527(.a(N1064), .b(N1063), .O(gate259inter2));
  inv1  gate1528(.a(s_92), .O(gate259inter3));
  inv1  gate1529(.a(s_93), .O(gate259inter4));
  nand2 gate1530(.a(gate259inter4), .b(gate259inter3), .O(gate259inter5));
  nor2  gate1531(.a(gate259inter5), .b(gate259inter2), .O(gate259inter6));
  inv1  gate1532(.a(N1063), .O(gate259inter7));
  inv1  gate1533(.a(N1064), .O(gate259inter8));
  nand2 gate1534(.a(gate259inter8), .b(gate259inter7), .O(gate259inter9));
  nand2 gate1535(.a(s_93), .b(gate259inter3), .O(gate259inter10));
  nor2  gate1536(.a(gate259inter10), .b(gate259inter9), .O(gate259inter11));
  nor2  gate1537(.a(gate259inter11), .b(gate259inter6), .O(gate259inter12));
  nand2 gate1538(.a(gate259inter12), .b(gate259inter1), .O(N1158));
inv1 gate260( .a(N985), .O(N1159) );
nand2 gate261( .a(N985), .b(N892), .O(N1160) );
inv1 gate262( .a(N998), .O(N1161) );
nand2 gate263( .a(N1067), .b(N1068), .O(N1162) );
inv1 gate264( .a(N899), .O(N1163) );
buf1 gate265( .a(N899), .O(N1164) );
inv1 gate266( .a(N903), .O(N1167) );
buf1 gate267( .a(N903), .O(N1168) );
nand2 gate268( .a(N921), .b(N923), .O(N1171) );

  xor2  gate1581(.a(N923), .b(N922), .O(gate269inter0));
  nand2 gate1582(.a(gate269inter0), .b(s_100), .O(gate269inter1));
  and2  gate1583(.a(N923), .b(N922), .O(gate269inter2));
  inv1  gate1584(.a(s_100), .O(gate269inter3));
  inv1  gate1585(.a(s_101), .O(gate269inter4));
  nand2 gate1586(.a(gate269inter4), .b(gate269inter3), .O(gate269inter5));
  nor2  gate1587(.a(gate269inter5), .b(gate269inter2), .O(gate269inter6));
  inv1  gate1588(.a(N922), .O(gate269inter7));
  inv1  gate1589(.a(N923), .O(gate269inter8));
  nand2 gate1590(.a(gate269inter8), .b(gate269inter7), .O(gate269inter9));
  nand2 gate1591(.a(s_101), .b(gate269inter3), .O(gate269inter10));
  nor2  gate1592(.a(gate269inter10), .b(gate269inter9), .O(gate269inter11));
  nor2  gate1593(.a(gate269inter11), .b(gate269inter6), .O(gate269inter12));
  nand2 gate1594(.a(gate269inter12), .b(gate269inter1), .O(N1188));
inv1 gate270( .a(N1010), .O(N1205) );
nand2 gate271( .a(N1010), .b(N938), .O(N1206) );
inv1 gate272( .a(N1013), .O(N1207) );

  xor2  gate1203(.a(N942), .b(N1013), .O(gate273inter0));
  nand2 gate1204(.a(gate273inter0), .b(s_46), .O(gate273inter1));
  and2  gate1205(.a(N942), .b(N1013), .O(gate273inter2));
  inv1  gate1206(.a(s_46), .O(gate273inter3));
  inv1  gate1207(.a(s_47), .O(gate273inter4));
  nand2 gate1208(.a(gate273inter4), .b(gate273inter3), .O(gate273inter5));
  nor2  gate1209(.a(gate273inter5), .b(gate273inter2), .O(gate273inter6));
  inv1  gate1210(.a(N1013), .O(gate273inter7));
  inv1  gate1211(.a(N942), .O(gate273inter8));
  nand2 gate1212(.a(gate273inter8), .b(gate273inter7), .O(gate273inter9));
  nand2 gate1213(.a(s_47), .b(gate273inter3), .O(gate273inter10));
  nor2  gate1214(.a(gate273inter10), .b(gate273inter9), .O(gate273inter11));
  nor2  gate1215(.a(gate273inter11), .b(gate273inter6), .O(gate273inter12));
  nand2 gate1216(.a(gate273inter12), .b(gate273inter1), .O(N1208));
inv1 gate274( .a(N1016), .O(N1209) );
nand2 gate275( .a(N1016), .b(N946), .O(N1210) );
inv1 gate276( .a(N1019), .O(N1211) );

  xor2  gate951(.a(N950), .b(N1019), .O(gate277inter0));
  nand2 gate952(.a(gate277inter0), .b(s_10), .O(gate277inter1));
  and2  gate953(.a(N950), .b(N1019), .O(gate277inter2));
  inv1  gate954(.a(s_10), .O(gate277inter3));
  inv1  gate955(.a(s_11), .O(gate277inter4));
  nand2 gate956(.a(gate277inter4), .b(gate277inter3), .O(gate277inter5));
  nor2  gate957(.a(gate277inter5), .b(gate277inter2), .O(gate277inter6));
  inv1  gate958(.a(N1019), .O(gate277inter7));
  inv1  gate959(.a(N950), .O(gate277inter8));
  nand2 gate960(.a(gate277inter8), .b(gate277inter7), .O(gate277inter9));
  nand2 gate961(.a(s_11), .b(gate277inter3), .O(gate277inter10));
  nor2  gate962(.a(gate277inter10), .b(gate277inter9), .O(gate277inter11));
  nor2  gate963(.a(gate277inter11), .b(gate277inter6), .O(gate277inter12));
  nand2 gate964(.a(gate277inter12), .b(gate277inter1), .O(N1212));
inv1 gate278( .a(N1022), .O(N1213) );
nand2 gate279( .a(N1022), .b(N954), .O(N1214) );
inv1 gate280( .a(N1025), .O(N1215) );

  xor2  gate2337(.a(N958), .b(N1025), .O(gate281inter0));
  nand2 gate2338(.a(gate281inter0), .b(s_208), .O(gate281inter1));
  and2  gate2339(.a(N958), .b(N1025), .O(gate281inter2));
  inv1  gate2340(.a(s_208), .O(gate281inter3));
  inv1  gate2341(.a(s_209), .O(gate281inter4));
  nand2 gate2342(.a(gate281inter4), .b(gate281inter3), .O(gate281inter5));
  nor2  gate2343(.a(gate281inter5), .b(gate281inter2), .O(gate281inter6));
  inv1  gate2344(.a(N1025), .O(gate281inter7));
  inv1  gate2345(.a(N958), .O(gate281inter8));
  nand2 gate2346(.a(gate281inter8), .b(gate281inter7), .O(gate281inter9));
  nand2 gate2347(.a(s_209), .b(gate281inter3), .O(gate281inter10));
  nor2  gate2348(.a(gate281inter10), .b(gate281inter9), .O(gate281inter11));
  nor2  gate2349(.a(gate281inter11), .b(gate281inter6), .O(gate281inter12));
  nand2 gate2350(.a(gate281inter12), .b(gate281inter1), .O(N1216));
inv1 gate282( .a(N1028), .O(N1217) );
inv1 gate283( .a(N959), .O(N1218) );
inv1 gate284( .a(N1031), .O(N1219) );
inv1 gate285( .a(N1034), .O(N1220) );

  xor2  gate2323(.a(N968), .b(N1034), .O(gate286inter0));
  nand2 gate2324(.a(gate286inter0), .b(s_206), .O(gate286inter1));
  and2  gate2325(.a(N968), .b(N1034), .O(gate286inter2));
  inv1  gate2326(.a(s_206), .O(gate286inter3));
  inv1  gate2327(.a(s_207), .O(gate286inter4));
  nand2 gate2328(.a(gate286inter4), .b(gate286inter3), .O(gate286inter5));
  nor2  gate2329(.a(gate286inter5), .b(gate286inter2), .O(gate286inter6));
  inv1  gate2330(.a(N1034), .O(gate286inter7));
  inv1  gate2331(.a(N968), .O(gate286inter8));
  nand2 gate2332(.a(gate286inter8), .b(gate286inter7), .O(gate286inter9));
  nand2 gate2333(.a(s_207), .b(gate286inter3), .O(gate286inter10));
  nor2  gate2334(.a(gate286inter10), .b(gate286inter9), .O(gate286inter11));
  nor2  gate2335(.a(gate286inter11), .b(gate286inter6), .O(gate286inter12));
  nand2 gate2336(.a(gate286inter12), .b(gate286inter1), .O(N1221));
inv1 gate287( .a(N965), .O(N1222) );
inv1 gate288( .a(N1037), .O(N1223) );
nand2 gate289( .a(N1037), .b(N972), .O(N1224) );
inv1 gate290( .a(N1040), .O(N1225) );
nand2 gate291( .a(N1040), .b(N976), .O(N1226) );
inv1 gate292( .a(N973), .O(N1227) );
inv1 gate293( .a(N1043), .O(N1228) );
nand2 gate294( .a(N1043), .b(N980), .O(N1229) );
inv1 gate295( .a(N981), .O(N1230) );
nand2 gate296( .a(N981), .b(N984), .O(N1231) );
nand2 gate297( .a(N1119), .b(N1120), .O(N1232) );
nand2 gate298( .a(N1121), .b(N1122), .O(N1235) );
inv1 gate299( .a(N1046), .O(N1238) );

  xor2  gate881(.a(N997), .b(N1046), .O(gate300inter0));
  nand2 gate882(.a(gate300inter0), .b(s_0), .O(gate300inter1));
  and2  gate883(.a(N997), .b(N1046), .O(gate300inter2));
  inv1  gate884(.a(s_0), .O(gate300inter3));
  inv1  gate885(.a(s_1), .O(gate300inter4));
  nand2 gate886(.a(gate300inter4), .b(gate300inter3), .O(gate300inter5));
  nor2  gate887(.a(gate300inter5), .b(gate300inter2), .O(gate300inter6));
  inv1  gate888(.a(N1046), .O(gate300inter7));
  inv1  gate889(.a(N997), .O(gate300inter8));
  nand2 gate890(.a(gate300inter8), .b(gate300inter7), .O(gate300inter9));
  nand2 gate891(.a(s_1), .b(gate300inter3), .O(gate300inter10));
  nor2  gate892(.a(gate300inter10), .b(gate300inter9), .O(gate300inter11));
  nor2  gate893(.a(gate300inter11), .b(gate300inter6), .O(gate300inter12));
  nand2 gate894(.a(gate300inter12), .b(gate300inter1), .O(N1239));
inv1 gate301( .a(N994), .O(N1240) );
inv1 gate302( .a(N1049), .O(N1241) );

  xor2  gate1945(.a(N1001), .b(N1049), .O(gate303inter0));
  nand2 gate1946(.a(gate303inter0), .b(s_152), .O(gate303inter1));
  and2  gate1947(.a(N1001), .b(N1049), .O(gate303inter2));
  inv1  gate1948(.a(s_152), .O(gate303inter3));
  inv1  gate1949(.a(s_153), .O(gate303inter4));
  nand2 gate1950(.a(gate303inter4), .b(gate303inter3), .O(gate303inter5));
  nor2  gate1951(.a(gate303inter5), .b(gate303inter2), .O(gate303inter6));
  inv1  gate1952(.a(N1049), .O(gate303inter7));
  inv1  gate1953(.a(N1001), .O(gate303inter8));
  nand2 gate1954(.a(gate303inter8), .b(gate303inter7), .O(gate303inter9));
  nand2 gate1955(.a(s_153), .b(gate303inter3), .O(gate303inter10));
  nor2  gate1956(.a(gate303inter10), .b(gate303inter9), .O(gate303inter11));
  nor2  gate1957(.a(gate303inter11), .b(gate303inter6), .O(gate303inter12));
  nand2 gate1958(.a(gate303inter12), .b(gate303inter1), .O(N1242));

  xor2  gate1399(.a(N1129), .b(N1128), .O(gate304inter0));
  nand2 gate1400(.a(gate304inter0), .b(s_74), .O(gate304inter1));
  and2  gate1401(.a(N1129), .b(N1128), .O(gate304inter2));
  inv1  gate1402(.a(s_74), .O(gate304inter3));
  inv1  gate1403(.a(s_75), .O(gate304inter4));
  nand2 gate1404(.a(gate304inter4), .b(gate304inter3), .O(gate304inter5));
  nor2  gate1405(.a(gate304inter5), .b(gate304inter2), .O(gate304inter6));
  inv1  gate1406(.a(N1128), .O(gate304inter7));
  inv1  gate1407(.a(N1129), .O(gate304inter8));
  nand2 gate1408(.a(gate304inter8), .b(gate304inter7), .O(gate304inter9));
  nand2 gate1409(.a(s_75), .b(gate304inter3), .O(gate304inter10));
  nor2  gate1410(.a(gate304inter10), .b(gate304inter9), .O(gate304inter11));
  nor2  gate1411(.a(gate304inter11), .b(gate304inter6), .O(gate304inter12));
  nand2 gate1412(.a(gate304inter12), .b(gate304inter1), .O(N1243));

  xor2  gate2267(.a(N1131), .b(N1130), .O(gate305inter0));
  nand2 gate2268(.a(gate305inter0), .b(s_198), .O(gate305inter1));
  and2  gate2269(.a(N1131), .b(N1130), .O(gate305inter2));
  inv1  gate2270(.a(s_198), .O(gate305inter3));
  inv1  gate2271(.a(s_199), .O(gate305inter4));
  nand2 gate2272(.a(gate305inter4), .b(gate305inter3), .O(gate305inter5));
  nor2  gate2273(.a(gate305inter5), .b(gate305inter2), .O(gate305inter6));
  inv1  gate2274(.a(N1130), .O(gate305inter7));
  inv1  gate2275(.a(N1131), .O(gate305inter8));
  nand2 gate2276(.a(gate305inter8), .b(gate305inter7), .O(gate305inter9));
  nand2 gate2277(.a(s_199), .b(gate305inter3), .O(gate305inter10));
  nor2  gate2278(.a(gate305inter10), .b(gate305inter9), .O(gate305inter11));
  nor2  gate2279(.a(gate305inter11), .b(gate305inter6), .O(gate305inter12));
  nand2 gate2280(.a(gate305inter12), .b(gate305inter1), .O(N1246));

  xor2  gate1231(.a(N1133), .b(N1132), .O(gate306inter0));
  nand2 gate1232(.a(gate306inter0), .b(s_50), .O(gate306inter1));
  and2  gate1233(.a(N1133), .b(N1132), .O(gate306inter2));
  inv1  gate1234(.a(s_50), .O(gate306inter3));
  inv1  gate1235(.a(s_51), .O(gate306inter4));
  nand2 gate1236(.a(gate306inter4), .b(gate306inter3), .O(gate306inter5));
  nor2  gate1237(.a(gate306inter5), .b(gate306inter2), .O(gate306inter6));
  inv1  gate1238(.a(N1132), .O(gate306inter7));
  inv1  gate1239(.a(N1133), .O(gate306inter8));
  nand2 gate1240(.a(gate306inter8), .b(gate306inter7), .O(gate306inter9));
  nand2 gate1241(.a(s_51), .b(gate306inter3), .O(gate306inter10));
  nor2  gate1242(.a(gate306inter10), .b(gate306inter9), .O(gate306inter11));
  nor2  gate1243(.a(gate306inter11), .b(gate306inter6), .O(gate306inter12));
  nand2 gate1244(.a(gate306inter12), .b(gate306inter1), .O(N1249));
buf1 gate307( .a(N907), .O(N1252) );
buf1 gate308( .a(N907), .O(N1255) );
buf1 gate309( .a(N910), .O(N1258) );
buf1 gate310( .a(N910), .O(N1261) );
inv1 gate311( .a(N1150), .O(N1264) );
nand2 gate312( .a(N631), .b(N1159), .O(N1267) );
nand2 gate313( .a(N688), .b(N1205), .O(N1309) );

  xor2  gate1049(.a(N1207), .b(N691), .O(gate314inter0));
  nand2 gate1050(.a(gate314inter0), .b(s_24), .O(gate314inter1));
  and2  gate1051(.a(N1207), .b(N691), .O(gate314inter2));
  inv1  gate1052(.a(s_24), .O(gate314inter3));
  inv1  gate1053(.a(s_25), .O(gate314inter4));
  nand2 gate1054(.a(gate314inter4), .b(gate314inter3), .O(gate314inter5));
  nor2  gate1055(.a(gate314inter5), .b(gate314inter2), .O(gate314inter6));
  inv1  gate1056(.a(N691), .O(gate314inter7));
  inv1  gate1057(.a(N1207), .O(gate314inter8));
  nand2 gate1058(.a(gate314inter8), .b(gate314inter7), .O(gate314inter9));
  nand2 gate1059(.a(s_25), .b(gate314inter3), .O(gate314inter10));
  nor2  gate1060(.a(gate314inter10), .b(gate314inter9), .O(gate314inter11));
  nor2  gate1061(.a(gate314inter11), .b(gate314inter6), .O(gate314inter12));
  nand2 gate1062(.a(gate314inter12), .b(gate314inter1), .O(N1310));
nand2 gate315( .a(N694), .b(N1209), .O(N1311) );

  xor2  gate1693(.a(N1211), .b(N697), .O(gate316inter0));
  nand2 gate1694(.a(gate316inter0), .b(s_116), .O(gate316inter1));
  and2  gate1695(.a(N1211), .b(N697), .O(gate316inter2));
  inv1  gate1696(.a(s_116), .O(gate316inter3));
  inv1  gate1697(.a(s_117), .O(gate316inter4));
  nand2 gate1698(.a(gate316inter4), .b(gate316inter3), .O(gate316inter5));
  nor2  gate1699(.a(gate316inter5), .b(gate316inter2), .O(gate316inter6));
  inv1  gate1700(.a(N697), .O(gate316inter7));
  inv1  gate1701(.a(N1211), .O(gate316inter8));
  nand2 gate1702(.a(gate316inter8), .b(gate316inter7), .O(gate316inter9));
  nand2 gate1703(.a(s_117), .b(gate316inter3), .O(gate316inter10));
  nor2  gate1704(.a(gate316inter10), .b(gate316inter9), .O(gate316inter11));
  nor2  gate1705(.a(gate316inter11), .b(gate316inter6), .O(gate316inter12));
  nand2 gate1706(.a(gate316inter12), .b(gate316inter1), .O(N1312));
nand2 gate317( .a(N700), .b(N1213), .O(N1313) );
nand2 gate318( .a(N703), .b(N1215), .O(N1314) );

  xor2  gate1595(.a(N1220), .b(N706), .O(gate319inter0));
  nand2 gate1596(.a(gate319inter0), .b(s_102), .O(gate319inter1));
  and2  gate1597(.a(N1220), .b(N706), .O(gate319inter2));
  inv1  gate1598(.a(s_102), .O(gate319inter3));
  inv1  gate1599(.a(s_103), .O(gate319inter4));
  nand2 gate1600(.a(gate319inter4), .b(gate319inter3), .O(gate319inter5));
  nor2  gate1601(.a(gate319inter5), .b(gate319inter2), .O(gate319inter6));
  inv1  gate1602(.a(N706), .O(gate319inter7));
  inv1  gate1603(.a(N1220), .O(gate319inter8));
  nand2 gate1604(.a(gate319inter8), .b(gate319inter7), .O(gate319inter9));
  nand2 gate1605(.a(s_103), .b(gate319inter3), .O(gate319inter10));
  nor2  gate1606(.a(gate319inter10), .b(gate319inter9), .O(gate319inter11));
  nor2  gate1607(.a(gate319inter11), .b(gate319inter6), .O(gate319inter12));
  nand2 gate1608(.a(gate319inter12), .b(gate319inter1), .O(N1315));
nand2 gate320( .a(N709), .b(N1223), .O(N1316) );
nand2 gate321( .a(N712), .b(N1225), .O(N1317) );

  xor2  gate923(.a(N1228), .b(N715), .O(gate322inter0));
  nand2 gate924(.a(gate322inter0), .b(s_6), .O(gate322inter1));
  and2  gate925(.a(N1228), .b(N715), .O(gate322inter2));
  inv1  gate926(.a(s_6), .O(gate322inter3));
  inv1  gate927(.a(s_7), .O(gate322inter4));
  nand2 gate928(.a(gate322inter4), .b(gate322inter3), .O(gate322inter5));
  nor2  gate929(.a(gate322inter5), .b(gate322inter2), .O(gate322inter6));
  inv1  gate930(.a(N715), .O(gate322inter7));
  inv1  gate931(.a(N1228), .O(gate322inter8));
  nand2 gate932(.a(gate322inter8), .b(gate322inter7), .O(gate322inter9));
  nand2 gate933(.a(s_7), .b(gate322inter3), .O(gate322inter10));
  nor2  gate934(.a(gate322inter10), .b(gate322inter9), .O(gate322inter11));
  nor2  gate935(.a(gate322inter11), .b(gate322inter6), .O(gate322inter12));
  nand2 gate936(.a(gate322inter12), .b(gate322inter1), .O(N1318));
inv1 gate323( .a(N1158), .O(N1319) );
nand2 gate324( .a(N628), .b(N1230), .O(N1322) );

  xor2  gate1455(.a(N1238), .b(N730), .O(gate325inter0));
  nand2 gate1456(.a(gate325inter0), .b(s_82), .O(gate325inter1));
  and2  gate1457(.a(N1238), .b(N730), .O(gate325inter2));
  inv1  gate1458(.a(s_82), .O(gate325inter3));
  inv1  gate1459(.a(s_83), .O(gate325inter4));
  nand2 gate1460(.a(gate325inter4), .b(gate325inter3), .O(gate325inter5));
  nor2  gate1461(.a(gate325inter5), .b(gate325inter2), .O(gate325inter6));
  inv1  gate1462(.a(N730), .O(gate325inter7));
  inv1  gate1463(.a(N1238), .O(gate325inter8));
  nand2 gate1464(.a(gate325inter8), .b(gate325inter7), .O(gate325inter9));
  nand2 gate1465(.a(s_83), .b(gate325inter3), .O(gate325inter10));
  nor2  gate1466(.a(gate325inter10), .b(gate325inter9), .O(gate325inter11));
  nor2  gate1467(.a(gate325inter11), .b(gate325inter6), .O(gate325inter12));
  nand2 gate1468(.a(gate325inter12), .b(gate325inter1), .O(N1327));

  xor2  gate2225(.a(N1241), .b(N733), .O(gate326inter0));
  nand2 gate2226(.a(gate326inter0), .b(s_192), .O(gate326inter1));
  and2  gate2227(.a(N1241), .b(N733), .O(gate326inter2));
  inv1  gate2228(.a(s_192), .O(gate326inter3));
  inv1  gate2229(.a(s_193), .O(gate326inter4));
  nand2 gate2230(.a(gate326inter4), .b(gate326inter3), .O(gate326inter5));
  nor2  gate2231(.a(gate326inter5), .b(gate326inter2), .O(gate326inter6));
  inv1  gate2232(.a(N733), .O(gate326inter7));
  inv1  gate2233(.a(N1241), .O(gate326inter8));
  nand2 gate2234(.a(gate326inter8), .b(gate326inter7), .O(gate326inter9));
  nand2 gate2235(.a(s_193), .b(gate326inter3), .O(gate326inter10));
  nor2  gate2236(.a(gate326inter10), .b(gate326inter9), .O(gate326inter11));
  nor2  gate2237(.a(gate326inter11), .b(gate326inter6), .O(gate326inter12));
  nand2 gate2238(.a(gate326inter12), .b(gate326inter1), .O(N1328));
inv1 gate327( .a(N1162), .O(N1334) );

  xor2  gate1903(.a(N1160), .b(N1267), .O(gate328inter0));
  nand2 gate1904(.a(gate328inter0), .b(s_146), .O(gate328inter1));
  and2  gate1905(.a(N1160), .b(N1267), .O(gate328inter2));
  inv1  gate1906(.a(s_146), .O(gate328inter3));
  inv1  gate1907(.a(s_147), .O(gate328inter4));
  nand2 gate1908(.a(gate328inter4), .b(gate328inter3), .O(gate328inter5));
  nor2  gate1909(.a(gate328inter5), .b(gate328inter2), .O(gate328inter6));
  inv1  gate1910(.a(N1267), .O(gate328inter7));
  inv1  gate1911(.a(N1160), .O(gate328inter8));
  nand2 gate1912(.a(gate328inter8), .b(gate328inter7), .O(gate328inter9));
  nand2 gate1913(.a(s_147), .b(gate328inter3), .O(gate328inter10));
  nor2  gate1914(.a(gate328inter10), .b(gate328inter9), .O(gate328inter11));
  nor2  gate1915(.a(gate328inter11), .b(gate328inter6), .O(gate328inter12));
  nand2 gate1916(.a(gate328inter12), .b(gate328inter1), .O(N1344));
nand2 gate329( .a(N1249), .b(N894), .O(N1345) );
inv1 gate330( .a(N1249), .O(N1346) );
inv1 gate331( .a(N1255), .O(N1348) );
inv1 gate332( .a(N1252), .O(N1349) );
inv1 gate333( .a(N1261), .O(N1350) );
inv1 gate334( .a(N1258), .O(N1351) );
nand2 gate335( .a(N1309), .b(N1206), .O(N1352) );

  xor2  gate1889(.a(N1208), .b(N1310), .O(gate336inter0));
  nand2 gate1890(.a(gate336inter0), .b(s_144), .O(gate336inter1));
  and2  gate1891(.a(N1208), .b(N1310), .O(gate336inter2));
  inv1  gate1892(.a(s_144), .O(gate336inter3));
  inv1  gate1893(.a(s_145), .O(gate336inter4));
  nand2 gate1894(.a(gate336inter4), .b(gate336inter3), .O(gate336inter5));
  nor2  gate1895(.a(gate336inter5), .b(gate336inter2), .O(gate336inter6));
  inv1  gate1896(.a(N1310), .O(gate336inter7));
  inv1  gate1897(.a(N1208), .O(gate336inter8));
  nand2 gate1898(.a(gate336inter8), .b(gate336inter7), .O(gate336inter9));
  nand2 gate1899(.a(s_145), .b(gate336inter3), .O(gate336inter10));
  nor2  gate1900(.a(gate336inter10), .b(gate336inter9), .O(gate336inter11));
  nor2  gate1901(.a(gate336inter11), .b(gate336inter6), .O(gate336inter12));
  nand2 gate1902(.a(gate336inter12), .b(gate336inter1), .O(N1355));
nand2 gate337( .a(N1311), .b(N1210), .O(N1358) );
nand2 gate338( .a(N1312), .b(N1212), .O(N1361) );
nand2 gate339( .a(N1313), .b(N1214), .O(N1364) );
nand2 gate340( .a(N1314), .b(N1216), .O(N1367) );

  xor2  gate2127(.a(N1221), .b(N1315), .O(gate341inter0));
  nand2 gate2128(.a(gate341inter0), .b(s_178), .O(gate341inter1));
  and2  gate2129(.a(N1221), .b(N1315), .O(gate341inter2));
  inv1  gate2130(.a(s_178), .O(gate341inter3));
  inv1  gate2131(.a(s_179), .O(gate341inter4));
  nand2 gate2132(.a(gate341inter4), .b(gate341inter3), .O(gate341inter5));
  nor2  gate2133(.a(gate341inter5), .b(gate341inter2), .O(gate341inter6));
  inv1  gate2134(.a(N1315), .O(gate341inter7));
  inv1  gate2135(.a(N1221), .O(gate341inter8));
  nand2 gate2136(.a(gate341inter8), .b(gate341inter7), .O(gate341inter9));
  nand2 gate2137(.a(s_179), .b(gate341inter3), .O(gate341inter10));
  nor2  gate2138(.a(gate341inter10), .b(gate341inter9), .O(gate341inter11));
  nor2  gate2139(.a(gate341inter11), .b(gate341inter6), .O(gate341inter12));
  nand2 gate2140(.a(gate341inter12), .b(gate341inter1), .O(N1370));
nand2 gate342( .a(N1316), .b(N1224), .O(N1373) );

  xor2  gate2015(.a(N1226), .b(N1317), .O(gate343inter0));
  nand2 gate2016(.a(gate343inter0), .b(s_162), .O(gate343inter1));
  and2  gate2017(.a(N1226), .b(N1317), .O(gate343inter2));
  inv1  gate2018(.a(s_162), .O(gate343inter3));
  inv1  gate2019(.a(s_163), .O(gate343inter4));
  nand2 gate2020(.a(gate343inter4), .b(gate343inter3), .O(gate343inter5));
  nor2  gate2021(.a(gate343inter5), .b(gate343inter2), .O(gate343inter6));
  inv1  gate2022(.a(N1317), .O(gate343inter7));
  inv1  gate2023(.a(N1226), .O(gate343inter8));
  nand2 gate2024(.a(gate343inter8), .b(gate343inter7), .O(gate343inter9));
  nand2 gate2025(.a(s_163), .b(gate343inter3), .O(gate343inter10));
  nor2  gate2026(.a(gate343inter10), .b(gate343inter9), .O(gate343inter11));
  nor2  gate2027(.a(gate343inter11), .b(gate343inter6), .O(gate343inter12));
  nand2 gate2028(.a(gate343inter12), .b(gate343inter1), .O(N1376));

  xor2  gate1749(.a(N1229), .b(N1318), .O(gate344inter0));
  nand2 gate1750(.a(gate344inter0), .b(s_124), .O(gate344inter1));
  and2  gate1751(.a(N1229), .b(N1318), .O(gate344inter2));
  inv1  gate1752(.a(s_124), .O(gate344inter3));
  inv1  gate1753(.a(s_125), .O(gate344inter4));
  nand2 gate1754(.a(gate344inter4), .b(gate344inter3), .O(gate344inter5));
  nor2  gate1755(.a(gate344inter5), .b(gate344inter2), .O(gate344inter6));
  inv1  gate1756(.a(N1318), .O(gate344inter7));
  inv1  gate1757(.a(N1229), .O(gate344inter8));
  nand2 gate1758(.a(gate344inter8), .b(gate344inter7), .O(gate344inter9));
  nand2 gate1759(.a(s_125), .b(gate344inter3), .O(gate344inter10));
  nor2  gate1760(.a(gate344inter10), .b(gate344inter9), .O(gate344inter11));
  nor2  gate1761(.a(gate344inter11), .b(gate344inter6), .O(gate344inter12));
  nand2 gate1762(.a(gate344inter12), .b(gate344inter1), .O(N1379));

  xor2  gate1217(.a(N1231), .b(N1322), .O(gate345inter0));
  nand2 gate1218(.a(gate345inter0), .b(s_48), .O(gate345inter1));
  and2  gate1219(.a(N1231), .b(N1322), .O(gate345inter2));
  inv1  gate1220(.a(s_48), .O(gate345inter3));
  inv1  gate1221(.a(s_49), .O(gate345inter4));
  nand2 gate1222(.a(gate345inter4), .b(gate345inter3), .O(gate345inter5));
  nor2  gate1223(.a(gate345inter5), .b(gate345inter2), .O(gate345inter6));
  inv1  gate1224(.a(N1322), .O(gate345inter7));
  inv1  gate1225(.a(N1231), .O(gate345inter8));
  nand2 gate1226(.a(gate345inter8), .b(gate345inter7), .O(gate345inter9));
  nand2 gate1227(.a(s_49), .b(gate345inter3), .O(gate345inter10));
  nor2  gate1228(.a(gate345inter10), .b(gate345inter9), .O(gate345inter11));
  nor2  gate1229(.a(gate345inter11), .b(gate345inter6), .O(gate345inter12));
  nand2 gate1230(.a(gate345inter12), .b(gate345inter1), .O(N1383));
inv1 gate346( .a(N1232), .O(N1386) );
nand2 gate347( .a(N1232), .b(N990), .O(N1387) );
inv1 gate348( .a(N1235), .O(N1388) );
nand2 gate349( .a(N1235), .b(N993), .O(N1389) );
nand2 gate350( .a(N1327), .b(N1239), .O(N1390) );
nand2 gate351( .a(N1328), .b(N1242), .O(N1393) );
inv1 gate352( .a(N1243), .O(N1396) );
nand2 gate353( .a(N1243), .b(N1004), .O(N1397) );
inv1 gate354( .a(N1246), .O(N1398) );
nand2 gate355( .a(N1246), .b(N1007), .O(N1399) );
inv1 gate356( .a(N1319), .O(N1409) );
nand2 gate357( .a(N649), .b(N1346), .O(N1412) );
inv1 gate358( .a(N1334), .O(N1413) );
buf1 gate359( .a(N1264), .O(N1416) );
buf1 gate360( .a(N1264), .O(N1419) );
nand2 gate361( .a(N634), .b(N1386), .O(N1433) );
nand2 gate362( .a(N637), .b(N1388), .O(N1434) );
nand2 gate363( .a(N640), .b(N1396), .O(N1438) );

  xor2  gate1091(.a(N1398), .b(N646), .O(gate364inter0));
  nand2 gate1092(.a(gate364inter0), .b(s_30), .O(gate364inter1));
  and2  gate1093(.a(N1398), .b(N646), .O(gate364inter2));
  inv1  gate1094(.a(s_30), .O(gate364inter3));
  inv1  gate1095(.a(s_31), .O(gate364inter4));
  nand2 gate1096(.a(gate364inter4), .b(gate364inter3), .O(gate364inter5));
  nor2  gate1097(.a(gate364inter5), .b(gate364inter2), .O(gate364inter6));
  inv1  gate1098(.a(N646), .O(gate364inter7));
  inv1  gate1099(.a(N1398), .O(gate364inter8));
  nand2 gate1100(.a(gate364inter8), .b(gate364inter7), .O(gate364inter9));
  nand2 gate1101(.a(s_31), .b(gate364inter3), .O(gate364inter10));
  nor2  gate1102(.a(gate364inter10), .b(gate364inter9), .O(gate364inter11));
  nor2  gate1103(.a(gate364inter11), .b(gate364inter6), .O(gate364inter12));
  nand2 gate1104(.a(gate364inter12), .b(gate364inter1), .O(N1439));
inv1 gate365( .a(N1344), .O(N1440) );
nand2 gate366( .a(N1355), .b(N1148), .O(N1443) );
inv1 gate367( .a(N1355), .O(N1444) );

  xor2  gate2253(.a(N1149), .b(N1352), .O(gate368inter0));
  nand2 gate2254(.a(gate368inter0), .b(s_196), .O(gate368inter1));
  and2  gate2255(.a(N1149), .b(N1352), .O(gate368inter2));
  inv1  gate2256(.a(s_196), .O(gate368inter3));
  inv1  gate2257(.a(s_197), .O(gate368inter4));
  nand2 gate2258(.a(gate368inter4), .b(gate368inter3), .O(gate368inter5));
  nor2  gate2259(.a(gate368inter5), .b(gate368inter2), .O(gate368inter6));
  inv1  gate2260(.a(N1352), .O(gate368inter7));
  inv1  gate2261(.a(N1149), .O(gate368inter8));
  nand2 gate2262(.a(gate368inter8), .b(gate368inter7), .O(gate368inter9));
  nand2 gate2263(.a(s_197), .b(gate368inter3), .O(gate368inter10));
  nor2  gate2264(.a(gate368inter10), .b(gate368inter9), .O(gate368inter11));
  nor2  gate2265(.a(gate368inter11), .b(gate368inter6), .O(gate368inter12));
  nand2 gate2266(.a(gate368inter12), .b(gate368inter1), .O(N1445));
inv1 gate369( .a(N1352), .O(N1446) );
nand2 gate370( .a(N1358), .b(N1151), .O(N1447) );
inv1 gate371( .a(N1358), .O(N1448) );
nand2 gate372( .a(N1361), .b(N1152), .O(N1451) );
inv1 gate373( .a(N1361), .O(N1452) );
nand2 gate374( .a(N1367), .b(N1153), .O(N1453) );
inv1 gate375( .a(N1367), .O(N1454) );
nand2 gate376( .a(N1364), .b(N1154), .O(N1455) );
inv1 gate377( .a(N1364), .O(N1456) );
nand2 gate378( .a(N1373), .b(N1156), .O(N1457) );
inv1 gate379( .a(N1373), .O(N1458) );
nand2 gate380( .a(N1379), .b(N1157), .O(N1459) );
inv1 gate381( .a(N1379), .O(N1460) );
inv1 gate382( .a(N1383), .O(N1461) );
nand2 gate383( .a(N1393), .b(N1161), .O(N1462) );
inv1 gate384( .a(N1393), .O(N1463) );
nand2 gate385( .a(N1345), .b(N1412), .O(N1464) );
inv1 gate386( .a(N1370), .O(N1468) );
nand2 gate387( .a(N1370), .b(N1222), .O(N1469) );
inv1 gate388( .a(N1376), .O(N1470) );
nand2 gate389( .a(N1376), .b(N1227), .O(N1471) );
nand2 gate390( .a(N1387), .b(N1433), .O(N1472) );
inv1 gate391( .a(N1390), .O(N1475) );
nand2 gate392( .a(N1390), .b(N1240), .O(N1476) );
nand2 gate393( .a(N1389), .b(N1434), .O(N1478) );

  xor2  gate1679(.a(N1439), .b(N1399), .O(gate394inter0));
  nand2 gate1680(.a(gate394inter0), .b(s_114), .O(gate394inter1));
  and2  gate1681(.a(N1439), .b(N1399), .O(gate394inter2));
  inv1  gate1682(.a(s_114), .O(gate394inter3));
  inv1  gate1683(.a(s_115), .O(gate394inter4));
  nand2 gate1684(.a(gate394inter4), .b(gate394inter3), .O(gate394inter5));
  nor2  gate1685(.a(gate394inter5), .b(gate394inter2), .O(gate394inter6));
  inv1  gate1686(.a(N1399), .O(gate394inter7));
  inv1  gate1687(.a(N1439), .O(gate394inter8));
  nand2 gate1688(.a(gate394inter8), .b(gate394inter7), .O(gate394inter9));
  nand2 gate1689(.a(s_115), .b(gate394inter3), .O(gate394inter10));
  nor2  gate1690(.a(gate394inter10), .b(gate394inter9), .O(gate394inter11));
  nor2  gate1691(.a(gate394inter11), .b(gate394inter6), .O(gate394inter12));
  nand2 gate1692(.a(gate394inter12), .b(gate394inter1), .O(N1481));
nand2 gate395( .a(N1397), .b(N1438), .O(N1484) );
nand2 gate396( .a(N939), .b(N1444), .O(N1487) );
nand2 gate397( .a(N935), .b(N1446), .O(N1488) );
nand2 gate398( .a(N943), .b(N1448), .O(N1489) );
inv1 gate399( .a(N1419), .O(N1490) );
inv1 gate400( .a(N1416), .O(N1491) );
nand2 gate401( .a(N947), .b(N1452), .O(N1492) );

  xor2  gate1651(.a(N1454), .b(N955), .O(gate402inter0));
  nand2 gate1652(.a(gate402inter0), .b(s_110), .O(gate402inter1));
  and2  gate1653(.a(N1454), .b(N955), .O(gate402inter2));
  inv1  gate1654(.a(s_110), .O(gate402inter3));
  inv1  gate1655(.a(s_111), .O(gate402inter4));
  nand2 gate1656(.a(gate402inter4), .b(gate402inter3), .O(gate402inter5));
  nor2  gate1657(.a(gate402inter5), .b(gate402inter2), .O(gate402inter6));
  inv1  gate1658(.a(N955), .O(gate402inter7));
  inv1  gate1659(.a(N1454), .O(gate402inter8));
  nand2 gate1660(.a(gate402inter8), .b(gate402inter7), .O(gate402inter9));
  nand2 gate1661(.a(s_111), .b(gate402inter3), .O(gate402inter10));
  nor2  gate1662(.a(gate402inter10), .b(gate402inter9), .O(gate402inter11));
  nor2  gate1663(.a(gate402inter11), .b(gate402inter6), .O(gate402inter12));
  nand2 gate1664(.a(gate402inter12), .b(gate402inter1), .O(N1493));

  xor2  gate2351(.a(N1456), .b(N951), .O(gate403inter0));
  nand2 gate2352(.a(gate403inter0), .b(s_210), .O(gate403inter1));
  and2  gate2353(.a(N1456), .b(N951), .O(gate403inter2));
  inv1  gate2354(.a(s_210), .O(gate403inter3));
  inv1  gate2355(.a(s_211), .O(gate403inter4));
  nand2 gate2356(.a(gate403inter4), .b(gate403inter3), .O(gate403inter5));
  nor2  gate2357(.a(gate403inter5), .b(gate403inter2), .O(gate403inter6));
  inv1  gate2358(.a(N951), .O(gate403inter7));
  inv1  gate2359(.a(N1456), .O(gate403inter8));
  nand2 gate2360(.a(gate403inter8), .b(gate403inter7), .O(gate403inter9));
  nand2 gate2361(.a(s_211), .b(gate403inter3), .O(gate403inter10));
  nor2  gate2362(.a(gate403inter10), .b(gate403inter9), .O(gate403inter11));
  nor2  gate2363(.a(gate403inter11), .b(gate403inter6), .O(gate403inter12));
  nand2 gate2364(.a(gate403inter12), .b(gate403inter1), .O(N1494));
nand2 gate404( .a(N969), .b(N1458), .O(N1495) );

  xor2  gate1315(.a(N1460), .b(N977), .O(gate405inter0));
  nand2 gate1316(.a(gate405inter0), .b(s_62), .O(gate405inter1));
  and2  gate1317(.a(N1460), .b(N977), .O(gate405inter2));
  inv1  gate1318(.a(s_62), .O(gate405inter3));
  inv1  gate1319(.a(s_63), .O(gate405inter4));
  nand2 gate1320(.a(gate405inter4), .b(gate405inter3), .O(gate405inter5));
  nor2  gate1321(.a(gate405inter5), .b(gate405inter2), .O(gate405inter6));
  inv1  gate1322(.a(N977), .O(gate405inter7));
  inv1  gate1323(.a(N1460), .O(gate405inter8));
  nand2 gate1324(.a(gate405inter8), .b(gate405inter7), .O(gate405inter9));
  nand2 gate1325(.a(s_63), .b(gate405inter3), .O(gate405inter10));
  nor2  gate1326(.a(gate405inter10), .b(gate405inter9), .O(gate405inter11));
  nor2  gate1327(.a(gate405inter11), .b(gate405inter6), .O(gate405inter12));
  nand2 gate1328(.a(gate405inter12), .b(gate405inter1), .O(N1496));
nand2 gate406( .a(N998), .b(N1463), .O(N1498) );
inv1 gate407( .a(N1440), .O(N1499) );
nand2 gate408( .a(N965), .b(N1468), .O(N1500) );
nand2 gate409( .a(N973), .b(N1470), .O(N1501) );
nand2 gate410( .a(N994), .b(N1475), .O(N1504) );
inv1 gate411( .a(N1464), .O(N1510) );
nand2 gate412( .a(N1443), .b(N1487), .O(N1513) );
nand2 gate413( .a(N1445), .b(N1488), .O(N1514) );
nand2 gate414( .a(N1447), .b(N1489), .O(N1517) );

  xor2  gate1763(.a(N1492), .b(N1451), .O(gate415inter0));
  nand2 gate1764(.a(gate415inter0), .b(s_126), .O(gate415inter1));
  and2  gate1765(.a(N1492), .b(N1451), .O(gate415inter2));
  inv1  gate1766(.a(s_126), .O(gate415inter3));
  inv1  gate1767(.a(s_127), .O(gate415inter4));
  nand2 gate1768(.a(gate415inter4), .b(gate415inter3), .O(gate415inter5));
  nor2  gate1769(.a(gate415inter5), .b(gate415inter2), .O(gate415inter6));
  inv1  gate1770(.a(N1451), .O(gate415inter7));
  inv1  gate1771(.a(N1492), .O(gate415inter8));
  nand2 gate1772(.a(gate415inter8), .b(gate415inter7), .O(gate415inter9));
  nand2 gate1773(.a(s_127), .b(gate415inter3), .O(gate415inter10));
  nor2  gate1774(.a(gate415inter10), .b(gate415inter9), .O(gate415inter11));
  nor2  gate1775(.a(gate415inter11), .b(gate415inter6), .O(gate415inter12));
  nand2 gate1776(.a(gate415inter12), .b(gate415inter1), .O(N1520));

  xor2  gate2295(.a(N1493), .b(N1453), .O(gate416inter0));
  nand2 gate2296(.a(gate416inter0), .b(s_202), .O(gate416inter1));
  and2  gate2297(.a(N1493), .b(N1453), .O(gate416inter2));
  inv1  gate2298(.a(s_202), .O(gate416inter3));
  inv1  gate2299(.a(s_203), .O(gate416inter4));
  nand2 gate2300(.a(gate416inter4), .b(gate416inter3), .O(gate416inter5));
  nor2  gate2301(.a(gate416inter5), .b(gate416inter2), .O(gate416inter6));
  inv1  gate2302(.a(N1453), .O(gate416inter7));
  inv1  gate2303(.a(N1493), .O(gate416inter8));
  nand2 gate2304(.a(gate416inter8), .b(gate416inter7), .O(gate416inter9));
  nand2 gate2305(.a(s_203), .b(gate416inter3), .O(gate416inter10));
  nor2  gate2306(.a(gate416inter10), .b(gate416inter9), .O(gate416inter11));
  nor2  gate2307(.a(gate416inter11), .b(gate416inter6), .O(gate416inter12));
  nand2 gate2308(.a(gate416inter12), .b(gate416inter1), .O(N1521));
nand2 gate417( .a(N1455), .b(N1494), .O(N1522) );
nand2 gate418( .a(N1457), .b(N1495), .O(N1526) );
nand2 gate419( .a(N1459), .b(N1496), .O(N1527) );
inv1 gate420( .a(N1472), .O(N1528) );

  xor2  gate1735(.a(N1498), .b(N1462), .O(gate421inter0));
  nand2 gate1736(.a(gate421inter0), .b(s_122), .O(gate421inter1));
  and2  gate1737(.a(N1498), .b(N1462), .O(gate421inter2));
  inv1  gate1738(.a(s_122), .O(gate421inter3));
  inv1  gate1739(.a(s_123), .O(gate421inter4));
  nand2 gate1740(.a(gate421inter4), .b(gate421inter3), .O(gate421inter5));
  nor2  gate1741(.a(gate421inter5), .b(gate421inter2), .O(gate421inter6));
  inv1  gate1742(.a(N1462), .O(gate421inter7));
  inv1  gate1743(.a(N1498), .O(gate421inter8));
  nand2 gate1744(.a(gate421inter8), .b(gate421inter7), .O(gate421inter9));
  nand2 gate1745(.a(s_123), .b(gate421inter3), .O(gate421inter10));
  nor2  gate1746(.a(gate421inter10), .b(gate421inter9), .O(gate421inter11));
  nor2  gate1747(.a(gate421inter11), .b(gate421inter6), .O(gate421inter12));
  nand2 gate1748(.a(gate421inter12), .b(gate421inter1), .O(N1529));
inv1 gate422( .a(N1478), .O(N1530) );
inv1 gate423( .a(N1481), .O(N1531) );
inv1 gate424( .a(N1484), .O(N1532) );

  xor2  gate937(.a(N1501), .b(N1471), .O(gate425inter0));
  nand2 gate938(.a(gate425inter0), .b(s_8), .O(gate425inter1));
  and2  gate939(.a(N1501), .b(N1471), .O(gate425inter2));
  inv1  gate940(.a(s_8), .O(gate425inter3));
  inv1  gate941(.a(s_9), .O(gate425inter4));
  nand2 gate942(.a(gate425inter4), .b(gate425inter3), .O(gate425inter5));
  nor2  gate943(.a(gate425inter5), .b(gate425inter2), .O(gate425inter6));
  inv1  gate944(.a(N1471), .O(gate425inter7));
  inv1  gate945(.a(N1501), .O(gate425inter8));
  nand2 gate946(.a(gate425inter8), .b(gate425inter7), .O(gate425inter9));
  nand2 gate947(.a(s_9), .b(gate425inter3), .O(gate425inter10));
  nor2  gate948(.a(gate425inter10), .b(gate425inter9), .O(gate425inter11));
  nor2  gate949(.a(gate425inter11), .b(gate425inter6), .O(gate425inter12));
  nand2 gate950(.a(gate425inter12), .b(gate425inter1), .O(N1534));
nand2 gate426( .a(N1469), .b(N1500), .O(N1537) );
nand2 gate427( .a(N1476), .b(N1504), .O(N1540) );
inv1 gate428( .a(N1513), .O(N1546) );
inv1 gate429( .a(N1521), .O(N1554) );
inv1 gate430( .a(N1526), .O(N1557) );
inv1 gate431( .a(N1520), .O(N1561) );
nand2 gate432( .a(N1484), .b(N1531), .O(N1567) );
nand2 gate433( .a(N1481), .b(N1532), .O(N1568) );
inv1 gate434( .a(N1510), .O(N1569) );
inv1 gate435( .a(N1527), .O(N1571) );
inv1 gate436( .a(N1529), .O(N1576) );
buf1 gate437( .a(N1522), .O(N1588) );
inv1 gate438( .a(N1534), .O(N1591) );
inv1 gate439( .a(N1537), .O(N1593) );
nand2 gate440( .a(N1540), .b(N1530), .O(N1594) );
inv1 gate441( .a(N1540), .O(N1595) );
nand2 gate442( .a(N1567), .b(N1568), .O(N1596) );
buf1 gate443( .a(N1517), .O(N1600) );
buf1 gate444( .a(N1517), .O(N1603) );
buf1 gate445( .a(N1522), .O(N1606) );
buf1 gate446( .a(N1522), .O(N1609) );
buf1 gate447( .a(N1514), .O(N1612) );
buf1 gate448( .a(N1514), .O(N1615) );
buf1 gate449( .a(N1557), .O(N1620) );
buf1 gate450( .a(N1554), .O(N1623) );
inv1 gate451( .a(N1571), .O(N1635) );
nand2 gate452( .a(N1478), .b(N1595), .O(N1636) );
nand2 gate453( .a(N1576), .b(N1569), .O(N1638) );
inv1 gate454( .a(N1576), .O(N1639) );
buf1 gate455( .a(N1561), .O(N1640) );
buf1 gate456( .a(N1561), .O(N1643) );
buf1 gate457( .a(N1546), .O(N1647) );
buf1 gate458( .a(N1546), .O(N1651) );
buf1 gate459( .a(N1554), .O(N1658) );
buf1 gate460( .a(N1557), .O(N1661) );
buf1 gate461( .a(N1557), .O(N1664) );
nand2 gate462( .a(N1596), .b(N893), .O(N1671) );
inv1 gate463( .a(N1596), .O(N1672) );
inv1 gate464( .a(N1600), .O(N1675) );
inv1 gate465( .a(N1603), .O(N1677) );

  xor2  gate1273(.a(N1217), .b(N1606), .O(gate466inter0));
  nand2 gate1274(.a(gate466inter0), .b(s_56), .O(gate466inter1));
  and2  gate1275(.a(N1217), .b(N1606), .O(gate466inter2));
  inv1  gate1276(.a(s_56), .O(gate466inter3));
  inv1  gate1277(.a(s_57), .O(gate466inter4));
  nand2 gate1278(.a(gate466inter4), .b(gate466inter3), .O(gate466inter5));
  nor2  gate1279(.a(gate466inter5), .b(gate466inter2), .O(gate466inter6));
  inv1  gate1280(.a(N1606), .O(gate466inter7));
  inv1  gate1281(.a(N1217), .O(gate466inter8));
  nand2 gate1282(.a(gate466inter8), .b(gate466inter7), .O(gate466inter9));
  nand2 gate1283(.a(s_57), .b(gate466inter3), .O(gate466inter10));
  nor2  gate1284(.a(gate466inter10), .b(gate466inter9), .O(gate466inter11));
  nor2  gate1285(.a(gate466inter11), .b(gate466inter6), .O(gate466inter12));
  nand2 gate1286(.a(gate466inter12), .b(gate466inter1), .O(N1678));
inv1 gate467( .a(N1606), .O(N1679) );
nand2 gate468( .a(N1609), .b(N1219), .O(N1680) );
inv1 gate469( .a(N1609), .O(N1681) );
inv1 gate470( .a(N1612), .O(N1682) );
inv1 gate471( .a(N1615), .O(N1683) );
nand2 gate472( .a(N1594), .b(N1636), .O(N1685) );
nand2 gate473( .a(N1510), .b(N1639), .O(N1688) );
buf1 gate474( .a(N1588), .O(N1697) );
buf1 gate475( .a(N1588), .O(N1701) );
nand2 gate476( .a(N643), .b(N1672), .O(N1706) );
inv1 gate477( .a(N1643), .O(N1707) );
nand2 gate478( .a(N1647), .b(N1675), .O(N1708) );
inv1 gate479( .a(N1647), .O(N1709) );
nand2 gate480( .a(N1651), .b(N1677), .O(N1710) );
inv1 gate481( .a(N1651), .O(N1711) );
nand2 gate482( .a(N1028), .b(N1679), .O(N1712) );

  xor2  gate1175(.a(N1681), .b(N1031), .O(gate483inter0));
  nand2 gate1176(.a(gate483inter0), .b(s_42), .O(gate483inter1));
  and2  gate1177(.a(N1681), .b(N1031), .O(gate483inter2));
  inv1  gate1178(.a(s_42), .O(gate483inter3));
  inv1  gate1179(.a(s_43), .O(gate483inter4));
  nand2 gate1180(.a(gate483inter4), .b(gate483inter3), .O(gate483inter5));
  nor2  gate1181(.a(gate483inter5), .b(gate483inter2), .O(gate483inter6));
  inv1  gate1182(.a(N1031), .O(gate483inter7));
  inv1  gate1183(.a(N1681), .O(gate483inter8));
  nand2 gate1184(.a(gate483inter8), .b(gate483inter7), .O(gate483inter9));
  nand2 gate1185(.a(s_43), .b(gate483inter3), .O(gate483inter10));
  nor2  gate1186(.a(gate483inter10), .b(gate483inter9), .O(gate483inter11));
  nor2  gate1187(.a(gate483inter11), .b(gate483inter6), .O(gate483inter12));
  nand2 gate1188(.a(gate483inter12), .b(gate483inter1), .O(N1713));
buf1 gate484( .a(N1620), .O(N1714) );
buf1 gate485( .a(N1620), .O(N1717) );

  xor2  gate2169(.a(N1593), .b(N1658), .O(gate486inter0));
  nand2 gate2170(.a(gate486inter0), .b(s_184), .O(gate486inter1));
  and2  gate2171(.a(N1593), .b(N1658), .O(gate486inter2));
  inv1  gate2172(.a(s_184), .O(gate486inter3));
  inv1  gate2173(.a(s_185), .O(gate486inter4));
  nand2 gate2174(.a(gate486inter4), .b(gate486inter3), .O(gate486inter5));
  nor2  gate2175(.a(gate486inter5), .b(gate486inter2), .O(gate486inter6));
  inv1  gate2176(.a(N1658), .O(gate486inter7));
  inv1  gate2177(.a(N1593), .O(gate486inter8));
  nand2 gate2178(.a(gate486inter8), .b(gate486inter7), .O(gate486inter9));
  nand2 gate2179(.a(s_185), .b(gate486inter3), .O(gate486inter10));
  nor2  gate2180(.a(gate486inter10), .b(gate486inter9), .O(gate486inter11));
  nor2  gate2181(.a(gate486inter11), .b(gate486inter6), .O(gate486inter12));
  nand2 gate2182(.a(gate486inter12), .b(gate486inter1), .O(N1720));
inv1 gate487( .a(N1658), .O(N1721) );
nand2 gate488( .a(N1638), .b(N1688), .O(N1723) );
inv1 gate489( .a(N1661), .O(N1727) );
inv1 gate490( .a(N1640), .O(N1728) );
inv1 gate491( .a(N1664), .O(N1730) );
buf1 gate492( .a(N1623), .O(N1731) );
buf1 gate493( .a(N1623), .O(N1734) );
nand2 gate494( .a(N1685), .b(N1528), .O(N1740) );
inv1 gate495( .a(N1685), .O(N1741) );
nand2 gate496( .a(N1671), .b(N1706), .O(N1742) );
nand2 gate497( .a(N1600), .b(N1709), .O(N1746) );
nand2 gate498( .a(N1603), .b(N1711), .O(N1747) );
nand2 gate499( .a(N1678), .b(N1712), .O(N1748) );

  xor2  gate2183(.a(N1713), .b(N1680), .O(gate500inter0));
  nand2 gate2184(.a(gate500inter0), .b(s_186), .O(gate500inter1));
  and2  gate2185(.a(N1713), .b(N1680), .O(gate500inter2));
  inv1  gate2186(.a(s_186), .O(gate500inter3));
  inv1  gate2187(.a(s_187), .O(gate500inter4));
  nand2 gate2188(.a(gate500inter4), .b(gate500inter3), .O(gate500inter5));
  nor2  gate2189(.a(gate500inter5), .b(gate500inter2), .O(gate500inter6));
  inv1  gate2190(.a(N1680), .O(gate500inter7));
  inv1  gate2191(.a(N1713), .O(gate500inter8));
  nand2 gate2192(.a(gate500inter8), .b(gate500inter7), .O(gate500inter9));
  nand2 gate2193(.a(s_187), .b(gate500inter3), .O(gate500inter10));
  nor2  gate2194(.a(gate500inter10), .b(gate500inter9), .O(gate500inter11));
  nor2  gate2195(.a(gate500inter11), .b(gate500inter6), .O(gate500inter12));
  nand2 gate2196(.a(gate500inter12), .b(gate500inter1), .O(N1751));

  xor2  gate1665(.a(N1721), .b(N1537), .O(gate501inter0));
  nand2 gate1666(.a(gate501inter0), .b(s_112), .O(gate501inter1));
  and2  gate1667(.a(N1721), .b(N1537), .O(gate501inter2));
  inv1  gate1668(.a(s_112), .O(gate501inter3));
  inv1  gate1669(.a(s_113), .O(gate501inter4));
  nand2 gate1670(.a(gate501inter4), .b(gate501inter3), .O(gate501inter5));
  nor2  gate1671(.a(gate501inter5), .b(gate501inter2), .O(gate501inter6));
  inv1  gate1672(.a(N1537), .O(gate501inter7));
  inv1  gate1673(.a(N1721), .O(gate501inter8));
  nand2 gate1674(.a(gate501inter8), .b(gate501inter7), .O(gate501inter9));
  nand2 gate1675(.a(s_113), .b(gate501inter3), .O(gate501inter10));
  nor2  gate1676(.a(gate501inter10), .b(gate501inter9), .O(gate501inter11));
  nor2  gate1677(.a(gate501inter11), .b(gate501inter6), .O(gate501inter12));
  nand2 gate1678(.a(gate501inter12), .b(gate501inter1), .O(N1759));
inv1 gate502( .a(N1697), .O(N1761) );

  xor2  gate1875(.a(N1727), .b(N1697), .O(gate503inter0));
  nand2 gate1876(.a(gate503inter0), .b(s_142), .O(gate503inter1));
  and2  gate1877(.a(N1727), .b(N1697), .O(gate503inter2));
  inv1  gate1878(.a(s_142), .O(gate503inter3));
  inv1  gate1879(.a(s_143), .O(gate503inter4));
  nand2 gate1880(.a(gate503inter4), .b(gate503inter3), .O(gate503inter5));
  nor2  gate1881(.a(gate503inter5), .b(gate503inter2), .O(gate503inter6));
  inv1  gate1882(.a(N1697), .O(gate503inter7));
  inv1  gate1883(.a(N1727), .O(gate503inter8));
  nand2 gate1884(.a(gate503inter8), .b(gate503inter7), .O(gate503inter9));
  nand2 gate1885(.a(s_143), .b(gate503inter3), .O(gate503inter10));
  nor2  gate1886(.a(gate503inter10), .b(gate503inter9), .O(gate503inter11));
  nor2  gate1887(.a(gate503inter11), .b(gate503inter6), .O(gate503inter12));
  nand2 gate1888(.a(gate503inter12), .b(gate503inter1), .O(N1762));
inv1 gate504( .a(N1701), .O(N1763) );
nand2 gate505( .a(N1701), .b(N1730), .O(N1764) );
inv1 gate506( .a(N1717), .O(N1768) );
nand2 gate507( .a(N1472), .b(N1741), .O(N1769) );

  xor2  gate1357(.a(N1413), .b(N1723), .O(gate508inter0));
  nand2 gate1358(.a(gate508inter0), .b(s_68), .O(gate508inter1));
  and2  gate1359(.a(N1413), .b(N1723), .O(gate508inter2));
  inv1  gate1360(.a(s_68), .O(gate508inter3));
  inv1  gate1361(.a(s_69), .O(gate508inter4));
  nand2 gate1362(.a(gate508inter4), .b(gate508inter3), .O(gate508inter5));
  nor2  gate1363(.a(gate508inter5), .b(gate508inter2), .O(gate508inter6));
  inv1  gate1364(.a(N1723), .O(gate508inter7));
  inv1  gate1365(.a(N1413), .O(gate508inter8));
  nand2 gate1366(.a(gate508inter8), .b(gate508inter7), .O(gate508inter9));
  nand2 gate1367(.a(s_69), .b(gate508inter3), .O(gate508inter10));
  nor2  gate1368(.a(gate508inter10), .b(gate508inter9), .O(gate508inter11));
  nor2  gate1369(.a(gate508inter11), .b(gate508inter6), .O(gate508inter12));
  nand2 gate1370(.a(gate508inter12), .b(gate508inter1), .O(N1772));
inv1 gate509( .a(N1723), .O(N1773) );

  xor2  gate1721(.a(N1746), .b(N1708), .O(gate510inter0));
  nand2 gate1722(.a(gate510inter0), .b(s_120), .O(gate510inter1));
  and2  gate1723(.a(N1746), .b(N1708), .O(gate510inter2));
  inv1  gate1724(.a(s_120), .O(gate510inter3));
  inv1  gate1725(.a(s_121), .O(gate510inter4));
  nand2 gate1726(.a(gate510inter4), .b(gate510inter3), .O(gate510inter5));
  nor2  gate1727(.a(gate510inter5), .b(gate510inter2), .O(gate510inter6));
  inv1  gate1728(.a(N1708), .O(gate510inter7));
  inv1  gate1729(.a(N1746), .O(gate510inter8));
  nand2 gate1730(.a(gate510inter8), .b(gate510inter7), .O(gate510inter9));
  nand2 gate1731(.a(s_121), .b(gate510inter3), .O(gate510inter10));
  nor2  gate1732(.a(gate510inter10), .b(gate510inter9), .O(gate510inter11));
  nor2  gate1733(.a(gate510inter11), .b(gate510inter6), .O(gate510inter12));
  nand2 gate1734(.a(gate510inter12), .b(gate510inter1), .O(N1774));

  xor2  gate1511(.a(N1747), .b(N1710), .O(gate511inter0));
  nand2 gate1512(.a(gate511inter0), .b(s_90), .O(gate511inter1));
  and2  gate1513(.a(N1747), .b(N1710), .O(gate511inter2));
  inv1  gate1514(.a(s_90), .O(gate511inter3));
  inv1  gate1515(.a(s_91), .O(gate511inter4));
  nand2 gate1516(.a(gate511inter4), .b(gate511inter3), .O(gate511inter5));
  nor2  gate1517(.a(gate511inter5), .b(gate511inter2), .O(gate511inter6));
  inv1  gate1518(.a(N1710), .O(gate511inter7));
  inv1  gate1519(.a(N1747), .O(gate511inter8));
  nand2 gate1520(.a(gate511inter8), .b(gate511inter7), .O(gate511inter9));
  nand2 gate1521(.a(s_91), .b(gate511inter3), .O(gate511inter10));
  nor2  gate1522(.a(gate511inter10), .b(gate511inter9), .O(gate511inter11));
  nor2  gate1523(.a(gate511inter11), .b(gate511inter6), .O(gate511inter12));
  nand2 gate1524(.a(gate511inter12), .b(gate511inter1), .O(N1777));
inv1 gate512( .a(N1731), .O(N1783) );
nand2 gate513( .a(N1731), .b(N1682), .O(N1784) );
inv1 gate514( .a(N1714), .O(N1785) );
inv1 gate515( .a(N1734), .O(N1786) );
nand2 gate516( .a(N1734), .b(N1683), .O(N1787) );
nand2 gate517( .a(N1720), .b(N1759), .O(N1788) );
nand2 gate518( .a(N1661), .b(N1761), .O(N1791) );
nand2 gate519( .a(N1664), .b(N1763), .O(N1792) );
nand2 gate520( .a(N1751), .b(N1155), .O(N1795) );
inv1 gate521( .a(N1751), .O(N1796) );
nand2 gate522( .a(N1740), .b(N1769), .O(N1798) );
nand2 gate523( .a(N1334), .b(N1773), .O(N1801) );
nand2 gate524( .a(N1742), .b(N290), .O(N1802) );
inv1 gate525( .a(N1748), .O(N1807) );
nand2 gate526( .a(N1748), .b(N1218), .O(N1808) );
nand2 gate527( .a(N1612), .b(N1783), .O(N1809) );
nand2 gate528( .a(N1615), .b(N1786), .O(N1810) );
nand2 gate529( .a(N1791), .b(N1762), .O(N1812) );
nand2 gate530( .a(N1792), .b(N1764), .O(N1815) );
buf1 gate531( .a(N1742), .O(N1818) );
nand2 gate532( .a(N1777), .b(N1490), .O(N1821) );
inv1 gate533( .a(N1777), .O(N1822) );
nand2 gate534( .a(N1774), .b(N1491), .O(N1823) );
inv1 gate535( .a(N1774), .O(N1824) );
nand2 gate536( .a(N962), .b(N1796), .O(N1825) );
nand2 gate537( .a(N1788), .b(N1409), .O(N1826) );
inv1 gate538( .a(N1788), .O(N1827) );
nand2 gate539( .a(N1772), .b(N1801), .O(N1830) );

  xor2  gate909(.a(N1807), .b(N959), .O(gate540inter0));
  nand2 gate910(.a(gate540inter0), .b(s_4), .O(gate540inter1));
  and2  gate911(.a(N1807), .b(N959), .O(gate540inter2));
  inv1  gate912(.a(s_4), .O(gate540inter3));
  inv1  gate913(.a(s_5), .O(gate540inter4));
  nand2 gate914(.a(gate540inter4), .b(gate540inter3), .O(gate540inter5));
  nor2  gate915(.a(gate540inter5), .b(gate540inter2), .O(gate540inter6));
  inv1  gate916(.a(N959), .O(gate540inter7));
  inv1  gate917(.a(N1807), .O(gate540inter8));
  nand2 gate918(.a(gate540inter8), .b(gate540inter7), .O(gate540inter9));
  nand2 gate919(.a(s_5), .b(gate540inter3), .O(gate540inter10));
  nor2  gate920(.a(gate540inter10), .b(gate540inter9), .O(gate540inter11));
  nor2  gate921(.a(gate540inter11), .b(gate540inter6), .O(gate540inter12));
  nand2 gate922(.a(gate540inter12), .b(gate540inter1), .O(N1837));

  xor2  gate1119(.a(N1784), .b(N1809), .O(gate541inter0));
  nand2 gate1120(.a(gate541inter0), .b(s_34), .O(gate541inter1));
  and2  gate1121(.a(N1784), .b(N1809), .O(gate541inter2));
  inv1  gate1122(.a(s_34), .O(gate541inter3));
  inv1  gate1123(.a(s_35), .O(gate541inter4));
  nand2 gate1124(.a(gate541inter4), .b(gate541inter3), .O(gate541inter5));
  nor2  gate1125(.a(gate541inter5), .b(gate541inter2), .O(gate541inter6));
  inv1  gate1126(.a(N1809), .O(gate541inter7));
  inv1  gate1127(.a(N1784), .O(gate541inter8));
  nand2 gate1128(.a(gate541inter8), .b(gate541inter7), .O(gate541inter9));
  nand2 gate1129(.a(s_35), .b(gate541inter3), .O(gate541inter10));
  nor2  gate1130(.a(gate541inter10), .b(gate541inter9), .O(gate541inter11));
  nor2  gate1131(.a(gate541inter11), .b(gate541inter6), .O(gate541inter12));
  nand2 gate1132(.a(gate541inter12), .b(gate541inter1), .O(N1838));
nand2 gate542( .a(N1810), .b(N1787), .O(N1841) );
nand2 gate543( .a(N1419), .b(N1822), .O(N1848) );
nand2 gate544( .a(N1416), .b(N1824), .O(N1849) );
nand2 gate545( .a(N1795), .b(N1825), .O(N1850) );

  xor2  gate2155(.a(N1827), .b(N1319), .O(gate546inter0));
  nand2 gate2156(.a(gate546inter0), .b(s_182), .O(gate546inter1));
  and2  gate2157(.a(N1827), .b(N1319), .O(gate546inter2));
  inv1  gate2158(.a(s_182), .O(gate546inter3));
  inv1  gate2159(.a(s_183), .O(gate546inter4));
  nand2 gate2160(.a(gate546inter4), .b(gate546inter3), .O(gate546inter5));
  nor2  gate2161(.a(gate546inter5), .b(gate546inter2), .O(gate546inter6));
  inv1  gate2162(.a(N1319), .O(gate546inter7));
  inv1  gate2163(.a(N1827), .O(gate546inter8));
  nand2 gate2164(.a(gate546inter8), .b(gate546inter7), .O(gate546inter9));
  nand2 gate2165(.a(s_183), .b(gate546inter3), .O(gate546inter10));
  nor2  gate2166(.a(gate546inter10), .b(gate546inter9), .O(gate546inter11));
  nor2  gate2167(.a(gate546inter11), .b(gate546inter6), .O(gate546inter12));
  nand2 gate2168(.a(gate546inter12), .b(gate546inter1), .O(N1852));

  xor2  gate1791(.a(N1707), .b(N1815), .O(gate547inter0));
  nand2 gate1792(.a(gate547inter0), .b(s_130), .O(gate547inter1));
  and2  gate1793(.a(N1707), .b(N1815), .O(gate547inter2));
  inv1  gate1794(.a(s_130), .O(gate547inter3));
  inv1  gate1795(.a(s_131), .O(gate547inter4));
  nand2 gate1796(.a(gate547inter4), .b(gate547inter3), .O(gate547inter5));
  nor2  gate1797(.a(gate547inter5), .b(gate547inter2), .O(gate547inter6));
  inv1  gate1798(.a(N1815), .O(gate547inter7));
  inv1  gate1799(.a(N1707), .O(gate547inter8));
  nand2 gate1800(.a(gate547inter8), .b(gate547inter7), .O(gate547inter9));
  nand2 gate1801(.a(s_131), .b(gate547inter3), .O(gate547inter10));
  nor2  gate1802(.a(gate547inter10), .b(gate547inter9), .O(gate547inter11));
  nor2  gate1803(.a(gate547inter11), .b(gate547inter6), .O(gate547inter12));
  nand2 gate1804(.a(gate547inter12), .b(gate547inter1), .O(N1855));
inv1 gate548( .a(N1815), .O(N1856) );
inv1 gate549( .a(N1818), .O(N1857) );
nand2 gate550( .a(N1798), .b(N290), .O(N1858) );
inv1 gate551( .a(N1812), .O(N1864) );

  xor2  gate1805(.a(N1728), .b(N1812), .O(gate552inter0));
  nand2 gate1806(.a(gate552inter0), .b(s_132), .O(gate552inter1));
  and2  gate1807(.a(N1728), .b(N1812), .O(gate552inter2));
  inv1  gate1808(.a(s_132), .O(gate552inter3));
  inv1  gate1809(.a(s_133), .O(gate552inter4));
  nand2 gate1810(.a(gate552inter4), .b(gate552inter3), .O(gate552inter5));
  nor2  gate1811(.a(gate552inter5), .b(gate552inter2), .O(gate552inter6));
  inv1  gate1812(.a(N1812), .O(gate552inter7));
  inv1  gate1813(.a(N1728), .O(gate552inter8));
  nand2 gate1814(.a(gate552inter8), .b(gate552inter7), .O(gate552inter9));
  nand2 gate1815(.a(s_133), .b(gate552inter3), .O(gate552inter10));
  nor2  gate1816(.a(gate552inter10), .b(gate552inter9), .O(gate552inter11));
  nor2  gate1817(.a(gate552inter11), .b(gate552inter6), .O(gate552inter12));
  nand2 gate1818(.a(gate552inter12), .b(gate552inter1), .O(N1865));
buf1 gate553( .a(N1798), .O(N1866) );
buf1 gate554( .a(N1802), .O(N1869) );
buf1 gate555( .a(N1802), .O(N1872) );
nand2 gate556( .a(N1808), .b(N1837), .O(N1875) );
nand2 gate557( .a(N1821), .b(N1848), .O(N1878) );

  xor2  gate2057(.a(N1849), .b(N1823), .O(gate558inter0));
  nand2 gate2058(.a(gate558inter0), .b(s_168), .O(gate558inter1));
  and2  gate2059(.a(N1849), .b(N1823), .O(gate558inter2));
  inv1  gate2060(.a(s_168), .O(gate558inter3));
  inv1  gate2061(.a(s_169), .O(gate558inter4));
  nand2 gate2062(.a(gate558inter4), .b(gate558inter3), .O(gate558inter5));
  nor2  gate2063(.a(gate558inter5), .b(gate558inter2), .O(gate558inter6));
  inv1  gate2064(.a(N1823), .O(gate558inter7));
  inv1  gate2065(.a(N1849), .O(gate558inter8));
  nand2 gate2066(.a(gate558inter8), .b(gate558inter7), .O(gate558inter9));
  nand2 gate2067(.a(s_169), .b(gate558inter3), .O(gate558inter10));
  nor2  gate2068(.a(gate558inter10), .b(gate558inter9), .O(gate558inter11));
  nor2  gate2069(.a(gate558inter11), .b(gate558inter6), .O(gate558inter12));
  nand2 gate2070(.a(gate558inter12), .b(gate558inter1), .O(N1879));

  xor2  gate1553(.a(N1768), .b(N1841), .O(gate559inter0));
  nand2 gate1554(.a(gate559inter0), .b(s_96), .O(gate559inter1));
  and2  gate1555(.a(N1768), .b(N1841), .O(gate559inter2));
  inv1  gate1556(.a(s_96), .O(gate559inter3));
  inv1  gate1557(.a(s_97), .O(gate559inter4));
  nand2 gate1558(.a(gate559inter4), .b(gate559inter3), .O(gate559inter5));
  nor2  gate1559(.a(gate559inter5), .b(gate559inter2), .O(gate559inter6));
  inv1  gate1560(.a(N1841), .O(gate559inter7));
  inv1  gate1561(.a(N1768), .O(gate559inter8));
  nand2 gate1562(.a(gate559inter8), .b(gate559inter7), .O(gate559inter9));
  nand2 gate1563(.a(s_97), .b(gate559inter3), .O(gate559inter10));
  nor2  gate1564(.a(gate559inter10), .b(gate559inter9), .O(gate559inter11));
  nor2  gate1565(.a(gate559inter11), .b(gate559inter6), .O(gate559inter12));
  nand2 gate1566(.a(gate559inter12), .b(gate559inter1), .O(N1882));
inv1 gate560( .a(N1841), .O(N1883) );

  xor2  gate2211(.a(N1852), .b(N1826), .O(gate561inter0));
  nand2 gate2212(.a(gate561inter0), .b(s_190), .O(gate561inter1));
  and2  gate2213(.a(N1852), .b(N1826), .O(gate561inter2));
  inv1  gate2214(.a(s_190), .O(gate561inter3));
  inv1  gate2215(.a(s_191), .O(gate561inter4));
  nand2 gate2216(.a(gate561inter4), .b(gate561inter3), .O(gate561inter5));
  nor2  gate2217(.a(gate561inter5), .b(gate561inter2), .O(gate561inter6));
  inv1  gate2218(.a(N1826), .O(gate561inter7));
  inv1  gate2219(.a(N1852), .O(gate561inter8));
  nand2 gate2220(.a(gate561inter8), .b(gate561inter7), .O(gate561inter9));
  nand2 gate2221(.a(s_191), .b(gate561inter3), .O(gate561inter10));
  nor2  gate2222(.a(gate561inter10), .b(gate561inter9), .O(gate561inter11));
  nor2  gate2223(.a(gate561inter11), .b(gate561inter6), .O(gate561inter12));
  nand2 gate2224(.a(gate561inter12), .b(gate561inter1), .O(N1884));

  xor2  gate1287(.a(N1856), .b(N1643), .O(gate562inter0));
  nand2 gate1288(.a(gate562inter0), .b(s_58), .O(gate562inter1));
  and2  gate1289(.a(N1856), .b(N1643), .O(gate562inter2));
  inv1  gate1290(.a(s_58), .O(gate562inter3));
  inv1  gate1291(.a(s_59), .O(gate562inter4));
  nand2 gate1292(.a(gate562inter4), .b(gate562inter3), .O(gate562inter5));
  nor2  gate1293(.a(gate562inter5), .b(gate562inter2), .O(gate562inter6));
  inv1  gate1294(.a(N1643), .O(gate562inter7));
  inv1  gate1295(.a(N1856), .O(gate562inter8));
  nand2 gate1296(.a(gate562inter8), .b(gate562inter7), .O(gate562inter9));
  nand2 gate1297(.a(s_59), .b(gate562inter3), .O(gate562inter10));
  nor2  gate1298(.a(gate562inter10), .b(gate562inter9), .O(gate562inter11));
  nor2  gate1299(.a(gate562inter11), .b(gate562inter6), .O(gate562inter12));
  nand2 gate1300(.a(gate562inter12), .b(gate562inter1), .O(N1885));

  xor2  gate2071(.a(N290), .b(N1830), .O(gate563inter0));
  nand2 gate2072(.a(gate563inter0), .b(s_170), .O(gate563inter1));
  and2  gate2073(.a(N290), .b(N1830), .O(gate563inter2));
  inv1  gate2074(.a(s_170), .O(gate563inter3));
  inv1  gate2075(.a(s_171), .O(gate563inter4));
  nand2 gate2076(.a(gate563inter4), .b(gate563inter3), .O(gate563inter5));
  nor2  gate2077(.a(gate563inter5), .b(gate563inter2), .O(gate563inter6));
  inv1  gate2078(.a(N1830), .O(gate563inter7));
  inv1  gate2079(.a(N290), .O(gate563inter8));
  nand2 gate2080(.a(gate563inter8), .b(gate563inter7), .O(gate563inter9));
  nand2 gate2081(.a(s_171), .b(gate563inter3), .O(gate563inter10));
  nor2  gate2082(.a(gate563inter10), .b(gate563inter9), .O(gate563inter11));
  nor2  gate2083(.a(gate563inter11), .b(gate563inter6), .O(gate563inter12));
  nand2 gate2084(.a(gate563inter12), .b(gate563inter1), .O(N1889));
inv1 gate564( .a(N1838), .O(N1895) );

  xor2  gate1539(.a(N1785), .b(N1838), .O(gate565inter0));
  nand2 gate1540(.a(gate565inter0), .b(s_94), .O(gate565inter1));
  and2  gate1541(.a(N1785), .b(N1838), .O(gate565inter2));
  inv1  gate1542(.a(s_94), .O(gate565inter3));
  inv1  gate1543(.a(s_95), .O(gate565inter4));
  nand2 gate1544(.a(gate565inter4), .b(gate565inter3), .O(gate565inter5));
  nor2  gate1545(.a(gate565inter5), .b(gate565inter2), .O(gate565inter6));
  inv1  gate1546(.a(N1838), .O(gate565inter7));
  inv1  gate1547(.a(N1785), .O(gate565inter8));
  nand2 gate1548(.a(gate565inter8), .b(gate565inter7), .O(gate565inter9));
  nand2 gate1549(.a(s_95), .b(gate565inter3), .O(gate565inter10));
  nor2  gate1550(.a(gate565inter10), .b(gate565inter9), .O(gate565inter11));
  nor2  gate1551(.a(gate565inter11), .b(gate565inter6), .O(gate565inter12));
  nand2 gate1552(.a(gate565inter12), .b(gate565inter1), .O(N1896));
nand2 gate566( .a(N1640), .b(N1864), .O(N1897) );
inv1 gate567( .a(N1850), .O(N1898) );
buf1 gate568( .a(N1830), .O(N1902) );
inv1 gate569( .a(N1878), .O(N1910) );
nand2 gate570( .a(N1717), .b(N1883), .O(N1911) );
inv1 gate571( .a(N1884), .O(N1912) );
nand2 gate572( .a(N1855), .b(N1885), .O(N1913) );
inv1 gate573( .a(N1866), .O(N1915) );
nand2 gate574( .a(N1872), .b(N919), .O(N1919) );
inv1 gate575( .a(N1872), .O(N1920) );
nand2 gate576( .a(N1869), .b(N920), .O(N1921) );
inv1 gate577( .a(N1869), .O(N1922) );
inv1 gate578( .a(N1875), .O(N1923) );
nand2 gate579( .a(N1714), .b(N1895), .O(N1924) );
buf1 gate580( .a(N1858), .O(N1927) );
buf1 gate581( .a(N1858), .O(N1930) );

  xor2  gate1567(.a(N1897), .b(N1865), .O(gate582inter0));
  nand2 gate1568(.a(gate582inter0), .b(s_98), .O(gate582inter1));
  and2  gate1569(.a(N1897), .b(N1865), .O(gate582inter2));
  inv1  gate1570(.a(s_98), .O(gate582inter3));
  inv1  gate1571(.a(s_99), .O(gate582inter4));
  nand2 gate1572(.a(gate582inter4), .b(gate582inter3), .O(gate582inter5));
  nor2  gate1573(.a(gate582inter5), .b(gate582inter2), .O(gate582inter6));
  inv1  gate1574(.a(N1865), .O(gate582inter7));
  inv1  gate1575(.a(N1897), .O(gate582inter8));
  nand2 gate1576(.a(gate582inter8), .b(gate582inter7), .O(gate582inter9));
  nand2 gate1577(.a(s_99), .b(gate582inter3), .O(gate582inter10));
  nor2  gate1578(.a(gate582inter10), .b(gate582inter9), .O(gate582inter11));
  nor2  gate1579(.a(gate582inter11), .b(gate582inter6), .O(gate582inter12));
  nand2 gate1580(.a(gate582inter12), .b(gate582inter1), .O(N1933));
nand2 gate583( .a(N1882), .b(N1911), .O(N1936) );
inv1 gate584( .a(N1898), .O(N1937) );
inv1 gate585( .a(N1902), .O(N1938) );
nand2 gate586( .a(N679), .b(N1920), .O(N1941) );

  xor2  gate1707(.a(N1922), .b(N676), .O(gate587inter0));
  nand2 gate1708(.a(gate587inter0), .b(s_118), .O(gate587inter1));
  and2  gate1709(.a(N1922), .b(N676), .O(gate587inter2));
  inv1  gate1710(.a(s_118), .O(gate587inter3));
  inv1  gate1711(.a(s_119), .O(gate587inter4));
  nand2 gate1712(.a(gate587inter4), .b(gate587inter3), .O(gate587inter5));
  nor2  gate1713(.a(gate587inter5), .b(gate587inter2), .O(gate587inter6));
  inv1  gate1714(.a(N676), .O(gate587inter7));
  inv1  gate1715(.a(N1922), .O(gate587inter8));
  nand2 gate1716(.a(gate587inter8), .b(gate587inter7), .O(gate587inter9));
  nand2 gate1717(.a(s_119), .b(gate587inter3), .O(gate587inter10));
  nor2  gate1718(.a(gate587inter10), .b(gate587inter9), .O(gate587inter11));
  nor2  gate1719(.a(gate587inter11), .b(gate587inter6), .O(gate587inter12));
  nand2 gate1720(.a(gate587inter12), .b(gate587inter1), .O(N1942));
buf1 gate588( .a(N1879), .O(N1944) );
inv1 gate589( .a(N1913), .O(N1947) );
buf1 gate590( .a(N1889), .O(N1950) );
buf1 gate591( .a(N1889), .O(N1953) );
buf1 gate592( .a(N1879), .O(N1958) );
nand2 gate593( .a(N1896), .b(N1924), .O(N1961) );
and2 gate594( .a(N1910), .b(N601), .O(N1965) );
and2 gate595( .a(N602), .b(N1912), .O(N1968) );

  xor2  gate979(.a(N917), .b(N1930), .O(gate596inter0));
  nand2 gate980(.a(gate596inter0), .b(s_14), .O(gate596inter1));
  and2  gate981(.a(N917), .b(N1930), .O(gate596inter2));
  inv1  gate982(.a(s_14), .O(gate596inter3));
  inv1  gate983(.a(s_15), .O(gate596inter4));
  nand2 gate984(.a(gate596inter4), .b(gate596inter3), .O(gate596inter5));
  nor2  gate985(.a(gate596inter5), .b(gate596inter2), .O(gate596inter6));
  inv1  gate986(.a(N1930), .O(gate596inter7));
  inv1  gate987(.a(N917), .O(gate596inter8));
  nand2 gate988(.a(gate596inter8), .b(gate596inter7), .O(gate596inter9));
  nand2 gate989(.a(s_15), .b(gate596inter3), .O(gate596inter10));
  nor2  gate990(.a(gate596inter10), .b(gate596inter9), .O(gate596inter11));
  nor2  gate991(.a(gate596inter11), .b(gate596inter6), .O(gate596inter12));
  nand2 gate992(.a(gate596inter12), .b(gate596inter1), .O(N1975));
inv1 gate597( .a(N1930), .O(N1976) );
nand2 gate598( .a(N1927), .b(N918), .O(N1977) );
inv1 gate599( .a(N1927), .O(N1978) );

  xor2  gate1483(.a(N1941), .b(N1919), .O(gate600inter0));
  nand2 gate1484(.a(gate600inter0), .b(s_86), .O(gate600inter1));
  and2  gate1485(.a(N1941), .b(N1919), .O(gate600inter2));
  inv1  gate1486(.a(s_86), .O(gate600inter3));
  inv1  gate1487(.a(s_87), .O(gate600inter4));
  nand2 gate1488(.a(gate600inter4), .b(gate600inter3), .O(gate600inter5));
  nor2  gate1489(.a(gate600inter5), .b(gate600inter2), .O(gate600inter6));
  inv1  gate1490(.a(N1919), .O(gate600inter7));
  inv1  gate1491(.a(N1941), .O(gate600inter8));
  nand2 gate1492(.a(gate600inter8), .b(gate600inter7), .O(gate600inter9));
  nand2 gate1493(.a(s_87), .b(gate600inter3), .O(gate600inter10));
  nor2  gate1494(.a(gate600inter10), .b(gate600inter9), .O(gate600inter11));
  nor2  gate1495(.a(gate600inter11), .b(gate600inter6), .O(gate600inter12));
  nand2 gate1496(.a(gate600inter12), .b(gate600inter1), .O(N1979));
nand2 gate601( .a(N1921), .b(N1942), .O(N1980) );
inv1 gate602( .a(N1933), .O(N1985) );
inv1 gate603( .a(N1936), .O(N1987) );
inv1 gate604( .a(N1944), .O(N1999) );
nand2 gate605( .a(N1944), .b(N1937), .O(N2000) );
inv1 gate606( .a(N1947), .O(N2002) );
nand2 gate607( .a(N1947), .b(N1499), .O(N2003) );
nand2 gate608( .a(N1953), .b(N1350), .O(N2004) );
inv1 gate609( .a(N1953), .O(N2005) );

  xor2  gate1007(.a(N1351), .b(N1950), .O(gate610inter0));
  nand2 gate1008(.a(gate610inter0), .b(s_18), .O(gate610inter1));
  and2  gate1009(.a(N1351), .b(N1950), .O(gate610inter2));
  inv1  gate1010(.a(s_18), .O(gate610inter3));
  inv1  gate1011(.a(s_19), .O(gate610inter4));
  nand2 gate1012(.a(gate610inter4), .b(gate610inter3), .O(gate610inter5));
  nor2  gate1013(.a(gate610inter5), .b(gate610inter2), .O(gate610inter6));
  inv1  gate1014(.a(N1950), .O(gate610inter7));
  inv1  gate1015(.a(N1351), .O(gate610inter8));
  nand2 gate1016(.a(gate610inter8), .b(gate610inter7), .O(gate610inter9));
  nand2 gate1017(.a(s_19), .b(gate610inter3), .O(gate610inter10));
  nor2  gate1018(.a(gate610inter10), .b(gate610inter9), .O(gate610inter11));
  nor2  gate1019(.a(gate610inter11), .b(gate610inter6), .O(gate610inter12));
  nand2 gate1020(.a(gate610inter12), .b(gate610inter1), .O(N2006));
inv1 gate611( .a(N1950), .O(N2007) );
nand2 gate612( .a(N673), .b(N1976), .O(N2008) );
nand2 gate613( .a(N670), .b(N1978), .O(N2009) );
inv1 gate614( .a(N1979), .O(N2012) );
inv1 gate615( .a(N1958), .O(N2013) );
nand2 gate616( .a(N1958), .b(N1923), .O(N2014) );
inv1 gate617( .a(N1961), .O(N2015) );
nand2 gate618( .a(N1961), .b(N1635), .O(N2016) );
inv1 gate619( .a(N1965), .O(N2018) );
inv1 gate620( .a(N1968), .O(N2019) );
nand2 gate621( .a(N1898), .b(N1999), .O(N2020) );
inv1 gate622( .a(N1987), .O(N2021) );
nand2 gate623( .a(N1987), .b(N1591), .O(N2022) );

  xor2  gate2281(.a(N2002), .b(N1440), .O(gate624inter0));
  nand2 gate2282(.a(gate624inter0), .b(s_200), .O(gate624inter1));
  and2  gate2283(.a(N2002), .b(N1440), .O(gate624inter2));
  inv1  gate2284(.a(s_200), .O(gate624inter3));
  inv1  gate2285(.a(s_201), .O(gate624inter4));
  nand2 gate2286(.a(gate624inter4), .b(gate624inter3), .O(gate624inter5));
  nor2  gate2287(.a(gate624inter5), .b(gate624inter2), .O(gate624inter6));
  inv1  gate2288(.a(N1440), .O(gate624inter7));
  inv1  gate2289(.a(N2002), .O(gate624inter8));
  nand2 gate2290(.a(gate624inter8), .b(gate624inter7), .O(gate624inter9));
  nand2 gate2291(.a(s_201), .b(gate624inter3), .O(gate624inter10));
  nor2  gate2292(.a(gate624inter10), .b(gate624inter9), .O(gate624inter11));
  nor2  gate2293(.a(gate624inter11), .b(gate624inter6), .O(gate624inter12));
  nand2 gate2294(.a(gate624inter12), .b(gate624inter1), .O(N2023));
nand2 gate625( .a(N1261), .b(N2005), .O(N2024) );
nand2 gate626( .a(N1258), .b(N2007), .O(N2025) );
nand2 gate627( .a(N1975), .b(N2008), .O(N2026) );

  xor2  gate1371(.a(N2009), .b(N1977), .O(gate628inter0));
  nand2 gate1372(.a(gate628inter0), .b(s_70), .O(gate628inter1));
  and2  gate1373(.a(N2009), .b(N1977), .O(gate628inter2));
  inv1  gate1374(.a(s_70), .O(gate628inter3));
  inv1  gate1375(.a(s_71), .O(gate628inter4));
  nand2 gate1376(.a(gate628inter4), .b(gate628inter3), .O(gate628inter5));
  nor2  gate1377(.a(gate628inter5), .b(gate628inter2), .O(gate628inter6));
  inv1  gate1378(.a(N1977), .O(gate628inter7));
  inv1  gate1379(.a(N2009), .O(gate628inter8));
  nand2 gate1380(.a(gate628inter8), .b(gate628inter7), .O(gate628inter9));
  nand2 gate1381(.a(s_71), .b(gate628inter3), .O(gate628inter10));
  nor2  gate1382(.a(gate628inter10), .b(gate628inter9), .O(gate628inter11));
  nor2  gate1383(.a(gate628inter11), .b(gate628inter6), .O(gate628inter12));
  nand2 gate1384(.a(gate628inter12), .b(gate628inter1), .O(N2027));
inv1 gate629( .a(N1980), .O(N2030) );
buf1 gate630( .a(N1980), .O(N2033) );
nand2 gate631( .a(N1875), .b(N2013), .O(N2036) );

  xor2  gate1385(.a(N2015), .b(N1571), .O(gate632inter0));
  nand2 gate1386(.a(gate632inter0), .b(s_72), .O(gate632inter1));
  and2  gate1387(.a(N2015), .b(N1571), .O(gate632inter2));
  inv1  gate1388(.a(s_72), .O(gate632inter3));
  inv1  gate1389(.a(s_73), .O(gate632inter4));
  nand2 gate1390(.a(gate632inter4), .b(gate632inter3), .O(gate632inter5));
  nor2  gate1391(.a(gate632inter5), .b(gate632inter2), .O(gate632inter6));
  inv1  gate1392(.a(N1571), .O(gate632inter7));
  inv1  gate1393(.a(N2015), .O(gate632inter8));
  nand2 gate1394(.a(gate632inter8), .b(gate632inter7), .O(gate632inter9));
  nand2 gate1395(.a(s_73), .b(gate632inter3), .O(gate632inter10));
  nor2  gate1396(.a(gate632inter10), .b(gate632inter9), .O(gate632inter11));
  nor2  gate1397(.a(gate632inter11), .b(gate632inter6), .O(gate632inter12));
  nand2 gate1398(.a(gate632inter12), .b(gate632inter1), .O(N2037));
nand2 gate633( .a(N2020), .b(N2000), .O(N2038) );
nand2 gate634( .a(N1534), .b(N2021), .O(N2039) );

  xor2  gate2001(.a(N2003), .b(N2023), .O(gate635inter0));
  nand2 gate2002(.a(gate635inter0), .b(s_160), .O(gate635inter1));
  and2  gate2003(.a(N2003), .b(N2023), .O(gate635inter2));
  inv1  gate2004(.a(s_160), .O(gate635inter3));
  inv1  gate2005(.a(s_161), .O(gate635inter4));
  nand2 gate2006(.a(gate635inter4), .b(gate635inter3), .O(gate635inter5));
  nor2  gate2007(.a(gate635inter5), .b(gate635inter2), .O(gate635inter6));
  inv1  gate2008(.a(N2023), .O(gate635inter7));
  inv1  gate2009(.a(N2003), .O(gate635inter8));
  nand2 gate2010(.a(gate635inter8), .b(gate635inter7), .O(gate635inter9));
  nand2 gate2011(.a(s_161), .b(gate635inter3), .O(gate635inter10));
  nor2  gate2012(.a(gate635inter10), .b(gate635inter9), .O(gate635inter11));
  nor2  gate2013(.a(gate635inter11), .b(gate635inter6), .O(gate635inter12));
  nand2 gate2014(.a(gate635inter12), .b(gate635inter1), .O(N2040));
nand2 gate636( .a(N2004), .b(N2024), .O(N2041) );

  xor2  gate1035(.a(N2025), .b(N2006), .O(gate637inter0));
  nand2 gate1036(.a(gate637inter0), .b(s_22), .O(gate637inter1));
  and2  gate1037(.a(N2025), .b(N2006), .O(gate637inter2));
  inv1  gate1038(.a(s_22), .O(gate637inter3));
  inv1  gate1039(.a(s_23), .O(gate637inter4));
  nand2 gate1040(.a(gate637inter4), .b(gate637inter3), .O(gate637inter5));
  nor2  gate1041(.a(gate637inter5), .b(gate637inter2), .O(gate637inter6));
  inv1  gate1042(.a(N2006), .O(gate637inter7));
  inv1  gate1043(.a(N2025), .O(gate637inter8));
  nand2 gate1044(.a(gate637inter8), .b(gate637inter7), .O(gate637inter9));
  nand2 gate1045(.a(s_23), .b(gate637inter3), .O(gate637inter10));
  nor2  gate1046(.a(gate637inter10), .b(gate637inter9), .O(gate637inter11));
  nor2  gate1047(.a(gate637inter11), .b(gate637inter6), .O(gate637inter12));
  nand2 gate1048(.a(gate637inter12), .b(gate637inter1), .O(N2042));
inv1 gate638( .a(N2026), .O(N2047) );
nand2 gate639( .a(N2036), .b(N2014), .O(N2052) );
nand2 gate640( .a(N2037), .b(N2016), .O(N2055) );
inv1 gate641( .a(N2038), .O(N2060) );
nand2 gate642( .a(N2039), .b(N2022), .O(N2061) );

  xor2  gate1245(.a(N290), .b(N2040), .O(gate643inter0));
  nand2 gate1246(.a(gate643inter0), .b(s_52), .O(gate643inter1));
  and2  gate1247(.a(N290), .b(N2040), .O(gate643inter2));
  inv1  gate1248(.a(s_52), .O(gate643inter3));
  inv1  gate1249(.a(s_53), .O(gate643inter4));
  nand2 gate1250(.a(gate643inter4), .b(gate643inter3), .O(gate643inter5));
  nor2  gate1251(.a(gate643inter5), .b(gate643inter2), .O(gate643inter6));
  inv1  gate1252(.a(N2040), .O(gate643inter7));
  inv1  gate1253(.a(N290), .O(gate643inter8));
  nand2 gate1254(.a(gate643inter8), .b(gate643inter7), .O(gate643inter9));
  nand2 gate1255(.a(s_53), .b(gate643inter3), .O(gate643inter10));
  nor2  gate1256(.a(gate643inter10), .b(gate643inter9), .O(gate643inter11));
  nor2  gate1257(.a(gate643inter11), .b(gate643inter6), .O(gate643inter12));
  nand2 gate1258(.a(gate643inter12), .b(gate643inter1), .O(N2062));
inv1 gate644( .a(N2041), .O(N2067) );
inv1 gate645( .a(N2027), .O(N2068) );
buf1 gate646( .a(N2027), .O(N2071) );
inv1 gate647( .a(N2052), .O(N2076) );
inv1 gate648( .a(N2055), .O(N2077) );

  xor2  gate1959(.a(N290), .b(N2060), .O(gate649inter0));
  nand2 gate1960(.a(gate649inter0), .b(s_154), .O(gate649inter1));
  and2  gate1961(.a(N290), .b(N2060), .O(gate649inter2));
  inv1  gate1962(.a(s_154), .O(gate649inter3));
  inv1  gate1963(.a(s_155), .O(gate649inter4));
  nand2 gate1964(.a(gate649inter4), .b(gate649inter3), .O(gate649inter5));
  nor2  gate1965(.a(gate649inter5), .b(gate649inter2), .O(gate649inter6));
  inv1  gate1966(.a(N2060), .O(gate649inter7));
  inv1  gate1967(.a(N290), .O(gate649inter8));
  nand2 gate1968(.a(gate649inter8), .b(gate649inter7), .O(gate649inter9));
  nand2 gate1969(.a(s_155), .b(gate649inter3), .O(gate649inter10));
  nor2  gate1970(.a(gate649inter10), .b(gate649inter9), .O(gate649inter11));
  nor2  gate1971(.a(gate649inter11), .b(gate649inter6), .O(gate649inter12));
  nand2 gate1972(.a(gate649inter12), .b(gate649inter1), .O(N2078));
nand2 gate650( .a(N2061), .b(N290), .O(N2081) );
inv1 gate651( .a(N2042), .O(N2086) );
buf1 gate652( .a(N2042), .O(N2089) );
and2 gate653( .a(N2030), .b(N2068), .O(N2104) );
and2 gate654( .a(N2033), .b(N2068), .O(N2119) );
and2 gate655( .a(N2030), .b(N2071), .O(N2129) );
and2 gate656( .a(N2033), .b(N2071), .O(N2143) );
buf1 gate657( .a(N2062), .O(N2148) );
buf1 gate658( .a(N2062), .O(N2151) );
buf1 gate659( .a(N2078), .O(N2196) );
buf1 gate660( .a(N2078), .O(N2199) );
buf1 gate661( .a(N2081), .O(N2202) );
buf1 gate662( .a(N2081), .O(N2205) );

  xor2  gate1077(.a(N915), .b(N2151), .O(gate663inter0));
  nand2 gate1078(.a(gate663inter0), .b(s_28), .O(gate663inter1));
  and2  gate1079(.a(N915), .b(N2151), .O(gate663inter2));
  inv1  gate1080(.a(s_28), .O(gate663inter3));
  inv1  gate1081(.a(s_29), .O(gate663inter4));
  nand2 gate1082(.a(gate663inter4), .b(gate663inter3), .O(gate663inter5));
  nor2  gate1083(.a(gate663inter5), .b(gate663inter2), .O(gate663inter6));
  inv1  gate1084(.a(N2151), .O(gate663inter7));
  inv1  gate1085(.a(N915), .O(gate663inter8));
  nand2 gate1086(.a(gate663inter8), .b(gate663inter7), .O(gate663inter9));
  nand2 gate1087(.a(s_29), .b(gate663inter3), .O(gate663inter10));
  nor2  gate1088(.a(gate663inter10), .b(gate663inter9), .O(gate663inter11));
  nor2  gate1089(.a(gate663inter11), .b(gate663inter6), .O(gate663inter12));
  nand2 gate1090(.a(gate663inter12), .b(gate663inter1), .O(N2214));
inv1 gate664( .a(N2151), .O(N2215) );

  xor2  gate1343(.a(N916), .b(N2148), .O(gate665inter0));
  nand2 gate1344(.a(gate665inter0), .b(s_66), .O(gate665inter1));
  and2  gate1345(.a(N916), .b(N2148), .O(gate665inter2));
  inv1  gate1346(.a(s_66), .O(gate665inter3));
  inv1  gate1347(.a(s_67), .O(gate665inter4));
  nand2 gate1348(.a(gate665inter4), .b(gate665inter3), .O(gate665inter5));
  nor2  gate1349(.a(gate665inter5), .b(gate665inter2), .O(gate665inter6));
  inv1  gate1350(.a(N2148), .O(gate665inter7));
  inv1  gate1351(.a(N916), .O(gate665inter8));
  nand2 gate1352(.a(gate665inter8), .b(gate665inter7), .O(gate665inter9));
  nand2 gate1353(.a(s_67), .b(gate665inter3), .O(gate665inter10));
  nor2  gate1354(.a(gate665inter10), .b(gate665inter9), .O(gate665inter11));
  nor2  gate1355(.a(gate665inter11), .b(gate665inter6), .O(gate665inter12));
  nand2 gate1356(.a(gate665inter12), .b(gate665inter1), .O(N2216));
inv1 gate666( .a(N2148), .O(N2217) );
nand2 gate667( .a(N2199), .b(N1348), .O(N2222) );
inv1 gate668( .a(N2199), .O(N2223) );
nand2 gate669( .a(N2196), .b(N1349), .O(N2224) );
inv1 gate670( .a(N2196), .O(N2225) );
nand2 gate671( .a(N2205), .b(N913), .O(N2226) );
inv1 gate672( .a(N2205), .O(N2227) );

  xor2  gate1819(.a(N914), .b(N2202), .O(gate673inter0));
  nand2 gate1820(.a(gate673inter0), .b(s_134), .O(gate673inter1));
  and2  gate1821(.a(N914), .b(N2202), .O(gate673inter2));
  inv1  gate1822(.a(s_134), .O(gate673inter3));
  inv1  gate1823(.a(s_135), .O(gate673inter4));
  nand2 gate1824(.a(gate673inter4), .b(gate673inter3), .O(gate673inter5));
  nor2  gate1825(.a(gate673inter5), .b(gate673inter2), .O(gate673inter6));
  inv1  gate1826(.a(N2202), .O(gate673inter7));
  inv1  gate1827(.a(N914), .O(gate673inter8));
  nand2 gate1828(.a(gate673inter8), .b(gate673inter7), .O(gate673inter9));
  nand2 gate1829(.a(s_135), .b(gate673inter3), .O(gate673inter10));
  nor2  gate1830(.a(gate673inter10), .b(gate673inter9), .O(gate673inter11));
  nor2  gate1831(.a(gate673inter11), .b(gate673inter6), .O(gate673inter12));
  nand2 gate1832(.a(gate673inter12), .b(gate673inter1), .O(N2228));
inv1 gate674( .a(N2202), .O(N2229) );

  xor2  gate2141(.a(N2215), .b(N667), .O(gate675inter0));
  nand2 gate2142(.a(gate675inter0), .b(s_180), .O(gate675inter1));
  and2  gate2143(.a(N2215), .b(N667), .O(gate675inter2));
  inv1  gate2144(.a(s_180), .O(gate675inter3));
  inv1  gate2145(.a(s_181), .O(gate675inter4));
  nand2 gate2146(.a(gate675inter4), .b(gate675inter3), .O(gate675inter5));
  nor2  gate2147(.a(gate675inter5), .b(gate675inter2), .O(gate675inter6));
  inv1  gate2148(.a(N667), .O(gate675inter7));
  inv1  gate2149(.a(N2215), .O(gate675inter8));
  nand2 gate2150(.a(gate675inter8), .b(gate675inter7), .O(gate675inter9));
  nand2 gate2151(.a(s_181), .b(gate675inter3), .O(gate675inter10));
  nor2  gate2152(.a(gate675inter10), .b(gate675inter9), .O(gate675inter11));
  nor2  gate2153(.a(gate675inter11), .b(gate675inter6), .O(gate675inter12));
  nand2 gate2154(.a(gate675inter12), .b(gate675inter1), .O(N2230));
nand2 gate676( .a(N664), .b(N2217), .O(N2231) );
nand2 gate677( .a(N1255), .b(N2223), .O(N2232) );
nand2 gate678( .a(N1252), .b(N2225), .O(N2233) );
nand2 gate679( .a(N661), .b(N2227), .O(N2234) );
nand2 gate680( .a(N658), .b(N2229), .O(N2235) );
nand2 gate681( .a(N2214), .b(N2230), .O(N2236) );
nand2 gate682( .a(N2216), .b(N2231), .O(N2237) );
nand2 gate683( .a(N2222), .b(N2232), .O(N2240) );

  xor2  gate1189(.a(N2233), .b(N2224), .O(gate684inter0));
  nand2 gate1190(.a(gate684inter0), .b(s_44), .O(gate684inter1));
  and2  gate1191(.a(N2233), .b(N2224), .O(gate684inter2));
  inv1  gate1192(.a(s_44), .O(gate684inter3));
  inv1  gate1193(.a(s_45), .O(gate684inter4));
  nand2 gate1194(.a(gate684inter4), .b(gate684inter3), .O(gate684inter5));
  nor2  gate1195(.a(gate684inter5), .b(gate684inter2), .O(gate684inter6));
  inv1  gate1196(.a(N2224), .O(gate684inter7));
  inv1  gate1197(.a(N2233), .O(gate684inter8));
  nand2 gate1198(.a(gate684inter8), .b(gate684inter7), .O(gate684inter9));
  nand2 gate1199(.a(s_45), .b(gate684inter3), .O(gate684inter10));
  nor2  gate1200(.a(gate684inter10), .b(gate684inter9), .O(gate684inter11));
  nor2  gate1201(.a(gate684inter11), .b(gate684inter6), .O(gate684inter12));
  nand2 gate1202(.a(gate684inter12), .b(gate684inter1), .O(N2241));
nand2 gate685( .a(N2226), .b(N2234), .O(N2244) );
nand2 gate686( .a(N2228), .b(N2235), .O(N2245) );
inv1 gate687( .a(N2236), .O(N2250) );
inv1 gate688( .a(N2240), .O(N2253) );
inv1 gate689( .a(N2244), .O(N2256) );
inv1 gate690( .a(N2237), .O(N2257) );
buf1 gate691( .a(N2237), .O(N2260) );
inv1 gate692( .a(N2241), .O(N2263) );
and2 gate693( .a(N1164), .b(N2241), .O(N2266) );
inv1 gate694( .a(N2245), .O(N2269) );
and2 gate695( .a(N1168), .b(N2245), .O(N2272) );
nand8 gate696( .a(N2067), .b(N2012), .c(N2047), .d(N2250), .e(N899), .f(N2256), .g(N2253), .h(N903), .O(N2279) );
buf1 gate697( .a(N2266), .O(N2286) );
buf1 gate698( .a(N2266), .O(N2297) );
buf1 gate699( .a(N2272), .O(N2315) );
buf1 gate700( .a(N2272), .O(N2326) );
and2 gate701( .a(N2086), .b(N2257), .O(N2340) );
and2 gate702( .a(N2089), .b(N2257), .O(N2353) );
and2 gate703( .a(N2086), .b(N2260), .O(N2361) );
and2 gate704( .a(N2089), .b(N2260), .O(N2375) );
and4 gate705( .a(N338), .b(N2279), .c(N313), .d(N313), .O(N2384) );
and2 gate706( .a(N1163), .b(N2263), .O(N2385) );
and2 gate707( .a(N1164), .b(N2263), .O(N2386) );
and2 gate708( .a(N1167), .b(N2269), .O(N2426) );
and2 gate709( .a(N1168), .b(N2269), .O(N2427) );
nand5 gate710( .a(N2286), .b(N2315), .c(N2361), .d(N2104), .e(N1171), .O(N2537) );
nand5 gate711( .a(N2286), .b(N2315), .c(N2340), .d(N2129), .e(N1171), .O(N2540) );
nand5 gate712( .a(N2286), .b(N2315), .c(N2340), .d(N2119), .e(N1171), .O(N2543) );
nand5 gate713( .a(N2286), .b(N2315), .c(N2353), .d(N2104), .e(N1171), .O(N2546) );
nand5 gate714( .a(N2297), .b(N2315), .c(N2375), .d(N2119), .e(N1188), .O(N2549) );
nand5 gate715( .a(N2297), .b(N2326), .c(N2361), .d(N2143), .e(N1188), .O(N2552) );
nand5 gate716( .a(N2297), .b(N2326), .c(N2375), .d(N2129), .e(N1188), .O(N2555) );
and5 gate717( .a(N2286), .b(N2315), .c(N2361), .d(N2104), .e(N1171), .O(N2558) );
and5 gate718( .a(N2286), .b(N2315), .c(N2340), .d(N2129), .e(N1171), .O(N2561) );
and5 gate719( .a(N2286), .b(N2315), .c(N2340), .d(N2119), .e(N1171), .O(N2564) );
and5 gate720( .a(N2286), .b(N2315), .c(N2353), .d(N2104), .e(N1171), .O(N2567) );
and5 gate721( .a(N2297), .b(N2315), .c(N2375), .d(N2119), .e(N1188), .O(N2570) );
and5 gate722( .a(N2297), .b(N2326), .c(N2361), .d(N2143), .e(N1188), .O(N2573) );
and5 gate723( .a(N2297), .b(N2326), .c(N2375), .d(N2129), .e(N1188), .O(N2576) );
nand5 gate724( .a(N2286), .b(N2427), .c(N2361), .d(N2129), .e(N1171), .O(N2594) );
nand5 gate725( .a(N2297), .b(N2427), .c(N2361), .d(N2119), .e(N1171), .O(N2597) );
nand5 gate726( .a(N2297), .b(N2427), .c(N2375), .d(N2104), .e(N1171), .O(N2600) );
nand5 gate727( .a(N2297), .b(N2427), .c(N2340), .d(N2143), .e(N1171), .O(N2603) );
nand5 gate728( .a(N2297), .b(N2427), .c(N2353), .d(N2129), .e(N1188), .O(N2606) );
nand5 gate729( .a(N2386), .b(N2326), .c(N2361), .d(N2129), .e(N1188), .O(N2611) );
nand5 gate730( .a(N2386), .b(N2326), .c(N2361), .d(N2119), .e(N1188), .O(N2614) );
nand5 gate731( .a(N2386), .b(N2326), .c(N2375), .d(N2104), .e(N1188), .O(N2617) );
nand5 gate732( .a(N2386), .b(N2326), .c(N2353), .d(N2129), .e(N1188), .O(N2620) );
nand5 gate733( .a(N2297), .b(N2427), .c(N2340), .d(N2104), .e(N926), .O(N2627) );
nand5 gate734( .a(N2386), .b(N2326), .c(N2340), .d(N2104), .e(N926), .O(N2628) );
nand5 gate735( .a(N2386), .b(N2427), .c(N2361), .d(N2104), .e(N926), .O(N2629) );
nand5 gate736( .a(N2386), .b(N2427), .c(N2340), .d(N2129), .e(N926), .O(N2630) );
nand5 gate737( .a(N2386), .b(N2427), .c(N2340), .d(N2119), .e(N926), .O(N2631) );
nand5 gate738( .a(N2386), .b(N2427), .c(N2353), .d(N2104), .e(N926), .O(N2632) );
nand5 gate739( .a(N2386), .b(N2426), .c(N2340), .d(N2104), .e(N926), .O(N2633) );
nand5 gate740( .a(N2385), .b(N2427), .c(N2340), .d(N2104), .e(N926), .O(N2634) );
and5 gate741( .a(N2286), .b(N2427), .c(N2361), .d(N2129), .e(N1171), .O(N2639) );
and5 gate742( .a(N2297), .b(N2427), .c(N2361), .d(N2119), .e(N1171), .O(N2642) );
and5 gate743( .a(N2297), .b(N2427), .c(N2375), .d(N2104), .e(N1171), .O(N2645) );
and5 gate744( .a(N2297), .b(N2427), .c(N2340), .d(N2143), .e(N1171), .O(N2648) );
and5 gate745( .a(N2297), .b(N2427), .c(N2353), .d(N2129), .e(N1188), .O(N2651) );
and5 gate746( .a(N2386), .b(N2326), .c(N2361), .d(N2129), .e(N1188), .O(N2655) );
and5 gate747( .a(N2386), .b(N2326), .c(N2361), .d(N2119), .e(N1188), .O(N2658) );
and5 gate748( .a(N2386), .b(N2326), .c(N2375), .d(N2104), .e(N1188), .O(N2661) );
and5 gate749( .a(N2386), .b(N2326), .c(N2353), .d(N2129), .e(N1188), .O(N2664) );
nand2 gate750( .a(N2558), .b(N534), .O(N2669) );
inv1 gate751( .a(N2558), .O(N2670) );
nand2 gate752( .a(N2561), .b(N535), .O(N2671) );
inv1 gate753( .a(N2561), .O(N2672) );

  xor2  gate2099(.a(N536), .b(N2564), .O(gate754inter0));
  nand2 gate2100(.a(gate754inter0), .b(s_174), .O(gate754inter1));
  and2  gate2101(.a(N536), .b(N2564), .O(gate754inter2));
  inv1  gate2102(.a(s_174), .O(gate754inter3));
  inv1  gate2103(.a(s_175), .O(gate754inter4));
  nand2 gate2104(.a(gate754inter4), .b(gate754inter3), .O(gate754inter5));
  nor2  gate2105(.a(gate754inter5), .b(gate754inter2), .O(gate754inter6));
  inv1  gate2106(.a(N2564), .O(gate754inter7));
  inv1  gate2107(.a(N536), .O(gate754inter8));
  nand2 gate2108(.a(gate754inter8), .b(gate754inter7), .O(gate754inter9));
  nand2 gate2109(.a(s_175), .b(gate754inter3), .O(gate754inter10));
  nor2  gate2110(.a(gate754inter10), .b(gate754inter9), .O(gate754inter11));
  nor2  gate2111(.a(gate754inter11), .b(gate754inter6), .O(gate754inter12));
  nand2 gate2112(.a(gate754inter12), .b(gate754inter1), .O(N2673));
inv1 gate755( .a(N2564), .O(N2674) );
nand2 gate756( .a(N2567), .b(N537), .O(N2675) );
inv1 gate757( .a(N2567), .O(N2676) );
nand2 gate758( .a(N2570), .b(N543), .O(N2682) );
inv1 gate759( .a(N2570), .O(N2683) );
nand2 gate760( .a(N2573), .b(N548), .O(N2688) );
inv1 gate761( .a(N2573), .O(N2689) );

  xor2  gate1063(.a(N549), .b(N2576), .O(gate762inter0));
  nand2 gate1064(.a(gate762inter0), .b(s_26), .O(gate762inter1));
  and2  gate1065(.a(N549), .b(N2576), .O(gate762inter2));
  inv1  gate1066(.a(s_26), .O(gate762inter3));
  inv1  gate1067(.a(s_27), .O(gate762inter4));
  nand2 gate1068(.a(gate762inter4), .b(gate762inter3), .O(gate762inter5));
  nor2  gate1069(.a(gate762inter5), .b(gate762inter2), .O(gate762inter6));
  inv1  gate1070(.a(N2576), .O(gate762inter7));
  inv1  gate1071(.a(N549), .O(gate762inter8));
  nand2 gate1072(.a(gate762inter8), .b(gate762inter7), .O(gate762inter9));
  nand2 gate1073(.a(s_27), .b(gate762inter3), .O(gate762inter10));
  nor2  gate1074(.a(gate762inter10), .b(gate762inter9), .O(gate762inter11));
  nor2  gate1075(.a(gate762inter11), .b(gate762inter6), .O(gate762inter12));
  nand2 gate1076(.a(gate762inter12), .b(gate762inter1), .O(N2690));
inv1 gate763( .a(N2576), .O(N2691) );
and8 gate764( .a(N2627), .b(N2628), .c(N2629), .d(N2630), .e(N2631), .f(N2632), .g(N2633), .h(N2634), .O(N2710) );
nand2 gate765( .a(N343), .b(N2670), .O(N2720) );
nand2 gate766( .a(N346), .b(N2672), .O(N2721) );
nand2 gate767( .a(N349), .b(N2674), .O(N2722) );
nand2 gate768( .a(N352), .b(N2676), .O(N2723) );
nand2 gate769( .a(N2639), .b(N538), .O(N2724) );
inv1 gate770( .a(N2639), .O(N2725) );
nand2 gate771( .a(N2642), .b(N539), .O(N2726) );
inv1 gate772( .a(N2642), .O(N2727) );
nand2 gate773( .a(N2645), .b(N540), .O(N2728) );
inv1 gate774( .a(N2645), .O(N2729) );
nand2 gate775( .a(N2648), .b(N541), .O(N2730) );
inv1 gate776( .a(N2648), .O(N2731) );
nand2 gate777( .a(N2651), .b(N542), .O(N2732) );
inv1 gate778( .a(N2651), .O(N2733) );
nand2 gate779( .a(N370), .b(N2683), .O(N2734) );
nand2 gate780( .a(N2655), .b(N544), .O(N2735) );
inv1 gate781( .a(N2655), .O(N2736) );

  xor2  gate1609(.a(N545), .b(N2658), .O(gate782inter0));
  nand2 gate1610(.a(gate782inter0), .b(s_104), .O(gate782inter1));
  and2  gate1611(.a(N545), .b(N2658), .O(gate782inter2));
  inv1  gate1612(.a(s_104), .O(gate782inter3));
  inv1  gate1613(.a(s_105), .O(gate782inter4));
  nand2 gate1614(.a(gate782inter4), .b(gate782inter3), .O(gate782inter5));
  nor2  gate1615(.a(gate782inter5), .b(gate782inter2), .O(gate782inter6));
  inv1  gate1616(.a(N2658), .O(gate782inter7));
  inv1  gate1617(.a(N545), .O(gate782inter8));
  nand2 gate1618(.a(gate782inter8), .b(gate782inter7), .O(gate782inter9));
  nand2 gate1619(.a(s_105), .b(gate782inter3), .O(gate782inter10));
  nor2  gate1620(.a(gate782inter10), .b(gate782inter9), .O(gate782inter11));
  nor2  gate1621(.a(gate782inter11), .b(gate782inter6), .O(gate782inter12));
  nand2 gate1622(.a(gate782inter12), .b(gate782inter1), .O(N2737));
inv1 gate783( .a(N2658), .O(N2738) );

  xor2  gate1623(.a(N546), .b(N2661), .O(gate784inter0));
  nand2 gate1624(.a(gate784inter0), .b(s_106), .O(gate784inter1));
  and2  gate1625(.a(N546), .b(N2661), .O(gate784inter2));
  inv1  gate1626(.a(s_106), .O(gate784inter3));
  inv1  gate1627(.a(s_107), .O(gate784inter4));
  nand2 gate1628(.a(gate784inter4), .b(gate784inter3), .O(gate784inter5));
  nor2  gate1629(.a(gate784inter5), .b(gate784inter2), .O(gate784inter6));
  inv1  gate1630(.a(N2661), .O(gate784inter7));
  inv1  gate1631(.a(N546), .O(gate784inter8));
  nand2 gate1632(.a(gate784inter8), .b(gate784inter7), .O(gate784inter9));
  nand2 gate1633(.a(s_107), .b(gate784inter3), .O(gate784inter10));
  nor2  gate1634(.a(gate784inter10), .b(gate784inter9), .O(gate784inter11));
  nor2  gate1635(.a(gate784inter11), .b(gate784inter6), .O(gate784inter12));
  nand2 gate1636(.a(gate784inter12), .b(gate784inter1), .O(N2739));
inv1 gate785( .a(N2661), .O(N2740) );
nand2 gate786( .a(N2664), .b(N547), .O(N2741) );
inv1 gate787( .a(N2664), .O(N2742) );

  xor2  gate895(.a(N2689), .b(N385), .O(gate788inter0));
  nand2 gate896(.a(gate788inter0), .b(s_2), .O(gate788inter1));
  and2  gate897(.a(N2689), .b(N385), .O(gate788inter2));
  inv1  gate898(.a(s_2), .O(gate788inter3));
  inv1  gate899(.a(s_3), .O(gate788inter4));
  nand2 gate900(.a(gate788inter4), .b(gate788inter3), .O(gate788inter5));
  nor2  gate901(.a(gate788inter5), .b(gate788inter2), .O(gate788inter6));
  inv1  gate902(.a(N385), .O(gate788inter7));
  inv1  gate903(.a(N2689), .O(gate788inter8));
  nand2 gate904(.a(gate788inter8), .b(gate788inter7), .O(gate788inter9));
  nand2 gate905(.a(s_3), .b(gate788inter3), .O(gate788inter10));
  nor2  gate906(.a(gate788inter10), .b(gate788inter9), .O(gate788inter11));
  nor2  gate907(.a(gate788inter11), .b(gate788inter6), .O(gate788inter12));
  nand2 gate908(.a(gate788inter12), .b(gate788inter1), .O(N2743));
nand2 gate789( .a(N388), .b(N2691), .O(N2744) );
nand8 gate790( .a(N2537), .b(N2540), .c(N2543), .d(N2546), .e(N2594), .f(N2597), .g(N2600), .h(N2603), .O(N2745) );
nand8 gate791( .a(N2606), .b(N2549), .c(N2611), .d(N2614), .e(N2617), .f(N2620), .g(N2552), .h(N2555), .O(N2746) );
and8 gate792( .a(N2537), .b(N2540), .c(N2543), .d(N2546), .e(N2594), .f(N2597), .g(N2600), .h(N2603), .O(N2747) );
and8 gate793( .a(N2606), .b(N2549), .c(N2611), .d(N2614), .e(N2617), .f(N2620), .g(N2552), .h(N2555), .O(N2750) );
nand2 gate794( .a(N2669), .b(N2720), .O(N2753) );
nand2 gate795( .a(N2671), .b(N2721), .O(N2754) );
nand2 gate796( .a(N2673), .b(N2722), .O(N2755) );
nand2 gate797( .a(N2675), .b(N2723), .O(N2756) );
nand2 gate798( .a(N355), .b(N2725), .O(N2757) );

  xor2  gate1105(.a(N2727), .b(N358), .O(gate799inter0));
  nand2 gate1106(.a(gate799inter0), .b(s_32), .O(gate799inter1));
  and2  gate1107(.a(N2727), .b(N358), .O(gate799inter2));
  inv1  gate1108(.a(s_32), .O(gate799inter3));
  inv1  gate1109(.a(s_33), .O(gate799inter4));
  nand2 gate1110(.a(gate799inter4), .b(gate799inter3), .O(gate799inter5));
  nor2  gate1111(.a(gate799inter5), .b(gate799inter2), .O(gate799inter6));
  inv1  gate1112(.a(N358), .O(gate799inter7));
  inv1  gate1113(.a(N2727), .O(gate799inter8));
  nand2 gate1114(.a(gate799inter8), .b(gate799inter7), .O(gate799inter9));
  nand2 gate1115(.a(s_33), .b(gate799inter3), .O(gate799inter10));
  nor2  gate1116(.a(gate799inter10), .b(gate799inter9), .O(gate799inter11));
  nor2  gate1117(.a(gate799inter11), .b(gate799inter6), .O(gate799inter12));
  nand2 gate1118(.a(gate799inter12), .b(gate799inter1), .O(N2758));
nand2 gate800( .a(N361), .b(N2729), .O(N2759) );
nand2 gate801( .a(N364), .b(N2731), .O(N2760) );
nand2 gate802( .a(N367), .b(N2733), .O(N2761) );
nand2 gate803( .a(N2682), .b(N2734), .O(N2762) );
nand2 gate804( .a(N373), .b(N2736), .O(N2763) );
nand2 gate805( .a(N376), .b(N2738), .O(N2764) );
nand2 gate806( .a(N379), .b(N2740), .O(N2765) );
nand2 gate807( .a(N382), .b(N2742), .O(N2766) );
nand2 gate808( .a(N2688), .b(N2743), .O(N2767) );

  xor2  gate1497(.a(N2744), .b(N2690), .O(gate809inter0));
  nand2 gate1498(.a(gate809inter0), .b(s_88), .O(gate809inter1));
  and2  gate1499(.a(N2744), .b(N2690), .O(gate809inter2));
  inv1  gate1500(.a(s_88), .O(gate809inter3));
  inv1  gate1501(.a(s_89), .O(gate809inter4));
  nand2 gate1502(.a(gate809inter4), .b(gate809inter3), .O(gate809inter5));
  nor2  gate1503(.a(gate809inter5), .b(gate809inter2), .O(gate809inter6));
  inv1  gate1504(.a(N2690), .O(gate809inter7));
  inv1  gate1505(.a(N2744), .O(gate809inter8));
  nand2 gate1506(.a(gate809inter8), .b(gate809inter7), .O(gate809inter9));
  nand2 gate1507(.a(s_89), .b(gate809inter3), .O(gate809inter10));
  nor2  gate1508(.a(gate809inter10), .b(gate809inter9), .O(gate809inter11));
  nor2  gate1509(.a(gate809inter11), .b(gate809inter6), .O(gate809inter12));
  nand2 gate1510(.a(gate809inter12), .b(gate809inter1), .O(N2768));
and2 gate810( .a(N2745), .b(N275), .O(N2773) );
and2 gate811( .a(N2746), .b(N276), .O(N2776) );

  xor2  gate1637(.a(N2757), .b(N2724), .O(gate812inter0));
  nand2 gate1638(.a(gate812inter0), .b(s_108), .O(gate812inter1));
  and2  gate1639(.a(N2757), .b(N2724), .O(gate812inter2));
  inv1  gate1640(.a(s_108), .O(gate812inter3));
  inv1  gate1641(.a(s_109), .O(gate812inter4));
  nand2 gate1642(.a(gate812inter4), .b(gate812inter3), .O(gate812inter5));
  nor2  gate1643(.a(gate812inter5), .b(gate812inter2), .O(gate812inter6));
  inv1  gate1644(.a(N2724), .O(gate812inter7));
  inv1  gate1645(.a(N2757), .O(gate812inter8));
  nand2 gate1646(.a(gate812inter8), .b(gate812inter7), .O(gate812inter9));
  nand2 gate1647(.a(s_109), .b(gate812inter3), .O(gate812inter10));
  nor2  gate1648(.a(gate812inter10), .b(gate812inter9), .O(gate812inter11));
  nor2  gate1649(.a(gate812inter11), .b(gate812inter6), .O(gate812inter12));
  nand2 gate1650(.a(gate812inter12), .b(gate812inter1), .O(N2779));
nand2 gate813( .a(N2726), .b(N2758), .O(N2780) );
nand2 gate814( .a(N2728), .b(N2759), .O(N2781) );
nand2 gate815( .a(N2730), .b(N2760), .O(N2782) );

  xor2  gate1441(.a(N2761), .b(N2732), .O(gate816inter0));
  nand2 gate1442(.a(gate816inter0), .b(s_80), .O(gate816inter1));
  and2  gate1443(.a(N2761), .b(N2732), .O(gate816inter2));
  inv1  gate1444(.a(s_80), .O(gate816inter3));
  inv1  gate1445(.a(s_81), .O(gate816inter4));
  nand2 gate1446(.a(gate816inter4), .b(gate816inter3), .O(gate816inter5));
  nor2  gate1447(.a(gate816inter5), .b(gate816inter2), .O(gate816inter6));
  inv1  gate1448(.a(N2732), .O(gate816inter7));
  inv1  gate1449(.a(N2761), .O(gate816inter8));
  nand2 gate1450(.a(gate816inter8), .b(gate816inter7), .O(gate816inter9));
  nand2 gate1451(.a(s_81), .b(gate816inter3), .O(gate816inter10));
  nor2  gate1452(.a(gate816inter10), .b(gate816inter9), .O(gate816inter11));
  nor2  gate1453(.a(gate816inter11), .b(gate816inter6), .O(gate816inter12));
  nand2 gate1454(.a(gate816inter12), .b(gate816inter1), .O(N2783));
nand2 gate817( .a(N2735), .b(N2763), .O(N2784) );
nand2 gate818( .a(N2737), .b(N2764), .O(N2785) );

  xor2  gate1301(.a(N2765), .b(N2739), .O(gate819inter0));
  nand2 gate1302(.a(gate819inter0), .b(s_60), .O(gate819inter1));
  and2  gate1303(.a(N2765), .b(N2739), .O(gate819inter2));
  inv1  gate1304(.a(s_60), .O(gate819inter3));
  inv1  gate1305(.a(s_61), .O(gate819inter4));
  nand2 gate1306(.a(gate819inter4), .b(gate819inter3), .O(gate819inter5));
  nor2  gate1307(.a(gate819inter5), .b(gate819inter2), .O(gate819inter6));
  inv1  gate1308(.a(N2739), .O(gate819inter7));
  inv1  gate1309(.a(N2765), .O(gate819inter8));
  nand2 gate1310(.a(gate819inter8), .b(gate819inter7), .O(gate819inter9));
  nand2 gate1311(.a(s_61), .b(gate819inter3), .O(gate819inter10));
  nor2  gate1312(.a(gate819inter10), .b(gate819inter9), .O(gate819inter11));
  nor2  gate1313(.a(gate819inter11), .b(gate819inter6), .O(gate819inter12));
  nand2 gate1314(.a(gate819inter12), .b(gate819inter1), .O(N2786));
nand2 gate820( .a(N2741), .b(N2766), .O(N2787) );
and3 gate821( .a(N2747), .b(N2750), .c(N2710), .O(N2788) );

  xor2  gate2197(.a(N2750), .b(N2747), .O(gate822inter0));
  nand2 gate2198(.a(gate822inter0), .b(s_188), .O(gate822inter1));
  and2  gate2199(.a(N2750), .b(N2747), .O(gate822inter2));
  inv1  gate2200(.a(s_188), .O(gate822inter3));
  inv1  gate2201(.a(s_189), .O(gate822inter4));
  nand2 gate2202(.a(gate822inter4), .b(gate822inter3), .O(gate822inter5));
  nor2  gate2203(.a(gate822inter5), .b(gate822inter2), .O(gate822inter6));
  inv1  gate2204(.a(N2747), .O(gate822inter7));
  inv1  gate2205(.a(N2750), .O(gate822inter8));
  nand2 gate2206(.a(gate822inter8), .b(gate822inter7), .O(gate822inter9));
  nand2 gate2207(.a(s_189), .b(gate822inter3), .O(gate822inter10));
  nor2  gate2208(.a(gate822inter10), .b(gate822inter9), .O(gate822inter11));
  nor2  gate2209(.a(gate822inter11), .b(gate822inter6), .O(gate822inter12));
  nand2 gate2210(.a(gate822inter12), .b(gate822inter1), .O(N2789));
and4 gate823( .a(N338), .b(N2279), .c(N99), .d(N2788), .O(N2800) );

  xor2  gate1259(.a(N2018), .b(N2773), .O(gate824inter0));
  nand2 gate1260(.a(gate824inter0), .b(s_54), .O(gate824inter1));
  and2  gate1261(.a(N2018), .b(N2773), .O(gate824inter2));
  inv1  gate1262(.a(s_54), .O(gate824inter3));
  inv1  gate1263(.a(s_55), .O(gate824inter4));
  nand2 gate1264(.a(gate824inter4), .b(gate824inter3), .O(gate824inter5));
  nor2  gate1265(.a(gate824inter5), .b(gate824inter2), .O(gate824inter6));
  inv1  gate1266(.a(N2773), .O(gate824inter7));
  inv1  gate1267(.a(N2018), .O(gate824inter8));
  nand2 gate1268(.a(gate824inter8), .b(gate824inter7), .O(gate824inter9));
  nand2 gate1269(.a(s_55), .b(gate824inter3), .O(gate824inter10));
  nor2  gate1270(.a(gate824inter10), .b(gate824inter9), .O(gate824inter11));
  nor2  gate1271(.a(gate824inter11), .b(gate824inter6), .O(gate824inter12));
  nand2 gate1272(.a(gate824inter12), .b(gate824inter1), .O(N2807));
inv1 gate825( .a(N2773), .O(N2808) );

  xor2  gate1861(.a(N2019), .b(N2776), .O(gate826inter0));
  nand2 gate1862(.a(gate826inter0), .b(s_140), .O(gate826inter1));
  and2  gate1863(.a(N2019), .b(N2776), .O(gate826inter2));
  inv1  gate1864(.a(s_140), .O(gate826inter3));
  inv1  gate1865(.a(s_141), .O(gate826inter4));
  nand2 gate1866(.a(gate826inter4), .b(gate826inter3), .O(gate826inter5));
  nor2  gate1867(.a(gate826inter5), .b(gate826inter2), .O(gate826inter6));
  inv1  gate1868(.a(N2776), .O(gate826inter7));
  inv1  gate1869(.a(N2019), .O(gate826inter8));
  nand2 gate1870(.a(gate826inter8), .b(gate826inter7), .O(gate826inter9));
  nand2 gate1871(.a(s_141), .b(gate826inter3), .O(gate826inter10));
  nor2  gate1872(.a(gate826inter10), .b(gate826inter9), .O(gate826inter11));
  nor2  gate1873(.a(gate826inter11), .b(gate826inter6), .O(gate826inter12));
  nand2 gate1874(.a(gate826inter12), .b(gate826inter1), .O(N2809));
inv1 gate827( .a(N2776), .O(N2810) );
nor2 gate828( .a(N2384), .b(N2800), .O(N2811) );
and3 gate829( .a(N897), .b(N283), .c(N2789), .O(N2812) );
and3 gate830( .a(N76), .b(N283), .c(N2789), .O(N2815) );
and3 gate831( .a(N82), .b(N283), .c(N2789), .O(N2818) );
and3 gate832( .a(N85), .b(N283), .c(N2789), .O(N2821) );
and3 gate833( .a(N898), .b(N283), .c(N2789), .O(N2824) );
nand2 gate834( .a(N1965), .b(N2808), .O(N2827) );

  xor2  gate2029(.a(N2810), .b(N1968), .O(gate835inter0));
  nand2 gate2030(.a(gate835inter0), .b(s_164), .O(gate835inter1));
  and2  gate2031(.a(N2810), .b(N1968), .O(gate835inter2));
  inv1  gate2032(.a(s_164), .O(gate835inter3));
  inv1  gate2033(.a(s_165), .O(gate835inter4));
  nand2 gate2034(.a(gate835inter4), .b(gate835inter3), .O(gate835inter5));
  nor2  gate2035(.a(gate835inter5), .b(gate835inter2), .O(gate835inter6));
  inv1  gate2036(.a(N1968), .O(gate835inter7));
  inv1  gate2037(.a(N2810), .O(gate835inter8));
  nand2 gate2038(.a(gate835inter8), .b(gate835inter7), .O(gate835inter9));
  nand2 gate2039(.a(s_165), .b(gate835inter3), .O(gate835inter10));
  nor2  gate2040(.a(gate835inter10), .b(gate835inter9), .O(gate835inter11));
  nor2  gate2041(.a(gate835inter11), .b(gate835inter6), .O(gate835inter12));
  nand2 gate2042(.a(gate835inter12), .b(gate835inter1), .O(N2828));
and3 gate836( .a(N79), .b(N283), .c(N2789), .O(N2829) );
nand2 gate837( .a(N2807), .b(N2827), .O(N2843) );
nand2 gate838( .a(N2809), .b(N2828), .O(N2846) );

  xor2  gate1987(.a(N2076), .b(N2812), .O(gate839inter0));
  nand2 gate1988(.a(gate839inter0), .b(s_158), .O(gate839inter1));
  and2  gate1989(.a(N2076), .b(N2812), .O(gate839inter2));
  inv1  gate1990(.a(s_158), .O(gate839inter3));
  inv1  gate1991(.a(s_159), .O(gate839inter4));
  nand2 gate1992(.a(gate839inter4), .b(gate839inter3), .O(gate839inter5));
  nor2  gate1993(.a(gate839inter5), .b(gate839inter2), .O(gate839inter6));
  inv1  gate1994(.a(N2812), .O(gate839inter7));
  inv1  gate1995(.a(N2076), .O(gate839inter8));
  nand2 gate1996(.a(gate839inter8), .b(gate839inter7), .O(gate839inter9));
  nand2 gate1997(.a(s_159), .b(gate839inter3), .O(gate839inter10));
  nor2  gate1998(.a(gate839inter10), .b(gate839inter9), .O(gate839inter11));
  nor2  gate1999(.a(gate839inter11), .b(gate839inter6), .O(gate839inter12));
  nand2 gate2000(.a(gate839inter12), .b(gate839inter1), .O(N2850));

  xor2  gate1777(.a(N2077), .b(N2815), .O(gate840inter0));
  nand2 gate1778(.a(gate840inter0), .b(s_128), .O(gate840inter1));
  and2  gate1779(.a(N2077), .b(N2815), .O(gate840inter2));
  inv1  gate1780(.a(s_128), .O(gate840inter3));
  inv1  gate1781(.a(s_129), .O(gate840inter4));
  nand2 gate1782(.a(gate840inter4), .b(gate840inter3), .O(gate840inter5));
  nor2  gate1783(.a(gate840inter5), .b(gate840inter2), .O(gate840inter6));
  inv1  gate1784(.a(N2815), .O(gate840inter7));
  inv1  gate1785(.a(N2077), .O(gate840inter8));
  nand2 gate1786(.a(gate840inter8), .b(gate840inter7), .O(gate840inter9));
  nand2 gate1787(.a(s_129), .b(gate840inter3), .O(gate840inter10));
  nor2  gate1788(.a(gate840inter10), .b(gate840inter9), .O(gate840inter11));
  nor2  gate1789(.a(gate840inter11), .b(gate840inter6), .O(gate840inter12));
  nand2 gate1790(.a(gate840inter12), .b(gate840inter1), .O(N2851));
nand2 gate841( .a(N2818), .b(N1915), .O(N2852) );
nand2 gate842( .a(N2821), .b(N1857), .O(N2853) );

  xor2  gate1161(.a(N1938), .b(N2824), .O(gate843inter0));
  nand2 gate1162(.a(gate843inter0), .b(s_40), .O(gate843inter1));
  and2  gate1163(.a(N1938), .b(N2824), .O(gate843inter2));
  inv1  gate1164(.a(s_40), .O(gate843inter3));
  inv1  gate1165(.a(s_41), .O(gate843inter4));
  nand2 gate1166(.a(gate843inter4), .b(gate843inter3), .O(gate843inter5));
  nor2  gate1167(.a(gate843inter5), .b(gate843inter2), .O(gate843inter6));
  inv1  gate1168(.a(N2824), .O(gate843inter7));
  inv1  gate1169(.a(N1938), .O(gate843inter8));
  nand2 gate1170(.a(gate843inter8), .b(gate843inter7), .O(gate843inter9));
  nand2 gate1171(.a(s_41), .b(gate843inter3), .O(gate843inter10));
  nor2  gate1172(.a(gate843inter10), .b(gate843inter9), .O(gate843inter11));
  nor2  gate1173(.a(gate843inter11), .b(gate843inter6), .O(gate843inter12));
  nand2 gate1174(.a(gate843inter12), .b(gate843inter1), .O(N2854));
inv1 gate844( .a(N2812), .O(N2857) );
inv1 gate845( .a(N2815), .O(N2858) );
inv1 gate846( .a(N2818), .O(N2859) );
inv1 gate847( .a(N2821), .O(N2860) );
inv1 gate848( .a(N2824), .O(N2861) );
inv1 gate849( .a(N2829), .O(N2862) );
nand2 gate850( .a(N2829), .b(N1985), .O(N2863) );
nand2 gate851( .a(N2052), .b(N2857), .O(N2866) );
nand2 gate852( .a(N2055), .b(N2858), .O(N2867) );

  xor2  gate1329(.a(N2859), .b(N1866), .O(gate853inter0));
  nand2 gate1330(.a(gate853inter0), .b(s_64), .O(gate853inter1));
  and2  gate1331(.a(N2859), .b(N1866), .O(gate853inter2));
  inv1  gate1332(.a(s_64), .O(gate853inter3));
  inv1  gate1333(.a(s_65), .O(gate853inter4));
  nand2 gate1334(.a(gate853inter4), .b(gate853inter3), .O(gate853inter5));
  nor2  gate1335(.a(gate853inter5), .b(gate853inter2), .O(gate853inter6));
  inv1  gate1336(.a(N1866), .O(gate853inter7));
  inv1  gate1337(.a(N2859), .O(gate853inter8));
  nand2 gate1338(.a(gate853inter8), .b(gate853inter7), .O(gate853inter9));
  nand2 gate1339(.a(s_65), .b(gate853inter3), .O(gate853inter10));
  nor2  gate1340(.a(gate853inter10), .b(gate853inter9), .O(gate853inter11));
  nor2  gate1341(.a(gate853inter11), .b(gate853inter6), .O(gate853inter12));
  nand2 gate1342(.a(gate853inter12), .b(gate853inter1), .O(N2868));
nand2 gate854( .a(N1818), .b(N2860), .O(N2869) );
nand2 gate855( .a(N1902), .b(N2861), .O(N2870) );

  xor2  gate1973(.a(N886), .b(N2843), .O(gate856inter0));
  nand2 gate1974(.a(gate856inter0), .b(s_156), .O(gate856inter1));
  and2  gate1975(.a(N886), .b(N2843), .O(gate856inter2));
  inv1  gate1976(.a(s_156), .O(gate856inter3));
  inv1  gate1977(.a(s_157), .O(gate856inter4));
  nand2 gate1978(.a(gate856inter4), .b(gate856inter3), .O(gate856inter5));
  nor2  gate1979(.a(gate856inter5), .b(gate856inter2), .O(gate856inter6));
  inv1  gate1980(.a(N2843), .O(gate856inter7));
  inv1  gate1981(.a(N886), .O(gate856inter8));
  nand2 gate1982(.a(gate856inter8), .b(gate856inter7), .O(gate856inter9));
  nand2 gate1983(.a(s_157), .b(gate856inter3), .O(gate856inter10));
  nor2  gate1984(.a(gate856inter10), .b(gate856inter9), .O(gate856inter11));
  nor2  gate1985(.a(gate856inter11), .b(gate856inter6), .O(gate856inter12));
  nand2 gate1986(.a(gate856inter12), .b(gate856inter1), .O(N2871));
inv1 gate857( .a(N2843), .O(N2872) );
nand2 gate858( .a(N2846), .b(N887), .O(N2873) );
inv1 gate859( .a(N2846), .O(N2874) );
nand2 gate860( .a(N1933), .b(N2862), .O(N2875) );
nand2 gate861( .a(N2866), .b(N2850), .O(N2876) );

  xor2  gate1133(.a(N2851), .b(N2867), .O(gate862inter0));
  nand2 gate1134(.a(gate862inter0), .b(s_36), .O(gate862inter1));
  and2  gate1135(.a(N2851), .b(N2867), .O(gate862inter2));
  inv1  gate1136(.a(s_36), .O(gate862inter3));
  inv1  gate1137(.a(s_37), .O(gate862inter4));
  nand2 gate1138(.a(gate862inter4), .b(gate862inter3), .O(gate862inter5));
  nor2  gate1139(.a(gate862inter5), .b(gate862inter2), .O(gate862inter6));
  inv1  gate1140(.a(N2867), .O(gate862inter7));
  inv1  gate1141(.a(N2851), .O(gate862inter8));
  nand2 gate1142(.a(gate862inter8), .b(gate862inter7), .O(gate862inter9));
  nand2 gate1143(.a(s_37), .b(gate862inter3), .O(gate862inter10));
  nor2  gate1144(.a(gate862inter10), .b(gate862inter9), .O(gate862inter11));
  nor2  gate1145(.a(gate862inter11), .b(gate862inter6), .O(gate862inter12));
  nand2 gate1146(.a(gate862inter12), .b(gate862inter1), .O(N2877));
nand2 gate863( .a(N2868), .b(N2852), .O(N2878) );
nand2 gate864( .a(N2869), .b(N2853), .O(N2879) );

  xor2  gate2309(.a(N2854), .b(N2870), .O(gate865inter0));
  nand2 gate2310(.a(gate865inter0), .b(s_204), .O(gate865inter1));
  and2  gate2311(.a(N2854), .b(N2870), .O(gate865inter2));
  inv1  gate2312(.a(s_204), .O(gate865inter3));
  inv1  gate2313(.a(s_205), .O(gate865inter4));
  nand2 gate2314(.a(gate865inter4), .b(gate865inter3), .O(gate865inter5));
  nor2  gate2315(.a(gate865inter5), .b(gate865inter2), .O(gate865inter6));
  inv1  gate2316(.a(N2870), .O(gate865inter7));
  inv1  gate2317(.a(N2854), .O(gate865inter8));
  nand2 gate2318(.a(gate865inter8), .b(gate865inter7), .O(gate865inter9));
  nand2 gate2319(.a(s_205), .b(gate865inter3), .O(gate865inter10));
  nor2  gate2320(.a(gate865inter10), .b(gate865inter9), .O(gate865inter11));
  nor2  gate2321(.a(gate865inter11), .b(gate865inter6), .O(gate865inter12));
  nand2 gate2322(.a(gate865inter12), .b(gate865inter1), .O(N2880));
nand2 gate866( .a(N682), .b(N2872), .O(N2881) );
nand2 gate867( .a(N685), .b(N2874), .O(N2882) );
nand2 gate868( .a(N2875), .b(N2863), .O(N2883) );
and2 gate869( .a(N2876), .b(N550), .O(N2886) );
and2 gate870( .a(N551), .b(N2877), .O(N2887) );
and2 gate871( .a(N553), .b(N2878), .O(N2888) );
and2 gate872( .a(N2879), .b(N554), .O(N2889) );
and2 gate873( .a(N555), .b(N2880), .O(N2890) );

  xor2  gate1147(.a(N2881), .b(N2871), .O(gate874inter0));
  nand2 gate1148(.a(gate874inter0), .b(s_38), .O(gate874inter1));
  and2  gate1149(.a(N2881), .b(N2871), .O(gate874inter2));
  inv1  gate1150(.a(s_38), .O(gate874inter3));
  inv1  gate1151(.a(s_39), .O(gate874inter4));
  nand2 gate1152(.a(gate874inter4), .b(gate874inter3), .O(gate874inter5));
  nor2  gate1153(.a(gate874inter5), .b(gate874inter2), .O(gate874inter6));
  inv1  gate1154(.a(N2871), .O(gate874inter7));
  inv1  gate1155(.a(N2881), .O(gate874inter8));
  nand2 gate1156(.a(gate874inter8), .b(gate874inter7), .O(gate874inter9));
  nand2 gate1157(.a(s_39), .b(gate874inter3), .O(gate874inter10));
  nor2  gate1158(.a(gate874inter10), .b(gate874inter9), .O(gate874inter11));
  nor2  gate1159(.a(gate874inter11), .b(gate874inter6), .O(gate874inter12));
  nand2 gate1160(.a(gate874inter12), .b(gate874inter1), .O(N2891));
nand2 gate875( .a(N2873), .b(N2882), .O(N2892) );

  xor2  gate2085(.a(N1461), .b(N2883), .O(gate876inter0));
  nand2 gate2086(.a(gate876inter0), .b(s_172), .O(gate876inter1));
  and2  gate2087(.a(N1461), .b(N2883), .O(gate876inter2));
  inv1  gate2088(.a(s_172), .O(gate876inter3));
  inv1  gate2089(.a(s_173), .O(gate876inter4));
  nand2 gate2090(.a(gate876inter4), .b(gate876inter3), .O(gate876inter5));
  nor2  gate2091(.a(gate876inter5), .b(gate876inter2), .O(gate876inter6));
  inv1  gate2092(.a(N2883), .O(gate876inter7));
  inv1  gate2093(.a(N1461), .O(gate876inter8));
  nand2 gate2094(.a(gate876inter8), .b(gate876inter7), .O(gate876inter9));
  nand2 gate2095(.a(s_173), .b(gate876inter3), .O(gate876inter10));
  nor2  gate2096(.a(gate876inter10), .b(gate876inter9), .O(gate876inter11));
  nor2  gate2097(.a(gate876inter11), .b(gate876inter6), .O(gate876inter12));
  nand2 gate2098(.a(gate876inter12), .b(gate876inter1), .O(N2895));
inv1 gate877( .a(N2883), .O(N2896) );
nand2 gate878( .a(N1383), .b(N2896), .O(N2897) );
nand2 gate879( .a(N2895), .b(N2897), .O(N2898) );
and2 gate880( .a(N2898), .b(N552), .O(N2899) );

endmodule