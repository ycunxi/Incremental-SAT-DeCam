module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);

input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;//RE__PI;

input s_0,s_1;//RE__ALLOW(00,01,10,11);
input s_2,s_3;//RE__ALLOW(00,01,10,11);
input s_4,s_5;//RE__ALLOW(00,01,10,11);
input s_6,s_7;//RE__ALLOW(00,01,10,11);
input s_8,s_9;//RE__ALLOW(00,01,10,11);
input s_10,s_11;//RE__ALLOW(00,01,10,11);
input s_12,s_13;//RE__ALLOW(00,01,10,11);
input s_14,s_15;//RE__ALLOW(00,01,10,11);
input s_16,s_17;//RE__ALLOW(00,01,10,11);
input s_18,s_19;//RE__ALLOW(00,01,10,11);
input s_20,s_21;//RE__ALLOW(00,01,10,11);
input s_22,s_23;//RE__ALLOW(00,01,10,11);
input s_24,s_25;//RE__ALLOW(00,01,10,11);
input s_26,s_27;//RE__ALLOW(00,01,10,11);
input s_28,s_29;//RE__ALLOW(00,01,10,11);
input s_30,s_31;//RE__ALLOW(00,01,10,11);
input s_32,s_33;//RE__ALLOW(00,01,10,11);
input s_34,s_35;//RE__ALLOW(00,01,10,11);
input s_36,s_37;//RE__ALLOW(00,01,10,11);
input s_38,s_39;//RE__ALLOW(00,01,10,11);
input s_40,s_41;//RE__ALLOW(00,01,10,11);
input s_42,s_43;//RE__ALLOW(00,01,10,11);
input s_44,s_45;//RE__ALLOW(00,01,10,11);
input s_46,s_47;//RE__ALLOW(00,01,10,11);
input s_48,s_49;//RE__ALLOW(00,01,10,11);
input s_50,s_51;//RE__ALLOW(00,01,10,11);
input s_52,s_53;//RE__ALLOW(00,01,10,11);
input s_54,s_55;//RE__ALLOW(00,01,10,11);
input s_56,s_57;//RE__ALLOW(00,01,10,11);
input s_58,s_59;//RE__ALLOW(00,01,10,11);
input s_60,s_61;//RE__ALLOW(00,01,10,11);
input s_62,s_63;//RE__ALLOW(00,01,10,11);
input s_64,s_65;//RE__ALLOW(00,01,10,11);
input s_66,s_67;//RE__ALLOW(00,01,10,11);
input s_68,s_69;//RE__ALLOW(00,01,10,11);
input s_70,s_71;//RE__ALLOW(00,01,10,11);
input s_72,s_73;//RE__ALLOW(00,01,10,11);
input s_74,s_75;//RE__ALLOW(00,01,10,11);
input s_76,s_77;//RE__ALLOW(00,01,10,11);
input s_78,s_79;//RE__ALLOW(00,01,10,11);
input s_80,s_81;//RE__ALLOW(00,01,10,11);
input s_82,s_83;//RE__ALLOW(00,01,10,11);
input s_84,s_85;//RE__ALLOW(00,01,10,11);
input s_86,s_87;//RE__ALLOW(00,01,10,11);
input s_88,s_89;//RE__ALLOW(00,01,10,11);
input s_90,s_91;//RE__ALLOW(00,01,10,11);
input s_92,s_93;//RE__ALLOW(00,01,10,11);
input s_94,s_95;//RE__ALLOW(00,01,10,11);
input s_96,s_97;//RE__ALLOW(00,01,10,11);
input s_98,s_99;//RE__ALLOW(00,01,10,11);
input s_100,s_101;//RE__ALLOW(00,01,10,11);
input s_102,s_103;//RE__ALLOW(00,01,10,11);
input s_104,s_105;//RE__ALLOW(00,01,10,11);
input s_106,s_107;//RE__ALLOW(00,01,10,11);
input s_108,s_109;//RE__ALLOW(00,01,10,11);
input s_110,s_111;//RE__ALLOW(00,01,10,11);
input s_112,s_113;//RE__ALLOW(00,01,10,11);
input s_114,s_115;//RE__ALLOW(00,01,10,11);
input s_116,s_117;//RE__ALLOW(00,01,10,11);
input s_118,s_119;//RE__ALLOW(00,01,10,11);
input s_120,s_121;//RE__ALLOW(00,01,10,11);
input s_122,s_123;//RE__ALLOW(00,01,10,11);
input s_124,s_125;//RE__ALLOW(00,01,10,11);
input s_126,s_127;//RE__ALLOW(00,01,10,11);
input s_128,s_129;//RE__ALLOW(00,01,10,11);
input s_130,s_131;//RE__ALLOW(00,01,10,11);
input s_132,s_133;//RE__ALLOW(00,01,10,11);
input s_134,s_135;//RE__ALLOW(00,01,10,11);
input s_136,s_137;//RE__ALLOW(00,01,10,11);
input s_138,s_139;//RE__ALLOW(00,01,10,11);
input s_140,s_141;//RE__ALLOW(00,01,10,11);
input s_142,s_143;//RE__ALLOW(00,01,10,11);
input s_144,s_145;//RE__ALLOW(00,01,10,11);
input s_146,s_147;//RE__ALLOW(00,01,10,11);
input s_148,s_149;//RE__ALLOW(00,01,10,11);
input s_150,s_151;//RE__ALLOW(00,01,10,11);
input s_152,s_153;//RE__ALLOW(00,01,10,11);
input s_154,s_155;//RE__ALLOW(00,01,10,11);
input s_156,s_157;//RE__ALLOW(00,01,10,11);
input s_158,s_159;//RE__ALLOW(00,01,10,11);
input s_160,s_161;//RE__ALLOW(00,01,10,11);
input s_162,s_163;//RE__ALLOW(00,01,10,11);
input s_164,s_165;//RE__ALLOW(00,01,10,11);
input s_166,s_167;//RE__ALLOW(00,01,10,11);
input s_168,s_169;//RE__ALLOW(00,01,10,11);
input s_170,s_171;//RE__ALLOW(00,01,10,11);
input s_172,s_173;//RE__ALLOW(00,01,10,11);
input s_174,s_175;//RE__ALLOW(00,01,10,11);
input s_176,s_177;//RE__ALLOW(00,01,10,11);
input s_178,s_179;//RE__ALLOW(00,01,10,11);
input s_180,s_181;//RE__ALLOW(00,01,10,11);
input s_182,s_183;//RE__ALLOW(00,01,10,11);
input s_184,s_185;//RE__ALLOW(00,01,10,11);
input s_186,s_187;//RE__ALLOW(00,01,10,11);
input s_188,s_189;//RE__ALLOW(00,01,10,11);
input s_190,s_191;//RE__ALLOW(00,01,10,11);
input s_192,s_193;//RE__ALLOW(00,01,10,11);
input s_194,s_195;//RE__ALLOW(00,01,10,11);
input s_196,s_197;//RE__ALLOW(00,01,10,11);
input s_198,s_199;//RE__ALLOW(00,01,10,11);
input s_200,s_201;//RE__ALLOW(00,01,10,11);
input s_202,s_203;//RE__ALLOW(00,01,10,11);
input s_204,s_205;//RE__ALLOW(00,01,10,11);
input s_206,s_207;//RE__ALLOW(00,01,10,11);
input s_208,s_209;//RE__ALLOW(00,01,10,11);
input s_210,s_211;//RE__ALLOW(00,01,10,11);
input s_212,s_213;//RE__ALLOW(00,01,10,11);
input s_214,s_215;//RE__ALLOW(00,01,10,11);
input s_216,s_217;//RE__ALLOW(00,01,10,11);
input s_218,s_219;//RE__ALLOW(00,01,10,11);
input s_220,s_221;//RE__ALLOW(00,01,10,11);
input s_222,s_223;//RE__ALLOW(00,01,10,11);
input s_224,s_225;//RE__ALLOW(00,01,10,11);
input s_226,s_227;//RE__ALLOW(00,01,10,11);
input s_228,s_229;//RE__ALLOW(00,01,10,11);
input s_230,s_231;//RE__ALLOW(00,01,10,11);
input s_232,s_233;//RE__ALLOW(00,01,10,11);
input s_234,s_235;//RE__ALLOW(00,01,10,11);
input s_236,s_237;//RE__ALLOW(00,01,10,11);
input s_238,s_239;//RE__ALLOW(00,01,10,11);
input s_240,s_241;//RE__ALLOW(00,01,10,11);
input s_242,s_243;//RE__ALLOW(00,01,10,11);
input s_244,s_245;//RE__ALLOW(00,01,10,11);
input s_246,s_247;//RE__ALLOW(00,01,10,11);
input s_248,s_249;//RE__ALLOW(00,01,10,11);
input s_250,s_251;//RE__ALLOW(00,01,10,11);
input s_252,s_253;//RE__ALLOW(00,01,10,11);
input s_254,s_255;//RE__ALLOW(00,01,10,11);
input s_256,s_257;//RE__ALLOW(00,01,10,11);
input s_258,s_259;//RE__ALLOW(00,01,10,11);
input s_260,s_261;//RE__ALLOW(00,01,10,11);
input s_262,s_263;//RE__ALLOW(00,01,10,11);
input s_264,s_265;//RE__ALLOW(00,01,10,11);
input s_266,s_267;//RE__ALLOW(00,01,10,11);
input s_268,s_269;//RE__ALLOW(00,01,10,11);
input s_270,s_271;//RE__ALLOW(00,01,10,11);
input s_272,s_273;//RE__ALLOW(00,01,10,11);
input s_274,s_275;//RE__ALLOW(00,01,10,11);
input s_276,s_277;//RE__ALLOW(00,01,10,11);
input s_278,s_279;//RE__ALLOW(00,01,10,11);
input s_280,s_281;//RE__ALLOW(00,01,10,11);
input s_282,s_283;//RE__ALLOW(00,01,10,11);
input s_284,s_285;//RE__ALLOW(00,01,10,11);
input s_286,s_287;//RE__ALLOW(00,01,10,11);
input s_288,s_289;//RE__ALLOW(00,01,10,11);
input s_290,s_291;//RE__ALLOW(00,01,10,11);
input s_292,s_293;//RE__ALLOW(00,01,10,11);
input s_294,s_295;//RE__ALLOW(00,01,10,11);
input s_296,s_297;//RE__ALLOW(00,01,10,11);
input s_298,s_299;//RE__ALLOW(00,01,10,11);
input s_300,s_301;//RE__ALLOW(00,01,10,11);
input s_302,s_303;//RE__ALLOW(00,01,10,11);
input s_304,s_305;//RE__ALLOW(00,01,10,11);
input s_306,s_307;//RE__ALLOW(00,01,10,11);
input s_308,s_309;//RE__ALLOW(00,01,10,11);
input s_310,s_311;//RE__ALLOW(00,01,10,11);
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;

  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate45inter0, gate45inter1, gate45inter2, gate45inter3, gate45inter4, gate45inter5, gate45inter6, gate45inter7, gate45inter8, gate45inter9, gate45inter10, gate45inter11, gate45inter12, gate164inter0, gate164inter1, gate164inter2, gate164inter3, gate164inter4, gate164inter5, gate164inter6, gate164inter7, gate164inter8, gate164inter9, gate164inter10, gate164inter11, gate164inter12, gate503inter0, gate503inter1, gate503inter2, gate503inter3, gate503inter4, gate503inter5, gate503inter6, gate503inter7, gate503inter8, gate503inter9, gate503inter10, gate503inter11, gate503inter12, gate51inter0, gate51inter1, gate51inter2, gate51inter3, gate51inter4, gate51inter5, gate51inter6, gate51inter7, gate51inter8, gate51inter9, gate51inter10, gate51inter11, gate51inter12, gate387inter0, gate387inter1, gate387inter2, gate387inter3, gate387inter4, gate387inter5, gate387inter6, gate387inter7, gate387inter8, gate387inter9, gate387inter10, gate387inter11, gate387inter12, gate73inter0, gate73inter1, gate73inter2, gate73inter3, gate73inter4, gate73inter5, gate73inter6, gate73inter7, gate73inter8, gate73inter9, gate73inter10, gate73inter11, gate73inter12, gate58inter0, gate58inter1, gate58inter2, gate58inter3, gate58inter4, gate58inter5, gate58inter6, gate58inter7, gate58inter8, gate58inter9, gate58inter10, gate58inter11, gate58inter12, gate172inter0, gate172inter1, gate172inter2, gate172inter3, gate172inter4, gate172inter5, gate172inter6, gate172inter7, gate172inter8, gate172inter9, gate172inter10, gate172inter11, gate172inter12, gate86inter0, gate86inter1, gate86inter2, gate86inter3, gate86inter4, gate86inter5, gate86inter6, gate86inter7, gate86inter8, gate86inter9, gate86inter10, gate86inter11, gate86inter12, gate391inter0, gate391inter1, gate391inter2, gate391inter3, gate391inter4, gate391inter5, gate391inter6, gate391inter7, gate391inter8, gate391inter9, gate391inter10, gate391inter11, gate391inter12, gate226inter0, gate226inter1, gate226inter2, gate226inter3, gate226inter4, gate226inter5, gate226inter6, gate226inter7, gate226inter8, gate226inter9, gate226inter10, gate226inter11, gate226inter12, gate48inter0, gate48inter1, gate48inter2, gate48inter3, gate48inter4, gate48inter5, gate48inter6, gate48inter7, gate48inter8, gate48inter9, gate48inter10, gate48inter11, gate48inter12, gate106inter0, gate106inter1, gate106inter2, gate106inter3, gate106inter4, gate106inter5, gate106inter6, gate106inter7, gate106inter8, gate106inter9, gate106inter10, gate106inter11, gate106inter12, gate455inter0, gate455inter1, gate455inter2, gate455inter3, gate455inter4, gate455inter5, gate455inter6, gate455inter7, gate455inter8, gate455inter9, gate455inter10, gate455inter11, gate455inter12, gate239inter0, gate239inter1, gate239inter2, gate239inter3, gate239inter4, gate239inter5, gate239inter6, gate239inter7, gate239inter8, gate239inter9, gate239inter10, gate239inter11, gate239inter12, gate490inter0, gate490inter1, gate490inter2, gate490inter3, gate490inter4, gate490inter5, gate490inter6, gate490inter7, gate490inter8, gate490inter9, gate490inter10, gate490inter11, gate490inter12, gate417inter0, gate417inter1, gate417inter2, gate417inter3, gate417inter4, gate417inter5, gate417inter6, gate417inter7, gate417inter8, gate417inter9, gate417inter10, gate417inter11, gate417inter12, gate427inter0, gate427inter1, gate427inter2, gate427inter3, gate427inter4, gate427inter5, gate427inter6, gate427inter7, gate427inter8, gate427inter9, gate427inter10, gate427inter11, gate427inter12, gate56inter0, gate56inter1, gate56inter2, gate56inter3, gate56inter4, gate56inter5, gate56inter6, gate56inter7, gate56inter8, gate56inter9, gate56inter10, gate56inter11, gate56inter12, gate499inter0, gate499inter1, gate499inter2, gate499inter3, gate499inter4, gate499inter5, gate499inter6, gate499inter7, gate499inter8, gate499inter9, gate499inter10, gate499inter11, gate499inter12, gate115inter0, gate115inter1, gate115inter2, gate115inter3, gate115inter4, gate115inter5, gate115inter6, gate115inter7, gate115inter8, gate115inter9, gate115inter10, gate115inter11, gate115inter12, gate228inter0, gate228inter1, gate228inter2, gate228inter3, gate228inter4, gate228inter5, gate228inter6, gate228inter7, gate228inter8, gate228inter9, gate228inter10, gate228inter11, gate228inter12, gate137inter0, gate137inter1, gate137inter2, gate137inter3, gate137inter4, gate137inter5, gate137inter6, gate137inter7, gate137inter8, gate137inter9, gate137inter10, gate137inter11, gate137inter12, gate53inter0, gate53inter1, gate53inter2, gate53inter3, gate53inter4, gate53inter5, gate53inter6, gate53inter7, gate53inter8, gate53inter9, gate53inter10, gate53inter11, gate53inter12, gate255inter0, gate255inter1, gate255inter2, gate255inter3, gate255inter4, gate255inter5, gate255inter6, gate255inter7, gate255inter8, gate255inter9, gate255inter10, gate255inter11, gate255inter12, gate388inter0, gate388inter1, gate388inter2, gate388inter3, gate388inter4, gate388inter5, gate388inter6, gate388inter7, gate388inter8, gate388inter9, gate388inter10, gate388inter11, gate388inter12, gate416inter0, gate416inter1, gate416inter2, gate416inter3, gate416inter4, gate416inter5, gate416inter6, gate416inter7, gate416inter8, gate416inter9, gate416inter10, gate416inter11, gate416inter12, gate408inter0, gate408inter1, gate408inter2, gate408inter3, gate408inter4, gate408inter5, gate408inter6, gate408inter7, gate408inter8, gate408inter9, gate408inter10, gate408inter11, gate408inter12, gate113inter0, gate113inter1, gate113inter2, gate113inter3, gate113inter4, gate113inter5, gate113inter6, gate113inter7, gate113inter8, gate113inter9, gate113inter10, gate113inter11, gate113inter12, gate473inter0, gate473inter1, gate473inter2, gate473inter3, gate473inter4, gate473inter5, gate473inter6, gate473inter7, gate473inter8, gate473inter9, gate473inter10, gate473inter11, gate473inter12, gate509inter0, gate509inter1, gate509inter2, gate509inter3, gate509inter4, gate509inter5, gate509inter6, gate509inter7, gate509inter8, gate509inter9, gate509inter10, gate509inter11, gate509inter12, gate111inter0, gate111inter1, gate111inter2, gate111inter3, gate111inter4, gate111inter5, gate111inter6, gate111inter7, gate111inter8, gate111inter9, gate111inter10, gate111inter11, gate111inter12, gate460inter0, gate460inter1, gate460inter2, gate460inter3, gate460inter4, gate460inter5, gate460inter6, gate460inter7, gate460inter8, gate460inter9, gate460inter10, gate460inter11, gate460inter12, gate83inter0, gate83inter1, gate83inter2, gate83inter3, gate83inter4, gate83inter5, gate83inter6, gate83inter7, gate83inter8, gate83inter9, gate83inter10, gate83inter11, gate83inter12, gate91inter0, gate91inter1, gate91inter2, gate91inter3, gate91inter4, gate91inter5, gate91inter6, gate91inter7, gate91inter8, gate91inter9, gate91inter10, gate91inter11, gate91inter12, gate98inter0, gate98inter1, gate98inter2, gate98inter3, gate98inter4, gate98inter5, gate98inter6, gate98inter7, gate98inter8, gate98inter9, gate98inter10, gate98inter11, gate98inter12, gate117inter0, gate117inter1, gate117inter2, gate117inter3, gate117inter4, gate117inter5, gate117inter6, gate117inter7, gate117inter8, gate117inter9, gate117inter10, gate117inter11, gate117inter12, gate394inter0, gate394inter1, gate394inter2, gate394inter3, gate394inter4, gate394inter5, gate394inter6, gate394inter7, gate394inter8, gate394inter9, gate394inter10, gate394inter11, gate394inter12, gate510inter0, gate510inter1, gate510inter2, gate510inter3, gate510inter4, gate510inter5, gate510inter6, gate510inter7, gate510inter8, gate510inter9, gate510inter10, gate510inter11, gate510inter12, gate188inter0, gate188inter1, gate188inter2, gate188inter3, gate188inter4, gate188inter5, gate188inter6, gate188inter7, gate188inter8, gate188inter9, gate188inter10, gate188inter11, gate188inter12, gate35inter0, gate35inter1, gate35inter2, gate35inter3, gate35inter4, gate35inter5, gate35inter6, gate35inter7, gate35inter8, gate35inter9, gate35inter10, gate35inter11, gate35inter12, gate174inter0, gate174inter1, gate174inter2, gate174inter3, gate174inter4, gate174inter5, gate174inter6, gate174inter7, gate174inter8, gate174inter9, gate174inter10, gate174inter11, gate174inter12, gate27inter0, gate27inter1, gate27inter2, gate27inter3, gate27inter4, gate27inter5, gate27inter6, gate27inter7, gate27inter8, gate27inter9, gate27inter10, gate27inter11, gate27inter12, gate119inter0, gate119inter1, gate119inter2, gate119inter3, gate119inter4, gate119inter5, gate119inter6, gate119inter7, gate119inter8, gate119inter9, gate119inter10, gate119inter11, gate119inter12, gate18inter0, gate18inter1, gate18inter2, gate18inter3, gate18inter4, gate18inter5, gate18inter6, gate18inter7, gate18inter8, gate18inter9, gate18inter10, gate18inter11, gate18inter12, gate225inter0, gate225inter1, gate225inter2, gate225inter3, gate225inter4, gate225inter5, gate225inter6, gate225inter7, gate225inter8, gate225inter9, gate225inter10, gate225inter11, gate225inter12, gate190inter0, gate190inter1, gate190inter2, gate190inter3, gate190inter4, gate190inter5, gate190inter6, gate190inter7, gate190inter8, gate190inter9, gate190inter10, gate190inter11, gate190inter12, gate153inter0, gate153inter1, gate153inter2, gate153inter3, gate153inter4, gate153inter5, gate153inter6, gate153inter7, gate153inter8, gate153inter9, gate153inter10, gate153inter11, gate153inter12, gate72inter0, gate72inter1, gate72inter2, gate72inter3, gate72inter4, gate72inter5, gate72inter6, gate72inter7, gate72inter8, gate72inter9, gate72inter10, gate72inter11, gate72inter12, gate59inter0, gate59inter1, gate59inter2, gate59inter3, gate59inter4, gate59inter5, gate59inter6, gate59inter7, gate59inter8, gate59inter9, gate59inter10, gate59inter11, gate59inter12, gate487inter0, gate487inter1, gate487inter2, gate487inter3, gate487inter4, gate487inter5, gate487inter6, gate487inter7, gate487inter8, gate487inter9, gate487inter10, gate487inter11, gate487inter12, gate511inter0, gate511inter1, gate511inter2, gate511inter3, gate511inter4, gate511inter5, gate511inter6, gate511inter7, gate511inter8, gate511inter9, gate511inter10, gate511inter11, gate511inter12, gate447inter0, gate447inter1, gate447inter2, gate447inter3, gate447inter4, gate447inter5, gate447inter6, gate447inter7, gate447inter8, gate447inter9, gate447inter10, gate447inter11, gate447inter12, gate476inter0, gate476inter1, gate476inter2, gate476inter3, gate476inter4, gate476inter5, gate476inter6, gate476inter7, gate476inter8, gate476inter9, gate476inter10, gate476inter11, gate476inter12, gate94inter0, gate94inter1, gate94inter2, gate94inter3, gate94inter4, gate94inter5, gate94inter6, gate94inter7, gate94inter8, gate94inter9, gate94inter10, gate94inter11, gate94inter12, gate469inter0, gate469inter1, gate469inter2, gate469inter3, gate469inter4, gate469inter5, gate469inter6, gate469inter7, gate469inter8, gate469inter9, gate469inter10, gate469inter11, gate469inter12, gate235inter0, gate235inter1, gate235inter2, gate235inter3, gate235inter4, gate235inter5, gate235inter6, gate235inter7, gate235inter8, gate235inter9, gate235inter10, gate235inter11, gate235inter12, gate206inter0, gate206inter1, gate206inter2, gate206inter3, gate206inter4, gate206inter5, gate206inter6, gate206inter7, gate206inter8, gate206inter9, gate206inter10, gate206inter11, gate206inter12, gate54inter0, gate54inter1, gate54inter2, gate54inter3, gate54inter4, gate54inter5, gate54inter6, gate54inter7, gate54inter8, gate54inter9, gate54inter10, gate54inter11, gate54inter12, gate265inter0, gate265inter1, gate265inter2, gate265inter3, gate265inter4, gate265inter5, gate265inter6, gate265inter7, gate265inter8, gate265inter9, gate265inter10, gate265inter11, gate265inter12, gate140inter0, gate140inter1, gate140inter2, gate140inter3, gate140inter4, gate140inter5, gate140inter6, gate140inter7, gate140inter8, gate140inter9, gate140inter10, gate140inter11, gate140inter12, gate100inter0, gate100inter1, gate100inter2, gate100inter3, gate100inter4, gate100inter5, gate100inter6, gate100inter7, gate100inter8, gate100inter9, gate100inter10, gate100inter11, gate100inter12, gate95inter0, gate95inter1, gate95inter2, gate95inter3, gate95inter4, gate95inter5, gate95inter6, gate95inter7, gate95inter8, gate95inter9, gate95inter10, gate95inter11, gate95inter12, gate389inter0, gate389inter1, gate389inter2, gate389inter3, gate389inter4, gate389inter5, gate389inter6, gate389inter7, gate389inter8, gate389inter9, gate389inter10, gate389inter11, gate389inter12, gate26inter0, gate26inter1, gate26inter2, gate26inter3, gate26inter4, gate26inter5, gate26inter6, gate26inter7, gate26inter8, gate26inter9, gate26inter10, gate26inter11, gate26inter12, gate245inter0, gate245inter1, gate245inter2, gate245inter3, gate245inter4, gate245inter5, gate245inter6, gate245inter7, gate245inter8, gate245inter9, gate245inter10, gate245inter11, gate245inter12, gate201inter0, gate201inter1, gate201inter2, gate201inter3, gate201inter4, gate201inter5, gate201inter6, gate201inter7, gate201inter8, gate201inter9, gate201inter10, gate201inter11, gate201inter12, gate183inter0, gate183inter1, gate183inter2, gate183inter3, gate183inter4, gate183inter5, gate183inter6, gate183inter7, gate183inter8, gate183inter9, gate183inter10, gate183inter11, gate183inter12, gate285inter0, gate285inter1, gate285inter2, gate285inter3, gate285inter4, gate285inter5, gate285inter6, gate285inter7, gate285inter8, gate285inter9, gate285inter10, gate285inter11, gate285inter12, gate293inter0, gate293inter1, gate293inter2, gate293inter3, gate293inter4, gate293inter5, gate293inter6, gate293inter7, gate293inter8, gate293inter9, gate293inter10, gate293inter11, gate293inter12, gate211inter0, gate211inter1, gate211inter2, gate211inter3, gate211inter4, gate211inter5, gate211inter6, gate211inter7, gate211inter8, gate211inter9, gate211inter10, gate211inter11, gate211inter12, gate456inter0, gate456inter1, gate456inter2, gate456inter3, gate456inter4, gate456inter5, gate456inter6, gate456inter7, gate456inter8, gate456inter9, gate456inter10, gate456inter11, gate456inter12, gate227inter0, gate227inter1, gate227inter2, gate227inter3, gate227inter4, gate227inter5, gate227inter6, gate227inter7, gate227inter8, gate227inter9, gate227inter10, gate227inter11, gate227inter12, gate409inter0, gate409inter1, gate409inter2, gate409inter3, gate409inter4, gate409inter5, gate409inter6, gate409inter7, gate409inter8, gate409inter9, gate409inter10, gate409inter11, gate409inter12, gate158inter0, gate158inter1, gate158inter2, gate158inter3, gate158inter4, gate158inter5, gate158inter6, gate158inter7, gate158inter8, gate158inter9, gate158inter10, gate158inter11, gate158inter12, gate185inter0, gate185inter1, gate185inter2, gate185inter3, gate185inter4, gate185inter5, gate185inter6, gate185inter7, gate185inter8, gate185inter9, gate185inter10, gate185inter11, gate185inter12, gate434inter0, gate434inter1, gate434inter2, gate434inter3, gate434inter4, gate434inter5, gate434inter6, gate434inter7, gate434inter8, gate434inter9, gate434inter10, gate434inter11, gate434inter12, gate97inter0, gate97inter1, gate97inter2, gate97inter3, gate97inter4, gate97inter5, gate97inter6, gate97inter7, gate97inter8, gate97inter9, gate97inter10, gate97inter11, gate97inter12, gate237inter0, gate237inter1, gate237inter2, gate237inter3, gate237inter4, gate237inter5, gate237inter6, gate237inter7, gate237inter8, gate237inter9, gate237inter10, gate237inter11, gate237inter12, gate261inter0, gate261inter1, gate261inter2, gate261inter3, gate261inter4, gate261inter5, gate261inter6, gate261inter7, gate261inter8, gate261inter9, gate261inter10, gate261inter11, gate261inter12, gate218inter0, gate218inter1, gate218inter2, gate218inter3, gate218inter4, gate218inter5, gate218inter6, gate218inter7, gate218inter8, gate218inter9, gate218inter10, gate218inter11, gate218inter12, gate223inter0, gate223inter1, gate223inter2, gate223inter3, gate223inter4, gate223inter5, gate223inter6, gate223inter7, gate223inter8, gate223inter9, gate223inter10, gate223inter11, gate223inter12, gate289inter0, gate289inter1, gate289inter2, gate289inter3, gate289inter4, gate289inter5, gate289inter6, gate289inter7, gate289inter8, gate289inter9, gate289inter10, gate289inter11, gate289inter12, gate399inter0, gate399inter1, gate399inter2, gate399inter3, gate399inter4, gate399inter5, gate399inter6, gate399inter7, gate399inter8, gate399inter9, gate399inter10, gate399inter11, gate399inter12, gate112inter0, gate112inter1, gate112inter2, gate112inter3, gate112inter4, gate112inter5, gate112inter6, gate112inter7, gate112inter8, gate112inter9, gate112inter10, gate112inter11, gate112inter12, gate425inter0, gate425inter1, gate425inter2, gate425inter3, gate425inter4, gate425inter5, gate425inter6, gate425inter7, gate425inter8, gate425inter9, gate425inter10, gate425inter11, gate425inter12, gate63inter0, gate63inter1, gate63inter2, gate63inter3, gate63inter4, gate63inter5, gate63inter6, gate63inter7, gate63inter8, gate63inter9, gate63inter10, gate63inter11, gate63inter12, gate123inter0, gate123inter1, gate123inter2, gate123inter3, gate123inter4, gate123inter5, gate123inter6, gate123inter7, gate123inter8, gate123inter9, gate123inter10, gate123inter11, gate123inter12, gate69inter0, gate69inter1, gate69inter2, gate69inter3, gate69inter4, gate69inter5, gate69inter6, gate69inter7, gate69inter8, gate69inter9, gate69inter10, gate69inter11, gate69inter12, gate214inter0, gate214inter1, gate214inter2, gate214inter3, gate214inter4, gate214inter5, gate214inter6, gate214inter7, gate214inter8, gate214inter9, gate214inter10, gate214inter11, gate214inter12, gate222inter0, gate222inter1, gate222inter2, gate222inter3, gate222inter4, gate222inter5, gate222inter6, gate222inter7, gate222inter8, gate222inter9, gate222inter10, gate222inter11, gate222inter12, gate291inter0, gate291inter1, gate291inter2, gate291inter3, gate291inter4, gate291inter5, gate291inter6, gate291inter7, gate291inter8, gate291inter9, gate291inter10, gate291inter11, gate291inter12, gate133inter0, gate133inter1, gate133inter2, gate133inter3, gate133inter4, gate133inter5, gate133inter6, gate133inter7, gate133inter8, gate133inter9, gate133inter10, gate133inter11, gate133inter12, gate431inter0, gate431inter1, gate431inter2, gate431inter3, gate431inter4, gate431inter5, gate431inter6, gate431inter7, gate431inter8, gate431inter9, gate431inter10, gate431inter11, gate431inter12, gate131inter0, gate131inter1, gate131inter2, gate131inter3, gate131inter4, gate131inter5, gate131inter6, gate131inter7, gate131inter8, gate131inter9, gate131inter10, gate131inter11, gate131inter12, gate210inter0, gate210inter1, gate210inter2, gate210inter3, gate210inter4, gate210inter5, gate210inter6, gate210inter7, gate210inter8, gate210inter9, gate210inter10, gate210inter11, gate210inter12, gate209inter0, gate209inter1, gate209inter2, gate209inter3, gate209inter4, gate209inter5, gate209inter6, gate209inter7, gate209inter8, gate209inter9, gate209inter10, gate209inter11, gate209inter12, gate196inter0, gate196inter1, gate196inter2, gate196inter3, gate196inter4, gate196inter5, gate196inter6, gate196inter7, gate196inter8, gate196inter9, gate196inter10, gate196inter11, gate196inter12, gate233inter0, gate233inter1, gate233inter2, gate233inter3, gate233inter4, gate233inter5, gate233inter6, gate233inter7, gate233inter8, gate233inter9, gate233inter10, gate233inter11, gate233inter12, gate254inter0, gate254inter1, gate254inter2, gate254inter3, gate254inter4, gate254inter5, gate254inter6, gate254inter7, gate254inter8, gate254inter9, gate254inter10, gate254inter11, gate254inter12, gate203inter0, gate203inter1, gate203inter2, gate203inter3, gate203inter4, gate203inter5, gate203inter6, gate203inter7, gate203inter8, gate203inter9, gate203inter10, gate203inter11, gate203inter12, gate396inter0, gate396inter1, gate396inter2, gate396inter3, gate396inter4, gate396inter5, gate396inter6, gate396inter7, gate396inter8, gate396inter9, gate396inter10, gate396inter11, gate396inter12, gate180inter0, gate180inter1, gate180inter2, gate180inter3, gate180inter4, gate180inter5, gate180inter6, gate180inter7, gate180inter8, gate180inter9, gate180inter10, gate180inter11, gate180inter12, gate464inter0, gate464inter1, gate464inter2, gate464inter3, gate464inter4, gate464inter5, gate464inter6, gate464inter7, gate464inter8, gate464inter9, gate464inter10, gate464inter11, gate464inter12, gate212inter0, gate212inter1, gate212inter2, gate212inter3, gate212inter4, gate212inter5, gate212inter6, gate212inter7, gate212inter8, gate212inter9, gate212inter10, gate212inter11, gate212inter12, gate20inter0, gate20inter1, gate20inter2, gate20inter3, gate20inter4, gate20inter5, gate20inter6, gate20inter7, gate20inter8, gate20inter9, gate20inter10, gate20inter11, gate20inter12, gate74inter0, gate74inter1, gate74inter2, gate74inter3, gate74inter4, gate74inter5, gate74inter6, gate74inter7, gate74inter8, gate74inter9, gate74inter10, gate74inter11, gate74inter12, gate286inter0, gate286inter1, gate286inter2, gate286inter3, gate286inter4, gate286inter5, gate286inter6, gate286inter7, gate286inter8, gate286inter9, gate286inter10, gate286inter11, gate286inter12, gate262inter0, gate262inter1, gate262inter2, gate262inter3, gate262inter4, gate262inter5, gate262inter6, gate262inter7, gate262inter8, gate262inter9, gate262inter10, gate262inter11, gate262inter12, gate208inter0, gate208inter1, gate208inter2, gate208inter3, gate208inter4, gate208inter5, gate208inter6, gate208inter7, gate208inter8, gate208inter9, gate208inter10, gate208inter11, gate208inter12, gate67inter0, gate67inter1, gate67inter2, gate67inter3, gate67inter4, gate67inter5, gate67inter6, gate67inter7, gate67inter8, gate67inter9, gate67inter10, gate67inter11, gate67inter12, gate242inter0, gate242inter1, gate242inter2, gate242inter3, gate242inter4, gate242inter5, gate242inter6, gate242inter7, gate242inter8, gate242inter9, gate242inter10, gate242inter11, gate242inter12, gate401inter0, gate401inter1, gate401inter2, gate401inter3, gate401inter4, gate401inter5, gate401inter6, gate401inter7, gate401inter8, gate401inter9, gate401inter10, gate401inter11, gate401inter12, gate463inter0, gate463inter1, gate463inter2, gate463inter3, gate463inter4, gate463inter5, gate463inter6, gate463inter7, gate463inter8, gate463inter9, gate463inter10, gate463inter11, gate463inter12, gate139inter0, gate139inter1, gate139inter2, gate139inter3, gate139inter4, gate139inter5, gate139inter6, gate139inter7, gate139inter8, gate139inter9, gate139inter10, gate139inter11, gate139inter12, gate23inter0, gate23inter1, gate23inter2, gate23inter3, gate23inter4, gate23inter5, gate23inter6, gate23inter7, gate23inter8, gate23inter9, gate23inter10, gate23inter11, gate23inter12, gate411inter0, gate411inter1, gate411inter2, gate411inter3, gate411inter4, gate411inter5, gate411inter6, gate411inter7, gate411inter8, gate411inter9, gate411inter10, gate411inter11, gate411inter12, gate17inter0, gate17inter1, gate17inter2, gate17inter3, gate17inter4, gate17inter5, gate17inter6, gate17inter7, gate17inter8, gate17inter9, gate17inter10, gate17inter11, gate17inter12, gate75inter0, gate75inter1, gate75inter2, gate75inter3, gate75inter4, gate75inter5, gate75inter6, gate75inter7, gate75inter8, gate75inter9, gate75inter10, gate75inter11, gate75inter12, gate34inter0, gate34inter1, gate34inter2, gate34inter3, gate34inter4, gate34inter5, gate34inter6, gate34inter7, gate34inter8, gate34inter9, gate34inter10, gate34inter11, gate34inter12, gate426inter0, gate426inter1, gate426inter2, gate426inter3, gate426inter4, gate426inter5, gate426inter6, gate426inter7, gate426inter8, gate426inter9, gate426inter10, gate426inter11, gate426inter12, gate220inter0, gate220inter1, gate220inter2, gate220inter3, gate220inter4, gate220inter5, gate220inter6, gate220inter7, gate220inter8, gate220inter9, gate220inter10, gate220inter11, gate220inter12, gate454inter0, gate454inter1, gate454inter2, gate454inter3, gate454inter4, gate454inter5, gate454inter6, gate454inter7, gate454inter8, gate454inter9, gate454inter10, gate454inter11, gate454inter12, gate184inter0, gate184inter1, gate184inter2, gate184inter3, gate184inter4, gate184inter5, gate184inter6, gate184inter7, gate184inter8, gate184inter9, gate184inter10, gate184inter11, gate184inter12, gate257inter0, gate257inter1, gate257inter2, gate257inter3, gate257inter4, gate257inter5, gate257inter6, gate257inter7, gate257inter8, gate257inter9, gate257inter10, gate257inter11, gate257inter12, gate108inter0, gate108inter1, gate108inter2, gate108inter3, gate108inter4, gate108inter5, gate108inter6, gate108inter7, gate108inter8, gate108inter9, gate108inter10, gate108inter11, gate108inter12, gate448inter0, gate448inter1, gate448inter2, gate448inter3, gate448inter4, gate448inter5, gate448inter6, gate448inter7, gate448inter8, gate448inter9, gate448inter10, gate448inter11, gate448inter12, gate397inter0, gate397inter1, gate397inter2, gate397inter3, gate397inter4, gate397inter5, gate397inter6, gate397inter7, gate397inter8, gate397inter9, gate397inter10, gate397inter11, gate397inter12, gate232inter0, gate232inter1, gate232inter2, gate232inter3, gate232inter4, gate232inter5, gate232inter6, gate232inter7, gate232inter8, gate232inter9, gate232inter10, gate232inter11, gate232inter12, gate39inter0, gate39inter1, gate39inter2, gate39inter3, gate39inter4, gate39inter5, gate39inter6, gate39inter7, gate39inter8, gate39inter9, gate39inter10, gate39inter11, gate39inter12, gate479inter0, gate479inter1, gate479inter2, gate479inter3, gate479inter4, gate479inter5, gate479inter6, gate479inter7, gate479inter8, gate479inter9, gate479inter10, gate479inter11, gate479inter12, gate276inter0, gate276inter1, gate276inter2, gate276inter3, gate276inter4, gate276inter5, gate276inter6, gate276inter7, gate276inter8, gate276inter9, gate276inter10, gate276inter11, gate276inter12, gate77inter0, gate77inter1, gate77inter2, gate77inter3, gate77inter4, gate77inter5, gate77inter6, gate77inter7, gate77inter8, gate77inter9, gate77inter10, gate77inter11, gate77inter12, gate485inter0, gate485inter1, gate485inter2, gate485inter3, gate485inter4, gate485inter5, gate485inter6, gate485inter7, gate485inter8, gate485inter9, gate485inter10, gate485inter11, gate485inter12, gate70inter0, gate70inter1, gate70inter2, gate70inter3, gate70inter4, gate70inter5, gate70inter6, gate70inter7, gate70inter8, gate70inter9, gate70inter10, gate70inter11, gate70inter12, gate241inter0, gate241inter1, gate241inter2, gate241inter3, gate241inter4, gate241inter5, gate241inter6, gate241inter7, gate241inter8, gate241inter9, gate241inter10, gate241inter11, gate241inter12, gate404inter0, gate404inter1, gate404inter2, gate404inter3, gate404inter4, gate404inter5, gate404inter6, gate404inter7, gate404inter8, gate404inter9, gate404inter10, gate404inter11, gate404inter12, gate483inter0, gate483inter1, gate483inter2, gate483inter3, gate483inter4, gate483inter5, gate483inter6, gate483inter7, gate483inter8, gate483inter9, gate483inter10, gate483inter11, gate483inter12, gate421inter0, gate421inter1, gate421inter2, gate421inter3, gate421inter4, gate421inter5, gate421inter6, gate421inter7, gate421inter8, gate421inter9, gate421inter10, gate421inter11, gate421inter12, gate295inter0, gate295inter1, gate295inter2, gate295inter3, gate295inter4, gate295inter5, gate295inter6, gate295inter7, gate295inter8, gate295inter9, gate295inter10, gate295inter11, gate295inter12, gate13inter0, gate13inter1, gate13inter2, gate13inter3, gate13inter4, gate13inter5, gate13inter6, gate13inter7, gate13inter8, gate13inter9, gate13inter10, gate13inter11, gate13inter12, gate21inter0, gate21inter1, gate21inter2, gate21inter3, gate21inter4, gate21inter5, gate21inter6, gate21inter7, gate21inter8, gate21inter9, gate21inter10, gate21inter11, gate21inter12, gate256inter0, gate256inter1, gate256inter2, gate256inter3, gate256inter4, gate256inter5, gate256inter6, gate256inter7, gate256inter8, gate256inter9, gate256inter10, gate256inter11, gate256inter12, gate253inter0, gate253inter1, gate253inter2, gate253inter3, gate253inter4, gate253inter5, gate253inter6, gate253inter7, gate253inter8, gate253inter9, gate253inter10, gate253inter11, gate253inter12, gate260inter0, gate260inter1, gate260inter2, gate260inter3, gate260inter4, gate260inter5, gate260inter6, gate260inter7, gate260inter8, gate260inter9, gate260inter10, gate260inter11, gate260inter12, gate159inter0, gate159inter1, gate159inter2, gate159inter3, gate159inter4, gate159inter5, gate159inter6, gate159inter7, gate159inter8, gate159inter9, gate159inter10, gate159inter11, gate159inter12, gate217inter0, gate217inter1, gate217inter2, gate217inter3, gate217inter4, gate217inter5, gate217inter6, gate217inter7, gate217inter8, gate217inter9, gate217inter10, gate217inter11, gate217inter12, gate64inter0, gate64inter1, gate64inter2, gate64inter3, gate64inter4, gate64inter5, gate64inter6, gate64inter7, gate64inter8, gate64inter9, gate64inter10, gate64inter11, gate64inter12, gate280inter0, gate280inter1, gate280inter2, gate280inter3, gate280inter4, gate280inter5, gate280inter6, gate280inter7, gate280inter8, gate280inter9, gate280inter10, gate280inter11, gate280inter12, gate270inter0, gate270inter1, gate270inter2, gate270inter3, gate270inter4, gate270inter5, gate270inter6, gate270inter7, gate270inter8, gate270inter9, gate270inter10, gate270inter11, gate270inter12, gate79inter0, gate79inter1, gate79inter2, gate79inter3, gate79inter4, gate79inter5, gate79inter6, gate79inter7, gate79inter8, gate79inter9, gate79inter10, gate79inter11, gate79inter12, gate19inter0, gate19inter1, gate19inter2, gate19inter3, gate19inter4, gate19inter5, gate19inter6, gate19inter7, gate19inter8, gate19inter9, gate19inter10, gate19inter11, gate19inter12, gate496inter0, gate496inter1, gate496inter2, gate496inter3, gate496inter4, gate496inter5, gate496inter6, gate496inter7, gate496inter8, gate496inter9, gate496inter10, gate496inter11, gate496inter12, gate44inter0, gate44inter1, gate44inter2, gate44inter3, gate44inter4, gate44inter5, gate44inter6, gate44inter7, gate44inter8, gate44inter9, gate44inter10, gate44inter11, gate44inter12, gate250inter0, gate250inter1, gate250inter2, gate250inter3, gate250inter4, gate250inter5, gate250inter6, gate250inter7, gate250inter8, gate250inter9, gate250inter10, gate250inter11, gate250inter12, gate249inter0, gate249inter1, gate249inter2, gate249inter3, gate249inter4, gate249inter5, gate249inter6, gate249inter7, gate249inter8, gate249inter9, gate249inter10, gate249inter11, gate249inter12;



and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );
nand2 gate9( .a(G1), .b(G2), .O(G266) );
nand2 gate10( .a(G3), .b(G4), .O(G269) );
nand2 gate11( .a(G5), .b(G6), .O(G272) );
nand2 gate12( .a(G7), .b(G8), .O(G275) );

  xor2  gate2507(.a(G10), .b(G9), .O(gate13inter0));
  nand2 gate2508(.a(gate13inter0), .b(s_280), .O(gate13inter1));
  and2  gate2509(.a(G10), .b(G9), .O(gate13inter2));
  inv1  gate2510(.a(s_280), .O(gate13inter3));
  inv1  gate2511(.a(s_281), .O(gate13inter4));
  nand2 gate2512(.a(gate13inter4), .b(gate13inter3), .O(gate13inter5));
  nor2  gate2513(.a(gate13inter5), .b(gate13inter2), .O(gate13inter6));
  inv1  gate2514(.a(G9), .O(gate13inter7));
  inv1  gate2515(.a(G10), .O(gate13inter8));
  nand2 gate2516(.a(gate13inter8), .b(gate13inter7), .O(gate13inter9));
  nand2 gate2517(.a(s_281), .b(gate13inter3), .O(gate13inter10));
  nor2  gate2518(.a(gate13inter10), .b(gate13inter9), .O(gate13inter11));
  nor2  gate2519(.a(gate13inter11), .b(gate13inter6), .O(gate13inter12));
  nand2 gate2520(.a(gate13inter12), .b(gate13inter1), .O(G278));
nand2 gate14( .a(G11), .b(G12), .O(G281) );
nand2 gate15( .a(G13), .b(G14), .O(G284) );
nand2 gate16( .a(G15), .b(G16), .O(G287) );

  xor2  gate2185(.a(G18), .b(G17), .O(gate17inter0));
  nand2 gate2186(.a(gate17inter0), .b(s_234), .O(gate17inter1));
  and2  gate2187(.a(G18), .b(G17), .O(gate17inter2));
  inv1  gate2188(.a(s_234), .O(gate17inter3));
  inv1  gate2189(.a(s_235), .O(gate17inter4));
  nand2 gate2190(.a(gate17inter4), .b(gate17inter3), .O(gate17inter5));
  nor2  gate2191(.a(gate17inter5), .b(gate17inter2), .O(gate17inter6));
  inv1  gate2192(.a(G17), .O(gate17inter7));
  inv1  gate2193(.a(G18), .O(gate17inter8));
  nand2 gate2194(.a(gate17inter8), .b(gate17inter7), .O(gate17inter9));
  nand2 gate2195(.a(s_235), .b(gate17inter3), .O(gate17inter10));
  nor2  gate2196(.a(gate17inter10), .b(gate17inter9), .O(gate17inter11));
  nor2  gate2197(.a(gate17inter11), .b(gate17inter6), .O(gate17inter12));
  nand2 gate2198(.a(gate17inter12), .b(gate17inter1), .O(G290));

  xor2  gate1163(.a(G20), .b(G19), .O(gate18inter0));
  nand2 gate1164(.a(gate18inter0), .b(s_88), .O(gate18inter1));
  and2  gate1165(.a(G20), .b(G19), .O(gate18inter2));
  inv1  gate1166(.a(s_88), .O(gate18inter3));
  inv1  gate1167(.a(s_89), .O(gate18inter4));
  nand2 gate1168(.a(gate18inter4), .b(gate18inter3), .O(gate18inter5));
  nor2  gate1169(.a(gate18inter5), .b(gate18inter2), .O(gate18inter6));
  inv1  gate1170(.a(G19), .O(gate18inter7));
  inv1  gate1171(.a(G20), .O(gate18inter8));
  nand2 gate1172(.a(gate18inter8), .b(gate18inter7), .O(gate18inter9));
  nand2 gate1173(.a(s_89), .b(gate18inter3), .O(gate18inter10));
  nor2  gate1174(.a(gate18inter10), .b(gate18inter9), .O(gate18inter11));
  nor2  gate1175(.a(gate18inter11), .b(gate18inter6), .O(gate18inter12));
  nand2 gate1176(.a(gate18inter12), .b(gate18inter1), .O(G293));

  xor2  gate2661(.a(G22), .b(G21), .O(gate19inter0));
  nand2 gate2662(.a(gate19inter0), .b(s_302), .O(gate19inter1));
  and2  gate2663(.a(G22), .b(G21), .O(gate19inter2));
  inv1  gate2664(.a(s_302), .O(gate19inter3));
  inv1  gate2665(.a(s_303), .O(gate19inter4));
  nand2 gate2666(.a(gate19inter4), .b(gate19inter3), .O(gate19inter5));
  nor2  gate2667(.a(gate19inter5), .b(gate19inter2), .O(gate19inter6));
  inv1  gate2668(.a(G21), .O(gate19inter7));
  inv1  gate2669(.a(G22), .O(gate19inter8));
  nand2 gate2670(.a(gate19inter8), .b(gate19inter7), .O(gate19inter9));
  nand2 gate2671(.a(s_303), .b(gate19inter3), .O(gate19inter10));
  nor2  gate2672(.a(gate19inter10), .b(gate19inter9), .O(gate19inter11));
  nor2  gate2673(.a(gate19inter11), .b(gate19inter6), .O(gate19inter12));
  nand2 gate2674(.a(gate19inter12), .b(gate19inter1), .O(G296));

  xor2  gate2017(.a(G24), .b(G23), .O(gate20inter0));
  nand2 gate2018(.a(gate20inter0), .b(s_210), .O(gate20inter1));
  and2  gate2019(.a(G24), .b(G23), .O(gate20inter2));
  inv1  gate2020(.a(s_210), .O(gate20inter3));
  inv1  gate2021(.a(s_211), .O(gate20inter4));
  nand2 gate2022(.a(gate20inter4), .b(gate20inter3), .O(gate20inter5));
  nor2  gate2023(.a(gate20inter5), .b(gate20inter2), .O(gate20inter6));
  inv1  gate2024(.a(G23), .O(gate20inter7));
  inv1  gate2025(.a(G24), .O(gate20inter8));
  nand2 gate2026(.a(gate20inter8), .b(gate20inter7), .O(gate20inter9));
  nand2 gate2027(.a(s_211), .b(gate20inter3), .O(gate20inter10));
  nor2  gate2028(.a(gate20inter10), .b(gate20inter9), .O(gate20inter11));
  nor2  gate2029(.a(gate20inter11), .b(gate20inter6), .O(gate20inter12));
  nand2 gate2030(.a(gate20inter12), .b(gate20inter1), .O(G299));

  xor2  gate2521(.a(G26), .b(G25), .O(gate21inter0));
  nand2 gate2522(.a(gate21inter0), .b(s_282), .O(gate21inter1));
  and2  gate2523(.a(G26), .b(G25), .O(gate21inter2));
  inv1  gate2524(.a(s_282), .O(gate21inter3));
  inv1  gate2525(.a(s_283), .O(gate21inter4));
  nand2 gate2526(.a(gate21inter4), .b(gate21inter3), .O(gate21inter5));
  nor2  gate2527(.a(gate21inter5), .b(gate21inter2), .O(gate21inter6));
  inv1  gate2528(.a(G25), .O(gate21inter7));
  inv1  gate2529(.a(G26), .O(gate21inter8));
  nand2 gate2530(.a(gate21inter8), .b(gate21inter7), .O(gate21inter9));
  nand2 gate2531(.a(s_283), .b(gate21inter3), .O(gate21inter10));
  nor2  gate2532(.a(gate21inter10), .b(gate21inter9), .O(gate21inter11));
  nor2  gate2533(.a(gate21inter11), .b(gate21inter6), .O(gate21inter12));
  nand2 gate2534(.a(gate21inter12), .b(gate21inter1), .O(G302));
nand2 gate22( .a(G27), .b(G28), .O(G305) );

  xor2  gate2157(.a(G30), .b(G29), .O(gate23inter0));
  nand2 gate2158(.a(gate23inter0), .b(s_230), .O(gate23inter1));
  and2  gate2159(.a(G30), .b(G29), .O(gate23inter2));
  inv1  gate2160(.a(s_230), .O(gate23inter3));
  inv1  gate2161(.a(s_231), .O(gate23inter4));
  nand2 gate2162(.a(gate23inter4), .b(gate23inter3), .O(gate23inter5));
  nor2  gate2163(.a(gate23inter5), .b(gate23inter2), .O(gate23inter6));
  inv1  gate2164(.a(G29), .O(gate23inter7));
  inv1  gate2165(.a(G30), .O(gate23inter8));
  nand2 gate2166(.a(gate23inter8), .b(gate23inter7), .O(gate23inter9));
  nand2 gate2167(.a(s_231), .b(gate23inter3), .O(gate23inter10));
  nor2  gate2168(.a(gate23inter10), .b(gate23inter9), .O(gate23inter11));
  nor2  gate2169(.a(gate23inter11), .b(gate23inter6), .O(gate23inter12));
  nand2 gate2170(.a(gate23inter12), .b(gate23inter1), .O(G308));
nand2 gate24( .a(G31), .b(G32), .O(G311) );
nand2 gate25( .a(G1), .b(G5), .O(G314) );

  xor2  gate1443(.a(G13), .b(G9), .O(gate26inter0));
  nand2 gate1444(.a(gate26inter0), .b(s_128), .O(gate26inter1));
  and2  gate1445(.a(G13), .b(G9), .O(gate26inter2));
  inv1  gate1446(.a(s_128), .O(gate26inter3));
  inv1  gate1447(.a(s_129), .O(gate26inter4));
  nand2 gate1448(.a(gate26inter4), .b(gate26inter3), .O(gate26inter5));
  nor2  gate1449(.a(gate26inter5), .b(gate26inter2), .O(gate26inter6));
  inv1  gate1450(.a(G9), .O(gate26inter7));
  inv1  gate1451(.a(G13), .O(gate26inter8));
  nand2 gate1452(.a(gate26inter8), .b(gate26inter7), .O(gate26inter9));
  nand2 gate1453(.a(s_129), .b(gate26inter3), .O(gate26inter10));
  nor2  gate1454(.a(gate26inter10), .b(gate26inter9), .O(gate26inter11));
  nor2  gate1455(.a(gate26inter11), .b(gate26inter6), .O(gate26inter12));
  nand2 gate1456(.a(gate26inter12), .b(gate26inter1), .O(G317));

  xor2  gate1135(.a(G6), .b(G2), .O(gate27inter0));
  nand2 gate1136(.a(gate27inter0), .b(s_84), .O(gate27inter1));
  and2  gate1137(.a(G6), .b(G2), .O(gate27inter2));
  inv1  gate1138(.a(s_84), .O(gate27inter3));
  inv1  gate1139(.a(s_85), .O(gate27inter4));
  nand2 gate1140(.a(gate27inter4), .b(gate27inter3), .O(gate27inter5));
  nor2  gate1141(.a(gate27inter5), .b(gate27inter2), .O(gate27inter6));
  inv1  gate1142(.a(G2), .O(gate27inter7));
  inv1  gate1143(.a(G6), .O(gate27inter8));
  nand2 gate1144(.a(gate27inter8), .b(gate27inter7), .O(gate27inter9));
  nand2 gate1145(.a(s_85), .b(gate27inter3), .O(gate27inter10));
  nor2  gate1146(.a(gate27inter10), .b(gate27inter9), .O(gate27inter11));
  nor2  gate1147(.a(gate27inter11), .b(gate27inter6), .O(gate27inter12));
  nand2 gate1148(.a(gate27inter12), .b(gate27inter1), .O(G320));
nand2 gate28( .a(G10), .b(G14), .O(G323) );
nand2 gate29( .a(G3), .b(G7), .O(G326) );
nand2 gate30( .a(G11), .b(G15), .O(G329) );
nand2 gate31( .a(G4), .b(G8), .O(G332) );
nand2 gate32( .a(G12), .b(G16), .O(G335) );
nand2 gate33( .a(G17), .b(G21), .O(G338) );

  xor2  gate2213(.a(G29), .b(G25), .O(gate34inter0));
  nand2 gate2214(.a(gate34inter0), .b(s_238), .O(gate34inter1));
  and2  gate2215(.a(G29), .b(G25), .O(gate34inter2));
  inv1  gate2216(.a(s_238), .O(gate34inter3));
  inv1  gate2217(.a(s_239), .O(gate34inter4));
  nand2 gate2218(.a(gate34inter4), .b(gate34inter3), .O(gate34inter5));
  nor2  gate2219(.a(gate34inter5), .b(gate34inter2), .O(gate34inter6));
  inv1  gate2220(.a(G25), .O(gate34inter7));
  inv1  gate2221(.a(G29), .O(gate34inter8));
  nand2 gate2222(.a(gate34inter8), .b(gate34inter7), .O(gate34inter9));
  nand2 gate2223(.a(s_239), .b(gate34inter3), .O(gate34inter10));
  nor2  gate2224(.a(gate34inter10), .b(gate34inter9), .O(gate34inter11));
  nor2  gate2225(.a(gate34inter11), .b(gate34inter6), .O(gate34inter12));
  nand2 gate2226(.a(gate34inter12), .b(gate34inter1), .O(G341));

  xor2  gate1107(.a(G22), .b(G18), .O(gate35inter0));
  nand2 gate1108(.a(gate35inter0), .b(s_80), .O(gate35inter1));
  and2  gate1109(.a(G22), .b(G18), .O(gate35inter2));
  inv1  gate1110(.a(s_80), .O(gate35inter3));
  inv1  gate1111(.a(s_81), .O(gate35inter4));
  nand2 gate1112(.a(gate35inter4), .b(gate35inter3), .O(gate35inter5));
  nor2  gate1113(.a(gate35inter5), .b(gate35inter2), .O(gate35inter6));
  inv1  gate1114(.a(G18), .O(gate35inter7));
  inv1  gate1115(.a(G22), .O(gate35inter8));
  nand2 gate1116(.a(gate35inter8), .b(gate35inter7), .O(gate35inter9));
  nand2 gate1117(.a(s_81), .b(gate35inter3), .O(gate35inter10));
  nor2  gate1118(.a(gate35inter10), .b(gate35inter9), .O(gate35inter11));
  nor2  gate1119(.a(gate35inter11), .b(gate35inter6), .O(gate35inter12));
  nand2 gate1120(.a(gate35inter12), .b(gate35inter1), .O(G344));
nand2 gate36( .a(G26), .b(G30), .O(G347) );
nand2 gate37( .a(G19), .b(G23), .O(G350) );
nand2 gate38( .a(G27), .b(G31), .O(G353) );

  xor2  gate2353(.a(G24), .b(G20), .O(gate39inter0));
  nand2 gate2354(.a(gate39inter0), .b(s_258), .O(gate39inter1));
  and2  gate2355(.a(G24), .b(G20), .O(gate39inter2));
  inv1  gate2356(.a(s_258), .O(gate39inter3));
  inv1  gate2357(.a(s_259), .O(gate39inter4));
  nand2 gate2358(.a(gate39inter4), .b(gate39inter3), .O(gate39inter5));
  nor2  gate2359(.a(gate39inter5), .b(gate39inter2), .O(gate39inter6));
  inv1  gate2360(.a(G20), .O(gate39inter7));
  inv1  gate2361(.a(G24), .O(gate39inter8));
  nand2 gate2362(.a(gate39inter8), .b(gate39inter7), .O(gate39inter9));
  nand2 gate2363(.a(s_259), .b(gate39inter3), .O(gate39inter10));
  nor2  gate2364(.a(gate39inter10), .b(gate39inter9), .O(gate39inter11));
  nor2  gate2365(.a(gate39inter11), .b(gate39inter6), .O(gate39inter12));
  nand2 gate2366(.a(gate39inter12), .b(gate39inter1), .O(G356));
nand2 gate40( .a(G28), .b(G32), .O(G359) );
nand2 gate41( .a(G1), .b(G266), .O(G362) );
nand2 gate42( .a(G2), .b(G266), .O(G363) );
nand2 gate43( .a(G3), .b(G269), .O(G364) );

  xor2  gate2689(.a(G269), .b(G4), .O(gate44inter0));
  nand2 gate2690(.a(gate44inter0), .b(s_306), .O(gate44inter1));
  and2  gate2691(.a(G269), .b(G4), .O(gate44inter2));
  inv1  gate2692(.a(s_306), .O(gate44inter3));
  inv1  gate2693(.a(s_307), .O(gate44inter4));
  nand2 gate2694(.a(gate44inter4), .b(gate44inter3), .O(gate44inter5));
  nor2  gate2695(.a(gate44inter5), .b(gate44inter2), .O(gate44inter6));
  inv1  gate2696(.a(G4), .O(gate44inter7));
  inv1  gate2697(.a(G269), .O(gate44inter8));
  nand2 gate2698(.a(gate44inter8), .b(gate44inter7), .O(gate44inter9));
  nand2 gate2699(.a(s_307), .b(gate44inter3), .O(gate44inter10));
  nor2  gate2700(.a(gate44inter10), .b(gate44inter9), .O(gate44inter11));
  nor2  gate2701(.a(gate44inter11), .b(gate44inter6), .O(gate44inter12));
  nand2 gate2702(.a(gate44inter12), .b(gate44inter1), .O(G365));

  xor2  gate547(.a(G272), .b(G5), .O(gate45inter0));
  nand2 gate548(.a(gate45inter0), .b(s_0), .O(gate45inter1));
  and2  gate549(.a(G272), .b(G5), .O(gate45inter2));
  inv1  gate550(.a(s_0), .O(gate45inter3));
  inv1  gate551(.a(s_1), .O(gate45inter4));
  nand2 gate552(.a(gate45inter4), .b(gate45inter3), .O(gate45inter5));
  nor2  gate553(.a(gate45inter5), .b(gate45inter2), .O(gate45inter6));
  inv1  gate554(.a(G5), .O(gate45inter7));
  inv1  gate555(.a(G272), .O(gate45inter8));
  nand2 gate556(.a(gate45inter8), .b(gate45inter7), .O(gate45inter9));
  nand2 gate557(.a(s_1), .b(gate45inter3), .O(gate45inter10));
  nor2  gate558(.a(gate45inter10), .b(gate45inter9), .O(gate45inter11));
  nor2  gate559(.a(gate45inter11), .b(gate45inter6), .O(gate45inter12));
  nand2 gate560(.a(gate45inter12), .b(gate45inter1), .O(G366));
nand2 gate46( .a(G6), .b(G272), .O(G367) );
nand2 gate47( .a(G7), .b(G275), .O(G368) );

  xor2  gate701(.a(G275), .b(G8), .O(gate48inter0));
  nand2 gate702(.a(gate48inter0), .b(s_22), .O(gate48inter1));
  and2  gate703(.a(G275), .b(G8), .O(gate48inter2));
  inv1  gate704(.a(s_22), .O(gate48inter3));
  inv1  gate705(.a(s_23), .O(gate48inter4));
  nand2 gate706(.a(gate48inter4), .b(gate48inter3), .O(gate48inter5));
  nor2  gate707(.a(gate48inter5), .b(gate48inter2), .O(gate48inter6));
  inv1  gate708(.a(G8), .O(gate48inter7));
  inv1  gate709(.a(G275), .O(gate48inter8));
  nand2 gate710(.a(gate48inter8), .b(gate48inter7), .O(gate48inter9));
  nand2 gate711(.a(s_23), .b(gate48inter3), .O(gate48inter10));
  nor2  gate712(.a(gate48inter10), .b(gate48inter9), .O(gate48inter11));
  nor2  gate713(.a(gate48inter11), .b(gate48inter6), .O(gate48inter12));
  nand2 gate714(.a(gate48inter12), .b(gate48inter1), .O(G369));
nand2 gate49( .a(G9), .b(G278), .O(G370) );
nand2 gate50( .a(G10), .b(G278), .O(G371) );

  xor2  gate589(.a(G281), .b(G11), .O(gate51inter0));
  nand2 gate590(.a(gate51inter0), .b(s_6), .O(gate51inter1));
  and2  gate591(.a(G281), .b(G11), .O(gate51inter2));
  inv1  gate592(.a(s_6), .O(gate51inter3));
  inv1  gate593(.a(s_7), .O(gate51inter4));
  nand2 gate594(.a(gate51inter4), .b(gate51inter3), .O(gate51inter5));
  nor2  gate595(.a(gate51inter5), .b(gate51inter2), .O(gate51inter6));
  inv1  gate596(.a(G11), .O(gate51inter7));
  inv1  gate597(.a(G281), .O(gate51inter8));
  nand2 gate598(.a(gate51inter8), .b(gate51inter7), .O(gate51inter9));
  nand2 gate599(.a(s_7), .b(gate51inter3), .O(gate51inter10));
  nor2  gate600(.a(gate51inter10), .b(gate51inter9), .O(gate51inter11));
  nor2  gate601(.a(gate51inter11), .b(gate51inter6), .O(gate51inter12));
  nand2 gate602(.a(gate51inter12), .b(gate51inter1), .O(G372));
nand2 gate52( .a(G12), .b(G281), .O(G373) );

  xor2  gate869(.a(G284), .b(G13), .O(gate53inter0));
  nand2 gate870(.a(gate53inter0), .b(s_46), .O(gate53inter1));
  and2  gate871(.a(G284), .b(G13), .O(gate53inter2));
  inv1  gate872(.a(s_46), .O(gate53inter3));
  inv1  gate873(.a(s_47), .O(gate53inter4));
  nand2 gate874(.a(gate53inter4), .b(gate53inter3), .O(gate53inter5));
  nor2  gate875(.a(gate53inter5), .b(gate53inter2), .O(gate53inter6));
  inv1  gate876(.a(G13), .O(gate53inter7));
  inv1  gate877(.a(G284), .O(gate53inter8));
  nand2 gate878(.a(gate53inter8), .b(gate53inter7), .O(gate53inter9));
  nand2 gate879(.a(s_47), .b(gate53inter3), .O(gate53inter10));
  nor2  gate880(.a(gate53inter10), .b(gate53inter9), .O(gate53inter11));
  nor2  gate881(.a(gate53inter11), .b(gate53inter6), .O(gate53inter12));
  nand2 gate882(.a(gate53inter12), .b(gate53inter1), .O(G374));

  xor2  gate1359(.a(G284), .b(G14), .O(gate54inter0));
  nand2 gate1360(.a(gate54inter0), .b(s_116), .O(gate54inter1));
  and2  gate1361(.a(G284), .b(G14), .O(gate54inter2));
  inv1  gate1362(.a(s_116), .O(gate54inter3));
  inv1  gate1363(.a(s_117), .O(gate54inter4));
  nand2 gate1364(.a(gate54inter4), .b(gate54inter3), .O(gate54inter5));
  nor2  gate1365(.a(gate54inter5), .b(gate54inter2), .O(gate54inter6));
  inv1  gate1366(.a(G14), .O(gate54inter7));
  inv1  gate1367(.a(G284), .O(gate54inter8));
  nand2 gate1368(.a(gate54inter8), .b(gate54inter7), .O(gate54inter9));
  nand2 gate1369(.a(s_117), .b(gate54inter3), .O(gate54inter10));
  nor2  gate1370(.a(gate54inter10), .b(gate54inter9), .O(gate54inter11));
  nor2  gate1371(.a(gate54inter11), .b(gate54inter6), .O(gate54inter12));
  nand2 gate1372(.a(gate54inter12), .b(gate54inter1), .O(G375));
nand2 gate55( .a(G15), .b(G287), .O(G376) );

  xor2  gate799(.a(G287), .b(G16), .O(gate56inter0));
  nand2 gate800(.a(gate56inter0), .b(s_36), .O(gate56inter1));
  and2  gate801(.a(G287), .b(G16), .O(gate56inter2));
  inv1  gate802(.a(s_36), .O(gate56inter3));
  inv1  gate803(.a(s_37), .O(gate56inter4));
  nand2 gate804(.a(gate56inter4), .b(gate56inter3), .O(gate56inter5));
  nor2  gate805(.a(gate56inter5), .b(gate56inter2), .O(gate56inter6));
  inv1  gate806(.a(G16), .O(gate56inter7));
  inv1  gate807(.a(G287), .O(gate56inter8));
  nand2 gate808(.a(gate56inter8), .b(gate56inter7), .O(gate56inter9));
  nand2 gate809(.a(s_37), .b(gate56inter3), .O(gate56inter10));
  nor2  gate810(.a(gate56inter10), .b(gate56inter9), .O(gate56inter11));
  nor2  gate811(.a(gate56inter11), .b(gate56inter6), .O(gate56inter12));
  nand2 gate812(.a(gate56inter12), .b(gate56inter1), .O(G377));
nand2 gate57( .a(G17), .b(G290), .O(G378) );

  xor2  gate631(.a(G290), .b(G18), .O(gate58inter0));
  nand2 gate632(.a(gate58inter0), .b(s_12), .O(gate58inter1));
  and2  gate633(.a(G290), .b(G18), .O(gate58inter2));
  inv1  gate634(.a(s_12), .O(gate58inter3));
  inv1  gate635(.a(s_13), .O(gate58inter4));
  nand2 gate636(.a(gate58inter4), .b(gate58inter3), .O(gate58inter5));
  nor2  gate637(.a(gate58inter5), .b(gate58inter2), .O(gate58inter6));
  inv1  gate638(.a(G18), .O(gate58inter7));
  inv1  gate639(.a(G290), .O(gate58inter8));
  nand2 gate640(.a(gate58inter8), .b(gate58inter7), .O(gate58inter9));
  nand2 gate641(.a(s_13), .b(gate58inter3), .O(gate58inter10));
  nor2  gate642(.a(gate58inter10), .b(gate58inter9), .O(gate58inter11));
  nor2  gate643(.a(gate58inter11), .b(gate58inter6), .O(gate58inter12));
  nand2 gate644(.a(gate58inter12), .b(gate58inter1), .O(G379));

  xor2  gate1233(.a(G293), .b(G19), .O(gate59inter0));
  nand2 gate1234(.a(gate59inter0), .b(s_98), .O(gate59inter1));
  and2  gate1235(.a(G293), .b(G19), .O(gate59inter2));
  inv1  gate1236(.a(s_98), .O(gate59inter3));
  inv1  gate1237(.a(s_99), .O(gate59inter4));
  nand2 gate1238(.a(gate59inter4), .b(gate59inter3), .O(gate59inter5));
  nor2  gate1239(.a(gate59inter5), .b(gate59inter2), .O(gate59inter6));
  inv1  gate1240(.a(G19), .O(gate59inter7));
  inv1  gate1241(.a(G293), .O(gate59inter8));
  nand2 gate1242(.a(gate59inter8), .b(gate59inter7), .O(gate59inter9));
  nand2 gate1243(.a(s_99), .b(gate59inter3), .O(gate59inter10));
  nor2  gate1244(.a(gate59inter10), .b(gate59inter9), .O(gate59inter11));
  nor2  gate1245(.a(gate59inter11), .b(gate59inter6), .O(gate59inter12));
  nand2 gate1246(.a(gate59inter12), .b(gate59inter1), .O(G380));
nand2 gate60( .a(G20), .b(G293), .O(G381) );
nand2 gate61( .a(G21), .b(G296), .O(G382) );
nand2 gate62( .a(G22), .b(G296), .O(G383) );

  xor2  gate1751(.a(G299), .b(G23), .O(gate63inter0));
  nand2 gate1752(.a(gate63inter0), .b(s_172), .O(gate63inter1));
  and2  gate1753(.a(G299), .b(G23), .O(gate63inter2));
  inv1  gate1754(.a(s_172), .O(gate63inter3));
  inv1  gate1755(.a(s_173), .O(gate63inter4));
  nand2 gate1756(.a(gate63inter4), .b(gate63inter3), .O(gate63inter5));
  nor2  gate1757(.a(gate63inter5), .b(gate63inter2), .O(gate63inter6));
  inv1  gate1758(.a(G23), .O(gate63inter7));
  inv1  gate1759(.a(G299), .O(gate63inter8));
  nand2 gate1760(.a(gate63inter8), .b(gate63inter7), .O(gate63inter9));
  nand2 gate1761(.a(s_173), .b(gate63inter3), .O(gate63inter10));
  nor2  gate1762(.a(gate63inter10), .b(gate63inter9), .O(gate63inter11));
  nor2  gate1763(.a(gate63inter11), .b(gate63inter6), .O(gate63inter12));
  nand2 gate1764(.a(gate63inter12), .b(gate63inter1), .O(G384));

  xor2  gate2605(.a(G299), .b(G24), .O(gate64inter0));
  nand2 gate2606(.a(gate64inter0), .b(s_294), .O(gate64inter1));
  and2  gate2607(.a(G299), .b(G24), .O(gate64inter2));
  inv1  gate2608(.a(s_294), .O(gate64inter3));
  inv1  gate2609(.a(s_295), .O(gate64inter4));
  nand2 gate2610(.a(gate64inter4), .b(gate64inter3), .O(gate64inter5));
  nor2  gate2611(.a(gate64inter5), .b(gate64inter2), .O(gate64inter6));
  inv1  gate2612(.a(G24), .O(gate64inter7));
  inv1  gate2613(.a(G299), .O(gate64inter8));
  nand2 gate2614(.a(gate64inter8), .b(gate64inter7), .O(gate64inter9));
  nand2 gate2615(.a(s_295), .b(gate64inter3), .O(gate64inter10));
  nor2  gate2616(.a(gate64inter10), .b(gate64inter9), .O(gate64inter11));
  nor2  gate2617(.a(gate64inter11), .b(gate64inter6), .O(gate64inter12));
  nand2 gate2618(.a(gate64inter12), .b(gate64inter1), .O(G385));
nand2 gate65( .a(G25), .b(G302), .O(G386) );
nand2 gate66( .a(G26), .b(G302), .O(G387) );

  xor2  gate2087(.a(G305), .b(G27), .O(gate67inter0));
  nand2 gate2088(.a(gate67inter0), .b(s_220), .O(gate67inter1));
  and2  gate2089(.a(G305), .b(G27), .O(gate67inter2));
  inv1  gate2090(.a(s_220), .O(gate67inter3));
  inv1  gate2091(.a(s_221), .O(gate67inter4));
  nand2 gate2092(.a(gate67inter4), .b(gate67inter3), .O(gate67inter5));
  nor2  gate2093(.a(gate67inter5), .b(gate67inter2), .O(gate67inter6));
  inv1  gate2094(.a(G27), .O(gate67inter7));
  inv1  gate2095(.a(G305), .O(gate67inter8));
  nand2 gate2096(.a(gate67inter8), .b(gate67inter7), .O(gate67inter9));
  nand2 gate2097(.a(s_221), .b(gate67inter3), .O(gate67inter10));
  nor2  gate2098(.a(gate67inter10), .b(gate67inter9), .O(gate67inter11));
  nor2  gate2099(.a(gate67inter11), .b(gate67inter6), .O(gate67inter12));
  nand2 gate2100(.a(gate67inter12), .b(gate67inter1), .O(G388));
nand2 gate68( .a(G28), .b(G305), .O(G389) );

  xor2  gate1779(.a(G308), .b(G29), .O(gate69inter0));
  nand2 gate1780(.a(gate69inter0), .b(s_176), .O(gate69inter1));
  and2  gate1781(.a(G308), .b(G29), .O(gate69inter2));
  inv1  gate1782(.a(s_176), .O(gate69inter3));
  inv1  gate1783(.a(s_177), .O(gate69inter4));
  nand2 gate1784(.a(gate69inter4), .b(gate69inter3), .O(gate69inter5));
  nor2  gate1785(.a(gate69inter5), .b(gate69inter2), .O(gate69inter6));
  inv1  gate1786(.a(G29), .O(gate69inter7));
  inv1  gate1787(.a(G308), .O(gate69inter8));
  nand2 gate1788(.a(gate69inter8), .b(gate69inter7), .O(gate69inter9));
  nand2 gate1789(.a(s_177), .b(gate69inter3), .O(gate69inter10));
  nor2  gate1790(.a(gate69inter10), .b(gate69inter9), .O(gate69inter11));
  nor2  gate1791(.a(gate69inter11), .b(gate69inter6), .O(gate69inter12));
  nand2 gate1792(.a(gate69inter12), .b(gate69inter1), .O(G390));

  xor2  gate2423(.a(G308), .b(G30), .O(gate70inter0));
  nand2 gate2424(.a(gate70inter0), .b(s_268), .O(gate70inter1));
  and2  gate2425(.a(G308), .b(G30), .O(gate70inter2));
  inv1  gate2426(.a(s_268), .O(gate70inter3));
  inv1  gate2427(.a(s_269), .O(gate70inter4));
  nand2 gate2428(.a(gate70inter4), .b(gate70inter3), .O(gate70inter5));
  nor2  gate2429(.a(gate70inter5), .b(gate70inter2), .O(gate70inter6));
  inv1  gate2430(.a(G30), .O(gate70inter7));
  inv1  gate2431(.a(G308), .O(gate70inter8));
  nand2 gate2432(.a(gate70inter8), .b(gate70inter7), .O(gate70inter9));
  nand2 gate2433(.a(s_269), .b(gate70inter3), .O(gate70inter10));
  nor2  gate2434(.a(gate70inter10), .b(gate70inter9), .O(gate70inter11));
  nor2  gate2435(.a(gate70inter11), .b(gate70inter6), .O(gate70inter12));
  nand2 gate2436(.a(gate70inter12), .b(gate70inter1), .O(G391));
nand2 gate71( .a(G31), .b(G311), .O(G392) );

  xor2  gate1219(.a(G311), .b(G32), .O(gate72inter0));
  nand2 gate1220(.a(gate72inter0), .b(s_96), .O(gate72inter1));
  and2  gate1221(.a(G311), .b(G32), .O(gate72inter2));
  inv1  gate1222(.a(s_96), .O(gate72inter3));
  inv1  gate1223(.a(s_97), .O(gate72inter4));
  nand2 gate1224(.a(gate72inter4), .b(gate72inter3), .O(gate72inter5));
  nor2  gate1225(.a(gate72inter5), .b(gate72inter2), .O(gate72inter6));
  inv1  gate1226(.a(G32), .O(gate72inter7));
  inv1  gate1227(.a(G311), .O(gate72inter8));
  nand2 gate1228(.a(gate72inter8), .b(gate72inter7), .O(gate72inter9));
  nand2 gate1229(.a(s_97), .b(gate72inter3), .O(gate72inter10));
  nor2  gate1230(.a(gate72inter10), .b(gate72inter9), .O(gate72inter11));
  nor2  gate1231(.a(gate72inter11), .b(gate72inter6), .O(gate72inter12));
  nand2 gate1232(.a(gate72inter12), .b(gate72inter1), .O(G393));

  xor2  gate617(.a(G314), .b(G1), .O(gate73inter0));
  nand2 gate618(.a(gate73inter0), .b(s_10), .O(gate73inter1));
  and2  gate619(.a(G314), .b(G1), .O(gate73inter2));
  inv1  gate620(.a(s_10), .O(gate73inter3));
  inv1  gate621(.a(s_11), .O(gate73inter4));
  nand2 gate622(.a(gate73inter4), .b(gate73inter3), .O(gate73inter5));
  nor2  gate623(.a(gate73inter5), .b(gate73inter2), .O(gate73inter6));
  inv1  gate624(.a(G1), .O(gate73inter7));
  inv1  gate625(.a(G314), .O(gate73inter8));
  nand2 gate626(.a(gate73inter8), .b(gate73inter7), .O(gate73inter9));
  nand2 gate627(.a(s_11), .b(gate73inter3), .O(gate73inter10));
  nor2  gate628(.a(gate73inter10), .b(gate73inter9), .O(gate73inter11));
  nor2  gate629(.a(gate73inter11), .b(gate73inter6), .O(gate73inter12));
  nand2 gate630(.a(gate73inter12), .b(gate73inter1), .O(G394));

  xor2  gate2031(.a(G314), .b(G5), .O(gate74inter0));
  nand2 gate2032(.a(gate74inter0), .b(s_212), .O(gate74inter1));
  and2  gate2033(.a(G314), .b(G5), .O(gate74inter2));
  inv1  gate2034(.a(s_212), .O(gate74inter3));
  inv1  gate2035(.a(s_213), .O(gate74inter4));
  nand2 gate2036(.a(gate74inter4), .b(gate74inter3), .O(gate74inter5));
  nor2  gate2037(.a(gate74inter5), .b(gate74inter2), .O(gate74inter6));
  inv1  gate2038(.a(G5), .O(gate74inter7));
  inv1  gate2039(.a(G314), .O(gate74inter8));
  nand2 gate2040(.a(gate74inter8), .b(gate74inter7), .O(gate74inter9));
  nand2 gate2041(.a(s_213), .b(gate74inter3), .O(gate74inter10));
  nor2  gate2042(.a(gate74inter10), .b(gate74inter9), .O(gate74inter11));
  nor2  gate2043(.a(gate74inter11), .b(gate74inter6), .O(gate74inter12));
  nand2 gate2044(.a(gate74inter12), .b(gate74inter1), .O(G395));

  xor2  gate2199(.a(G317), .b(G9), .O(gate75inter0));
  nand2 gate2200(.a(gate75inter0), .b(s_236), .O(gate75inter1));
  and2  gate2201(.a(G317), .b(G9), .O(gate75inter2));
  inv1  gate2202(.a(s_236), .O(gate75inter3));
  inv1  gate2203(.a(s_237), .O(gate75inter4));
  nand2 gate2204(.a(gate75inter4), .b(gate75inter3), .O(gate75inter5));
  nor2  gate2205(.a(gate75inter5), .b(gate75inter2), .O(gate75inter6));
  inv1  gate2206(.a(G9), .O(gate75inter7));
  inv1  gate2207(.a(G317), .O(gate75inter8));
  nand2 gate2208(.a(gate75inter8), .b(gate75inter7), .O(gate75inter9));
  nand2 gate2209(.a(s_237), .b(gate75inter3), .O(gate75inter10));
  nor2  gate2210(.a(gate75inter10), .b(gate75inter9), .O(gate75inter11));
  nor2  gate2211(.a(gate75inter11), .b(gate75inter6), .O(gate75inter12));
  nand2 gate2212(.a(gate75inter12), .b(gate75inter1), .O(G396));
nand2 gate76( .a(G13), .b(G317), .O(G397) );

  xor2  gate2395(.a(G320), .b(G2), .O(gate77inter0));
  nand2 gate2396(.a(gate77inter0), .b(s_264), .O(gate77inter1));
  and2  gate2397(.a(G320), .b(G2), .O(gate77inter2));
  inv1  gate2398(.a(s_264), .O(gate77inter3));
  inv1  gate2399(.a(s_265), .O(gate77inter4));
  nand2 gate2400(.a(gate77inter4), .b(gate77inter3), .O(gate77inter5));
  nor2  gate2401(.a(gate77inter5), .b(gate77inter2), .O(gate77inter6));
  inv1  gate2402(.a(G2), .O(gate77inter7));
  inv1  gate2403(.a(G320), .O(gate77inter8));
  nand2 gate2404(.a(gate77inter8), .b(gate77inter7), .O(gate77inter9));
  nand2 gate2405(.a(s_265), .b(gate77inter3), .O(gate77inter10));
  nor2  gate2406(.a(gate77inter10), .b(gate77inter9), .O(gate77inter11));
  nor2  gate2407(.a(gate77inter11), .b(gate77inter6), .O(gate77inter12));
  nand2 gate2408(.a(gate77inter12), .b(gate77inter1), .O(G398));
nand2 gate78( .a(G6), .b(G320), .O(G399) );

  xor2  gate2647(.a(G323), .b(G10), .O(gate79inter0));
  nand2 gate2648(.a(gate79inter0), .b(s_300), .O(gate79inter1));
  and2  gate2649(.a(G323), .b(G10), .O(gate79inter2));
  inv1  gate2650(.a(s_300), .O(gate79inter3));
  inv1  gate2651(.a(s_301), .O(gate79inter4));
  nand2 gate2652(.a(gate79inter4), .b(gate79inter3), .O(gate79inter5));
  nor2  gate2653(.a(gate79inter5), .b(gate79inter2), .O(gate79inter6));
  inv1  gate2654(.a(G10), .O(gate79inter7));
  inv1  gate2655(.a(G323), .O(gate79inter8));
  nand2 gate2656(.a(gate79inter8), .b(gate79inter7), .O(gate79inter9));
  nand2 gate2657(.a(s_301), .b(gate79inter3), .O(gate79inter10));
  nor2  gate2658(.a(gate79inter10), .b(gate79inter9), .O(gate79inter11));
  nor2  gate2659(.a(gate79inter11), .b(gate79inter6), .O(gate79inter12));
  nand2 gate2660(.a(gate79inter12), .b(gate79inter1), .O(G400));
nand2 gate80( .a(G14), .b(G323), .O(G401) );
nand2 gate81( .a(G3), .b(G326), .O(G402) );
nand2 gate82( .a(G7), .b(G326), .O(G403) );

  xor2  gate1009(.a(G329), .b(G11), .O(gate83inter0));
  nand2 gate1010(.a(gate83inter0), .b(s_66), .O(gate83inter1));
  and2  gate1011(.a(G329), .b(G11), .O(gate83inter2));
  inv1  gate1012(.a(s_66), .O(gate83inter3));
  inv1  gate1013(.a(s_67), .O(gate83inter4));
  nand2 gate1014(.a(gate83inter4), .b(gate83inter3), .O(gate83inter5));
  nor2  gate1015(.a(gate83inter5), .b(gate83inter2), .O(gate83inter6));
  inv1  gate1016(.a(G11), .O(gate83inter7));
  inv1  gate1017(.a(G329), .O(gate83inter8));
  nand2 gate1018(.a(gate83inter8), .b(gate83inter7), .O(gate83inter9));
  nand2 gate1019(.a(s_67), .b(gate83inter3), .O(gate83inter10));
  nor2  gate1020(.a(gate83inter10), .b(gate83inter9), .O(gate83inter11));
  nor2  gate1021(.a(gate83inter11), .b(gate83inter6), .O(gate83inter12));
  nand2 gate1022(.a(gate83inter12), .b(gate83inter1), .O(G404));
nand2 gate84( .a(G15), .b(G329), .O(G405) );
nand2 gate85( .a(G4), .b(G332), .O(G406) );

  xor2  gate659(.a(G332), .b(G8), .O(gate86inter0));
  nand2 gate660(.a(gate86inter0), .b(s_16), .O(gate86inter1));
  and2  gate661(.a(G332), .b(G8), .O(gate86inter2));
  inv1  gate662(.a(s_16), .O(gate86inter3));
  inv1  gate663(.a(s_17), .O(gate86inter4));
  nand2 gate664(.a(gate86inter4), .b(gate86inter3), .O(gate86inter5));
  nor2  gate665(.a(gate86inter5), .b(gate86inter2), .O(gate86inter6));
  inv1  gate666(.a(G8), .O(gate86inter7));
  inv1  gate667(.a(G332), .O(gate86inter8));
  nand2 gate668(.a(gate86inter8), .b(gate86inter7), .O(gate86inter9));
  nand2 gate669(.a(s_17), .b(gate86inter3), .O(gate86inter10));
  nor2  gate670(.a(gate86inter10), .b(gate86inter9), .O(gate86inter11));
  nor2  gate671(.a(gate86inter11), .b(gate86inter6), .O(gate86inter12));
  nand2 gate672(.a(gate86inter12), .b(gate86inter1), .O(G407));
nand2 gate87( .a(G12), .b(G335), .O(G408) );
nand2 gate88( .a(G16), .b(G335), .O(G409) );
nand2 gate89( .a(G17), .b(G338), .O(G410) );
nand2 gate90( .a(G21), .b(G338), .O(G411) );

  xor2  gate1023(.a(G341), .b(G25), .O(gate91inter0));
  nand2 gate1024(.a(gate91inter0), .b(s_68), .O(gate91inter1));
  and2  gate1025(.a(G341), .b(G25), .O(gate91inter2));
  inv1  gate1026(.a(s_68), .O(gate91inter3));
  inv1  gate1027(.a(s_69), .O(gate91inter4));
  nand2 gate1028(.a(gate91inter4), .b(gate91inter3), .O(gate91inter5));
  nor2  gate1029(.a(gate91inter5), .b(gate91inter2), .O(gate91inter6));
  inv1  gate1030(.a(G25), .O(gate91inter7));
  inv1  gate1031(.a(G341), .O(gate91inter8));
  nand2 gate1032(.a(gate91inter8), .b(gate91inter7), .O(gate91inter9));
  nand2 gate1033(.a(s_69), .b(gate91inter3), .O(gate91inter10));
  nor2  gate1034(.a(gate91inter10), .b(gate91inter9), .O(gate91inter11));
  nor2  gate1035(.a(gate91inter11), .b(gate91inter6), .O(gate91inter12));
  nand2 gate1036(.a(gate91inter12), .b(gate91inter1), .O(G412));
nand2 gate92( .a(G29), .b(G341), .O(G413) );
nand2 gate93( .a(G18), .b(G344), .O(G414) );

  xor2  gate1303(.a(G344), .b(G22), .O(gate94inter0));
  nand2 gate1304(.a(gate94inter0), .b(s_108), .O(gate94inter1));
  and2  gate1305(.a(G344), .b(G22), .O(gate94inter2));
  inv1  gate1306(.a(s_108), .O(gate94inter3));
  inv1  gate1307(.a(s_109), .O(gate94inter4));
  nand2 gate1308(.a(gate94inter4), .b(gate94inter3), .O(gate94inter5));
  nor2  gate1309(.a(gate94inter5), .b(gate94inter2), .O(gate94inter6));
  inv1  gate1310(.a(G22), .O(gate94inter7));
  inv1  gate1311(.a(G344), .O(gate94inter8));
  nand2 gate1312(.a(gate94inter8), .b(gate94inter7), .O(gate94inter9));
  nand2 gate1313(.a(s_109), .b(gate94inter3), .O(gate94inter10));
  nor2  gate1314(.a(gate94inter10), .b(gate94inter9), .O(gate94inter11));
  nor2  gate1315(.a(gate94inter11), .b(gate94inter6), .O(gate94inter12));
  nand2 gate1316(.a(gate94inter12), .b(gate94inter1), .O(G415));

  xor2  gate1415(.a(G347), .b(G26), .O(gate95inter0));
  nand2 gate1416(.a(gate95inter0), .b(s_124), .O(gate95inter1));
  and2  gate1417(.a(G347), .b(G26), .O(gate95inter2));
  inv1  gate1418(.a(s_124), .O(gate95inter3));
  inv1  gate1419(.a(s_125), .O(gate95inter4));
  nand2 gate1420(.a(gate95inter4), .b(gate95inter3), .O(gate95inter5));
  nor2  gate1421(.a(gate95inter5), .b(gate95inter2), .O(gate95inter6));
  inv1  gate1422(.a(G26), .O(gate95inter7));
  inv1  gate1423(.a(G347), .O(gate95inter8));
  nand2 gate1424(.a(gate95inter8), .b(gate95inter7), .O(gate95inter9));
  nand2 gate1425(.a(s_125), .b(gate95inter3), .O(gate95inter10));
  nor2  gate1426(.a(gate95inter10), .b(gate95inter9), .O(gate95inter11));
  nor2  gate1427(.a(gate95inter11), .b(gate95inter6), .O(gate95inter12));
  nand2 gate1428(.a(gate95inter12), .b(gate95inter1), .O(G416));
nand2 gate96( .a(G30), .b(G347), .O(G417) );

  xor2  gate1625(.a(G350), .b(G19), .O(gate97inter0));
  nand2 gate1626(.a(gate97inter0), .b(s_154), .O(gate97inter1));
  and2  gate1627(.a(G350), .b(G19), .O(gate97inter2));
  inv1  gate1628(.a(s_154), .O(gate97inter3));
  inv1  gate1629(.a(s_155), .O(gate97inter4));
  nand2 gate1630(.a(gate97inter4), .b(gate97inter3), .O(gate97inter5));
  nor2  gate1631(.a(gate97inter5), .b(gate97inter2), .O(gate97inter6));
  inv1  gate1632(.a(G19), .O(gate97inter7));
  inv1  gate1633(.a(G350), .O(gate97inter8));
  nand2 gate1634(.a(gate97inter8), .b(gate97inter7), .O(gate97inter9));
  nand2 gate1635(.a(s_155), .b(gate97inter3), .O(gate97inter10));
  nor2  gate1636(.a(gate97inter10), .b(gate97inter9), .O(gate97inter11));
  nor2  gate1637(.a(gate97inter11), .b(gate97inter6), .O(gate97inter12));
  nand2 gate1638(.a(gate97inter12), .b(gate97inter1), .O(G418));

  xor2  gate1037(.a(G350), .b(G23), .O(gate98inter0));
  nand2 gate1038(.a(gate98inter0), .b(s_70), .O(gate98inter1));
  and2  gate1039(.a(G350), .b(G23), .O(gate98inter2));
  inv1  gate1040(.a(s_70), .O(gate98inter3));
  inv1  gate1041(.a(s_71), .O(gate98inter4));
  nand2 gate1042(.a(gate98inter4), .b(gate98inter3), .O(gate98inter5));
  nor2  gate1043(.a(gate98inter5), .b(gate98inter2), .O(gate98inter6));
  inv1  gate1044(.a(G23), .O(gate98inter7));
  inv1  gate1045(.a(G350), .O(gate98inter8));
  nand2 gate1046(.a(gate98inter8), .b(gate98inter7), .O(gate98inter9));
  nand2 gate1047(.a(s_71), .b(gate98inter3), .O(gate98inter10));
  nor2  gate1048(.a(gate98inter10), .b(gate98inter9), .O(gate98inter11));
  nor2  gate1049(.a(gate98inter11), .b(gate98inter6), .O(gate98inter12));
  nand2 gate1050(.a(gate98inter12), .b(gate98inter1), .O(G419));
nand2 gate99( .a(G27), .b(G353), .O(G420) );

  xor2  gate1401(.a(G353), .b(G31), .O(gate100inter0));
  nand2 gate1402(.a(gate100inter0), .b(s_122), .O(gate100inter1));
  and2  gate1403(.a(G353), .b(G31), .O(gate100inter2));
  inv1  gate1404(.a(s_122), .O(gate100inter3));
  inv1  gate1405(.a(s_123), .O(gate100inter4));
  nand2 gate1406(.a(gate100inter4), .b(gate100inter3), .O(gate100inter5));
  nor2  gate1407(.a(gate100inter5), .b(gate100inter2), .O(gate100inter6));
  inv1  gate1408(.a(G31), .O(gate100inter7));
  inv1  gate1409(.a(G353), .O(gate100inter8));
  nand2 gate1410(.a(gate100inter8), .b(gate100inter7), .O(gate100inter9));
  nand2 gate1411(.a(s_123), .b(gate100inter3), .O(gate100inter10));
  nor2  gate1412(.a(gate100inter10), .b(gate100inter9), .O(gate100inter11));
  nor2  gate1413(.a(gate100inter11), .b(gate100inter6), .O(gate100inter12));
  nand2 gate1414(.a(gate100inter12), .b(gate100inter1), .O(G421));
nand2 gate101( .a(G20), .b(G356), .O(G422) );
nand2 gate102( .a(G24), .b(G356), .O(G423) );
nand2 gate103( .a(G28), .b(G359), .O(G424) );
nand2 gate104( .a(G32), .b(G359), .O(G425) );
nand2 gate105( .a(G362), .b(G363), .O(G426) );

  xor2  gate715(.a(G365), .b(G364), .O(gate106inter0));
  nand2 gate716(.a(gate106inter0), .b(s_24), .O(gate106inter1));
  and2  gate717(.a(G365), .b(G364), .O(gate106inter2));
  inv1  gate718(.a(s_24), .O(gate106inter3));
  inv1  gate719(.a(s_25), .O(gate106inter4));
  nand2 gate720(.a(gate106inter4), .b(gate106inter3), .O(gate106inter5));
  nor2  gate721(.a(gate106inter5), .b(gate106inter2), .O(gate106inter6));
  inv1  gate722(.a(G364), .O(gate106inter7));
  inv1  gate723(.a(G365), .O(gate106inter8));
  nand2 gate724(.a(gate106inter8), .b(gate106inter7), .O(gate106inter9));
  nand2 gate725(.a(s_25), .b(gate106inter3), .O(gate106inter10));
  nor2  gate726(.a(gate106inter10), .b(gate106inter9), .O(gate106inter11));
  nor2  gate727(.a(gate106inter11), .b(gate106inter6), .O(gate106inter12));
  nand2 gate728(.a(gate106inter12), .b(gate106inter1), .O(G429));
nand2 gate107( .a(G366), .b(G367), .O(G432) );

  xor2  gate2297(.a(G369), .b(G368), .O(gate108inter0));
  nand2 gate2298(.a(gate108inter0), .b(s_250), .O(gate108inter1));
  and2  gate2299(.a(G369), .b(G368), .O(gate108inter2));
  inv1  gate2300(.a(s_250), .O(gate108inter3));
  inv1  gate2301(.a(s_251), .O(gate108inter4));
  nand2 gate2302(.a(gate108inter4), .b(gate108inter3), .O(gate108inter5));
  nor2  gate2303(.a(gate108inter5), .b(gate108inter2), .O(gate108inter6));
  inv1  gate2304(.a(G368), .O(gate108inter7));
  inv1  gate2305(.a(G369), .O(gate108inter8));
  nand2 gate2306(.a(gate108inter8), .b(gate108inter7), .O(gate108inter9));
  nand2 gate2307(.a(s_251), .b(gate108inter3), .O(gate108inter10));
  nor2  gate2308(.a(gate108inter10), .b(gate108inter9), .O(gate108inter11));
  nor2  gate2309(.a(gate108inter11), .b(gate108inter6), .O(gate108inter12));
  nand2 gate2310(.a(gate108inter12), .b(gate108inter1), .O(G435));
nand2 gate109( .a(G370), .b(G371), .O(G438) );
nand2 gate110( .a(G372), .b(G373), .O(G441) );

  xor2  gate981(.a(G375), .b(G374), .O(gate111inter0));
  nand2 gate982(.a(gate111inter0), .b(s_62), .O(gate111inter1));
  and2  gate983(.a(G375), .b(G374), .O(gate111inter2));
  inv1  gate984(.a(s_62), .O(gate111inter3));
  inv1  gate985(.a(s_63), .O(gate111inter4));
  nand2 gate986(.a(gate111inter4), .b(gate111inter3), .O(gate111inter5));
  nor2  gate987(.a(gate111inter5), .b(gate111inter2), .O(gate111inter6));
  inv1  gate988(.a(G374), .O(gate111inter7));
  inv1  gate989(.a(G375), .O(gate111inter8));
  nand2 gate990(.a(gate111inter8), .b(gate111inter7), .O(gate111inter9));
  nand2 gate991(.a(s_63), .b(gate111inter3), .O(gate111inter10));
  nor2  gate992(.a(gate111inter10), .b(gate111inter9), .O(gate111inter11));
  nor2  gate993(.a(gate111inter11), .b(gate111inter6), .O(gate111inter12));
  nand2 gate994(.a(gate111inter12), .b(gate111inter1), .O(G444));

  xor2  gate1723(.a(G377), .b(G376), .O(gate112inter0));
  nand2 gate1724(.a(gate112inter0), .b(s_168), .O(gate112inter1));
  and2  gate1725(.a(G377), .b(G376), .O(gate112inter2));
  inv1  gate1726(.a(s_168), .O(gate112inter3));
  inv1  gate1727(.a(s_169), .O(gate112inter4));
  nand2 gate1728(.a(gate112inter4), .b(gate112inter3), .O(gate112inter5));
  nor2  gate1729(.a(gate112inter5), .b(gate112inter2), .O(gate112inter6));
  inv1  gate1730(.a(G376), .O(gate112inter7));
  inv1  gate1731(.a(G377), .O(gate112inter8));
  nand2 gate1732(.a(gate112inter8), .b(gate112inter7), .O(gate112inter9));
  nand2 gate1733(.a(s_169), .b(gate112inter3), .O(gate112inter10));
  nor2  gate1734(.a(gate112inter10), .b(gate112inter9), .O(gate112inter11));
  nor2  gate1735(.a(gate112inter11), .b(gate112inter6), .O(gate112inter12));
  nand2 gate1736(.a(gate112inter12), .b(gate112inter1), .O(G447));

  xor2  gate939(.a(G379), .b(G378), .O(gate113inter0));
  nand2 gate940(.a(gate113inter0), .b(s_56), .O(gate113inter1));
  and2  gate941(.a(G379), .b(G378), .O(gate113inter2));
  inv1  gate942(.a(s_56), .O(gate113inter3));
  inv1  gate943(.a(s_57), .O(gate113inter4));
  nand2 gate944(.a(gate113inter4), .b(gate113inter3), .O(gate113inter5));
  nor2  gate945(.a(gate113inter5), .b(gate113inter2), .O(gate113inter6));
  inv1  gate946(.a(G378), .O(gate113inter7));
  inv1  gate947(.a(G379), .O(gate113inter8));
  nand2 gate948(.a(gate113inter8), .b(gate113inter7), .O(gate113inter9));
  nand2 gate949(.a(s_57), .b(gate113inter3), .O(gate113inter10));
  nor2  gate950(.a(gate113inter10), .b(gate113inter9), .O(gate113inter11));
  nor2  gate951(.a(gate113inter11), .b(gate113inter6), .O(gate113inter12));
  nand2 gate952(.a(gate113inter12), .b(gate113inter1), .O(G450));
nand2 gate114( .a(G380), .b(G381), .O(G453) );

  xor2  gate827(.a(G383), .b(G382), .O(gate115inter0));
  nand2 gate828(.a(gate115inter0), .b(s_40), .O(gate115inter1));
  and2  gate829(.a(G383), .b(G382), .O(gate115inter2));
  inv1  gate830(.a(s_40), .O(gate115inter3));
  inv1  gate831(.a(s_41), .O(gate115inter4));
  nand2 gate832(.a(gate115inter4), .b(gate115inter3), .O(gate115inter5));
  nor2  gate833(.a(gate115inter5), .b(gate115inter2), .O(gate115inter6));
  inv1  gate834(.a(G382), .O(gate115inter7));
  inv1  gate835(.a(G383), .O(gate115inter8));
  nand2 gate836(.a(gate115inter8), .b(gate115inter7), .O(gate115inter9));
  nand2 gate837(.a(s_41), .b(gate115inter3), .O(gate115inter10));
  nor2  gate838(.a(gate115inter10), .b(gate115inter9), .O(gate115inter11));
  nor2  gate839(.a(gate115inter11), .b(gate115inter6), .O(gate115inter12));
  nand2 gate840(.a(gate115inter12), .b(gate115inter1), .O(G456));
nand2 gate116( .a(G384), .b(G385), .O(G459) );

  xor2  gate1051(.a(G387), .b(G386), .O(gate117inter0));
  nand2 gate1052(.a(gate117inter0), .b(s_72), .O(gate117inter1));
  and2  gate1053(.a(G387), .b(G386), .O(gate117inter2));
  inv1  gate1054(.a(s_72), .O(gate117inter3));
  inv1  gate1055(.a(s_73), .O(gate117inter4));
  nand2 gate1056(.a(gate117inter4), .b(gate117inter3), .O(gate117inter5));
  nor2  gate1057(.a(gate117inter5), .b(gate117inter2), .O(gate117inter6));
  inv1  gate1058(.a(G386), .O(gate117inter7));
  inv1  gate1059(.a(G387), .O(gate117inter8));
  nand2 gate1060(.a(gate117inter8), .b(gate117inter7), .O(gate117inter9));
  nand2 gate1061(.a(s_73), .b(gate117inter3), .O(gate117inter10));
  nor2  gate1062(.a(gate117inter10), .b(gate117inter9), .O(gate117inter11));
  nor2  gate1063(.a(gate117inter11), .b(gate117inter6), .O(gate117inter12));
  nand2 gate1064(.a(gate117inter12), .b(gate117inter1), .O(G462));
nand2 gate118( .a(G388), .b(G389), .O(G465) );

  xor2  gate1149(.a(G391), .b(G390), .O(gate119inter0));
  nand2 gate1150(.a(gate119inter0), .b(s_86), .O(gate119inter1));
  and2  gate1151(.a(G391), .b(G390), .O(gate119inter2));
  inv1  gate1152(.a(s_86), .O(gate119inter3));
  inv1  gate1153(.a(s_87), .O(gate119inter4));
  nand2 gate1154(.a(gate119inter4), .b(gate119inter3), .O(gate119inter5));
  nor2  gate1155(.a(gate119inter5), .b(gate119inter2), .O(gate119inter6));
  inv1  gate1156(.a(G390), .O(gate119inter7));
  inv1  gate1157(.a(G391), .O(gate119inter8));
  nand2 gate1158(.a(gate119inter8), .b(gate119inter7), .O(gate119inter9));
  nand2 gate1159(.a(s_87), .b(gate119inter3), .O(gate119inter10));
  nor2  gate1160(.a(gate119inter10), .b(gate119inter9), .O(gate119inter11));
  nor2  gate1161(.a(gate119inter11), .b(gate119inter6), .O(gate119inter12));
  nand2 gate1162(.a(gate119inter12), .b(gate119inter1), .O(G468));
nand2 gate120( .a(G392), .b(G393), .O(G471) );
nand2 gate121( .a(G394), .b(G395), .O(G474) );
nand2 gate122( .a(G396), .b(G397), .O(G477) );

  xor2  gate1765(.a(G399), .b(G398), .O(gate123inter0));
  nand2 gate1766(.a(gate123inter0), .b(s_174), .O(gate123inter1));
  and2  gate1767(.a(G399), .b(G398), .O(gate123inter2));
  inv1  gate1768(.a(s_174), .O(gate123inter3));
  inv1  gate1769(.a(s_175), .O(gate123inter4));
  nand2 gate1770(.a(gate123inter4), .b(gate123inter3), .O(gate123inter5));
  nor2  gate1771(.a(gate123inter5), .b(gate123inter2), .O(gate123inter6));
  inv1  gate1772(.a(G398), .O(gate123inter7));
  inv1  gate1773(.a(G399), .O(gate123inter8));
  nand2 gate1774(.a(gate123inter8), .b(gate123inter7), .O(gate123inter9));
  nand2 gate1775(.a(s_175), .b(gate123inter3), .O(gate123inter10));
  nor2  gate1776(.a(gate123inter10), .b(gate123inter9), .O(gate123inter11));
  nor2  gate1777(.a(gate123inter11), .b(gate123inter6), .O(gate123inter12));
  nand2 gate1778(.a(gate123inter12), .b(gate123inter1), .O(G480));
nand2 gate124( .a(G400), .b(G401), .O(G483) );
nand2 gate125( .a(G402), .b(G403), .O(G486) );
nand2 gate126( .a(G404), .b(G405), .O(G489) );
nand2 gate127( .a(G406), .b(G407), .O(G492) );
nand2 gate128( .a(G408), .b(G409), .O(G495) );
nand2 gate129( .a(G410), .b(G411), .O(G498) );
nand2 gate130( .a(G412), .b(G413), .O(G501) );

  xor2  gate1863(.a(G415), .b(G414), .O(gate131inter0));
  nand2 gate1864(.a(gate131inter0), .b(s_188), .O(gate131inter1));
  and2  gate1865(.a(G415), .b(G414), .O(gate131inter2));
  inv1  gate1866(.a(s_188), .O(gate131inter3));
  inv1  gate1867(.a(s_189), .O(gate131inter4));
  nand2 gate1868(.a(gate131inter4), .b(gate131inter3), .O(gate131inter5));
  nor2  gate1869(.a(gate131inter5), .b(gate131inter2), .O(gate131inter6));
  inv1  gate1870(.a(G414), .O(gate131inter7));
  inv1  gate1871(.a(G415), .O(gate131inter8));
  nand2 gate1872(.a(gate131inter8), .b(gate131inter7), .O(gate131inter9));
  nand2 gate1873(.a(s_189), .b(gate131inter3), .O(gate131inter10));
  nor2  gate1874(.a(gate131inter10), .b(gate131inter9), .O(gate131inter11));
  nor2  gate1875(.a(gate131inter11), .b(gate131inter6), .O(gate131inter12));
  nand2 gate1876(.a(gate131inter12), .b(gate131inter1), .O(G504));
nand2 gate132( .a(G416), .b(G417), .O(G507) );

  xor2  gate1835(.a(G419), .b(G418), .O(gate133inter0));
  nand2 gate1836(.a(gate133inter0), .b(s_184), .O(gate133inter1));
  and2  gate1837(.a(G419), .b(G418), .O(gate133inter2));
  inv1  gate1838(.a(s_184), .O(gate133inter3));
  inv1  gate1839(.a(s_185), .O(gate133inter4));
  nand2 gate1840(.a(gate133inter4), .b(gate133inter3), .O(gate133inter5));
  nor2  gate1841(.a(gate133inter5), .b(gate133inter2), .O(gate133inter6));
  inv1  gate1842(.a(G418), .O(gate133inter7));
  inv1  gate1843(.a(G419), .O(gate133inter8));
  nand2 gate1844(.a(gate133inter8), .b(gate133inter7), .O(gate133inter9));
  nand2 gate1845(.a(s_185), .b(gate133inter3), .O(gate133inter10));
  nor2  gate1846(.a(gate133inter10), .b(gate133inter9), .O(gate133inter11));
  nor2  gate1847(.a(gate133inter11), .b(gate133inter6), .O(gate133inter12));
  nand2 gate1848(.a(gate133inter12), .b(gate133inter1), .O(G510));
nand2 gate134( .a(G420), .b(G421), .O(G513) );
nand2 gate135( .a(G422), .b(G423), .O(G516) );
nand2 gate136( .a(G424), .b(G425), .O(G519) );

  xor2  gate855(.a(G429), .b(G426), .O(gate137inter0));
  nand2 gate856(.a(gate137inter0), .b(s_44), .O(gate137inter1));
  and2  gate857(.a(G429), .b(G426), .O(gate137inter2));
  inv1  gate858(.a(s_44), .O(gate137inter3));
  inv1  gate859(.a(s_45), .O(gate137inter4));
  nand2 gate860(.a(gate137inter4), .b(gate137inter3), .O(gate137inter5));
  nor2  gate861(.a(gate137inter5), .b(gate137inter2), .O(gate137inter6));
  inv1  gate862(.a(G426), .O(gate137inter7));
  inv1  gate863(.a(G429), .O(gate137inter8));
  nand2 gate864(.a(gate137inter8), .b(gate137inter7), .O(gate137inter9));
  nand2 gate865(.a(s_45), .b(gate137inter3), .O(gate137inter10));
  nor2  gate866(.a(gate137inter10), .b(gate137inter9), .O(gate137inter11));
  nor2  gate867(.a(gate137inter11), .b(gate137inter6), .O(gate137inter12));
  nand2 gate868(.a(gate137inter12), .b(gate137inter1), .O(G522));
nand2 gate138( .a(G432), .b(G435), .O(G525) );

  xor2  gate2143(.a(G441), .b(G438), .O(gate139inter0));
  nand2 gate2144(.a(gate139inter0), .b(s_228), .O(gate139inter1));
  and2  gate2145(.a(G441), .b(G438), .O(gate139inter2));
  inv1  gate2146(.a(s_228), .O(gate139inter3));
  inv1  gate2147(.a(s_229), .O(gate139inter4));
  nand2 gate2148(.a(gate139inter4), .b(gate139inter3), .O(gate139inter5));
  nor2  gate2149(.a(gate139inter5), .b(gate139inter2), .O(gate139inter6));
  inv1  gate2150(.a(G438), .O(gate139inter7));
  inv1  gate2151(.a(G441), .O(gate139inter8));
  nand2 gate2152(.a(gate139inter8), .b(gate139inter7), .O(gate139inter9));
  nand2 gate2153(.a(s_229), .b(gate139inter3), .O(gate139inter10));
  nor2  gate2154(.a(gate139inter10), .b(gate139inter9), .O(gate139inter11));
  nor2  gate2155(.a(gate139inter11), .b(gate139inter6), .O(gate139inter12));
  nand2 gate2156(.a(gate139inter12), .b(gate139inter1), .O(G528));

  xor2  gate1387(.a(G447), .b(G444), .O(gate140inter0));
  nand2 gate1388(.a(gate140inter0), .b(s_120), .O(gate140inter1));
  and2  gate1389(.a(G447), .b(G444), .O(gate140inter2));
  inv1  gate1390(.a(s_120), .O(gate140inter3));
  inv1  gate1391(.a(s_121), .O(gate140inter4));
  nand2 gate1392(.a(gate140inter4), .b(gate140inter3), .O(gate140inter5));
  nor2  gate1393(.a(gate140inter5), .b(gate140inter2), .O(gate140inter6));
  inv1  gate1394(.a(G444), .O(gate140inter7));
  inv1  gate1395(.a(G447), .O(gate140inter8));
  nand2 gate1396(.a(gate140inter8), .b(gate140inter7), .O(gate140inter9));
  nand2 gate1397(.a(s_121), .b(gate140inter3), .O(gate140inter10));
  nor2  gate1398(.a(gate140inter10), .b(gate140inter9), .O(gate140inter11));
  nor2  gate1399(.a(gate140inter11), .b(gate140inter6), .O(gate140inter12));
  nand2 gate1400(.a(gate140inter12), .b(gate140inter1), .O(G531));
nand2 gate141( .a(G450), .b(G453), .O(G534) );
nand2 gate142( .a(G456), .b(G459), .O(G537) );
nand2 gate143( .a(G462), .b(G465), .O(G540) );
nand2 gate144( .a(G468), .b(G471), .O(G543) );
nand2 gate145( .a(G474), .b(G477), .O(G546) );
nand2 gate146( .a(G480), .b(G483), .O(G549) );
nand2 gate147( .a(G486), .b(G489), .O(G552) );
nand2 gate148( .a(G492), .b(G495), .O(G555) );
nand2 gate149( .a(G498), .b(G501), .O(G558) );
nand2 gate150( .a(G504), .b(G507), .O(G561) );
nand2 gate151( .a(G510), .b(G513), .O(G564) );
nand2 gate152( .a(G516), .b(G519), .O(G567) );

  xor2  gate1205(.a(G522), .b(G426), .O(gate153inter0));
  nand2 gate1206(.a(gate153inter0), .b(s_94), .O(gate153inter1));
  and2  gate1207(.a(G522), .b(G426), .O(gate153inter2));
  inv1  gate1208(.a(s_94), .O(gate153inter3));
  inv1  gate1209(.a(s_95), .O(gate153inter4));
  nand2 gate1210(.a(gate153inter4), .b(gate153inter3), .O(gate153inter5));
  nor2  gate1211(.a(gate153inter5), .b(gate153inter2), .O(gate153inter6));
  inv1  gate1212(.a(G426), .O(gate153inter7));
  inv1  gate1213(.a(G522), .O(gate153inter8));
  nand2 gate1214(.a(gate153inter8), .b(gate153inter7), .O(gate153inter9));
  nand2 gate1215(.a(s_95), .b(gate153inter3), .O(gate153inter10));
  nor2  gate1216(.a(gate153inter10), .b(gate153inter9), .O(gate153inter11));
  nor2  gate1217(.a(gate153inter11), .b(gate153inter6), .O(gate153inter12));
  nand2 gate1218(.a(gate153inter12), .b(gate153inter1), .O(G570));
nand2 gate154( .a(G429), .b(G522), .O(G571) );
nand2 gate155( .a(G432), .b(G525), .O(G572) );
nand2 gate156( .a(G435), .b(G525), .O(G573) );
nand2 gate157( .a(G438), .b(G528), .O(G574) );

  xor2  gate1583(.a(G528), .b(G441), .O(gate158inter0));
  nand2 gate1584(.a(gate158inter0), .b(s_148), .O(gate158inter1));
  and2  gate1585(.a(G528), .b(G441), .O(gate158inter2));
  inv1  gate1586(.a(s_148), .O(gate158inter3));
  inv1  gate1587(.a(s_149), .O(gate158inter4));
  nand2 gate1588(.a(gate158inter4), .b(gate158inter3), .O(gate158inter5));
  nor2  gate1589(.a(gate158inter5), .b(gate158inter2), .O(gate158inter6));
  inv1  gate1590(.a(G441), .O(gate158inter7));
  inv1  gate1591(.a(G528), .O(gate158inter8));
  nand2 gate1592(.a(gate158inter8), .b(gate158inter7), .O(gate158inter9));
  nand2 gate1593(.a(s_149), .b(gate158inter3), .O(gate158inter10));
  nor2  gate1594(.a(gate158inter10), .b(gate158inter9), .O(gate158inter11));
  nor2  gate1595(.a(gate158inter11), .b(gate158inter6), .O(gate158inter12));
  nand2 gate1596(.a(gate158inter12), .b(gate158inter1), .O(G575));

  xor2  gate2577(.a(G531), .b(G444), .O(gate159inter0));
  nand2 gate2578(.a(gate159inter0), .b(s_290), .O(gate159inter1));
  and2  gate2579(.a(G531), .b(G444), .O(gate159inter2));
  inv1  gate2580(.a(s_290), .O(gate159inter3));
  inv1  gate2581(.a(s_291), .O(gate159inter4));
  nand2 gate2582(.a(gate159inter4), .b(gate159inter3), .O(gate159inter5));
  nor2  gate2583(.a(gate159inter5), .b(gate159inter2), .O(gate159inter6));
  inv1  gate2584(.a(G444), .O(gate159inter7));
  inv1  gate2585(.a(G531), .O(gate159inter8));
  nand2 gate2586(.a(gate159inter8), .b(gate159inter7), .O(gate159inter9));
  nand2 gate2587(.a(s_291), .b(gate159inter3), .O(gate159inter10));
  nor2  gate2588(.a(gate159inter10), .b(gate159inter9), .O(gate159inter11));
  nor2  gate2589(.a(gate159inter11), .b(gate159inter6), .O(gate159inter12));
  nand2 gate2590(.a(gate159inter12), .b(gate159inter1), .O(G576));
nand2 gate160( .a(G447), .b(G531), .O(G577) );
nand2 gate161( .a(G450), .b(G534), .O(G578) );
nand2 gate162( .a(G453), .b(G534), .O(G579) );
nand2 gate163( .a(G456), .b(G537), .O(G580) );

  xor2  gate561(.a(G537), .b(G459), .O(gate164inter0));
  nand2 gate562(.a(gate164inter0), .b(s_2), .O(gate164inter1));
  and2  gate563(.a(G537), .b(G459), .O(gate164inter2));
  inv1  gate564(.a(s_2), .O(gate164inter3));
  inv1  gate565(.a(s_3), .O(gate164inter4));
  nand2 gate566(.a(gate164inter4), .b(gate164inter3), .O(gate164inter5));
  nor2  gate567(.a(gate164inter5), .b(gate164inter2), .O(gate164inter6));
  inv1  gate568(.a(G459), .O(gate164inter7));
  inv1  gate569(.a(G537), .O(gate164inter8));
  nand2 gate570(.a(gate164inter8), .b(gate164inter7), .O(gate164inter9));
  nand2 gate571(.a(s_3), .b(gate164inter3), .O(gate164inter10));
  nor2  gate572(.a(gate164inter10), .b(gate164inter9), .O(gate164inter11));
  nor2  gate573(.a(gate164inter11), .b(gate164inter6), .O(gate164inter12));
  nand2 gate574(.a(gate164inter12), .b(gate164inter1), .O(G581));
nand2 gate165( .a(G462), .b(G540), .O(G582) );
nand2 gate166( .a(G465), .b(G540), .O(G583) );
nand2 gate167( .a(G468), .b(G543), .O(G584) );
nand2 gate168( .a(G471), .b(G543), .O(G585) );
nand2 gate169( .a(G474), .b(G546), .O(G586) );
nand2 gate170( .a(G477), .b(G546), .O(G587) );
nand2 gate171( .a(G480), .b(G549), .O(G588) );

  xor2  gate645(.a(G549), .b(G483), .O(gate172inter0));
  nand2 gate646(.a(gate172inter0), .b(s_14), .O(gate172inter1));
  and2  gate647(.a(G549), .b(G483), .O(gate172inter2));
  inv1  gate648(.a(s_14), .O(gate172inter3));
  inv1  gate649(.a(s_15), .O(gate172inter4));
  nand2 gate650(.a(gate172inter4), .b(gate172inter3), .O(gate172inter5));
  nor2  gate651(.a(gate172inter5), .b(gate172inter2), .O(gate172inter6));
  inv1  gate652(.a(G483), .O(gate172inter7));
  inv1  gate653(.a(G549), .O(gate172inter8));
  nand2 gate654(.a(gate172inter8), .b(gate172inter7), .O(gate172inter9));
  nand2 gate655(.a(s_15), .b(gate172inter3), .O(gate172inter10));
  nor2  gate656(.a(gate172inter10), .b(gate172inter9), .O(gate172inter11));
  nor2  gate657(.a(gate172inter11), .b(gate172inter6), .O(gate172inter12));
  nand2 gate658(.a(gate172inter12), .b(gate172inter1), .O(G589));
nand2 gate173( .a(G486), .b(G552), .O(G590) );

  xor2  gate1121(.a(G552), .b(G489), .O(gate174inter0));
  nand2 gate1122(.a(gate174inter0), .b(s_82), .O(gate174inter1));
  and2  gate1123(.a(G552), .b(G489), .O(gate174inter2));
  inv1  gate1124(.a(s_82), .O(gate174inter3));
  inv1  gate1125(.a(s_83), .O(gate174inter4));
  nand2 gate1126(.a(gate174inter4), .b(gate174inter3), .O(gate174inter5));
  nor2  gate1127(.a(gate174inter5), .b(gate174inter2), .O(gate174inter6));
  inv1  gate1128(.a(G489), .O(gate174inter7));
  inv1  gate1129(.a(G552), .O(gate174inter8));
  nand2 gate1130(.a(gate174inter8), .b(gate174inter7), .O(gate174inter9));
  nand2 gate1131(.a(s_83), .b(gate174inter3), .O(gate174inter10));
  nor2  gate1132(.a(gate174inter10), .b(gate174inter9), .O(gate174inter11));
  nor2  gate1133(.a(gate174inter11), .b(gate174inter6), .O(gate174inter12));
  nand2 gate1134(.a(gate174inter12), .b(gate174inter1), .O(G591));
nand2 gate175( .a(G492), .b(G555), .O(G592) );
nand2 gate176( .a(G495), .b(G555), .O(G593) );
nand2 gate177( .a(G498), .b(G558), .O(G594) );
nand2 gate178( .a(G501), .b(G558), .O(G595) );
nand2 gate179( .a(G504), .b(G561), .O(G596) );

  xor2  gate1975(.a(G561), .b(G507), .O(gate180inter0));
  nand2 gate1976(.a(gate180inter0), .b(s_204), .O(gate180inter1));
  and2  gate1977(.a(G561), .b(G507), .O(gate180inter2));
  inv1  gate1978(.a(s_204), .O(gate180inter3));
  inv1  gate1979(.a(s_205), .O(gate180inter4));
  nand2 gate1980(.a(gate180inter4), .b(gate180inter3), .O(gate180inter5));
  nor2  gate1981(.a(gate180inter5), .b(gate180inter2), .O(gate180inter6));
  inv1  gate1982(.a(G507), .O(gate180inter7));
  inv1  gate1983(.a(G561), .O(gate180inter8));
  nand2 gate1984(.a(gate180inter8), .b(gate180inter7), .O(gate180inter9));
  nand2 gate1985(.a(s_205), .b(gate180inter3), .O(gate180inter10));
  nor2  gate1986(.a(gate180inter10), .b(gate180inter9), .O(gate180inter11));
  nor2  gate1987(.a(gate180inter11), .b(gate180inter6), .O(gate180inter12));
  nand2 gate1988(.a(gate180inter12), .b(gate180inter1), .O(G597));
nand2 gate181( .a(G510), .b(G564), .O(G598) );
nand2 gate182( .a(G513), .b(G564), .O(G599) );

  xor2  gate1485(.a(G567), .b(G516), .O(gate183inter0));
  nand2 gate1486(.a(gate183inter0), .b(s_134), .O(gate183inter1));
  and2  gate1487(.a(G567), .b(G516), .O(gate183inter2));
  inv1  gate1488(.a(s_134), .O(gate183inter3));
  inv1  gate1489(.a(s_135), .O(gate183inter4));
  nand2 gate1490(.a(gate183inter4), .b(gate183inter3), .O(gate183inter5));
  nor2  gate1491(.a(gate183inter5), .b(gate183inter2), .O(gate183inter6));
  inv1  gate1492(.a(G516), .O(gate183inter7));
  inv1  gate1493(.a(G567), .O(gate183inter8));
  nand2 gate1494(.a(gate183inter8), .b(gate183inter7), .O(gate183inter9));
  nand2 gate1495(.a(s_135), .b(gate183inter3), .O(gate183inter10));
  nor2  gate1496(.a(gate183inter10), .b(gate183inter9), .O(gate183inter11));
  nor2  gate1497(.a(gate183inter11), .b(gate183inter6), .O(gate183inter12));
  nand2 gate1498(.a(gate183inter12), .b(gate183inter1), .O(G600));

  xor2  gate2269(.a(G567), .b(G519), .O(gate184inter0));
  nand2 gate2270(.a(gate184inter0), .b(s_246), .O(gate184inter1));
  and2  gate2271(.a(G567), .b(G519), .O(gate184inter2));
  inv1  gate2272(.a(s_246), .O(gate184inter3));
  inv1  gate2273(.a(s_247), .O(gate184inter4));
  nand2 gate2274(.a(gate184inter4), .b(gate184inter3), .O(gate184inter5));
  nor2  gate2275(.a(gate184inter5), .b(gate184inter2), .O(gate184inter6));
  inv1  gate2276(.a(G519), .O(gate184inter7));
  inv1  gate2277(.a(G567), .O(gate184inter8));
  nand2 gate2278(.a(gate184inter8), .b(gate184inter7), .O(gate184inter9));
  nand2 gate2279(.a(s_247), .b(gate184inter3), .O(gate184inter10));
  nor2  gate2280(.a(gate184inter10), .b(gate184inter9), .O(gate184inter11));
  nor2  gate2281(.a(gate184inter11), .b(gate184inter6), .O(gate184inter12));
  nand2 gate2282(.a(gate184inter12), .b(gate184inter1), .O(G601));

  xor2  gate1597(.a(G571), .b(G570), .O(gate185inter0));
  nand2 gate1598(.a(gate185inter0), .b(s_150), .O(gate185inter1));
  and2  gate1599(.a(G571), .b(G570), .O(gate185inter2));
  inv1  gate1600(.a(s_150), .O(gate185inter3));
  inv1  gate1601(.a(s_151), .O(gate185inter4));
  nand2 gate1602(.a(gate185inter4), .b(gate185inter3), .O(gate185inter5));
  nor2  gate1603(.a(gate185inter5), .b(gate185inter2), .O(gate185inter6));
  inv1  gate1604(.a(G570), .O(gate185inter7));
  inv1  gate1605(.a(G571), .O(gate185inter8));
  nand2 gate1606(.a(gate185inter8), .b(gate185inter7), .O(gate185inter9));
  nand2 gate1607(.a(s_151), .b(gate185inter3), .O(gate185inter10));
  nor2  gate1608(.a(gate185inter10), .b(gate185inter9), .O(gate185inter11));
  nor2  gate1609(.a(gate185inter11), .b(gate185inter6), .O(gate185inter12));
  nand2 gate1610(.a(gate185inter12), .b(gate185inter1), .O(G602));
nand2 gate186( .a(G572), .b(G573), .O(G607) );
nand2 gate187( .a(G574), .b(G575), .O(G612) );

  xor2  gate1093(.a(G577), .b(G576), .O(gate188inter0));
  nand2 gate1094(.a(gate188inter0), .b(s_78), .O(gate188inter1));
  and2  gate1095(.a(G577), .b(G576), .O(gate188inter2));
  inv1  gate1096(.a(s_78), .O(gate188inter3));
  inv1  gate1097(.a(s_79), .O(gate188inter4));
  nand2 gate1098(.a(gate188inter4), .b(gate188inter3), .O(gate188inter5));
  nor2  gate1099(.a(gate188inter5), .b(gate188inter2), .O(gate188inter6));
  inv1  gate1100(.a(G576), .O(gate188inter7));
  inv1  gate1101(.a(G577), .O(gate188inter8));
  nand2 gate1102(.a(gate188inter8), .b(gate188inter7), .O(gate188inter9));
  nand2 gate1103(.a(s_79), .b(gate188inter3), .O(gate188inter10));
  nor2  gate1104(.a(gate188inter10), .b(gate188inter9), .O(gate188inter11));
  nor2  gate1105(.a(gate188inter11), .b(gate188inter6), .O(gate188inter12));
  nand2 gate1106(.a(gate188inter12), .b(gate188inter1), .O(G617));
nand2 gate189( .a(G578), .b(G579), .O(G622) );

  xor2  gate1191(.a(G581), .b(G580), .O(gate190inter0));
  nand2 gate1192(.a(gate190inter0), .b(s_92), .O(gate190inter1));
  and2  gate1193(.a(G581), .b(G580), .O(gate190inter2));
  inv1  gate1194(.a(s_92), .O(gate190inter3));
  inv1  gate1195(.a(s_93), .O(gate190inter4));
  nand2 gate1196(.a(gate190inter4), .b(gate190inter3), .O(gate190inter5));
  nor2  gate1197(.a(gate190inter5), .b(gate190inter2), .O(gate190inter6));
  inv1  gate1198(.a(G580), .O(gate190inter7));
  inv1  gate1199(.a(G581), .O(gate190inter8));
  nand2 gate1200(.a(gate190inter8), .b(gate190inter7), .O(gate190inter9));
  nand2 gate1201(.a(s_93), .b(gate190inter3), .O(gate190inter10));
  nor2  gate1202(.a(gate190inter10), .b(gate190inter9), .O(gate190inter11));
  nor2  gate1203(.a(gate190inter11), .b(gate190inter6), .O(gate190inter12));
  nand2 gate1204(.a(gate190inter12), .b(gate190inter1), .O(G627));
nand2 gate191( .a(G582), .b(G583), .O(G632) );
nand2 gate192( .a(G584), .b(G585), .O(G637) );
nand2 gate193( .a(G586), .b(G587), .O(G642) );
nand2 gate194( .a(G588), .b(G589), .O(G645) );
nand2 gate195( .a(G590), .b(G591), .O(G648) );

  xor2  gate1905(.a(G593), .b(G592), .O(gate196inter0));
  nand2 gate1906(.a(gate196inter0), .b(s_194), .O(gate196inter1));
  and2  gate1907(.a(G593), .b(G592), .O(gate196inter2));
  inv1  gate1908(.a(s_194), .O(gate196inter3));
  inv1  gate1909(.a(s_195), .O(gate196inter4));
  nand2 gate1910(.a(gate196inter4), .b(gate196inter3), .O(gate196inter5));
  nor2  gate1911(.a(gate196inter5), .b(gate196inter2), .O(gate196inter6));
  inv1  gate1912(.a(G592), .O(gate196inter7));
  inv1  gate1913(.a(G593), .O(gate196inter8));
  nand2 gate1914(.a(gate196inter8), .b(gate196inter7), .O(gate196inter9));
  nand2 gate1915(.a(s_195), .b(gate196inter3), .O(gate196inter10));
  nor2  gate1916(.a(gate196inter10), .b(gate196inter9), .O(gate196inter11));
  nor2  gate1917(.a(gate196inter11), .b(gate196inter6), .O(gate196inter12));
  nand2 gate1918(.a(gate196inter12), .b(gate196inter1), .O(G651));
nand2 gate197( .a(G594), .b(G595), .O(G654) );
nand2 gate198( .a(G596), .b(G597), .O(G657) );
nand2 gate199( .a(G598), .b(G599), .O(G660) );
nand2 gate200( .a(G600), .b(G601), .O(G663) );

  xor2  gate1471(.a(G607), .b(G602), .O(gate201inter0));
  nand2 gate1472(.a(gate201inter0), .b(s_132), .O(gate201inter1));
  and2  gate1473(.a(G607), .b(G602), .O(gate201inter2));
  inv1  gate1474(.a(s_132), .O(gate201inter3));
  inv1  gate1475(.a(s_133), .O(gate201inter4));
  nand2 gate1476(.a(gate201inter4), .b(gate201inter3), .O(gate201inter5));
  nor2  gate1477(.a(gate201inter5), .b(gate201inter2), .O(gate201inter6));
  inv1  gate1478(.a(G602), .O(gate201inter7));
  inv1  gate1479(.a(G607), .O(gate201inter8));
  nand2 gate1480(.a(gate201inter8), .b(gate201inter7), .O(gate201inter9));
  nand2 gate1481(.a(s_133), .b(gate201inter3), .O(gate201inter10));
  nor2  gate1482(.a(gate201inter10), .b(gate201inter9), .O(gate201inter11));
  nor2  gate1483(.a(gate201inter11), .b(gate201inter6), .O(gate201inter12));
  nand2 gate1484(.a(gate201inter12), .b(gate201inter1), .O(G666));
nand2 gate202( .a(G612), .b(G617), .O(G669) );

  xor2  gate1947(.a(G612), .b(G602), .O(gate203inter0));
  nand2 gate1948(.a(gate203inter0), .b(s_200), .O(gate203inter1));
  and2  gate1949(.a(G612), .b(G602), .O(gate203inter2));
  inv1  gate1950(.a(s_200), .O(gate203inter3));
  inv1  gate1951(.a(s_201), .O(gate203inter4));
  nand2 gate1952(.a(gate203inter4), .b(gate203inter3), .O(gate203inter5));
  nor2  gate1953(.a(gate203inter5), .b(gate203inter2), .O(gate203inter6));
  inv1  gate1954(.a(G602), .O(gate203inter7));
  inv1  gate1955(.a(G612), .O(gate203inter8));
  nand2 gate1956(.a(gate203inter8), .b(gate203inter7), .O(gate203inter9));
  nand2 gate1957(.a(s_201), .b(gate203inter3), .O(gate203inter10));
  nor2  gate1958(.a(gate203inter10), .b(gate203inter9), .O(gate203inter11));
  nor2  gate1959(.a(gate203inter11), .b(gate203inter6), .O(gate203inter12));
  nand2 gate1960(.a(gate203inter12), .b(gate203inter1), .O(G672));
nand2 gate204( .a(G607), .b(G617), .O(G675) );
nand2 gate205( .a(G622), .b(G627), .O(G678) );

  xor2  gate1345(.a(G637), .b(G632), .O(gate206inter0));
  nand2 gate1346(.a(gate206inter0), .b(s_114), .O(gate206inter1));
  and2  gate1347(.a(G637), .b(G632), .O(gate206inter2));
  inv1  gate1348(.a(s_114), .O(gate206inter3));
  inv1  gate1349(.a(s_115), .O(gate206inter4));
  nand2 gate1350(.a(gate206inter4), .b(gate206inter3), .O(gate206inter5));
  nor2  gate1351(.a(gate206inter5), .b(gate206inter2), .O(gate206inter6));
  inv1  gate1352(.a(G632), .O(gate206inter7));
  inv1  gate1353(.a(G637), .O(gate206inter8));
  nand2 gate1354(.a(gate206inter8), .b(gate206inter7), .O(gate206inter9));
  nand2 gate1355(.a(s_115), .b(gate206inter3), .O(gate206inter10));
  nor2  gate1356(.a(gate206inter10), .b(gate206inter9), .O(gate206inter11));
  nor2  gate1357(.a(gate206inter11), .b(gate206inter6), .O(gate206inter12));
  nand2 gate1358(.a(gate206inter12), .b(gate206inter1), .O(G681));
nand2 gate207( .a(G622), .b(G632), .O(G684) );

  xor2  gate2073(.a(G637), .b(G627), .O(gate208inter0));
  nand2 gate2074(.a(gate208inter0), .b(s_218), .O(gate208inter1));
  and2  gate2075(.a(G637), .b(G627), .O(gate208inter2));
  inv1  gate2076(.a(s_218), .O(gate208inter3));
  inv1  gate2077(.a(s_219), .O(gate208inter4));
  nand2 gate2078(.a(gate208inter4), .b(gate208inter3), .O(gate208inter5));
  nor2  gate2079(.a(gate208inter5), .b(gate208inter2), .O(gate208inter6));
  inv1  gate2080(.a(G627), .O(gate208inter7));
  inv1  gate2081(.a(G637), .O(gate208inter8));
  nand2 gate2082(.a(gate208inter8), .b(gate208inter7), .O(gate208inter9));
  nand2 gate2083(.a(s_219), .b(gate208inter3), .O(gate208inter10));
  nor2  gate2084(.a(gate208inter10), .b(gate208inter9), .O(gate208inter11));
  nor2  gate2085(.a(gate208inter11), .b(gate208inter6), .O(gate208inter12));
  nand2 gate2086(.a(gate208inter12), .b(gate208inter1), .O(G687));

  xor2  gate1891(.a(G666), .b(G602), .O(gate209inter0));
  nand2 gate1892(.a(gate209inter0), .b(s_192), .O(gate209inter1));
  and2  gate1893(.a(G666), .b(G602), .O(gate209inter2));
  inv1  gate1894(.a(s_192), .O(gate209inter3));
  inv1  gate1895(.a(s_193), .O(gate209inter4));
  nand2 gate1896(.a(gate209inter4), .b(gate209inter3), .O(gate209inter5));
  nor2  gate1897(.a(gate209inter5), .b(gate209inter2), .O(gate209inter6));
  inv1  gate1898(.a(G602), .O(gate209inter7));
  inv1  gate1899(.a(G666), .O(gate209inter8));
  nand2 gate1900(.a(gate209inter8), .b(gate209inter7), .O(gate209inter9));
  nand2 gate1901(.a(s_193), .b(gate209inter3), .O(gate209inter10));
  nor2  gate1902(.a(gate209inter10), .b(gate209inter9), .O(gate209inter11));
  nor2  gate1903(.a(gate209inter11), .b(gate209inter6), .O(gate209inter12));
  nand2 gate1904(.a(gate209inter12), .b(gate209inter1), .O(G690));

  xor2  gate1877(.a(G666), .b(G607), .O(gate210inter0));
  nand2 gate1878(.a(gate210inter0), .b(s_190), .O(gate210inter1));
  and2  gate1879(.a(G666), .b(G607), .O(gate210inter2));
  inv1  gate1880(.a(s_190), .O(gate210inter3));
  inv1  gate1881(.a(s_191), .O(gate210inter4));
  nand2 gate1882(.a(gate210inter4), .b(gate210inter3), .O(gate210inter5));
  nor2  gate1883(.a(gate210inter5), .b(gate210inter2), .O(gate210inter6));
  inv1  gate1884(.a(G607), .O(gate210inter7));
  inv1  gate1885(.a(G666), .O(gate210inter8));
  nand2 gate1886(.a(gate210inter8), .b(gate210inter7), .O(gate210inter9));
  nand2 gate1887(.a(s_191), .b(gate210inter3), .O(gate210inter10));
  nor2  gate1888(.a(gate210inter10), .b(gate210inter9), .O(gate210inter11));
  nor2  gate1889(.a(gate210inter11), .b(gate210inter6), .O(gate210inter12));
  nand2 gate1890(.a(gate210inter12), .b(gate210inter1), .O(G691));

  xor2  gate1527(.a(G669), .b(G612), .O(gate211inter0));
  nand2 gate1528(.a(gate211inter0), .b(s_140), .O(gate211inter1));
  and2  gate1529(.a(G669), .b(G612), .O(gate211inter2));
  inv1  gate1530(.a(s_140), .O(gate211inter3));
  inv1  gate1531(.a(s_141), .O(gate211inter4));
  nand2 gate1532(.a(gate211inter4), .b(gate211inter3), .O(gate211inter5));
  nor2  gate1533(.a(gate211inter5), .b(gate211inter2), .O(gate211inter6));
  inv1  gate1534(.a(G612), .O(gate211inter7));
  inv1  gate1535(.a(G669), .O(gate211inter8));
  nand2 gate1536(.a(gate211inter8), .b(gate211inter7), .O(gate211inter9));
  nand2 gate1537(.a(s_141), .b(gate211inter3), .O(gate211inter10));
  nor2  gate1538(.a(gate211inter10), .b(gate211inter9), .O(gate211inter11));
  nor2  gate1539(.a(gate211inter11), .b(gate211inter6), .O(gate211inter12));
  nand2 gate1540(.a(gate211inter12), .b(gate211inter1), .O(G692));

  xor2  gate2003(.a(G669), .b(G617), .O(gate212inter0));
  nand2 gate2004(.a(gate212inter0), .b(s_208), .O(gate212inter1));
  and2  gate2005(.a(G669), .b(G617), .O(gate212inter2));
  inv1  gate2006(.a(s_208), .O(gate212inter3));
  inv1  gate2007(.a(s_209), .O(gate212inter4));
  nand2 gate2008(.a(gate212inter4), .b(gate212inter3), .O(gate212inter5));
  nor2  gate2009(.a(gate212inter5), .b(gate212inter2), .O(gate212inter6));
  inv1  gate2010(.a(G617), .O(gate212inter7));
  inv1  gate2011(.a(G669), .O(gate212inter8));
  nand2 gate2012(.a(gate212inter8), .b(gate212inter7), .O(gate212inter9));
  nand2 gate2013(.a(s_209), .b(gate212inter3), .O(gate212inter10));
  nor2  gate2014(.a(gate212inter10), .b(gate212inter9), .O(gate212inter11));
  nor2  gate2015(.a(gate212inter11), .b(gate212inter6), .O(gate212inter12));
  nand2 gate2016(.a(gate212inter12), .b(gate212inter1), .O(G693));
nand2 gate213( .a(G602), .b(G672), .O(G694) );

  xor2  gate1793(.a(G672), .b(G612), .O(gate214inter0));
  nand2 gate1794(.a(gate214inter0), .b(s_178), .O(gate214inter1));
  and2  gate1795(.a(G672), .b(G612), .O(gate214inter2));
  inv1  gate1796(.a(s_178), .O(gate214inter3));
  inv1  gate1797(.a(s_179), .O(gate214inter4));
  nand2 gate1798(.a(gate214inter4), .b(gate214inter3), .O(gate214inter5));
  nor2  gate1799(.a(gate214inter5), .b(gate214inter2), .O(gate214inter6));
  inv1  gate1800(.a(G612), .O(gate214inter7));
  inv1  gate1801(.a(G672), .O(gate214inter8));
  nand2 gate1802(.a(gate214inter8), .b(gate214inter7), .O(gate214inter9));
  nand2 gate1803(.a(s_179), .b(gate214inter3), .O(gate214inter10));
  nor2  gate1804(.a(gate214inter10), .b(gate214inter9), .O(gate214inter11));
  nor2  gate1805(.a(gate214inter11), .b(gate214inter6), .O(gate214inter12));
  nand2 gate1806(.a(gate214inter12), .b(gate214inter1), .O(G695));
nand2 gate215( .a(G607), .b(G675), .O(G696) );
nand2 gate216( .a(G617), .b(G675), .O(G697) );

  xor2  gate2591(.a(G678), .b(G622), .O(gate217inter0));
  nand2 gate2592(.a(gate217inter0), .b(s_292), .O(gate217inter1));
  and2  gate2593(.a(G678), .b(G622), .O(gate217inter2));
  inv1  gate2594(.a(s_292), .O(gate217inter3));
  inv1  gate2595(.a(s_293), .O(gate217inter4));
  nand2 gate2596(.a(gate217inter4), .b(gate217inter3), .O(gate217inter5));
  nor2  gate2597(.a(gate217inter5), .b(gate217inter2), .O(gate217inter6));
  inv1  gate2598(.a(G622), .O(gate217inter7));
  inv1  gate2599(.a(G678), .O(gate217inter8));
  nand2 gate2600(.a(gate217inter8), .b(gate217inter7), .O(gate217inter9));
  nand2 gate2601(.a(s_293), .b(gate217inter3), .O(gate217inter10));
  nor2  gate2602(.a(gate217inter10), .b(gate217inter9), .O(gate217inter11));
  nor2  gate2603(.a(gate217inter11), .b(gate217inter6), .O(gate217inter12));
  nand2 gate2604(.a(gate217inter12), .b(gate217inter1), .O(G698));

  xor2  gate1667(.a(G678), .b(G627), .O(gate218inter0));
  nand2 gate1668(.a(gate218inter0), .b(s_160), .O(gate218inter1));
  and2  gate1669(.a(G678), .b(G627), .O(gate218inter2));
  inv1  gate1670(.a(s_160), .O(gate218inter3));
  inv1  gate1671(.a(s_161), .O(gate218inter4));
  nand2 gate1672(.a(gate218inter4), .b(gate218inter3), .O(gate218inter5));
  nor2  gate1673(.a(gate218inter5), .b(gate218inter2), .O(gate218inter6));
  inv1  gate1674(.a(G627), .O(gate218inter7));
  inv1  gate1675(.a(G678), .O(gate218inter8));
  nand2 gate1676(.a(gate218inter8), .b(gate218inter7), .O(gate218inter9));
  nand2 gate1677(.a(s_161), .b(gate218inter3), .O(gate218inter10));
  nor2  gate1678(.a(gate218inter10), .b(gate218inter9), .O(gate218inter11));
  nor2  gate1679(.a(gate218inter11), .b(gate218inter6), .O(gate218inter12));
  nand2 gate1680(.a(gate218inter12), .b(gate218inter1), .O(G699));
nand2 gate219( .a(G632), .b(G681), .O(G700) );

  xor2  gate2241(.a(G681), .b(G637), .O(gate220inter0));
  nand2 gate2242(.a(gate220inter0), .b(s_242), .O(gate220inter1));
  and2  gate2243(.a(G681), .b(G637), .O(gate220inter2));
  inv1  gate2244(.a(s_242), .O(gate220inter3));
  inv1  gate2245(.a(s_243), .O(gate220inter4));
  nand2 gate2246(.a(gate220inter4), .b(gate220inter3), .O(gate220inter5));
  nor2  gate2247(.a(gate220inter5), .b(gate220inter2), .O(gate220inter6));
  inv1  gate2248(.a(G637), .O(gate220inter7));
  inv1  gate2249(.a(G681), .O(gate220inter8));
  nand2 gate2250(.a(gate220inter8), .b(gate220inter7), .O(gate220inter9));
  nand2 gate2251(.a(s_243), .b(gate220inter3), .O(gate220inter10));
  nor2  gate2252(.a(gate220inter10), .b(gate220inter9), .O(gate220inter11));
  nor2  gate2253(.a(gate220inter11), .b(gate220inter6), .O(gate220inter12));
  nand2 gate2254(.a(gate220inter12), .b(gate220inter1), .O(G701));
nand2 gate221( .a(G622), .b(G684), .O(G702) );

  xor2  gate1807(.a(G684), .b(G632), .O(gate222inter0));
  nand2 gate1808(.a(gate222inter0), .b(s_180), .O(gate222inter1));
  and2  gate1809(.a(G684), .b(G632), .O(gate222inter2));
  inv1  gate1810(.a(s_180), .O(gate222inter3));
  inv1  gate1811(.a(s_181), .O(gate222inter4));
  nand2 gate1812(.a(gate222inter4), .b(gate222inter3), .O(gate222inter5));
  nor2  gate1813(.a(gate222inter5), .b(gate222inter2), .O(gate222inter6));
  inv1  gate1814(.a(G632), .O(gate222inter7));
  inv1  gate1815(.a(G684), .O(gate222inter8));
  nand2 gate1816(.a(gate222inter8), .b(gate222inter7), .O(gate222inter9));
  nand2 gate1817(.a(s_181), .b(gate222inter3), .O(gate222inter10));
  nor2  gate1818(.a(gate222inter10), .b(gate222inter9), .O(gate222inter11));
  nor2  gate1819(.a(gate222inter11), .b(gate222inter6), .O(gate222inter12));
  nand2 gate1820(.a(gate222inter12), .b(gate222inter1), .O(G703));

  xor2  gate1681(.a(G687), .b(G627), .O(gate223inter0));
  nand2 gate1682(.a(gate223inter0), .b(s_162), .O(gate223inter1));
  and2  gate1683(.a(G687), .b(G627), .O(gate223inter2));
  inv1  gate1684(.a(s_162), .O(gate223inter3));
  inv1  gate1685(.a(s_163), .O(gate223inter4));
  nand2 gate1686(.a(gate223inter4), .b(gate223inter3), .O(gate223inter5));
  nor2  gate1687(.a(gate223inter5), .b(gate223inter2), .O(gate223inter6));
  inv1  gate1688(.a(G627), .O(gate223inter7));
  inv1  gate1689(.a(G687), .O(gate223inter8));
  nand2 gate1690(.a(gate223inter8), .b(gate223inter7), .O(gate223inter9));
  nand2 gate1691(.a(s_163), .b(gate223inter3), .O(gate223inter10));
  nor2  gate1692(.a(gate223inter10), .b(gate223inter9), .O(gate223inter11));
  nor2  gate1693(.a(gate223inter11), .b(gate223inter6), .O(gate223inter12));
  nand2 gate1694(.a(gate223inter12), .b(gate223inter1), .O(G704));
nand2 gate224( .a(G637), .b(G687), .O(G705) );

  xor2  gate1177(.a(G691), .b(G690), .O(gate225inter0));
  nand2 gate1178(.a(gate225inter0), .b(s_90), .O(gate225inter1));
  and2  gate1179(.a(G691), .b(G690), .O(gate225inter2));
  inv1  gate1180(.a(s_90), .O(gate225inter3));
  inv1  gate1181(.a(s_91), .O(gate225inter4));
  nand2 gate1182(.a(gate225inter4), .b(gate225inter3), .O(gate225inter5));
  nor2  gate1183(.a(gate225inter5), .b(gate225inter2), .O(gate225inter6));
  inv1  gate1184(.a(G690), .O(gate225inter7));
  inv1  gate1185(.a(G691), .O(gate225inter8));
  nand2 gate1186(.a(gate225inter8), .b(gate225inter7), .O(gate225inter9));
  nand2 gate1187(.a(s_91), .b(gate225inter3), .O(gate225inter10));
  nor2  gate1188(.a(gate225inter10), .b(gate225inter9), .O(gate225inter11));
  nor2  gate1189(.a(gate225inter11), .b(gate225inter6), .O(gate225inter12));
  nand2 gate1190(.a(gate225inter12), .b(gate225inter1), .O(G706));

  xor2  gate687(.a(G693), .b(G692), .O(gate226inter0));
  nand2 gate688(.a(gate226inter0), .b(s_20), .O(gate226inter1));
  and2  gate689(.a(G693), .b(G692), .O(gate226inter2));
  inv1  gate690(.a(s_20), .O(gate226inter3));
  inv1  gate691(.a(s_21), .O(gate226inter4));
  nand2 gate692(.a(gate226inter4), .b(gate226inter3), .O(gate226inter5));
  nor2  gate693(.a(gate226inter5), .b(gate226inter2), .O(gate226inter6));
  inv1  gate694(.a(G692), .O(gate226inter7));
  inv1  gate695(.a(G693), .O(gate226inter8));
  nand2 gate696(.a(gate226inter8), .b(gate226inter7), .O(gate226inter9));
  nand2 gate697(.a(s_21), .b(gate226inter3), .O(gate226inter10));
  nor2  gate698(.a(gate226inter10), .b(gate226inter9), .O(gate226inter11));
  nor2  gate699(.a(gate226inter11), .b(gate226inter6), .O(gate226inter12));
  nand2 gate700(.a(gate226inter12), .b(gate226inter1), .O(G709));

  xor2  gate1555(.a(G695), .b(G694), .O(gate227inter0));
  nand2 gate1556(.a(gate227inter0), .b(s_144), .O(gate227inter1));
  and2  gate1557(.a(G695), .b(G694), .O(gate227inter2));
  inv1  gate1558(.a(s_144), .O(gate227inter3));
  inv1  gate1559(.a(s_145), .O(gate227inter4));
  nand2 gate1560(.a(gate227inter4), .b(gate227inter3), .O(gate227inter5));
  nor2  gate1561(.a(gate227inter5), .b(gate227inter2), .O(gate227inter6));
  inv1  gate1562(.a(G694), .O(gate227inter7));
  inv1  gate1563(.a(G695), .O(gate227inter8));
  nand2 gate1564(.a(gate227inter8), .b(gate227inter7), .O(gate227inter9));
  nand2 gate1565(.a(s_145), .b(gate227inter3), .O(gate227inter10));
  nor2  gate1566(.a(gate227inter10), .b(gate227inter9), .O(gate227inter11));
  nor2  gate1567(.a(gate227inter11), .b(gate227inter6), .O(gate227inter12));
  nand2 gate1568(.a(gate227inter12), .b(gate227inter1), .O(G712));

  xor2  gate841(.a(G697), .b(G696), .O(gate228inter0));
  nand2 gate842(.a(gate228inter0), .b(s_42), .O(gate228inter1));
  and2  gate843(.a(G697), .b(G696), .O(gate228inter2));
  inv1  gate844(.a(s_42), .O(gate228inter3));
  inv1  gate845(.a(s_43), .O(gate228inter4));
  nand2 gate846(.a(gate228inter4), .b(gate228inter3), .O(gate228inter5));
  nor2  gate847(.a(gate228inter5), .b(gate228inter2), .O(gate228inter6));
  inv1  gate848(.a(G696), .O(gate228inter7));
  inv1  gate849(.a(G697), .O(gate228inter8));
  nand2 gate850(.a(gate228inter8), .b(gate228inter7), .O(gate228inter9));
  nand2 gate851(.a(s_43), .b(gate228inter3), .O(gate228inter10));
  nor2  gate852(.a(gate228inter10), .b(gate228inter9), .O(gate228inter11));
  nor2  gate853(.a(gate228inter11), .b(gate228inter6), .O(gate228inter12));
  nand2 gate854(.a(gate228inter12), .b(gate228inter1), .O(G715));
nand2 gate229( .a(G698), .b(G699), .O(G718) );
nand2 gate230( .a(G700), .b(G701), .O(G721) );
nand2 gate231( .a(G702), .b(G703), .O(G724) );

  xor2  gate2339(.a(G705), .b(G704), .O(gate232inter0));
  nand2 gate2340(.a(gate232inter0), .b(s_256), .O(gate232inter1));
  and2  gate2341(.a(G705), .b(G704), .O(gate232inter2));
  inv1  gate2342(.a(s_256), .O(gate232inter3));
  inv1  gate2343(.a(s_257), .O(gate232inter4));
  nand2 gate2344(.a(gate232inter4), .b(gate232inter3), .O(gate232inter5));
  nor2  gate2345(.a(gate232inter5), .b(gate232inter2), .O(gate232inter6));
  inv1  gate2346(.a(G704), .O(gate232inter7));
  inv1  gate2347(.a(G705), .O(gate232inter8));
  nand2 gate2348(.a(gate232inter8), .b(gate232inter7), .O(gate232inter9));
  nand2 gate2349(.a(s_257), .b(gate232inter3), .O(gate232inter10));
  nor2  gate2350(.a(gate232inter10), .b(gate232inter9), .O(gate232inter11));
  nor2  gate2351(.a(gate232inter11), .b(gate232inter6), .O(gate232inter12));
  nand2 gate2352(.a(gate232inter12), .b(gate232inter1), .O(G727));

  xor2  gate1919(.a(G718), .b(G242), .O(gate233inter0));
  nand2 gate1920(.a(gate233inter0), .b(s_196), .O(gate233inter1));
  and2  gate1921(.a(G718), .b(G242), .O(gate233inter2));
  inv1  gate1922(.a(s_196), .O(gate233inter3));
  inv1  gate1923(.a(s_197), .O(gate233inter4));
  nand2 gate1924(.a(gate233inter4), .b(gate233inter3), .O(gate233inter5));
  nor2  gate1925(.a(gate233inter5), .b(gate233inter2), .O(gate233inter6));
  inv1  gate1926(.a(G242), .O(gate233inter7));
  inv1  gate1927(.a(G718), .O(gate233inter8));
  nand2 gate1928(.a(gate233inter8), .b(gate233inter7), .O(gate233inter9));
  nand2 gate1929(.a(s_197), .b(gate233inter3), .O(gate233inter10));
  nor2  gate1930(.a(gate233inter10), .b(gate233inter9), .O(gate233inter11));
  nor2  gate1931(.a(gate233inter11), .b(gate233inter6), .O(gate233inter12));
  nand2 gate1932(.a(gate233inter12), .b(gate233inter1), .O(G730));
nand2 gate234( .a(G245), .b(G721), .O(G733) );

  xor2  gate1331(.a(G724), .b(G248), .O(gate235inter0));
  nand2 gate1332(.a(gate235inter0), .b(s_112), .O(gate235inter1));
  and2  gate1333(.a(G724), .b(G248), .O(gate235inter2));
  inv1  gate1334(.a(s_112), .O(gate235inter3));
  inv1  gate1335(.a(s_113), .O(gate235inter4));
  nand2 gate1336(.a(gate235inter4), .b(gate235inter3), .O(gate235inter5));
  nor2  gate1337(.a(gate235inter5), .b(gate235inter2), .O(gate235inter6));
  inv1  gate1338(.a(G248), .O(gate235inter7));
  inv1  gate1339(.a(G724), .O(gate235inter8));
  nand2 gate1340(.a(gate235inter8), .b(gate235inter7), .O(gate235inter9));
  nand2 gate1341(.a(s_113), .b(gate235inter3), .O(gate235inter10));
  nor2  gate1342(.a(gate235inter10), .b(gate235inter9), .O(gate235inter11));
  nor2  gate1343(.a(gate235inter11), .b(gate235inter6), .O(gate235inter12));
  nand2 gate1344(.a(gate235inter12), .b(gate235inter1), .O(G736));
nand2 gate236( .a(G251), .b(G727), .O(G739) );

  xor2  gate1639(.a(G706), .b(G254), .O(gate237inter0));
  nand2 gate1640(.a(gate237inter0), .b(s_156), .O(gate237inter1));
  and2  gate1641(.a(G706), .b(G254), .O(gate237inter2));
  inv1  gate1642(.a(s_156), .O(gate237inter3));
  inv1  gate1643(.a(s_157), .O(gate237inter4));
  nand2 gate1644(.a(gate237inter4), .b(gate237inter3), .O(gate237inter5));
  nor2  gate1645(.a(gate237inter5), .b(gate237inter2), .O(gate237inter6));
  inv1  gate1646(.a(G254), .O(gate237inter7));
  inv1  gate1647(.a(G706), .O(gate237inter8));
  nand2 gate1648(.a(gate237inter8), .b(gate237inter7), .O(gate237inter9));
  nand2 gate1649(.a(s_157), .b(gate237inter3), .O(gate237inter10));
  nor2  gate1650(.a(gate237inter10), .b(gate237inter9), .O(gate237inter11));
  nor2  gate1651(.a(gate237inter11), .b(gate237inter6), .O(gate237inter12));
  nand2 gate1652(.a(gate237inter12), .b(gate237inter1), .O(G742));
nand2 gate238( .a(G257), .b(G709), .O(G745) );

  xor2  gate743(.a(G712), .b(G260), .O(gate239inter0));
  nand2 gate744(.a(gate239inter0), .b(s_28), .O(gate239inter1));
  and2  gate745(.a(G712), .b(G260), .O(gate239inter2));
  inv1  gate746(.a(s_28), .O(gate239inter3));
  inv1  gate747(.a(s_29), .O(gate239inter4));
  nand2 gate748(.a(gate239inter4), .b(gate239inter3), .O(gate239inter5));
  nor2  gate749(.a(gate239inter5), .b(gate239inter2), .O(gate239inter6));
  inv1  gate750(.a(G260), .O(gate239inter7));
  inv1  gate751(.a(G712), .O(gate239inter8));
  nand2 gate752(.a(gate239inter8), .b(gate239inter7), .O(gate239inter9));
  nand2 gate753(.a(s_29), .b(gate239inter3), .O(gate239inter10));
  nor2  gate754(.a(gate239inter10), .b(gate239inter9), .O(gate239inter11));
  nor2  gate755(.a(gate239inter11), .b(gate239inter6), .O(gate239inter12));
  nand2 gate756(.a(gate239inter12), .b(gate239inter1), .O(G748));
nand2 gate240( .a(G263), .b(G715), .O(G751) );

  xor2  gate2437(.a(G730), .b(G242), .O(gate241inter0));
  nand2 gate2438(.a(gate241inter0), .b(s_270), .O(gate241inter1));
  and2  gate2439(.a(G730), .b(G242), .O(gate241inter2));
  inv1  gate2440(.a(s_270), .O(gate241inter3));
  inv1  gate2441(.a(s_271), .O(gate241inter4));
  nand2 gate2442(.a(gate241inter4), .b(gate241inter3), .O(gate241inter5));
  nor2  gate2443(.a(gate241inter5), .b(gate241inter2), .O(gate241inter6));
  inv1  gate2444(.a(G242), .O(gate241inter7));
  inv1  gate2445(.a(G730), .O(gate241inter8));
  nand2 gate2446(.a(gate241inter8), .b(gate241inter7), .O(gate241inter9));
  nand2 gate2447(.a(s_271), .b(gate241inter3), .O(gate241inter10));
  nor2  gate2448(.a(gate241inter10), .b(gate241inter9), .O(gate241inter11));
  nor2  gate2449(.a(gate241inter11), .b(gate241inter6), .O(gate241inter12));
  nand2 gate2450(.a(gate241inter12), .b(gate241inter1), .O(G754));

  xor2  gate2101(.a(G730), .b(G718), .O(gate242inter0));
  nand2 gate2102(.a(gate242inter0), .b(s_222), .O(gate242inter1));
  and2  gate2103(.a(G730), .b(G718), .O(gate242inter2));
  inv1  gate2104(.a(s_222), .O(gate242inter3));
  inv1  gate2105(.a(s_223), .O(gate242inter4));
  nand2 gate2106(.a(gate242inter4), .b(gate242inter3), .O(gate242inter5));
  nor2  gate2107(.a(gate242inter5), .b(gate242inter2), .O(gate242inter6));
  inv1  gate2108(.a(G718), .O(gate242inter7));
  inv1  gate2109(.a(G730), .O(gate242inter8));
  nand2 gate2110(.a(gate242inter8), .b(gate242inter7), .O(gate242inter9));
  nand2 gate2111(.a(s_223), .b(gate242inter3), .O(gate242inter10));
  nor2  gate2112(.a(gate242inter10), .b(gate242inter9), .O(gate242inter11));
  nor2  gate2113(.a(gate242inter11), .b(gate242inter6), .O(gate242inter12));
  nand2 gate2114(.a(gate242inter12), .b(gate242inter1), .O(G755));
nand2 gate243( .a(G245), .b(G733), .O(G756) );
nand2 gate244( .a(G721), .b(G733), .O(G757) );

  xor2  gate1457(.a(G736), .b(G248), .O(gate245inter0));
  nand2 gate1458(.a(gate245inter0), .b(s_130), .O(gate245inter1));
  and2  gate1459(.a(G736), .b(G248), .O(gate245inter2));
  inv1  gate1460(.a(s_130), .O(gate245inter3));
  inv1  gate1461(.a(s_131), .O(gate245inter4));
  nand2 gate1462(.a(gate245inter4), .b(gate245inter3), .O(gate245inter5));
  nor2  gate1463(.a(gate245inter5), .b(gate245inter2), .O(gate245inter6));
  inv1  gate1464(.a(G248), .O(gate245inter7));
  inv1  gate1465(.a(G736), .O(gate245inter8));
  nand2 gate1466(.a(gate245inter8), .b(gate245inter7), .O(gate245inter9));
  nand2 gate1467(.a(s_131), .b(gate245inter3), .O(gate245inter10));
  nor2  gate1468(.a(gate245inter10), .b(gate245inter9), .O(gate245inter11));
  nor2  gate1469(.a(gate245inter11), .b(gate245inter6), .O(gate245inter12));
  nand2 gate1470(.a(gate245inter12), .b(gate245inter1), .O(G758));
nand2 gate246( .a(G724), .b(G736), .O(G759) );
nand2 gate247( .a(G251), .b(G739), .O(G760) );
nand2 gate248( .a(G727), .b(G739), .O(G761) );

  xor2  gate2717(.a(G742), .b(G254), .O(gate249inter0));
  nand2 gate2718(.a(gate249inter0), .b(s_310), .O(gate249inter1));
  and2  gate2719(.a(G742), .b(G254), .O(gate249inter2));
  inv1  gate2720(.a(s_310), .O(gate249inter3));
  inv1  gate2721(.a(s_311), .O(gate249inter4));
  nand2 gate2722(.a(gate249inter4), .b(gate249inter3), .O(gate249inter5));
  nor2  gate2723(.a(gate249inter5), .b(gate249inter2), .O(gate249inter6));
  inv1  gate2724(.a(G254), .O(gate249inter7));
  inv1  gate2725(.a(G742), .O(gate249inter8));
  nand2 gate2726(.a(gate249inter8), .b(gate249inter7), .O(gate249inter9));
  nand2 gate2727(.a(s_311), .b(gate249inter3), .O(gate249inter10));
  nor2  gate2728(.a(gate249inter10), .b(gate249inter9), .O(gate249inter11));
  nor2  gate2729(.a(gate249inter11), .b(gate249inter6), .O(gate249inter12));
  nand2 gate2730(.a(gate249inter12), .b(gate249inter1), .O(G762));

  xor2  gate2703(.a(G742), .b(G706), .O(gate250inter0));
  nand2 gate2704(.a(gate250inter0), .b(s_308), .O(gate250inter1));
  and2  gate2705(.a(G742), .b(G706), .O(gate250inter2));
  inv1  gate2706(.a(s_308), .O(gate250inter3));
  inv1  gate2707(.a(s_309), .O(gate250inter4));
  nand2 gate2708(.a(gate250inter4), .b(gate250inter3), .O(gate250inter5));
  nor2  gate2709(.a(gate250inter5), .b(gate250inter2), .O(gate250inter6));
  inv1  gate2710(.a(G706), .O(gate250inter7));
  inv1  gate2711(.a(G742), .O(gate250inter8));
  nand2 gate2712(.a(gate250inter8), .b(gate250inter7), .O(gate250inter9));
  nand2 gate2713(.a(s_309), .b(gate250inter3), .O(gate250inter10));
  nor2  gate2714(.a(gate250inter10), .b(gate250inter9), .O(gate250inter11));
  nor2  gate2715(.a(gate250inter11), .b(gate250inter6), .O(gate250inter12));
  nand2 gate2716(.a(gate250inter12), .b(gate250inter1), .O(G763));
nand2 gate251( .a(G257), .b(G745), .O(G764) );
nand2 gate252( .a(G709), .b(G745), .O(G765) );

  xor2  gate2549(.a(G748), .b(G260), .O(gate253inter0));
  nand2 gate2550(.a(gate253inter0), .b(s_286), .O(gate253inter1));
  and2  gate2551(.a(G748), .b(G260), .O(gate253inter2));
  inv1  gate2552(.a(s_286), .O(gate253inter3));
  inv1  gate2553(.a(s_287), .O(gate253inter4));
  nand2 gate2554(.a(gate253inter4), .b(gate253inter3), .O(gate253inter5));
  nor2  gate2555(.a(gate253inter5), .b(gate253inter2), .O(gate253inter6));
  inv1  gate2556(.a(G260), .O(gate253inter7));
  inv1  gate2557(.a(G748), .O(gate253inter8));
  nand2 gate2558(.a(gate253inter8), .b(gate253inter7), .O(gate253inter9));
  nand2 gate2559(.a(s_287), .b(gate253inter3), .O(gate253inter10));
  nor2  gate2560(.a(gate253inter10), .b(gate253inter9), .O(gate253inter11));
  nor2  gate2561(.a(gate253inter11), .b(gate253inter6), .O(gate253inter12));
  nand2 gate2562(.a(gate253inter12), .b(gate253inter1), .O(G766));

  xor2  gate1933(.a(G748), .b(G712), .O(gate254inter0));
  nand2 gate1934(.a(gate254inter0), .b(s_198), .O(gate254inter1));
  and2  gate1935(.a(G748), .b(G712), .O(gate254inter2));
  inv1  gate1936(.a(s_198), .O(gate254inter3));
  inv1  gate1937(.a(s_199), .O(gate254inter4));
  nand2 gate1938(.a(gate254inter4), .b(gate254inter3), .O(gate254inter5));
  nor2  gate1939(.a(gate254inter5), .b(gate254inter2), .O(gate254inter6));
  inv1  gate1940(.a(G712), .O(gate254inter7));
  inv1  gate1941(.a(G748), .O(gate254inter8));
  nand2 gate1942(.a(gate254inter8), .b(gate254inter7), .O(gate254inter9));
  nand2 gate1943(.a(s_199), .b(gate254inter3), .O(gate254inter10));
  nor2  gate1944(.a(gate254inter10), .b(gate254inter9), .O(gate254inter11));
  nor2  gate1945(.a(gate254inter11), .b(gate254inter6), .O(gate254inter12));
  nand2 gate1946(.a(gate254inter12), .b(gate254inter1), .O(G767));

  xor2  gate883(.a(G751), .b(G263), .O(gate255inter0));
  nand2 gate884(.a(gate255inter0), .b(s_48), .O(gate255inter1));
  and2  gate885(.a(G751), .b(G263), .O(gate255inter2));
  inv1  gate886(.a(s_48), .O(gate255inter3));
  inv1  gate887(.a(s_49), .O(gate255inter4));
  nand2 gate888(.a(gate255inter4), .b(gate255inter3), .O(gate255inter5));
  nor2  gate889(.a(gate255inter5), .b(gate255inter2), .O(gate255inter6));
  inv1  gate890(.a(G263), .O(gate255inter7));
  inv1  gate891(.a(G751), .O(gate255inter8));
  nand2 gate892(.a(gate255inter8), .b(gate255inter7), .O(gate255inter9));
  nand2 gate893(.a(s_49), .b(gate255inter3), .O(gate255inter10));
  nor2  gate894(.a(gate255inter10), .b(gate255inter9), .O(gate255inter11));
  nor2  gate895(.a(gate255inter11), .b(gate255inter6), .O(gate255inter12));
  nand2 gate896(.a(gate255inter12), .b(gate255inter1), .O(G768));

  xor2  gate2535(.a(G751), .b(G715), .O(gate256inter0));
  nand2 gate2536(.a(gate256inter0), .b(s_284), .O(gate256inter1));
  and2  gate2537(.a(G751), .b(G715), .O(gate256inter2));
  inv1  gate2538(.a(s_284), .O(gate256inter3));
  inv1  gate2539(.a(s_285), .O(gate256inter4));
  nand2 gate2540(.a(gate256inter4), .b(gate256inter3), .O(gate256inter5));
  nor2  gate2541(.a(gate256inter5), .b(gate256inter2), .O(gate256inter6));
  inv1  gate2542(.a(G715), .O(gate256inter7));
  inv1  gate2543(.a(G751), .O(gate256inter8));
  nand2 gate2544(.a(gate256inter8), .b(gate256inter7), .O(gate256inter9));
  nand2 gate2545(.a(s_285), .b(gate256inter3), .O(gate256inter10));
  nor2  gate2546(.a(gate256inter10), .b(gate256inter9), .O(gate256inter11));
  nor2  gate2547(.a(gate256inter11), .b(gate256inter6), .O(gate256inter12));
  nand2 gate2548(.a(gate256inter12), .b(gate256inter1), .O(G769));

  xor2  gate2283(.a(G755), .b(G754), .O(gate257inter0));
  nand2 gate2284(.a(gate257inter0), .b(s_248), .O(gate257inter1));
  and2  gate2285(.a(G755), .b(G754), .O(gate257inter2));
  inv1  gate2286(.a(s_248), .O(gate257inter3));
  inv1  gate2287(.a(s_249), .O(gate257inter4));
  nand2 gate2288(.a(gate257inter4), .b(gate257inter3), .O(gate257inter5));
  nor2  gate2289(.a(gate257inter5), .b(gate257inter2), .O(gate257inter6));
  inv1  gate2290(.a(G754), .O(gate257inter7));
  inv1  gate2291(.a(G755), .O(gate257inter8));
  nand2 gate2292(.a(gate257inter8), .b(gate257inter7), .O(gate257inter9));
  nand2 gate2293(.a(s_249), .b(gate257inter3), .O(gate257inter10));
  nor2  gate2294(.a(gate257inter10), .b(gate257inter9), .O(gate257inter11));
  nor2  gate2295(.a(gate257inter11), .b(gate257inter6), .O(gate257inter12));
  nand2 gate2296(.a(gate257inter12), .b(gate257inter1), .O(G770));
nand2 gate258( .a(G756), .b(G757), .O(G773) );
nand2 gate259( .a(G758), .b(G759), .O(G776) );

  xor2  gate2563(.a(G761), .b(G760), .O(gate260inter0));
  nand2 gate2564(.a(gate260inter0), .b(s_288), .O(gate260inter1));
  and2  gate2565(.a(G761), .b(G760), .O(gate260inter2));
  inv1  gate2566(.a(s_288), .O(gate260inter3));
  inv1  gate2567(.a(s_289), .O(gate260inter4));
  nand2 gate2568(.a(gate260inter4), .b(gate260inter3), .O(gate260inter5));
  nor2  gate2569(.a(gate260inter5), .b(gate260inter2), .O(gate260inter6));
  inv1  gate2570(.a(G760), .O(gate260inter7));
  inv1  gate2571(.a(G761), .O(gate260inter8));
  nand2 gate2572(.a(gate260inter8), .b(gate260inter7), .O(gate260inter9));
  nand2 gate2573(.a(s_289), .b(gate260inter3), .O(gate260inter10));
  nor2  gate2574(.a(gate260inter10), .b(gate260inter9), .O(gate260inter11));
  nor2  gate2575(.a(gate260inter11), .b(gate260inter6), .O(gate260inter12));
  nand2 gate2576(.a(gate260inter12), .b(gate260inter1), .O(G779));

  xor2  gate1653(.a(G763), .b(G762), .O(gate261inter0));
  nand2 gate1654(.a(gate261inter0), .b(s_158), .O(gate261inter1));
  and2  gate1655(.a(G763), .b(G762), .O(gate261inter2));
  inv1  gate1656(.a(s_158), .O(gate261inter3));
  inv1  gate1657(.a(s_159), .O(gate261inter4));
  nand2 gate1658(.a(gate261inter4), .b(gate261inter3), .O(gate261inter5));
  nor2  gate1659(.a(gate261inter5), .b(gate261inter2), .O(gate261inter6));
  inv1  gate1660(.a(G762), .O(gate261inter7));
  inv1  gate1661(.a(G763), .O(gate261inter8));
  nand2 gate1662(.a(gate261inter8), .b(gate261inter7), .O(gate261inter9));
  nand2 gate1663(.a(s_159), .b(gate261inter3), .O(gate261inter10));
  nor2  gate1664(.a(gate261inter10), .b(gate261inter9), .O(gate261inter11));
  nor2  gate1665(.a(gate261inter11), .b(gate261inter6), .O(gate261inter12));
  nand2 gate1666(.a(gate261inter12), .b(gate261inter1), .O(G782));

  xor2  gate2059(.a(G765), .b(G764), .O(gate262inter0));
  nand2 gate2060(.a(gate262inter0), .b(s_216), .O(gate262inter1));
  and2  gate2061(.a(G765), .b(G764), .O(gate262inter2));
  inv1  gate2062(.a(s_216), .O(gate262inter3));
  inv1  gate2063(.a(s_217), .O(gate262inter4));
  nand2 gate2064(.a(gate262inter4), .b(gate262inter3), .O(gate262inter5));
  nor2  gate2065(.a(gate262inter5), .b(gate262inter2), .O(gate262inter6));
  inv1  gate2066(.a(G764), .O(gate262inter7));
  inv1  gate2067(.a(G765), .O(gate262inter8));
  nand2 gate2068(.a(gate262inter8), .b(gate262inter7), .O(gate262inter9));
  nand2 gate2069(.a(s_217), .b(gate262inter3), .O(gate262inter10));
  nor2  gate2070(.a(gate262inter10), .b(gate262inter9), .O(gate262inter11));
  nor2  gate2071(.a(gate262inter11), .b(gate262inter6), .O(gate262inter12));
  nand2 gate2072(.a(gate262inter12), .b(gate262inter1), .O(G785));
nand2 gate263( .a(G766), .b(G767), .O(G788) );
nand2 gate264( .a(G768), .b(G769), .O(G791) );

  xor2  gate1373(.a(G770), .b(G642), .O(gate265inter0));
  nand2 gate1374(.a(gate265inter0), .b(s_118), .O(gate265inter1));
  and2  gate1375(.a(G770), .b(G642), .O(gate265inter2));
  inv1  gate1376(.a(s_118), .O(gate265inter3));
  inv1  gate1377(.a(s_119), .O(gate265inter4));
  nand2 gate1378(.a(gate265inter4), .b(gate265inter3), .O(gate265inter5));
  nor2  gate1379(.a(gate265inter5), .b(gate265inter2), .O(gate265inter6));
  inv1  gate1380(.a(G642), .O(gate265inter7));
  inv1  gate1381(.a(G770), .O(gate265inter8));
  nand2 gate1382(.a(gate265inter8), .b(gate265inter7), .O(gate265inter9));
  nand2 gate1383(.a(s_119), .b(gate265inter3), .O(gate265inter10));
  nor2  gate1384(.a(gate265inter10), .b(gate265inter9), .O(gate265inter11));
  nor2  gate1385(.a(gate265inter11), .b(gate265inter6), .O(gate265inter12));
  nand2 gate1386(.a(gate265inter12), .b(gate265inter1), .O(G794));
nand2 gate266( .a(G645), .b(G773), .O(G797) );
nand2 gate267( .a(G648), .b(G776), .O(G800) );
nand2 gate268( .a(G651), .b(G779), .O(G803) );
nand2 gate269( .a(G654), .b(G782), .O(G806) );

  xor2  gate2633(.a(G785), .b(G657), .O(gate270inter0));
  nand2 gate2634(.a(gate270inter0), .b(s_298), .O(gate270inter1));
  and2  gate2635(.a(G785), .b(G657), .O(gate270inter2));
  inv1  gate2636(.a(s_298), .O(gate270inter3));
  inv1  gate2637(.a(s_299), .O(gate270inter4));
  nand2 gate2638(.a(gate270inter4), .b(gate270inter3), .O(gate270inter5));
  nor2  gate2639(.a(gate270inter5), .b(gate270inter2), .O(gate270inter6));
  inv1  gate2640(.a(G657), .O(gate270inter7));
  inv1  gate2641(.a(G785), .O(gate270inter8));
  nand2 gate2642(.a(gate270inter8), .b(gate270inter7), .O(gate270inter9));
  nand2 gate2643(.a(s_299), .b(gate270inter3), .O(gate270inter10));
  nor2  gate2644(.a(gate270inter10), .b(gate270inter9), .O(gate270inter11));
  nor2  gate2645(.a(gate270inter11), .b(gate270inter6), .O(gate270inter12));
  nand2 gate2646(.a(gate270inter12), .b(gate270inter1), .O(G809));
nand2 gate271( .a(G660), .b(G788), .O(G812) );
nand2 gate272( .a(G663), .b(G791), .O(G815) );
nand2 gate273( .a(G642), .b(G794), .O(G818) );
nand2 gate274( .a(G770), .b(G794), .O(G819) );
nand2 gate275( .a(G645), .b(G797), .O(G820) );

  xor2  gate2381(.a(G797), .b(G773), .O(gate276inter0));
  nand2 gate2382(.a(gate276inter0), .b(s_262), .O(gate276inter1));
  and2  gate2383(.a(G797), .b(G773), .O(gate276inter2));
  inv1  gate2384(.a(s_262), .O(gate276inter3));
  inv1  gate2385(.a(s_263), .O(gate276inter4));
  nand2 gate2386(.a(gate276inter4), .b(gate276inter3), .O(gate276inter5));
  nor2  gate2387(.a(gate276inter5), .b(gate276inter2), .O(gate276inter6));
  inv1  gate2388(.a(G773), .O(gate276inter7));
  inv1  gate2389(.a(G797), .O(gate276inter8));
  nand2 gate2390(.a(gate276inter8), .b(gate276inter7), .O(gate276inter9));
  nand2 gate2391(.a(s_263), .b(gate276inter3), .O(gate276inter10));
  nor2  gate2392(.a(gate276inter10), .b(gate276inter9), .O(gate276inter11));
  nor2  gate2393(.a(gate276inter11), .b(gate276inter6), .O(gate276inter12));
  nand2 gate2394(.a(gate276inter12), .b(gate276inter1), .O(G821));
nand2 gate277( .a(G648), .b(G800), .O(G822) );
nand2 gate278( .a(G776), .b(G800), .O(G823) );
nand2 gate279( .a(G651), .b(G803), .O(G824) );

  xor2  gate2619(.a(G803), .b(G779), .O(gate280inter0));
  nand2 gate2620(.a(gate280inter0), .b(s_296), .O(gate280inter1));
  and2  gate2621(.a(G803), .b(G779), .O(gate280inter2));
  inv1  gate2622(.a(s_296), .O(gate280inter3));
  inv1  gate2623(.a(s_297), .O(gate280inter4));
  nand2 gate2624(.a(gate280inter4), .b(gate280inter3), .O(gate280inter5));
  nor2  gate2625(.a(gate280inter5), .b(gate280inter2), .O(gate280inter6));
  inv1  gate2626(.a(G779), .O(gate280inter7));
  inv1  gate2627(.a(G803), .O(gate280inter8));
  nand2 gate2628(.a(gate280inter8), .b(gate280inter7), .O(gate280inter9));
  nand2 gate2629(.a(s_297), .b(gate280inter3), .O(gate280inter10));
  nor2  gate2630(.a(gate280inter10), .b(gate280inter9), .O(gate280inter11));
  nor2  gate2631(.a(gate280inter11), .b(gate280inter6), .O(gate280inter12));
  nand2 gate2632(.a(gate280inter12), .b(gate280inter1), .O(G825));
nand2 gate281( .a(G654), .b(G806), .O(G826) );
nand2 gate282( .a(G782), .b(G806), .O(G827) );
nand2 gate283( .a(G657), .b(G809), .O(G828) );
nand2 gate284( .a(G785), .b(G809), .O(G829) );

  xor2  gate1499(.a(G812), .b(G660), .O(gate285inter0));
  nand2 gate1500(.a(gate285inter0), .b(s_136), .O(gate285inter1));
  and2  gate1501(.a(G812), .b(G660), .O(gate285inter2));
  inv1  gate1502(.a(s_136), .O(gate285inter3));
  inv1  gate1503(.a(s_137), .O(gate285inter4));
  nand2 gate1504(.a(gate285inter4), .b(gate285inter3), .O(gate285inter5));
  nor2  gate1505(.a(gate285inter5), .b(gate285inter2), .O(gate285inter6));
  inv1  gate1506(.a(G660), .O(gate285inter7));
  inv1  gate1507(.a(G812), .O(gate285inter8));
  nand2 gate1508(.a(gate285inter8), .b(gate285inter7), .O(gate285inter9));
  nand2 gate1509(.a(s_137), .b(gate285inter3), .O(gate285inter10));
  nor2  gate1510(.a(gate285inter10), .b(gate285inter9), .O(gate285inter11));
  nor2  gate1511(.a(gate285inter11), .b(gate285inter6), .O(gate285inter12));
  nand2 gate1512(.a(gate285inter12), .b(gate285inter1), .O(G830));

  xor2  gate2045(.a(G812), .b(G788), .O(gate286inter0));
  nand2 gate2046(.a(gate286inter0), .b(s_214), .O(gate286inter1));
  and2  gate2047(.a(G812), .b(G788), .O(gate286inter2));
  inv1  gate2048(.a(s_214), .O(gate286inter3));
  inv1  gate2049(.a(s_215), .O(gate286inter4));
  nand2 gate2050(.a(gate286inter4), .b(gate286inter3), .O(gate286inter5));
  nor2  gate2051(.a(gate286inter5), .b(gate286inter2), .O(gate286inter6));
  inv1  gate2052(.a(G788), .O(gate286inter7));
  inv1  gate2053(.a(G812), .O(gate286inter8));
  nand2 gate2054(.a(gate286inter8), .b(gate286inter7), .O(gate286inter9));
  nand2 gate2055(.a(s_215), .b(gate286inter3), .O(gate286inter10));
  nor2  gate2056(.a(gate286inter10), .b(gate286inter9), .O(gate286inter11));
  nor2  gate2057(.a(gate286inter11), .b(gate286inter6), .O(gate286inter12));
  nand2 gate2058(.a(gate286inter12), .b(gate286inter1), .O(G831));
nand2 gate287( .a(G663), .b(G815), .O(G832) );
nand2 gate288( .a(G791), .b(G815), .O(G833) );

  xor2  gate1695(.a(G819), .b(G818), .O(gate289inter0));
  nand2 gate1696(.a(gate289inter0), .b(s_164), .O(gate289inter1));
  and2  gate1697(.a(G819), .b(G818), .O(gate289inter2));
  inv1  gate1698(.a(s_164), .O(gate289inter3));
  inv1  gate1699(.a(s_165), .O(gate289inter4));
  nand2 gate1700(.a(gate289inter4), .b(gate289inter3), .O(gate289inter5));
  nor2  gate1701(.a(gate289inter5), .b(gate289inter2), .O(gate289inter6));
  inv1  gate1702(.a(G818), .O(gate289inter7));
  inv1  gate1703(.a(G819), .O(gate289inter8));
  nand2 gate1704(.a(gate289inter8), .b(gate289inter7), .O(gate289inter9));
  nand2 gate1705(.a(s_165), .b(gate289inter3), .O(gate289inter10));
  nor2  gate1706(.a(gate289inter10), .b(gate289inter9), .O(gate289inter11));
  nor2  gate1707(.a(gate289inter11), .b(gate289inter6), .O(gate289inter12));
  nand2 gate1708(.a(gate289inter12), .b(gate289inter1), .O(G834));
nand2 gate290( .a(G820), .b(G821), .O(G847) );

  xor2  gate1821(.a(G823), .b(G822), .O(gate291inter0));
  nand2 gate1822(.a(gate291inter0), .b(s_182), .O(gate291inter1));
  and2  gate1823(.a(G823), .b(G822), .O(gate291inter2));
  inv1  gate1824(.a(s_182), .O(gate291inter3));
  inv1  gate1825(.a(s_183), .O(gate291inter4));
  nand2 gate1826(.a(gate291inter4), .b(gate291inter3), .O(gate291inter5));
  nor2  gate1827(.a(gate291inter5), .b(gate291inter2), .O(gate291inter6));
  inv1  gate1828(.a(G822), .O(gate291inter7));
  inv1  gate1829(.a(G823), .O(gate291inter8));
  nand2 gate1830(.a(gate291inter8), .b(gate291inter7), .O(gate291inter9));
  nand2 gate1831(.a(s_183), .b(gate291inter3), .O(gate291inter10));
  nor2  gate1832(.a(gate291inter10), .b(gate291inter9), .O(gate291inter11));
  nor2  gate1833(.a(gate291inter11), .b(gate291inter6), .O(gate291inter12));
  nand2 gate1834(.a(gate291inter12), .b(gate291inter1), .O(G860));
nand2 gate292( .a(G824), .b(G825), .O(G873) );

  xor2  gate1513(.a(G829), .b(G828), .O(gate293inter0));
  nand2 gate1514(.a(gate293inter0), .b(s_138), .O(gate293inter1));
  and2  gate1515(.a(G829), .b(G828), .O(gate293inter2));
  inv1  gate1516(.a(s_138), .O(gate293inter3));
  inv1  gate1517(.a(s_139), .O(gate293inter4));
  nand2 gate1518(.a(gate293inter4), .b(gate293inter3), .O(gate293inter5));
  nor2  gate1519(.a(gate293inter5), .b(gate293inter2), .O(gate293inter6));
  inv1  gate1520(.a(G828), .O(gate293inter7));
  inv1  gate1521(.a(G829), .O(gate293inter8));
  nand2 gate1522(.a(gate293inter8), .b(gate293inter7), .O(gate293inter9));
  nand2 gate1523(.a(s_139), .b(gate293inter3), .O(gate293inter10));
  nor2  gate1524(.a(gate293inter10), .b(gate293inter9), .O(gate293inter11));
  nor2  gate1525(.a(gate293inter11), .b(gate293inter6), .O(gate293inter12));
  nand2 gate1526(.a(gate293inter12), .b(gate293inter1), .O(G886));
nand2 gate294( .a(G832), .b(G833), .O(G899) );

  xor2  gate2493(.a(G831), .b(G830), .O(gate295inter0));
  nand2 gate2494(.a(gate295inter0), .b(s_278), .O(gate295inter1));
  and2  gate2495(.a(G831), .b(G830), .O(gate295inter2));
  inv1  gate2496(.a(s_278), .O(gate295inter3));
  inv1  gate2497(.a(s_279), .O(gate295inter4));
  nand2 gate2498(.a(gate295inter4), .b(gate295inter3), .O(gate295inter5));
  nor2  gate2499(.a(gate295inter5), .b(gate295inter2), .O(gate295inter6));
  inv1  gate2500(.a(G830), .O(gate295inter7));
  inv1  gate2501(.a(G831), .O(gate295inter8));
  nand2 gate2502(.a(gate295inter8), .b(gate295inter7), .O(gate295inter9));
  nand2 gate2503(.a(s_279), .b(gate295inter3), .O(gate295inter10));
  nor2  gate2504(.a(gate295inter10), .b(gate295inter9), .O(gate295inter11));
  nor2  gate2505(.a(gate295inter11), .b(gate295inter6), .O(gate295inter12));
  nand2 gate2506(.a(gate295inter12), .b(gate295inter1), .O(G912));
nand2 gate296( .a(G826), .b(G827), .O(G925) );
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );

  xor2  gate603(.a(G1036), .b(G1), .O(gate387inter0));
  nand2 gate604(.a(gate387inter0), .b(s_8), .O(gate387inter1));
  and2  gate605(.a(G1036), .b(G1), .O(gate387inter2));
  inv1  gate606(.a(s_8), .O(gate387inter3));
  inv1  gate607(.a(s_9), .O(gate387inter4));
  nand2 gate608(.a(gate387inter4), .b(gate387inter3), .O(gate387inter5));
  nor2  gate609(.a(gate387inter5), .b(gate387inter2), .O(gate387inter6));
  inv1  gate610(.a(G1), .O(gate387inter7));
  inv1  gate611(.a(G1036), .O(gate387inter8));
  nand2 gate612(.a(gate387inter8), .b(gate387inter7), .O(gate387inter9));
  nand2 gate613(.a(s_9), .b(gate387inter3), .O(gate387inter10));
  nor2  gate614(.a(gate387inter10), .b(gate387inter9), .O(gate387inter11));
  nor2  gate615(.a(gate387inter11), .b(gate387inter6), .O(gate387inter12));
  nand2 gate616(.a(gate387inter12), .b(gate387inter1), .O(G1132));

  xor2  gate897(.a(G1039), .b(G2), .O(gate388inter0));
  nand2 gate898(.a(gate388inter0), .b(s_50), .O(gate388inter1));
  and2  gate899(.a(G1039), .b(G2), .O(gate388inter2));
  inv1  gate900(.a(s_50), .O(gate388inter3));
  inv1  gate901(.a(s_51), .O(gate388inter4));
  nand2 gate902(.a(gate388inter4), .b(gate388inter3), .O(gate388inter5));
  nor2  gate903(.a(gate388inter5), .b(gate388inter2), .O(gate388inter6));
  inv1  gate904(.a(G2), .O(gate388inter7));
  inv1  gate905(.a(G1039), .O(gate388inter8));
  nand2 gate906(.a(gate388inter8), .b(gate388inter7), .O(gate388inter9));
  nand2 gate907(.a(s_51), .b(gate388inter3), .O(gate388inter10));
  nor2  gate908(.a(gate388inter10), .b(gate388inter9), .O(gate388inter11));
  nor2  gate909(.a(gate388inter11), .b(gate388inter6), .O(gate388inter12));
  nand2 gate910(.a(gate388inter12), .b(gate388inter1), .O(G1135));

  xor2  gate1429(.a(G1042), .b(G3), .O(gate389inter0));
  nand2 gate1430(.a(gate389inter0), .b(s_126), .O(gate389inter1));
  and2  gate1431(.a(G1042), .b(G3), .O(gate389inter2));
  inv1  gate1432(.a(s_126), .O(gate389inter3));
  inv1  gate1433(.a(s_127), .O(gate389inter4));
  nand2 gate1434(.a(gate389inter4), .b(gate389inter3), .O(gate389inter5));
  nor2  gate1435(.a(gate389inter5), .b(gate389inter2), .O(gate389inter6));
  inv1  gate1436(.a(G3), .O(gate389inter7));
  inv1  gate1437(.a(G1042), .O(gate389inter8));
  nand2 gate1438(.a(gate389inter8), .b(gate389inter7), .O(gate389inter9));
  nand2 gate1439(.a(s_127), .b(gate389inter3), .O(gate389inter10));
  nor2  gate1440(.a(gate389inter10), .b(gate389inter9), .O(gate389inter11));
  nor2  gate1441(.a(gate389inter11), .b(gate389inter6), .O(gate389inter12));
  nand2 gate1442(.a(gate389inter12), .b(gate389inter1), .O(G1138));
nand2 gate390( .a(G4), .b(G1045), .O(G1141) );

  xor2  gate673(.a(G1048), .b(G5), .O(gate391inter0));
  nand2 gate674(.a(gate391inter0), .b(s_18), .O(gate391inter1));
  and2  gate675(.a(G1048), .b(G5), .O(gate391inter2));
  inv1  gate676(.a(s_18), .O(gate391inter3));
  inv1  gate677(.a(s_19), .O(gate391inter4));
  nand2 gate678(.a(gate391inter4), .b(gate391inter3), .O(gate391inter5));
  nor2  gate679(.a(gate391inter5), .b(gate391inter2), .O(gate391inter6));
  inv1  gate680(.a(G5), .O(gate391inter7));
  inv1  gate681(.a(G1048), .O(gate391inter8));
  nand2 gate682(.a(gate391inter8), .b(gate391inter7), .O(gate391inter9));
  nand2 gate683(.a(s_19), .b(gate391inter3), .O(gate391inter10));
  nor2  gate684(.a(gate391inter10), .b(gate391inter9), .O(gate391inter11));
  nor2  gate685(.a(gate391inter11), .b(gate391inter6), .O(gate391inter12));
  nand2 gate686(.a(gate391inter12), .b(gate391inter1), .O(G1144));
nand2 gate392( .a(G6), .b(G1051), .O(G1147) );
nand2 gate393( .a(G7), .b(G1054), .O(G1150) );

  xor2  gate1065(.a(G1057), .b(G8), .O(gate394inter0));
  nand2 gate1066(.a(gate394inter0), .b(s_74), .O(gate394inter1));
  and2  gate1067(.a(G1057), .b(G8), .O(gate394inter2));
  inv1  gate1068(.a(s_74), .O(gate394inter3));
  inv1  gate1069(.a(s_75), .O(gate394inter4));
  nand2 gate1070(.a(gate394inter4), .b(gate394inter3), .O(gate394inter5));
  nor2  gate1071(.a(gate394inter5), .b(gate394inter2), .O(gate394inter6));
  inv1  gate1072(.a(G8), .O(gate394inter7));
  inv1  gate1073(.a(G1057), .O(gate394inter8));
  nand2 gate1074(.a(gate394inter8), .b(gate394inter7), .O(gate394inter9));
  nand2 gate1075(.a(s_75), .b(gate394inter3), .O(gate394inter10));
  nor2  gate1076(.a(gate394inter10), .b(gate394inter9), .O(gate394inter11));
  nor2  gate1077(.a(gate394inter11), .b(gate394inter6), .O(gate394inter12));
  nand2 gate1078(.a(gate394inter12), .b(gate394inter1), .O(G1153));
nand2 gate395( .a(G9), .b(G1060), .O(G1156) );

  xor2  gate1961(.a(G1063), .b(G10), .O(gate396inter0));
  nand2 gate1962(.a(gate396inter0), .b(s_202), .O(gate396inter1));
  and2  gate1963(.a(G1063), .b(G10), .O(gate396inter2));
  inv1  gate1964(.a(s_202), .O(gate396inter3));
  inv1  gate1965(.a(s_203), .O(gate396inter4));
  nand2 gate1966(.a(gate396inter4), .b(gate396inter3), .O(gate396inter5));
  nor2  gate1967(.a(gate396inter5), .b(gate396inter2), .O(gate396inter6));
  inv1  gate1968(.a(G10), .O(gate396inter7));
  inv1  gate1969(.a(G1063), .O(gate396inter8));
  nand2 gate1970(.a(gate396inter8), .b(gate396inter7), .O(gate396inter9));
  nand2 gate1971(.a(s_203), .b(gate396inter3), .O(gate396inter10));
  nor2  gate1972(.a(gate396inter10), .b(gate396inter9), .O(gate396inter11));
  nor2  gate1973(.a(gate396inter11), .b(gate396inter6), .O(gate396inter12));
  nand2 gate1974(.a(gate396inter12), .b(gate396inter1), .O(G1159));

  xor2  gate2325(.a(G1066), .b(G11), .O(gate397inter0));
  nand2 gate2326(.a(gate397inter0), .b(s_254), .O(gate397inter1));
  and2  gate2327(.a(G1066), .b(G11), .O(gate397inter2));
  inv1  gate2328(.a(s_254), .O(gate397inter3));
  inv1  gate2329(.a(s_255), .O(gate397inter4));
  nand2 gate2330(.a(gate397inter4), .b(gate397inter3), .O(gate397inter5));
  nor2  gate2331(.a(gate397inter5), .b(gate397inter2), .O(gate397inter6));
  inv1  gate2332(.a(G11), .O(gate397inter7));
  inv1  gate2333(.a(G1066), .O(gate397inter8));
  nand2 gate2334(.a(gate397inter8), .b(gate397inter7), .O(gate397inter9));
  nand2 gate2335(.a(s_255), .b(gate397inter3), .O(gate397inter10));
  nor2  gate2336(.a(gate397inter10), .b(gate397inter9), .O(gate397inter11));
  nor2  gate2337(.a(gate397inter11), .b(gate397inter6), .O(gate397inter12));
  nand2 gate2338(.a(gate397inter12), .b(gate397inter1), .O(G1162));
nand2 gate398( .a(G12), .b(G1069), .O(G1165) );

  xor2  gate1709(.a(G1072), .b(G13), .O(gate399inter0));
  nand2 gate1710(.a(gate399inter0), .b(s_166), .O(gate399inter1));
  and2  gate1711(.a(G1072), .b(G13), .O(gate399inter2));
  inv1  gate1712(.a(s_166), .O(gate399inter3));
  inv1  gate1713(.a(s_167), .O(gate399inter4));
  nand2 gate1714(.a(gate399inter4), .b(gate399inter3), .O(gate399inter5));
  nor2  gate1715(.a(gate399inter5), .b(gate399inter2), .O(gate399inter6));
  inv1  gate1716(.a(G13), .O(gate399inter7));
  inv1  gate1717(.a(G1072), .O(gate399inter8));
  nand2 gate1718(.a(gate399inter8), .b(gate399inter7), .O(gate399inter9));
  nand2 gate1719(.a(s_167), .b(gate399inter3), .O(gate399inter10));
  nor2  gate1720(.a(gate399inter10), .b(gate399inter9), .O(gate399inter11));
  nor2  gate1721(.a(gate399inter11), .b(gate399inter6), .O(gate399inter12));
  nand2 gate1722(.a(gate399inter12), .b(gate399inter1), .O(G1168));
nand2 gate400( .a(G14), .b(G1075), .O(G1171) );

  xor2  gate2115(.a(G1078), .b(G15), .O(gate401inter0));
  nand2 gate2116(.a(gate401inter0), .b(s_224), .O(gate401inter1));
  and2  gate2117(.a(G1078), .b(G15), .O(gate401inter2));
  inv1  gate2118(.a(s_224), .O(gate401inter3));
  inv1  gate2119(.a(s_225), .O(gate401inter4));
  nand2 gate2120(.a(gate401inter4), .b(gate401inter3), .O(gate401inter5));
  nor2  gate2121(.a(gate401inter5), .b(gate401inter2), .O(gate401inter6));
  inv1  gate2122(.a(G15), .O(gate401inter7));
  inv1  gate2123(.a(G1078), .O(gate401inter8));
  nand2 gate2124(.a(gate401inter8), .b(gate401inter7), .O(gate401inter9));
  nand2 gate2125(.a(s_225), .b(gate401inter3), .O(gate401inter10));
  nor2  gate2126(.a(gate401inter10), .b(gate401inter9), .O(gate401inter11));
  nor2  gate2127(.a(gate401inter11), .b(gate401inter6), .O(gate401inter12));
  nand2 gate2128(.a(gate401inter12), .b(gate401inter1), .O(G1174));
nand2 gate402( .a(G16), .b(G1081), .O(G1177) );
nand2 gate403( .a(G17), .b(G1084), .O(G1180) );

  xor2  gate2451(.a(G1087), .b(G18), .O(gate404inter0));
  nand2 gate2452(.a(gate404inter0), .b(s_272), .O(gate404inter1));
  and2  gate2453(.a(G1087), .b(G18), .O(gate404inter2));
  inv1  gate2454(.a(s_272), .O(gate404inter3));
  inv1  gate2455(.a(s_273), .O(gate404inter4));
  nand2 gate2456(.a(gate404inter4), .b(gate404inter3), .O(gate404inter5));
  nor2  gate2457(.a(gate404inter5), .b(gate404inter2), .O(gate404inter6));
  inv1  gate2458(.a(G18), .O(gate404inter7));
  inv1  gate2459(.a(G1087), .O(gate404inter8));
  nand2 gate2460(.a(gate404inter8), .b(gate404inter7), .O(gate404inter9));
  nand2 gate2461(.a(s_273), .b(gate404inter3), .O(gate404inter10));
  nor2  gate2462(.a(gate404inter10), .b(gate404inter9), .O(gate404inter11));
  nor2  gate2463(.a(gate404inter11), .b(gate404inter6), .O(gate404inter12));
  nand2 gate2464(.a(gate404inter12), .b(gate404inter1), .O(G1183));
nand2 gate405( .a(G19), .b(G1090), .O(G1186) );
nand2 gate406( .a(G20), .b(G1093), .O(G1189) );
nand2 gate407( .a(G21), .b(G1096), .O(G1192) );

  xor2  gate925(.a(G1099), .b(G22), .O(gate408inter0));
  nand2 gate926(.a(gate408inter0), .b(s_54), .O(gate408inter1));
  and2  gate927(.a(G1099), .b(G22), .O(gate408inter2));
  inv1  gate928(.a(s_54), .O(gate408inter3));
  inv1  gate929(.a(s_55), .O(gate408inter4));
  nand2 gate930(.a(gate408inter4), .b(gate408inter3), .O(gate408inter5));
  nor2  gate931(.a(gate408inter5), .b(gate408inter2), .O(gate408inter6));
  inv1  gate932(.a(G22), .O(gate408inter7));
  inv1  gate933(.a(G1099), .O(gate408inter8));
  nand2 gate934(.a(gate408inter8), .b(gate408inter7), .O(gate408inter9));
  nand2 gate935(.a(s_55), .b(gate408inter3), .O(gate408inter10));
  nor2  gate936(.a(gate408inter10), .b(gate408inter9), .O(gate408inter11));
  nor2  gate937(.a(gate408inter11), .b(gate408inter6), .O(gate408inter12));
  nand2 gate938(.a(gate408inter12), .b(gate408inter1), .O(G1195));

  xor2  gate1569(.a(G1102), .b(G23), .O(gate409inter0));
  nand2 gate1570(.a(gate409inter0), .b(s_146), .O(gate409inter1));
  and2  gate1571(.a(G1102), .b(G23), .O(gate409inter2));
  inv1  gate1572(.a(s_146), .O(gate409inter3));
  inv1  gate1573(.a(s_147), .O(gate409inter4));
  nand2 gate1574(.a(gate409inter4), .b(gate409inter3), .O(gate409inter5));
  nor2  gate1575(.a(gate409inter5), .b(gate409inter2), .O(gate409inter6));
  inv1  gate1576(.a(G23), .O(gate409inter7));
  inv1  gate1577(.a(G1102), .O(gate409inter8));
  nand2 gate1578(.a(gate409inter8), .b(gate409inter7), .O(gate409inter9));
  nand2 gate1579(.a(s_147), .b(gate409inter3), .O(gate409inter10));
  nor2  gate1580(.a(gate409inter10), .b(gate409inter9), .O(gate409inter11));
  nor2  gate1581(.a(gate409inter11), .b(gate409inter6), .O(gate409inter12));
  nand2 gate1582(.a(gate409inter12), .b(gate409inter1), .O(G1198));
nand2 gate410( .a(G24), .b(G1105), .O(G1201) );

  xor2  gate2171(.a(G1108), .b(G25), .O(gate411inter0));
  nand2 gate2172(.a(gate411inter0), .b(s_232), .O(gate411inter1));
  and2  gate2173(.a(G1108), .b(G25), .O(gate411inter2));
  inv1  gate2174(.a(s_232), .O(gate411inter3));
  inv1  gate2175(.a(s_233), .O(gate411inter4));
  nand2 gate2176(.a(gate411inter4), .b(gate411inter3), .O(gate411inter5));
  nor2  gate2177(.a(gate411inter5), .b(gate411inter2), .O(gate411inter6));
  inv1  gate2178(.a(G25), .O(gate411inter7));
  inv1  gate2179(.a(G1108), .O(gate411inter8));
  nand2 gate2180(.a(gate411inter8), .b(gate411inter7), .O(gate411inter9));
  nand2 gate2181(.a(s_233), .b(gate411inter3), .O(gate411inter10));
  nor2  gate2182(.a(gate411inter10), .b(gate411inter9), .O(gate411inter11));
  nor2  gate2183(.a(gate411inter11), .b(gate411inter6), .O(gate411inter12));
  nand2 gate2184(.a(gate411inter12), .b(gate411inter1), .O(G1204));
nand2 gate412( .a(G26), .b(G1111), .O(G1207) );
nand2 gate413( .a(G27), .b(G1114), .O(G1210) );
nand2 gate414( .a(G28), .b(G1117), .O(G1213) );
nand2 gate415( .a(G29), .b(G1120), .O(G1216) );

  xor2  gate911(.a(G1123), .b(G30), .O(gate416inter0));
  nand2 gate912(.a(gate416inter0), .b(s_52), .O(gate416inter1));
  and2  gate913(.a(G1123), .b(G30), .O(gate416inter2));
  inv1  gate914(.a(s_52), .O(gate416inter3));
  inv1  gate915(.a(s_53), .O(gate416inter4));
  nand2 gate916(.a(gate416inter4), .b(gate416inter3), .O(gate416inter5));
  nor2  gate917(.a(gate416inter5), .b(gate416inter2), .O(gate416inter6));
  inv1  gate918(.a(G30), .O(gate416inter7));
  inv1  gate919(.a(G1123), .O(gate416inter8));
  nand2 gate920(.a(gate416inter8), .b(gate416inter7), .O(gate416inter9));
  nand2 gate921(.a(s_53), .b(gate416inter3), .O(gate416inter10));
  nor2  gate922(.a(gate416inter10), .b(gate416inter9), .O(gate416inter11));
  nor2  gate923(.a(gate416inter11), .b(gate416inter6), .O(gate416inter12));
  nand2 gate924(.a(gate416inter12), .b(gate416inter1), .O(G1219));

  xor2  gate771(.a(G1126), .b(G31), .O(gate417inter0));
  nand2 gate772(.a(gate417inter0), .b(s_32), .O(gate417inter1));
  and2  gate773(.a(G1126), .b(G31), .O(gate417inter2));
  inv1  gate774(.a(s_32), .O(gate417inter3));
  inv1  gate775(.a(s_33), .O(gate417inter4));
  nand2 gate776(.a(gate417inter4), .b(gate417inter3), .O(gate417inter5));
  nor2  gate777(.a(gate417inter5), .b(gate417inter2), .O(gate417inter6));
  inv1  gate778(.a(G31), .O(gate417inter7));
  inv1  gate779(.a(G1126), .O(gate417inter8));
  nand2 gate780(.a(gate417inter8), .b(gate417inter7), .O(gate417inter9));
  nand2 gate781(.a(s_33), .b(gate417inter3), .O(gate417inter10));
  nor2  gate782(.a(gate417inter10), .b(gate417inter9), .O(gate417inter11));
  nor2  gate783(.a(gate417inter11), .b(gate417inter6), .O(gate417inter12));
  nand2 gate784(.a(gate417inter12), .b(gate417inter1), .O(G1222));
nand2 gate418( .a(G32), .b(G1129), .O(G1225) );
nand2 gate419( .a(G1), .b(G1132), .O(G1228) );
nand2 gate420( .a(G1036), .b(G1132), .O(G1229) );

  xor2  gate2479(.a(G1135), .b(G2), .O(gate421inter0));
  nand2 gate2480(.a(gate421inter0), .b(s_276), .O(gate421inter1));
  and2  gate2481(.a(G1135), .b(G2), .O(gate421inter2));
  inv1  gate2482(.a(s_276), .O(gate421inter3));
  inv1  gate2483(.a(s_277), .O(gate421inter4));
  nand2 gate2484(.a(gate421inter4), .b(gate421inter3), .O(gate421inter5));
  nor2  gate2485(.a(gate421inter5), .b(gate421inter2), .O(gate421inter6));
  inv1  gate2486(.a(G2), .O(gate421inter7));
  inv1  gate2487(.a(G1135), .O(gate421inter8));
  nand2 gate2488(.a(gate421inter8), .b(gate421inter7), .O(gate421inter9));
  nand2 gate2489(.a(s_277), .b(gate421inter3), .O(gate421inter10));
  nor2  gate2490(.a(gate421inter10), .b(gate421inter9), .O(gate421inter11));
  nor2  gate2491(.a(gate421inter11), .b(gate421inter6), .O(gate421inter12));
  nand2 gate2492(.a(gate421inter12), .b(gate421inter1), .O(G1230));
nand2 gate422( .a(G1039), .b(G1135), .O(G1231) );
nand2 gate423( .a(G3), .b(G1138), .O(G1232) );
nand2 gate424( .a(G1042), .b(G1138), .O(G1233) );

  xor2  gate1737(.a(G1141), .b(G4), .O(gate425inter0));
  nand2 gate1738(.a(gate425inter0), .b(s_170), .O(gate425inter1));
  and2  gate1739(.a(G1141), .b(G4), .O(gate425inter2));
  inv1  gate1740(.a(s_170), .O(gate425inter3));
  inv1  gate1741(.a(s_171), .O(gate425inter4));
  nand2 gate1742(.a(gate425inter4), .b(gate425inter3), .O(gate425inter5));
  nor2  gate1743(.a(gate425inter5), .b(gate425inter2), .O(gate425inter6));
  inv1  gate1744(.a(G4), .O(gate425inter7));
  inv1  gate1745(.a(G1141), .O(gate425inter8));
  nand2 gate1746(.a(gate425inter8), .b(gate425inter7), .O(gate425inter9));
  nand2 gate1747(.a(s_171), .b(gate425inter3), .O(gate425inter10));
  nor2  gate1748(.a(gate425inter10), .b(gate425inter9), .O(gate425inter11));
  nor2  gate1749(.a(gate425inter11), .b(gate425inter6), .O(gate425inter12));
  nand2 gate1750(.a(gate425inter12), .b(gate425inter1), .O(G1234));

  xor2  gate2227(.a(G1141), .b(G1045), .O(gate426inter0));
  nand2 gate2228(.a(gate426inter0), .b(s_240), .O(gate426inter1));
  and2  gate2229(.a(G1141), .b(G1045), .O(gate426inter2));
  inv1  gate2230(.a(s_240), .O(gate426inter3));
  inv1  gate2231(.a(s_241), .O(gate426inter4));
  nand2 gate2232(.a(gate426inter4), .b(gate426inter3), .O(gate426inter5));
  nor2  gate2233(.a(gate426inter5), .b(gate426inter2), .O(gate426inter6));
  inv1  gate2234(.a(G1045), .O(gate426inter7));
  inv1  gate2235(.a(G1141), .O(gate426inter8));
  nand2 gate2236(.a(gate426inter8), .b(gate426inter7), .O(gate426inter9));
  nand2 gate2237(.a(s_241), .b(gate426inter3), .O(gate426inter10));
  nor2  gate2238(.a(gate426inter10), .b(gate426inter9), .O(gate426inter11));
  nor2  gate2239(.a(gate426inter11), .b(gate426inter6), .O(gate426inter12));
  nand2 gate2240(.a(gate426inter12), .b(gate426inter1), .O(G1235));

  xor2  gate785(.a(G1144), .b(G5), .O(gate427inter0));
  nand2 gate786(.a(gate427inter0), .b(s_34), .O(gate427inter1));
  and2  gate787(.a(G1144), .b(G5), .O(gate427inter2));
  inv1  gate788(.a(s_34), .O(gate427inter3));
  inv1  gate789(.a(s_35), .O(gate427inter4));
  nand2 gate790(.a(gate427inter4), .b(gate427inter3), .O(gate427inter5));
  nor2  gate791(.a(gate427inter5), .b(gate427inter2), .O(gate427inter6));
  inv1  gate792(.a(G5), .O(gate427inter7));
  inv1  gate793(.a(G1144), .O(gate427inter8));
  nand2 gate794(.a(gate427inter8), .b(gate427inter7), .O(gate427inter9));
  nand2 gate795(.a(s_35), .b(gate427inter3), .O(gate427inter10));
  nor2  gate796(.a(gate427inter10), .b(gate427inter9), .O(gate427inter11));
  nor2  gate797(.a(gate427inter11), .b(gate427inter6), .O(gate427inter12));
  nand2 gate798(.a(gate427inter12), .b(gate427inter1), .O(G1236));
nand2 gate428( .a(G1048), .b(G1144), .O(G1237) );
nand2 gate429( .a(G6), .b(G1147), .O(G1238) );
nand2 gate430( .a(G1051), .b(G1147), .O(G1239) );

  xor2  gate1849(.a(G1150), .b(G7), .O(gate431inter0));
  nand2 gate1850(.a(gate431inter0), .b(s_186), .O(gate431inter1));
  and2  gate1851(.a(G1150), .b(G7), .O(gate431inter2));
  inv1  gate1852(.a(s_186), .O(gate431inter3));
  inv1  gate1853(.a(s_187), .O(gate431inter4));
  nand2 gate1854(.a(gate431inter4), .b(gate431inter3), .O(gate431inter5));
  nor2  gate1855(.a(gate431inter5), .b(gate431inter2), .O(gate431inter6));
  inv1  gate1856(.a(G7), .O(gate431inter7));
  inv1  gate1857(.a(G1150), .O(gate431inter8));
  nand2 gate1858(.a(gate431inter8), .b(gate431inter7), .O(gate431inter9));
  nand2 gate1859(.a(s_187), .b(gate431inter3), .O(gate431inter10));
  nor2  gate1860(.a(gate431inter10), .b(gate431inter9), .O(gate431inter11));
  nor2  gate1861(.a(gate431inter11), .b(gate431inter6), .O(gate431inter12));
  nand2 gate1862(.a(gate431inter12), .b(gate431inter1), .O(G1240));
nand2 gate432( .a(G1054), .b(G1150), .O(G1241) );
nand2 gate433( .a(G8), .b(G1153), .O(G1242) );

  xor2  gate1611(.a(G1153), .b(G1057), .O(gate434inter0));
  nand2 gate1612(.a(gate434inter0), .b(s_152), .O(gate434inter1));
  and2  gate1613(.a(G1153), .b(G1057), .O(gate434inter2));
  inv1  gate1614(.a(s_152), .O(gate434inter3));
  inv1  gate1615(.a(s_153), .O(gate434inter4));
  nand2 gate1616(.a(gate434inter4), .b(gate434inter3), .O(gate434inter5));
  nor2  gate1617(.a(gate434inter5), .b(gate434inter2), .O(gate434inter6));
  inv1  gate1618(.a(G1057), .O(gate434inter7));
  inv1  gate1619(.a(G1153), .O(gate434inter8));
  nand2 gate1620(.a(gate434inter8), .b(gate434inter7), .O(gate434inter9));
  nand2 gate1621(.a(s_153), .b(gate434inter3), .O(gate434inter10));
  nor2  gate1622(.a(gate434inter10), .b(gate434inter9), .O(gate434inter11));
  nor2  gate1623(.a(gate434inter11), .b(gate434inter6), .O(gate434inter12));
  nand2 gate1624(.a(gate434inter12), .b(gate434inter1), .O(G1243));
nand2 gate435( .a(G9), .b(G1156), .O(G1244) );
nand2 gate436( .a(G1060), .b(G1156), .O(G1245) );
nand2 gate437( .a(G10), .b(G1159), .O(G1246) );
nand2 gate438( .a(G1063), .b(G1159), .O(G1247) );
nand2 gate439( .a(G11), .b(G1162), .O(G1248) );
nand2 gate440( .a(G1066), .b(G1162), .O(G1249) );
nand2 gate441( .a(G12), .b(G1165), .O(G1250) );
nand2 gate442( .a(G1069), .b(G1165), .O(G1251) );
nand2 gate443( .a(G13), .b(G1168), .O(G1252) );
nand2 gate444( .a(G1072), .b(G1168), .O(G1253) );
nand2 gate445( .a(G14), .b(G1171), .O(G1254) );
nand2 gate446( .a(G1075), .b(G1171), .O(G1255) );

  xor2  gate1275(.a(G1174), .b(G15), .O(gate447inter0));
  nand2 gate1276(.a(gate447inter0), .b(s_104), .O(gate447inter1));
  and2  gate1277(.a(G1174), .b(G15), .O(gate447inter2));
  inv1  gate1278(.a(s_104), .O(gate447inter3));
  inv1  gate1279(.a(s_105), .O(gate447inter4));
  nand2 gate1280(.a(gate447inter4), .b(gate447inter3), .O(gate447inter5));
  nor2  gate1281(.a(gate447inter5), .b(gate447inter2), .O(gate447inter6));
  inv1  gate1282(.a(G15), .O(gate447inter7));
  inv1  gate1283(.a(G1174), .O(gate447inter8));
  nand2 gate1284(.a(gate447inter8), .b(gate447inter7), .O(gate447inter9));
  nand2 gate1285(.a(s_105), .b(gate447inter3), .O(gate447inter10));
  nor2  gate1286(.a(gate447inter10), .b(gate447inter9), .O(gate447inter11));
  nor2  gate1287(.a(gate447inter11), .b(gate447inter6), .O(gate447inter12));
  nand2 gate1288(.a(gate447inter12), .b(gate447inter1), .O(G1256));

  xor2  gate2311(.a(G1174), .b(G1078), .O(gate448inter0));
  nand2 gate2312(.a(gate448inter0), .b(s_252), .O(gate448inter1));
  and2  gate2313(.a(G1174), .b(G1078), .O(gate448inter2));
  inv1  gate2314(.a(s_252), .O(gate448inter3));
  inv1  gate2315(.a(s_253), .O(gate448inter4));
  nand2 gate2316(.a(gate448inter4), .b(gate448inter3), .O(gate448inter5));
  nor2  gate2317(.a(gate448inter5), .b(gate448inter2), .O(gate448inter6));
  inv1  gate2318(.a(G1078), .O(gate448inter7));
  inv1  gate2319(.a(G1174), .O(gate448inter8));
  nand2 gate2320(.a(gate448inter8), .b(gate448inter7), .O(gate448inter9));
  nand2 gate2321(.a(s_253), .b(gate448inter3), .O(gate448inter10));
  nor2  gate2322(.a(gate448inter10), .b(gate448inter9), .O(gate448inter11));
  nor2  gate2323(.a(gate448inter11), .b(gate448inter6), .O(gate448inter12));
  nand2 gate2324(.a(gate448inter12), .b(gate448inter1), .O(G1257));
nand2 gate449( .a(G16), .b(G1177), .O(G1258) );
nand2 gate450( .a(G1081), .b(G1177), .O(G1259) );
nand2 gate451( .a(G17), .b(G1180), .O(G1260) );
nand2 gate452( .a(G1084), .b(G1180), .O(G1261) );
nand2 gate453( .a(G18), .b(G1183), .O(G1262) );

  xor2  gate2255(.a(G1183), .b(G1087), .O(gate454inter0));
  nand2 gate2256(.a(gate454inter0), .b(s_244), .O(gate454inter1));
  and2  gate2257(.a(G1183), .b(G1087), .O(gate454inter2));
  inv1  gate2258(.a(s_244), .O(gate454inter3));
  inv1  gate2259(.a(s_245), .O(gate454inter4));
  nand2 gate2260(.a(gate454inter4), .b(gate454inter3), .O(gate454inter5));
  nor2  gate2261(.a(gate454inter5), .b(gate454inter2), .O(gate454inter6));
  inv1  gate2262(.a(G1087), .O(gate454inter7));
  inv1  gate2263(.a(G1183), .O(gate454inter8));
  nand2 gate2264(.a(gate454inter8), .b(gate454inter7), .O(gate454inter9));
  nand2 gate2265(.a(s_245), .b(gate454inter3), .O(gate454inter10));
  nor2  gate2266(.a(gate454inter10), .b(gate454inter9), .O(gate454inter11));
  nor2  gate2267(.a(gate454inter11), .b(gate454inter6), .O(gate454inter12));
  nand2 gate2268(.a(gate454inter12), .b(gate454inter1), .O(G1263));

  xor2  gate729(.a(G1186), .b(G19), .O(gate455inter0));
  nand2 gate730(.a(gate455inter0), .b(s_26), .O(gate455inter1));
  and2  gate731(.a(G1186), .b(G19), .O(gate455inter2));
  inv1  gate732(.a(s_26), .O(gate455inter3));
  inv1  gate733(.a(s_27), .O(gate455inter4));
  nand2 gate734(.a(gate455inter4), .b(gate455inter3), .O(gate455inter5));
  nor2  gate735(.a(gate455inter5), .b(gate455inter2), .O(gate455inter6));
  inv1  gate736(.a(G19), .O(gate455inter7));
  inv1  gate737(.a(G1186), .O(gate455inter8));
  nand2 gate738(.a(gate455inter8), .b(gate455inter7), .O(gate455inter9));
  nand2 gate739(.a(s_27), .b(gate455inter3), .O(gate455inter10));
  nor2  gate740(.a(gate455inter10), .b(gate455inter9), .O(gate455inter11));
  nor2  gate741(.a(gate455inter11), .b(gate455inter6), .O(gate455inter12));
  nand2 gate742(.a(gate455inter12), .b(gate455inter1), .O(G1264));

  xor2  gate1541(.a(G1186), .b(G1090), .O(gate456inter0));
  nand2 gate1542(.a(gate456inter0), .b(s_142), .O(gate456inter1));
  and2  gate1543(.a(G1186), .b(G1090), .O(gate456inter2));
  inv1  gate1544(.a(s_142), .O(gate456inter3));
  inv1  gate1545(.a(s_143), .O(gate456inter4));
  nand2 gate1546(.a(gate456inter4), .b(gate456inter3), .O(gate456inter5));
  nor2  gate1547(.a(gate456inter5), .b(gate456inter2), .O(gate456inter6));
  inv1  gate1548(.a(G1090), .O(gate456inter7));
  inv1  gate1549(.a(G1186), .O(gate456inter8));
  nand2 gate1550(.a(gate456inter8), .b(gate456inter7), .O(gate456inter9));
  nand2 gate1551(.a(s_143), .b(gate456inter3), .O(gate456inter10));
  nor2  gate1552(.a(gate456inter10), .b(gate456inter9), .O(gate456inter11));
  nor2  gate1553(.a(gate456inter11), .b(gate456inter6), .O(gate456inter12));
  nand2 gate1554(.a(gate456inter12), .b(gate456inter1), .O(G1265));
nand2 gate457( .a(G20), .b(G1189), .O(G1266) );
nand2 gate458( .a(G1093), .b(G1189), .O(G1267) );
nand2 gate459( .a(G21), .b(G1192), .O(G1268) );

  xor2  gate995(.a(G1192), .b(G1096), .O(gate460inter0));
  nand2 gate996(.a(gate460inter0), .b(s_64), .O(gate460inter1));
  and2  gate997(.a(G1192), .b(G1096), .O(gate460inter2));
  inv1  gate998(.a(s_64), .O(gate460inter3));
  inv1  gate999(.a(s_65), .O(gate460inter4));
  nand2 gate1000(.a(gate460inter4), .b(gate460inter3), .O(gate460inter5));
  nor2  gate1001(.a(gate460inter5), .b(gate460inter2), .O(gate460inter6));
  inv1  gate1002(.a(G1096), .O(gate460inter7));
  inv1  gate1003(.a(G1192), .O(gate460inter8));
  nand2 gate1004(.a(gate460inter8), .b(gate460inter7), .O(gate460inter9));
  nand2 gate1005(.a(s_65), .b(gate460inter3), .O(gate460inter10));
  nor2  gate1006(.a(gate460inter10), .b(gate460inter9), .O(gate460inter11));
  nor2  gate1007(.a(gate460inter11), .b(gate460inter6), .O(gate460inter12));
  nand2 gate1008(.a(gate460inter12), .b(gate460inter1), .O(G1269));
nand2 gate461( .a(G22), .b(G1195), .O(G1270) );
nand2 gate462( .a(G1099), .b(G1195), .O(G1271) );

  xor2  gate2129(.a(G1198), .b(G23), .O(gate463inter0));
  nand2 gate2130(.a(gate463inter0), .b(s_226), .O(gate463inter1));
  and2  gate2131(.a(G1198), .b(G23), .O(gate463inter2));
  inv1  gate2132(.a(s_226), .O(gate463inter3));
  inv1  gate2133(.a(s_227), .O(gate463inter4));
  nand2 gate2134(.a(gate463inter4), .b(gate463inter3), .O(gate463inter5));
  nor2  gate2135(.a(gate463inter5), .b(gate463inter2), .O(gate463inter6));
  inv1  gate2136(.a(G23), .O(gate463inter7));
  inv1  gate2137(.a(G1198), .O(gate463inter8));
  nand2 gate2138(.a(gate463inter8), .b(gate463inter7), .O(gate463inter9));
  nand2 gate2139(.a(s_227), .b(gate463inter3), .O(gate463inter10));
  nor2  gate2140(.a(gate463inter10), .b(gate463inter9), .O(gate463inter11));
  nor2  gate2141(.a(gate463inter11), .b(gate463inter6), .O(gate463inter12));
  nand2 gate2142(.a(gate463inter12), .b(gate463inter1), .O(G1272));

  xor2  gate1989(.a(G1198), .b(G1102), .O(gate464inter0));
  nand2 gate1990(.a(gate464inter0), .b(s_206), .O(gate464inter1));
  and2  gate1991(.a(G1198), .b(G1102), .O(gate464inter2));
  inv1  gate1992(.a(s_206), .O(gate464inter3));
  inv1  gate1993(.a(s_207), .O(gate464inter4));
  nand2 gate1994(.a(gate464inter4), .b(gate464inter3), .O(gate464inter5));
  nor2  gate1995(.a(gate464inter5), .b(gate464inter2), .O(gate464inter6));
  inv1  gate1996(.a(G1102), .O(gate464inter7));
  inv1  gate1997(.a(G1198), .O(gate464inter8));
  nand2 gate1998(.a(gate464inter8), .b(gate464inter7), .O(gate464inter9));
  nand2 gate1999(.a(s_207), .b(gate464inter3), .O(gate464inter10));
  nor2  gate2000(.a(gate464inter10), .b(gate464inter9), .O(gate464inter11));
  nor2  gate2001(.a(gate464inter11), .b(gate464inter6), .O(gate464inter12));
  nand2 gate2002(.a(gate464inter12), .b(gate464inter1), .O(G1273));
nand2 gate465( .a(G24), .b(G1201), .O(G1274) );
nand2 gate466( .a(G1105), .b(G1201), .O(G1275) );
nand2 gate467( .a(G25), .b(G1204), .O(G1276) );
nand2 gate468( .a(G1108), .b(G1204), .O(G1277) );

  xor2  gate1317(.a(G1207), .b(G26), .O(gate469inter0));
  nand2 gate1318(.a(gate469inter0), .b(s_110), .O(gate469inter1));
  and2  gate1319(.a(G1207), .b(G26), .O(gate469inter2));
  inv1  gate1320(.a(s_110), .O(gate469inter3));
  inv1  gate1321(.a(s_111), .O(gate469inter4));
  nand2 gate1322(.a(gate469inter4), .b(gate469inter3), .O(gate469inter5));
  nor2  gate1323(.a(gate469inter5), .b(gate469inter2), .O(gate469inter6));
  inv1  gate1324(.a(G26), .O(gate469inter7));
  inv1  gate1325(.a(G1207), .O(gate469inter8));
  nand2 gate1326(.a(gate469inter8), .b(gate469inter7), .O(gate469inter9));
  nand2 gate1327(.a(s_111), .b(gate469inter3), .O(gate469inter10));
  nor2  gate1328(.a(gate469inter10), .b(gate469inter9), .O(gate469inter11));
  nor2  gate1329(.a(gate469inter11), .b(gate469inter6), .O(gate469inter12));
  nand2 gate1330(.a(gate469inter12), .b(gate469inter1), .O(G1278));
nand2 gate470( .a(G1111), .b(G1207), .O(G1279) );
nand2 gate471( .a(G27), .b(G1210), .O(G1280) );
nand2 gate472( .a(G1114), .b(G1210), .O(G1281) );

  xor2  gate953(.a(G1213), .b(G28), .O(gate473inter0));
  nand2 gate954(.a(gate473inter0), .b(s_58), .O(gate473inter1));
  and2  gate955(.a(G1213), .b(G28), .O(gate473inter2));
  inv1  gate956(.a(s_58), .O(gate473inter3));
  inv1  gate957(.a(s_59), .O(gate473inter4));
  nand2 gate958(.a(gate473inter4), .b(gate473inter3), .O(gate473inter5));
  nor2  gate959(.a(gate473inter5), .b(gate473inter2), .O(gate473inter6));
  inv1  gate960(.a(G28), .O(gate473inter7));
  inv1  gate961(.a(G1213), .O(gate473inter8));
  nand2 gate962(.a(gate473inter8), .b(gate473inter7), .O(gate473inter9));
  nand2 gate963(.a(s_59), .b(gate473inter3), .O(gate473inter10));
  nor2  gate964(.a(gate473inter10), .b(gate473inter9), .O(gate473inter11));
  nor2  gate965(.a(gate473inter11), .b(gate473inter6), .O(gate473inter12));
  nand2 gate966(.a(gate473inter12), .b(gate473inter1), .O(G1282));
nand2 gate474( .a(G1117), .b(G1213), .O(G1283) );
nand2 gate475( .a(G29), .b(G1216), .O(G1284) );

  xor2  gate1289(.a(G1216), .b(G1120), .O(gate476inter0));
  nand2 gate1290(.a(gate476inter0), .b(s_106), .O(gate476inter1));
  and2  gate1291(.a(G1216), .b(G1120), .O(gate476inter2));
  inv1  gate1292(.a(s_106), .O(gate476inter3));
  inv1  gate1293(.a(s_107), .O(gate476inter4));
  nand2 gate1294(.a(gate476inter4), .b(gate476inter3), .O(gate476inter5));
  nor2  gate1295(.a(gate476inter5), .b(gate476inter2), .O(gate476inter6));
  inv1  gate1296(.a(G1120), .O(gate476inter7));
  inv1  gate1297(.a(G1216), .O(gate476inter8));
  nand2 gate1298(.a(gate476inter8), .b(gate476inter7), .O(gate476inter9));
  nand2 gate1299(.a(s_107), .b(gate476inter3), .O(gate476inter10));
  nor2  gate1300(.a(gate476inter10), .b(gate476inter9), .O(gate476inter11));
  nor2  gate1301(.a(gate476inter11), .b(gate476inter6), .O(gate476inter12));
  nand2 gate1302(.a(gate476inter12), .b(gate476inter1), .O(G1285));
nand2 gate477( .a(G30), .b(G1219), .O(G1286) );
nand2 gate478( .a(G1123), .b(G1219), .O(G1287) );

  xor2  gate2367(.a(G1222), .b(G31), .O(gate479inter0));
  nand2 gate2368(.a(gate479inter0), .b(s_260), .O(gate479inter1));
  and2  gate2369(.a(G1222), .b(G31), .O(gate479inter2));
  inv1  gate2370(.a(s_260), .O(gate479inter3));
  inv1  gate2371(.a(s_261), .O(gate479inter4));
  nand2 gate2372(.a(gate479inter4), .b(gate479inter3), .O(gate479inter5));
  nor2  gate2373(.a(gate479inter5), .b(gate479inter2), .O(gate479inter6));
  inv1  gate2374(.a(G31), .O(gate479inter7));
  inv1  gate2375(.a(G1222), .O(gate479inter8));
  nand2 gate2376(.a(gate479inter8), .b(gate479inter7), .O(gate479inter9));
  nand2 gate2377(.a(s_261), .b(gate479inter3), .O(gate479inter10));
  nor2  gate2378(.a(gate479inter10), .b(gate479inter9), .O(gate479inter11));
  nor2  gate2379(.a(gate479inter11), .b(gate479inter6), .O(gate479inter12));
  nand2 gate2380(.a(gate479inter12), .b(gate479inter1), .O(G1288));
nand2 gate480( .a(G1126), .b(G1222), .O(G1289) );
nand2 gate481( .a(G32), .b(G1225), .O(G1290) );
nand2 gate482( .a(G1129), .b(G1225), .O(G1291) );

  xor2  gate2465(.a(G1229), .b(G1228), .O(gate483inter0));
  nand2 gate2466(.a(gate483inter0), .b(s_274), .O(gate483inter1));
  and2  gate2467(.a(G1229), .b(G1228), .O(gate483inter2));
  inv1  gate2468(.a(s_274), .O(gate483inter3));
  inv1  gate2469(.a(s_275), .O(gate483inter4));
  nand2 gate2470(.a(gate483inter4), .b(gate483inter3), .O(gate483inter5));
  nor2  gate2471(.a(gate483inter5), .b(gate483inter2), .O(gate483inter6));
  inv1  gate2472(.a(G1228), .O(gate483inter7));
  inv1  gate2473(.a(G1229), .O(gate483inter8));
  nand2 gate2474(.a(gate483inter8), .b(gate483inter7), .O(gate483inter9));
  nand2 gate2475(.a(s_275), .b(gate483inter3), .O(gate483inter10));
  nor2  gate2476(.a(gate483inter10), .b(gate483inter9), .O(gate483inter11));
  nor2  gate2477(.a(gate483inter11), .b(gate483inter6), .O(gate483inter12));
  nand2 gate2478(.a(gate483inter12), .b(gate483inter1), .O(G1292));
nand2 gate484( .a(G1230), .b(G1231), .O(G1293) );

  xor2  gate2409(.a(G1233), .b(G1232), .O(gate485inter0));
  nand2 gate2410(.a(gate485inter0), .b(s_266), .O(gate485inter1));
  and2  gate2411(.a(G1233), .b(G1232), .O(gate485inter2));
  inv1  gate2412(.a(s_266), .O(gate485inter3));
  inv1  gate2413(.a(s_267), .O(gate485inter4));
  nand2 gate2414(.a(gate485inter4), .b(gate485inter3), .O(gate485inter5));
  nor2  gate2415(.a(gate485inter5), .b(gate485inter2), .O(gate485inter6));
  inv1  gate2416(.a(G1232), .O(gate485inter7));
  inv1  gate2417(.a(G1233), .O(gate485inter8));
  nand2 gate2418(.a(gate485inter8), .b(gate485inter7), .O(gate485inter9));
  nand2 gate2419(.a(s_267), .b(gate485inter3), .O(gate485inter10));
  nor2  gate2420(.a(gate485inter10), .b(gate485inter9), .O(gate485inter11));
  nor2  gate2421(.a(gate485inter11), .b(gate485inter6), .O(gate485inter12));
  nand2 gate2422(.a(gate485inter12), .b(gate485inter1), .O(G1294));
nand2 gate486( .a(G1234), .b(G1235), .O(G1295) );

  xor2  gate1247(.a(G1237), .b(G1236), .O(gate487inter0));
  nand2 gate1248(.a(gate487inter0), .b(s_100), .O(gate487inter1));
  and2  gate1249(.a(G1237), .b(G1236), .O(gate487inter2));
  inv1  gate1250(.a(s_100), .O(gate487inter3));
  inv1  gate1251(.a(s_101), .O(gate487inter4));
  nand2 gate1252(.a(gate487inter4), .b(gate487inter3), .O(gate487inter5));
  nor2  gate1253(.a(gate487inter5), .b(gate487inter2), .O(gate487inter6));
  inv1  gate1254(.a(G1236), .O(gate487inter7));
  inv1  gate1255(.a(G1237), .O(gate487inter8));
  nand2 gate1256(.a(gate487inter8), .b(gate487inter7), .O(gate487inter9));
  nand2 gate1257(.a(s_101), .b(gate487inter3), .O(gate487inter10));
  nor2  gate1258(.a(gate487inter10), .b(gate487inter9), .O(gate487inter11));
  nor2  gate1259(.a(gate487inter11), .b(gate487inter6), .O(gate487inter12));
  nand2 gate1260(.a(gate487inter12), .b(gate487inter1), .O(G1296));
nand2 gate488( .a(G1238), .b(G1239), .O(G1297) );
nand2 gate489( .a(G1240), .b(G1241), .O(G1298) );

  xor2  gate757(.a(G1243), .b(G1242), .O(gate490inter0));
  nand2 gate758(.a(gate490inter0), .b(s_30), .O(gate490inter1));
  and2  gate759(.a(G1243), .b(G1242), .O(gate490inter2));
  inv1  gate760(.a(s_30), .O(gate490inter3));
  inv1  gate761(.a(s_31), .O(gate490inter4));
  nand2 gate762(.a(gate490inter4), .b(gate490inter3), .O(gate490inter5));
  nor2  gate763(.a(gate490inter5), .b(gate490inter2), .O(gate490inter6));
  inv1  gate764(.a(G1242), .O(gate490inter7));
  inv1  gate765(.a(G1243), .O(gate490inter8));
  nand2 gate766(.a(gate490inter8), .b(gate490inter7), .O(gate490inter9));
  nand2 gate767(.a(s_31), .b(gate490inter3), .O(gate490inter10));
  nor2  gate768(.a(gate490inter10), .b(gate490inter9), .O(gate490inter11));
  nor2  gate769(.a(gate490inter11), .b(gate490inter6), .O(gate490inter12));
  nand2 gate770(.a(gate490inter12), .b(gate490inter1), .O(G1299));
nand2 gate491( .a(G1244), .b(G1245), .O(G1300) );
nand2 gate492( .a(G1246), .b(G1247), .O(G1301) );
nand2 gate493( .a(G1248), .b(G1249), .O(G1302) );
nand2 gate494( .a(G1250), .b(G1251), .O(G1303) );
nand2 gate495( .a(G1252), .b(G1253), .O(G1304) );

  xor2  gate2675(.a(G1255), .b(G1254), .O(gate496inter0));
  nand2 gate2676(.a(gate496inter0), .b(s_304), .O(gate496inter1));
  and2  gate2677(.a(G1255), .b(G1254), .O(gate496inter2));
  inv1  gate2678(.a(s_304), .O(gate496inter3));
  inv1  gate2679(.a(s_305), .O(gate496inter4));
  nand2 gate2680(.a(gate496inter4), .b(gate496inter3), .O(gate496inter5));
  nor2  gate2681(.a(gate496inter5), .b(gate496inter2), .O(gate496inter6));
  inv1  gate2682(.a(G1254), .O(gate496inter7));
  inv1  gate2683(.a(G1255), .O(gate496inter8));
  nand2 gate2684(.a(gate496inter8), .b(gate496inter7), .O(gate496inter9));
  nand2 gate2685(.a(s_305), .b(gate496inter3), .O(gate496inter10));
  nor2  gate2686(.a(gate496inter10), .b(gate496inter9), .O(gate496inter11));
  nor2  gate2687(.a(gate496inter11), .b(gate496inter6), .O(gate496inter12));
  nand2 gate2688(.a(gate496inter12), .b(gate496inter1), .O(G1305));
nand2 gate497( .a(G1256), .b(G1257), .O(G1306) );
nand2 gate498( .a(G1258), .b(G1259), .O(G1307) );

  xor2  gate813(.a(G1261), .b(G1260), .O(gate499inter0));
  nand2 gate814(.a(gate499inter0), .b(s_38), .O(gate499inter1));
  and2  gate815(.a(G1261), .b(G1260), .O(gate499inter2));
  inv1  gate816(.a(s_38), .O(gate499inter3));
  inv1  gate817(.a(s_39), .O(gate499inter4));
  nand2 gate818(.a(gate499inter4), .b(gate499inter3), .O(gate499inter5));
  nor2  gate819(.a(gate499inter5), .b(gate499inter2), .O(gate499inter6));
  inv1  gate820(.a(G1260), .O(gate499inter7));
  inv1  gate821(.a(G1261), .O(gate499inter8));
  nand2 gate822(.a(gate499inter8), .b(gate499inter7), .O(gate499inter9));
  nand2 gate823(.a(s_39), .b(gate499inter3), .O(gate499inter10));
  nor2  gate824(.a(gate499inter10), .b(gate499inter9), .O(gate499inter11));
  nor2  gate825(.a(gate499inter11), .b(gate499inter6), .O(gate499inter12));
  nand2 gate826(.a(gate499inter12), .b(gate499inter1), .O(G1308));
nand2 gate500( .a(G1262), .b(G1263), .O(G1309) );
nand2 gate501( .a(G1264), .b(G1265), .O(G1310) );
nand2 gate502( .a(G1266), .b(G1267), .O(G1311) );

  xor2  gate575(.a(G1269), .b(G1268), .O(gate503inter0));
  nand2 gate576(.a(gate503inter0), .b(s_4), .O(gate503inter1));
  and2  gate577(.a(G1269), .b(G1268), .O(gate503inter2));
  inv1  gate578(.a(s_4), .O(gate503inter3));
  inv1  gate579(.a(s_5), .O(gate503inter4));
  nand2 gate580(.a(gate503inter4), .b(gate503inter3), .O(gate503inter5));
  nor2  gate581(.a(gate503inter5), .b(gate503inter2), .O(gate503inter6));
  inv1  gate582(.a(G1268), .O(gate503inter7));
  inv1  gate583(.a(G1269), .O(gate503inter8));
  nand2 gate584(.a(gate503inter8), .b(gate503inter7), .O(gate503inter9));
  nand2 gate585(.a(s_5), .b(gate503inter3), .O(gate503inter10));
  nor2  gate586(.a(gate503inter10), .b(gate503inter9), .O(gate503inter11));
  nor2  gate587(.a(gate503inter11), .b(gate503inter6), .O(gate503inter12));
  nand2 gate588(.a(gate503inter12), .b(gate503inter1), .O(G1312));
nand2 gate504( .a(G1270), .b(G1271), .O(G1313) );
nand2 gate505( .a(G1272), .b(G1273), .O(G1314) );
nand2 gate506( .a(G1274), .b(G1275), .O(G1315) );
nand2 gate507( .a(G1276), .b(G1277), .O(G1316) );
nand2 gate508( .a(G1278), .b(G1279), .O(G1317) );

  xor2  gate967(.a(G1281), .b(G1280), .O(gate509inter0));
  nand2 gate968(.a(gate509inter0), .b(s_60), .O(gate509inter1));
  and2  gate969(.a(G1281), .b(G1280), .O(gate509inter2));
  inv1  gate970(.a(s_60), .O(gate509inter3));
  inv1  gate971(.a(s_61), .O(gate509inter4));
  nand2 gate972(.a(gate509inter4), .b(gate509inter3), .O(gate509inter5));
  nor2  gate973(.a(gate509inter5), .b(gate509inter2), .O(gate509inter6));
  inv1  gate974(.a(G1280), .O(gate509inter7));
  inv1  gate975(.a(G1281), .O(gate509inter8));
  nand2 gate976(.a(gate509inter8), .b(gate509inter7), .O(gate509inter9));
  nand2 gate977(.a(s_61), .b(gate509inter3), .O(gate509inter10));
  nor2  gate978(.a(gate509inter10), .b(gate509inter9), .O(gate509inter11));
  nor2  gate979(.a(gate509inter11), .b(gate509inter6), .O(gate509inter12));
  nand2 gate980(.a(gate509inter12), .b(gate509inter1), .O(G1318));

  xor2  gate1079(.a(G1283), .b(G1282), .O(gate510inter0));
  nand2 gate1080(.a(gate510inter0), .b(s_76), .O(gate510inter1));
  and2  gate1081(.a(G1283), .b(G1282), .O(gate510inter2));
  inv1  gate1082(.a(s_76), .O(gate510inter3));
  inv1  gate1083(.a(s_77), .O(gate510inter4));
  nand2 gate1084(.a(gate510inter4), .b(gate510inter3), .O(gate510inter5));
  nor2  gate1085(.a(gate510inter5), .b(gate510inter2), .O(gate510inter6));
  inv1  gate1086(.a(G1282), .O(gate510inter7));
  inv1  gate1087(.a(G1283), .O(gate510inter8));
  nand2 gate1088(.a(gate510inter8), .b(gate510inter7), .O(gate510inter9));
  nand2 gate1089(.a(s_77), .b(gate510inter3), .O(gate510inter10));
  nor2  gate1090(.a(gate510inter10), .b(gate510inter9), .O(gate510inter11));
  nor2  gate1091(.a(gate510inter11), .b(gate510inter6), .O(gate510inter12));
  nand2 gate1092(.a(gate510inter12), .b(gate510inter1), .O(G1319));

  xor2  gate1261(.a(G1285), .b(G1284), .O(gate511inter0));
  nand2 gate1262(.a(gate511inter0), .b(s_102), .O(gate511inter1));
  and2  gate1263(.a(G1285), .b(G1284), .O(gate511inter2));
  inv1  gate1264(.a(s_102), .O(gate511inter3));
  inv1  gate1265(.a(s_103), .O(gate511inter4));
  nand2 gate1266(.a(gate511inter4), .b(gate511inter3), .O(gate511inter5));
  nor2  gate1267(.a(gate511inter5), .b(gate511inter2), .O(gate511inter6));
  inv1  gate1268(.a(G1284), .O(gate511inter7));
  inv1  gate1269(.a(G1285), .O(gate511inter8));
  nand2 gate1270(.a(gate511inter8), .b(gate511inter7), .O(gate511inter9));
  nand2 gate1271(.a(s_103), .b(gate511inter3), .O(gate511inter10));
  nor2  gate1272(.a(gate511inter10), .b(gate511inter9), .O(gate511inter11));
  nor2  gate1273(.a(gate511inter11), .b(gate511inter6), .O(gate511inter12));
  nand2 gate1274(.a(gate511inter12), .b(gate511inter1), .O(G1320));
nand2 gate512( .a(G1286), .b(G1287), .O(G1321) );
nand2 gate513( .a(G1288), .b(G1289), .O(G1322) );
nand2 gate514( .a(G1290), .b(G1291), .O(G1323) );
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule