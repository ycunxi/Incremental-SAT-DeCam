module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);

input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;//RE__PI;

input s_0,s_1;//RE__ALLOW(00,01,10,11);
input s_2,s_3;//RE__ALLOW(00,01,10,11);
input s_4,s_5;//RE__ALLOW(00,01,10,11);
input s_6,s_7;//RE__ALLOW(00,01,10,11);
input s_8,s_9;//RE__ALLOW(00,01,10,11);
input s_10,s_11;//RE__ALLOW(00,01,10,11);
input s_12,s_13;//RE__ALLOW(00,01,10,11);
input s_14,s_15;//RE__ALLOW(00,01,10,11);
input s_16,s_17;//RE__ALLOW(00,01,10,11);
input s_18,s_19;//RE__ALLOW(00,01,10,11);
input s_20,s_21;//RE__ALLOW(00,01,10,11);
input s_22,s_23;//RE__ALLOW(00,01,10,11);
input s_24,s_25;//RE__ALLOW(00,01,10,11);
input s_26,s_27;//RE__ALLOW(00,01,10,11);
input s_28,s_29;//RE__ALLOW(00,01,10,11);
input s_30,s_31;//RE__ALLOW(00,01,10,11);
input s_32,s_33;//RE__ALLOW(00,01,10,11);
input s_34,s_35;//RE__ALLOW(00,01,10,11);
input s_36,s_37;//RE__ALLOW(00,01,10,11);
input s_38,s_39;//RE__ALLOW(00,01,10,11);
input s_40,s_41;//RE__ALLOW(00,01,10,11);
input s_42,s_43;//RE__ALLOW(00,01,10,11);
input s_44,s_45;//RE__ALLOW(00,01,10,11);
input s_46,s_47;//RE__ALLOW(00,01,10,11);
input s_48,s_49;//RE__ALLOW(00,01,10,11);
input s_50,s_51;//RE__ALLOW(00,01,10,11);
input s_52,s_53;//RE__ALLOW(00,01,10,11);
input s_54,s_55;//RE__ALLOW(00,01,10,11);
input s_56,s_57;//RE__ALLOW(00,01,10,11);
input s_58,s_59;//RE__ALLOW(00,01,10,11);
input s_60,s_61;//RE__ALLOW(00,01,10,11);
input s_62,s_63;//RE__ALLOW(00,01,10,11);
input s_64,s_65;//RE__ALLOW(00,01,10,11);
input s_66,s_67;//RE__ALLOW(00,01,10,11);
input s_68,s_69;//RE__ALLOW(00,01,10,11);
input s_70,s_71;//RE__ALLOW(00,01,10,11);
input s_72,s_73;//RE__ALLOW(00,01,10,11);
input s_74,s_75;//RE__ALLOW(00,01,10,11);
input s_76,s_77;//RE__ALLOW(00,01,10,11);
input s_78,s_79;//RE__ALLOW(00,01,10,11);
input s_80,s_81;//RE__ALLOW(00,01,10,11);
input s_82,s_83;//RE__ALLOW(00,01,10,11);
input s_84,s_85;//RE__ALLOW(00,01,10,11);
input s_86,s_87;//RE__ALLOW(00,01,10,11);
input s_88,s_89;//RE__ALLOW(00,01,10,11);
input s_90,s_91;//RE__ALLOW(00,01,10,11);
input s_92,s_93;//RE__ALLOW(00,01,10,11);
input s_94,s_95;//RE__ALLOW(00,01,10,11);
input s_96,s_97;//RE__ALLOW(00,01,10,11);
input s_98,s_99;//RE__ALLOW(00,01,10,11);
input s_100,s_101;//RE__ALLOW(00,01,10,11);
input s_102,s_103;//RE__ALLOW(00,01,10,11);
input s_104,s_105;//RE__ALLOW(00,01,10,11);
input s_106,s_107;//RE__ALLOW(00,01,10,11);
input s_108,s_109;//RE__ALLOW(00,01,10,11);
input s_110,s_111;//RE__ALLOW(00,01,10,11);
input s_112,s_113;//RE__ALLOW(00,01,10,11);
input s_114,s_115;//RE__ALLOW(00,01,10,11);
input s_116,s_117;//RE__ALLOW(00,01,10,11);
input s_118,s_119;//RE__ALLOW(00,01,10,11);
input s_120,s_121;//RE__ALLOW(00,01,10,11);
input s_122,s_123;//RE__ALLOW(00,01,10,11);
input s_124,s_125;//RE__ALLOW(00,01,10,11);
input s_126,s_127;//RE__ALLOW(00,01,10,11);
input s_128,s_129;//RE__ALLOW(00,01,10,11);
input s_130,s_131;//RE__ALLOW(00,01,10,11);
input s_132,s_133;//RE__ALLOW(00,01,10,11);
input s_134,s_135;//RE__ALLOW(00,01,10,11);
input s_136,s_137;//RE__ALLOW(00,01,10,11);
input s_138,s_139;//RE__ALLOW(00,01,10,11);
input s_140,s_141;//RE__ALLOW(00,01,10,11);
input s_142,s_143;//RE__ALLOW(00,01,10,11);
input s_144,s_145;//RE__ALLOW(00,01,10,11);
input s_146,s_147;//RE__ALLOW(00,01,10,11);
input s_148,s_149;//RE__ALLOW(00,01,10,11);
input s_150,s_151;//RE__ALLOW(00,01,10,11);
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;

  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate48inter0, gate48inter1, gate48inter2, gate48inter3, gate48inter4, gate48inter5, gate48inter6, gate48inter7, gate48inter8, gate48inter9, gate48inter10, gate48inter11, gate48inter12, gate464inter0, gate464inter1, gate464inter2, gate464inter3, gate464inter4, gate464inter5, gate464inter6, gate464inter7, gate464inter8, gate464inter9, gate464inter10, gate464inter11, gate464inter12, gate436inter0, gate436inter1, gate436inter2, gate436inter3, gate436inter4, gate436inter5, gate436inter6, gate436inter7, gate436inter8, gate436inter9, gate436inter10, gate436inter11, gate436inter12, gate142inter0, gate142inter1, gate142inter2, gate142inter3, gate142inter4, gate142inter5, gate142inter6, gate142inter7, gate142inter8, gate142inter9, gate142inter10, gate142inter11, gate142inter12, gate36inter0, gate36inter1, gate36inter2, gate36inter3, gate36inter4, gate36inter5, gate36inter6, gate36inter7, gate36inter8, gate36inter9, gate36inter10, gate36inter11, gate36inter12, gate157inter0, gate157inter1, gate157inter2, gate157inter3, gate157inter4, gate157inter5, gate157inter6, gate157inter7, gate157inter8, gate157inter9, gate157inter10, gate157inter11, gate157inter12, gate467inter0, gate467inter1, gate467inter2, gate467inter3, gate467inter4, gate467inter5, gate467inter6, gate467inter7, gate467inter8, gate467inter9, gate467inter10, gate467inter11, gate467inter12, gate223inter0, gate223inter1, gate223inter2, gate223inter3, gate223inter4, gate223inter5, gate223inter6, gate223inter7, gate223inter8, gate223inter9, gate223inter10, gate223inter11, gate223inter12, gate462inter0, gate462inter1, gate462inter2, gate462inter3, gate462inter4, gate462inter5, gate462inter6, gate462inter7, gate462inter8, gate462inter9, gate462inter10, gate462inter11, gate462inter12, gate476inter0, gate476inter1, gate476inter2, gate476inter3, gate476inter4, gate476inter5, gate476inter6, gate476inter7, gate476inter8, gate476inter9, gate476inter10, gate476inter11, gate476inter12, gate459inter0, gate459inter1, gate459inter2, gate459inter3, gate459inter4, gate459inter5, gate459inter6, gate459inter7, gate459inter8, gate459inter9, gate459inter10, gate459inter11, gate459inter12, gate433inter0, gate433inter1, gate433inter2, gate433inter3, gate433inter4, gate433inter5, gate433inter6, gate433inter7, gate433inter8, gate433inter9, gate433inter10, gate433inter11, gate433inter12, gate212inter0, gate212inter1, gate212inter2, gate212inter3, gate212inter4, gate212inter5, gate212inter6, gate212inter7, gate212inter8, gate212inter9, gate212inter10, gate212inter11, gate212inter12, gate276inter0, gate276inter1, gate276inter2, gate276inter3, gate276inter4, gate276inter5, gate276inter6, gate276inter7, gate276inter8, gate276inter9, gate276inter10, gate276inter11, gate276inter12, gate135inter0, gate135inter1, gate135inter2, gate135inter3, gate135inter4, gate135inter5, gate135inter6, gate135inter7, gate135inter8, gate135inter9, gate135inter10, gate135inter11, gate135inter12, gate284inter0, gate284inter1, gate284inter2, gate284inter3, gate284inter4, gate284inter5, gate284inter6, gate284inter7, gate284inter8, gate284inter9, gate284inter10, gate284inter11, gate284inter12, gate163inter0, gate163inter1, gate163inter2, gate163inter3, gate163inter4, gate163inter5, gate163inter6, gate163inter7, gate163inter8, gate163inter9, gate163inter10, gate163inter11, gate163inter12, gate58inter0, gate58inter1, gate58inter2, gate58inter3, gate58inter4, gate58inter5, gate58inter6, gate58inter7, gate58inter8, gate58inter9, gate58inter10, gate58inter11, gate58inter12, gate292inter0, gate292inter1, gate292inter2, gate292inter3, gate292inter4, gate292inter5, gate292inter6, gate292inter7, gate292inter8, gate292inter9, gate292inter10, gate292inter11, gate292inter12, gate31inter0, gate31inter1, gate31inter2, gate31inter3, gate31inter4, gate31inter5, gate31inter6, gate31inter7, gate31inter8, gate31inter9, gate31inter10, gate31inter11, gate31inter12, gate24inter0, gate24inter1, gate24inter2, gate24inter3, gate24inter4, gate24inter5, gate24inter6, gate24inter7, gate24inter8, gate24inter9, gate24inter10, gate24inter11, gate24inter12, gate508inter0, gate508inter1, gate508inter2, gate508inter3, gate508inter4, gate508inter5, gate508inter6, gate508inter7, gate508inter8, gate508inter9, gate508inter10, gate508inter11, gate508inter12, gate39inter0, gate39inter1, gate39inter2, gate39inter3, gate39inter4, gate39inter5, gate39inter6, gate39inter7, gate39inter8, gate39inter9, gate39inter10, gate39inter11, gate39inter12, gate274inter0, gate274inter1, gate274inter2, gate274inter3, gate274inter4, gate274inter5, gate274inter6, gate274inter7, gate274inter8, gate274inter9, gate274inter10, gate274inter11, gate274inter12, gate164inter0, gate164inter1, gate164inter2, gate164inter3, gate164inter4, gate164inter5, gate164inter6, gate164inter7, gate164inter8, gate164inter9, gate164inter10, gate164inter11, gate164inter12, gate435inter0, gate435inter1, gate435inter2, gate435inter3, gate435inter4, gate435inter5, gate435inter6, gate435inter7, gate435inter8, gate435inter9, gate435inter10, gate435inter11, gate435inter12, gate458inter0, gate458inter1, gate458inter2, gate458inter3, gate458inter4, gate458inter5, gate458inter6, gate458inter7, gate458inter8, gate458inter9, gate458inter10, gate458inter11, gate458inter12, gate188inter0, gate188inter1, gate188inter2, gate188inter3, gate188inter4, gate188inter5, gate188inter6, gate188inter7, gate188inter8, gate188inter9, gate188inter10, gate188inter11, gate188inter12, gate181inter0, gate181inter1, gate181inter2, gate181inter3, gate181inter4, gate181inter5, gate181inter6, gate181inter7, gate181inter8, gate181inter9, gate181inter10, gate181inter11, gate181inter12, gate451inter0, gate451inter1, gate451inter2, gate451inter3, gate451inter4, gate451inter5, gate451inter6, gate451inter7, gate451inter8, gate451inter9, gate451inter10, gate451inter11, gate451inter12, gate118inter0, gate118inter1, gate118inter2, gate118inter3, gate118inter4, gate118inter5, gate118inter6, gate118inter7, gate118inter8, gate118inter9, gate118inter10, gate118inter11, gate118inter12, gate217inter0, gate217inter1, gate217inter2, gate217inter3, gate217inter4, gate217inter5, gate217inter6, gate217inter7, gate217inter8, gate217inter9, gate217inter10, gate217inter11, gate217inter12, gate294inter0, gate294inter1, gate294inter2, gate294inter3, gate294inter4, gate294inter5, gate294inter6, gate294inter7, gate294inter8, gate294inter9, gate294inter10, gate294inter11, gate294inter12, gate393inter0, gate393inter1, gate393inter2, gate393inter3, gate393inter4, gate393inter5, gate393inter6, gate393inter7, gate393inter8, gate393inter9, gate393inter10, gate393inter11, gate393inter12, gate199inter0, gate199inter1, gate199inter2, gate199inter3, gate199inter4, gate199inter5, gate199inter6, gate199inter7, gate199inter8, gate199inter9, gate199inter10, gate199inter11, gate199inter12, gate111inter0, gate111inter1, gate111inter2, gate111inter3, gate111inter4, gate111inter5, gate111inter6, gate111inter7, gate111inter8, gate111inter9, gate111inter10, gate111inter11, gate111inter12, gate100inter0, gate100inter1, gate100inter2, gate100inter3, gate100inter4, gate100inter5, gate100inter6, gate100inter7, gate100inter8, gate100inter9, gate100inter10, gate100inter11, gate100inter12, gate510inter0, gate510inter1, gate510inter2, gate510inter3, gate510inter4, gate510inter5, gate510inter6, gate510inter7, gate510inter8, gate510inter9, gate510inter10, gate510inter11, gate510inter12, gate457inter0, gate457inter1, gate457inter2, gate457inter3, gate457inter4, gate457inter5, gate457inter6, gate457inter7, gate457inter8, gate457inter9, gate457inter10, gate457inter11, gate457inter12, gate441inter0, gate441inter1, gate441inter2, gate441inter3, gate441inter4, gate441inter5, gate441inter6, gate441inter7, gate441inter8, gate441inter9, gate441inter10, gate441inter11, gate441inter12, gate117inter0, gate117inter1, gate117inter2, gate117inter3, gate117inter4, gate117inter5, gate117inter6, gate117inter7, gate117inter8, gate117inter9, gate117inter10, gate117inter11, gate117inter12, gate469inter0, gate469inter1, gate469inter2, gate469inter3, gate469inter4, gate469inter5, gate469inter6, gate469inter7, gate469inter8, gate469inter9, gate469inter10, gate469inter11, gate469inter12, gate34inter0, gate34inter1, gate34inter2, gate34inter3, gate34inter4, gate34inter5, gate34inter6, gate34inter7, gate34inter8, gate34inter9, gate34inter10, gate34inter11, gate34inter12, gate173inter0, gate173inter1, gate173inter2, gate173inter3, gate173inter4, gate173inter5, gate173inter6, gate173inter7, gate173inter8, gate173inter9, gate173inter10, gate173inter11, gate173inter12, gate20inter0, gate20inter1, gate20inter2, gate20inter3, gate20inter4, gate20inter5, gate20inter6, gate20inter7, gate20inter8, gate20inter9, gate20inter10, gate20inter11, gate20inter12, gate291inter0, gate291inter1, gate291inter2, gate291inter3, gate291inter4, gate291inter5, gate291inter6, gate291inter7, gate291inter8, gate291inter9, gate291inter10, gate291inter11, gate291inter12, gate23inter0, gate23inter1, gate23inter2, gate23inter3, gate23inter4, gate23inter5, gate23inter6, gate23inter7, gate23inter8, gate23inter9, gate23inter10, gate23inter11, gate23inter12, gate89inter0, gate89inter1, gate89inter2, gate89inter3, gate89inter4, gate89inter5, gate89inter6, gate89inter7, gate89inter8, gate89inter9, gate89inter10, gate89inter11, gate89inter12, gate506inter0, gate506inter1, gate506inter2, gate506inter3, gate506inter4, gate506inter5, gate506inter6, gate506inter7, gate506inter8, gate506inter9, gate506inter10, gate506inter11, gate506inter12, gate94inter0, gate94inter1, gate94inter2, gate94inter3, gate94inter4, gate94inter5, gate94inter6, gate94inter7, gate94inter8, gate94inter9, gate94inter10, gate94inter11, gate94inter12, gate147inter0, gate147inter1, gate147inter2, gate147inter3, gate147inter4, gate147inter5, gate147inter6, gate147inter7, gate147inter8, gate147inter9, gate147inter10, gate147inter11, gate147inter12, gate460inter0, gate460inter1, gate460inter2, gate460inter3, gate460inter4, gate460inter5, gate460inter6, gate460inter7, gate460inter8, gate460inter9, gate460inter10, gate460inter11, gate460inter12, gate439inter0, gate439inter1, gate439inter2, gate439inter3, gate439inter4, gate439inter5, gate439inter6, gate439inter7, gate439inter8, gate439inter9, gate439inter10, gate439inter11, gate439inter12, gate152inter0, gate152inter1, gate152inter2, gate152inter3, gate152inter4, gate152inter5, gate152inter6, gate152inter7, gate152inter8, gate152inter9, gate152inter10, gate152inter11, gate152inter12, gate423inter0, gate423inter1, gate423inter2, gate423inter3, gate423inter4, gate423inter5, gate423inter6, gate423inter7, gate423inter8, gate423inter9, gate423inter10, gate423inter11, gate423inter12, gate51inter0, gate51inter1, gate51inter2, gate51inter3, gate51inter4, gate51inter5, gate51inter6, gate51inter7, gate51inter8, gate51inter9, gate51inter10, gate51inter11, gate51inter12, gate44inter0, gate44inter1, gate44inter2, gate44inter3, gate44inter4, gate44inter5, gate44inter6, gate44inter7, gate44inter8, gate44inter9, gate44inter10, gate44inter11, gate44inter12, gate93inter0, gate93inter1, gate93inter2, gate93inter3, gate93inter4, gate93inter5, gate93inter6, gate93inter7, gate93inter8, gate93inter9, gate93inter10, gate93inter11, gate93inter12, gate501inter0, gate501inter1, gate501inter2, gate501inter3, gate501inter4, gate501inter5, gate501inter6, gate501inter7, gate501inter8, gate501inter9, gate501inter10, gate501inter11, gate501inter12, gate86inter0, gate86inter1, gate86inter2, gate86inter3, gate86inter4, gate86inter5, gate86inter6, gate86inter7, gate86inter8, gate86inter9, gate86inter10, gate86inter11, gate86inter12, gate66inter0, gate66inter1, gate66inter2, gate66inter3, gate66inter4, gate66inter5, gate66inter6, gate66inter7, gate66inter8, gate66inter9, gate66inter10, gate66inter11, gate66inter12, gate22inter0, gate22inter1, gate22inter2, gate22inter3, gate22inter4, gate22inter5, gate22inter6, gate22inter7, gate22inter8, gate22inter9, gate22inter10, gate22inter11, gate22inter12, gate448inter0, gate448inter1, gate448inter2, gate448inter3, gate448inter4, gate448inter5, gate448inter6, gate448inter7, gate448inter8, gate448inter9, gate448inter10, gate448inter11, gate448inter12, gate182inter0, gate182inter1, gate182inter2, gate182inter3, gate182inter4, gate182inter5, gate182inter6, gate182inter7, gate182inter8, gate182inter9, gate182inter10, gate182inter11, gate182inter12, gate397inter0, gate397inter1, gate397inter2, gate397inter3, gate397inter4, gate397inter5, gate397inter6, gate397inter7, gate397inter8, gate397inter9, gate397inter10, gate397inter11, gate397inter12, gate180inter0, gate180inter1, gate180inter2, gate180inter3, gate180inter4, gate180inter5, gate180inter6, gate180inter7, gate180inter8, gate180inter9, gate180inter10, gate180inter11, gate180inter12, gate17inter0, gate17inter1, gate17inter2, gate17inter3, gate17inter4, gate17inter5, gate17inter6, gate17inter7, gate17inter8, gate17inter9, gate17inter10, gate17inter11, gate17inter12, gate161inter0, gate161inter1, gate161inter2, gate161inter3, gate161inter4, gate161inter5, gate161inter6, gate161inter7, gate161inter8, gate161inter9, gate161inter10, gate161inter11, gate161inter12, gate148inter0, gate148inter1, gate148inter2, gate148inter3, gate148inter4, gate148inter5, gate148inter6, gate148inter7, gate148inter8, gate148inter9, gate148inter10, gate148inter11, gate148inter12, gate103inter0, gate103inter1, gate103inter2, gate103inter3, gate103inter4, gate103inter5, gate103inter6, gate103inter7, gate103inter8, gate103inter9, gate103inter10, gate103inter11, gate103inter12, gate285inter0, gate285inter1, gate285inter2, gate285inter3, gate285inter4, gate285inter5, gate285inter6, gate285inter7, gate285inter8, gate285inter9, gate285inter10, gate285inter11, gate285inter12, gate119inter0, gate119inter1, gate119inter2, gate119inter3, gate119inter4, gate119inter5, gate119inter6, gate119inter7, gate119inter8, gate119inter9, gate119inter10, gate119inter11, gate119inter12, gate29inter0, gate29inter1, gate29inter2, gate29inter3, gate29inter4, gate29inter5, gate29inter6, gate29inter7, gate29inter8, gate29inter9, gate29inter10, gate29inter11, gate29inter12, gate232inter0, gate232inter1, gate232inter2, gate232inter3, gate232inter4, gate232inter5, gate232inter6, gate232inter7, gate232inter8, gate232inter9, gate232inter10, gate232inter11, gate232inter12, gate184inter0, gate184inter1, gate184inter2, gate184inter3, gate184inter4, gate184inter5, gate184inter6, gate184inter7, gate184inter8, gate184inter9, gate184inter10, gate184inter11, gate184inter12, gate130inter0, gate130inter1, gate130inter2, gate130inter3, gate130inter4, gate130inter5, gate130inter6, gate130inter7, gate130inter8, gate130inter9, gate130inter10, gate130inter11, gate130inter12;



and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );
nand2 gate9( .a(G1), .b(G2), .O(G266) );
nand2 gate10( .a(G3), .b(G4), .O(G269) );
nand2 gate11( .a(G5), .b(G6), .O(G272) );
nand2 gate12( .a(G7), .b(G8), .O(G275) );
nand2 gate13( .a(G9), .b(G10), .O(G278) );
nand2 gate14( .a(G11), .b(G12), .O(G281) );
nand2 gate15( .a(G13), .b(G14), .O(G284) );
nand2 gate16( .a(G15), .b(G16), .O(G287) );

  xor2  gate1471(.a(G18), .b(G17), .O(gate17inter0));
  nand2 gate1472(.a(gate17inter0), .b(s_132), .O(gate17inter1));
  and2  gate1473(.a(G18), .b(G17), .O(gate17inter2));
  inv1  gate1474(.a(s_132), .O(gate17inter3));
  inv1  gate1475(.a(s_133), .O(gate17inter4));
  nand2 gate1476(.a(gate17inter4), .b(gate17inter3), .O(gate17inter5));
  nor2  gate1477(.a(gate17inter5), .b(gate17inter2), .O(gate17inter6));
  inv1  gate1478(.a(G17), .O(gate17inter7));
  inv1  gate1479(.a(G18), .O(gate17inter8));
  nand2 gate1480(.a(gate17inter8), .b(gate17inter7), .O(gate17inter9));
  nand2 gate1481(.a(s_133), .b(gate17inter3), .O(gate17inter10));
  nor2  gate1482(.a(gate17inter10), .b(gate17inter9), .O(gate17inter11));
  nor2  gate1483(.a(gate17inter11), .b(gate17inter6), .O(gate17inter12));
  nand2 gate1484(.a(gate17inter12), .b(gate17inter1), .O(G290));
nand2 gate18( .a(G19), .b(G20), .O(G293) );
nand2 gate19( .a(G21), .b(G22), .O(G296) );

  xor2  gate1163(.a(G24), .b(G23), .O(gate20inter0));
  nand2 gate1164(.a(gate20inter0), .b(s_88), .O(gate20inter1));
  and2  gate1165(.a(G24), .b(G23), .O(gate20inter2));
  inv1  gate1166(.a(s_88), .O(gate20inter3));
  inv1  gate1167(.a(s_89), .O(gate20inter4));
  nand2 gate1168(.a(gate20inter4), .b(gate20inter3), .O(gate20inter5));
  nor2  gate1169(.a(gate20inter5), .b(gate20inter2), .O(gate20inter6));
  inv1  gate1170(.a(G23), .O(gate20inter7));
  inv1  gate1171(.a(G24), .O(gate20inter8));
  nand2 gate1172(.a(gate20inter8), .b(gate20inter7), .O(gate20inter9));
  nand2 gate1173(.a(s_89), .b(gate20inter3), .O(gate20inter10));
  nor2  gate1174(.a(gate20inter10), .b(gate20inter9), .O(gate20inter11));
  nor2  gate1175(.a(gate20inter11), .b(gate20inter6), .O(gate20inter12));
  nand2 gate1176(.a(gate20inter12), .b(gate20inter1), .O(G299));
nand2 gate21( .a(G25), .b(G26), .O(G302) );

  xor2  gate1401(.a(G28), .b(G27), .O(gate22inter0));
  nand2 gate1402(.a(gate22inter0), .b(s_122), .O(gate22inter1));
  and2  gate1403(.a(G28), .b(G27), .O(gate22inter2));
  inv1  gate1404(.a(s_122), .O(gate22inter3));
  inv1  gate1405(.a(s_123), .O(gate22inter4));
  nand2 gate1406(.a(gate22inter4), .b(gate22inter3), .O(gate22inter5));
  nor2  gate1407(.a(gate22inter5), .b(gate22inter2), .O(gate22inter6));
  inv1  gate1408(.a(G27), .O(gate22inter7));
  inv1  gate1409(.a(G28), .O(gate22inter8));
  nand2 gate1410(.a(gate22inter8), .b(gate22inter7), .O(gate22inter9));
  nand2 gate1411(.a(s_123), .b(gate22inter3), .O(gate22inter10));
  nor2  gate1412(.a(gate22inter10), .b(gate22inter9), .O(gate22inter11));
  nor2  gate1413(.a(gate22inter11), .b(gate22inter6), .O(gate22inter12));
  nand2 gate1414(.a(gate22inter12), .b(gate22inter1), .O(G305));

  xor2  gate1191(.a(G30), .b(G29), .O(gate23inter0));
  nand2 gate1192(.a(gate23inter0), .b(s_92), .O(gate23inter1));
  and2  gate1193(.a(G30), .b(G29), .O(gate23inter2));
  inv1  gate1194(.a(s_92), .O(gate23inter3));
  inv1  gate1195(.a(s_93), .O(gate23inter4));
  nand2 gate1196(.a(gate23inter4), .b(gate23inter3), .O(gate23inter5));
  nor2  gate1197(.a(gate23inter5), .b(gate23inter2), .O(gate23inter6));
  inv1  gate1198(.a(G29), .O(gate23inter7));
  inv1  gate1199(.a(G30), .O(gate23inter8));
  nand2 gate1200(.a(gate23inter8), .b(gate23inter7), .O(gate23inter9));
  nand2 gate1201(.a(s_93), .b(gate23inter3), .O(gate23inter10));
  nor2  gate1202(.a(gate23inter10), .b(gate23inter9), .O(gate23inter11));
  nor2  gate1203(.a(gate23inter11), .b(gate23inter6), .O(gate23inter12));
  nand2 gate1204(.a(gate23inter12), .b(gate23inter1), .O(G308));

  xor2  gate827(.a(G32), .b(G31), .O(gate24inter0));
  nand2 gate828(.a(gate24inter0), .b(s_40), .O(gate24inter1));
  and2  gate829(.a(G32), .b(G31), .O(gate24inter2));
  inv1  gate830(.a(s_40), .O(gate24inter3));
  inv1  gate831(.a(s_41), .O(gate24inter4));
  nand2 gate832(.a(gate24inter4), .b(gate24inter3), .O(gate24inter5));
  nor2  gate833(.a(gate24inter5), .b(gate24inter2), .O(gate24inter6));
  inv1  gate834(.a(G31), .O(gate24inter7));
  inv1  gate835(.a(G32), .O(gate24inter8));
  nand2 gate836(.a(gate24inter8), .b(gate24inter7), .O(gate24inter9));
  nand2 gate837(.a(s_41), .b(gate24inter3), .O(gate24inter10));
  nor2  gate838(.a(gate24inter10), .b(gate24inter9), .O(gate24inter11));
  nor2  gate839(.a(gate24inter11), .b(gate24inter6), .O(gate24inter12));
  nand2 gate840(.a(gate24inter12), .b(gate24inter1), .O(G311));
nand2 gate25( .a(G1), .b(G5), .O(G314) );
nand2 gate26( .a(G9), .b(G13), .O(G317) );
nand2 gate27( .a(G2), .b(G6), .O(G320) );
nand2 gate28( .a(G10), .b(G14), .O(G323) );

  xor2  gate1555(.a(G7), .b(G3), .O(gate29inter0));
  nand2 gate1556(.a(gate29inter0), .b(s_144), .O(gate29inter1));
  and2  gate1557(.a(G7), .b(G3), .O(gate29inter2));
  inv1  gate1558(.a(s_144), .O(gate29inter3));
  inv1  gate1559(.a(s_145), .O(gate29inter4));
  nand2 gate1560(.a(gate29inter4), .b(gate29inter3), .O(gate29inter5));
  nor2  gate1561(.a(gate29inter5), .b(gate29inter2), .O(gate29inter6));
  inv1  gate1562(.a(G3), .O(gate29inter7));
  inv1  gate1563(.a(G7), .O(gate29inter8));
  nand2 gate1564(.a(gate29inter8), .b(gate29inter7), .O(gate29inter9));
  nand2 gate1565(.a(s_145), .b(gate29inter3), .O(gate29inter10));
  nor2  gate1566(.a(gate29inter10), .b(gate29inter9), .O(gate29inter11));
  nor2  gate1567(.a(gate29inter11), .b(gate29inter6), .O(gate29inter12));
  nand2 gate1568(.a(gate29inter12), .b(gate29inter1), .O(G326));
nand2 gate30( .a(G11), .b(G15), .O(G329) );

  xor2  gate813(.a(G8), .b(G4), .O(gate31inter0));
  nand2 gate814(.a(gate31inter0), .b(s_38), .O(gate31inter1));
  and2  gate815(.a(G8), .b(G4), .O(gate31inter2));
  inv1  gate816(.a(s_38), .O(gate31inter3));
  inv1  gate817(.a(s_39), .O(gate31inter4));
  nand2 gate818(.a(gate31inter4), .b(gate31inter3), .O(gate31inter5));
  nor2  gate819(.a(gate31inter5), .b(gate31inter2), .O(gate31inter6));
  inv1  gate820(.a(G4), .O(gate31inter7));
  inv1  gate821(.a(G8), .O(gate31inter8));
  nand2 gate822(.a(gate31inter8), .b(gate31inter7), .O(gate31inter9));
  nand2 gate823(.a(s_39), .b(gate31inter3), .O(gate31inter10));
  nor2  gate824(.a(gate31inter10), .b(gate31inter9), .O(gate31inter11));
  nor2  gate825(.a(gate31inter11), .b(gate31inter6), .O(gate31inter12));
  nand2 gate826(.a(gate31inter12), .b(gate31inter1), .O(G332));
nand2 gate32( .a(G12), .b(G16), .O(G335) );
nand2 gate33( .a(G17), .b(G21), .O(G338) );

  xor2  gate1135(.a(G29), .b(G25), .O(gate34inter0));
  nand2 gate1136(.a(gate34inter0), .b(s_84), .O(gate34inter1));
  and2  gate1137(.a(G29), .b(G25), .O(gate34inter2));
  inv1  gate1138(.a(s_84), .O(gate34inter3));
  inv1  gate1139(.a(s_85), .O(gate34inter4));
  nand2 gate1140(.a(gate34inter4), .b(gate34inter3), .O(gate34inter5));
  nor2  gate1141(.a(gate34inter5), .b(gate34inter2), .O(gate34inter6));
  inv1  gate1142(.a(G25), .O(gate34inter7));
  inv1  gate1143(.a(G29), .O(gate34inter8));
  nand2 gate1144(.a(gate34inter8), .b(gate34inter7), .O(gate34inter9));
  nand2 gate1145(.a(s_85), .b(gate34inter3), .O(gate34inter10));
  nor2  gate1146(.a(gate34inter10), .b(gate34inter9), .O(gate34inter11));
  nor2  gate1147(.a(gate34inter11), .b(gate34inter6), .O(gate34inter12));
  nand2 gate1148(.a(gate34inter12), .b(gate34inter1), .O(G341));
nand2 gate35( .a(G18), .b(G22), .O(G344) );

  xor2  gate603(.a(G30), .b(G26), .O(gate36inter0));
  nand2 gate604(.a(gate36inter0), .b(s_8), .O(gate36inter1));
  and2  gate605(.a(G30), .b(G26), .O(gate36inter2));
  inv1  gate606(.a(s_8), .O(gate36inter3));
  inv1  gate607(.a(s_9), .O(gate36inter4));
  nand2 gate608(.a(gate36inter4), .b(gate36inter3), .O(gate36inter5));
  nor2  gate609(.a(gate36inter5), .b(gate36inter2), .O(gate36inter6));
  inv1  gate610(.a(G26), .O(gate36inter7));
  inv1  gate611(.a(G30), .O(gate36inter8));
  nand2 gate612(.a(gate36inter8), .b(gate36inter7), .O(gate36inter9));
  nand2 gate613(.a(s_9), .b(gate36inter3), .O(gate36inter10));
  nor2  gate614(.a(gate36inter10), .b(gate36inter9), .O(gate36inter11));
  nor2  gate615(.a(gate36inter11), .b(gate36inter6), .O(gate36inter12));
  nand2 gate616(.a(gate36inter12), .b(gate36inter1), .O(G347));
nand2 gate37( .a(G19), .b(G23), .O(G350) );
nand2 gate38( .a(G27), .b(G31), .O(G353) );

  xor2  gate855(.a(G24), .b(G20), .O(gate39inter0));
  nand2 gate856(.a(gate39inter0), .b(s_44), .O(gate39inter1));
  and2  gate857(.a(G24), .b(G20), .O(gate39inter2));
  inv1  gate858(.a(s_44), .O(gate39inter3));
  inv1  gate859(.a(s_45), .O(gate39inter4));
  nand2 gate860(.a(gate39inter4), .b(gate39inter3), .O(gate39inter5));
  nor2  gate861(.a(gate39inter5), .b(gate39inter2), .O(gate39inter6));
  inv1  gate862(.a(G20), .O(gate39inter7));
  inv1  gate863(.a(G24), .O(gate39inter8));
  nand2 gate864(.a(gate39inter8), .b(gate39inter7), .O(gate39inter9));
  nand2 gate865(.a(s_45), .b(gate39inter3), .O(gate39inter10));
  nor2  gate866(.a(gate39inter10), .b(gate39inter9), .O(gate39inter11));
  nor2  gate867(.a(gate39inter11), .b(gate39inter6), .O(gate39inter12));
  nand2 gate868(.a(gate39inter12), .b(gate39inter1), .O(G356));
nand2 gate40( .a(G28), .b(G32), .O(G359) );
nand2 gate41( .a(G1), .b(G266), .O(G362) );
nand2 gate42( .a(G2), .b(G266), .O(G363) );
nand2 gate43( .a(G3), .b(G269), .O(G364) );

  xor2  gate1331(.a(G269), .b(G4), .O(gate44inter0));
  nand2 gate1332(.a(gate44inter0), .b(s_112), .O(gate44inter1));
  and2  gate1333(.a(G269), .b(G4), .O(gate44inter2));
  inv1  gate1334(.a(s_112), .O(gate44inter3));
  inv1  gate1335(.a(s_113), .O(gate44inter4));
  nand2 gate1336(.a(gate44inter4), .b(gate44inter3), .O(gate44inter5));
  nor2  gate1337(.a(gate44inter5), .b(gate44inter2), .O(gate44inter6));
  inv1  gate1338(.a(G4), .O(gate44inter7));
  inv1  gate1339(.a(G269), .O(gate44inter8));
  nand2 gate1340(.a(gate44inter8), .b(gate44inter7), .O(gate44inter9));
  nand2 gate1341(.a(s_113), .b(gate44inter3), .O(gate44inter10));
  nor2  gate1342(.a(gate44inter10), .b(gate44inter9), .O(gate44inter11));
  nor2  gate1343(.a(gate44inter11), .b(gate44inter6), .O(gate44inter12));
  nand2 gate1344(.a(gate44inter12), .b(gate44inter1), .O(G365));
nand2 gate45( .a(G5), .b(G272), .O(G366) );
nand2 gate46( .a(G6), .b(G272), .O(G367) );
nand2 gate47( .a(G7), .b(G275), .O(G368) );

  xor2  gate547(.a(G275), .b(G8), .O(gate48inter0));
  nand2 gate548(.a(gate48inter0), .b(s_0), .O(gate48inter1));
  and2  gate549(.a(G275), .b(G8), .O(gate48inter2));
  inv1  gate550(.a(s_0), .O(gate48inter3));
  inv1  gate551(.a(s_1), .O(gate48inter4));
  nand2 gate552(.a(gate48inter4), .b(gate48inter3), .O(gate48inter5));
  nor2  gate553(.a(gate48inter5), .b(gate48inter2), .O(gate48inter6));
  inv1  gate554(.a(G8), .O(gate48inter7));
  inv1  gate555(.a(G275), .O(gate48inter8));
  nand2 gate556(.a(gate48inter8), .b(gate48inter7), .O(gate48inter9));
  nand2 gate557(.a(s_1), .b(gate48inter3), .O(gate48inter10));
  nor2  gate558(.a(gate48inter10), .b(gate48inter9), .O(gate48inter11));
  nor2  gate559(.a(gate48inter11), .b(gate48inter6), .O(gate48inter12));
  nand2 gate560(.a(gate48inter12), .b(gate48inter1), .O(G369));
nand2 gate49( .a(G9), .b(G278), .O(G370) );
nand2 gate50( .a(G10), .b(G278), .O(G371) );

  xor2  gate1317(.a(G281), .b(G11), .O(gate51inter0));
  nand2 gate1318(.a(gate51inter0), .b(s_110), .O(gate51inter1));
  and2  gate1319(.a(G281), .b(G11), .O(gate51inter2));
  inv1  gate1320(.a(s_110), .O(gate51inter3));
  inv1  gate1321(.a(s_111), .O(gate51inter4));
  nand2 gate1322(.a(gate51inter4), .b(gate51inter3), .O(gate51inter5));
  nor2  gate1323(.a(gate51inter5), .b(gate51inter2), .O(gate51inter6));
  inv1  gate1324(.a(G11), .O(gate51inter7));
  inv1  gate1325(.a(G281), .O(gate51inter8));
  nand2 gate1326(.a(gate51inter8), .b(gate51inter7), .O(gate51inter9));
  nand2 gate1327(.a(s_111), .b(gate51inter3), .O(gate51inter10));
  nor2  gate1328(.a(gate51inter10), .b(gate51inter9), .O(gate51inter11));
  nor2  gate1329(.a(gate51inter11), .b(gate51inter6), .O(gate51inter12));
  nand2 gate1330(.a(gate51inter12), .b(gate51inter1), .O(G372));
nand2 gate52( .a(G12), .b(G281), .O(G373) );
nand2 gate53( .a(G13), .b(G284), .O(G374) );
nand2 gate54( .a(G14), .b(G284), .O(G375) );
nand2 gate55( .a(G15), .b(G287), .O(G376) );
nand2 gate56( .a(G16), .b(G287), .O(G377) );
nand2 gate57( .a(G17), .b(G290), .O(G378) );

  xor2  gate785(.a(G290), .b(G18), .O(gate58inter0));
  nand2 gate786(.a(gate58inter0), .b(s_34), .O(gate58inter1));
  and2  gate787(.a(G290), .b(G18), .O(gate58inter2));
  inv1  gate788(.a(s_34), .O(gate58inter3));
  inv1  gate789(.a(s_35), .O(gate58inter4));
  nand2 gate790(.a(gate58inter4), .b(gate58inter3), .O(gate58inter5));
  nor2  gate791(.a(gate58inter5), .b(gate58inter2), .O(gate58inter6));
  inv1  gate792(.a(G18), .O(gate58inter7));
  inv1  gate793(.a(G290), .O(gate58inter8));
  nand2 gate794(.a(gate58inter8), .b(gate58inter7), .O(gate58inter9));
  nand2 gate795(.a(s_35), .b(gate58inter3), .O(gate58inter10));
  nor2  gate796(.a(gate58inter10), .b(gate58inter9), .O(gate58inter11));
  nor2  gate797(.a(gate58inter11), .b(gate58inter6), .O(gate58inter12));
  nand2 gate798(.a(gate58inter12), .b(gate58inter1), .O(G379));
nand2 gate59( .a(G19), .b(G293), .O(G380) );
nand2 gate60( .a(G20), .b(G293), .O(G381) );
nand2 gate61( .a(G21), .b(G296), .O(G382) );
nand2 gate62( .a(G22), .b(G296), .O(G383) );
nand2 gate63( .a(G23), .b(G299), .O(G384) );
nand2 gate64( .a(G24), .b(G299), .O(G385) );
nand2 gate65( .a(G25), .b(G302), .O(G386) );

  xor2  gate1387(.a(G302), .b(G26), .O(gate66inter0));
  nand2 gate1388(.a(gate66inter0), .b(s_120), .O(gate66inter1));
  and2  gate1389(.a(G302), .b(G26), .O(gate66inter2));
  inv1  gate1390(.a(s_120), .O(gate66inter3));
  inv1  gate1391(.a(s_121), .O(gate66inter4));
  nand2 gate1392(.a(gate66inter4), .b(gate66inter3), .O(gate66inter5));
  nor2  gate1393(.a(gate66inter5), .b(gate66inter2), .O(gate66inter6));
  inv1  gate1394(.a(G26), .O(gate66inter7));
  inv1  gate1395(.a(G302), .O(gate66inter8));
  nand2 gate1396(.a(gate66inter8), .b(gate66inter7), .O(gate66inter9));
  nand2 gate1397(.a(s_121), .b(gate66inter3), .O(gate66inter10));
  nor2  gate1398(.a(gate66inter10), .b(gate66inter9), .O(gate66inter11));
  nor2  gate1399(.a(gate66inter11), .b(gate66inter6), .O(gate66inter12));
  nand2 gate1400(.a(gate66inter12), .b(gate66inter1), .O(G387));
nand2 gate67( .a(G27), .b(G305), .O(G388) );
nand2 gate68( .a(G28), .b(G305), .O(G389) );
nand2 gate69( .a(G29), .b(G308), .O(G390) );
nand2 gate70( .a(G30), .b(G308), .O(G391) );
nand2 gate71( .a(G31), .b(G311), .O(G392) );
nand2 gate72( .a(G32), .b(G311), .O(G393) );
nand2 gate73( .a(G1), .b(G314), .O(G394) );
nand2 gate74( .a(G5), .b(G314), .O(G395) );
nand2 gate75( .a(G9), .b(G317), .O(G396) );
nand2 gate76( .a(G13), .b(G317), .O(G397) );
nand2 gate77( .a(G2), .b(G320), .O(G398) );
nand2 gate78( .a(G6), .b(G320), .O(G399) );
nand2 gate79( .a(G10), .b(G323), .O(G400) );
nand2 gate80( .a(G14), .b(G323), .O(G401) );
nand2 gate81( .a(G3), .b(G326), .O(G402) );
nand2 gate82( .a(G7), .b(G326), .O(G403) );
nand2 gate83( .a(G11), .b(G329), .O(G404) );
nand2 gate84( .a(G15), .b(G329), .O(G405) );
nand2 gate85( .a(G4), .b(G332), .O(G406) );

  xor2  gate1373(.a(G332), .b(G8), .O(gate86inter0));
  nand2 gate1374(.a(gate86inter0), .b(s_118), .O(gate86inter1));
  and2  gate1375(.a(G332), .b(G8), .O(gate86inter2));
  inv1  gate1376(.a(s_118), .O(gate86inter3));
  inv1  gate1377(.a(s_119), .O(gate86inter4));
  nand2 gate1378(.a(gate86inter4), .b(gate86inter3), .O(gate86inter5));
  nor2  gate1379(.a(gate86inter5), .b(gate86inter2), .O(gate86inter6));
  inv1  gate1380(.a(G8), .O(gate86inter7));
  inv1  gate1381(.a(G332), .O(gate86inter8));
  nand2 gate1382(.a(gate86inter8), .b(gate86inter7), .O(gate86inter9));
  nand2 gate1383(.a(s_119), .b(gate86inter3), .O(gate86inter10));
  nor2  gate1384(.a(gate86inter10), .b(gate86inter9), .O(gate86inter11));
  nor2  gate1385(.a(gate86inter11), .b(gate86inter6), .O(gate86inter12));
  nand2 gate1386(.a(gate86inter12), .b(gate86inter1), .O(G407));
nand2 gate87( .a(G12), .b(G335), .O(G408) );
nand2 gate88( .a(G16), .b(G335), .O(G409) );

  xor2  gate1205(.a(G338), .b(G17), .O(gate89inter0));
  nand2 gate1206(.a(gate89inter0), .b(s_94), .O(gate89inter1));
  and2  gate1207(.a(G338), .b(G17), .O(gate89inter2));
  inv1  gate1208(.a(s_94), .O(gate89inter3));
  inv1  gate1209(.a(s_95), .O(gate89inter4));
  nand2 gate1210(.a(gate89inter4), .b(gate89inter3), .O(gate89inter5));
  nor2  gate1211(.a(gate89inter5), .b(gate89inter2), .O(gate89inter6));
  inv1  gate1212(.a(G17), .O(gate89inter7));
  inv1  gate1213(.a(G338), .O(gate89inter8));
  nand2 gate1214(.a(gate89inter8), .b(gate89inter7), .O(gate89inter9));
  nand2 gate1215(.a(s_95), .b(gate89inter3), .O(gate89inter10));
  nor2  gate1216(.a(gate89inter10), .b(gate89inter9), .O(gate89inter11));
  nor2  gate1217(.a(gate89inter11), .b(gate89inter6), .O(gate89inter12));
  nand2 gate1218(.a(gate89inter12), .b(gate89inter1), .O(G410));
nand2 gate90( .a(G21), .b(G338), .O(G411) );
nand2 gate91( .a(G25), .b(G341), .O(G412) );
nand2 gate92( .a(G29), .b(G341), .O(G413) );

  xor2  gate1345(.a(G344), .b(G18), .O(gate93inter0));
  nand2 gate1346(.a(gate93inter0), .b(s_114), .O(gate93inter1));
  and2  gate1347(.a(G344), .b(G18), .O(gate93inter2));
  inv1  gate1348(.a(s_114), .O(gate93inter3));
  inv1  gate1349(.a(s_115), .O(gate93inter4));
  nand2 gate1350(.a(gate93inter4), .b(gate93inter3), .O(gate93inter5));
  nor2  gate1351(.a(gate93inter5), .b(gate93inter2), .O(gate93inter6));
  inv1  gate1352(.a(G18), .O(gate93inter7));
  inv1  gate1353(.a(G344), .O(gate93inter8));
  nand2 gate1354(.a(gate93inter8), .b(gate93inter7), .O(gate93inter9));
  nand2 gate1355(.a(s_115), .b(gate93inter3), .O(gate93inter10));
  nor2  gate1356(.a(gate93inter10), .b(gate93inter9), .O(gate93inter11));
  nor2  gate1357(.a(gate93inter11), .b(gate93inter6), .O(gate93inter12));
  nand2 gate1358(.a(gate93inter12), .b(gate93inter1), .O(G414));

  xor2  gate1233(.a(G344), .b(G22), .O(gate94inter0));
  nand2 gate1234(.a(gate94inter0), .b(s_98), .O(gate94inter1));
  and2  gate1235(.a(G344), .b(G22), .O(gate94inter2));
  inv1  gate1236(.a(s_98), .O(gate94inter3));
  inv1  gate1237(.a(s_99), .O(gate94inter4));
  nand2 gate1238(.a(gate94inter4), .b(gate94inter3), .O(gate94inter5));
  nor2  gate1239(.a(gate94inter5), .b(gate94inter2), .O(gate94inter6));
  inv1  gate1240(.a(G22), .O(gate94inter7));
  inv1  gate1241(.a(G344), .O(gate94inter8));
  nand2 gate1242(.a(gate94inter8), .b(gate94inter7), .O(gate94inter9));
  nand2 gate1243(.a(s_99), .b(gate94inter3), .O(gate94inter10));
  nor2  gate1244(.a(gate94inter10), .b(gate94inter9), .O(gate94inter11));
  nor2  gate1245(.a(gate94inter11), .b(gate94inter6), .O(gate94inter12));
  nand2 gate1246(.a(gate94inter12), .b(gate94inter1), .O(G415));
nand2 gate95( .a(G26), .b(G347), .O(G416) );
nand2 gate96( .a(G30), .b(G347), .O(G417) );
nand2 gate97( .a(G19), .b(G350), .O(G418) );
nand2 gate98( .a(G23), .b(G350), .O(G419) );
nand2 gate99( .a(G27), .b(G353), .O(G420) );

  xor2  gate1051(.a(G353), .b(G31), .O(gate100inter0));
  nand2 gate1052(.a(gate100inter0), .b(s_72), .O(gate100inter1));
  and2  gate1053(.a(G353), .b(G31), .O(gate100inter2));
  inv1  gate1054(.a(s_72), .O(gate100inter3));
  inv1  gate1055(.a(s_73), .O(gate100inter4));
  nand2 gate1056(.a(gate100inter4), .b(gate100inter3), .O(gate100inter5));
  nor2  gate1057(.a(gate100inter5), .b(gate100inter2), .O(gate100inter6));
  inv1  gate1058(.a(G31), .O(gate100inter7));
  inv1  gate1059(.a(G353), .O(gate100inter8));
  nand2 gate1060(.a(gate100inter8), .b(gate100inter7), .O(gate100inter9));
  nand2 gate1061(.a(s_73), .b(gate100inter3), .O(gate100inter10));
  nor2  gate1062(.a(gate100inter10), .b(gate100inter9), .O(gate100inter11));
  nor2  gate1063(.a(gate100inter11), .b(gate100inter6), .O(gate100inter12));
  nand2 gate1064(.a(gate100inter12), .b(gate100inter1), .O(G421));
nand2 gate101( .a(G20), .b(G356), .O(G422) );
nand2 gate102( .a(G24), .b(G356), .O(G423) );

  xor2  gate1513(.a(G359), .b(G28), .O(gate103inter0));
  nand2 gate1514(.a(gate103inter0), .b(s_138), .O(gate103inter1));
  and2  gate1515(.a(G359), .b(G28), .O(gate103inter2));
  inv1  gate1516(.a(s_138), .O(gate103inter3));
  inv1  gate1517(.a(s_139), .O(gate103inter4));
  nand2 gate1518(.a(gate103inter4), .b(gate103inter3), .O(gate103inter5));
  nor2  gate1519(.a(gate103inter5), .b(gate103inter2), .O(gate103inter6));
  inv1  gate1520(.a(G28), .O(gate103inter7));
  inv1  gate1521(.a(G359), .O(gate103inter8));
  nand2 gate1522(.a(gate103inter8), .b(gate103inter7), .O(gate103inter9));
  nand2 gate1523(.a(s_139), .b(gate103inter3), .O(gate103inter10));
  nor2  gate1524(.a(gate103inter10), .b(gate103inter9), .O(gate103inter11));
  nor2  gate1525(.a(gate103inter11), .b(gate103inter6), .O(gate103inter12));
  nand2 gate1526(.a(gate103inter12), .b(gate103inter1), .O(G424));
nand2 gate104( .a(G32), .b(G359), .O(G425) );
nand2 gate105( .a(G362), .b(G363), .O(G426) );
nand2 gate106( .a(G364), .b(G365), .O(G429) );
nand2 gate107( .a(G366), .b(G367), .O(G432) );
nand2 gate108( .a(G368), .b(G369), .O(G435) );
nand2 gate109( .a(G370), .b(G371), .O(G438) );
nand2 gate110( .a(G372), .b(G373), .O(G441) );

  xor2  gate1037(.a(G375), .b(G374), .O(gate111inter0));
  nand2 gate1038(.a(gate111inter0), .b(s_70), .O(gate111inter1));
  and2  gate1039(.a(G375), .b(G374), .O(gate111inter2));
  inv1  gate1040(.a(s_70), .O(gate111inter3));
  inv1  gate1041(.a(s_71), .O(gate111inter4));
  nand2 gate1042(.a(gate111inter4), .b(gate111inter3), .O(gate111inter5));
  nor2  gate1043(.a(gate111inter5), .b(gate111inter2), .O(gate111inter6));
  inv1  gate1044(.a(G374), .O(gate111inter7));
  inv1  gate1045(.a(G375), .O(gate111inter8));
  nand2 gate1046(.a(gate111inter8), .b(gate111inter7), .O(gate111inter9));
  nand2 gate1047(.a(s_71), .b(gate111inter3), .O(gate111inter10));
  nor2  gate1048(.a(gate111inter10), .b(gate111inter9), .O(gate111inter11));
  nor2  gate1049(.a(gate111inter11), .b(gate111inter6), .O(gate111inter12));
  nand2 gate1050(.a(gate111inter12), .b(gate111inter1), .O(G444));
nand2 gate112( .a(G376), .b(G377), .O(G447) );
nand2 gate113( .a(G378), .b(G379), .O(G450) );
nand2 gate114( .a(G380), .b(G381), .O(G453) );
nand2 gate115( .a(G382), .b(G383), .O(G456) );
nand2 gate116( .a(G384), .b(G385), .O(G459) );

  xor2  gate1107(.a(G387), .b(G386), .O(gate117inter0));
  nand2 gate1108(.a(gate117inter0), .b(s_80), .O(gate117inter1));
  and2  gate1109(.a(G387), .b(G386), .O(gate117inter2));
  inv1  gate1110(.a(s_80), .O(gate117inter3));
  inv1  gate1111(.a(s_81), .O(gate117inter4));
  nand2 gate1112(.a(gate117inter4), .b(gate117inter3), .O(gate117inter5));
  nor2  gate1113(.a(gate117inter5), .b(gate117inter2), .O(gate117inter6));
  inv1  gate1114(.a(G386), .O(gate117inter7));
  inv1  gate1115(.a(G387), .O(gate117inter8));
  nand2 gate1116(.a(gate117inter8), .b(gate117inter7), .O(gate117inter9));
  nand2 gate1117(.a(s_81), .b(gate117inter3), .O(gate117inter10));
  nor2  gate1118(.a(gate117inter10), .b(gate117inter9), .O(gate117inter11));
  nor2  gate1119(.a(gate117inter11), .b(gate117inter6), .O(gate117inter12));
  nand2 gate1120(.a(gate117inter12), .b(gate117inter1), .O(G462));

  xor2  gate967(.a(G389), .b(G388), .O(gate118inter0));
  nand2 gate968(.a(gate118inter0), .b(s_60), .O(gate118inter1));
  and2  gate969(.a(G389), .b(G388), .O(gate118inter2));
  inv1  gate970(.a(s_60), .O(gate118inter3));
  inv1  gate971(.a(s_61), .O(gate118inter4));
  nand2 gate972(.a(gate118inter4), .b(gate118inter3), .O(gate118inter5));
  nor2  gate973(.a(gate118inter5), .b(gate118inter2), .O(gate118inter6));
  inv1  gate974(.a(G388), .O(gate118inter7));
  inv1  gate975(.a(G389), .O(gate118inter8));
  nand2 gate976(.a(gate118inter8), .b(gate118inter7), .O(gate118inter9));
  nand2 gate977(.a(s_61), .b(gate118inter3), .O(gate118inter10));
  nor2  gate978(.a(gate118inter10), .b(gate118inter9), .O(gate118inter11));
  nor2  gate979(.a(gate118inter11), .b(gate118inter6), .O(gate118inter12));
  nand2 gate980(.a(gate118inter12), .b(gate118inter1), .O(G465));

  xor2  gate1541(.a(G391), .b(G390), .O(gate119inter0));
  nand2 gate1542(.a(gate119inter0), .b(s_142), .O(gate119inter1));
  and2  gate1543(.a(G391), .b(G390), .O(gate119inter2));
  inv1  gate1544(.a(s_142), .O(gate119inter3));
  inv1  gate1545(.a(s_143), .O(gate119inter4));
  nand2 gate1546(.a(gate119inter4), .b(gate119inter3), .O(gate119inter5));
  nor2  gate1547(.a(gate119inter5), .b(gate119inter2), .O(gate119inter6));
  inv1  gate1548(.a(G390), .O(gate119inter7));
  inv1  gate1549(.a(G391), .O(gate119inter8));
  nand2 gate1550(.a(gate119inter8), .b(gate119inter7), .O(gate119inter9));
  nand2 gate1551(.a(s_143), .b(gate119inter3), .O(gate119inter10));
  nor2  gate1552(.a(gate119inter10), .b(gate119inter9), .O(gate119inter11));
  nor2  gate1553(.a(gate119inter11), .b(gate119inter6), .O(gate119inter12));
  nand2 gate1554(.a(gate119inter12), .b(gate119inter1), .O(G468));
nand2 gate120( .a(G392), .b(G393), .O(G471) );
nand2 gate121( .a(G394), .b(G395), .O(G474) );
nand2 gate122( .a(G396), .b(G397), .O(G477) );
nand2 gate123( .a(G398), .b(G399), .O(G480) );
nand2 gate124( .a(G400), .b(G401), .O(G483) );
nand2 gate125( .a(G402), .b(G403), .O(G486) );
nand2 gate126( .a(G404), .b(G405), .O(G489) );
nand2 gate127( .a(G406), .b(G407), .O(G492) );
nand2 gate128( .a(G408), .b(G409), .O(G495) );
nand2 gate129( .a(G410), .b(G411), .O(G498) );

  xor2  gate1597(.a(G413), .b(G412), .O(gate130inter0));
  nand2 gate1598(.a(gate130inter0), .b(s_150), .O(gate130inter1));
  and2  gate1599(.a(G413), .b(G412), .O(gate130inter2));
  inv1  gate1600(.a(s_150), .O(gate130inter3));
  inv1  gate1601(.a(s_151), .O(gate130inter4));
  nand2 gate1602(.a(gate130inter4), .b(gate130inter3), .O(gate130inter5));
  nor2  gate1603(.a(gate130inter5), .b(gate130inter2), .O(gate130inter6));
  inv1  gate1604(.a(G412), .O(gate130inter7));
  inv1  gate1605(.a(G413), .O(gate130inter8));
  nand2 gate1606(.a(gate130inter8), .b(gate130inter7), .O(gate130inter9));
  nand2 gate1607(.a(s_151), .b(gate130inter3), .O(gate130inter10));
  nor2  gate1608(.a(gate130inter10), .b(gate130inter9), .O(gate130inter11));
  nor2  gate1609(.a(gate130inter11), .b(gate130inter6), .O(gate130inter12));
  nand2 gate1610(.a(gate130inter12), .b(gate130inter1), .O(G501));
nand2 gate131( .a(G414), .b(G415), .O(G504) );
nand2 gate132( .a(G416), .b(G417), .O(G507) );
nand2 gate133( .a(G418), .b(G419), .O(G510) );
nand2 gate134( .a(G420), .b(G421), .O(G513) );

  xor2  gate743(.a(G423), .b(G422), .O(gate135inter0));
  nand2 gate744(.a(gate135inter0), .b(s_28), .O(gate135inter1));
  and2  gate745(.a(G423), .b(G422), .O(gate135inter2));
  inv1  gate746(.a(s_28), .O(gate135inter3));
  inv1  gate747(.a(s_29), .O(gate135inter4));
  nand2 gate748(.a(gate135inter4), .b(gate135inter3), .O(gate135inter5));
  nor2  gate749(.a(gate135inter5), .b(gate135inter2), .O(gate135inter6));
  inv1  gate750(.a(G422), .O(gate135inter7));
  inv1  gate751(.a(G423), .O(gate135inter8));
  nand2 gate752(.a(gate135inter8), .b(gate135inter7), .O(gate135inter9));
  nand2 gate753(.a(s_29), .b(gate135inter3), .O(gate135inter10));
  nor2  gate754(.a(gate135inter10), .b(gate135inter9), .O(gate135inter11));
  nor2  gate755(.a(gate135inter11), .b(gate135inter6), .O(gate135inter12));
  nand2 gate756(.a(gate135inter12), .b(gate135inter1), .O(G516));
nand2 gate136( .a(G424), .b(G425), .O(G519) );
nand2 gate137( .a(G426), .b(G429), .O(G522) );
nand2 gate138( .a(G432), .b(G435), .O(G525) );
nand2 gate139( .a(G438), .b(G441), .O(G528) );
nand2 gate140( .a(G444), .b(G447), .O(G531) );
nand2 gate141( .a(G450), .b(G453), .O(G534) );

  xor2  gate589(.a(G459), .b(G456), .O(gate142inter0));
  nand2 gate590(.a(gate142inter0), .b(s_6), .O(gate142inter1));
  and2  gate591(.a(G459), .b(G456), .O(gate142inter2));
  inv1  gate592(.a(s_6), .O(gate142inter3));
  inv1  gate593(.a(s_7), .O(gate142inter4));
  nand2 gate594(.a(gate142inter4), .b(gate142inter3), .O(gate142inter5));
  nor2  gate595(.a(gate142inter5), .b(gate142inter2), .O(gate142inter6));
  inv1  gate596(.a(G456), .O(gate142inter7));
  inv1  gate597(.a(G459), .O(gate142inter8));
  nand2 gate598(.a(gate142inter8), .b(gate142inter7), .O(gate142inter9));
  nand2 gate599(.a(s_7), .b(gate142inter3), .O(gate142inter10));
  nor2  gate600(.a(gate142inter10), .b(gate142inter9), .O(gate142inter11));
  nor2  gate601(.a(gate142inter11), .b(gate142inter6), .O(gate142inter12));
  nand2 gate602(.a(gate142inter12), .b(gate142inter1), .O(G537));
nand2 gate143( .a(G462), .b(G465), .O(G540) );
nand2 gate144( .a(G468), .b(G471), .O(G543) );
nand2 gate145( .a(G474), .b(G477), .O(G546) );
nand2 gate146( .a(G480), .b(G483), .O(G549) );

  xor2  gate1247(.a(G489), .b(G486), .O(gate147inter0));
  nand2 gate1248(.a(gate147inter0), .b(s_100), .O(gate147inter1));
  and2  gate1249(.a(G489), .b(G486), .O(gate147inter2));
  inv1  gate1250(.a(s_100), .O(gate147inter3));
  inv1  gate1251(.a(s_101), .O(gate147inter4));
  nand2 gate1252(.a(gate147inter4), .b(gate147inter3), .O(gate147inter5));
  nor2  gate1253(.a(gate147inter5), .b(gate147inter2), .O(gate147inter6));
  inv1  gate1254(.a(G486), .O(gate147inter7));
  inv1  gate1255(.a(G489), .O(gate147inter8));
  nand2 gate1256(.a(gate147inter8), .b(gate147inter7), .O(gate147inter9));
  nand2 gate1257(.a(s_101), .b(gate147inter3), .O(gate147inter10));
  nor2  gate1258(.a(gate147inter10), .b(gate147inter9), .O(gate147inter11));
  nor2  gate1259(.a(gate147inter11), .b(gate147inter6), .O(gate147inter12));
  nand2 gate1260(.a(gate147inter12), .b(gate147inter1), .O(G552));

  xor2  gate1499(.a(G495), .b(G492), .O(gate148inter0));
  nand2 gate1500(.a(gate148inter0), .b(s_136), .O(gate148inter1));
  and2  gate1501(.a(G495), .b(G492), .O(gate148inter2));
  inv1  gate1502(.a(s_136), .O(gate148inter3));
  inv1  gate1503(.a(s_137), .O(gate148inter4));
  nand2 gate1504(.a(gate148inter4), .b(gate148inter3), .O(gate148inter5));
  nor2  gate1505(.a(gate148inter5), .b(gate148inter2), .O(gate148inter6));
  inv1  gate1506(.a(G492), .O(gate148inter7));
  inv1  gate1507(.a(G495), .O(gate148inter8));
  nand2 gate1508(.a(gate148inter8), .b(gate148inter7), .O(gate148inter9));
  nand2 gate1509(.a(s_137), .b(gate148inter3), .O(gate148inter10));
  nor2  gate1510(.a(gate148inter10), .b(gate148inter9), .O(gate148inter11));
  nor2  gate1511(.a(gate148inter11), .b(gate148inter6), .O(gate148inter12));
  nand2 gate1512(.a(gate148inter12), .b(gate148inter1), .O(G555));
nand2 gate149( .a(G498), .b(G501), .O(G558) );
nand2 gate150( .a(G504), .b(G507), .O(G561) );
nand2 gate151( .a(G510), .b(G513), .O(G564) );

  xor2  gate1289(.a(G519), .b(G516), .O(gate152inter0));
  nand2 gate1290(.a(gate152inter0), .b(s_106), .O(gate152inter1));
  and2  gate1291(.a(G519), .b(G516), .O(gate152inter2));
  inv1  gate1292(.a(s_106), .O(gate152inter3));
  inv1  gate1293(.a(s_107), .O(gate152inter4));
  nand2 gate1294(.a(gate152inter4), .b(gate152inter3), .O(gate152inter5));
  nor2  gate1295(.a(gate152inter5), .b(gate152inter2), .O(gate152inter6));
  inv1  gate1296(.a(G516), .O(gate152inter7));
  inv1  gate1297(.a(G519), .O(gate152inter8));
  nand2 gate1298(.a(gate152inter8), .b(gate152inter7), .O(gate152inter9));
  nand2 gate1299(.a(s_107), .b(gate152inter3), .O(gate152inter10));
  nor2  gate1300(.a(gate152inter10), .b(gate152inter9), .O(gate152inter11));
  nor2  gate1301(.a(gate152inter11), .b(gate152inter6), .O(gate152inter12));
  nand2 gate1302(.a(gate152inter12), .b(gate152inter1), .O(G567));
nand2 gate153( .a(G426), .b(G522), .O(G570) );
nand2 gate154( .a(G429), .b(G522), .O(G571) );
nand2 gate155( .a(G432), .b(G525), .O(G572) );
nand2 gate156( .a(G435), .b(G525), .O(G573) );

  xor2  gate617(.a(G528), .b(G438), .O(gate157inter0));
  nand2 gate618(.a(gate157inter0), .b(s_10), .O(gate157inter1));
  and2  gate619(.a(G528), .b(G438), .O(gate157inter2));
  inv1  gate620(.a(s_10), .O(gate157inter3));
  inv1  gate621(.a(s_11), .O(gate157inter4));
  nand2 gate622(.a(gate157inter4), .b(gate157inter3), .O(gate157inter5));
  nor2  gate623(.a(gate157inter5), .b(gate157inter2), .O(gate157inter6));
  inv1  gate624(.a(G438), .O(gate157inter7));
  inv1  gate625(.a(G528), .O(gate157inter8));
  nand2 gate626(.a(gate157inter8), .b(gate157inter7), .O(gate157inter9));
  nand2 gate627(.a(s_11), .b(gate157inter3), .O(gate157inter10));
  nor2  gate628(.a(gate157inter10), .b(gate157inter9), .O(gate157inter11));
  nor2  gate629(.a(gate157inter11), .b(gate157inter6), .O(gate157inter12));
  nand2 gate630(.a(gate157inter12), .b(gate157inter1), .O(G574));
nand2 gate158( .a(G441), .b(G528), .O(G575) );
nand2 gate159( .a(G444), .b(G531), .O(G576) );
nand2 gate160( .a(G447), .b(G531), .O(G577) );

  xor2  gate1485(.a(G534), .b(G450), .O(gate161inter0));
  nand2 gate1486(.a(gate161inter0), .b(s_134), .O(gate161inter1));
  and2  gate1487(.a(G534), .b(G450), .O(gate161inter2));
  inv1  gate1488(.a(s_134), .O(gate161inter3));
  inv1  gate1489(.a(s_135), .O(gate161inter4));
  nand2 gate1490(.a(gate161inter4), .b(gate161inter3), .O(gate161inter5));
  nor2  gate1491(.a(gate161inter5), .b(gate161inter2), .O(gate161inter6));
  inv1  gate1492(.a(G450), .O(gate161inter7));
  inv1  gate1493(.a(G534), .O(gate161inter8));
  nand2 gate1494(.a(gate161inter8), .b(gate161inter7), .O(gate161inter9));
  nand2 gate1495(.a(s_135), .b(gate161inter3), .O(gate161inter10));
  nor2  gate1496(.a(gate161inter10), .b(gate161inter9), .O(gate161inter11));
  nor2  gate1497(.a(gate161inter11), .b(gate161inter6), .O(gate161inter12));
  nand2 gate1498(.a(gate161inter12), .b(gate161inter1), .O(G578));
nand2 gate162( .a(G453), .b(G534), .O(G579) );

  xor2  gate771(.a(G537), .b(G456), .O(gate163inter0));
  nand2 gate772(.a(gate163inter0), .b(s_32), .O(gate163inter1));
  and2  gate773(.a(G537), .b(G456), .O(gate163inter2));
  inv1  gate774(.a(s_32), .O(gate163inter3));
  inv1  gate775(.a(s_33), .O(gate163inter4));
  nand2 gate776(.a(gate163inter4), .b(gate163inter3), .O(gate163inter5));
  nor2  gate777(.a(gate163inter5), .b(gate163inter2), .O(gate163inter6));
  inv1  gate778(.a(G456), .O(gate163inter7));
  inv1  gate779(.a(G537), .O(gate163inter8));
  nand2 gate780(.a(gate163inter8), .b(gate163inter7), .O(gate163inter9));
  nand2 gate781(.a(s_33), .b(gate163inter3), .O(gate163inter10));
  nor2  gate782(.a(gate163inter10), .b(gate163inter9), .O(gate163inter11));
  nor2  gate783(.a(gate163inter11), .b(gate163inter6), .O(gate163inter12));
  nand2 gate784(.a(gate163inter12), .b(gate163inter1), .O(G580));

  xor2  gate883(.a(G537), .b(G459), .O(gate164inter0));
  nand2 gate884(.a(gate164inter0), .b(s_48), .O(gate164inter1));
  and2  gate885(.a(G537), .b(G459), .O(gate164inter2));
  inv1  gate886(.a(s_48), .O(gate164inter3));
  inv1  gate887(.a(s_49), .O(gate164inter4));
  nand2 gate888(.a(gate164inter4), .b(gate164inter3), .O(gate164inter5));
  nor2  gate889(.a(gate164inter5), .b(gate164inter2), .O(gate164inter6));
  inv1  gate890(.a(G459), .O(gate164inter7));
  inv1  gate891(.a(G537), .O(gate164inter8));
  nand2 gate892(.a(gate164inter8), .b(gate164inter7), .O(gate164inter9));
  nand2 gate893(.a(s_49), .b(gate164inter3), .O(gate164inter10));
  nor2  gate894(.a(gate164inter10), .b(gate164inter9), .O(gate164inter11));
  nor2  gate895(.a(gate164inter11), .b(gate164inter6), .O(gate164inter12));
  nand2 gate896(.a(gate164inter12), .b(gate164inter1), .O(G581));
nand2 gate165( .a(G462), .b(G540), .O(G582) );
nand2 gate166( .a(G465), .b(G540), .O(G583) );
nand2 gate167( .a(G468), .b(G543), .O(G584) );
nand2 gate168( .a(G471), .b(G543), .O(G585) );
nand2 gate169( .a(G474), .b(G546), .O(G586) );
nand2 gate170( .a(G477), .b(G546), .O(G587) );
nand2 gate171( .a(G480), .b(G549), .O(G588) );
nand2 gate172( .a(G483), .b(G549), .O(G589) );

  xor2  gate1149(.a(G552), .b(G486), .O(gate173inter0));
  nand2 gate1150(.a(gate173inter0), .b(s_86), .O(gate173inter1));
  and2  gate1151(.a(G552), .b(G486), .O(gate173inter2));
  inv1  gate1152(.a(s_86), .O(gate173inter3));
  inv1  gate1153(.a(s_87), .O(gate173inter4));
  nand2 gate1154(.a(gate173inter4), .b(gate173inter3), .O(gate173inter5));
  nor2  gate1155(.a(gate173inter5), .b(gate173inter2), .O(gate173inter6));
  inv1  gate1156(.a(G486), .O(gate173inter7));
  inv1  gate1157(.a(G552), .O(gate173inter8));
  nand2 gate1158(.a(gate173inter8), .b(gate173inter7), .O(gate173inter9));
  nand2 gate1159(.a(s_87), .b(gate173inter3), .O(gate173inter10));
  nor2  gate1160(.a(gate173inter10), .b(gate173inter9), .O(gate173inter11));
  nor2  gate1161(.a(gate173inter11), .b(gate173inter6), .O(gate173inter12));
  nand2 gate1162(.a(gate173inter12), .b(gate173inter1), .O(G590));
nand2 gate174( .a(G489), .b(G552), .O(G591) );
nand2 gate175( .a(G492), .b(G555), .O(G592) );
nand2 gate176( .a(G495), .b(G555), .O(G593) );
nand2 gate177( .a(G498), .b(G558), .O(G594) );
nand2 gate178( .a(G501), .b(G558), .O(G595) );
nand2 gate179( .a(G504), .b(G561), .O(G596) );

  xor2  gate1457(.a(G561), .b(G507), .O(gate180inter0));
  nand2 gate1458(.a(gate180inter0), .b(s_130), .O(gate180inter1));
  and2  gate1459(.a(G561), .b(G507), .O(gate180inter2));
  inv1  gate1460(.a(s_130), .O(gate180inter3));
  inv1  gate1461(.a(s_131), .O(gate180inter4));
  nand2 gate1462(.a(gate180inter4), .b(gate180inter3), .O(gate180inter5));
  nor2  gate1463(.a(gate180inter5), .b(gate180inter2), .O(gate180inter6));
  inv1  gate1464(.a(G507), .O(gate180inter7));
  inv1  gate1465(.a(G561), .O(gate180inter8));
  nand2 gate1466(.a(gate180inter8), .b(gate180inter7), .O(gate180inter9));
  nand2 gate1467(.a(s_131), .b(gate180inter3), .O(gate180inter10));
  nor2  gate1468(.a(gate180inter10), .b(gate180inter9), .O(gate180inter11));
  nor2  gate1469(.a(gate180inter11), .b(gate180inter6), .O(gate180inter12));
  nand2 gate1470(.a(gate180inter12), .b(gate180inter1), .O(G597));

  xor2  gate939(.a(G564), .b(G510), .O(gate181inter0));
  nand2 gate940(.a(gate181inter0), .b(s_56), .O(gate181inter1));
  and2  gate941(.a(G564), .b(G510), .O(gate181inter2));
  inv1  gate942(.a(s_56), .O(gate181inter3));
  inv1  gate943(.a(s_57), .O(gate181inter4));
  nand2 gate944(.a(gate181inter4), .b(gate181inter3), .O(gate181inter5));
  nor2  gate945(.a(gate181inter5), .b(gate181inter2), .O(gate181inter6));
  inv1  gate946(.a(G510), .O(gate181inter7));
  inv1  gate947(.a(G564), .O(gate181inter8));
  nand2 gate948(.a(gate181inter8), .b(gate181inter7), .O(gate181inter9));
  nand2 gate949(.a(s_57), .b(gate181inter3), .O(gate181inter10));
  nor2  gate950(.a(gate181inter10), .b(gate181inter9), .O(gate181inter11));
  nor2  gate951(.a(gate181inter11), .b(gate181inter6), .O(gate181inter12));
  nand2 gate952(.a(gate181inter12), .b(gate181inter1), .O(G598));

  xor2  gate1429(.a(G564), .b(G513), .O(gate182inter0));
  nand2 gate1430(.a(gate182inter0), .b(s_126), .O(gate182inter1));
  and2  gate1431(.a(G564), .b(G513), .O(gate182inter2));
  inv1  gate1432(.a(s_126), .O(gate182inter3));
  inv1  gate1433(.a(s_127), .O(gate182inter4));
  nand2 gate1434(.a(gate182inter4), .b(gate182inter3), .O(gate182inter5));
  nor2  gate1435(.a(gate182inter5), .b(gate182inter2), .O(gate182inter6));
  inv1  gate1436(.a(G513), .O(gate182inter7));
  inv1  gate1437(.a(G564), .O(gate182inter8));
  nand2 gate1438(.a(gate182inter8), .b(gate182inter7), .O(gate182inter9));
  nand2 gate1439(.a(s_127), .b(gate182inter3), .O(gate182inter10));
  nor2  gate1440(.a(gate182inter10), .b(gate182inter9), .O(gate182inter11));
  nor2  gate1441(.a(gate182inter11), .b(gate182inter6), .O(gate182inter12));
  nand2 gate1442(.a(gate182inter12), .b(gate182inter1), .O(G599));
nand2 gate183( .a(G516), .b(G567), .O(G600) );

  xor2  gate1583(.a(G567), .b(G519), .O(gate184inter0));
  nand2 gate1584(.a(gate184inter0), .b(s_148), .O(gate184inter1));
  and2  gate1585(.a(G567), .b(G519), .O(gate184inter2));
  inv1  gate1586(.a(s_148), .O(gate184inter3));
  inv1  gate1587(.a(s_149), .O(gate184inter4));
  nand2 gate1588(.a(gate184inter4), .b(gate184inter3), .O(gate184inter5));
  nor2  gate1589(.a(gate184inter5), .b(gate184inter2), .O(gate184inter6));
  inv1  gate1590(.a(G519), .O(gate184inter7));
  inv1  gate1591(.a(G567), .O(gate184inter8));
  nand2 gate1592(.a(gate184inter8), .b(gate184inter7), .O(gate184inter9));
  nand2 gate1593(.a(s_149), .b(gate184inter3), .O(gate184inter10));
  nor2  gate1594(.a(gate184inter10), .b(gate184inter9), .O(gate184inter11));
  nor2  gate1595(.a(gate184inter11), .b(gate184inter6), .O(gate184inter12));
  nand2 gate1596(.a(gate184inter12), .b(gate184inter1), .O(G601));
nand2 gate185( .a(G570), .b(G571), .O(G602) );
nand2 gate186( .a(G572), .b(G573), .O(G607) );
nand2 gate187( .a(G574), .b(G575), .O(G612) );

  xor2  gate925(.a(G577), .b(G576), .O(gate188inter0));
  nand2 gate926(.a(gate188inter0), .b(s_54), .O(gate188inter1));
  and2  gate927(.a(G577), .b(G576), .O(gate188inter2));
  inv1  gate928(.a(s_54), .O(gate188inter3));
  inv1  gate929(.a(s_55), .O(gate188inter4));
  nand2 gate930(.a(gate188inter4), .b(gate188inter3), .O(gate188inter5));
  nor2  gate931(.a(gate188inter5), .b(gate188inter2), .O(gate188inter6));
  inv1  gate932(.a(G576), .O(gate188inter7));
  inv1  gate933(.a(G577), .O(gate188inter8));
  nand2 gate934(.a(gate188inter8), .b(gate188inter7), .O(gate188inter9));
  nand2 gate935(.a(s_55), .b(gate188inter3), .O(gate188inter10));
  nor2  gate936(.a(gate188inter10), .b(gate188inter9), .O(gate188inter11));
  nor2  gate937(.a(gate188inter11), .b(gate188inter6), .O(gate188inter12));
  nand2 gate938(.a(gate188inter12), .b(gate188inter1), .O(G617));
nand2 gate189( .a(G578), .b(G579), .O(G622) );
nand2 gate190( .a(G580), .b(G581), .O(G627) );
nand2 gate191( .a(G582), .b(G583), .O(G632) );
nand2 gate192( .a(G584), .b(G585), .O(G637) );
nand2 gate193( .a(G586), .b(G587), .O(G642) );
nand2 gate194( .a(G588), .b(G589), .O(G645) );
nand2 gate195( .a(G590), .b(G591), .O(G648) );
nand2 gate196( .a(G592), .b(G593), .O(G651) );
nand2 gate197( .a(G594), .b(G595), .O(G654) );
nand2 gate198( .a(G596), .b(G597), .O(G657) );

  xor2  gate1023(.a(G599), .b(G598), .O(gate199inter0));
  nand2 gate1024(.a(gate199inter0), .b(s_68), .O(gate199inter1));
  and2  gate1025(.a(G599), .b(G598), .O(gate199inter2));
  inv1  gate1026(.a(s_68), .O(gate199inter3));
  inv1  gate1027(.a(s_69), .O(gate199inter4));
  nand2 gate1028(.a(gate199inter4), .b(gate199inter3), .O(gate199inter5));
  nor2  gate1029(.a(gate199inter5), .b(gate199inter2), .O(gate199inter6));
  inv1  gate1030(.a(G598), .O(gate199inter7));
  inv1  gate1031(.a(G599), .O(gate199inter8));
  nand2 gate1032(.a(gate199inter8), .b(gate199inter7), .O(gate199inter9));
  nand2 gate1033(.a(s_69), .b(gate199inter3), .O(gate199inter10));
  nor2  gate1034(.a(gate199inter10), .b(gate199inter9), .O(gate199inter11));
  nor2  gate1035(.a(gate199inter11), .b(gate199inter6), .O(gate199inter12));
  nand2 gate1036(.a(gate199inter12), .b(gate199inter1), .O(G660));
nand2 gate200( .a(G600), .b(G601), .O(G663) );
nand2 gate201( .a(G602), .b(G607), .O(G666) );
nand2 gate202( .a(G612), .b(G617), .O(G669) );
nand2 gate203( .a(G602), .b(G612), .O(G672) );
nand2 gate204( .a(G607), .b(G617), .O(G675) );
nand2 gate205( .a(G622), .b(G627), .O(G678) );
nand2 gate206( .a(G632), .b(G637), .O(G681) );
nand2 gate207( .a(G622), .b(G632), .O(G684) );
nand2 gate208( .a(G627), .b(G637), .O(G687) );
nand2 gate209( .a(G602), .b(G666), .O(G690) );
nand2 gate210( .a(G607), .b(G666), .O(G691) );
nand2 gate211( .a(G612), .b(G669), .O(G692) );

  xor2  gate715(.a(G669), .b(G617), .O(gate212inter0));
  nand2 gate716(.a(gate212inter0), .b(s_24), .O(gate212inter1));
  and2  gate717(.a(G669), .b(G617), .O(gate212inter2));
  inv1  gate718(.a(s_24), .O(gate212inter3));
  inv1  gate719(.a(s_25), .O(gate212inter4));
  nand2 gate720(.a(gate212inter4), .b(gate212inter3), .O(gate212inter5));
  nor2  gate721(.a(gate212inter5), .b(gate212inter2), .O(gate212inter6));
  inv1  gate722(.a(G617), .O(gate212inter7));
  inv1  gate723(.a(G669), .O(gate212inter8));
  nand2 gate724(.a(gate212inter8), .b(gate212inter7), .O(gate212inter9));
  nand2 gate725(.a(s_25), .b(gate212inter3), .O(gate212inter10));
  nor2  gate726(.a(gate212inter10), .b(gate212inter9), .O(gate212inter11));
  nor2  gate727(.a(gate212inter11), .b(gate212inter6), .O(gate212inter12));
  nand2 gate728(.a(gate212inter12), .b(gate212inter1), .O(G693));
nand2 gate213( .a(G602), .b(G672), .O(G694) );
nand2 gate214( .a(G612), .b(G672), .O(G695) );
nand2 gate215( .a(G607), .b(G675), .O(G696) );
nand2 gate216( .a(G617), .b(G675), .O(G697) );

  xor2  gate981(.a(G678), .b(G622), .O(gate217inter0));
  nand2 gate982(.a(gate217inter0), .b(s_62), .O(gate217inter1));
  and2  gate983(.a(G678), .b(G622), .O(gate217inter2));
  inv1  gate984(.a(s_62), .O(gate217inter3));
  inv1  gate985(.a(s_63), .O(gate217inter4));
  nand2 gate986(.a(gate217inter4), .b(gate217inter3), .O(gate217inter5));
  nor2  gate987(.a(gate217inter5), .b(gate217inter2), .O(gate217inter6));
  inv1  gate988(.a(G622), .O(gate217inter7));
  inv1  gate989(.a(G678), .O(gate217inter8));
  nand2 gate990(.a(gate217inter8), .b(gate217inter7), .O(gate217inter9));
  nand2 gate991(.a(s_63), .b(gate217inter3), .O(gate217inter10));
  nor2  gate992(.a(gate217inter10), .b(gate217inter9), .O(gate217inter11));
  nor2  gate993(.a(gate217inter11), .b(gate217inter6), .O(gate217inter12));
  nand2 gate994(.a(gate217inter12), .b(gate217inter1), .O(G698));
nand2 gate218( .a(G627), .b(G678), .O(G699) );
nand2 gate219( .a(G632), .b(G681), .O(G700) );
nand2 gate220( .a(G637), .b(G681), .O(G701) );
nand2 gate221( .a(G622), .b(G684), .O(G702) );
nand2 gate222( .a(G632), .b(G684), .O(G703) );

  xor2  gate645(.a(G687), .b(G627), .O(gate223inter0));
  nand2 gate646(.a(gate223inter0), .b(s_14), .O(gate223inter1));
  and2  gate647(.a(G687), .b(G627), .O(gate223inter2));
  inv1  gate648(.a(s_14), .O(gate223inter3));
  inv1  gate649(.a(s_15), .O(gate223inter4));
  nand2 gate650(.a(gate223inter4), .b(gate223inter3), .O(gate223inter5));
  nor2  gate651(.a(gate223inter5), .b(gate223inter2), .O(gate223inter6));
  inv1  gate652(.a(G627), .O(gate223inter7));
  inv1  gate653(.a(G687), .O(gate223inter8));
  nand2 gate654(.a(gate223inter8), .b(gate223inter7), .O(gate223inter9));
  nand2 gate655(.a(s_15), .b(gate223inter3), .O(gate223inter10));
  nor2  gate656(.a(gate223inter10), .b(gate223inter9), .O(gate223inter11));
  nor2  gate657(.a(gate223inter11), .b(gate223inter6), .O(gate223inter12));
  nand2 gate658(.a(gate223inter12), .b(gate223inter1), .O(G704));
nand2 gate224( .a(G637), .b(G687), .O(G705) );
nand2 gate225( .a(G690), .b(G691), .O(G706) );
nand2 gate226( .a(G692), .b(G693), .O(G709) );
nand2 gate227( .a(G694), .b(G695), .O(G712) );
nand2 gate228( .a(G696), .b(G697), .O(G715) );
nand2 gate229( .a(G698), .b(G699), .O(G718) );
nand2 gate230( .a(G700), .b(G701), .O(G721) );
nand2 gate231( .a(G702), .b(G703), .O(G724) );

  xor2  gate1569(.a(G705), .b(G704), .O(gate232inter0));
  nand2 gate1570(.a(gate232inter0), .b(s_146), .O(gate232inter1));
  and2  gate1571(.a(G705), .b(G704), .O(gate232inter2));
  inv1  gate1572(.a(s_146), .O(gate232inter3));
  inv1  gate1573(.a(s_147), .O(gate232inter4));
  nand2 gate1574(.a(gate232inter4), .b(gate232inter3), .O(gate232inter5));
  nor2  gate1575(.a(gate232inter5), .b(gate232inter2), .O(gate232inter6));
  inv1  gate1576(.a(G704), .O(gate232inter7));
  inv1  gate1577(.a(G705), .O(gate232inter8));
  nand2 gate1578(.a(gate232inter8), .b(gate232inter7), .O(gate232inter9));
  nand2 gate1579(.a(s_147), .b(gate232inter3), .O(gate232inter10));
  nor2  gate1580(.a(gate232inter10), .b(gate232inter9), .O(gate232inter11));
  nor2  gate1581(.a(gate232inter11), .b(gate232inter6), .O(gate232inter12));
  nand2 gate1582(.a(gate232inter12), .b(gate232inter1), .O(G727));
nand2 gate233( .a(G242), .b(G718), .O(G730) );
nand2 gate234( .a(G245), .b(G721), .O(G733) );
nand2 gate235( .a(G248), .b(G724), .O(G736) );
nand2 gate236( .a(G251), .b(G727), .O(G739) );
nand2 gate237( .a(G254), .b(G706), .O(G742) );
nand2 gate238( .a(G257), .b(G709), .O(G745) );
nand2 gate239( .a(G260), .b(G712), .O(G748) );
nand2 gate240( .a(G263), .b(G715), .O(G751) );
nand2 gate241( .a(G242), .b(G730), .O(G754) );
nand2 gate242( .a(G718), .b(G730), .O(G755) );
nand2 gate243( .a(G245), .b(G733), .O(G756) );
nand2 gate244( .a(G721), .b(G733), .O(G757) );
nand2 gate245( .a(G248), .b(G736), .O(G758) );
nand2 gate246( .a(G724), .b(G736), .O(G759) );
nand2 gate247( .a(G251), .b(G739), .O(G760) );
nand2 gate248( .a(G727), .b(G739), .O(G761) );
nand2 gate249( .a(G254), .b(G742), .O(G762) );
nand2 gate250( .a(G706), .b(G742), .O(G763) );
nand2 gate251( .a(G257), .b(G745), .O(G764) );
nand2 gate252( .a(G709), .b(G745), .O(G765) );
nand2 gate253( .a(G260), .b(G748), .O(G766) );
nand2 gate254( .a(G712), .b(G748), .O(G767) );
nand2 gate255( .a(G263), .b(G751), .O(G768) );
nand2 gate256( .a(G715), .b(G751), .O(G769) );
nand2 gate257( .a(G754), .b(G755), .O(G770) );
nand2 gate258( .a(G756), .b(G757), .O(G773) );
nand2 gate259( .a(G758), .b(G759), .O(G776) );
nand2 gate260( .a(G760), .b(G761), .O(G779) );
nand2 gate261( .a(G762), .b(G763), .O(G782) );
nand2 gate262( .a(G764), .b(G765), .O(G785) );
nand2 gate263( .a(G766), .b(G767), .O(G788) );
nand2 gate264( .a(G768), .b(G769), .O(G791) );
nand2 gate265( .a(G642), .b(G770), .O(G794) );
nand2 gate266( .a(G645), .b(G773), .O(G797) );
nand2 gate267( .a(G648), .b(G776), .O(G800) );
nand2 gate268( .a(G651), .b(G779), .O(G803) );
nand2 gate269( .a(G654), .b(G782), .O(G806) );
nand2 gate270( .a(G657), .b(G785), .O(G809) );
nand2 gate271( .a(G660), .b(G788), .O(G812) );
nand2 gate272( .a(G663), .b(G791), .O(G815) );
nand2 gate273( .a(G642), .b(G794), .O(G818) );

  xor2  gate869(.a(G794), .b(G770), .O(gate274inter0));
  nand2 gate870(.a(gate274inter0), .b(s_46), .O(gate274inter1));
  and2  gate871(.a(G794), .b(G770), .O(gate274inter2));
  inv1  gate872(.a(s_46), .O(gate274inter3));
  inv1  gate873(.a(s_47), .O(gate274inter4));
  nand2 gate874(.a(gate274inter4), .b(gate274inter3), .O(gate274inter5));
  nor2  gate875(.a(gate274inter5), .b(gate274inter2), .O(gate274inter6));
  inv1  gate876(.a(G770), .O(gate274inter7));
  inv1  gate877(.a(G794), .O(gate274inter8));
  nand2 gate878(.a(gate274inter8), .b(gate274inter7), .O(gate274inter9));
  nand2 gate879(.a(s_47), .b(gate274inter3), .O(gate274inter10));
  nor2  gate880(.a(gate274inter10), .b(gate274inter9), .O(gate274inter11));
  nor2  gate881(.a(gate274inter11), .b(gate274inter6), .O(gate274inter12));
  nand2 gate882(.a(gate274inter12), .b(gate274inter1), .O(G819));
nand2 gate275( .a(G645), .b(G797), .O(G820) );

  xor2  gate729(.a(G797), .b(G773), .O(gate276inter0));
  nand2 gate730(.a(gate276inter0), .b(s_26), .O(gate276inter1));
  and2  gate731(.a(G797), .b(G773), .O(gate276inter2));
  inv1  gate732(.a(s_26), .O(gate276inter3));
  inv1  gate733(.a(s_27), .O(gate276inter4));
  nand2 gate734(.a(gate276inter4), .b(gate276inter3), .O(gate276inter5));
  nor2  gate735(.a(gate276inter5), .b(gate276inter2), .O(gate276inter6));
  inv1  gate736(.a(G773), .O(gate276inter7));
  inv1  gate737(.a(G797), .O(gate276inter8));
  nand2 gate738(.a(gate276inter8), .b(gate276inter7), .O(gate276inter9));
  nand2 gate739(.a(s_27), .b(gate276inter3), .O(gate276inter10));
  nor2  gate740(.a(gate276inter10), .b(gate276inter9), .O(gate276inter11));
  nor2  gate741(.a(gate276inter11), .b(gate276inter6), .O(gate276inter12));
  nand2 gate742(.a(gate276inter12), .b(gate276inter1), .O(G821));
nand2 gate277( .a(G648), .b(G800), .O(G822) );
nand2 gate278( .a(G776), .b(G800), .O(G823) );
nand2 gate279( .a(G651), .b(G803), .O(G824) );
nand2 gate280( .a(G779), .b(G803), .O(G825) );
nand2 gate281( .a(G654), .b(G806), .O(G826) );
nand2 gate282( .a(G782), .b(G806), .O(G827) );
nand2 gate283( .a(G657), .b(G809), .O(G828) );

  xor2  gate757(.a(G809), .b(G785), .O(gate284inter0));
  nand2 gate758(.a(gate284inter0), .b(s_30), .O(gate284inter1));
  and2  gate759(.a(G809), .b(G785), .O(gate284inter2));
  inv1  gate760(.a(s_30), .O(gate284inter3));
  inv1  gate761(.a(s_31), .O(gate284inter4));
  nand2 gate762(.a(gate284inter4), .b(gate284inter3), .O(gate284inter5));
  nor2  gate763(.a(gate284inter5), .b(gate284inter2), .O(gate284inter6));
  inv1  gate764(.a(G785), .O(gate284inter7));
  inv1  gate765(.a(G809), .O(gate284inter8));
  nand2 gate766(.a(gate284inter8), .b(gate284inter7), .O(gate284inter9));
  nand2 gate767(.a(s_31), .b(gate284inter3), .O(gate284inter10));
  nor2  gate768(.a(gate284inter10), .b(gate284inter9), .O(gate284inter11));
  nor2  gate769(.a(gate284inter11), .b(gate284inter6), .O(gate284inter12));
  nand2 gate770(.a(gate284inter12), .b(gate284inter1), .O(G829));

  xor2  gate1527(.a(G812), .b(G660), .O(gate285inter0));
  nand2 gate1528(.a(gate285inter0), .b(s_140), .O(gate285inter1));
  and2  gate1529(.a(G812), .b(G660), .O(gate285inter2));
  inv1  gate1530(.a(s_140), .O(gate285inter3));
  inv1  gate1531(.a(s_141), .O(gate285inter4));
  nand2 gate1532(.a(gate285inter4), .b(gate285inter3), .O(gate285inter5));
  nor2  gate1533(.a(gate285inter5), .b(gate285inter2), .O(gate285inter6));
  inv1  gate1534(.a(G660), .O(gate285inter7));
  inv1  gate1535(.a(G812), .O(gate285inter8));
  nand2 gate1536(.a(gate285inter8), .b(gate285inter7), .O(gate285inter9));
  nand2 gate1537(.a(s_141), .b(gate285inter3), .O(gate285inter10));
  nor2  gate1538(.a(gate285inter10), .b(gate285inter9), .O(gate285inter11));
  nor2  gate1539(.a(gate285inter11), .b(gate285inter6), .O(gate285inter12));
  nand2 gate1540(.a(gate285inter12), .b(gate285inter1), .O(G830));
nand2 gate286( .a(G788), .b(G812), .O(G831) );
nand2 gate287( .a(G663), .b(G815), .O(G832) );
nand2 gate288( .a(G791), .b(G815), .O(G833) );
nand2 gate289( .a(G818), .b(G819), .O(G834) );
nand2 gate290( .a(G820), .b(G821), .O(G847) );

  xor2  gate1177(.a(G823), .b(G822), .O(gate291inter0));
  nand2 gate1178(.a(gate291inter0), .b(s_90), .O(gate291inter1));
  and2  gate1179(.a(G823), .b(G822), .O(gate291inter2));
  inv1  gate1180(.a(s_90), .O(gate291inter3));
  inv1  gate1181(.a(s_91), .O(gate291inter4));
  nand2 gate1182(.a(gate291inter4), .b(gate291inter3), .O(gate291inter5));
  nor2  gate1183(.a(gate291inter5), .b(gate291inter2), .O(gate291inter6));
  inv1  gate1184(.a(G822), .O(gate291inter7));
  inv1  gate1185(.a(G823), .O(gate291inter8));
  nand2 gate1186(.a(gate291inter8), .b(gate291inter7), .O(gate291inter9));
  nand2 gate1187(.a(s_91), .b(gate291inter3), .O(gate291inter10));
  nor2  gate1188(.a(gate291inter10), .b(gate291inter9), .O(gate291inter11));
  nor2  gate1189(.a(gate291inter11), .b(gate291inter6), .O(gate291inter12));
  nand2 gate1190(.a(gate291inter12), .b(gate291inter1), .O(G860));

  xor2  gate799(.a(G825), .b(G824), .O(gate292inter0));
  nand2 gate800(.a(gate292inter0), .b(s_36), .O(gate292inter1));
  and2  gate801(.a(G825), .b(G824), .O(gate292inter2));
  inv1  gate802(.a(s_36), .O(gate292inter3));
  inv1  gate803(.a(s_37), .O(gate292inter4));
  nand2 gate804(.a(gate292inter4), .b(gate292inter3), .O(gate292inter5));
  nor2  gate805(.a(gate292inter5), .b(gate292inter2), .O(gate292inter6));
  inv1  gate806(.a(G824), .O(gate292inter7));
  inv1  gate807(.a(G825), .O(gate292inter8));
  nand2 gate808(.a(gate292inter8), .b(gate292inter7), .O(gate292inter9));
  nand2 gate809(.a(s_37), .b(gate292inter3), .O(gate292inter10));
  nor2  gate810(.a(gate292inter10), .b(gate292inter9), .O(gate292inter11));
  nor2  gate811(.a(gate292inter11), .b(gate292inter6), .O(gate292inter12));
  nand2 gate812(.a(gate292inter12), .b(gate292inter1), .O(G873));
nand2 gate293( .a(G828), .b(G829), .O(G886) );

  xor2  gate995(.a(G833), .b(G832), .O(gate294inter0));
  nand2 gate996(.a(gate294inter0), .b(s_64), .O(gate294inter1));
  and2  gate997(.a(G833), .b(G832), .O(gate294inter2));
  inv1  gate998(.a(s_64), .O(gate294inter3));
  inv1  gate999(.a(s_65), .O(gate294inter4));
  nand2 gate1000(.a(gate294inter4), .b(gate294inter3), .O(gate294inter5));
  nor2  gate1001(.a(gate294inter5), .b(gate294inter2), .O(gate294inter6));
  inv1  gate1002(.a(G832), .O(gate294inter7));
  inv1  gate1003(.a(G833), .O(gate294inter8));
  nand2 gate1004(.a(gate294inter8), .b(gate294inter7), .O(gate294inter9));
  nand2 gate1005(.a(s_65), .b(gate294inter3), .O(gate294inter10));
  nor2  gate1006(.a(gate294inter10), .b(gate294inter9), .O(gate294inter11));
  nor2  gate1007(.a(gate294inter11), .b(gate294inter6), .O(gate294inter12));
  nand2 gate1008(.a(gate294inter12), .b(gate294inter1), .O(G899));
nand2 gate295( .a(G830), .b(G831), .O(G912) );
nand2 gate296( .a(G826), .b(G827), .O(G925) );
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );
nand2 gate387( .a(G1), .b(G1036), .O(G1132) );
nand2 gate388( .a(G2), .b(G1039), .O(G1135) );
nand2 gate389( .a(G3), .b(G1042), .O(G1138) );
nand2 gate390( .a(G4), .b(G1045), .O(G1141) );
nand2 gate391( .a(G5), .b(G1048), .O(G1144) );
nand2 gate392( .a(G6), .b(G1051), .O(G1147) );

  xor2  gate1009(.a(G1054), .b(G7), .O(gate393inter0));
  nand2 gate1010(.a(gate393inter0), .b(s_66), .O(gate393inter1));
  and2  gate1011(.a(G1054), .b(G7), .O(gate393inter2));
  inv1  gate1012(.a(s_66), .O(gate393inter3));
  inv1  gate1013(.a(s_67), .O(gate393inter4));
  nand2 gate1014(.a(gate393inter4), .b(gate393inter3), .O(gate393inter5));
  nor2  gate1015(.a(gate393inter5), .b(gate393inter2), .O(gate393inter6));
  inv1  gate1016(.a(G7), .O(gate393inter7));
  inv1  gate1017(.a(G1054), .O(gate393inter8));
  nand2 gate1018(.a(gate393inter8), .b(gate393inter7), .O(gate393inter9));
  nand2 gate1019(.a(s_67), .b(gate393inter3), .O(gate393inter10));
  nor2  gate1020(.a(gate393inter10), .b(gate393inter9), .O(gate393inter11));
  nor2  gate1021(.a(gate393inter11), .b(gate393inter6), .O(gate393inter12));
  nand2 gate1022(.a(gate393inter12), .b(gate393inter1), .O(G1150));
nand2 gate394( .a(G8), .b(G1057), .O(G1153) );
nand2 gate395( .a(G9), .b(G1060), .O(G1156) );
nand2 gate396( .a(G10), .b(G1063), .O(G1159) );

  xor2  gate1443(.a(G1066), .b(G11), .O(gate397inter0));
  nand2 gate1444(.a(gate397inter0), .b(s_128), .O(gate397inter1));
  and2  gate1445(.a(G1066), .b(G11), .O(gate397inter2));
  inv1  gate1446(.a(s_128), .O(gate397inter3));
  inv1  gate1447(.a(s_129), .O(gate397inter4));
  nand2 gate1448(.a(gate397inter4), .b(gate397inter3), .O(gate397inter5));
  nor2  gate1449(.a(gate397inter5), .b(gate397inter2), .O(gate397inter6));
  inv1  gate1450(.a(G11), .O(gate397inter7));
  inv1  gate1451(.a(G1066), .O(gate397inter8));
  nand2 gate1452(.a(gate397inter8), .b(gate397inter7), .O(gate397inter9));
  nand2 gate1453(.a(s_129), .b(gate397inter3), .O(gate397inter10));
  nor2  gate1454(.a(gate397inter10), .b(gate397inter9), .O(gate397inter11));
  nor2  gate1455(.a(gate397inter11), .b(gate397inter6), .O(gate397inter12));
  nand2 gate1456(.a(gate397inter12), .b(gate397inter1), .O(G1162));
nand2 gate398( .a(G12), .b(G1069), .O(G1165) );
nand2 gate399( .a(G13), .b(G1072), .O(G1168) );
nand2 gate400( .a(G14), .b(G1075), .O(G1171) );
nand2 gate401( .a(G15), .b(G1078), .O(G1174) );
nand2 gate402( .a(G16), .b(G1081), .O(G1177) );
nand2 gate403( .a(G17), .b(G1084), .O(G1180) );
nand2 gate404( .a(G18), .b(G1087), .O(G1183) );
nand2 gate405( .a(G19), .b(G1090), .O(G1186) );
nand2 gate406( .a(G20), .b(G1093), .O(G1189) );
nand2 gate407( .a(G21), .b(G1096), .O(G1192) );
nand2 gate408( .a(G22), .b(G1099), .O(G1195) );
nand2 gate409( .a(G23), .b(G1102), .O(G1198) );
nand2 gate410( .a(G24), .b(G1105), .O(G1201) );
nand2 gate411( .a(G25), .b(G1108), .O(G1204) );
nand2 gate412( .a(G26), .b(G1111), .O(G1207) );
nand2 gate413( .a(G27), .b(G1114), .O(G1210) );
nand2 gate414( .a(G28), .b(G1117), .O(G1213) );
nand2 gate415( .a(G29), .b(G1120), .O(G1216) );
nand2 gate416( .a(G30), .b(G1123), .O(G1219) );
nand2 gate417( .a(G31), .b(G1126), .O(G1222) );
nand2 gate418( .a(G32), .b(G1129), .O(G1225) );
nand2 gate419( .a(G1), .b(G1132), .O(G1228) );
nand2 gate420( .a(G1036), .b(G1132), .O(G1229) );
nand2 gate421( .a(G2), .b(G1135), .O(G1230) );
nand2 gate422( .a(G1039), .b(G1135), .O(G1231) );

  xor2  gate1303(.a(G1138), .b(G3), .O(gate423inter0));
  nand2 gate1304(.a(gate423inter0), .b(s_108), .O(gate423inter1));
  and2  gate1305(.a(G1138), .b(G3), .O(gate423inter2));
  inv1  gate1306(.a(s_108), .O(gate423inter3));
  inv1  gate1307(.a(s_109), .O(gate423inter4));
  nand2 gate1308(.a(gate423inter4), .b(gate423inter3), .O(gate423inter5));
  nor2  gate1309(.a(gate423inter5), .b(gate423inter2), .O(gate423inter6));
  inv1  gate1310(.a(G3), .O(gate423inter7));
  inv1  gate1311(.a(G1138), .O(gate423inter8));
  nand2 gate1312(.a(gate423inter8), .b(gate423inter7), .O(gate423inter9));
  nand2 gate1313(.a(s_109), .b(gate423inter3), .O(gate423inter10));
  nor2  gate1314(.a(gate423inter10), .b(gate423inter9), .O(gate423inter11));
  nor2  gate1315(.a(gate423inter11), .b(gate423inter6), .O(gate423inter12));
  nand2 gate1316(.a(gate423inter12), .b(gate423inter1), .O(G1232));
nand2 gate424( .a(G1042), .b(G1138), .O(G1233) );
nand2 gate425( .a(G4), .b(G1141), .O(G1234) );
nand2 gate426( .a(G1045), .b(G1141), .O(G1235) );
nand2 gate427( .a(G5), .b(G1144), .O(G1236) );
nand2 gate428( .a(G1048), .b(G1144), .O(G1237) );
nand2 gate429( .a(G6), .b(G1147), .O(G1238) );
nand2 gate430( .a(G1051), .b(G1147), .O(G1239) );
nand2 gate431( .a(G7), .b(G1150), .O(G1240) );
nand2 gate432( .a(G1054), .b(G1150), .O(G1241) );

  xor2  gate701(.a(G1153), .b(G8), .O(gate433inter0));
  nand2 gate702(.a(gate433inter0), .b(s_22), .O(gate433inter1));
  and2  gate703(.a(G1153), .b(G8), .O(gate433inter2));
  inv1  gate704(.a(s_22), .O(gate433inter3));
  inv1  gate705(.a(s_23), .O(gate433inter4));
  nand2 gate706(.a(gate433inter4), .b(gate433inter3), .O(gate433inter5));
  nor2  gate707(.a(gate433inter5), .b(gate433inter2), .O(gate433inter6));
  inv1  gate708(.a(G8), .O(gate433inter7));
  inv1  gate709(.a(G1153), .O(gate433inter8));
  nand2 gate710(.a(gate433inter8), .b(gate433inter7), .O(gate433inter9));
  nand2 gate711(.a(s_23), .b(gate433inter3), .O(gate433inter10));
  nor2  gate712(.a(gate433inter10), .b(gate433inter9), .O(gate433inter11));
  nor2  gate713(.a(gate433inter11), .b(gate433inter6), .O(gate433inter12));
  nand2 gate714(.a(gate433inter12), .b(gate433inter1), .O(G1242));
nand2 gate434( .a(G1057), .b(G1153), .O(G1243) );

  xor2  gate897(.a(G1156), .b(G9), .O(gate435inter0));
  nand2 gate898(.a(gate435inter0), .b(s_50), .O(gate435inter1));
  and2  gate899(.a(G1156), .b(G9), .O(gate435inter2));
  inv1  gate900(.a(s_50), .O(gate435inter3));
  inv1  gate901(.a(s_51), .O(gate435inter4));
  nand2 gate902(.a(gate435inter4), .b(gate435inter3), .O(gate435inter5));
  nor2  gate903(.a(gate435inter5), .b(gate435inter2), .O(gate435inter6));
  inv1  gate904(.a(G9), .O(gate435inter7));
  inv1  gate905(.a(G1156), .O(gate435inter8));
  nand2 gate906(.a(gate435inter8), .b(gate435inter7), .O(gate435inter9));
  nand2 gate907(.a(s_51), .b(gate435inter3), .O(gate435inter10));
  nor2  gate908(.a(gate435inter10), .b(gate435inter9), .O(gate435inter11));
  nor2  gate909(.a(gate435inter11), .b(gate435inter6), .O(gate435inter12));
  nand2 gate910(.a(gate435inter12), .b(gate435inter1), .O(G1244));

  xor2  gate575(.a(G1156), .b(G1060), .O(gate436inter0));
  nand2 gate576(.a(gate436inter0), .b(s_4), .O(gate436inter1));
  and2  gate577(.a(G1156), .b(G1060), .O(gate436inter2));
  inv1  gate578(.a(s_4), .O(gate436inter3));
  inv1  gate579(.a(s_5), .O(gate436inter4));
  nand2 gate580(.a(gate436inter4), .b(gate436inter3), .O(gate436inter5));
  nor2  gate581(.a(gate436inter5), .b(gate436inter2), .O(gate436inter6));
  inv1  gate582(.a(G1060), .O(gate436inter7));
  inv1  gate583(.a(G1156), .O(gate436inter8));
  nand2 gate584(.a(gate436inter8), .b(gate436inter7), .O(gate436inter9));
  nand2 gate585(.a(s_5), .b(gate436inter3), .O(gate436inter10));
  nor2  gate586(.a(gate436inter10), .b(gate436inter9), .O(gate436inter11));
  nor2  gate587(.a(gate436inter11), .b(gate436inter6), .O(gate436inter12));
  nand2 gate588(.a(gate436inter12), .b(gate436inter1), .O(G1245));
nand2 gate437( .a(G10), .b(G1159), .O(G1246) );
nand2 gate438( .a(G1063), .b(G1159), .O(G1247) );

  xor2  gate1275(.a(G1162), .b(G11), .O(gate439inter0));
  nand2 gate1276(.a(gate439inter0), .b(s_104), .O(gate439inter1));
  and2  gate1277(.a(G1162), .b(G11), .O(gate439inter2));
  inv1  gate1278(.a(s_104), .O(gate439inter3));
  inv1  gate1279(.a(s_105), .O(gate439inter4));
  nand2 gate1280(.a(gate439inter4), .b(gate439inter3), .O(gate439inter5));
  nor2  gate1281(.a(gate439inter5), .b(gate439inter2), .O(gate439inter6));
  inv1  gate1282(.a(G11), .O(gate439inter7));
  inv1  gate1283(.a(G1162), .O(gate439inter8));
  nand2 gate1284(.a(gate439inter8), .b(gate439inter7), .O(gate439inter9));
  nand2 gate1285(.a(s_105), .b(gate439inter3), .O(gate439inter10));
  nor2  gate1286(.a(gate439inter10), .b(gate439inter9), .O(gate439inter11));
  nor2  gate1287(.a(gate439inter11), .b(gate439inter6), .O(gate439inter12));
  nand2 gate1288(.a(gate439inter12), .b(gate439inter1), .O(G1248));
nand2 gate440( .a(G1066), .b(G1162), .O(G1249) );

  xor2  gate1093(.a(G1165), .b(G12), .O(gate441inter0));
  nand2 gate1094(.a(gate441inter0), .b(s_78), .O(gate441inter1));
  and2  gate1095(.a(G1165), .b(G12), .O(gate441inter2));
  inv1  gate1096(.a(s_78), .O(gate441inter3));
  inv1  gate1097(.a(s_79), .O(gate441inter4));
  nand2 gate1098(.a(gate441inter4), .b(gate441inter3), .O(gate441inter5));
  nor2  gate1099(.a(gate441inter5), .b(gate441inter2), .O(gate441inter6));
  inv1  gate1100(.a(G12), .O(gate441inter7));
  inv1  gate1101(.a(G1165), .O(gate441inter8));
  nand2 gate1102(.a(gate441inter8), .b(gate441inter7), .O(gate441inter9));
  nand2 gate1103(.a(s_79), .b(gate441inter3), .O(gate441inter10));
  nor2  gate1104(.a(gate441inter10), .b(gate441inter9), .O(gate441inter11));
  nor2  gate1105(.a(gate441inter11), .b(gate441inter6), .O(gate441inter12));
  nand2 gate1106(.a(gate441inter12), .b(gate441inter1), .O(G1250));
nand2 gate442( .a(G1069), .b(G1165), .O(G1251) );
nand2 gate443( .a(G13), .b(G1168), .O(G1252) );
nand2 gate444( .a(G1072), .b(G1168), .O(G1253) );
nand2 gate445( .a(G14), .b(G1171), .O(G1254) );
nand2 gate446( .a(G1075), .b(G1171), .O(G1255) );
nand2 gate447( .a(G15), .b(G1174), .O(G1256) );

  xor2  gate1415(.a(G1174), .b(G1078), .O(gate448inter0));
  nand2 gate1416(.a(gate448inter0), .b(s_124), .O(gate448inter1));
  and2  gate1417(.a(G1174), .b(G1078), .O(gate448inter2));
  inv1  gate1418(.a(s_124), .O(gate448inter3));
  inv1  gate1419(.a(s_125), .O(gate448inter4));
  nand2 gate1420(.a(gate448inter4), .b(gate448inter3), .O(gate448inter5));
  nor2  gate1421(.a(gate448inter5), .b(gate448inter2), .O(gate448inter6));
  inv1  gate1422(.a(G1078), .O(gate448inter7));
  inv1  gate1423(.a(G1174), .O(gate448inter8));
  nand2 gate1424(.a(gate448inter8), .b(gate448inter7), .O(gate448inter9));
  nand2 gate1425(.a(s_125), .b(gate448inter3), .O(gate448inter10));
  nor2  gate1426(.a(gate448inter10), .b(gate448inter9), .O(gate448inter11));
  nor2  gate1427(.a(gate448inter11), .b(gate448inter6), .O(gate448inter12));
  nand2 gate1428(.a(gate448inter12), .b(gate448inter1), .O(G1257));
nand2 gate449( .a(G16), .b(G1177), .O(G1258) );
nand2 gate450( .a(G1081), .b(G1177), .O(G1259) );

  xor2  gate953(.a(G1180), .b(G17), .O(gate451inter0));
  nand2 gate954(.a(gate451inter0), .b(s_58), .O(gate451inter1));
  and2  gate955(.a(G1180), .b(G17), .O(gate451inter2));
  inv1  gate956(.a(s_58), .O(gate451inter3));
  inv1  gate957(.a(s_59), .O(gate451inter4));
  nand2 gate958(.a(gate451inter4), .b(gate451inter3), .O(gate451inter5));
  nor2  gate959(.a(gate451inter5), .b(gate451inter2), .O(gate451inter6));
  inv1  gate960(.a(G17), .O(gate451inter7));
  inv1  gate961(.a(G1180), .O(gate451inter8));
  nand2 gate962(.a(gate451inter8), .b(gate451inter7), .O(gate451inter9));
  nand2 gate963(.a(s_59), .b(gate451inter3), .O(gate451inter10));
  nor2  gate964(.a(gate451inter10), .b(gate451inter9), .O(gate451inter11));
  nor2  gate965(.a(gate451inter11), .b(gate451inter6), .O(gate451inter12));
  nand2 gate966(.a(gate451inter12), .b(gate451inter1), .O(G1260));
nand2 gate452( .a(G1084), .b(G1180), .O(G1261) );
nand2 gate453( .a(G18), .b(G1183), .O(G1262) );
nand2 gate454( .a(G1087), .b(G1183), .O(G1263) );
nand2 gate455( .a(G19), .b(G1186), .O(G1264) );
nand2 gate456( .a(G1090), .b(G1186), .O(G1265) );

  xor2  gate1079(.a(G1189), .b(G20), .O(gate457inter0));
  nand2 gate1080(.a(gate457inter0), .b(s_76), .O(gate457inter1));
  and2  gate1081(.a(G1189), .b(G20), .O(gate457inter2));
  inv1  gate1082(.a(s_76), .O(gate457inter3));
  inv1  gate1083(.a(s_77), .O(gate457inter4));
  nand2 gate1084(.a(gate457inter4), .b(gate457inter3), .O(gate457inter5));
  nor2  gate1085(.a(gate457inter5), .b(gate457inter2), .O(gate457inter6));
  inv1  gate1086(.a(G20), .O(gate457inter7));
  inv1  gate1087(.a(G1189), .O(gate457inter8));
  nand2 gate1088(.a(gate457inter8), .b(gate457inter7), .O(gate457inter9));
  nand2 gate1089(.a(s_77), .b(gate457inter3), .O(gate457inter10));
  nor2  gate1090(.a(gate457inter10), .b(gate457inter9), .O(gate457inter11));
  nor2  gate1091(.a(gate457inter11), .b(gate457inter6), .O(gate457inter12));
  nand2 gate1092(.a(gate457inter12), .b(gate457inter1), .O(G1266));

  xor2  gate911(.a(G1189), .b(G1093), .O(gate458inter0));
  nand2 gate912(.a(gate458inter0), .b(s_52), .O(gate458inter1));
  and2  gate913(.a(G1189), .b(G1093), .O(gate458inter2));
  inv1  gate914(.a(s_52), .O(gate458inter3));
  inv1  gate915(.a(s_53), .O(gate458inter4));
  nand2 gate916(.a(gate458inter4), .b(gate458inter3), .O(gate458inter5));
  nor2  gate917(.a(gate458inter5), .b(gate458inter2), .O(gate458inter6));
  inv1  gate918(.a(G1093), .O(gate458inter7));
  inv1  gate919(.a(G1189), .O(gate458inter8));
  nand2 gate920(.a(gate458inter8), .b(gate458inter7), .O(gate458inter9));
  nand2 gate921(.a(s_53), .b(gate458inter3), .O(gate458inter10));
  nor2  gate922(.a(gate458inter10), .b(gate458inter9), .O(gate458inter11));
  nor2  gate923(.a(gate458inter11), .b(gate458inter6), .O(gate458inter12));
  nand2 gate924(.a(gate458inter12), .b(gate458inter1), .O(G1267));

  xor2  gate687(.a(G1192), .b(G21), .O(gate459inter0));
  nand2 gate688(.a(gate459inter0), .b(s_20), .O(gate459inter1));
  and2  gate689(.a(G1192), .b(G21), .O(gate459inter2));
  inv1  gate690(.a(s_20), .O(gate459inter3));
  inv1  gate691(.a(s_21), .O(gate459inter4));
  nand2 gate692(.a(gate459inter4), .b(gate459inter3), .O(gate459inter5));
  nor2  gate693(.a(gate459inter5), .b(gate459inter2), .O(gate459inter6));
  inv1  gate694(.a(G21), .O(gate459inter7));
  inv1  gate695(.a(G1192), .O(gate459inter8));
  nand2 gate696(.a(gate459inter8), .b(gate459inter7), .O(gate459inter9));
  nand2 gate697(.a(s_21), .b(gate459inter3), .O(gate459inter10));
  nor2  gate698(.a(gate459inter10), .b(gate459inter9), .O(gate459inter11));
  nor2  gate699(.a(gate459inter11), .b(gate459inter6), .O(gate459inter12));
  nand2 gate700(.a(gate459inter12), .b(gate459inter1), .O(G1268));

  xor2  gate1261(.a(G1192), .b(G1096), .O(gate460inter0));
  nand2 gate1262(.a(gate460inter0), .b(s_102), .O(gate460inter1));
  and2  gate1263(.a(G1192), .b(G1096), .O(gate460inter2));
  inv1  gate1264(.a(s_102), .O(gate460inter3));
  inv1  gate1265(.a(s_103), .O(gate460inter4));
  nand2 gate1266(.a(gate460inter4), .b(gate460inter3), .O(gate460inter5));
  nor2  gate1267(.a(gate460inter5), .b(gate460inter2), .O(gate460inter6));
  inv1  gate1268(.a(G1096), .O(gate460inter7));
  inv1  gate1269(.a(G1192), .O(gate460inter8));
  nand2 gate1270(.a(gate460inter8), .b(gate460inter7), .O(gate460inter9));
  nand2 gate1271(.a(s_103), .b(gate460inter3), .O(gate460inter10));
  nor2  gate1272(.a(gate460inter10), .b(gate460inter9), .O(gate460inter11));
  nor2  gate1273(.a(gate460inter11), .b(gate460inter6), .O(gate460inter12));
  nand2 gate1274(.a(gate460inter12), .b(gate460inter1), .O(G1269));
nand2 gate461( .a(G22), .b(G1195), .O(G1270) );

  xor2  gate659(.a(G1195), .b(G1099), .O(gate462inter0));
  nand2 gate660(.a(gate462inter0), .b(s_16), .O(gate462inter1));
  and2  gate661(.a(G1195), .b(G1099), .O(gate462inter2));
  inv1  gate662(.a(s_16), .O(gate462inter3));
  inv1  gate663(.a(s_17), .O(gate462inter4));
  nand2 gate664(.a(gate462inter4), .b(gate462inter3), .O(gate462inter5));
  nor2  gate665(.a(gate462inter5), .b(gate462inter2), .O(gate462inter6));
  inv1  gate666(.a(G1099), .O(gate462inter7));
  inv1  gate667(.a(G1195), .O(gate462inter8));
  nand2 gate668(.a(gate462inter8), .b(gate462inter7), .O(gate462inter9));
  nand2 gate669(.a(s_17), .b(gate462inter3), .O(gate462inter10));
  nor2  gate670(.a(gate462inter10), .b(gate462inter9), .O(gate462inter11));
  nor2  gate671(.a(gate462inter11), .b(gate462inter6), .O(gate462inter12));
  nand2 gate672(.a(gate462inter12), .b(gate462inter1), .O(G1271));
nand2 gate463( .a(G23), .b(G1198), .O(G1272) );

  xor2  gate561(.a(G1198), .b(G1102), .O(gate464inter0));
  nand2 gate562(.a(gate464inter0), .b(s_2), .O(gate464inter1));
  and2  gate563(.a(G1198), .b(G1102), .O(gate464inter2));
  inv1  gate564(.a(s_2), .O(gate464inter3));
  inv1  gate565(.a(s_3), .O(gate464inter4));
  nand2 gate566(.a(gate464inter4), .b(gate464inter3), .O(gate464inter5));
  nor2  gate567(.a(gate464inter5), .b(gate464inter2), .O(gate464inter6));
  inv1  gate568(.a(G1102), .O(gate464inter7));
  inv1  gate569(.a(G1198), .O(gate464inter8));
  nand2 gate570(.a(gate464inter8), .b(gate464inter7), .O(gate464inter9));
  nand2 gate571(.a(s_3), .b(gate464inter3), .O(gate464inter10));
  nor2  gate572(.a(gate464inter10), .b(gate464inter9), .O(gate464inter11));
  nor2  gate573(.a(gate464inter11), .b(gate464inter6), .O(gate464inter12));
  nand2 gate574(.a(gate464inter12), .b(gate464inter1), .O(G1273));
nand2 gate465( .a(G24), .b(G1201), .O(G1274) );
nand2 gate466( .a(G1105), .b(G1201), .O(G1275) );

  xor2  gate631(.a(G1204), .b(G25), .O(gate467inter0));
  nand2 gate632(.a(gate467inter0), .b(s_12), .O(gate467inter1));
  and2  gate633(.a(G1204), .b(G25), .O(gate467inter2));
  inv1  gate634(.a(s_12), .O(gate467inter3));
  inv1  gate635(.a(s_13), .O(gate467inter4));
  nand2 gate636(.a(gate467inter4), .b(gate467inter3), .O(gate467inter5));
  nor2  gate637(.a(gate467inter5), .b(gate467inter2), .O(gate467inter6));
  inv1  gate638(.a(G25), .O(gate467inter7));
  inv1  gate639(.a(G1204), .O(gate467inter8));
  nand2 gate640(.a(gate467inter8), .b(gate467inter7), .O(gate467inter9));
  nand2 gate641(.a(s_13), .b(gate467inter3), .O(gate467inter10));
  nor2  gate642(.a(gate467inter10), .b(gate467inter9), .O(gate467inter11));
  nor2  gate643(.a(gate467inter11), .b(gate467inter6), .O(gate467inter12));
  nand2 gate644(.a(gate467inter12), .b(gate467inter1), .O(G1276));
nand2 gate468( .a(G1108), .b(G1204), .O(G1277) );

  xor2  gate1121(.a(G1207), .b(G26), .O(gate469inter0));
  nand2 gate1122(.a(gate469inter0), .b(s_82), .O(gate469inter1));
  and2  gate1123(.a(G1207), .b(G26), .O(gate469inter2));
  inv1  gate1124(.a(s_82), .O(gate469inter3));
  inv1  gate1125(.a(s_83), .O(gate469inter4));
  nand2 gate1126(.a(gate469inter4), .b(gate469inter3), .O(gate469inter5));
  nor2  gate1127(.a(gate469inter5), .b(gate469inter2), .O(gate469inter6));
  inv1  gate1128(.a(G26), .O(gate469inter7));
  inv1  gate1129(.a(G1207), .O(gate469inter8));
  nand2 gate1130(.a(gate469inter8), .b(gate469inter7), .O(gate469inter9));
  nand2 gate1131(.a(s_83), .b(gate469inter3), .O(gate469inter10));
  nor2  gate1132(.a(gate469inter10), .b(gate469inter9), .O(gate469inter11));
  nor2  gate1133(.a(gate469inter11), .b(gate469inter6), .O(gate469inter12));
  nand2 gate1134(.a(gate469inter12), .b(gate469inter1), .O(G1278));
nand2 gate470( .a(G1111), .b(G1207), .O(G1279) );
nand2 gate471( .a(G27), .b(G1210), .O(G1280) );
nand2 gate472( .a(G1114), .b(G1210), .O(G1281) );
nand2 gate473( .a(G28), .b(G1213), .O(G1282) );
nand2 gate474( .a(G1117), .b(G1213), .O(G1283) );
nand2 gate475( .a(G29), .b(G1216), .O(G1284) );

  xor2  gate673(.a(G1216), .b(G1120), .O(gate476inter0));
  nand2 gate674(.a(gate476inter0), .b(s_18), .O(gate476inter1));
  and2  gate675(.a(G1216), .b(G1120), .O(gate476inter2));
  inv1  gate676(.a(s_18), .O(gate476inter3));
  inv1  gate677(.a(s_19), .O(gate476inter4));
  nand2 gate678(.a(gate476inter4), .b(gate476inter3), .O(gate476inter5));
  nor2  gate679(.a(gate476inter5), .b(gate476inter2), .O(gate476inter6));
  inv1  gate680(.a(G1120), .O(gate476inter7));
  inv1  gate681(.a(G1216), .O(gate476inter8));
  nand2 gate682(.a(gate476inter8), .b(gate476inter7), .O(gate476inter9));
  nand2 gate683(.a(s_19), .b(gate476inter3), .O(gate476inter10));
  nor2  gate684(.a(gate476inter10), .b(gate476inter9), .O(gate476inter11));
  nor2  gate685(.a(gate476inter11), .b(gate476inter6), .O(gate476inter12));
  nand2 gate686(.a(gate476inter12), .b(gate476inter1), .O(G1285));
nand2 gate477( .a(G30), .b(G1219), .O(G1286) );
nand2 gate478( .a(G1123), .b(G1219), .O(G1287) );
nand2 gate479( .a(G31), .b(G1222), .O(G1288) );
nand2 gate480( .a(G1126), .b(G1222), .O(G1289) );
nand2 gate481( .a(G32), .b(G1225), .O(G1290) );
nand2 gate482( .a(G1129), .b(G1225), .O(G1291) );
nand2 gate483( .a(G1228), .b(G1229), .O(G1292) );
nand2 gate484( .a(G1230), .b(G1231), .O(G1293) );
nand2 gate485( .a(G1232), .b(G1233), .O(G1294) );
nand2 gate486( .a(G1234), .b(G1235), .O(G1295) );
nand2 gate487( .a(G1236), .b(G1237), .O(G1296) );
nand2 gate488( .a(G1238), .b(G1239), .O(G1297) );
nand2 gate489( .a(G1240), .b(G1241), .O(G1298) );
nand2 gate490( .a(G1242), .b(G1243), .O(G1299) );
nand2 gate491( .a(G1244), .b(G1245), .O(G1300) );
nand2 gate492( .a(G1246), .b(G1247), .O(G1301) );
nand2 gate493( .a(G1248), .b(G1249), .O(G1302) );
nand2 gate494( .a(G1250), .b(G1251), .O(G1303) );
nand2 gate495( .a(G1252), .b(G1253), .O(G1304) );
nand2 gate496( .a(G1254), .b(G1255), .O(G1305) );
nand2 gate497( .a(G1256), .b(G1257), .O(G1306) );
nand2 gate498( .a(G1258), .b(G1259), .O(G1307) );
nand2 gate499( .a(G1260), .b(G1261), .O(G1308) );
nand2 gate500( .a(G1262), .b(G1263), .O(G1309) );

  xor2  gate1359(.a(G1265), .b(G1264), .O(gate501inter0));
  nand2 gate1360(.a(gate501inter0), .b(s_116), .O(gate501inter1));
  and2  gate1361(.a(G1265), .b(G1264), .O(gate501inter2));
  inv1  gate1362(.a(s_116), .O(gate501inter3));
  inv1  gate1363(.a(s_117), .O(gate501inter4));
  nand2 gate1364(.a(gate501inter4), .b(gate501inter3), .O(gate501inter5));
  nor2  gate1365(.a(gate501inter5), .b(gate501inter2), .O(gate501inter6));
  inv1  gate1366(.a(G1264), .O(gate501inter7));
  inv1  gate1367(.a(G1265), .O(gate501inter8));
  nand2 gate1368(.a(gate501inter8), .b(gate501inter7), .O(gate501inter9));
  nand2 gate1369(.a(s_117), .b(gate501inter3), .O(gate501inter10));
  nor2  gate1370(.a(gate501inter10), .b(gate501inter9), .O(gate501inter11));
  nor2  gate1371(.a(gate501inter11), .b(gate501inter6), .O(gate501inter12));
  nand2 gate1372(.a(gate501inter12), .b(gate501inter1), .O(G1310));
nand2 gate502( .a(G1266), .b(G1267), .O(G1311) );
nand2 gate503( .a(G1268), .b(G1269), .O(G1312) );
nand2 gate504( .a(G1270), .b(G1271), .O(G1313) );
nand2 gate505( .a(G1272), .b(G1273), .O(G1314) );

  xor2  gate1219(.a(G1275), .b(G1274), .O(gate506inter0));
  nand2 gate1220(.a(gate506inter0), .b(s_96), .O(gate506inter1));
  and2  gate1221(.a(G1275), .b(G1274), .O(gate506inter2));
  inv1  gate1222(.a(s_96), .O(gate506inter3));
  inv1  gate1223(.a(s_97), .O(gate506inter4));
  nand2 gate1224(.a(gate506inter4), .b(gate506inter3), .O(gate506inter5));
  nor2  gate1225(.a(gate506inter5), .b(gate506inter2), .O(gate506inter6));
  inv1  gate1226(.a(G1274), .O(gate506inter7));
  inv1  gate1227(.a(G1275), .O(gate506inter8));
  nand2 gate1228(.a(gate506inter8), .b(gate506inter7), .O(gate506inter9));
  nand2 gate1229(.a(s_97), .b(gate506inter3), .O(gate506inter10));
  nor2  gate1230(.a(gate506inter10), .b(gate506inter9), .O(gate506inter11));
  nor2  gate1231(.a(gate506inter11), .b(gate506inter6), .O(gate506inter12));
  nand2 gate1232(.a(gate506inter12), .b(gate506inter1), .O(G1315));
nand2 gate507( .a(G1276), .b(G1277), .O(G1316) );

  xor2  gate841(.a(G1279), .b(G1278), .O(gate508inter0));
  nand2 gate842(.a(gate508inter0), .b(s_42), .O(gate508inter1));
  and2  gate843(.a(G1279), .b(G1278), .O(gate508inter2));
  inv1  gate844(.a(s_42), .O(gate508inter3));
  inv1  gate845(.a(s_43), .O(gate508inter4));
  nand2 gate846(.a(gate508inter4), .b(gate508inter3), .O(gate508inter5));
  nor2  gate847(.a(gate508inter5), .b(gate508inter2), .O(gate508inter6));
  inv1  gate848(.a(G1278), .O(gate508inter7));
  inv1  gate849(.a(G1279), .O(gate508inter8));
  nand2 gate850(.a(gate508inter8), .b(gate508inter7), .O(gate508inter9));
  nand2 gate851(.a(s_43), .b(gate508inter3), .O(gate508inter10));
  nor2  gate852(.a(gate508inter10), .b(gate508inter9), .O(gate508inter11));
  nor2  gate853(.a(gate508inter11), .b(gate508inter6), .O(gate508inter12));
  nand2 gate854(.a(gate508inter12), .b(gate508inter1), .O(G1317));
nand2 gate509( .a(G1280), .b(G1281), .O(G1318) );

  xor2  gate1065(.a(G1283), .b(G1282), .O(gate510inter0));
  nand2 gate1066(.a(gate510inter0), .b(s_74), .O(gate510inter1));
  and2  gate1067(.a(G1283), .b(G1282), .O(gate510inter2));
  inv1  gate1068(.a(s_74), .O(gate510inter3));
  inv1  gate1069(.a(s_75), .O(gate510inter4));
  nand2 gate1070(.a(gate510inter4), .b(gate510inter3), .O(gate510inter5));
  nor2  gate1071(.a(gate510inter5), .b(gate510inter2), .O(gate510inter6));
  inv1  gate1072(.a(G1282), .O(gate510inter7));
  inv1  gate1073(.a(G1283), .O(gate510inter8));
  nand2 gate1074(.a(gate510inter8), .b(gate510inter7), .O(gate510inter9));
  nand2 gate1075(.a(s_75), .b(gate510inter3), .O(gate510inter10));
  nor2  gate1076(.a(gate510inter10), .b(gate510inter9), .O(gate510inter11));
  nor2  gate1077(.a(gate510inter11), .b(gate510inter6), .O(gate510inter12));
  nand2 gate1078(.a(gate510inter12), .b(gate510inter1), .O(G1319));
nand2 gate511( .a(G1284), .b(G1285), .O(G1320) );
nand2 gate512( .a(G1286), .b(G1287), .O(G1321) );
nand2 gate513( .a(G1288), .b(G1289), .O(G1322) );
nand2 gate514( .a(G1290), .b(G1291), .O(G1323) );
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule