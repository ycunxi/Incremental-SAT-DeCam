module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);

input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;//RE__PI;

input s_0,s_1;//RE__ALLOW(00,01,10,11);
input s_2,s_3;//RE__ALLOW(00,01,10,11);
input s_4,s_5;//RE__ALLOW(00,01,10,11);
input s_6,s_7;//RE__ALLOW(00,01,10,11);
input s_8,s_9;//RE__ALLOW(00,01,10,11);
input s_10,s_11;//RE__ALLOW(00,01,10,11);
input s_12,s_13;//RE__ALLOW(00,01,10,11);
input s_14,s_15;//RE__ALLOW(00,01,10,11);
input s_16,s_17;//RE__ALLOW(00,01,10,11);
input s_18,s_19;//RE__ALLOW(00,01,10,11);
input s_20,s_21;//RE__ALLOW(00,01,10,11);
input s_22,s_23;//RE__ALLOW(00,01,10,11);
input s_24,s_25;//RE__ALLOW(00,01,10,11);
input s_26,s_27;//RE__ALLOW(00,01,10,11);
input s_28,s_29;//RE__ALLOW(00,01,10,11);
input s_30,s_31;//RE__ALLOW(00,01,10,11);
input s_32,s_33;//RE__ALLOW(00,01,10,11);
input s_34,s_35;//RE__ALLOW(00,01,10,11);
input s_36,s_37;//RE__ALLOW(00,01,10,11);
input s_38,s_39;//RE__ALLOW(00,01,10,11);
input s_40,s_41;//RE__ALLOW(00,01,10,11);
input s_42,s_43;//RE__ALLOW(00,01,10,11);
input s_44,s_45;//RE__ALLOW(00,01,10,11);
input s_46,s_47;//RE__ALLOW(00,01,10,11);
input s_48,s_49;//RE__ALLOW(00,01,10,11);
input s_50,s_51;//RE__ALLOW(00,01,10,11);
input s_52,s_53;//RE__ALLOW(00,01,10,11);
input s_54,s_55;//RE__ALLOW(00,01,10,11);
input s_56,s_57;//RE__ALLOW(00,01,10,11);
input s_58,s_59;//RE__ALLOW(00,01,10,11);
input s_60,s_61;//RE__ALLOW(00,01,10,11);
input s_62,s_63;//RE__ALLOW(00,01,10,11);
input s_64,s_65;//RE__ALLOW(00,01,10,11);
input s_66,s_67;//RE__ALLOW(00,01,10,11);
input s_68,s_69;//RE__ALLOW(00,01,10,11);
input s_70,s_71;//RE__ALLOW(00,01,10,11);
input s_72,s_73;//RE__ALLOW(00,01,10,11);
input s_74,s_75;//RE__ALLOW(00,01,10,11);
input s_76,s_77;//RE__ALLOW(00,01,10,11);
input s_78,s_79;//RE__ALLOW(00,01,10,11);
input s_80,s_81;//RE__ALLOW(00,01,10,11);
input s_82,s_83;//RE__ALLOW(00,01,10,11);
input s_84,s_85;//RE__ALLOW(00,01,10,11);
input s_86,s_87;//RE__ALLOW(00,01,10,11);
input s_88,s_89;//RE__ALLOW(00,01,10,11);
input s_90,s_91;//RE__ALLOW(00,01,10,11);
input s_92,s_93;//RE__ALLOW(00,01,10,11);
input s_94,s_95;//RE__ALLOW(00,01,10,11);
input s_96,s_97;//RE__ALLOW(00,01,10,11);
input s_98,s_99;//RE__ALLOW(00,01,10,11);
input s_100,s_101;//RE__ALLOW(00,01,10,11);
input s_102,s_103;//RE__ALLOW(00,01,10,11);
input s_104,s_105;//RE__ALLOW(00,01,10,11);
input s_106,s_107;//RE__ALLOW(00,01,10,11);
input s_108,s_109;//RE__ALLOW(00,01,10,11);
input s_110,s_111;//RE__ALLOW(00,01,10,11);
input s_112,s_113;//RE__ALLOW(00,01,10,11);
input s_114,s_115;//RE__ALLOW(00,01,10,11);
input s_116,s_117;//RE__ALLOW(00,01,10,11);
input s_118,s_119;//RE__ALLOW(00,01,10,11);
input s_120,s_121;//RE__ALLOW(00,01,10,11);
input s_122,s_123;//RE__ALLOW(00,01,10,11);
input s_124,s_125;//RE__ALLOW(00,01,10,11);
input s_126,s_127;//RE__ALLOW(00,01,10,11);
input s_128,s_129;//RE__ALLOW(00,01,10,11);
input s_130,s_131;//RE__ALLOW(00,01,10,11);
input s_132,s_133;//RE__ALLOW(00,01,10,11);
input s_134,s_135;//RE__ALLOW(00,01,10,11);
input s_136,s_137;//RE__ALLOW(00,01,10,11);
input s_138,s_139;//RE__ALLOW(00,01,10,11);
input s_140,s_141;//RE__ALLOW(00,01,10,11);
input s_142,s_143;//RE__ALLOW(00,01,10,11);
input s_144,s_145;//RE__ALLOW(00,01,10,11);
input s_146,s_147;//RE__ALLOW(00,01,10,11);
input s_148,s_149;//RE__ALLOW(00,01,10,11);
input s_150,s_151;//RE__ALLOW(00,01,10,11);
input s_152,s_153;//RE__ALLOW(00,01,10,11);
input s_154,s_155;//RE__ALLOW(00,01,10,11);
input s_156,s_157;//RE__ALLOW(00,01,10,11);
input s_158,s_159;//RE__ALLOW(00,01,10,11);
input s_160,s_161;//RE__ALLOW(00,01,10,11);
input s_162,s_163;//RE__ALLOW(00,01,10,11);
input s_164,s_165;//RE__ALLOW(00,01,10,11);
input s_166,s_167;//RE__ALLOW(00,01,10,11);
input s_168,s_169;//RE__ALLOW(00,01,10,11);
input s_170,s_171;//RE__ALLOW(00,01,10,11);
input s_172,s_173;//RE__ALLOW(00,01,10,11);
input s_174,s_175;//RE__ALLOW(00,01,10,11);
input s_176,s_177;//RE__ALLOW(00,01,10,11);
input s_178,s_179;//RE__ALLOW(00,01,10,11);
input s_180,s_181;//RE__ALLOW(00,01,10,11);
input s_182,s_183;//RE__ALLOW(00,01,10,11);
input s_184,s_185;//RE__ALLOW(00,01,10,11);
input s_186,s_187;//RE__ALLOW(00,01,10,11);
input s_188,s_189;//RE__ALLOW(00,01,10,11);
input s_190,s_191;//RE__ALLOW(00,01,10,11);
input s_192,s_193;//RE__ALLOW(00,01,10,11);
input s_194,s_195;//RE__ALLOW(00,01,10,11);
input s_196,s_197;//RE__ALLOW(00,01,10,11);
input s_198,s_199;//RE__ALLOW(00,01,10,11);
input s_200,s_201;//RE__ALLOW(00,01,10,11);
input s_202,s_203;//RE__ALLOW(00,01,10,11);
input s_204,s_205;//RE__ALLOW(00,01,10,11);
input s_206,s_207;//RE__ALLOW(00,01,10,11);
input s_208,s_209;//RE__ALLOW(00,01,10,11);
input s_210,s_211;//RE__ALLOW(00,01,10,11);
input s_212,s_213;//RE__ALLOW(00,01,10,11);
input s_214,s_215;//RE__ALLOW(00,01,10,11);
input s_216,s_217;//RE__ALLOW(00,01,10,11);
input s_218,s_219;//RE__ALLOW(00,01,10,11);
input s_220,s_221;//RE__ALLOW(00,01,10,11);
input s_222,s_223;//RE__ALLOW(00,01,10,11);
input s_224,s_225;//RE__ALLOW(00,01,10,11);
input s_226,s_227;//RE__ALLOW(00,01,10,11);
input s_228,s_229;//RE__ALLOW(00,01,10,11);
input s_230,s_231;//RE__ALLOW(00,01,10,11);
input s_232,s_233;//RE__ALLOW(00,01,10,11);
input s_234,s_235;//RE__ALLOW(00,01,10,11);
input s_236,s_237;//RE__ALLOW(00,01,10,11);
input s_238,s_239;//RE__ALLOW(00,01,10,11);
input s_240,s_241;//RE__ALLOW(00,01,10,11);
input s_242,s_243;//RE__ALLOW(00,01,10,11);
input s_244,s_245;//RE__ALLOW(00,01,10,11);
input s_246,s_247;//RE__ALLOW(00,01,10,11);
input s_248,s_249;//RE__ALLOW(00,01,10,11);
input s_250,s_251;//RE__ALLOW(00,01,10,11);
input s_252,s_253;//RE__ALLOW(00,01,10,11);
input s_254,s_255;//RE__ALLOW(00,01,10,11);
input s_256,s_257;//RE__ALLOW(00,01,10,11);
input s_258,s_259;//RE__ALLOW(00,01,10,11);
input s_260,s_261;//RE__ALLOW(00,01,10,11);
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;

  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate465inter0, gate465inter1, gate465inter2, gate465inter3, gate465inter4, gate465inter5, gate465inter6, gate465inter7, gate465inter8, gate465inter9, gate465inter10, gate465inter11, gate465inter12, gate161inter0, gate161inter1, gate161inter2, gate161inter3, gate161inter4, gate161inter5, gate161inter6, gate161inter7, gate161inter8, gate161inter9, gate161inter10, gate161inter11, gate161inter12, gate450inter0, gate450inter1, gate450inter2, gate450inter3, gate450inter4, gate450inter5, gate450inter6, gate450inter7, gate450inter8, gate450inter9, gate450inter10, gate450inter11, gate450inter12, gate262inter0, gate262inter1, gate262inter2, gate262inter3, gate262inter4, gate262inter5, gate262inter6, gate262inter7, gate262inter8, gate262inter9, gate262inter10, gate262inter11, gate262inter12, gate464inter0, gate464inter1, gate464inter2, gate464inter3, gate464inter4, gate464inter5, gate464inter6, gate464inter7, gate464inter8, gate464inter9, gate464inter10, gate464inter11, gate464inter12, gate18inter0, gate18inter1, gate18inter2, gate18inter3, gate18inter4, gate18inter5, gate18inter6, gate18inter7, gate18inter8, gate18inter9, gate18inter10, gate18inter11, gate18inter12, gate432inter0, gate432inter1, gate432inter2, gate432inter3, gate432inter4, gate432inter5, gate432inter6, gate432inter7, gate432inter8, gate432inter9, gate432inter10, gate432inter11, gate432inter12, gate45inter0, gate45inter1, gate45inter2, gate45inter3, gate45inter4, gate45inter5, gate45inter6, gate45inter7, gate45inter8, gate45inter9, gate45inter10, gate45inter11, gate45inter12, gate148inter0, gate148inter1, gate148inter2, gate148inter3, gate148inter4, gate148inter5, gate148inter6, gate148inter7, gate148inter8, gate148inter9, gate148inter10, gate148inter11, gate148inter12, gate231inter0, gate231inter1, gate231inter2, gate231inter3, gate231inter4, gate231inter5, gate231inter6, gate231inter7, gate231inter8, gate231inter9, gate231inter10, gate231inter11, gate231inter12, gate187inter0, gate187inter1, gate187inter2, gate187inter3, gate187inter4, gate187inter5, gate187inter6, gate187inter7, gate187inter8, gate187inter9, gate187inter10, gate187inter11, gate187inter12, gate495inter0, gate495inter1, gate495inter2, gate495inter3, gate495inter4, gate495inter5, gate495inter6, gate495inter7, gate495inter8, gate495inter9, gate495inter10, gate495inter11, gate495inter12, gate95inter0, gate95inter1, gate95inter2, gate95inter3, gate95inter4, gate95inter5, gate95inter6, gate95inter7, gate95inter8, gate95inter9, gate95inter10, gate95inter11, gate95inter12, gate241inter0, gate241inter1, gate241inter2, gate241inter3, gate241inter4, gate241inter5, gate241inter6, gate241inter7, gate241inter8, gate241inter9, gate241inter10, gate241inter11, gate241inter12, gate236inter0, gate236inter1, gate236inter2, gate236inter3, gate236inter4, gate236inter5, gate236inter6, gate236inter7, gate236inter8, gate236inter9, gate236inter10, gate236inter11, gate236inter12, gate509inter0, gate509inter1, gate509inter2, gate509inter3, gate509inter4, gate509inter5, gate509inter6, gate509inter7, gate509inter8, gate509inter9, gate509inter10, gate509inter11, gate509inter12, gate153inter0, gate153inter1, gate153inter2, gate153inter3, gate153inter4, gate153inter5, gate153inter6, gate153inter7, gate153inter8, gate153inter9, gate153inter10, gate153inter11, gate153inter12, gate41inter0, gate41inter1, gate41inter2, gate41inter3, gate41inter4, gate41inter5, gate41inter6, gate41inter7, gate41inter8, gate41inter9, gate41inter10, gate41inter11, gate41inter12, gate189inter0, gate189inter1, gate189inter2, gate189inter3, gate189inter4, gate189inter5, gate189inter6, gate189inter7, gate189inter8, gate189inter9, gate189inter10, gate189inter11, gate189inter12, gate68inter0, gate68inter1, gate68inter2, gate68inter3, gate68inter4, gate68inter5, gate68inter6, gate68inter7, gate68inter8, gate68inter9, gate68inter10, gate68inter11, gate68inter12, gate426inter0, gate426inter1, gate426inter2, gate426inter3, gate426inter4, gate426inter5, gate426inter6, gate426inter7, gate426inter8, gate426inter9, gate426inter10, gate426inter11, gate426inter12, gate407inter0, gate407inter1, gate407inter2, gate407inter3, gate407inter4, gate407inter5, gate407inter6, gate407inter7, gate407inter8, gate407inter9, gate407inter10, gate407inter11, gate407inter12, gate497inter0, gate497inter1, gate497inter2, gate497inter3, gate497inter4, gate497inter5, gate497inter6, gate497inter7, gate497inter8, gate497inter9, gate497inter10, gate497inter11, gate497inter12, gate446inter0, gate446inter1, gate446inter2, gate446inter3, gate446inter4, gate446inter5, gate446inter6, gate446inter7, gate446inter8, gate446inter9, gate446inter10, gate446inter11, gate446inter12, gate208inter0, gate208inter1, gate208inter2, gate208inter3, gate208inter4, gate208inter5, gate208inter6, gate208inter7, gate208inter8, gate208inter9, gate208inter10, gate208inter11, gate208inter12, gate213inter0, gate213inter1, gate213inter2, gate213inter3, gate213inter4, gate213inter5, gate213inter6, gate213inter7, gate213inter8, gate213inter9, gate213inter10, gate213inter11, gate213inter12, gate445inter0, gate445inter1, gate445inter2, gate445inter3, gate445inter4, gate445inter5, gate445inter6, gate445inter7, gate445inter8, gate445inter9, gate445inter10, gate445inter11, gate445inter12, gate491inter0, gate491inter1, gate491inter2, gate491inter3, gate491inter4, gate491inter5, gate491inter6, gate491inter7, gate491inter8, gate491inter9, gate491inter10, gate491inter11, gate491inter12, gate239inter0, gate239inter1, gate239inter2, gate239inter3, gate239inter4, gate239inter5, gate239inter6, gate239inter7, gate239inter8, gate239inter9, gate239inter10, gate239inter11, gate239inter12, gate417inter0, gate417inter1, gate417inter2, gate417inter3, gate417inter4, gate417inter5, gate417inter6, gate417inter7, gate417inter8, gate417inter9, gate417inter10, gate417inter11, gate417inter12, gate31inter0, gate31inter1, gate31inter2, gate31inter3, gate31inter4, gate31inter5, gate31inter6, gate31inter7, gate31inter8, gate31inter9, gate31inter10, gate31inter11, gate31inter12, gate281inter0, gate281inter1, gate281inter2, gate281inter3, gate281inter4, gate281inter5, gate281inter6, gate281inter7, gate281inter8, gate281inter9, gate281inter10, gate281inter11, gate281inter12, gate130inter0, gate130inter1, gate130inter2, gate130inter3, gate130inter4, gate130inter5, gate130inter6, gate130inter7, gate130inter8, gate130inter9, gate130inter10, gate130inter11, gate130inter12, gate155inter0, gate155inter1, gate155inter2, gate155inter3, gate155inter4, gate155inter5, gate155inter6, gate155inter7, gate155inter8, gate155inter9, gate155inter10, gate155inter11, gate155inter12, gate395inter0, gate395inter1, gate395inter2, gate395inter3, gate395inter4, gate395inter5, gate395inter6, gate395inter7, gate395inter8, gate395inter9, gate395inter10, gate395inter11, gate395inter12, gate106inter0, gate106inter1, gate106inter2, gate106inter3, gate106inter4, gate106inter5, gate106inter6, gate106inter7, gate106inter8, gate106inter9, gate106inter10, gate106inter11, gate106inter12, gate233inter0, gate233inter1, gate233inter2, gate233inter3, gate233inter4, gate233inter5, gate233inter6, gate233inter7, gate233inter8, gate233inter9, gate233inter10, gate233inter11, gate233inter12, gate512inter0, gate512inter1, gate512inter2, gate512inter3, gate512inter4, gate512inter5, gate512inter6, gate512inter7, gate512inter8, gate512inter9, gate512inter10, gate512inter11, gate512inter12, gate461inter0, gate461inter1, gate461inter2, gate461inter3, gate461inter4, gate461inter5, gate461inter6, gate461inter7, gate461inter8, gate461inter9, gate461inter10, gate461inter11, gate461inter12, gate63inter0, gate63inter1, gate63inter2, gate63inter3, gate63inter4, gate63inter5, gate63inter6, gate63inter7, gate63inter8, gate63inter9, gate63inter10, gate63inter11, gate63inter12, gate36inter0, gate36inter1, gate36inter2, gate36inter3, gate36inter4, gate36inter5, gate36inter6, gate36inter7, gate36inter8, gate36inter9, gate36inter10, gate36inter11, gate36inter12, gate503inter0, gate503inter1, gate503inter2, gate503inter3, gate503inter4, gate503inter5, gate503inter6, gate503inter7, gate503inter8, gate503inter9, gate503inter10, gate503inter11, gate503inter12, gate457inter0, gate457inter1, gate457inter2, gate457inter3, gate457inter4, gate457inter5, gate457inter6, gate457inter7, gate457inter8, gate457inter9, gate457inter10, gate457inter11, gate457inter12, gate37inter0, gate37inter1, gate37inter2, gate37inter3, gate37inter4, gate37inter5, gate37inter6, gate37inter7, gate37inter8, gate37inter9, gate37inter10, gate37inter11, gate37inter12, gate25inter0, gate25inter1, gate25inter2, gate25inter3, gate25inter4, gate25inter5, gate25inter6, gate25inter7, gate25inter8, gate25inter9, gate25inter10, gate25inter11, gate25inter12, gate74inter0, gate74inter1, gate74inter2, gate74inter3, gate74inter4, gate74inter5, gate74inter6, gate74inter7, gate74inter8, gate74inter9, gate74inter10, gate74inter11, gate74inter12, gate200inter0, gate200inter1, gate200inter2, gate200inter3, gate200inter4, gate200inter5, gate200inter6, gate200inter7, gate200inter8, gate200inter9, gate200inter10, gate200inter11, gate200inter12, gate131inter0, gate131inter1, gate131inter2, gate131inter3, gate131inter4, gate131inter5, gate131inter6, gate131inter7, gate131inter8, gate131inter9, gate131inter10, gate131inter11, gate131inter12, gate272inter0, gate272inter1, gate272inter2, gate272inter3, gate272inter4, gate272inter5, gate272inter6, gate272inter7, gate272inter8, gate272inter9, gate272inter10, gate272inter11, gate272inter12, gate289inter0, gate289inter1, gate289inter2, gate289inter3, gate289inter4, gate289inter5, gate289inter6, gate289inter7, gate289inter8, gate289inter9, gate289inter10, gate289inter11, gate289inter12, gate455inter0, gate455inter1, gate455inter2, gate455inter3, gate455inter4, gate455inter5, gate455inter6, gate455inter7, gate455inter8, gate455inter9, gate455inter10, gate455inter11, gate455inter12, gate115inter0, gate115inter1, gate115inter2, gate115inter3, gate115inter4, gate115inter5, gate115inter6, gate115inter7, gate115inter8, gate115inter9, gate115inter10, gate115inter11, gate115inter12, gate228inter0, gate228inter1, gate228inter2, gate228inter3, gate228inter4, gate228inter5, gate228inter6, gate228inter7, gate228inter8, gate228inter9, gate228inter10, gate228inter11, gate228inter12, gate222inter0, gate222inter1, gate222inter2, gate222inter3, gate222inter4, gate222inter5, gate222inter6, gate222inter7, gate222inter8, gate222inter9, gate222inter10, gate222inter11, gate222inter12, gate401inter0, gate401inter1, gate401inter2, gate401inter3, gate401inter4, gate401inter5, gate401inter6, gate401inter7, gate401inter8, gate401inter9, gate401inter10, gate401inter11, gate401inter12, gate264inter0, gate264inter1, gate264inter2, gate264inter3, gate264inter4, gate264inter5, gate264inter6, gate264inter7, gate264inter8, gate264inter9, gate264inter10, gate264inter11, gate264inter12, gate99inter0, gate99inter1, gate99inter2, gate99inter3, gate99inter4, gate99inter5, gate99inter6, gate99inter7, gate99inter8, gate99inter9, gate99inter10, gate99inter11, gate99inter12, gate507inter0, gate507inter1, gate507inter2, gate507inter3, gate507inter4, gate507inter5, gate507inter6, gate507inter7, gate507inter8, gate507inter9, gate507inter10, gate507inter11, gate507inter12, gate181inter0, gate181inter1, gate181inter2, gate181inter3, gate181inter4, gate181inter5, gate181inter6, gate181inter7, gate181inter8, gate181inter9, gate181inter10, gate181inter11, gate181inter12, gate126inter0, gate126inter1, gate126inter2, gate126inter3, gate126inter4, gate126inter5, gate126inter6, gate126inter7, gate126inter8, gate126inter9, gate126inter10, gate126inter11, gate126inter12, gate467inter0, gate467inter1, gate467inter2, gate467inter3, gate467inter4, gate467inter5, gate467inter6, gate467inter7, gate467inter8, gate467inter9, gate467inter10, gate467inter11, gate467inter12, gate218inter0, gate218inter1, gate218inter2, gate218inter3, gate218inter4, gate218inter5, gate218inter6, gate218inter7, gate218inter8, gate218inter9, gate218inter10, gate218inter11, gate218inter12, gate471inter0, gate471inter1, gate471inter2, gate471inter3, gate471inter4, gate471inter5, gate471inter6, gate471inter7, gate471inter8, gate471inter9, gate471inter10, gate471inter11, gate471inter12, gate144inter0, gate144inter1, gate144inter2, gate144inter3, gate144inter4, gate144inter5, gate144inter6, gate144inter7, gate144inter8, gate144inter9, gate144inter10, gate144inter11, gate144inter12, gate276inter0, gate276inter1, gate276inter2, gate276inter3, gate276inter4, gate276inter5, gate276inter6, gate276inter7, gate276inter8, gate276inter9, gate276inter10, gate276inter11, gate276inter12, gate398inter0, gate398inter1, gate398inter2, gate398inter3, gate398inter4, gate398inter5, gate398inter6, gate398inter7, gate398inter8, gate398inter9, gate398inter10, gate398inter11, gate398inter12, gate101inter0, gate101inter1, gate101inter2, gate101inter3, gate101inter4, gate101inter5, gate101inter6, gate101inter7, gate101inter8, gate101inter9, gate101inter10, gate101inter11, gate101inter12, gate260inter0, gate260inter1, gate260inter2, gate260inter3, gate260inter4, gate260inter5, gate260inter6, gate260inter7, gate260inter8, gate260inter9, gate260inter10, gate260inter11, gate260inter12, gate188inter0, gate188inter1, gate188inter2, gate188inter3, gate188inter4, gate188inter5, gate188inter6, gate188inter7, gate188inter8, gate188inter9, gate188inter10, gate188inter11, gate188inter12, gate52inter0, gate52inter1, gate52inter2, gate52inter3, gate52inter4, gate52inter5, gate52inter6, gate52inter7, gate52inter8, gate52inter9, gate52inter10, gate52inter11, gate52inter12, gate215inter0, gate215inter1, gate215inter2, gate215inter3, gate215inter4, gate215inter5, gate215inter6, gate215inter7, gate215inter8, gate215inter9, gate215inter10, gate215inter11, gate215inter12, gate49inter0, gate49inter1, gate49inter2, gate49inter3, gate49inter4, gate49inter5, gate49inter6, gate49inter7, gate49inter8, gate49inter9, gate49inter10, gate49inter11, gate49inter12, gate55inter0, gate55inter1, gate55inter2, gate55inter3, gate55inter4, gate55inter5, gate55inter6, gate55inter7, gate55inter8, gate55inter9, gate55inter10, gate55inter11, gate55inter12, gate44inter0, gate44inter1, gate44inter2, gate44inter3, gate44inter4, gate44inter5, gate44inter6, gate44inter7, gate44inter8, gate44inter9, gate44inter10, gate44inter11, gate44inter12, gate393inter0, gate393inter1, gate393inter2, gate393inter3, gate393inter4, gate393inter5, gate393inter6, gate393inter7, gate393inter8, gate393inter9, gate393inter10, gate393inter11, gate393inter12, gate496inter0, gate496inter1, gate496inter2, gate496inter3, gate496inter4, gate496inter5, gate496inter6, gate496inter7, gate496inter8, gate496inter9, gate496inter10, gate496inter11, gate496inter12, gate511inter0, gate511inter1, gate511inter2, gate511inter3, gate511inter4, gate511inter5, gate511inter6, gate511inter7, gate511inter8, gate511inter9, gate511inter10, gate511inter11, gate511inter12, gate87inter0, gate87inter1, gate87inter2, gate87inter3, gate87inter4, gate87inter5, gate87inter6, gate87inter7, gate87inter8, gate87inter9, gate87inter10, gate87inter11, gate87inter12, gate170inter0, gate170inter1, gate170inter2, gate170inter3, gate170inter4, gate170inter5, gate170inter6, gate170inter7, gate170inter8, gate170inter9, gate170inter10, gate170inter11, gate170inter12, gate46inter0, gate46inter1, gate46inter2, gate46inter3, gate46inter4, gate46inter5, gate46inter6, gate46inter7, gate46inter8, gate46inter9, gate46inter10, gate46inter11, gate46inter12, gate190inter0, gate190inter1, gate190inter2, gate190inter3, gate190inter4, gate190inter5, gate190inter6, gate190inter7, gate190inter8, gate190inter9, gate190inter10, gate190inter11, gate190inter12, gate428inter0, gate428inter1, gate428inter2, gate428inter3, gate428inter4, gate428inter5, gate428inter6, gate428inter7, gate428inter8, gate428inter9, gate428inter10, gate428inter11, gate428inter12, gate174inter0, gate174inter1, gate174inter2, gate174inter3, gate174inter4, gate174inter5, gate174inter6, gate174inter7, gate174inter8, gate174inter9, gate174inter10, gate174inter11, gate174inter12, gate431inter0, gate431inter1, gate431inter2, gate431inter3, gate431inter4, gate431inter5, gate431inter6, gate431inter7, gate431inter8, gate431inter9, gate431inter10, gate431inter11, gate431inter12, gate410inter0, gate410inter1, gate410inter2, gate410inter3, gate410inter4, gate410inter5, gate410inter6, gate410inter7, gate410inter8, gate410inter9, gate410inter10, gate410inter11, gate410inter12, gate473inter0, gate473inter1, gate473inter2, gate473inter3, gate473inter4, gate473inter5, gate473inter6, gate473inter7, gate473inter8, gate473inter9, gate473inter10, gate473inter11, gate473inter12, gate165inter0, gate165inter1, gate165inter2, gate165inter3, gate165inter4, gate165inter5, gate165inter6, gate165inter7, gate165inter8, gate165inter9, gate165inter10, gate165inter11, gate165inter12, gate259inter0, gate259inter1, gate259inter2, gate259inter3, gate259inter4, gate259inter5, gate259inter6, gate259inter7, gate259inter8, gate259inter9, gate259inter10, gate259inter11, gate259inter12, gate146inter0, gate146inter1, gate146inter2, gate146inter3, gate146inter4, gate146inter5, gate146inter6, gate146inter7, gate146inter8, gate146inter9, gate146inter10, gate146inter11, gate146inter12, gate237inter0, gate237inter1, gate237inter2, gate237inter3, gate237inter4, gate237inter5, gate237inter6, gate237inter7, gate237inter8, gate237inter9, gate237inter10, gate237inter11, gate237inter12, gate394inter0, gate394inter1, gate394inter2, gate394inter3, gate394inter4, gate394inter5, gate394inter6, gate394inter7, gate394inter8, gate394inter9, gate394inter10, gate394inter11, gate394inter12, gate242inter0, gate242inter1, gate242inter2, gate242inter3, gate242inter4, gate242inter5, gate242inter6, gate242inter7, gate242inter8, gate242inter9, gate242inter10, gate242inter11, gate242inter12, gate293inter0, gate293inter1, gate293inter2, gate293inter3, gate293inter4, gate293inter5, gate293inter6, gate293inter7, gate293inter8, gate293inter9, gate293inter10, gate293inter11, gate293inter12, gate86inter0, gate86inter1, gate86inter2, gate86inter3, gate86inter4, gate86inter5, gate86inter6, gate86inter7, gate86inter8, gate86inter9, gate86inter10, gate86inter11, gate86inter12, gate292inter0, gate292inter1, gate292inter2, gate292inter3, gate292inter4, gate292inter5, gate292inter6, gate292inter7, gate292inter8, gate292inter9, gate292inter10, gate292inter11, gate292inter12, gate487inter0, gate487inter1, gate487inter2, gate487inter3, gate487inter4, gate487inter5, gate487inter6, gate487inter7, gate487inter8, gate487inter9, gate487inter10, gate487inter11, gate487inter12, gate194inter0, gate194inter1, gate194inter2, gate194inter3, gate194inter4, gate194inter5, gate194inter6, gate194inter7, gate194inter8, gate194inter9, gate194inter10, gate194inter11, gate194inter12, gate478inter0, gate478inter1, gate478inter2, gate478inter3, gate478inter4, gate478inter5, gate478inter6, gate478inter7, gate478inter8, gate478inter9, gate478inter10, gate478inter11, gate478inter12, gate274inter0, gate274inter1, gate274inter2, gate274inter3, gate274inter4, gate274inter5, gate274inter6, gate274inter7, gate274inter8, gate274inter9, gate274inter10, gate274inter11, gate274inter12, gate397inter0, gate397inter1, gate397inter2, gate397inter3, gate397inter4, gate397inter5, gate397inter6, gate397inter7, gate397inter8, gate397inter9, gate397inter10, gate397inter11, gate397inter12, gate266inter0, gate266inter1, gate266inter2, gate266inter3, gate266inter4, gate266inter5, gate266inter6, gate266inter7, gate266inter8, gate266inter9, gate266inter10, gate266inter11, gate266inter12, gate157inter0, gate157inter1, gate157inter2, gate157inter3, gate157inter4, gate157inter5, gate157inter6, gate157inter7, gate157inter8, gate157inter9, gate157inter10, gate157inter11, gate157inter12, gate296inter0, gate296inter1, gate296inter2, gate296inter3, gate296inter4, gate296inter5, gate296inter6, gate296inter7, gate296inter8, gate296inter9, gate296inter10, gate296inter11, gate296inter12, gate145inter0, gate145inter1, gate145inter2, gate145inter3, gate145inter4, gate145inter5, gate145inter6, gate145inter7, gate145inter8, gate145inter9, gate145inter10, gate145inter11, gate145inter12, gate429inter0, gate429inter1, gate429inter2, gate429inter3, gate429inter4, gate429inter5, gate429inter6, gate429inter7, gate429inter8, gate429inter9, gate429inter10, gate429inter11, gate429inter12, gate220inter0, gate220inter1, gate220inter2, gate220inter3, gate220inter4, gate220inter5, gate220inter6, gate220inter7, gate220inter8, gate220inter9, gate220inter10, gate220inter11, gate220inter12, gate13inter0, gate13inter1, gate13inter2, gate13inter3, gate13inter4, gate13inter5, gate13inter6, gate13inter7, gate13inter8, gate13inter9, gate13inter10, gate13inter11, gate13inter12, gate399inter0, gate399inter1, gate399inter2, gate399inter3, gate399inter4, gate399inter5, gate399inter6, gate399inter7, gate399inter8, gate399inter9, gate399inter10, gate399inter11, gate399inter12, gate514inter0, gate514inter1, gate514inter2, gate514inter3, gate514inter4, gate514inter5, gate514inter6, gate514inter7, gate514inter8, gate514inter9, gate514inter10, gate514inter11, gate514inter12, gate127inter0, gate127inter1, gate127inter2, gate127inter3, gate127inter4, gate127inter5, gate127inter6, gate127inter7, gate127inter8, gate127inter9, gate127inter10, gate127inter11, gate127inter12, gate451inter0, gate451inter1, gate451inter2, gate451inter3, gate451inter4, gate451inter5, gate451inter6, gate451inter7, gate451inter8, gate451inter9, gate451inter10, gate451inter11, gate451inter12, gate472inter0, gate472inter1, gate472inter2, gate472inter3, gate472inter4, gate472inter5, gate472inter6, gate472inter7, gate472inter8, gate472inter9, gate472inter10, gate472inter11, gate472inter12, gate122inter0, gate122inter1, gate122inter2, gate122inter3, gate122inter4, gate122inter5, gate122inter6, gate122inter7, gate122inter8, gate122inter9, gate122inter10, gate122inter11, gate122inter12, gate191inter0, gate191inter1, gate191inter2, gate191inter3, gate191inter4, gate191inter5, gate191inter6, gate191inter7, gate191inter8, gate191inter9, gate191inter10, gate191inter11, gate191inter12, gate192inter0, gate192inter1, gate192inter2, gate192inter3, gate192inter4, gate192inter5, gate192inter6, gate192inter7, gate192inter8, gate192inter9, gate192inter10, gate192inter11, gate192inter12, gate162inter0, gate162inter1, gate162inter2, gate162inter3, gate162inter4, gate162inter5, gate162inter6, gate162inter7, gate162inter8, gate162inter9, gate162inter10, gate162inter11, gate162inter12, gate493inter0, gate493inter1, gate493inter2, gate493inter3, gate493inter4, gate493inter5, gate493inter6, gate493inter7, gate493inter8, gate493inter9, gate493inter10, gate493inter11, gate493inter12, gate79inter0, gate79inter1, gate79inter2, gate79inter3, gate79inter4, gate79inter5, gate79inter6, gate79inter7, gate79inter8, gate79inter9, gate79inter10, gate79inter11, gate79inter12, gate47inter0, gate47inter1, gate47inter2, gate47inter3, gate47inter4, gate47inter5, gate47inter6, gate47inter7, gate47inter8, gate47inter9, gate47inter10, gate47inter11, gate47inter12, gate23inter0, gate23inter1, gate23inter2, gate23inter3, gate23inter4, gate23inter5, gate23inter6, gate23inter7, gate23inter8, gate23inter9, gate23inter10, gate23inter11, gate23inter12, gate201inter0, gate201inter1, gate201inter2, gate201inter3, gate201inter4, gate201inter5, gate201inter6, gate201inter7, gate201inter8, gate201inter9, gate201inter10, gate201inter11, gate201inter12, gate470inter0, gate470inter1, gate470inter2, gate470inter3, gate470inter4, gate470inter5, gate470inter6, gate470inter7, gate470inter8, gate470inter9, gate470inter10, gate470inter11, gate470inter12, gate254inter0, gate254inter1, gate254inter2, gate254inter3, gate254inter4, gate254inter5, gate254inter6, gate254inter7, gate254inter8, gate254inter9, gate254inter10, gate254inter11, gate254inter12, gate415inter0, gate415inter1, gate415inter2, gate415inter3, gate415inter4, gate415inter5, gate415inter6, gate415inter7, gate415inter8, gate415inter9, gate415inter10, gate415inter11, gate415inter12, gate169inter0, gate169inter1, gate169inter2, gate169inter3, gate169inter4, gate169inter5, gate169inter6, gate169inter7, gate169inter8, gate169inter9, gate169inter10, gate169inter11, gate169inter12, gate43inter0, gate43inter1, gate43inter2, gate43inter3, gate43inter4, gate43inter5, gate43inter6, gate43inter7, gate43inter8, gate43inter9, gate43inter10, gate43inter11, gate43inter12, gate406inter0, gate406inter1, gate406inter2, gate406inter3, gate406inter4, gate406inter5, gate406inter6, gate406inter7, gate406inter8, gate406inter9, gate406inter10, gate406inter11, gate406inter12, gate50inter0, gate50inter1, gate50inter2, gate50inter3, gate50inter4, gate50inter5, gate50inter6, gate50inter7, gate50inter8, gate50inter9, gate50inter10, gate50inter11, gate50inter12, gate66inter0, gate66inter1, gate66inter2, gate66inter3, gate66inter4, gate66inter5, gate66inter6, gate66inter7, gate66inter8, gate66inter9, gate66inter10, gate66inter11, gate66inter12, gate76inter0, gate76inter1, gate76inter2, gate76inter3, gate76inter4, gate76inter5, gate76inter6, gate76inter7, gate76inter8, gate76inter9, gate76inter10, gate76inter11, gate76inter12, gate212inter0, gate212inter1, gate212inter2, gate212inter3, gate212inter4, gate212inter5, gate212inter6, gate212inter7, gate212inter8, gate212inter9, gate212inter10, gate212inter11, gate212inter12;



and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );
nand2 gate9( .a(G1), .b(G2), .O(G266) );
nand2 gate10( .a(G3), .b(G4), .O(G269) );
nand2 gate11( .a(G5), .b(G6), .O(G272) );
nand2 gate12( .a(G7), .b(G8), .O(G275) );

  xor2  gate2031(.a(G10), .b(G9), .O(gate13inter0));
  nand2 gate2032(.a(gate13inter0), .b(s_212), .O(gate13inter1));
  and2  gate2033(.a(G10), .b(G9), .O(gate13inter2));
  inv1  gate2034(.a(s_212), .O(gate13inter3));
  inv1  gate2035(.a(s_213), .O(gate13inter4));
  nand2 gate2036(.a(gate13inter4), .b(gate13inter3), .O(gate13inter5));
  nor2  gate2037(.a(gate13inter5), .b(gate13inter2), .O(gate13inter6));
  inv1  gate2038(.a(G9), .O(gate13inter7));
  inv1  gate2039(.a(G10), .O(gate13inter8));
  nand2 gate2040(.a(gate13inter8), .b(gate13inter7), .O(gate13inter9));
  nand2 gate2041(.a(s_213), .b(gate13inter3), .O(gate13inter10));
  nor2  gate2042(.a(gate13inter10), .b(gate13inter9), .O(gate13inter11));
  nor2  gate2043(.a(gate13inter11), .b(gate13inter6), .O(gate13inter12));
  nand2 gate2044(.a(gate13inter12), .b(gate13inter1), .O(G278));
nand2 gate14( .a(G11), .b(G12), .O(G281) );
nand2 gate15( .a(G13), .b(G14), .O(G284) );
nand2 gate16( .a(G15), .b(G16), .O(G287) );
nand2 gate17( .a(G17), .b(G18), .O(G290) );

  xor2  gate617(.a(G20), .b(G19), .O(gate18inter0));
  nand2 gate618(.a(gate18inter0), .b(s_10), .O(gate18inter1));
  and2  gate619(.a(G20), .b(G19), .O(gate18inter2));
  inv1  gate620(.a(s_10), .O(gate18inter3));
  inv1  gate621(.a(s_11), .O(gate18inter4));
  nand2 gate622(.a(gate18inter4), .b(gate18inter3), .O(gate18inter5));
  nor2  gate623(.a(gate18inter5), .b(gate18inter2), .O(gate18inter6));
  inv1  gate624(.a(G19), .O(gate18inter7));
  inv1  gate625(.a(G20), .O(gate18inter8));
  nand2 gate626(.a(gate18inter8), .b(gate18inter7), .O(gate18inter9));
  nand2 gate627(.a(s_11), .b(gate18inter3), .O(gate18inter10));
  nor2  gate628(.a(gate18inter10), .b(gate18inter9), .O(gate18inter11));
  nor2  gate629(.a(gate18inter11), .b(gate18inter6), .O(gate18inter12));
  nand2 gate630(.a(gate18inter12), .b(gate18inter1), .O(G293));
nand2 gate19( .a(G21), .b(G22), .O(G296) );
nand2 gate20( .a(G23), .b(G24), .O(G299) );
nand2 gate21( .a(G25), .b(G26), .O(G302) );
nand2 gate22( .a(G27), .b(G28), .O(G305) );

  xor2  gate2213(.a(G30), .b(G29), .O(gate23inter0));
  nand2 gate2214(.a(gate23inter0), .b(s_238), .O(gate23inter1));
  and2  gate2215(.a(G30), .b(G29), .O(gate23inter2));
  inv1  gate2216(.a(s_238), .O(gate23inter3));
  inv1  gate2217(.a(s_239), .O(gate23inter4));
  nand2 gate2218(.a(gate23inter4), .b(gate23inter3), .O(gate23inter5));
  nor2  gate2219(.a(gate23inter5), .b(gate23inter2), .O(gate23inter6));
  inv1  gate2220(.a(G29), .O(gate23inter7));
  inv1  gate2221(.a(G30), .O(gate23inter8));
  nand2 gate2222(.a(gate23inter8), .b(gate23inter7), .O(gate23inter9));
  nand2 gate2223(.a(s_239), .b(gate23inter3), .O(gate23inter10));
  nor2  gate2224(.a(gate23inter10), .b(gate23inter9), .O(gate23inter11));
  nor2  gate2225(.a(gate23inter11), .b(gate23inter6), .O(gate23inter12));
  nand2 gate2226(.a(gate23inter12), .b(gate23inter1), .O(G308));
nand2 gate24( .a(G31), .b(G32), .O(G311) );

  xor2  gate1163(.a(G5), .b(G1), .O(gate25inter0));
  nand2 gate1164(.a(gate25inter0), .b(s_88), .O(gate25inter1));
  and2  gate1165(.a(G5), .b(G1), .O(gate25inter2));
  inv1  gate1166(.a(s_88), .O(gate25inter3));
  inv1  gate1167(.a(s_89), .O(gate25inter4));
  nand2 gate1168(.a(gate25inter4), .b(gate25inter3), .O(gate25inter5));
  nor2  gate1169(.a(gate25inter5), .b(gate25inter2), .O(gate25inter6));
  inv1  gate1170(.a(G1), .O(gate25inter7));
  inv1  gate1171(.a(G5), .O(gate25inter8));
  nand2 gate1172(.a(gate25inter8), .b(gate25inter7), .O(gate25inter9));
  nand2 gate1173(.a(s_89), .b(gate25inter3), .O(gate25inter10));
  nor2  gate1174(.a(gate25inter10), .b(gate25inter9), .O(gate25inter11));
  nor2  gate1175(.a(gate25inter11), .b(gate25inter6), .O(gate25inter12));
  nand2 gate1176(.a(gate25inter12), .b(gate25inter1), .O(G314));
nand2 gate26( .a(G9), .b(G13), .O(G317) );
nand2 gate27( .a(G2), .b(G6), .O(G320) );
nand2 gate28( .a(G10), .b(G14), .O(G323) );
nand2 gate29( .a(G3), .b(G7), .O(G326) );
nand2 gate30( .a(G11), .b(G15), .O(G329) );

  xor2  gate967(.a(G8), .b(G4), .O(gate31inter0));
  nand2 gate968(.a(gate31inter0), .b(s_60), .O(gate31inter1));
  and2  gate969(.a(G8), .b(G4), .O(gate31inter2));
  inv1  gate970(.a(s_60), .O(gate31inter3));
  inv1  gate971(.a(s_61), .O(gate31inter4));
  nand2 gate972(.a(gate31inter4), .b(gate31inter3), .O(gate31inter5));
  nor2  gate973(.a(gate31inter5), .b(gate31inter2), .O(gate31inter6));
  inv1  gate974(.a(G4), .O(gate31inter7));
  inv1  gate975(.a(G8), .O(gate31inter8));
  nand2 gate976(.a(gate31inter8), .b(gate31inter7), .O(gate31inter9));
  nand2 gate977(.a(s_61), .b(gate31inter3), .O(gate31inter10));
  nor2  gate978(.a(gate31inter10), .b(gate31inter9), .O(gate31inter11));
  nor2  gate979(.a(gate31inter11), .b(gate31inter6), .O(gate31inter12));
  nand2 gate980(.a(gate31inter12), .b(gate31inter1), .O(G332));
nand2 gate32( .a(G12), .b(G16), .O(G335) );
nand2 gate33( .a(G17), .b(G21), .O(G338) );
nand2 gate34( .a(G25), .b(G29), .O(G341) );
nand2 gate35( .a(G18), .b(G22), .O(G344) );

  xor2  gate1107(.a(G30), .b(G26), .O(gate36inter0));
  nand2 gate1108(.a(gate36inter0), .b(s_80), .O(gate36inter1));
  and2  gate1109(.a(G30), .b(G26), .O(gate36inter2));
  inv1  gate1110(.a(s_80), .O(gate36inter3));
  inv1  gate1111(.a(s_81), .O(gate36inter4));
  nand2 gate1112(.a(gate36inter4), .b(gate36inter3), .O(gate36inter5));
  nor2  gate1113(.a(gate36inter5), .b(gate36inter2), .O(gate36inter6));
  inv1  gate1114(.a(G26), .O(gate36inter7));
  inv1  gate1115(.a(G30), .O(gate36inter8));
  nand2 gate1116(.a(gate36inter8), .b(gate36inter7), .O(gate36inter9));
  nand2 gate1117(.a(s_81), .b(gate36inter3), .O(gate36inter10));
  nor2  gate1118(.a(gate36inter10), .b(gate36inter9), .O(gate36inter11));
  nor2  gate1119(.a(gate36inter11), .b(gate36inter6), .O(gate36inter12));
  nand2 gate1120(.a(gate36inter12), .b(gate36inter1), .O(G347));

  xor2  gate1149(.a(G23), .b(G19), .O(gate37inter0));
  nand2 gate1150(.a(gate37inter0), .b(s_86), .O(gate37inter1));
  and2  gate1151(.a(G23), .b(G19), .O(gate37inter2));
  inv1  gate1152(.a(s_86), .O(gate37inter3));
  inv1  gate1153(.a(s_87), .O(gate37inter4));
  nand2 gate1154(.a(gate37inter4), .b(gate37inter3), .O(gate37inter5));
  nor2  gate1155(.a(gate37inter5), .b(gate37inter2), .O(gate37inter6));
  inv1  gate1156(.a(G19), .O(gate37inter7));
  inv1  gate1157(.a(G23), .O(gate37inter8));
  nand2 gate1158(.a(gate37inter8), .b(gate37inter7), .O(gate37inter9));
  nand2 gate1159(.a(s_87), .b(gate37inter3), .O(gate37inter10));
  nor2  gate1160(.a(gate37inter10), .b(gate37inter9), .O(gate37inter11));
  nor2  gate1161(.a(gate37inter11), .b(gate37inter6), .O(gate37inter12));
  nand2 gate1162(.a(gate37inter12), .b(gate37inter1), .O(G350));
nand2 gate38( .a(G27), .b(G31), .O(G353) );
nand2 gate39( .a(G20), .b(G24), .O(G356) );
nand2 gate40( .a(G28), .b(G32), .O(G359) );

  xor2  gate785(.a(G266), .b(G1), .O(gate41inter0));
  nand2 gate786(.a(gate41inter0), .b(s_34), .O(gate41inter1));
  and2  gate787(.a(G266), .b(G1), .O(gate41inter2));
  inv1  gate788(.a(s_34), .O(gate41inter3));
  inv1  gate789(.a(s_35), .O(gate41inter4));
  nand2 gate790(.a(gate41inter4), .b(gate41inter3), .O(gate41inter5));
  nor2  gate791(.a(gate41inter5), .b(gate41inter2), .O(gate41inter6));
  inv1  gate792(.a(G1), .O(gate41inter7));
  inv1  gate793(.a(G266), .O(gate41inter8));
  nand2 gate794(.a(gate41inter8), .b(gate41inter7), .O(gate41inter9));
  nand2 gate795(.a(s_35), .b(gate41inter3), .O(gate41inter10));
  nor2  gate796(.a(gate41inter10), .b(gate41inter9), .O(gate41inter11));
  nor2  gate797(.a(gate41inter11), .b(gate41inter6), .O(gate41inter12));
  nand2 gate798(.a(gate41inter12), .b(gate41inter1), .O(G362));
nand2 gate42( .a(G2), .b(G266), .O(G363) );

  xor2  gate2297(.a(G269), .b(G3), .O(gate43inter0));
  nand2 gate2298(.a(gate43inter0), .b(s_250), .O(gate43inter1));
  and2  gate2299(.a(G269), .b(G3), .O(gate43inter2));
  inv1  gate2300(.a(s_250), .O(gate43inter3));
  inv1  gate2301(.a(s_251), .O(gate43inter4));
  nand2 gate2302(.a(gate43inter4), .b(gate43inter3), .O(gate43inter5));
  nor2  gate2303(.a(gate43inter5), .b(gate43inter2), .O(gate43inter6));
  inv1  gate2304(.a(G3), .O(gate43inter7));
  inv1  gate2305(.a(G269), .O(gate43inter8));
  nand2 gate2306(.a(gate43inter8), .b(gate43inter7), .O(gate43inter9));
  nand2 gate2307(.a(s_251), .b(gate43inter3), .O(gate43inter10));
  nor2  gate2308(.a(gate43inter10), .b(gate43inter9), .O(gate43inter11));
  nor2  gate2309(.a(gate43inter11), .b(gate43inter6), .O(gate43inter12));
  nand2 gate2310(.a(gate43inter12), .b(gate43inter1), .O(G364));

  xor2  gate1569(.a(G269), .b(G4), .O(gate44inter0));
  nand2 gate1570(.a(gate44inter0), .b(s_146), .O(gate44inter1));
  and2  gate1571(.a(G269), .b(G4), .O(gate44inter2));
  inv1  gate1572(.a(s_146), .O(gate44inter3));
  inv1  gate1573(.a(s_147), .O(gate44inter4));
  nand2 gate1574(.a(gate44inter4), .b(gate44inter3), .O(gate44inter5));
  nor2  gate1575(.a(gate44inter5), .b(gate44inter2), .O(gate44inter6));
  inv1  gate1576(.a(G4), .O(gate44inter7));
  inv1  gate1577(.a(G269), .O(gate44inter8));
  nand2 gate1578(.a(gate44inter8), .b(gate44inter7), .O(gate44inter9));
  nand2 gate1579(.a(s_147), .b(gate44inter3), .O(gate44inter10));
  nor2  gate1580(.a(gate44inter10), .b(gate44inter9), .O(gate44inter11));
  nor2  gate1581(.a(gate44inter11), .b(gate44inter6), .O(gate44inter12));
  nand2 gate1582(.a(gate44inter12), .b(gate44inter1), .O(G365));

  xor2  gate645(.a(G272), .b(G5), .O(gate45inter0));
  nand2 gate646(.a(gate45inter0), .b(s_14), .O(gate45inter1));
  and2  gate647(.a(G272), .b(G5), .O(gate45inter2));
  inv1  gate648(.a(s_14), .O(gate45inter3));
  inv1  gate649(.a(s_15), .O(gate45inter4));
  nand2 gate650(.a(gate45inter4), .b(gate45inter3), .O(gate45inter5));
  nor2  gate651(.a(gate45inter5), .b(gate45inter2), .O(gate45inter6));
  inv1  gate652(.a(G5), .O(gate45inter7));
  inv1  gate653(.a(G272), .O(gate45inter8));
  nand2 gate654(.a(gate45inter8), .b(gate45inter7), .O(gate45inter9));
  nand2 gate655(.a(s_15), .b(gate45inter3), .O(gate45inter10));
  nor2  gate656(.a(gate45inter10), .b(gate45inter9), .O(gate45inter11));
  nor2  gate657(.a(gate45inter11), .b(gate45inter6), .O(gate45inter12));
  nand2 gate658(.a(gate45inter12), .b(gate45inter1), .O(G366));

  xor2  gate1653(.a(G272), .b(G6), .O(gate46inter0));
  nand2 gate1654(.a(gate46inter0), .b(s_158), .O(gate46inter1));
  and2  gate1655(.a(G272), .b(G6), .O(gate46inter2));
  inv1  gate1656(.a(s_158), .O(gate46inter3));
  inv1  gate1657(.a(s_159), .O(gate46inter4));
  nand2 gate1658(.a(gate46inter4), .b(gate46inter3), .O(gate46inter5));
  nor2  gate1659(.a(gate46inter5), .b(gate46inter2), .O(gate46inter6));
  inv1  gate1660(.a(G6), .O(gate46inter7));
  inv1  gate1661(.a(G272), .O(gate46inter8));
  nand2 gate1662(.a(gate46inter8), .b(gate46inter7), .O(gate46inter9));
  nand2 gate1663(.a(s_159), .b(gate46inter3), .O(gate46inter10));
  nor2  gate1664(.a(gate46inter10), .b(gate46inter9), .O(gate46inter11));
  nor2  gate1665(.a(gate46inter11), .b(gate46inter6), .O(gate46inter12));
  nand2 gate1666(.a(gate46inter12), .b(gate46inter1), .O(G367));

  xor2  gate2199(.a(G275), .b(G7), .O(gate47inter0));
  nand2 gate2200(.a(gate47inter0), .b(s_236), .O(gate47inter1));
  and2  gate2201(.a(G275), .b(G7), .O(gate47inter2));
  inv1  gate2202(.a(s_236), .O(gate47inter3));
  inv1  gate2203(.a(s_237), .O(gate47inter4));
  nand2 gate2204(.a(gate47inter4), .b(gate47inter3), .O(gate47inter5));
  nor2  gate2205(.a(gate47inter5), .b(gate47inter2), .O(gate47inter6));
  inv1  gate2206(.a(G7), .O(gate47inter7));
  inv1  gate2207(.a(G275), .O(gate47inter8));
  nand2 gate2208(.a(gate47inter8), .b(gate47inter7), .O(gate47inter9));
  nand2 gate2209(.a(s_237), .b(gate47inter3), .O(gate47inter10));
  nor2  gate2210(.a(gate47inter10), .b(gate47inter9), .O(gate47inter11));
  nor2  gate2211(.a(gate47inter11), .b(gate47inter6), .O(gate47inter12));
  nand2 gate2212(.a(gate47inter12), .b(gate47inter1), .O(G368));
nand2 gate48( .a(G8), .b(G275), .O(G369) );

  xor2  gate1541(.a(G278), .b(G9), .O(gate49inter0));
  nand2 gate1542(.a(gate49inter0), .b(s_142), .O(gate49inter1));
  and2  gate1543(.a(G278), .b(G9), .O(gate49inter2));
  inv1  gate1544(.a(s_142), .O(gate49inter3));
  inv1  gate1545(.a(s_143), .O(gate49inter4));
  nand2 gate1546(.a(gate49inter4), .b(gate49inter3), .O(gate49inter5));
  nor2  gate1547(.a(gate49inter5), .b(gate49inter2), .O(gate49inter6));
  inv1  gate1548(.a(G9), .O(gate49inter7));
  inv1  gate1549(.a(G278), .O(gate49inter8));
  nand2 gate1550(.a(gate49inter8), .b(gate49inter7), .O(gate49inter9));
  nand2 gate1551(.a(s_143), .b(gate49inter3), .O(gate49inter10));
  nor2  gate1552(.a(gate49inter10), .b(gate49inter9), .O(gate49inter11));
  nor2  gate1553(.a(gate49inter11), .b(gate49inter6), .O(gate49inter12));
  nand2 gate1554(.a(gate49inter12), .b(gate49inter1), .O(G370));

  xor2  gate2325(.a(G278), .b(G10), .O(gate50inter0));
  nand2 gate2326(.a(gate50inter0), .b(s_254), .O(gate50inter1));
  and2  gate2327(.a(G278), .b(G10), .O(gate50inter2));
  inv1  gate2328(.a(s_254), .O(gate50inter3));
  inv1  gate2329(.a(s_255), .O(gate50inter4));
  nand2 gate2330(.a(gate50inter4), .b(gate50inter3), .O(gate50inter5));
  nor2  gate2331(.a(gate50inter5), .b(gate50inter2), .O(gate50inter6));
  inv1  gate2332(.a(G10), .O(gate50inter7));
  inv1  gate2333(.a(G278), .O(gate50inter8));
  nand2 gate2334(.a(gate50inter8), .b(gate50inter7), .O(gate50inter9));
  nand2 gate2335(.a(s_255), .b(gate50inter3), .O(gate50inter10));
  nor2  gate2336(.a(gate50inter10), .b(gate50inter9), .O(gate50inter11));
  nor2  gate2337(.a(gate50inter11), .b(gate50inter6), .O(gate50inter12));
  nand2 gate2338(.a(gate50inter12), .b(gate50inter1), .O(G371));
nand2 gate51( .a(G11), .b(G281), .O(G372) );

  xor2  gate1513(.a(G281), .b(G12), .O(gate52inter0));
  nand2 gate1514(.a(gate52inter0), .b(s_138), .O(gate52inter1));
  and2  gate1515(.a(G281), .b(G12), .O(gate52inter2));
  inv1  gate1516(.a(s_138), .O(gate52inter3));
  inv1  gate1517(.a(s_139), .O(gate52inter4));
  nand2 gate1518(.a(gate52inter4), .b(gate52inter3), .O(gate52inter5));
  nor2  gate1519(.a(gate52inter5), .b(gate52inter2), .O(gate52inter6));
  inv1  gate1520(.a(G12), .O(gate52inter7));
  inv1  gate1521(.a(G281), .O(gate52inter8));
  nand2 gate1522(.a(gate52inter8), .b(gate52inter7), .O(gate52inter9));
  nand2 gate1523(.a(s_139), .b(gate52inter3), .O(gate52inter10));
  nor2  gate1524(.a(gate52inter10), .b(gate52inter9), .O(gate52inter11));
  nor2  gate1525(.a(gate52inter11), .b(gate52inter6), .O(gate52inter12));
  nand2 gate1526(.a(gate52inter12), .b(gate52inter1), .O(G373));
nand2 gate53( .a(G13), .b(G284), .O(G374) );
nand2 gate54( .a(G14), .b(G284), .O(G375) );

  xor2  gate1555(.a(G287), .b(G15), .O(gate55inter0));
  nand2 gate1556(.a(gate55inter0), .b(s_144), .O(gate55inter1));
  and2  gate1557(.a(G287), .b(G15), .O(gate55inter2));
  inv1  gate1558(.a(s_144), .O(gate55inter3));
  inv1  gate1559(.a(s_145), .O(gate55inter4));
  nand2 gate1560(.a(gate55inter4), .b(gate55inter3), .O(gate55inter5));
  nor2  gate1561(.a(gate55inter5), .b(gate55inter2), .O(gate55inter6));
  inv1  gate1562(.a(G15), .O(gate55inter7));
  inv1  gate1563(.a(G287), .O(gate55inter8));
  nand2 gate1564(.a(gate55inter8), .b(gate55inter7), .O(gate55inter9));
  nand2 gate1565(.a(s_145), .b(gate55inter3), .O(gate55inter10));
  nor2  gate1566(.a(gate55inter10), .b(gate55inter9), .O(gate55inter11));
  nor2  gate1567(.a(gate55inter11), .b(gate55inter6), .O(gate55inter12));
  nand2 gate1568(.a(gate55inter12), .b(gate55inter1), .O(G376));
nand2 gate56( .a(G16), .b(G287), .O(G377) );
nand2 gate57( .a(G17), .b(G290), .O(G378) );
nand2 gate58( .a(G18), .b(G290), .O(G379) );
nand2 gate59( .a(G19), .b(G293), .O(G380) );
nand2 gate60( .a(G20), .b(G293), .O(G381) );
nand2 gate61( .a(G21), .b(G296), .O(G382) );
nand2 gate62( .a(G22), .b(G296), .O(G383) );

  xor2  gate1093(.a(G299), .b(G23), .O(gate63inter0));
  nand2 gate1094(.a(gate63inter0), .b(s_78), .O(gate63inter1));
  and2  gate1095(.a(G299), .b(G23), .O(gate63inter2));
  inv1  gate1096(.a(s_78), .O(gate63inter3));
  inv1  gate1097(.a(s_79), .O(gate63inter4));
  nand2 gate1098(.a(gate63inter4), .b(gate63inter3), .O(gate63inter5));
  nor2  gate1099(.a(gate63inter5), .b(gate63inter2), .O(gate63inter6));
  inv1  gate1100(.a(G23), .O(gate63inter7));
  inv1  gate1101(.a(G299), .O(gate63inter8));
  nand2 gate1102(.a(gate63inter8), .b(gate63inter7), .O(gate63inter9));
  nand2 gate1103(.a(s_79), .b(gate63inter3), .O(gate63inter10));
  nor2  gate1104(.a(gate63inter10), .b(gate63inter9), .O(gate63inter11));
  nor2  gate1105(.a(gate63inter11), .b(gate63inter6), .O(gate63inter12));
  nand2 gate1106(.a(gate63inter12), .b(gate63inter1), .O(G384));
nand2 gate64( .a(G24), .b(G299), .O(G385) );
nand2 gate65( .a(G25), .b(G302), .O(G386) );

  xor2  gate2339(.a(G302), .b(G26), .O(gate66inter0));
  nand2 gate2340(.a(gate66inter0), .b(s_256), .O(gate66inter1));
  and2  gate2341(.a(G302), .b(G26), .O(gate66inter2));
  inv1  gate2342(.a(s_256), .O(gate66inter3));
  inv1  gate2343(.a(s_257), .O(gate66inter4));
  nand2 gate2344(.a(gate66inter4), .b(gate66inter3), .O(gate66inter5));
  nor2  gate2345(.a(gate66inter5), .b(gate66inter2), .O(gate66inter6));
  inv1  gate2346(.a(G26), .O(gate66inter7));
  inv1  gate2347(.a(G302), .O(gate66inter8));
  nand2 gate2348(.a(gate66inter8), .b(gate66inter7), .O(gate66inter9));
  nand2 gate2349(.a(s_257), .b(gate66inter3), .O(gate66inter10));
  nor2  gate2350(.a(gate66inter10), .b(gate66inter9), .O(gate66inter11));
  nor2  gate2351(.a(gate66inter11), .b(gate66inter6), .O(gate66inter12));
  nand2 gate2352(.a(gate66inter12), .b(gate66inter1), .O(G387));
nand2 gate67( .a(G27), .b(G305), .O(G388) );

  xor2  gate813(.a(G305), .b(G28), .O(gate68inter0));
  nand2 gate814(.a(gate68inter0), .b(s_38), .O(gate68inter1));
  and2  gate815(.a(G305), .b(G28), .O(gate68inter2));
  inv1  gate816(.a(s_38), .O(gate68inter3));
  inv1  gate817(.a(s_39), .O(gate68inter4));
  nand2 gate818(.a(gate68inter4), .b(gate68inter3), .O(gate68inter5));
  nor2  gate819(.a(gate68inter5), .b(gate68inter2), .O(gate68inter6));
  inv1  gate820(.a(G28), .O(gate68inter7));
  inv1  gate821(.a(G305), .O(gate68inter8));
  nand2 gate822(.a(gate68inter8), .b(gate68inter7), .O(gate68inter9));
  nand2 gate823(.a(s_39), .b(gate68inter3), .O(gate68inter10));
  nor2  gate824(.a(gate68inter10), .b(gate68inter9), .O(gate68inter11));
  nor2  gate825(.a(gate68inter11), .b(gate68inter6), .O(gate68inter12));
  nand2 gate826(.a(gate68inter12), .b(gate68inter1), .O(G389));
nand2 gate69( .a(G29), .b(G308), .O(G390) );
nand2 gate70( .a(G30), .b(G308), .O(G391) );
nand2 gate71( .a(G31), .b(G311), .O(G392) );
nand2 gate72( .a(G32), .b(G311), .O(G393) );
nand2 gate73( .a(G1), .b(G314), .O(G394) );

  xor2  gate1177(.a(G314), .b(G5), .O(gate74inter0));
  nand2 gate1178(.a(gate74inter0), .b(s_90), .O(gate74inter1));
  and2  gate1179(.a(G314), .b(G5), .O(gate74inter2));
  inv1  gate1180(.a(s_90), .O(gate74inter3));
  inv1  gate1181(.a(s_91), .O(gate74inter4));
  nand2 gate1182(.a(gate74inter4), .b(gate74inter3), .O(gate74inter5));
  nor2  gate1183(.a(gate74inter5), .b(gate74inter2), .O(gate74inter6));
  inv1  gate1184(.a(G5), .O(gate74inter7));
  inv1  gate1185(.a(G314), .O(gate74inter8));
  nand2 gate1186(.a(gate74inter8), .b(gate74inter7), .O(gate74inter9));
  nand2 gate1187(.a(s_91), .b(gate74inter3), .O(gate74inter10));
  nor2  gate1188(.a(gate74inter10), .b(gate74inter9), .O(gate74inter11));
  nor2  gate1189(.a(gate74inter11), .b(gate74inter6), .O(gate74inter12));
  nand2 gate1190(.a(gate74inter12), .b(gate74inter1), .O(G395));
nand2 gate75( .a(G9), .b(G317), .O(G396) );

  xor2  gate2353(.a(G317), .b(G13), .O(gate76inter0));
  nand2 gate2354(.a(gate76inter0), .b(s_258), .O(gate76inter1));
  and2  gate2355(.a(G317), .b(G13), .O(gate76inter2));
  inv1  gate2356(.a(s_258), .O(gate76inter3));
  inv1  gate2357(.a(s_259), .O(gate76inter4));
  nand2 gate2358(.a(gate76inter4), .b(gate76inter3), .O(gate76inter5));
  nor2  gate2359(.a(gate76inter5), .b(gate76inter2), .O(gate76inter6));
  inv1  gate2360(.a(G13), .O(gate76inter7));
  inv1  gate2361(.a(G317), .O(gate76inter8));
  nand2 gate2362(.a(gate76inter8), .b(gate76inter7), .O(gate76inter9));
  nand2 gate2363(.a(s_259), .b(gate76inter3), .O(gate76inter10));
  nor2  gate2364(.a(gate76inter10), .b(gate76inter9), .O(gate76inter11));
  nor2  gate2365(.a(gate76inter11), .b(gate76inter6), .O(gate76inter12));
  nand2 gate2366(.a(gate76inter12), .b(gate76inter1), .O(G397));
nand2 gate77( .a(G2), .b(G320), .O(G398) );
nand2 gate78( .a(G6), .b(G320), .O(G399) );

  xor2  gate2185(.a(G323), .b(G10), .O(gate79inter0));
  nand2 gate2186(.a(gate79inter0), .b(s_234), .O(gate79inter1));
  and2  gate2187(.a(G323), .b(G10), .O(gate79inter2));
  inv1  gate2188(.a(s_234), .O(gate79inter3));
  inv1  gate2189(.a(s_235), .O(gate79inter4));
  nand2 gate2190(.a(gate79inter4), .b(gate79inter3), .O(gate79inter5));
  nor2  gate2191(.a(gate79inter5), .b(gate79inter2), .O(gate79inter6));
  inv1  gate2192(.a(G10), .O(gate79inter7));
  inv1  gate2193(.a(G323), .O(gate79inter8));
  nand2 gate2194(.a(gate79inter8), .b(gate79inter7), .O(gate79inter9));
  nand2 gate2195(.a(s_235), .b(gate79inter3), .O(gate79inter10));
  nor2  gate2196(.a(gate79inter10), .b(gate79inter9), .O(gate79inter11));
  nor2  gate2197(.a(gate79inter11), .b(gate79inter6), .O(gate79inter12));
  nand2 gate2198(.a(gate79inter12), .b(gate79inter1), .O(G400));
nand2 gate80( .a(G14), .b(G323), .O(G401) );
nand2 gate81( .a(G3), .b(G326), .O(G402) );
nand2 gate82( .a(G7), .b(G326), .O(G403) );
nand2 gate83( .a(G11), .b(G329), .O(G404) );
nand2 gate84( .a(G15), .b(G329), .O(G405) );
nand2 gate85( .a(G4), .b(G332), .O(G406) );

  xor2  gate1849(.a(G332), .b(G8), .O(gate86inter0));
  nand2 gate1850(.a(gate86inter0), .b(s_186), .O(gate86inter1));
  and2  gate1851(.a(G332), .b(G8), .O(gate86inter2));
  inv1  gate1852(.a(s_186), .O(gate86inter3));
  inv1  gate1853(.a(s_187), .O(gate86inter4));
  nand2 gate1854(.a(gate86inter4), .b(gate86inter3), .O(gate86inter5));
  nor2  gate1855(.a(gate86inter5), .b(gate86inter2), .O(gate86inter6));
  inv1  gate1856(.a(G8), .O(gate86inter7));
  inv1  gate1857(.a(G332), .O(gate86inter8));
  nand2 gate1858(.a(gate86inter8), .b(gate86inter7), .O(gate86inter9));
  nand2 gate1859(.a(s_187), .b(gate86inter3), .O(gate86inter10));
  nor2  gate1860(.a(gate86inter10), .b(gate86inter9), .O(gate86inter11));
  nor2  gate1861(.a(gate86inter11), .b(gate86inter6), .O(gate86inter12));
  nand2 gate1862(.a(gate86inter12), .b(gate86inter1), .O(G407));

  xor2  gate1625(.a(G335), .b(G12), .O(gate87inter0));
  nand2 gate1626(.a(gate87inter0), .b(s_154), .O(gate87inter1));
  and2  gate1627(.a(G335), .b(G12), .O(gate87inter2));
  inv1  gate1628(.a(s_154), .O(gate87inter3));
  inv1  gate1629(.a(s_155), .O(gate87inter4));
  nand2 gate1630(.a(gate87inter4), .b(gate87inter3), .O(gate87inter5));
  nor2  gate1631(.a(gate87inter5), .b(gate87inter2), .O(gate87inter6));
  inv1  gate1632(.a(G12), .O(gate87inter7));
  inv1  gate1633(.a(G335), .O(gate87inter8));
  nand2 gate1634(.a(gate87inter8), .b(gate87inter7), .O(gate87inter9));
  nand2 gate1635(.a(s_155), .b(gate87inter3), .O(gate87inter10));
  nor2  gate1636(.a(gate87inter10), .b(gate87inter9), .O(gate87inter11));
  nor2  gate1637(.a(gate87inter11), .b(gate87inter6), .O(gate87inter12));
  nand2 gate1638(.a(gate87inter12), .b(gate87inter1), .O(G408));
nand2 gate88( .a(G16), .b(G335), .O(G409) );
nand2 gate89( .a(G17), .b(G338), .O(G410) );
nand2 gate90( .a(G21), .b(G338), .O(G411) );
nand2 gate91( .a(G25), .b(G341), .O(G412) );
nand2 gate92( .a(G29), .b(G341), .O(G413) );
nand2 gate93( .a(G18), .b(G344), .O(G414) );
nand2 gate94( .a(G22), .b(G344), .O(G415) );

  xor2  gate715(.a(G347), .b(G26), .O(gate95inter0));
  nand2 gate716(.a(gate95inter0), .b(s_24), .O(gate95inter1));
  and2  gate717(.a(G347), .b(G26), .O(gate95inter2));
  inv1  gate718(.a(s_24), .O(gate95inter3));
  inv1  gate719(.a(s_25), .O(gate95inter4));
  nand2 gate720(.a(gate95inter4), .b(gate95inter3), .O(gate95inter5));
  nor2  gate721(.a(gate95inter5), .b(gate95inter2), .O(gate95inter6));
  inv1  gate722(.a(G26), .O(gate95inter7));
  inv1  gate723(.a(G347), .O(gate95inter8));
  nand2 gate724(.a(gate95inter8), .b(gate95inter7), .O(gate95inter9));
  nand2 gate725(.a(s_25), .b(gate95inter3), .O(gate95inter10));
  nor2  gate726(.a(gate95inter10), .b(gate95inter9), .O(gate95inter11));
  nor2  gate727(.a(gate95inter11), .b(gate95inter6), .O(gate95inter12));
  nand2 gate728(.a(gate95inter12), .b(gate95inter1), .O(G416));
nand2 gate96( .a(G30), .b(G347), .O(G417) );
nand2 gate97( .a(G19), .b(G350), .O(G418) );
nand2 gate98( .a(G23), .b(G350), .O(G419) );

  xor2  gate1331(.a(G353), .b(G27), .O(gate99inter0));
  nand2 gate1332(.a(gate99inter0), .b(s_112), .O(gate99inter1));
  and2  gate1333(.a(G353), .b(G27), .O(gate99inter2));
  inv1  gate1334(.a(s_112), .O(gate99inter3));
  inv1  gate1335(.a(s_113), .O(gate99inter4));
  nand2 gate1336(.a(gate99inter4), .b(gate99inter3), .O(gate99inter5));
  nor2  gate1337(.a(gate99inter5), .b(gate99inter2), .O(gate99inter6));
  inv1  gate1338(.a(G27), .O(gate99inter7));
  inv1  gate1339(.a(G353), .O(gate99inter8));
  nand2 gate1340(.a(gate99inter8), .b(gate99inter7), .O(gate99inter9));
  nand2 gate1341(.a(s_113), .b(gate99inter3), .O(gate99inter10));
  nor2  gate1342(.a(gate99inter10), .b(gate99inter9), .O(gate99inter11));
  nor2  gate1343(.a(gate99inter11), .b(gate99inter6), .O(gate99inter12));
  nand2 gate1344(.a(gate99inter12), .b(gate99inter1), .O(G420));
nand2 gate100( .a(G31), .b(G353), .O(G421) );

  xor2  gate1471(.a(G356), .b(G20), .O(gate101inter0));
  nand2 gate1472(.a(gate101inter0), .b(s_132), .O(gate101inter1));
  and2  gate1473(.a(G356), .b(G20), .O(gate101inter2));
  inv1  gate1474(.a(s_132), .O(gate101inter3));
  inv1  gate1475(.a(s_133), .O(gate101inter4));
  nand2 gate1476(.a(gate101inter4), .b(gate101inter3), .O(gate101inter5));
  nor2  gate1477(.a(gate101inter5), .b(gate101inter2), .O(gate101inter6));
  inv1  gate1478(.a(G20), .O(gate101inter7));
  inv1  gate1479(.a(G356), .O(gate101inter8));
  nand2 gate1480(.a(gate101inter8), .b(gate101inter7), .O(gate101inter9));
  nand2 gate1481(.a(s_133), .b(gate101inter3), .O(gate101inter10));
  nor2  gate1482(.a(gate101inter10), .b(gate101inter9), .O(gate101inter11));
  nor2  gate1483(.a(gate101inter11), .b(gate101inter6), .O(gate101inter12));
  nand2 gate1484(.a(gate101inter12), .b(gate101inter1), .O(G422));
nand2 gate102( .a(G24), .b(G356), .O(G423) );
nand2 gate103( .a(G28), .b(G359), .O(G424) );
nand2 gate104( .a(G32), .b(G359), .O(G425) );
nand2 gate105( .a(G362), .b(G363), .O(G426) );

  xor2  gate1037(.a(G365), .b(G364), .O(gate106inter0));
  nand2 gate1038(.a(gate106inter0), .b(s_70), .O(gate106inter1));
  and2  gate1039(.a(G365), .b(G364), .O(gate106inter2));
  inv1  gate1040(.a(s_70), .O(gate106inter3));
  inv1  gate1041(.a(s_71), .O(gate106inter4));
  nand2 gate1042(.a(gate106inter4), .b(gate106inter3), .O(gate106inter5));
  nor2  gate1043(.a(gate106inter5), .b(gate106inter2), .O(gate106inter6));
  inv1  gate1044(.a(G364), .O(gate106inter7));
  inv1  gate1045(.a(G365), .O(gate106inter8));
  nand2 gate1046(.a(gate106inter8), .b(gate106inter7), .O(gate106inter9));
  nand2 gate1047(.a(s_71), .b(gate106inter3), .O(gate106inter10));
  nor2  gate1048(.a(gate106inter10), .b(gate106inter9), .O(gate106inter11));
  nor2  gate1049(.a(gate106inter11), .b(gate106inter6), .O(gate106inter12));
  nand2 gate1050(.a(gate106inter12), .b(gate106inter1), .O(G429));
nand2 gate107( .a(G366), .b(G367), .O(G432) );
nand2 gate108( .a(G368), .b(G369), .O(G435) );
nand2 gate109( .a(G370), .b(G371), .O(G438) );
nand2 gate110( .a(G372), .b(G373), .O(G441) );
nand2 gate111( .a(G374), .b(G375), .O(G444) );
nand2 gate112( .a(G376), .b(G377), .O(G447) );
nand2 gate113( .a(G378), .b(G379), .O(G450) );
nand2 gate114( .a(G380), .b(G381), .O(G453) );

  xor2  gate1261(.a(G383), .b(G382), .O(gate115inter0));
  nand2 gate1262(.a(gate115inter0), .b(s_102), .O(gate115inter1));
  and2  gate1263(.a(G383), .b(G382), .O(gate115inter2));
  inv1  gate1264(.a(s_102), .O(gate115inter3));
  inv1  gate1265(.a(s_103), .O(gate115inter4));
  nand2 gate1266(.a(gate115inter4), .b(gate115inter3), .O(gate115inter5));
  nor2  gate1267(.a(gate115inter5), .b(gate115inter2), .O(gate115inter6));
  inv1  gate1268(.a(G382), .O(gate115inter7));
  inv1  gate1269(.a(G383), .O(gate115inter8));
  nand2 gate1270(.a(gate115inter8), .b(gate115inter7), .O(gate115inter9));
  nand2 gate1271(.a(s_103), .b(gate115inter3), .O(gate115inter10));
  nor2  gate1272(.a(gate115inter10), .b(gate115inter9), .O(gate115inter11));
  nor2  gate1273(.a(gate115inter11), .b(gate115inter6), .O(gate115inter12));
  nand2 gate1274(.a(gate115inter12), .b(gate115inter1), .O(G456));
nand2 gate116( .a(G384), .b(G385), .O(G459) );
nand2 gate117( .a(G386), .b(G387), .O(G462) );
nand2 gate118( .a(G388), .b(G389), .O(G465) );
nand2 gate119( .a(G390), .b(G391), .O(G468) );
nand2 gate120( .a(G392), .b(G393), .O(G471) );
nand2 gate121( .a(G394), .b(G395), .O(G474) );

  xor2  gate2115(.a(G397), .b(G396), .O(gate122inter0));
  nand2 gate2116(.a(gate122inter0), .b(s_224), .O(gate122inter1));
  and2  gate2117(.a(G397), .b(G396), .O(gate122inter2));
  inv1  gate2118(.a(s_224), .O(gate122inter3));
  inv1  gate2119(.a(s_225), .O(gate122inter4));
  nand2 gate2120(.a(gate122inter4), .b(gate122inter3), .O(gate122inter5));
  nor2  gate2121(.a(gate122inter5), .b(gate122inter2), .O(gate122inter6));
  inv1  gate2122(.a(G396), .O(gate122inter7));
  inv1  gate2123(.a(G397), .O(gate122inter8));
  nand2 gate2124(.a(gate122inter8), .b(gate122inter7), .O(gate122inter9));
  nand2 gate2125(.a(s_225), .b(gate122inter3), .O(gate122inter10));
  nor2  gate2126(.a(gate122inter10), .b(gate122inter9), .O(gate122inter11));
  nor2  gate2127(.a(gate122inter11), .b(gate122inter6), .O(gate122inter12));
  nand2 gate2128(.a(gate122inter12), .b(gate122inter1), .O(G477));
nand2 gate123( .a(G398), .b(G399), .O(G480) );
nand2 gate124( .a(G400), .b(G401), .O(G483) );
nand2 gate125( .a(G402), .b(G403), .O(G486) );

  xor2  gate1373(.a(G405), .b(G404), .O(gate126inter0));
  nand2 gate1374(.a(gate126inter0), .b(s_118), .O(gate126inter1));
  and2  gate1375(.a(G405), .b(G404), .O(gate126inter2));
  inv1  gate1376(.a(s_118), .O(gate126inter3));
  inv1  gate1377(.a(s_119), .O(gate126inter4));
  nand2 gate1378(.a(gate126inter4), .b(gate126inter3), .O(gate126inter5));
  nor2  gate1379(.a(gate126inter5), .b(gate126inter2), .O(gate126inter6));
  inv1  gate1380(.a(G404), .O(gate126inter7));
  inv1  gate1381(.a(G405), .O(gate126inter8));
  nand2 gate1382(.a(gate126inter8), .b(gate126inter7), .O(gate126inter9));
  nand2 gate1383(.a(s_119), .b(gate126inter3), .O(gate126inter10));
  nor2  gate1384(.a(gate126inter10), .b(gate126inter9), .O(gate126inter11));
  nor2  gate1385(.a(gate126inter11), .b(gate126inter6), .O(gate126inter12));
  nand2 gate1386(.a(gate126inter12), .b(gate126inter1), .O(G489));

  xor2  gate2073(.a(G407), .b(G406), .O(gate127inter0));
  nand2 gate2074(.a(gate127inter0), .b(s_218), .O(gate127inter1));
  and2  gate2075(.a(G407), .b(G406), .O(gate127inter2));
  inv1  gate2076(.a(s_218), .O(gate127inter3));
  inv1  gate2077(.a(s_219), .O(gate127inter4));
  nand2 gate2078(.a(gate127inter4), .b(gate127inter3), .O(gate127inter5));
  nor2  gate2079(.a(gate127inter5), .b(gate127inter2), .O(gate127inter6));
  inv1  gate2080(.a(G406), .O(gate127inter7));
  inv1  gate2081(.a(G407), .O(gate127inter8));
  nand2 gate2082(.a(gate127inter8), .b(gate127inter7), .O(gate127inter9));
  nand2 gate2083(.a(s_219), .b(gate127inter3), .O(gate127inter10));
  nor2  gate2084(.a(gate127inter10), .b(gate127inter9), .O(gate127inter11));
  nor2  gate2085(.a(gate127inter11), .b(gate127inter6), .O(gate127inter12));
  nand2 gate2086(.a(gate127inter12), .b(gate127inter1), .O(G492));
nand2 gate128( .a(G408), .b(G409), .O(G495) );
nand2 gate129( .a(G410), .b(G411), .O(G498) );

  xor2  gate995(.a(G413), .b(G412), .O(gate130inter0));
  nand2 gate996(.a(gate130inter0), .b(s_64), .O(gate130inter1));
  and2  gate997(.a(G413), .b(G412), .O(gate130inter2));
  inv1  gate998(.a(s_64), .O(gate130inter3));
  inv1  gate999(.a(s_65), .O(gate130inter4));
  nand2 gate1000(.a(gate130inter4), .b(gate130inter3), .O(gate130inter5));
  nor2  gate1001(.a(gate130inter5), .b(gate130inter2), .O(gate130inter6));
  inv1  gate1002(.a(G412), .O(gate130inter7));
  inv1  gate1003(.a(G413), .O(gate130inter8));
  nand2 gate1004(.a(gate130inter8), .b(gate130inter7), .O(gate130inter9));
  nand2 gate1005(.a(s_65), .b(gate130inter3), .O(gate130inter10));
  nor2  gate1006(.a(gate130inter10), .b(gate130inter9), .O(gate130inter11));
  nor2  gate1007(.a(gate130inter11), .b(gate130inter6), .O(gate130inter12));
  nand2 gate1008(.a(gate130inter12), .b(gate130inter1), .O(G501));

  xor2  gate1205(.a(G415), .b(G414), .O(gate131inter0));
  nand2 gate1206(.a(gate131inter0), .b(s_94), .O(gate131inter1));
  and2  gate1207(.a(G415), .b(G414), .O(gate131inter2));
  inv1  gate1208(.a(s_94), .O(gate131inter3));
  inv1  gate1209(.a(s_95), .O(gate131inter4));
  nand2 gate1210(.a(gate131inter4), .b(gate131inter3), .O(gate131inter5));
  nor2  gate1211(.a(gate131inter5), .b(gate131inter2), .O(gate131inter6));
  inv1  gate1212(.a(G414), .O(gate131inter7));
  inv1  gate1213(.a(G415), .O(gate131inter8));
  nand2 gate1214(.a(gate131inter8), .b(gate131inter7), .O(gate131inter9));
  nand2 gate1215(.a(s_95), .b(gate131inter3), .O(gate131inter10));
  nor2  gate1216(.a(gate131inter10), .b(gate131inter9), .O(gate131inter11));
  nor2  gate1217(.a(gate131inter11), .b(gate131inter6), .O(gate131inter12));
  nand2 gate1218(.a(gate131inter12), .b(gate131inter1), .O(G504));
nand2 gate132( .a(G416), .b(G417), .O(G507) );
nand2 gate133( .a(G418), .b(G419), .O(G510) );
nand2 gate134( .a(G420), .b(G421), .O(G513) );
nand2 gate135( .a(G422), .b(G423), .O(G516) );
nand2 gate136( .a(G424), .b(G425), .O(G519) );
nand2 gate137( .a(G426), .b(G429), .O(G522) );
nand2 gate138( .a(G432), .b(G435), .O(G525) );
nand2 gate139( .a(G438), .b(G441), .O(G528) );
nand2 gate140( .a(G444), .b(G447), .O(G531) );
nand2 gate141( .a(G450), .b(G453), .O(G534) );
nand2 gate142( .a(G456), .b(G459), .O(G537) );
nand2 gate143( .a(G462), .b(G465), .O(G540) );

  xor2  gate1429(.a(G471), .b(G468), .O(gate144inter0));
  nand2 gate1430(.a(gate144inter0), .b(s_126), .O(gate144inter1));
  and2  gate1431(.a(G471), .b(G468), .O(gate144inter2));
  inv1  gate1432(.a(s_126), .O(gate144inter3));
  inv1  gate1433(.a(s_127), .O(gate144inter4));
  nand2 gate1434(.a(gate144inter4), .b(gate144inter3), .O(gate144inter5));
  nor2  gate1435(.a(gate144inter5), .b(gate144inter2), .O(gate144inter6));
  inv1  gate1436(.a(G468), .O(gate144inter7));
  inv1  gate1437(.a(G471), .O(gate144inter8));
  nand2 gate1438(.a(gate144inter8), .b(gate144inter7), .O(gate144inter9));
  nand2 gate1439(.a(s_127), .b(gate144inter3), .O(gate144inter10));
  nor2  gate1440(.a(gate144inter10), .b(gate144inter9), .O(gate144inter11));
  nor2  gate1441(.a(gate144inter11), .b(gate144inter6), .O(gate144inter12));
  nand2 gate1442(.a(gate144inter12), .b(gate144inter1), .O(G543));

  xor2  gate1989(.a(G477), .b(G474), .O(gate145inter0));
  nand2 gate1990(.a(gate145inter0), .b(s_206), .O(gate145inter1));
  and2  gate1991(.a(G477), .b(G474), .O(gate145inter2));
  inv1  gate1992(.a(s_206), .O(gate145inter3));
  inv1  gate1993(.a(s_207), .O(gate145inter4));
  nand2 gate1994(.a(gate145inter4), .b(gate145inter3), .O(gate145inter5));
  nor2  gate1995(.a(gate145inter5), .b(gate145inter2), .O(gate145inter6));
  inv1  gate1996(.a(G474), .O(gate145inter7));
  inv1  gate1997(.a(G477), .O(gate145inter8));
  nand2 gate1998(.a(gate145inter8), .b(gate145inter7), .O(gate145inter9));
  nand2 gate1999(.a(s_207), .b(gate145inter3), .O(gate145inter10));
  nor2  gate2000(.a(gate145inter10), .b(gate145inter9), .O(gate145inter11));
  nor2  gate2001(.a(gate145inter11), .b(gate145inter6), .O(gate145inter12));
  nand2 gate2002(.a(gate145inter12), .b(gate145inter1), .O(G546));

  xor2  gate1779(.a(G483), .b(G480), .O(gate146inter0));
  nand2 gate1780(.a(gate146inter0), .b(s_176), .O(gate146inter1));
  and2  gate1781(.a(G483), .b(G480), .O(gate146inter2));
  inv1  gate1782(.a(s_176), .O(gate146inter3));
  inv1  gate1783(.a(s_177), .O(gate146inter4));
  nand2 gate1784(.a(gate146inter4), .b(gate146inter3), .O(gate146inter5));
  nor2  gate1785(.a(gate146inter5), .b(gate146inter2), .O(gate146inter6));
  inv1  gate1786(.a(G480), .O(gate146inter7));
  inv1  gate1787(.a(G483), .O(gate146inter8));
  nand2 gate1788(.a(gate146inter8), .b(gate146inter7), .O(gate146inter9));
  nand2 gate1789(.a(s_177), .b(gate146inter3), .O(gate146inter10));
  nor2  gate1790(.a(gate146inter10), .b(gate146inter9), .O(gate146inter11));
  nor2  gate1791(.a(gate146inter11), .b(gate146inter6), .O(gate146inter12));
  nand2 gate1792(.a(gate146inter12), .b(gate146inter1), .O(G549));
nand2 gate147( .a(G486), .b(G489), .O(G552) );

  xor2  gate659(.a(G495), .b(G492), .O(gate148inter0));
  nand2 gate660(.a(gate148inter0), .b(s_16), .O(gate148inter1));
  and2  gate661(.a(G495), .b(G492), .O(gate148inter2));
  inv1  gate662(.a(s_16), .O(gate148inter3));
  inv1  gate663(.a(s_17), .O(gate148inter4));
  nand2 gate664(.a(gate148inter4), .b(gate148inter3), .O(gate148inter5));
  nor2  gate665(.a(gate148inter5), .b(gate148inter2), .O(gate148inter6));
  inv1  gate666(.a(G492), .O(gate148inter7));
  inv1  gate667(.a(G495), .O(gate148inter8));
  nand2 gate668(.a(gate148inter8), .b(gate148inter7), .O(gate148inter9));
  nand2 gate669(.a(s_17), .b(gate148inter3), .O(gate148inter10));
  nor2  gate670(.a(gate148inter10), .b(gate148inter9), .O(gate148inter11));
  nor2  gate671(.a(gate148inter11), .b(gate148inter6), .O(gate148inter12));
  nand2 gate672(.a(gate148inter12), .b(gate148inter1), .O(G555));
nand2 gate149( .a(G498), .b(G501), .O(G558) );
nand2 gate150( .a(G504), .b(G507), .O(G561) );
nand2 gate151( .a(G510), .b(G513), .O(G564) );
nand2 gate152( .a(G516), .b(G519), .O(G567) );

  xor2  gate771(.a(G522), .b(G426), .O(gate153inter0));
  nand2 gate772(.a(gate153inter0), .b(s_32), .O(gate153inter1));
  and2  gate773(.a(G522), .b(G426), .O(gate153inter2));
  inv1  gate774(.a(s_32), .O(gate153inter3));
  inv1  gate775(.a(s_33), .O(gate153inter4));
  nand2 gate776(.a(gate153inter4), .b(gate153inter3), .O(gate153inter5));
  nor2  gate777(.a(gate153inter5), .b(gate153inter2), .O(gate153inter6));
  inv1  gate778(.a(G426), .O(gate153inter7));
  inv1  gate779(.a(G522), .O(gate153inter8));
  nand2 gate780(.a(gate153inter8), .b(gate153inter7), .O(gate153inter9));
  nand2 gate781(.a(s_33), .b(gate153inter3), .O(gate153inter10));
  nor2  gate782(.a(gate153inter10), .b(gate153inter9), .O(gate153inter11));
  nor2  gate783(.a(gate153inter11), .b(gate153inter6), .O(gate153inter12));
  nand2 gate784(.a(gate153inter12), .b(gate153inter1), .O(G570));
nand2 gate154( .a(G429), .b(G522), .O(G571) );

  xor2  gate1009(.a(G525), .b(G432), .O(gate155inter0));
  nand2 gate1010(.a(gate155inter0), .b(s_66), .O(gate155inter1));
  and2  gate1011(.a(G525), .b(G432), .O(gate155inter2));
  inv1  gate1012(.a(s_66), .O(gate155inter3));
  inv1  gate1013(.a(s_67), .O(gate155inter4));
  nand2 gate1014(.a(gate155inter4), .b(gate155inter3), .O(gate155inter5));
  nor2  gate1015(.a(gate155inter5), .b(gate155inter2), .O(gate155inter6));
  inv1  gate1016(.a(G432), .O(gate155inter7));
  inv1  gate1017(.a(G525), .O(gate155inter8));
  nand2 gate1018(.a(gate155inter8), .b(gate155inter7), .O(gate155inter9));
  nand2 gate1019(.a(s_67), .b(gate155inter3), .O(gate155inter10));
  nor2  gate1020(.a(gate155inter10), .b(gate155inter9), .O(gate155inter11));
  nor2  gate1021(.a(gate155inter11), .b(gate155inter6), .O(gate155inter12));
  nand2 gate1022(.a(gate155inter12), .b(gate155inter1), .O(G572));
nand2 gate156( .a(G435), .b(G525), .O(G573) );

  xor2  gate1961(.a(G528), .b(G438), .O(gate157inter0));
  nand2 gate1962(.a(gate157inter0), .b(s_202), .O(gate157inter1));
  and2  gate1963(.a(G528), .b(G438), .O(gate157inter2));
  inv1  gate1964(.a(s_202), .O(gate157inter3));
  inv1  gate1965(.a(s_203), .O(gate157inter4));
  nand2 gate1966(.a(gate157inter4), .b(gate157inter3), .O(gate157inter5));
  nor2  gate1967(.a(gate157inter5), .b(gate157inter2), .O(gate157inter6));
  inv1  gate1968(.a(G438), .O(gate157inter7));
  inv1  gate1969(.a(G528), .O(gate157inter8));
  nand2 gate1970(.a(gate157inter8), .b(gate157inter7), .O(gate157inter9));
  nand2 gate1971(.a(s_203), .b(gate157inter3), .O(gate157inter10));
  nor2  gate1972(.a(gate157inter10), .b(gate157inter9), .O(gate157inter11));
  nor2  gate1973(.a(gate157inter11), .b(gate157inter6), .O(gate157inter12));
  nand2 gate1974(.a(gate157inter12), .b(gate157inter1), .O(G574));
nand2 gate158( .a(G441), .b(G528), .O(G575) );
nand2 gate159( .a(G444), .b(G531), .O(G576) );
nand2 gate160( .a(G447), .b(G531), .O(G577) );

  xor2  gate561(.a(G534), .b(G450), .O(gate161inter0));
  nand2 gate562(.a(gate161inter0), .b(s_2), .O(gate161inter1));
  and2  gate563(.a(G534), .b(G450), .O(gate161inter2));
  inv1  gate564(.a(s_2), .O(gate161inter3));
  inv1  gate565(.a(s_3), .O(gate161inter4));
  nand2 gate566(.a(gate161inter4), .b(gate161inter3), .O(gate161inter5));
  nor2  gate567(.a(gate161inter5), .b(gate161inter2), .O(gate161inter6));
  inv1  gate568(.a(G450), .O(gate161inter7));
  inv1  gate569(.a(G534), .O(gate161inter8));
  nand2 gate570(.a(gate161inter8), .b(gate161inter7), .O(gate161inter9));
  nand2 gate571(.a(s_3), .b(gate161inter3), .O(gate161inter10));
  nor2  gate572(.a(gate161inter10), .b(gate161inter9), .O(gate161inter11));
  nor2  gate573(.a(gate161inter11), .b(gate161inter6), .O(gate161inter12));
  nand2 gate574(.a(gate161inter12), .b(gate161inter1), .O(G578));

  xor2  gate2157(.a(G534), .b(G453), .O(gate162inter0));
  nand2 gate2158(.a(gate162inter0), .b(s_230), .O(gate162inter1));
  and2  gate2159(.a(G534), .b(G453), .O(gate162inter2));
  inv1  gate2160(.a(s_230), .O(gate162inter3));
  inv1  gate2161(.a(s_231), .O(gate162inter4));
  nand2 gate2162(.a(gate162inter4), .b(gate162inter3), .O(gate162inter5));
  nor2  gate2163(.a(gate162inter5), .b(gate162inter2), .O(gate162inter6));
  inv1  gate2164(.a(G453), .O(gate162inter7));
  inv1  gate2165(.a(G534), .O(gate162inter8));
  nand2 gate2166(.a(gate162inter8), .b(gate162inter7), .O(gate162inter9));
  nand2 gate2167(.a(s_231), .b(gate162inter3), .O(gate162inter10));
  nor2  gate2168(.a(gate162inter10), .b(gate162inter9), .O(gate162inter11));
  nor2  gate2169(.a(gate162inter11), .b(gate162inter6), .O(gate162inter12));
  nand2 gate2170(.a(gate162inter12), .b(gate162inter1), .O(G579));
nand2 gate163( .a(G456), .b(G537), .O(G580) );
nand2 gate164( .a(G459), .b(G537), .O(G581) );

  xor2  gate1751(.a(G540), .b(G462), .O(gate165inter0));
  nand2 gate1752(.a(gate165inter0), .b(s_172), .O(gate165inter1));
  and2  gate1753(.a(G540), .b(G462), .O(gate165inter2));
  inv1  gate1754(.a(s_172), .O(gate165inter3));
  inv1  gate1755(.a(s_173), .O(gate165inter4));
  nand2 gate1756(.a(gate165inter4), .b(gate165inter3), .O(gate165inter5));
  nor2  gate1757(.a(gate165inter5), .b(gate165inter2), .O(gate165inter6));
  inv1  gate1758(.a(G462), .O(gate165inter7));
  inv1  gate1759(.a(G540), .O(gate165inter8));
  nand2 gate1760(.a(gate165inter8), .b(gate165inter7), .O(gate165inter9));
  nand2 gate1761(.a(s_173), .b(gate165inter3), .O(gate165inter10));
  nor2  gate1762(.a(gate165inter10), .b(gate165inter9), .O(gate165inter11));
  nor2  gate1763(.a(gate165inter11), .b(gate165inter6), .O(gate165inter12));
  nand2 gate1764(.a(gate165inter12), .b(gate165inter1), .O(G582));
nand2 gate166( .a(G465), .b(G540), .O(G583) );
nand2 gate167( .a(G468), .b(G543), .O(G584) );
nand2 gate168( .a(G471), .b(G543), .O(G585) );

  xor2  gate2283(.a(G546), .b(G474), .O(gate169inter0));
  nand2 gate2284(.a(gate169inter0), .b(s_248), .O(gate169inter1));
  and2  gate2285(.a(G546), .b(G474), .O(gate169inter2));
  inv1  gate2286(.a(s_248), .O(gate169inter3));
  inv1  gate2287(.a(s_249), .O(gate169inter4));
  nand2 gate2288(.a(gate169inter4), .b(gate169inter3), .O(gate169inter5));
  nor2  gate2289(.a(gate169inter5), .b(gate169inter2), .O(gate169inter6));
  inv1  gate2290(.a(G474), .O(gate169inter7));
  inv1  gate2291(.a(G546), .O(gate169inter8));
  nand2 gate2292(.a(gate169inter8), .b(gate169inter7), .O(gate169inter9));
  nand2 gate2293(.a(s_249), .b(gate169inter3), .O(gate169inter10));
  nor2  gate2294(.a(gate169inter10), .b(gate169inter9), .O(gate169inter11));
  nor2  gate2295(.a(gate169inter11), .b(gate169inter6), .O(gate169inter12));
  nand2 gate2296(.a(gate169inter12), .b(gate169inter1), .O(G586));

  xor2  gate1639(.a(G546), .b(G477), .O(gate170inter0));
  nand2 gate1640(.a(gate170inter0), .b(s_156), .O(gate170inter1));
  and2  gate1641(.a(G546), .b(G477), .O(gate170inter2));
  inv1  gate1642(.a(s_156), .O(gate170inter3));
  inv1  gate1643(.a(s_157), .O(gate170inter4));
  nand2 gate1644(.a(gate170inter4), .b(gate170inter3), .O(gate170inter5));
  nor2  gate1645(.a(gate170inter5), .b(gate170inter2), .O(gate170inter6));
  inv1  gate1646(.a(G477), .O(gate170inter7));
  inv1  gate1647(.a(G546), .O(gate170inter8));
  nand2 gate1648(.a(gate170inter8), .b(gate170inter7), .O(gate170inter9));
  nand2 gate1649(.a(s_157), .b(gate170inter3), .O(gate170inter10));
  nor2  gate1650(.a(gate170inter10), .b(gate170inter9), .O(gate170inter11));
  nor2  gate1651(.a(gate170inter11), .b(gate170inter6), .O(gate170inter12));
  nand2 gate1652(.a(gate170inter12), .b(gate170inter1), .O(G587));
nand2 gate171( .a(G480), .b(G549), .O(G588) );
nand2 gate172( .a(G483), .b(G549), .O(G589) );
nand2 gate173( .a(G486), .b(G552), .O(G590) );

  xor2  gate1695(.a(G552), .b(G489), .O(gate174inter0));
  nand2 gate1696(.a(gate174inter0), .b(s_164), .O(gate174inter1));
  and2  gate1697(.a(G552), .b(G489), .O(gate174inter2));
  inv1  gate1698(.a(s_164), .O(gate174inter3));
  inv1  gate1699(.a(s_165), .O(gate174inter4));
  nand2 gate1700(.a(gate174inter4), .b(gate174inter3), .O(gate174inter5));
  nor2  gate1701(.a(gate174inter5), .b(gate174inter2), .O(gate174inter6));
  inv1  gate1702(.a(G489), .O(gate174inter7));
  inv1  gate1703(.a(G552), .O(gate174inter8));
  nand2 gate1704(.a(gate174inter8), .b(gate174inter7), .O(gate174inter9));
  nand2 gate1705(.a(s_165), .b(gate174inter3), .O(gate174inter10));
  nor2  gate1706(.a(gate174inter10), .b(gate174inter9), .O(gate174inter11));
  nor2  gate1707(.a(gate174inter11), .b(gate174inter6), .O(gate174inter12));
  nand2 gate1708(.a(gate174inter12), .b(gate174inter1), .O(G591));
nand2 gate175( .a(G492), .b(G555), .O(G592) );
nand2 gate176( .a(G495), .b(G555), .O(G593) );
nand2 gate177( .a(G498), .b(G558), .O(G594) );
nand2 gate178( .a(G501), .b(G558), .O(G595) );
nand2 gate179( .a(G504), .b(G561), .O(G596) );
nand2 gate180( .a(G507), .b(G561), .O(G597) );

  xor2  gate1359(.a(G564), .b(G510), .O(gate181inter0));
  nand2 gate1360(.a(gate181inter0), .b(s_116), .O(gate181inter1));
  and2  gate1361(.a(G564), .b(G510), .O(gate181inter2));
  inv1  gate1362(.a(s_116), .O(gate181inter3));
  inv1  gate1363(.a(s_117), .O(gate181inter4));
  nand2 gate1364(.a(gate181inter4), .b(gate181inter3), .O(gate181inter5));
  nor2  gate1365(.a(gate181inter5), .b(gate181inter2), .O(gate181inter6));
  inv1  gate1366(.a(G510), .O(gate181inter7));
  inv1  gate1367(.a(G564), .O(gate181inter8));
  nand2 gate1368(.a(gate181inter8), .b(gate181inter7), .O(gate181inter9));
  nand2 gate1369(.a(s_117), .b(gate181inter3), .O(gate181inter10));
  nor2  gate1370(.a(gate181inter10), .b(gate181inter9), .O(gate181inter11));
  nor2  gate1371(.a(gate181inter11), .b(gate181inter6), .O(gate181inter12));
  nand2 gate1372(.a(gate181inter12), .b(gate181inter1), .O(G598));
nand2 gate182( .a(G513), .b(G564), .O(G599) );
nand2 gate183( .a(G516), .b(G567), .O(G600) );
nand2 gate184( .a(G519), .b(G567), .O(G601) );
nand2 gate185( .a(G570), .b(G571), .O(G602) );
nand2 gate186( .a(G572), .b(G573), .O(G607) );

  xor2  gate687(.a(G575), .b(G574), .O(gate187inter0));
  nand2 gate688(.a(gate187inter0), .b(s_20), .O(gate187inter1));
  and2  gate689(.a(G575), .b(G574), .O(gate187inter2));
  inv1  gate690(.a(s_20), .O(gate187inter3));
  inv1  gate691(.a(s_21), .O(gate187inter4));
  nand2 gate692(.a(gate187inter4), .b(gate187inter3), .O(gate187inter5));
  nor2  gate693(.a(gate187inter5), .b(gate187inter2), .O(gate187inter6));
  inv1  gate694(.a(G574), .O(gate187inter7));
  inv1  gate695(.a(G575), .O(gate187inter8));
  nand2 gate696(.a(gate187inter8), .b(gate187inter7), .O(gate187inter9));
  nand2 gate697(.a(s_21), .b(gate187inter3), .O(gate187inter10));
  nor2  gate698(.a(gate187inter10), .b(gate187inter9), .O(gate187inter11));
  nor2  gate699(.a(gate187inter11), .b(gate187inter6), .O(gate187inter12));
  nand2 gate700(.a(gate187inter12), .b(gate187inter1), .O(G612));

  xor2  gate1499(.a(G577), .b(G576), .O(gate188inter0));
  nand2 gate1500(.a(gate188inter0), .b(s_136), .O(gate188inter1));
  and2  gate1501(.a(G577), .b(G576), .O(gate188inter2));
  inv1  gate1502(.a(s_136), .O(gate188inter3));
  inv1  gate1503(.a(s_137), .O(gate188inter4));
  nand2 gate1504(.a(gate188inter4), .b(gate188inter3), .O(gate188inter5));
  nor2  gate1505(.a(gate188inter5), .b(gate188inter2), .O(gate188inter6));
  inv1  gate1506(.a(G576), .O(gate188inter7));
  inv1  gate1507(.a(G577), .O(gate188inter8));
  nand2 gate1508(.a(gate188inter8), .b(gate188inter7), .O(gate188inter9));
  nand2 gate1509(.a(s_137), .b(gate188inter3), .O(gate188inter10));
  nor2  gate1510(.a(gate188inter10), .b(gate188inter9), .O(gate188inter11));
  nor2  gate1511(.a(gate188inter11), .b(gate188inter6), .O(gate188inter12));
  nand2 gate1512(.a(gate188inter12), .b(gate188inter1), .O(G617));

  xor2  gate799(.a(G579), .b(G578), .O(gate189inter0));
  nand2 gate800(.a(gate189inter0), .b(s_36), .O(gate189inter1));
  and2  gate801(.a(G579), .b(G578), .O(gate189inter2));
  inv1  gate802(.a(s_36), .O(gate189inter3));
  inv1  gate803(.a(s_37), .O(gate189inter4));
  nand2 gate804(.a(gate189inter4), .b(gate189inter3), .O(gate189inter5));
  nor2  gate805(.a(gate189inter5), .b(gate189inter2), .O(gate189inter6));
  inv1  gate806(.a(G578), .O(gate189inter7));
  inv1  gate807(.a(G579), .O(gate189inter8));
  nand2 gate808(.a(gate189inter8), .b(gate189inter7), .O(gate189inter9));
  nand2 gate809(.a(s_37), .b(gate189inter3), .O(gate189inter10));
  nor2  gate810(.a(gate189inter10), .b(gate189inter9), .O(gate189inter11));
  nor2  gate811(.a(gate189inter11), .b(gate189inter6), .O(gate189inter12));
  nand2 gate812(.a(gate189inter12), .b(gate189inter1), .O(G622));

  xor2  gate1667(.a(G581), .b(G580), .O(gate190inter0));
  nand2 gate1668(.a(gate190inter0), .b(s_160), .O(gate190inter1));
  and2  gate1669(.a(G581), .b(G580), .O(gate190inter2));
  inv1  gate1670(.a(s_160), .O(gate190inter3));
  inv1  gate1671(.a(s_161), .O(gate190inter4));
  nand2 gate1672(.a(gate190inter4), .b(gate190inter3), .O(gate190inter5));
  nor2  gate1673(.a(gate190inter5), .b(gate190inter2), .O(gate190inter6));
  inv1  gate1674(.a(G580), .O(gate190inter7));
  inv1  gate1675(.a(G581), .O(gate190inter8));
  nand2 gate1676(.a(gate190inter8), .b(gate190inter7), .O(gate190inter9));
  nand2 gate1677(.a(s_161), .b(gate190inter3), .O(gate190inter10));
  nor2  gate1678(.a(gate190inter10), .b(gate190inter9), .O(gate190inter11));
  nor2  gate1679(.a(gate190inter11), .b(gate190inter6), .O(gate190inter12));
  nand2 gate1680(.a(gate190inter12), .b(gate190inter1), .O(G627));

  xor2  gate2129(.a(G583), .b(G582), .O(gate191inter0));
  nand2 gate2130(.a(gate191inter0), .b(s_226), .O(gate191inter1));
  and2  gate2131(.a(G583), .b(G582), .O(gate191inter2));
  inv1  gate2132(.a(s_226), .O(gate191inter3));
  inv1  gate2133(.a(s_227), .O(gate191inter4));
  nand2 gate2134(.a(gate191inter4), .b(gate191inter3), .O(gate191inter5));
  nor2  gate2135(.a(gate191inter5), .b(gate191inter2), .O(gate191inter6));
  inv1  gate2136(.a(G582), .O(gate191inter7));
  inv1  gate2137(.a(G583), .O(gate191inter8));
  nand2 gate2138(.a(gate191inter8), .b(gate191inter7), .O(gate191inter9));
  nand2 gate2139(.a(s_227), .b(gate191inter3), .O(gate191inter10));
  nor2  gate2140(.a(gate191inter10), .b(gate191inter9), .O(gate191inter11));
  nor2  gate2141(.a(gate191inter11), .b(gate191inter6), .O(gate191inter12));
  nand2 gate2142(.a(gate191inter12), .b(gate191inter1), .O(G632));

  xor2  gate2143(.a(G585), .b(G584), .O(gate192inter0));
  nand2 gate2144(.a(gate192inter0), .b(s_228), .O(gate192inter1));
  and2  gate2145(.a(G585), .b(G584), .O(gate192inter2));
  inv1  gate2146(.a(s_228), .O(gate192inter3));
  inv1  gate2147(.a(s_229), .O(gate192inter4));
  nand2 gate2148(.a(gate192inter4), .b(gate192inter3), .O(gate192inter5));
  nor2  gate2149(.a(gate192inter5), .b(gate192inter2), .O(gate192inter6));
  inv1  gate2150(.a(G584), .O(gate192inter7));
  inv1  gate2151(.a(G585), .O(gate192inter8));
  nand2 gate2152(.a(gate192inter8), .b(gate192inter7), .O(gate192inter9));
  nand2 gate2153(.a(s_229), .b(gate192inter3), .O(gate192inter10));
  nor2  gate2154(.a(gate192inter10), .b(gate192inter9), .O(gate192inter11));
  nor2  gate2155(.a(gate192inter11), .b(gate192inter6), .O(gate192inter12));
  nand2 gate2156(.a(gate192inter12), .b(gate192inter1), .O(G637));
nand2 gate193( .a(G586), .b(G587), .O(G642) );

  xor2  gate1891(.a(G589), .b(G588), .O(gate194inter0));
  nand2 gate1892(.a(gate194inter0), .b(s_192), .O(gate194inter1));
  and2  gate1893(.a(G589), .b(G588), .O(gate194inter2));
  inv1  gate1894(.a(s_192), .O(gate194inter3));
  inv1  gate1895(.a(s_193), .O(gate194inter4));
  nand2 gate1896(.a(gate194inter4), .b(gate194inter3), .O(gate194inter5));
  nor2  gate1897(.a(gate194inter5), .b(gate194inter2), .O(gate194inter6));
  inv1  gate1898(.a(G588), .O(gate194inter7));
  inv1  gate1899(.a(G589), .O(gate194inter8));
  nand2 gate1900(.a(gate194inter8), .b(gate194inter7), .O(gate194inter9));
  nand2 gate1901(.a(s_193), .b(gate194inter3), .O(gate194inter10));
  nor2  gate1902(.a(gate194inter10), .b(gate194inter9), .O(gate194inter11));
  nor2  gate1903(.a(gate194inter11), .b(gate194inter6), .O(gate194inter12));
  nand2 gate1904(.a(gate194inter12), .b(gate194inter1), .O(G645));
nand2 gate195( .a(G590), .b(G591), .O(G648) );
nand2 gate196( .a(G592), .b(G593), .O(G651) );
nand2 gate197( .a(G594), .b(G595), .O(G654) );
nand2 gate198( .a(G596), .b(G597), .O(G657) );
nand2 gate199( .a(G598), .b(G599), .O(G660) );

  xor2  gate1191(.a(G601), .b(G600), .O(gate200inter0));
  nand2 gate1192(.a(gate200inter0), .b(s_92), .O(gate200inter1));
  and2  gate1193(.a(G601), .b(G600), .O(gate200inter2));
  inv1  gate1194(.a(s_92), .O(gate200inter3));
  inv1  gate1195(.a(s_93), .O(gate200inter4));
  nand2 gate1196(.a(gate200inter4), .b(gate200inter3), .O(gate200inter5));
  nor2  gate1197(.a(gate200inter5), .b(gate200inter2), .O(gate200inter6));
  inv1  gate1198(.a(G600), .O(gate200inter7));
  inv1  gate1199(.a(G601), .O(gate200inter8));
  nand2 gate1200(.a(gate200inter8), .b(gate200inter7), .O(gate200inter9));
  nand2 gate1201(.a(s_93), .b(gate200inter3), .O(gate200inter10));
  nor2  gate1202(.a(gate200inter10), .b(gate200inter9), .O(gate200inter11));
  nor2  gate1203(.a(gate200inter11), .b(gate200inter6), .O(gate200inter12));
  nand2 gate1204(.a(gate200inter12), .b(gate200inter1), .O(G663));

  xor2  gate2227(.a(G607), .b(G602), .O(gate201inter0));
  nand2 gate2228(.a(gate201inter0), .b(s_240), .O(gate201inter1));
  and2  gate2229(.a(G607), .b(G602), .O(gate201inter2));
  inv1  gate2230(.a(s_240), .O(gate201inter3));
  inv1  gate2231(.a(s_241), .O(gate201inter4));
  nand2 gate2232(.a(gate201inter4), .b(gate201inter3), .O(gate201inter5));
  nor2  gate2233(.a(gate201inter5), .b(gate201inter2), .O(gate201inter6));
  inv1  gate2234(.a(G602), .O(gate201inter7));
  inv1  gate2235(.a(G607), .O(gate201inter8));
  nand2 gate2236(.a(gate201inter8), .b(gate201inter7), .O(gate201inter9));
  nand2 gate2237(.a(s_241), .b(gate201inter3), .O(gate201inter10));
  nor2  gate2238(.a(gate201inter10), .b(gate201inter9), .O(gate201inter11));
  nor2  gate2239(.a(gate201inter11), .b(gate201inter6), .O(gate201inter12));
  nand2 gate2240(.a(gate201inter12), .b(gate201inter1), .O(G666));
nand2 gate202( .a(G612), .b(G617), .O(G669) );
nand2 gate203( .a(G602), .b(G612), .O(G672) );
nand2 gate204( .a(G607), .b(G617), .O(G675) );
nand2 gate205( .a(G622), .b(G627), .O(G678) );
nand2 gate206( .a(G632), .b(G637), .O(G681) );
nand2 gate207( .a(G622), .b(G632), .O(G684) );

  xor2  gate883(.a(G637), .b(G627), .O(gate208inter0));
  nand2 gate884(.a(gate208inter0), .b(s_48), .O(gate208inter1));
  and2  gate885(.a(G637), .b(G627), .O(gate208inter2));
  inv1  gate886(.a(s_48), .O(gate208inter3));
  inv1  gate887(.a(s_49), .O(gate208inter4));
  nand2 gate888(.a(gate208inter4), .b(gate208inter3), .O(gate208inter5));
  nor2  gate889(.a(gate208inter5), .b(gate208inter2), .O(gate208inter6));
  inv1  gate890(.a(G627), .O(gate208inter7));
  inv1  gate891(.a(G637), .O(gate208inter8));
  nand2 gate892(.a(gate208inter8), .b(gate208inter7), .O(gate208inter9));
  nand2 gate893(.a(s_49), .b(gate208inter3), .O(gate208inter10));
  nor2  gate894(.a(gate208inter10), .b(gate208inter9), .O(gate208inter11));
  nor2  gate895(.a(gate208inter11), .b(gate208inter6), .O(gate208inter12));
  nand2 gate896(.a(gate208inter12), .b(gate208inter1), .O(G687));
nand2 gate209( .a(G602), .b(G666), .O(G690) );
nand2 gate210( .a(G607), .b(G666), .O(G691) );
nand2 gate211( .a(G612), .b(G669), .O(G692) );

  xor2  gate2367(.a(G669), .b(G617), .O(gate212inter0));
  nand2 gate2368(.a(gate212inter0), .b(s_260), .O(gate212inter1));
  and2  gate2369(.a(G669), .b(G617), .O(gate212inter2));
  inv1  gate2370(.a(s_260), .O(gate212inter3));
  inv1  gate2371(.a(s_261), .O(gate212inter4));
  nand2 gate2372(.a(gate212inter4), .b(gate212inter3), .O(gate212inter5));
  nor2  gate2373(.a(gate212inter5), .b(gate212inter2), .O(gate212inter6));
  inv1  gate2374(.a(G617), .O(gate212inter7));
  inv1  gate2375(.a(G669), .O(gate212inter8));
  nand2 gate2376(.a(gate212inter8), .b(gate212inter7), .O(gate212inter9));
  nand2 gate2377(.a(s_261), .b(gate212inter3), .O(gate212inter10));
  nor2  gate2378(.a(gate212inter10), .b(gate212inter9), .O(gate212inter11));
  nor2  gate2379(.a(gate212inter11), .b(gate212inter6), .O(gate212inter12));
  nand2 gate2380(.a(gate212inter12), .b(gate212inter1), .O(G693));

  xor2  gate897(.a(G672), .b(G602), .O(gate213inter0));
  nand2 gate898(.a(gate213inter0), .b(s_50), .O(gate213inter1));
  and2  gate899(.a(G672), .b(G602), .O(gate213inter2));
  inv1  gate900(.a(s_50), .O(gate213inter3));
  inv1  gate901(.a(s_51), .O(gate213inter4));
  nand2 gate902(.a(gate213inter4), .b(gate213inter3), .O(gate213inter5));
  nor2  gate903(.a(gate213inter5), .b(gate213inter2), .O(gate213inter6));
  inv1  gate904(.a(G602), .O(gate213inter7));
  inv1  gate905(.a(G672), .O(gate213inter8));
  nand2 gate906(.a(gate213inter8), .b(gate213inter7), .O(gate213inter9));
  nand2 gate907(.a(s_51), .b(gate213inter3), .O(gate213inter10));
  nor2  gate908(.a(gate213inter10), .b(gate213inter9), .O(gate213inter11));
  nor2  gate909(.a(gate213inter11), .b(gate213inter6), .O(gate213inter12));
  nand2 gate910(.a(gate213inter12), .b(gate213inter1), .O(G694));
nand2 gate214( .a(G612), .b(G672), .O(G695) );

  xor2  gate1527(.a(G675), .b(G607), .O(gate215inter0));
  nand2 gate1528(.a(gate215inter0), .b(s_140), .O(gate215inter1));
  and2  gate1529(.a(G675), .b(G607), .O(gate215inter2));
  inv1  gate1530(.a(s_140), .O(gate215inter3));
  inv1  gate1531(.a(s_141), .O(gate215inter4));
  nand2 gate1532(.a(gate215inter4), .b(gate215inter3), .O(gate215inter5));
  nor2  gate1533(.a(gate215inter5), .b(gate215inter2), .O(gate215inter6));
  inv1  gate1534(.a(G607), .O(gate215inter7));
  inv1  gate1535(.a(G675), .O(gate215inter8));
  nand2 gate1536(.a(gate215inter8), .b(gate215inter7), .O(gate215inter9));
  nand2 gate1537(.a(s_141), .b(gate215inter3), .O(gate215inter10));
  nor2  gate1538(.a(gate215inter10), .b(gate215inter9), .O(gate215inter11));
  nor2  gate1539(.a(gate215inter11), .b(gate215inter6), .O(gate215inter12));
  nand2 gate1540(.a(gate215inter12), .b(gate215inter1), .O(G696));
nand2 gate216( .a(G617), .b(G675), .O(G697) );
nand2 gate217( .a(G622), .b(G678), .O(G698) );

  xor2  gate1401(.a(G678), .b(G627), .O(gate218inter0));
  nand2 gate1402(.a(gate218inter0), .b(s_122), .O(gate218inter1));
  and2  gate1403(.a(G678), .b(G627), .O(gate218inter2));
  inv1  gate1404(.a(s_122), .O(gate218inter3));
  inv1  gate1405(.a(s_123), .O(gate218inter4));
  nand2 gate1406(.a(gate218inter4), .b(gate218inter3), .O(gate218inter5));
  nor2  gate1407(.a(gate218inter5), .b(gate218inter2), .O(gate218inter6));
  inv1  gate1408(.a(G627), .O(gate218inter7));
  inv1  gate1409(.a(G678), .O(gate218inter8));
  nand2 gate1410(.a(gate218inter8), .b(gate218inter7), .O(gate218inter9));
  nand2 gate1411(.a(s_123), .b(gate218inter3), .O(gate218inter10));
  nor2  gate1412(.a(gate218inter10), .b(gate218inter9), .O(gate218inter11));
  nor2  gate1413(.a(gate218inter11), .b(gate218inter6), .O(gate218inter12));
  nand2 gate1414(.a(gate218inter12), .b(gate218inter1), .O(G699));
nand2 gate219( .a(G632), .b(G681), .O(G700) );

  xor2  gate2017(.a(G681), .b(G637), .O(gate220inter0));
  nand2 gate2018(.a(gate220inter0), .b(s_210), .O(gate220inter1));
  and2  gate2019(.a(G681), .b(G637), .O(gate220inter2));
  inv1  gate2020(.a(s_210), .O(gate220inter3));
  inv1  gate2021(.a(s_211), .O(gate220inter4));
  nand2 gate2022(.a(gate220inter4), .b(gate220inter3), .O(gate220inter5));
  nor2  gate2023(.a(gate220inter5), .b(gate220inter2), .O(gate220inter6));
  inv1  gate2024(.a(G637), .O(gate220inter7));
  inv1  gate2025(.a(G681), .O(gate220inter8));
  nand2 gate2026(.a(gate220inter8), .b(gate220inter7), .O(gate220inter9));
  nand2 gate2027(.a(s_211), .b(gate220inter3), .O(gate220inter10));
  nor2  gate2028(.a(gate220inter10), .b(gate220inter9), .O(gate220inter11));
  nor2  gate2029(.a(gate220inter11), .b(gate220inter6), .O(gate220inter12));
  nand2 gate2030(.a(gate220inter12), .b(gate220inter1), .O(G701));
nand2 gate221( .a(G622), .b(G684), .O(G702) );

  xor2  gate1289(.a(G684), .b(G632), .O(gate222inter0));
  nand2 gate1290(.a(gate222inter0), .b(s_106), .O(gate222inter1));
  and2  gate1291(.a(G684), .b(G632), .O(gate222inter2));
  inv1  gate1292(.a(s_106), .O(gate222inter3));
  inv1  gate1293(.a(s_107), .O(gate222inter4));
  nand2 gate1294(.a(gate222inter4), .b(gate222inter3), .O(gate222inter5));
  nor2  gate1295(.a(gate222inter5), .b(gate222inter2), .O(gate222inter6));
  inv1  gate1296(.a(G632), .O(gate222inter7));
  inv1  gate1297(.a(G684), .O(gate222inter8));
  nand2 gate1298(.a(gate222inter8), .b(gate222inter7), .O(gate222inter9));
  nand2 gate1299(.a(s_107), .b(gate222inter3), .O(gate222inter10));
  nor2  gate1300(.a(gate222inter10), .b(gate222inter9), .O(gate222inter11));
  nor2  gate1301(.a(gate222inter11), .b(gate222inter6), .O(gate222inter12));
  nand2 gate1302(.a(gate222inter12), .b(gate222inter1), .O(G703));
nand2 gate223( .a(G627), .b(G687), .O(G704) );
nand2 gate224( .a(G637), .b(G687), .O(G705) );
nand2 gate225( .a(G690), .b(G691), .O(G706) );
nand2 gate226( .a(G692), .b(G693), .O(G709) );
nand2 gate227( .a(G694), .b(G695), .O(G712) );

  xor2  gate1275(.a(G697), .b(G696), .O(gate228inter0));
  nand2 gate1276(.a(gate228inter0), .b(s_104), .O(gate228inter1));
  and2  gate1277(.a(G697), .b(G696), .O(gate228inter2));
  inv1  gate1278(.a(s_104), .O(gate228inter3));
  inv1  gate1279(.a(s_105), .O(gate228inter4));
  nand2 gate1280(.a(gate228inter4), .b(gate228inter3), .O(gate228inter5));
  nor2  gate1281(.a(gate228inter5), .b(gate228inter2), .O(gate228inter6));
  inv1  gate1282(.a(G696), .O(gate228inter7));
  inv1  gate1283(.a(G697), .O(gate228inter8));
  nand2 gate1284(.a(gate228inter8), .b(gate228inter7), .O(gate228inter9));
  nand2 gate1285(.a(s_105), .b(gate228inter3), .O(gate228inter10));
  nor2  gate1286(.a(gate228inter10), .b(gate228inter9), .O(gate228inter11));
  nor2  gate1287(.a(gate228inter11), .b(gate228inter6), .O(gate228inter12));
  nand2 gate1288(.a(gate228inter12), .b(gate228inter1), .O(G715));
nand2 gate229( .a(G698), .b(G699), .O(G718) );
nand2 gate230( .a(G700), .b(G701), .O(G721) );

  xor2  gate673(.a(G703), .b(G702), .O(gate231inter0));
  nand2 gate674(.a(gate231inter0), .b(s_18), .O(gate231inter1));
  and2  gate675(.a(G703), .b(G702), .O(gate231inter2));
  inv1  gate676(.a(s_18), .O(gate231inter3));
  inv1  gate677(.a(s_19), .O(gate231inter4));
  nand2 gate678(.a(gate231inter4), .b(gate231inter3), .O(gate231inter5));
  nor2  gate679(.a(gate231inter5), .b(gate231inter2), .O(gate231inter6));
  inv1  gate680(.a(G702), .O(gate231inter7));
  inv1  gate681(.a(G703), .O(gate231inter8));
  nand2 gate682(.a(gate231inter8), .b(gate231inter7), .O(gate231inter9));
  nand2 gate683(.a(s_19), .b(gate231inter3), .O(gate231inter10));
  nor2  gate684(.a(gate231inter10), .b(gate231inter9), .O(gate231inter11));
  nor2  gate685(.a(gate231inter11), .b(gate231inter6), .O(gate231inter12));
  nand2 gate686(.a(gate231inter12), .b(gate231inter1), .O(G724));
nand2 gate232( .a(G704), .b(G705), .O(G727) );

  xor2  gate1051(.a(G718), .b(G242), .O(gate233inter0));
  nand2 gate1052(.a(gate233inter0), .b(s_72), .O(gate233inter1));
  and2  gate1053(.a(G718), .b(G242), .O(gate233inter2));
  inv1  gate1054(.a(s_72), .O(gate233inter3));
  inv1  gate1055(.a(s_73), .O(gate233inter4));
  nand2 gate1056(.a(gate233inter4), .b(gate233inter3), .O(gate233inter5));
  nor2  gate1057(.a(gate233inter5), .b(gate233inter2), .O(gate233inter6));
  inv1  gate1058(.a(G242), .O(gate233inter7));
  inv1  gate1059(.a(G718), .O(gate233inter8));
  nand2 gate1060(.a(gate233inter8), .b(gate233inter7), .O(gate233inter9));
  nand2 gate1061(.a(s_73), .b(gate233inter3), .O(gate233inter10));
  nor2  gate1062(.a(gate233inter10), .b(gate233inter9), .O(gate233inter11));
  nor2  gate1063(.a(gate233inter11), .b(gate233inter6), .O(gate233inter12));
  nand2 gate1064(.a(gate233inter12), .b(gate233inter1), .O(G730));
nand2 gate234( .a(G245), .b(G721), .O(G733) );
nand2 gate235( .a(G248), .b(G724), .O(G736) );

  xor2  gate743(.a(G727), .b(G251), .O(gate236inter0));
  nand2 gate744(.a(gate236inter0), .b(s_28), .O(gate236inter1));
  and2  gate745(.a(G727), .b(G251), .O(gate236inter2));
  inv1  gate746(.a(s_28), .O(gate236inter3));
  inv1  gate747(.a(s_29), .O(gate236inter4));
  nand2 gate748(.a(gate236inter4), .b(gate236inter3), .O(gate236inter5));
  nor2  gate749(.a(gate236inter5), .b(gate236inter2), .O(gate236inter6));
  inv1  gate750(.a(G251), .O(gate236inter7));
  inv1  gate751(.a(G727), .O(gate236inter8));
  nand2 gate752(.a(gate236inter8), .b(gate236inter7), .O(gate236inter9));
  nand2 gate753(.a(s_29), .b(gate236inter3), .O(gate236inter10));
  nor2  gate754(.a(gate236inter10), .b(gate236inter9), .O(gate236inter11));
  nor2  gate755(.a(gate236inter11), .b(gate236inter6), .O(gate236inter12));
  nand2 gate756(.a(gate236inter12), .b(gate236inter1), .O(G739));

  xor2  gate1793(.a(G706), .b(G254), .O(gate237inter0));
  nand2 gate1794(.a(gate237inter0), .b(s_178), .O(gate237inter1));
  and2  gate1795(.a(G706), .b(G254), .O(gate237inter2));
  inv1  gate1796(.a(s_178), .O(gate237inter3));
  inv1  gate1797(.a(s_179), .O(gate237inter4));
  nand2 gate1798(.a(gate237inter4), .b(gate237inter3), .O(gate237inter5));
  nor2  gate1799(.a(gate237inter5), .b(gate237inter2), .O(gate237inter6));
  inv1  gate1800(.a(G254), .O(gate237inter7));
  inv1  gate1801(.a(G706), .O(gate237inter8));
  nand2 gate1802(.a(gate237inter8), .b(gate237inter7), .O(gate237inter9));
  nand2 gate1803(.a(s_179), .b(gate237inter3), .O(gate237inter10));
  nor2  gate1804(.a(gate237inter10), .b(gate237inter9), .O(gate237inter11));
  nor2  gate1805(.a(gate237inter11), .b(gate237inter6), .O(gate237inter12));
  nand2 gate1806(.a(gate237inter12), .b(gate237inter1), .O(G742));
nand2 gate238( .a(G257), .b(G709), .O(G745) );

  xor2  gate939(.a(G712), .b(G260), .O(gate239inter0));
  nand2 gate940(.a(gate239inter0), .b(s_56), .O(gate239inter1));
  and2  gate941(.a(G712), .b(G260), .O(gate239inter2));
  inv1  gate942(.a(s_56), .O(gate239inter3));
  inv1  gate943(.a(s_57), .O(gate239inter4));
  nand2 gate944(.a(gate239inter4), .b(gate239inter3), .O(gate239inter5));
  nor2  gate945(.a(gate239inter5), .b(gate239inter2), .O(gate239inter6));
  inv1  gate946(.a(G260), .O(gate239inter7));
  inv1  gate947(.a(G712), .O(gate239inter8));
  nand2 gate948(.a(gate239inter8), .b(gate239inter7), .O(gate239inter9));
  nand2 gate949(.a(s_57), .b(gate239inter3), .O(gate239inter10));
  nor2  gate950(.a(gate239inter10), .b(gate239inter9), .O(gate239inter11));
  nor2  gate951(.a(gate239inter11), .b(gate239inter6), .O(gate239inter12));
  nand2 gate952(.a(gate239inter12), .b(gate239inter1), .O(G748));
nand2 gate240( .a(G263), .b(G715), .O(G751) );

  xor2  gate729(.a(G730), .b(G242), .O(gate241inter0));
  nand2 gate730(.a(gate241inter0), .b(s_26), .O(gate241inter1));
  and2  gate731(.a(G730), .b(G242), .O(gate241inter2));
  inv1  gate732(.a(s_26), .O(gate241inter3));
  inv1  gate733(.a(s_27), .O(gate241inter4));
  nand2 gate734(.a(gate241inter4), .b(gate241inter3), .O(gate241inter5));
  nor2  gate735(.a(gate241inter5), .b(gate241inter2), .O(gate241inter6));
  inv1  gate736(.a(G242), .O(gate241inter7));
  inv1  gate737(.a(G730), .O(gate241inter8));
  nand2 gate738(.a(gate241inter8), .b(gate241inter7), .O(gate241inter9));
  nand2 gate739(.a(s_27), .b(gate241inter3), .O(gate241inter10));
  nor2  gate740(.a(gate241inter10), .b(gate241inter9), .O(gate241inter11));
  nor2  gate741(.a(gate241inter11), .b(gate241inter6), .O(gate241inter12));
  nand2 gate742(.a(gate241inter12), .b(gate241inter1), .O(G754));

  xor2  gate1821(.a(G730), .b(G718), .O(gate242inter0));
  nand2 gate1822(.a(gate242inter0), .b(s_182), .O(gate242inter1));
  and2  gate1823(.a(G730), .b(G718), .O(gate242inter2));
  inv1  gate1824(.a(s_182), .O(gate242inter3));
  inv1  gate1825(.a(s_183), .O(gate242inter4));
  nand2 gate1826(.a(gate242inter4), .b(gate242inter3), .O(gate242inter5));
  nor2  gate1827(.a(gate242inter5), .b(gate242inter2), .O(gate242inter6));
  inv1  gate1828(.a(G718), .O(gate242inter7));
  inv1  gate1829(.a(G730), .O(gate242inter8));
  nand2 gate1830(.a(gate242inter8), .b(gate242inter7), .O(gate242inter9));
  nand2 gate1831(.a(s_183), .b(gate242inter3), .O(gate242inter10));
  nor2  gate1832(.a(gate242inter10), .b(gate242inter9), .O(gate242inter11));
  nor2  gate1833(.a(gate242inter11), .b(gate242inter6), .O(gate242inter12));
  nand2 gate1834(.a(gate242inter12), .b(gate242inter1), .O(G755));
nand2 gate243( .a(G245), .b(G733), .O(G756) );
nand2 gate244( .a(G721), .b(G733), .O(G757) );
nand2 gate245( .a(G248), .b(G736), .O(G758) );
nand2 gate246( .a(G724), .b(G736), .O(G759) );
nand2 gate247( .a(G251), .b(G739), .O(G760) );
nand2 gate248( .a(G727), .b(G739), .O(G761) );
nand2 gate249( .a(G254), .b(G742), .O(G762) );
nand2 gate250( .a(G706), .b(G742), .O(G763) );
nand2 gate251( .a(G257), .b(G745), .O(G764) );
nand2 gate252( .a(G709), .b(G745), .O(G765) );
nand2 gate253( .a(G260), .b(G748), .O(G766) );

  xor2  gate2255(.a(G748), .b(G712), .O(gate254inter0));
  nand2 gate2256(.a(gate254inter0), .b(s_244), .O(gate254inter1));
  and2  gate2257(.a(G748), .b(G712), .O(gate254inter2));
  inv1  gate2258(.a(s_244), .O(gate254inter3));
  inv1  gate2259(.a(s_245), .O(gate254inter4));
  nand2 gate2260(.a(gate254inter4), .b(gate254inter3), .O(gate254inter5));
  nor2  gate2261(.a(gate254inter5), .b(gate254inter2), .O(gate254inter6));
  inv1  gate2262(.a(G712), .O(gate254inter7));
  inv1  gate2263(.a(G748), .O(gate254inter8));
  nand2 gate2264(.a(gate254inter8), .b(gate254inter7), .O(gate254inter9));
  nand2 gate2265(.a(s_245), .b(gate254inter3), .O(gate254inter10));
  nor2  gate2266(.a(gate254inter10), .b(gate254inter9), .O(gate254inter11));
  nor2  gate2267(.a(gate254inter11), .b(gate254inter6), .O(gate254inter12));
  nand2 gate2268(.a(gate254inter12), .b(gate254inter1), .O(G767));
nand2 gate255( .a(G263), .b(G751), .O(G768) );
nand2 gate256( .a(G715), .b(G751), .O(G769) );
nand2 gate257( .a(G754), .b(G755), .O(G770) );
nand2 gate258( .a(G756), .b(G757), .O(G773) );

  xor2  gate1765(.a(G759), .b(G758), .O(gate259inter0));
  nand2 gate1766(.a(gate259inter0), .b(s_174), .O(gate259inter1));
  and2  gate1767(.a(G759), .b(G758), .O(gate259inter2));
  inv1  gate1768(.a(s_174), .O(gate259inter3));
  inv1  gate1769(.a(s_175), .O(gate259inter4));
  nand2 gate1770(.a(gate259inter4), .b(gate259inter3), .O(gate259inter5));
  nor2  gate1771(.a(gate259inter5), .b(gate259inter2), .O(gate259inter6));
  inv1  gate1772(.a(G758), .O(gate259inter7));
  inv1  gate1773(.a(G759), .O(gate259inter8));
  nand2 gate1774(.a(gate259inter8), .b(gate259inter7), .O(gate259inter9));
  nand2 gate1775(.a(s_175), .b(gate259inter3), .O(gate259inter10));
  nor2  gate1776(.a(gate259inter10), .b(gate259inter9), .O(gate259inter11));
  nor2  gate1777(.a(gate259inter11), .b(gate259inter6), .O(gate259inter12));
  nand2 gate1778(.a(gate259inter12), .b(gate259inter1), .O(G776));

  xor2  gate1485(.a(G761), .b(G760), .O(gate260inter0));
  nand2 gate1486(.a(gate260inter0), .b(s_134), .O(gate260inter1));
  and2  gate1487(.a(G761), .b(G760), .O(gate260inter2));
  inv1  gate1488(.a(s_134), .O(gate260inter3));
  inv1  gate1489(.a(s_135), .O(gate260inter4));
  nand2 gate1490(.a(gate260inter4), .b(gate260inter3), .O(gate260inter5));
  nor2  gate1491(.a(gate260inter5), .b(gate260inter2), .O(gate260inter6));
  inv1  gate1492(.a(G760), .O(gate260inter7));
  inv1  gate1493(.a(G761), .O(gate260inter8));
  nand2 gate1494(.a(gate260inter8), .b(gate260inter7), .O(gate260inter9));
  nand2 gate1495(.a(s_135), .b(gate260inter3), .O(gate260inter10));
  nor2  gate1496(.a(gate260inter10), .b(gate260inter9), .O(gate260inter11));
  nor2  gate1497(.a(gate260inter11), .b(gate260inter6), .O(gate260inter12));
  nand2 gate1498(.a(gate260inter12), .b(gate260inter1), .O(G779));
nand2 gate261( .a(G762), .b(G763), .O(G782) );

  xor2  gate589(.a(G765), .b(G764), .O(gate262inter0));
  nand2 gate590(.a(gate262inter0), .b(s_6), .O(gate262inter1));
  and2  gate591(.a(G765), .b(G764), .O(gate262inter2));
  inv1  gate592(.a(s_6), .O(gate262inter3));
  inv1  gate593(.a(s_7), .O(gate262inter4));
  nand2 gate594(.a(gate262inter4), .b(gate262inter3), .O(gate262inter5));
  nor2  gate595(.a(gate262inter5), .b(gate262inter2), .O(gate262inter6));
  inv1  gate596(.a(G764), .O(gate262inter7));
  inv1  gate597(.a(G765), .O(gate262inter8));
  nand2 gate598(.a(gate262inter8), .b(gate262inter7), .O(gate262inter9));
  nand2 gate599(.a(s_7), .b(gate262inter3), .O(gate262inter10));
  nor2  gate600(.a(gate262inter10), .b(gate262inter9), .O(gate262inter11));
  nor2  gate601(.a(gate262inter11), .b(gate262inter6), .O(gate262inter12));
  nand2 gate602(.a(gate262inter12), .b(gate262inter1), .O(G785));
nand2 gate263( .a(G766), .b(G767), .O(G788) );

  xor2  gate1317(.a(G769), .b(G768), .O(gate264inter0));
  nand2 gate1318(.a(gate264inter0), .b(s_110), .O(gate264inter1));
  and2  gate1319(.a(G769), .b(G768), .O(gate264inter2));
  inv1  gate1320(.a(s_110), .O(gate264inter3));
  inv1  gate1321(.a(s_111), .O(gate264inter4));
  nand2 gate1322(.a(gate264inter4), .b(gate264inter3), .O(gate264inter5));
  nor2  gate1323(.a(gate264inter5), .b(gate264inter2), .O(gate264inter6));
  inv1  gate1324(.a(G768), .O(gate264inter7));
  inv1  gate1325(.a(G769), .O(gate264inter8));
  nand2 gate1326(.a(gate264inter8), .b(gate264inter7), .O(gate264inter9));
  nand2 gate1327(.a(s_111), .b(gate264inter3), .O(gate264inter10));
  nor2  gate1328(.a(gate264inter10), .b(gate264inter9), .O(gate264inter11));
  nor2  gate1329(.a(gate264inter11), .b(gate264inter6), .O(gate264inter12));
  nand2 gate1330(.a(gate264inter12), .b(gate264inter1), .O(G791));
nand2 gate265( .a(G642), .b(G770), .O(G794) );

  xor2  gate1947(.a(G773), .b(G645), .O(gate266inter0));
  nand2 gate1948(.a(gate266inter0), .b(s_200), .O(gate266inter1));
  and2  gate1949(.a(G773), .b(G645), .O(gate266inter2));
  inv1  gate1950(.a(s_200), .O(gate266inter3));
  inv1  gate1951(.a(s_201), .O(gate266inter4));
  nand2 gate1952(.a(gate266inter4), .b(gate266inter3), .O(gate266inter5));
  nor2  gate1953(.a(gate266inter5), .b(gate266inter2), .O(gate266inter6));
  inv1  gate1954(.a(G645), .O(gate266inter7));
  inv1  gate1955(.a(G773), .O(gate266inter8));
  nand2 gate1956(.a(gate266inter8), .b(gate266inter7), .O(gate266inter9));
  nand2 gate1957(.a(s_201), .b(gate266inter3), .O(gate266inter10));
  nor2  gate1958(.a(gate266inter10), .b(gate266inter9), .O(gate266inter11));
  nor2  gate1959(.a(gate266inter11), .b(gate266inter6), .O(gate266inter12));
  nand2 gate1960(.a(gate266inter12), .b(gate266inter1), .O(G797));
nand2 gate267( .a(G648), .b(G776), .O(G800) );
nand2 gate268( .a(G651), .b(G779), .O(G803) );
nand2 gate269( .a(G654), .b(G782), .O(G806) );
nand2 gate270( .a(G657), .b(G785), .O(G809) );
nand2 gate271( .a(G660), .b(G788), .O(G812) );

  xor2  gate1219(.a(G791), .b(G663), .O(gate272inter0));
  nand2 gate1220(.a(gate272inter0), .b(s_96), .O(gate272inter1));
  and2  gate1221(.a(G791), .b(G663), .O(gate272inter2));
  inv1  gate1222(.a(s_96), .O(gate272inter3));
  inv1  gate1223(.a(s_97), .O(gate272inter4));
  nand2 gate1224(.a(gate272inter4), .b(gate272inter3), .O(gate272inter5));
  nor2  gate1225(.a(gate272inter5), .b(gate272inter2), .O(gate272inter6));
  inv1  gate1226(.a(G663), .O(gate272inter7));
  inv1  gate1227(.a(G791), .O(gate272inter8));
  nand2 gate1228(.a(gate272inter8), .b(gate272inter7), .O(gate272inter9));
  nand2 gate1229(.a(s_97), .b(gate272inter3), .O(gate272inter10));
  nor2  gate1230(.a(gate272inter10), .b(gate272inter9), .O(gate272inter11));
  nor2  gate1231(.a(gate272inter11), .b(gate272inter6), .O(gate272inter12));
  nand2 gate1232(.a(gate272inter12), .b(gate272inter1), .O(G815));
nand2 gate273( .a(G642), .b(G794), .O(G818) );

  xor2  gate1919(.a(G794), .b(G770), .O(gate274inter0));
  nand2 gate1920(.a(gate274inter0), .b(s_196), .O(gate274inter1));
  and2  gate1921(.a(G794), .b(G770), .O(gate274inter2));
  inv1  gate1922(.a(s_196), .O(gate274inter3));
  inv1  gate1923(.a(s_197), .O(gate274inter4));
  nand2 gate1924(.a(gate274inter4), .b(gate274inter3), .O(gate274inter5));
  nor2  gate1925(.a(gate274inter5), .b(gate274inter2), .O(gate274inter6));
  inv1  gate1926(.a(G770), .O(gate274inter7));
  inv1  gate1927(.a(G794), .O(gate274inter8));
  nand2 gate1928(.a(gate274inter8), .b(gate274inter7), .O(gate274inter9));
  nand2 gate1929(.a(s_197), .b(gate274inter3), .O(gate274inter10));
  nor2  gate1930(.a(gate274inter10), .b(gate274inter9), .O(gate274inter11));
  nor2  gate1931(.a(gate274inter11), .b(gate274inter6), .O(gate274inter12));
  nand2 gate1932(.a(gate274inter12), .b(gate274inter1), .O(G819));
nand2 gate275( .a(G645), .b(G797), .O(G820) );

  xor2  gate1443(.a(G797), .b(G773), .O(gate276inter0));
  nand2 gate1444(.a(gate276inter0), .b(s_128), .O(gate276inter1));
  and2  gate1445(.a(G797), .b(G773), .O(gate276inter2));
  inv1  gate1446(.a(s_128), .O(gate276inter3));
  inv1  gate1447(.a(s_129), .O(gate276inter4));
  nand2 gate1448(.a(gate276inter4), .b(gate276inter3), .O(gate276inter5));
  nor2  gate1449(.a(gate276inter5), .b(gate276inter2), .O(gate276inter6));
  inv1  gate1450(.a(G773), .O(gate276inter7));
  inv1  gate1451(.a(G797), .O(gate276inter8));
  nand2 gate1452(.a(gate276inter8), .b(gate276inter7), .O(gate276inter9));
  nand2 gate1453(.a(s_129), .b(gate276inter3), .O(gate276inter10));
  nor2  gate1454(.a(gate276inter10), .b(gate276inter9), .O(gate276inter11));
  nor2  gate1455(.a(gate276inter11), .b(gate276inter6), .O(gate276inter12));
  nand2 gate1456(.a(gate276inter12), .b(gate276inter1), .O(G821));
nand2 gate277( .a(G648), .b(G800), .O(G822) );
nand2 gate278( .a(G776), .b(G800), .O(G823) );
nand2 gate279( .a(G651), .b(G803), .O(G824) );
nand2 gate280( .a(G779), .b(G803), .O(G825) );

  xor2  gate981(.a(G806), .b(G654), .O(gate281inter0));
  nand2 gate982(.a(gate281inter0), .b(s_62), .O(gate281inter1));
  and2  gate983(.a(G806), .b(G654), .O(gate281inter2));
  inv1  gate984(.a(s_62), .O(gate281inter3));
  inv1  gate985(.a(s_63), .O(gate281inter4));
  nand2 gate986(.a(gate281inter4), .b(gate281inter3), .O(gate281inter5));
  nor2  gate987(.a(gate281inter5), .b(gate281inter2), .O(gate281inter6));
  inv1  gate988(.a(G654), .O(gate281inter7));
  inv1  gate989(.a(G806), .O(gate281inter8));
  nand2 gate990(.a(gate281inter8), .b(gate281inter7), .O(gate281inter9));
  nand2 gate991(.a(s_63), .b(gate281inter3), .O(gate281inter10));
  nor2  gate992(.a(gate281inter10), .b(gate281inter9), .O(gate281inter11));
  nor2  gate993(.a(gate281inter11), .b(gate281inter6), .O(gate281inter12));
  nand2 gate994(.a(gate281inter12), .b(gate281inter1), .O(G826));
nand2 gate282( .a(G782), .b(G806), .O(G827) );
nand2 gate283( .a(G657), .b(G809), .O(G828) );
nand2 gate284( .a(G785), .b(G809), .O(G829) );
nand2 gate285( .a(G660), .b(G812), .O(G830) );
nand2 gate286( .a(G788), .b(G812), .O(G831) );
nand2 gate287( .a(G663), .b(G815), .O(G832) );
nand2 gate288( .a(G791), .b(G815), .O(G833) );

  xor2  gate1233(.a(G819), .b(G818), .O(gate289inter0));
  nand2 gate1234(.a(gate289inter0), .b(s_98), .O(gate289inter1));
  and2  gate1235(.a(G819), .b(G818), .O(gate289inter2));
  inv1  gate1236(.a(s_98), .O(gate289inter3));
  inv1  gate1237(.a(s_99), .O(gate289inter4));
  nand2 gate1238(.a(gate289inter4), .b(gate289inter3), .O(gate289inter5));
  nor2  gate1239(.a(gate289inter5), .b(gate289inter2), .O(gate289inter6));
  inv1  gate1240(.a(G818), .O(gate289inter7));
  inv1  gate1241(.a(G819), .O(gate289inter8));
  nand2 gate1242(.a(gate289inter8), .b(gate289inter7), .O(gate289inter9));
  nand2 gate1243(.a(s_99), .b(gate289inter3), .O(gate289inter10));
  nor2  gate1244(.a(gate289inter10), .b(gate289inter9), .O(gate289inter11));
  nor2  gate1245(.a(gate289inter11), .b(gate289inter6), .O(gate289inter12));
  nand2 gate1246(.a(gate289inter12), .b(gate289inter1), .O(G834));
nand2 gate290( .a(G820), .b(G821), .O(G847) );
nand2 gate291( .a(G822), .b(G823), .O(G860) );

  xor2  gate1863(.a(G825), .b(G824), .O(gate292inter0));
  nand2 gate1864(.a(gate292inter0), .b(s_188), .O(gate292inter1));
  and2  gate1865(.a(G825), .b(G824), .O(gate292inter2));
  inv1  gate1866(.a(s_188), .O(gate292inter3));
  inv1  gate1867(.a(s_189), .O(gate292inter4));
  nand2 gate1868(.a(gate292inter4), .b(gate292inter3), .O(gate292inter5));
  nor2  gate1869(.a(gate292inter5), .b(gate292inter2), .O(gate292inter6));
  inv1  gate1870(.a(G824), .O(gate292inter7));
  inv1  gate1871(.a(G825), .O(gate292inter8));
  nand2 gate1872(.a(gate292inter8), .b(gate292inter7), .O(gate292inter9));
  nand2 gate1873(.a(s_189), .b(gate292inter3), .O(gate292inter10));
  nor2  gate1874(.a(gate292inter10), .b(gate292inter9), .O(gate292inter11));
  nor2  gate1875(.a(gate292inter11), .b(gate292inter6), .O(gate292inter12));
  nand2 gate1876(.a(gate292inter12), .b(gate292inter1), .O(G873));

  xor2  gate1835(.a(G829), .b(G828), .O(gate293inter0));
  nand2 gate1836(.a(gate293inter0), .b(s_184), .O(gate293inter1));
  and2  gate1837(.a(G829), .b(G828), .O(gate293inter2));
  inv1  gate1838(.a(s_184), .O(gate293inter3));
  inv1  gate1839(.a(s_185), .O(gate293inter4));
  nand2 gate1840(.a(gate293inter4), .b(gate293inter3), .O(gate293inter5));
  nor2  gate1841(.a(gate293inter5), .b(gate293inter2), .O(gate293inter6));
  inv1  gate1842(.a(G828), .O(gate293inter7));
  inv1  gate1843(.a(G829), .O(gate293inter8));
  nand2 gate1844(.a(gate293inter8), .b(gate293inter7), .O(gate293inter9));
  nand2 gate1845(.a(s_185), .b(gate293inter3), .O(gate293inter10));
  nor2  gate1846(.a(gate293inter10), .b(gate293inter9), .O(gate293inter11));
  nor2  gate1847(.a(gate293inter11), .b(gate293inter6), .O(gate293inter12));
  nand2 gate1848(.a(gate293inter12), .b(gate293inter1), .O(G886));
nand2 gate294( .a(G832), .b(G833), .O(G899) );
nand2 gate295( .a(G830), .b(G831), .O(G912) );

  xor2  gate1975(.a(G827), .b(G826), .O(gate296inter0));
  nand2 gate1976(.a(gate296inter0), .b(s_204), .O(gate296inter1));
  and2  gate1977(.a(G827), .b(G826), .O(gate296inter2));
  inv1  gate1978(.a(s_204), .O(gate296inter3));
  inv1  gate1979(.a(s_205), .O(gate296inter4));
  nand2 gate1980(.a(gate296inter4), .b(gate296inter3), .O(gate296inter5));
  nor2  gate1981(.a(gate296inter5), .b(gate296inter2), .O(gate296inter6));
  inv1  gate1982(.a(G826), .O(gate296inter7));
  inv1  gate1983(.a(G827), .O(gate296inter8));
  nand2 gate1984(.a(gate296inter8), .b(gate296inter7), .O(gate296inter9));
  nand2 gate1985(.a(s_205), .b(gate296inter3), .O(gate296inter10));
  nor2  gate1986(.a(gate296inter10), .b(gate296inter9), .O(gate296inter11));
  nor2  gate1987(.a(gate296inter11), .b(gate296inter6), .O(gate296inter12));
  nand2 gate1988(.a(gate296inter12), .b(gate296inter1), .O(G925));
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );
nand2 gate387( .a(G1), .b(G1036), .O(G1132) );
nand2 gate388( .a(G2), .b(G1039), .O(G1135) );
nand2 gate389( .a(G3), .b(G1042), .O(G1138) );
nand2 gate390( .a(G4), .b(G1045), .O(G1141) );
nand2 gate391( .a(G5), .b(G1048), .O(G1144) );
nand2 gate392( .a(G6), .b(G1051), .O(G1147) );

  xor2  gate1583(.a(G1054), .b(G7), .O(gate393inter0));
  nand2 gate1584(.a(gate393inter0), .b(s_148), .O(gate393inter1));
  and2  gate1585(.a(G1054), .b(G7), .O(gate393inter2));
  inv1  gate1586(.a(s_148), .O(gate393inter3));
  inv1  gate1587(.a(s_149), .O(gate393inter4));
  nand2 gate1588(.a(gate393inter4), .b(gate393inter3), .O(gate393inter5));
  nor2  gate1589(.a(gate393inter5), .b(gate393inter2), .O(gate393inter6));
  inv1  gate1590(.a(G7), .O(gate393inter7));
  inv1  gate1591(.a(G1054), .O(gate393inter8));
  nand2 gate1592(.a(gate393inter8), .b(gate393inter7), .O(gate393inter9));
  nand2 gate1593(.a(s_149), .b(gate393inter3), .O(gate393inter10));
  nor2  gate1594(.a(gate393inter10), .b(gate393inter9), .O(gate393inter11));
  nor2  gate1595(.a(gate393inter11), .b(gate393inter6), .O(gate393inter12));
  nand2 gate1596(.a(gate393inter12), .b(gate393inter1), .O(G1150));

  xor2  gate1807(.a(G1057), .b(G8), .O(gate394inter0));
  nand2 gate1808(.a(gate394inter0), .b(s_180), .O(gate394inter1));
  and2  gate1809(.a(G1057), .b(G8), .O(gate394inter2));
  inv1  gate1810(.a(s_180), .O(gate394inter3));
  inv1  gate1811(.a(s_181), .O(gate394inter4));
  nand2 gate1812(.a(gate394inter4), .b(gate394inter3), .O(gate394inter5));
  nor2  gate1813(.a(gate394inter5), .b(gate394inter2), .O(gate394inter6));
  inv1  gate1814(.a(G8), .O(gate394inter7));
  inv1  gate1815(.a(G1057), .O(gate394inter8));
  nand2 gate1816(.a(gate394inter8), .b(gate394inter7), .O(gate394inter9));
  nand2 gate1817(.a(s_181), .b(gate394inter3), .O(gate394inter10));
  nor2  gate1818(.a(gate394inter10), .b(gate394inter9), .O(gate394inter11));
  nor2  gate1819(.a(gate394inter11), .b(gate394inter6), .O(gate394inter12));
  nand2 gate1820(.a(gate394inter12), .b(gate394inter1), .O(G1153));

  xor2  gate1023(.a(G1060), .b(G9), .O(gate395inter0));
  nand2 gate1024(.a(gate395inter0), .b(s_68), .O(gate395inter1));
  and2  gate1025(.a(G1060), .b(G9), .O(gate395inter2));
  inv1  gate1026(.a(s_68), .O(gate395inter3));
  inv1  gate1027(.a(s_69), .O(gate395inter4));
  nand2 gate1028(.a(gate395inter4), .b(gate395inter3), .O(gate395inter5));
  nor2  gate1029(.a(gate395inter5), .b(gate395inter2), .O(gate395inter6));
  inv1  gate1030(.a(G9), .O(gate395inter7));
  inv1  gate1031(.a(G1060), .O(gate395inter8));
  nand2 gate1032(.a(gate395inter8), .b(gate395inter7), .O(gate395inter9));
  nand2 gate1033(.a(s_69), .b(gate395inter3), .O(gate395inter10));
  nor2  gate1034(.a(gate395inter10), .b(gate395inter9), .O(gate395inter11));
  nor2  gate1035(.a(gate395inter11), .b(gate395inter6), .O(gate395inter12));
  nand2 gate1036(.a(gate395inter12), .b(gate395inter1), .O(G1156));
nand2 gate396( .a(G10), .b(G1063), .O(G1159) );

  xor2  gate1933(.a(G1066), .b(G11), .O(gate397inter0));
  nand2 gate1934(.a(gate397inter0), .b(s_198), .O(gate397inter1));
  and2  gate1935(.a(G1066), .b(G11), .O(gate397inter2));
  inv1  gate1936(.a(s_198), .O(gate397inter3));
  inv1  gate1937(.a(s_199), .O(gate397inter4));
  nand2 gate1938(.a(gate397inter4), .b(gate397inter3), .O(gate397inter5));
  nor2  gate1939(.a(gate397inter5), .b(gate397inter2), .O(gate397inter6));
  inv1  gate1940(.a(G11), .O(gate397inter7));
  inv1  gate1941(.a(G1066), .O(gate397inter8));
  nand2 gate1942(.a(gate397inter8), .b(gate397inter7), .O(gate397inter9));
  nand2 gate1943(.a(s_199), .b(gate397inter3), .O(gate397inter10));
  nor2  gate1944(.a(gate397inter10), .b(gate397inter9), .O(gate397inter11));
  nor2  gate1945(.a(gate397inter11), .b(gate397inter6), .O(gate397inter12));
  nand2 gate1946(.a(gate397inter12), .b(gate397inter1), .O(G1162));

  xor2  gate1457(.a(G1069), .b(G12), .O(gate398inter0));
  nand2 gate1458(.a(gate398inter0), .b(s_130), .O(gate398inter1));
  and2  gate1459(.a(G1069), .b(G12), .O(gate398inter2));
  inv1  gate1460(.a(s_130), .O(gate398inter3));
  inv1  gate1461(.a(s_131), .O(gate398inter4));
  nand2 gate1462(.a(gate398inter4), .b(gate398inter3), .O(gate398inter5));
  nor2  gate1463(.a(gate398inter5), .b(gate398inter2), .O(gate398inter6));
  inv1  gate1464(.a(G12), .O(gate398inter7));
  inv1  gate1465(.a(G1069), .O(gate398inter8));
  nand2 gate1466(.a(gate398inter8), .b(gate398inter7), .O(gate398inter9));
  nand2 gate1467(.a(s_131), .b(gate398inter3), .O(gate398inter10));
  nor2  gate1468(.a(gate398inter10), .b(gate398inter9), .O(gate398inter11));
  nor2  gate1469(.a(gate398inter11), .b(gate398inter6), .O(gate398inter12));
  nand2 gate1470(.a(gate398inter12), .b(gate398inter1), .O(G1165));

  xor2  gate2045(.a(G1072), .b(G13), .O(gate399inter0));
  nand2 gate2046(.a(gate399inter0), .b(s_214), .O(gate399inter1));
  and2  gate2047(.a(G1072), .b(G13), .O(gate399inter2));
  inv1  gate2048(.a(s_214), .O(gate399inter3));
  inv1  gate2049(.a(s_215), .O(gate399inter4));
  nand2 gate2050(.a(gate399inter4), .b(gate399inter3), .O(gate399inter5));
  nor2  gate2051(.a(gate399inter5), .b(gate399inter2), .O(gate399inter6));
  inv1  gate2052(.a(G13), .O(gate399inter7));
  inv1  gate2053(.a(G1072), .O(gate399inter8));
  nand2 gate2054(.a(gate399inter8), .b(gate399inter7), .O(gate399inter9));
  nand2 gate2055(.a(s_215), .b(gate399inter3), .O(gate399inter10));
  nor2  gate2056(.a(gate399inter10), .b(gate399inter9), .O(gate399inter11));
  nor2  gate2057(.a(gate399inter11), .b(gate399inter6), .O(gate399inter12));
  nand2 gate2058(.a(gate399inter12), .b(gate399inter1), .O(G1168));
nand2 gate400( .a(G14), .b(G1075), .O(G1171) );

  xor2  gate1303(.a(G1078), .b(G15), .O(gate401inter0));
  nand2 gate1304(.a(gate401inter0), .b(s_108), .O(gate401inter1));
  and2  gate1305(.a(G1078), .b(G15), .O(gate401inter2));
  inv1  gate1306(.a(s_108), .O(gate401inter3));
  inv1  gate1307(.a(s_109), .O(gate401inter4));
  nand2 gate1308(.a(gate401inter4), .b(gate401inter3), .O(gate401inter5));
  nor2  gate1309(.a(gate401inter5), .b(gate401inter2), .O(gate401inter6));
  inv1  gate1310(.a(G15), .O(gate401inter7));
  inv1  gate1311(.a(G1078), .O(gate401inter8));
  nand2 gate1312(.a(gate401inter8), .b(gate401inter7), .O(gate401inter9));
  nand2 gate1313(.a(s_109), .b(gate401inter3), .O(gate401inter10));
  nor2  gate1314(.a(gate401inter10), .b(gate401inter9), .O(gate401inter11));
  nor2  gate1315(.a(gate401inter11), .b(gate401inter6), .O(gate401inter12));
  nand2 gate1316(.a(gate401inter12), .b(gate401inter1), .O(G1174));
nand2 gate402( .a(G16), .b(G1081), .O(G1177) );
nand2 gate403( .a(G17), .b(G1084), .O(G1180) );
nand2 gate404( .a(G18), .b(G1087), .O(G1183) );
nand2 gate405( .a(G19), .b(G1090), .O(G1186) );

  xor2  gate2311(.a(G1093), .b(G20), .O(gate406inter0));
  nand2 gate2312(.a(gate406inter0), .b(s_252), .O(gate406inter1));
  and2  gate2313(.a(G1093), .b(G20), .O(gate406inter2));
  inv1  gate2314(.a(s_252), .O(gate406inter3));
  inv1  gate2315(.a(s_253), .O(gate406inter4));
  nand2 gate2316(.a(gate406inter4), .b(gate406inter3), .O(gate406inter5));
  nor2  gate2317(.a(gate406inter5), .b(gate406inter2), .O(gate406inter6));
  inv1  gate2318(.a(G20), .O(gate406inter7));
  inv1  gate2319(.a(G1093), .O(gate406inter8));
  nand2 gate2320(.a(gate406inter8), .b(gate406inter7), .O(gate406inter9));
  nand2 gate2321(.a(s_253), .b(gate406inter3), .O(gate406inter10));
  nor2  gate2322(.a(gate406inter10), .b(gate406inter9), .O(gate406inter11));
  nor2  gate2323(.a(gate406inter11), .b(gate406inter6), .O(gate406inter12));
  nand2 gate2324(.a(gate406inter12), .b(gate406inter1), .O(G1189));

  xor2  gate841(.a(G1096), .b(G21), .O(gate407inter0));
  nand2 gate842(.a(gate407inter0), .b(s_42), .O(gate407inter1));
  and2  gate843(.a(G1096), .b(G21), .O(gate407inter2));
  inv1  gate844(.a(s_42), .O(gate407inter3));
  inv1  gate845(.a(s_43), .O(gate407inter4));
  nand2 gate846(.a(gate407inter4), .b(gate407inter3), .O(gate407inter5));
  nor2  gate847(.a(gate407inter5), .b(gate407inter2), .O(gate407inter6));
  inv1  gate848(.a(G21), .O(gate407inter7));
  inv1  gate849(.a(G1096), .O(gate407inter8));
  nand2 gate850(.a(gate407inter8), .b(gate407inter7), .O(gate407inter9));
  nand2 gate851(.a(s_43), .b(gate407inter3), .O(gate407inter10));
  nor2  gate852(.a(gate407inter10), .b(gate407inter9), .O(gate407inter11));
  nor2  gate853(.a(gate407inter11), .b(gate407inter6), .O(gate407inter12));
  nand2 gate854(.a(gate407inter12), .b(gate407inter1), .O(G1192));
nand2 gate408( .a(G22), .b(G1099), .O(G1195) );
nand2 gate409( .a(G23), .b(G1102), .O(G1198) );

  xor2  gate1723(.a(G1105), .b(G24), .O(gate410inter0));
  nand2 gate1724(.a(gate410inter0), .b(s_168), .O(gate410inter1));
  and2  gate1725(.a(G1105), .b(G24), .O(gate410inter2));
  inv1  gate1726(.a(s_168), .O(gate410inter3));
  inv1  gate1727(.a(s_169), .O(gate410inter4));
  nand2 gate1728(.a(gate410inter4), .b(gate410inter3), .O(gate410inter5));
  nor2  gate1729(.a(gate410inter5), .b(gate410inter2), .O(gate410inter6));
  inv1  gate1730(.a(G24), .O(gate410inter7));
  inv1  gate1731(.a(G1105), .O(gate410inter8));
  nand2 gate1732(.a(gate410inter8), .b(gate410inter7), .O(gate410inter9));
  nand2 gate1733(.a(s_169), .b(gate410inter3), .O(gate410inter10));
  nor2  gate1734(.a(gate410inter10), .b(gate410inter9), .O(gate410inter11));
  nor2  gate1735(.a(gate410inter11), .b(gate410inter6), .O(gate410inter12));
  nand2 gate1736(.a(gate410inter12), .b(gate410inter1), .O(G1201));
nand2 gate411( .a(G25), .b(G1108), .O(G1204) );
nand2 gate412( .a(G26), .b(G1111), .O(G1207) );
nand2 gate413( .a(G27), .b(G1114), .O(G1210) );
nand2 gate414( .a(G28), .b(G1117), .O(G1213) );

  xor2  gate2269(.a(G1120), .b(G29), .O(gate415inter0));
  nand2 gate2270(.a(gate415inter0), .b(s_246), .O(gate415inter1));
  and2  gate2271(.a(G1120), .b(G29), .O(gate415inter2));
  inv1  gate2272(.a(s_246), .O(gate415inter3));
  inv1  gate2273(.a(s_247), .O(gate415inter4));
  nand2 gate2274(.a(gate415inter4), .b(gate415inter3), .O(gate415inter5));
  nor2  gate2275(.a(gate415inter5), .b(gate415inter2), .O(gate415inter6));
  inv1  gate2276(.a(G29), .O(gate415inter7));
  inv1  gate2277(.a(G1120), .O(gate415inter8));
  nand2 gate2278(.a(gate415inter8), .b(gate415inter7), .O(gate415inter9));
  nand2 gate2279(.a(s_247), .b(gate415inter3), .O(gate415inter10));
  nor2  gate2280(.a(gate415inter10), .b(gate415inter9), .O(gate415inter11));
  nor2  gate2281(.a(gate415inter11), .b(gate415inter6), .O(gate415inter12));
  nand2 gate2282(.a(gate415inter12), .b(gate415inter1), .O(G1216));
nand2 gate416( .a(G30), .b(G1123), .O(G1219) );

  xor2  gate953(.a(G1126), .b(G31), .O(gate417inter0));
  nand2 gate954(.a(gate417inter0), .b(s_58), .O(gate417inter1));
  and2  gate955(.a(G1126), .b(G31), .O(gate417inter2));
  inv1  gate956(.a(s_58), .O(gate417inter3));
  inv1  gate957(.a(s_59), .O(gate417inter4));
  nand2 gate958(.a(gate417inter4), .b(gate417inter3), .O(gate417inter5));
  nor2  gate959(.a(gate417inter5), .b(gate417inter2), .O(gate417inter6));
  inv1  gate960(.a(G31), .O(gate417inter7));
  inv1  gate961(.a(G1126), .O(gate417inter8));
  nand2 gate962(.a(gate417inter8), .b(gate417inter7), .O(gate417inter9));
  nand2 gate963(.a(s_59), .b(gate417inter3), .O(gate417inter10));
  nor2  gate964(.a(gate417inter10), .b(gate417inter9), .O(gate417inter11));
  nor2  gate965(.a(gate417inter11), .b(gate417inter6), .O(gate417inter12));
  nand2 gate966(.a(gate417inter12), .b(gate417inter1), .O(G1222));
nand2 gate418( .a(G32), .b(G1129), .O(G1225) );
nand2 gate419( .a(G1), .b(G1132), .O(G1228) );
nand2 gate420( .a(G1036), .b(G1132), .O(G1229) );
nand2 gate421( .a(G2), .b(G1135), .O(G1230) );
nand2 gate422( .a(G1039), .b(G1135), .O(G1231) );
nand2 gate423( .a(G3), .b(G1138), .O(G1232) );
nand2 gate424( .a(G1042), .b(G1138), .O(G1233) );
nand2 gate425( .a(G4), .b(G1141), .O(G1234) );

  xor2  gate827(.a(G1141), .b(G1045), .O(gate426inter0));
  nand2 gate828(.a(gate426inter0), .b(s_40), .O(gate426inter1));
  and2  gate829(.a(G1141), .b(G1045), .O(gate426inter2));
  inv1  gate830(.a(s_40), .O(gate426inter3));
  inv1  gate831(.a(s_41), .O(gate426inter4));
  nand2 gate832(.a(gate426inter4), .b(gate426inter3), .O(gate426inter5));
  nor2  gate833(.a(gate426inter5), .b(gate426inter2), .O(gate426inter6));
  inv1  gate834(.a(G1045), .O(gate426inter7));
  inv1  gate835(.a(G1141), .O(gate426inter8));
  nand2 gate836(.a(gate426inter8), .b(gate426inter7), .O(gate426inter9));
  nand2 gate837(.a(s_41), .b(gate426inter3), .O(gate426inter10));
  nor2  gate838(.a(gate426inter10), .b(gate426inter9), .O(gate426inter11));
  nor2  gate839(.a(gate426inter11), .b(gate426inter6), .O(gate426inter12));
  nand2 gate840(.a(gate426inter12), .b(gate426inter1), .O(G1235));
nand2 gate427( .a(G5), .b(G1144), .O(G1236) );

  xor2  gate1681(.a(G1144), .b(G1048), .O(gate428inter0));
  nand2 gate1682(.a(gate428inter0), .b(s_162), .O(gate428inter1));
  and2  gate1683(.a(G1144), .b(G1048), .O(gate428inter2));
  inv1  gate1684(.a(s_162), .O(gate428inter3));
  inv1  gate1685(.a(s_163), .O(gate428inter4));
  nand2 gate1686(.a(gate428inter4), .b(gate428inter3), .O(gate428inter5));
  nor2  gate1687(.a(gate428inter5), .b(gate428inter2), .O(gate428inter6));
  inv1  gate1688(.a(G1048), .O(gate428inter7));
  inv1  gate1689(.a(G1144), .O(gate428inter8));
  nand2 gate1690(.a(gate428inter8), .b(gate428inter7), .O(gate428inter9));
  nand2 gate1691(.a(s_163), .b(gate428inter3), .O(gate428inter10));
  nor2  gate1692(.a(gate428inter10), .b(gate428inter9), .O(gate428inter11));
  nor2  gate1693(.a(gate428inter11), .b(gate428inter6), .O(gate428inter12));
  nand2 gate1694(.a(gate428inter12), .b(gate428inter1), .O(G1237));

  xor2  gate2003(.a(G1147), .b(G6), .O(gate429inter0));
  nand2 gate2004(.a(gate429inter0), .b(s_208), .O(gate429inter1));
  and2  gate2005(.a(G1147), .b(G6), .O(gate429inter2));
  inv1  gate2006(.a(s_208), .O(gate429inter3));
  inv1  gate2007(.a(s_209), .O(gate429inter4));
  nand2 gate2008(.a(gate429inter4), .b(gate429inter3), .O(gate429inter5));
  nor2  gate2009(.a(gate429inter5), .b(gate429inter2), .O(gate429inter6));
  inv1  gate2010(.a(G6), .O(gate429inter7));
  inv1  gate2011(.a(G1147), .O(gate429inter8));
  nand2 gate2012(.a(gate429inter8), .b(gate429inter7), .O(gate429inter9));
  nand2 gate2013(.a(s_209), .b(gate429inter3), .O(gate429inter10));
  nor2  gate2014(.a(gate429inter10), .b(gate429inter9), .O(gate429inter11));
  nor2  gate2015(.a(gate429inter11), .b(gate429inter6), .O(gate429inter12));
  nand2 gate2016(.a(gate429inter12), .b(gate429inter1), .O(G1238));
nand2 gate430( .a(G1051), .b(G1147), .O(G1239) );

  xor2  gate1709(.a(G1150), .b(G7), .O(gate431inter0));
  nand2 gate1710(.a(gate431inter0), .b(s_166), .O(gate431inter1));
  and2  gate1711(.a(G1150), .b(G7), .O(gate431inter2));
  inv1  gate1712(.a(s_166), .O(gate431inter3));
  inv1  gate1713(.a(s_167), .O(gate431inter4));
  nand2 gate1714(.a(gate431inter4), .b(gate431inter3), .O(gate431inter5));
  nor2  gate1715(.a(gate431inter5), .b(gate431inter2), .O(gate431inter6));
  inv1  gate1716(.a(G7), .O(gate431inter7));
  inv1  gate1717(.a(G1150), .O(gate431inter8));
  nand2 gate1718(.a(gate431inter8), .b(gate431inter7), .O(gate431inter9));
  nand2 gate1719(.a(s_167), .b(gate431inter3), .O(gate431inter10));
  nor2  gate1720(.a(gate431inter10), .b(gate431inter9), .O(gate431inter11));
  nor2  gate1721(.a(gate431inter11), .b(gate431inter6), .O(gate431inter12));
  nand2 gate1722(.a(gate431inter12), .b(gate431inter1), .O(G1240));

  xor2  gate631(.a(G1150), .b(G1054), .O(gate432inter0));
  nand2 gate632(.a(gate432inter0), .b(s_12), .O(gate432inter1));
  and2  gate633(.a(G1150), .b(G1054), .O(gate432inter2));
  inv1  gate634(.a(s_12), .O(gate432inter3));
  inv1  gate635(.a(s_13), .O(gate432inter4));
  nand2 gate636(.a(gate432inter4), .b(gate432inter3), .O(gate432inter5));
  nor2  gate637(.a(gate432inter5), .b(gate432inter2), .O(gate432inter6));
  inv1  gate638(.a(G1054), .O(gate432inter7));
  inv1  gate639(.a(G1150), .O(gate432inter8));
  nand2 gate640(.a(gate432inter8), .b(gate432inter7), .O(gate432inter9));
  nand2 gate641(.a(s_13), .b(gate432inter3), .O(gate432inter10));
  nor2  gate642(.a(gate432inter10), .b(gate432inter9), .O(gate432inter11));
  nor2  gate643(.a(gate432inter11), .b(gate432inter6), .O(gate432inter12));
  nand2 gate644(.a(gate432inter12), .b(gate432inter1), .O(G1241));
nand2 gate433( .a(G8), .b(G1153), .O(G1242) );
nand2 gate434( .a(G1057), .b(G1153), .O(G1243) );
nand2 gate435( .a(G9), .b(G1156), .O(G1244) );
nand2 gate436( .a(G1060), .b(G1156), .O(G1245) );
nand2 gate437( .a(G10), .b(G1159), .O(G1246) );
nand2 gate438( .a(G1063), .b(G1159), .O(G1247) );
nand2 gate439( .a(G11), .b(G1162), .O(G1248) );
nand2 gate440( .a(G1066), .b(G1162), .O(G1249) );
nand2 gate441( .a(G12), .b(G1165), .O(G1250) );
nand2 gate442( .a(G1069), .b(G1165), .O(G1251) );
nand2 gate443( .a(G13), .b(G1168), .O(G1252) );
nand2 gate444( .a(G1072), .b(G1168), .O(G1253) );

  xor2  gate911(.a(G1171), .b(G14), .O(gate445inter0));
  nand2 gate912(.a(gate445inter0), .b(s_52), .O(gate445inter1));
  and2  gate913(.a(G1171), .b(G14), .O(gate445inter2));
  inv1  gate914(.a(s_52), .O(gate445inter3));
  inv1  gate915(.a(s_53), .O(gate445inter4));
  nand2 gate916(.a(gate445inter4), .b(gate445inter3), .O(gate445inter5));
  nor2  gate917(.a(gate445inter5), .b(gate445inter2), .O(gate445inter6));
  inv1  gate918(.a(G14), .O(gate445inter7));
  inv1  gate919(.a(G1171), .O(gate445inter8));
  nand2 gate920(.a(gate445inter8), .b(gate445inter7), .O(gate445inter9));
  nand2 gate921(.a(s_53), .b(gate445inter3), .O(gate445inter10));
  nor2  gate922(.a(gate445inter10), .b(gate445inter9), .O(gate445inter11));
  nor2  gate923(.a(gate445inter11), .b(gate445inter6), .O(gate445inter12));
  nand2 gate924(.a(gate445inter12), .b(gate445inter1), .O(G1254));

  xor2  gate869(.a(G1171), .b(G1075), .O(gate446inter0));
  nand2 gate870(.a(gate446inter0), .b(s_46), .O(gate446inter1));
  and2  gate871(.a(G1171), .b(G1075), .O(gate446inter2));
  inv1  gate872(.a(s_46), .O(gate446inter3));
  inv1  gate873(.a(s_47), .O(gate446inter4));
  nand2 gate874(.a(gate446inter4), .b(gate446inter3), .O(gate446inter5));
  nor2  gate875(.a(gate446inter5), .b(gate446inter2), .O(gate446inter6));
  inv1  gate876(.a(G1075), .O(gate446inter7));
  inv1  gate877(.a(G1171), .O(gate446inter8));
  nand2 gate878(.a(gate446inter8), .b(gate446inter7), .O(gate446inter9));
  nand2 gate879(.a(s_47), .b(gate446inter3), .O(gate446inter10));
  nor2  gate880(.a(gate446inter10), .b(gate446inter9), .O(gate446inter11));
  nor2  gate881(.a(gate446inter11), .b(gate446inter6), .O(gate446inter12));
  nand2 gate882(.a(gate446inter12), .b(gate446inter1), .O(G1255));
nand2 gate447( .a(G15), .b(G1174), .O(G1256) );
nand2 gate448( .a(G1078), .b(G1174), .O(G1257) );
nand2 gate449( .a(G16), .b(G1177), .O(G1258) );

  xor2  gate575(.a(G1177), .b(G1081), .O(gate450inter0));
  nand2 gate576(.a(gate450inter0), .b(s_4), .O(gate450inter1));
  and2  gate577(.a(G1177), .b(G1081), .O(gate450inter2));
  inv1  gate578(.a(s_4), .O(gate450inter3));
  inv1  gate579(.a(s_5), .O(gate450inter4));
  nand2 gate580(.a(gate450inter4), .b(gate450inter3), .O(gate450inter5));
  nor2  gate581(.a(gate450inter5), .b(gate450inter2), .O(gate450inter6));
  inv1  gate582(.a(G1081), .O(gate450inter7));
  inv1  gate583(.a(G1177), .O(gate450inter8));
  nand2 gate584(.a(gate450inter8), .b(gate450inter7), .O(gate450inter9));
  nand2 gate585(.a(s_5), .b(gate450inter3), .O(gate450inter10));
  nor2  gate586(.a(gate450inter10), .b(gate450inter9), .O(gate450inter11));
  nor2  gate587(.a(gate450inter11), .b(gate450inter6), .O(gate450inter12));
  nand2 gate588(.a(gate450inter12), .b(gate450inter1), .O(G1259));

  xor2  gate2087(.a(G1180), .b(G17), .O(gate451inter0));
  nand2 gate2088(.a(gate451inter0), .b(s_220), .O(gate451inter1));
  and2  gate2089(.a(G1180), .b(G17), .O(gate451inter2));
  inv1  gate2090(.a(s_220), .O(gate451inter3));
  inv1  gate2091(.a(s_221), .O(gate451inter4));
  nand2 gate2092(.a(gate451inter4), .b(gate451inter3), .O(gate451inter5));
  nor2  gate2093(.a(gate451inter5), .b(gate451inter2), .O(gate451inter6));
  inv1  gate2094(.a(G17), .O(gate451inter7));
  inv1  gate2095(.a(G1180), .O(gate451inter8));
  nand2 gate2096(.a(gate451inter8), .b(gate451inter7), .O(gate451inter9));
  nand2 gate2097(.a(s_221), .b(gate451inter3), .O(gate451inter10));
  nor2  gate2098(.a(gate451inter10), .b(gate451inter9), .O(gate451inter11));
  nor2  gate2099(.a(gate451inter11), .b(gate451inter6), .O(gate451inter12));
  nand2 gate2100(.a(gate451inter12), .b(gate451inter1), .O(G1260));
nand2 gate452( .a(G1084), .b(G1180), .O(G1261) );
nand2 gate453( .a(G18), .b(G1183), .O(G1262) );
nand2 gate454( .a(G1087), .b(G1183), .O(G1263) );

  xor2  gate1247(.a(G1186), .b(G19), .O(gate455inter0));
  nand2 gate1248(.a(gate455inter0), .b(s_100), .O(gate455inter1));
  and2  gate1249(.a(G1186), .b(G19), .O(gate455inter2));
  inv1  gate1250(.a(s_100), .O(gate455inter3));
  inv1  gate1251(.a(s_101), .O(gate455inter4));
  nand2 gate1252(.a(gate455inter4), .b(gate455inter3), .O(gate455inter5));
  nor2  gate1253(.a(gate455inter5), .b(gate455inter2), .O(gate455inter6));
  inv1  gate1254(.a(G19), .O(gate455inter7));
  inv1  gate1255(.a(G1186), .O(gate455inter8));
  nand2 gate1256(.a(gate455inter8), .b(gate455inter7), .O(gate455inter9));
  nand2 gate1257(.a(s_101), .b(gate455inter3), .O(gate455inter10));
  nor2  gate1258(.a(gate455inter10), .b(gate455inter9), .O(gate455inter11));
  nor2  gate1259(.a(gate455inter11), .b(gate455inter6), .O(gate455inter12));
  nand2 gate1260(.a(gate455inter12), .b(gate455inter1), .O(G1264));
nand2 gate456( .a(G1090), .b(G1186), .O(G1265) );

  xor2  gate1135(.a(G1189), .b(G20), .O(gate457inter0));
  nand2 gate1136(.a(gate457inter0), .b(s_84), .O(gate457inter1));
  and2  gate1137(.a(G1189), .b(G20), .O(gate457inter2));
  inv1  gate1138(.a(s_84), .O(gate457inter3));
  inv1  gate1139(.a(s_85), .O(gate457inter4));
  nand2 gate1140(.a(gate457inter4), .b(gate457inter3), .O(gate457inter5));
  nor2  gate1141(.a(gate457inter5), .b(gate457inter2), .O(gate457inter6));
  inv1  gate1142(.a(G20), .O(gate457inter7));
  inv1  gate1143(.a(G1189), .O(gate457inter8));
  nand2 gate1144(.a(gate457inter8), .b(gate457inter7), .O(gate457inter9));
  nand2 gate1145(.a(s_85), .b(gate457inter3), .O(gate457inter10));
  nor2  gate1146(.a(gate457inter10), .b(gate457inter9), .O(gate457inter11));
  nor2  gate1147(.a(gate457inter11), .b(gate457inter6), .O(gate457inter12));
  nand2 gate1148(.a(gate457inter12), .b(gate457inter1), .O(G1266));
nand2 gate458( .a(G1093), .b(G1189), .O(G1267) );
nand2 gate459( .a(G21), .b(G1192), .O(G1268) );
nand2 gate460( .a(G1096), .b(G1192), .O(G1269) );

  xor2  gate1079(.a(G1195), .b(G22), .O(gate461inter0));
  nand2 gate1080(.a(gate461inter0), .b(s_76), .O(gate461inter1));
  and2  gate1081(.a(G1195), .b(G22), .O(gate461inter2));
  inv1  gate1082(.a(s_76), .O(gate461inter3));
  inv1  gate1083(.a(s_77), .O(gate461inter4));
  nand2 gate1084(.a(gate461inter4), .b(gate461inter3), .O(gate461inter5));
  nor2  gate1085(.a(gate461inter5), .b(gate461inter2), .O(gate461inter6));
  inv1  gate1086(.a(G22), .O(gate461inter7));
  inv1  gate1087(.a(G1195), .O(gate461inter8));
  nand2 gate1088(.a(gate461inter8), .b(gate461inter7), .O(gate461inter9));
  nand2 gate1089(.a(s_77), .b(gate461inter3), .O(gate461inter10));
  nor2  gate1090(.a(gate461inter10), .b(gate461inter9), .O(gate461inter11));
  nor2  gate1091(.a(gate461inter11), .b(gate461inter6), .O(gate461inter12));
  nand2 gate1092(.a(gate461inter12), .b(gate461inter1), .O(G1270));
nand2 gate462( .a(G1099), .b(G1195), .O(G1271) );
nand2 gate463( .a(G23), .b(G1198), .O(G1272) );

  xor2  gate603(.a(G1198), .b(G1102), .O(gate464inter0));
  nand2 gate604(.a(gate464inter0), .b(s_8), .O(gate464inter1));
  and2  gate605(.a(G1198), .b(G1102), .O(gate464inter2));
  inv1  gate606(.a(s_8), .O(gate464inter3));
  inv1  gate607(.a(s_9), .O(gate464inter4));
  nand2 gate608(.a(gate464inter4), .b(gate464inter3), .O(gate464inter5));
  nor2  gate609(.a(gate464inter5), .b(gate464inter2), .O(gate464inter6));
  inv1  gate610(.a(G1102), .O(gate464inter7));
  inv1  gate611(.a(G1198), .O(gate464inter8));
  nand2 gate612(.a(gate464inter8), .b(gate464inter7), .O(gate464inter9));
  nand2 gate613(.a(s_9), .b(gate464inter3), .O(gate464inter10));
  nor2  gate614(.a(gate464inter10), .b(gate464inter9), .O(gate464inter11));
  nor2  gate615(.a(gate464inter11), .b(gate464inter6), .O(gate464inter12));
  nand2 gate616(.a(gate464inter12), .b(gate464inter1), .O(G1273));

  xor2  gate547(.a(G1201), .b(G24), .O(gate465inter0));
  nand2 gate548(.a(gate465inter0), .b(s_0), .O(gate465inter1));
  and2  gate549(.a(G1201), .b(G24), .O(gate465inter2));
  inv1  gate550(.a(s_0), .O(gate465inter3));
  inv1  gate551(.a(s_1), .O(gate465inter4));
  nand2 gate552(.a(gate465inter4), .b(gate465inter3), .O(gate465inter5));
  nor2  gate553(.a(gate465inter5), .b(gate465inter2), .O(gate465inter6));
  inv1  gate554(.a(G24), .O(gate465inter7));
  inv1  gate555(.a(G1201), .O(gate465inter8));
  nand2 gate556(.a(gate465inter8), .b(gate465inter7), .O(gate465inter9));
  nand2 gate557(.a(s_1), .b(gate465inter3), .O(gate465inter10));
  nor2  gate558(.a(gate465inter10), .b(gate465inter9), .O(gate465inter11));
  nor2  gate559(.a(gate465inter11), .b(gate465inter6), .O(gate465inter12));
  nand2 gate560(.a(gate465inter12), .b(gate465inter1), .O(G1274));
nand2 gate466( .a(G1105), .b(G1201), .O(G1275) );

  xor2  gate1387(.a(G1204), .b(G25), .O(gate467inter0));
  nand2 gate1388(.a(gate467inter0), .b(s_120), .O(gate467inter1));
  and2  gate1389(.a(G1204), .b(G25), .O(gate467inter2));
  inv1  gate1390(.a(s_120), .O(gate467inter3));
  inv1  gate1391(.a(s_121), .O(gate467inter4));
  nand2 gate1392(.a(gate467inter4), .b(gate467inter3), .O(gate467inter5));
  nor2  gate1393(.a(gate467inter5), .b(gate467inter2), .O(gate467inter6));
  inv1  gate1394(.a(G25), .O(gate467inter7));
  inv1  gate1395(.a(G1204), .O(gate467inter8));
  nand2 gate1396(.a(gate467inter8), .b(gate467inter7), .O(gate467inter9));
  nand2 gate1397(.a(s_121), .b(gate467inter3), .O(gate467inter10));
  nor2  gate1398(.a(gate467inter10), .b(gate467inter9), .O(gate467inter11));
  nor2  gate1399(.a(gate467inter11), .b(gate467inter6), .O(gate467inter12));
  nand2 gate1400(.a(gate467inter12), .b(gate467inter1), .O(G1276));
nand2 gate468( .a(G1108), .b(G1204), .O(G1277) );
nand2 gate469( .a(G26), .b(G1207), .O(G1278) );

  xor2  gate2241(.a(G1207), .b(G1111), .O(gate470inter0));
  nand2 gate2242(.a(gate470inter0), .b(s_242), .O(gate470inter1));
  and2  gate2243(.a(G1207), .b(G1111), .O(gate470inter2));
  inv1  gate2244(.a(s_242), .O(gate470inter3));
  inv1  gate2245(.a(s_243), .O(gate470inter4));
  nand2 gate2246(.a(gate470inter4), .b(gate470inter3), .O(gate470inter5));
  nor2  gate2247(.a(gate470inter5), .b(gate470inter2), .O(gate470inter6));
  inv1  gate2248(.a(G1111), .O(gate470inter7));
  inv1  gate2249(.a(G1207), .O(gate470inter8));
  nand2 gate2250(.a(gate470inter8), .b(gate470inter7), .O(gate470inter9));
  nand2 gate2251(.a(s_243), .b(gate470inter3), .O(gate470inter10));
  nor2  gate2252(.a(gate470inter10), .b(gate470inter9), .O(gate470inter11));
  nor2  gate2253(.a(gate470inter11), .b(gate470inter6), .O(gate470inter12));
  nand2 gate2254(.a(gate470inter12), .b(gate470inter1), .O(G1279));

  xor2  gate1415(.a(G1210), .b(G27), .O(gate471inter0));
  nand2 gate1416(.a(gate471inter0), .b(s_124), .O(gate471inter1));
  and2  gate1417(.a(G1210), .b(G27), .O(gate471inter2));
  inv1  gate1418(.a(s_124), .O(gate471inter3));
  inv1  gate1419(.a(s_125), .O(gate471inter4));
  nand2 gate1420(.a(gate471inter4), .b(gate471inter3), .O(gate471inter5));
  nor2  gate1421(.a(gate471inter5), .b(gate471inter2), .O(gate471inter6));
  inv1  gate1422(.a(G27), .O(gate471inter7));
  inv1  gate1423(.a(G1210), .O(gate471inter8));
  nand2 gate1424(.a(gate471inter8), .b(gate471inter7), .O(gate471inter9));
  nand2 gate1425(.a(s_125), .b(gate471inter3), .O(gate471inter10));
  nor2  gate1426(.a(gate471inter10), .b(gate471inter9), .O(gate471inter11));
  nor2  gate1427(.a(gate471inter11), .b(gate471inter6), .O(gate471inter12));
  nand2 gate1428(.a(gate471inter12), .b(gate471inter1), .O(G1280));

  xor2  gate2101(.a(G1210), .b(G1114), .O(gate472inter0));
  nand2 gate2102(.a(gate472inter0), .b(s_222), .O(gate472inter1));
  and2  gate2103(.a(G1210), .b(G1114), .O(gate472inter2));
  inv1  gate2104(.a(s_222), .O(gate472inter3));
  inv1  gate2105(.a(s_223), .O(gate472inter4));
  nand2 gate2106(.a(gate472inter4), .b(gate472inter3), .O(gate472inter5));
  nor2  gate2107(.a(gate472inter5), .b(gate472inter2), .O(gate472inter6));
  inv1  gate2108(.a(G1114), .O(gate472inter7));
  inv1  gate2109(.a(G1210), .O(gate472inter8));
  nand2 gate2110(.a(gate472inter8), .b(gate472inter7), .O(gate472inter9));
  nand2 gate2111(.a(s_223), .b(gate472inter3), .O(gate472inter10));
  nor2  gate2112(.a(gate472inter10), .b(gate472inter9), .O(gate472inter11));
  nor2  gate2113(.a(gate472inter11), .b(gate472inter6), .O(gate472inter12));
  nand2 gate2114(.a(gate472inter12), .b(gate472inter1), .O(G1281));

  xor2  gate1737(.a(G1213), .b(G28), .O(gate473inter0));
  nand2 gate1738(.a(gate473inter0), .b(s_170), .O(gate473inter1));
  and2  gate1739(.a(G1213), .b(G28), .O(gate473inter2));
  inv1  gate1740(.a(s_170), .O(gate473inter3));
  inv1  gate1741(.a(s_171), .O(gate473inter4));
  nand2 gate1742(.a(gate473inter4), .b(gate473inter3), .O(gate473inter5));
  nor2  gate1743(.a(gate473inter5), .b(gate473inter2), .O(gate473inter6));
  inv1  gate1744(.a(G28), .O(gate473inter7));
  inv1  gate1745(.a(G1213), .O(gate473inter8));
  nand2 gate1746(.a(gate473inter8), .b(gate473inter7), .O(gate473inter9));
  nand2 gate1747(.a(s_171), .b(gate473inter3), .O(gate473inter10));
  nor2  gate1748(.a(gate473inter10), .b(gate473inter9), .O(gate473inter11));
  nor2  gate1749(.a(gate473inter11), .b(gate473inter6), .O(gate473inter12));
  nand2 gate1750(.a(gate473inter12), .b(gate473inter1), .O(G1282));
nand2 gate474( .a(G1117), .b(G1213), .O(G1283) );
nand2 gate475( .a(G29), .b(G1216), .O(G1284) );
nand2 gate476( .a(G1120), .b(G1216), .O(G1285) );
nand2 gate477( .a(G30), .b(G1219), .O(G1286) );

  xor2  gate1905(.a(G1219), .b(G1123), .O(gate478inter0));
  nand2 gate1906(.a(gate478inter0), .b(s_194), .O(gate478inter1));
  and2  gate1907(.a(G1219), .b(G1123), .O(gate478inter2));
  inv1  gate1908(.a(s_194), .O(gate478inter3));
  inv1  gate1909(.a(s_195), .O(gate478inter4));
  nand2 gate1910(.a(gate478inter4), .b(gate478inter3), .O(gate478inter5));
  nor2  gate1911(.a(gate478inter5), .b(gate478inter2), .O(gate478inter6));
  inv1  gate1912(.a(G1123), .O(gate478inter7));
  inv1  gate1913(.a(G1219), .O(gate478inter8));
  nand2 gate1914(.a(gate478inter8), .b(gate478inter7), .O(gate478inter9));
  nand2 gate1915(.a(s_195), .b(gate478inter3), .O(gate478inter10));
  nor2  gate1916(.a(gate478inter10), .b(gate478inter9), .O(gate478inter11));
  nor2  gate1917(.a(gate478inter11), .b(gate478inter6), .O(gate478inter12));
  nand2 gate1918(.a(gate478inter12), .b(gate478inter1), .O(G1287));
nand2 gate479( .a(G31), .b(G1222), .O(G1288) );
nand2 gate480( .a(G1126), .b(G1222), .O(G1289) );
nand2 gate481( .a(G32), .b(G1225), .O(G1290) );
nand2 gate482( .a(G1129), .b(G1225), .O(G1291) );
nand2 gate483( .a(G1228), .b(G1229), .O(G1292) );
nand2 gate484( .a(G1230), .b(G1231), .O(G1293) );
nand2 gate485( .a(G1232), .b(G1233), .O(G1294) );
nand2 gate486( .a(G1234), .b(G1235), .O(G1295) );

  xor2  gate1877(.a(G1237), .b(G1236), .O(gate487inter0));
  nand2 gate1878(.a(gate487inter0), .b(s_190), .O(gate487inter1));
  and2  gate1879(.a(G1237), .b(G1236), .O(gate487inter2));
  inv1  gate1880(.a(s_190), .O(gate487inter3));
  inv1  gate1881(.a(s_191), .O(gate487inter4));
  nand2 gate1882(.a(gate487inter4), .b(gate487inter3), .O(gate487inter5));
  nor2  gate1883(.a(gate487inter5), .b(gate487inter2), .O(gate487inter6));
  inv1  gate1884(.a(G1236), .O(gate487inter7));
  inv1  gate1885(.a(G1237), .O(gate487inter8));
  nand2 gate1886(.a(gate487inter8), .b(gate487inter7), .O(gate487inter9));
  nand2 gate1887(.a(s_191), .b(gate487inter3), .O(gate487inter10));
  nor2  gate1888(.a(gate487inter10), .b(gate487inter9), .O(gate487inter11));
  nor2  gate1889(.a(gate487inter11), .b(gate487inter6), .O(gate487inter12));
  nand2 gate1890(.a(gate487inter12), .b(gate487inter1), .O(G1296));
nand2 gate488( .a(G1238), .b(G1239), .O(G1297) );
nand2 gate489( .a(G1240), .b(G1241), .O(G1298) );
nand2 gate490( .a(G1242), .b(G1243), .O(G1299) );

  xor2  gate925(.a(G1245), .b(G1244), .O(gate491inter0));
  nand2 gate926(.a(gate491inter0), .b(s_54), .O(gate491inter1));
  and2  gate927(.a(G1245), .b(G1244), .O(gate491inter2));
  inv1  gate928(.a(s_54), .O(gate491inter3));
  inv1  gate929(.a(s_55), .O(gate491inter4));
  nand2 gate930(.a(gate491inter4), .b(gate491inter3), .O(gate491inter5));
  nor2  gate931(.a(gate491inter5), .b(gate491inter2), .O(gate491inter6));
  inv1  gate932(.a(G1244), .O(gate491inter7));
  inv1  gate933(.a(G1245), .O(gate491inter8));
  nand2 gate934(.a(gate491inter8), .b(gate491inter7), .O(gate491inter9));
  nand2 gate935(.a(s_55), .b(gate491inter3), .O(gate491inter10));
  nor2  gate936(.a(gate491inter10), .b(gate491inter9), .O(gate491inter11));
  nor2  gate937(.a(gate491inter11), .b(gate491inter6), .O(gate491inter12));
  nand2 gate938(.a(gate491inter12), .b(gate491inter1), .O(G1300));
nand2 gate492( .a(G1246), .b(G1247), .O(G1301) );

  xor2  gate2171(.a(G1249), .b(G1248), .O(gate493inter0));
  nand2 gate2172(.a(gate493inter0), .b(s_232), .O(gate493inter1));
  and2  gate2173(.a(G1249), .b(G1248), .O(gate493inter2));
  inv1  gate2174(.a(s_232), .O(gate493inter3));
  inv1  gate2175(.a(s_233), .O(gate493inter4));
  nand2 gate2176(.a(gate493inter4), .b(gate493inter3), .O(gate493inter5));
  nor2  gate2177(.a(gate493inter5), .b(gate493inter2), .O(gate493inter6));
  inv1  gate2178(.a(G1248), .O(gate493inter7));
  inv1  gate2179(.a(G1249), .O(gate493inter8));
  nand2 gate2180(.a(gate493inter8), .b(gate493inter7), .O(gate493inter9));
  nand2 gate2181(.a(s_233), .b(gate493inter3), .O(gate493inter10));
  nor2  gate2182(.a(gate493inter10), .b(gate493inter9), .O(gate493inter11));
  nor2  gate2183(.a(gate493inter11), .b(gate493inter6), .O(gate493inter12));
  nand2 gate2184(.a(gate493inter12), .b(gate493inter1), .O(G1302));
nand2 gate494( .a(G1250), .b(G1251), .O(G1303) );

  xor2  gate701(.a(G1253), .b(G1252), .O(gate495inter0));
  nand2 gate702(.a(gate495inter0), .b(s_22), .O(gate495inter1));
  and2  gate703(.a(G1253), .b(G1252), .O(gate495inter2));
  inv1  gate704(.a(s_22), .O(gate495inter3));
  inv1  gate705(.a(s_23), .O(gate495inter4));
  nand2 gate706(.a(gate495inter4), .b(gate495inter3), .O(gate495inter5));
  nor2  gate707(.a(gate495inter5), .b(gate495inter2), .O(gate495inter6));
  inv1  gate708(.a(G1252), .O(gate495inter7));
  inv1  gate709(.a(G1253), .O(gate495inter8));
  nand2 gate710(.a(gate495inter8), .b(gate495inter7), .O(gate495inter9));
  nand2 gate711(.a(s_23), .b(gate495inter3), .O(gate495inter10));
  nor2  gate712(.a(gate495inter10), .b(gate495inter9), .O(gate495inter11));
  nor2  gate713(.a(gate495inter11), .b(gate495inter6), .O(gate495inter12));
  nand2 gate714(.a(gate495inter12), .b(gate495inter1), .O(G1304));

  xor2  gate1597(.a(G1255), .b(G1254), .O(gate496inter0));
  nand2 gate1598(.a(gate496inter0), .b(s_150), .O(gate496inter1));
  and2  gate1599(.a(G1255), .b(G1254), .O(gate496inter2));
  inv1  gate1600(.a(s_150), .O(gate496inter3));
  inv1  gate1601(.a(s_151), .O(gate496inter4));
  nand2 gate1602(.a(gate496inter4), .b(gate496inter3), .O(gate496inter5));
  nor2  gate1603(.a(gate496inter5), .b(gate496inter2), .O(gate496inter6));
  inv1  gate1604(.a(G1254), .O(gate496inter7));
  inv1  gate1605(.a(G1255), .O(gate496inter8));
  nand2 gate1606(.a(gate496inter8), .b(gate496inter7), .O(gate496inter9));
  nand2 gate1607(.a(s_151), .b(gate496inter3), .O(gate496inter10));
  nor2  gate1608(.a(gate496inter10), .b(gate496inter9), .O(gate496inter11));
  nor2  gate1609(.a(gate496inter11), .b(gate496inter6), .O(gate496inter12));
  nand2 gate1610(.a(gate496inter12), .b(gate496inter1), .O(G1305));

  xor2  gate855(.a(G1257), .b(G1256), .O(gate497inter0));
  nand2 gate856(.a(gate497inter0), .b(s_44), .O(gate497inter1));
  and2  gate857(.a(G1257), .b(G1256), .O(gate497inter2));
  inv1  gate858(.a(s_44), .O(gate497inter3));
  inv1  gate859(.a(s_45), .O(gate497inter4));
  nand2 gate860(.a(gate497inter4), .b(gate497inter3), .O(gate497inter5));
  nor2  gate861(.a(gate497inter5), .b(gate497inter2), .O(gate497inter6));
  inv1  gate862(.a(G1256), .O(gate497inter7));
  inv1  gate863(.a(G1257), .O(gate497inter8));
  nand2 gate864(.a(gate497inter8), .b(gate497inter7), .O(gate497inter9));
  nand2 gate865(.a(s_45), .b(gate497inter3), .O(gate497inter10));
  nor2  gate866(.a(gate497inter10), .b(gate497inter9), .O(gate497inter11));
  nor2  gate867(.a(gate497inter11), .b(gate497inter6), .O(gate497inter12));
  nand2 gate868(.a(gate497inter12), .b(gate497inter1), .O(G1306));
nand2 gate498( .a(G1258), .b(G1259), .O(G1307) );
nand2 gate499( .a(G1260), .b(G1261), .O(G1308) );
nand2 gate500( .a(G1262), .b(G1263), .O(G1309) );
nand2 gate501( .a(G1264), .b(G1265), .O(G1310) );
nand2 gate502( .a(G1266), .b(G1267), .O(G1311) );

  xor2  gate1121(.a(G1269), .b(G1268), .O(gate503inter0));
  nand2 gate1122(.a(gate503inter0), .b(s_82), .O(gate503inter1));
  and2  gate1123(.a(G1269), .b(G1268), .O(gate503inter2));
  inv1  gate1124(.a(s_82), .O(gate503inter3));
  inv1  gate1125(.a(s_83), .O(gate503inter4));
  nand2 gate1126(.a(gate503inter4), .b(gate503inter3), .O(gate503inter5));
  nor2  gate1127(.a(gate503inter5), .b(gate503inter2), .O(gate503inter6));
  inv1  gate1128(.a(G1268), .O(gate503inter7));
  inv1  gate1129(.a(G1269), .O(gate503inter8));
  nand2 gate1130(.a(gate503inter8), .b(gate503inter7), .O(gate503inter9));
  nand2 gate1131(.a(s_83), .b(gate503inter3), .O(gate503inter10));
  nor2  gate1132(.a(gate503inter10), .b(gate503inter9), .O(gate503inter11));
  nor2  gate1133(.a(gate503inter11), .b(gate503inter6), .O(gate503inter12));
  nand2 gate1134(.a(gate503inter12), .b(gate503inter1), .O(G1312));
nand2 gate504( .a(G1270), .b(G1271), .O(G1313) );
nand2 gate505( .a(G1272), .b(G1273), .O(G1314) );
nand2 gate506( .a(G1274), .b(G1275), .O(G1315) );

  xor2  gate1345(.a(G1277), .b(G1276), .O(gate507inter0));
  nand2 gate1346(.a(gate507inter0), .b(s_114), .O(gate507inter1));
  and2  gate1347(.a(G1277), .b(G1276), .O(gate507inter2));
  inv1  gate1348(.a(s_114), .O(gate507inter3));
  inv1  gate1349(.a(s_115), .O(gate507inter4));
  nand2 gate1350(.a(gate507inter4), .b(gate507inter3), .O(gate507inter5));
  nor2  gate1351(.a(gate507inter5), .b(gate507inter2), .O(gate507inter6));
  inv1  gate1352(.a(G1276), .O(gate507inter7));
  inv1  gate1353(.a(G1277), .O(gate507inter8));
  nand2 gate1354(.a(gate507inter8), .b(gate507inter7), .O(gate507inter9));
  nand2 gate1355(.a(s_115), .b(gate507inter3), .O(gate507inter10));
  nor2  gate1356(.a(gate507inter10), .b(gate507inter9), .O(gate507inter11));
  nor2  gate1357(.a(gate507inter11), .b(gate507inter6), .O(gate507inter12));
  nand2 gate1358(.a(gate507inter12), .b(gate507inter1), .O(G1316));
nand2 gate508( .a(G1278), .b(G1279), .O(G1317) );

  xor2  gate757(.a(G1281), .b(G1280), .O(gate509inter0));
  nand2 gate758(.a(gate509inter0), .b(s_30), .O(gate509inter1));
  and2  gate759(.a(G1281), .b(G1280), .O(gate509inter2));
  inv1  gate760(.a(s_30), .O(gate509inter3));
  inv1  gate761(.a(s_31), .O(gate509inter4));
  nand2 gate762(.a(gate509inter4), .b(gate509inter3), .O(gate509inter5));
  nor2  gate763(.a(gate509inter5), .b(gate509inter2), .O(gate509inter6));
  inv1  gate764(.a(G1280), .O(gate509inter7));
  inv1  gate765(.a(G1281), .O(gate509inter8));
  nand2 gate766(.a(gate509inter8), .b(gate509inter7), .O(gate509inter9));
  nand2 gate767(.a(s_31), .b(gate509inter3), .O(gate509inter10));
  nor2  gate768(.a(gate509inter10), .b(gate509inter9), .O(gate509inter11));
  nor2  gate769(.a(gate509inter11), .b(gate509inter6), .O(gate509inter12));
  nand2 gate770(.a(gate509inter12), .b(gate509inter1), .O(G1318));
nand2 gate510( .a(G1282), .b(G1283), .O(G1319) );

  xor2  gate1611(.a(G1285), .b(G1284), .O(gate511inter0));
  nand2 gate1612(.a(gate511inter0), .b(s_152), .O(gate511inter1));
  and2  gate1613(.a(G1285), .b(G1284), .O(gate511inter2));
  inv1  gate1614(.a(s_152), .O(gate511inter3));
  inv1  gate1615(.a(s_153), .O(gate511inter4));
  nand2 gate1616(.a(gate511inter4), .b(gate511inter3), .O(gate511inter5));
  nor2  gate1617(.a(gate511inter5), .b(gate511inter2), .O(gate511inter6));
  inv1  gate1618(.a(G1284), .O(gate511inter7));
  inv1  gate1619(.a(G1285), .O(gate511inter8));
  nand2 gate1620(.a(gate511inter8), .b(gate511inter7), .O(gate511inter9));
  nand2 gate1621(.a(s_153), .b(gate511inter3), .O(gate511inter10));
  nor2  gate1622(.a(gate511inter10), .b(gate511inter9), .O(gate511inter11));
  nor2  gate1623(.a(gate511inter11), .b(gate511inter6), .O(gate511inter12));
  nand2 gate1624(.a(gate511inter12), .b(gate511inter1), .O(G1320));

  xor2  gate1065(.a(G1287), .b(G1286), .O(gate512inter0));
  nand2 gate1066(.a(gate512inter0), .b(s_74), .O(gate512inter1));
  and2  gate1067(.a(G1287), .b(G1286), .O(gate512inter2));
  inv1  gate1068(.a(s_74), .O(gate512inter3));
  inv1  gate1069(.a(s_75), .O(gate512inter4));
  nand2 gate1070(.a(gate512inter4), .b(gate512inter3), .O(gate512inter5));
  nor2  gate1071(.a(gate512inter5), .b(gate512inter2), .O(gate512inter6));
  inv1  gate1072(.a(G1286), .O(gate512inter7));
  inv1  gate1073(.a(G1287), .O(gate512inter8));
  nand2 gate1074(.a(gate512inter8), .b(gate512inter7), .O(gate512inter9));
  nand2 gate1075(.a(s_75), .b(gate512inter3), .O(gate512inter10));
  nor2  gate1076(.a(gate512inter10), .b(gate512inter9), .O(gate512inter11));
  nor2  gate1077(.a(gate512inter11), .b(gate512inter6), .O(gate512inter12));
  nand2 gate1078(.a(gate512inter12), .b(gate512inter1), .O(G1321));
nand2 gate513( .a(G1288), .b(G1289), .O(G1322) );

  xor2  gate2059(.a(G1291), .b(G1290), .O(gate514inter0));
  nand2 gate2060(.a(gate514inter0), .b(s_216), .O(gate514inter1));
  and2  gate2061(.a(G1291), .b(G1290), .O(gate514inter2));
  inv1  gate2062(.a(s_216), .O(gate514inter3));
  inv1  gate2063(.a(s_217), .O(gate514inter4));
  nand2 gate2064(.a(gate514inter4), .b(gate514inter3), .O(gate514inter5));
  nor2  gate2065(.a(gate514inter5), .b(gate514inter2), .O(gate514inter6));
  inv1  gate2066(.a(G1290), .O(gate514inter7));
  inv1  gate2067(.a(G1291), .O(gate514inter8));
  nand2 gate2068(.a(gate514inter8), .b(gate514inter7), .O(gate514inter9));
  nand2 gate2069(.a(s_217), .b(gate514inter3), .O(gate514inter10));
  nor2  gate2070(.a(gate514inter10), .b(gate514inter9), .O(gate514inter11));
  nor2  gate2071(.a(gate514inter11), .b(gate514inter6), .O(gate514inter12));
  nand2 gate2072(.a(gate514inter12), .b(gate514inter1), .O(G1323));
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule