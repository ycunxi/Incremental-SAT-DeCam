module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);

input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;//RE__PI;

input s_0,s_1;//RE__ALLOW(00,01,10,11);
input s_2,s_3;//RE__ALLOW(00,01,10,11);
input s_4,s_5;//RE__ALLOW(00,01,10,11);
input s_6,s_7;//RE__ALLOW(00,01,10,11);
input s_8,s_9;//RE__ALLOW(00,01,10,11);
input s_10,s_11;//RE__ALLOW(00,01,10,11);
input s_12,s_13;//RE__ALLOW(00,01,10,11);
input s_14,s_15;//RE__ALLOW(00,01,10,11);
input s_16,s_17;//RE__ALLOW(00,01,10,11);
input s_18,s_19;//RE__ALLOW(00,01,10,11);
input s_20,s_21;//RE__ALLOW(00,01,10,11);
input s_22,s_23;//RE__ALLOW(00,01,10,11);
input s_24,s_25;//RE__ALLOW(00,01,10,11);
input s_26,s_27;//RE__ALLOW(00,01,10,11);
input s_28,s_29;//RE__ALLOW(00,01,10,11);
input s_30,s_31;//RE__ALLOW(00,01,10,11);
input s_32,s_33;//RE__ALLOW(00,01,10,11);
input s_34,s_35;//RE__ALLOW(00,01,10,11);
input s_36,s_37;//RE__ALLOW(00,01,10,11);
input s_38,s_39;//RE__ALLOW(00,01,10,11);
input s_40,s_41;//RE__ALLOW(00,01,10,11);
input s_42,s_43;//RE__ALLOW(00,01,10,11);
input s_44,s_45;//RE__ALLOW(00,01,10,11);
input s_46,s_47;//RE__ALLOW(00,01,10,11);
input s_48,s_49;//RE__ALLOW(00,01,10,11);
input s_50,s_51;//RE__ALLOW(00,01,10,11);
input s_52,s_53;//RE__ALLOW(00,01,10,11);
input s_54,s_55;//RE__ALLOW(00,01,10,11);
input s_56,s_57;//RE__ALLOW(00,01,10,11);
input s_58,s_59;//RE__ALLOW(00,01,10,11);
input s_60,s_61;//RE__ALLOW(00,01,10,11);
input s_62,s_63;//RE__ALLOW(00,01,10,11);
input s_64,s_65;//RE__ALLOW(00,01,10,11);
input s_66,s_67;//RE__ALLOW(00,01,10,11);
input s_68,s_69;//RE__ALLOW(00,01,10,11);
input s_70,s_71;//RE__ALLOW(00,01,10,11);
input s_72,s_73;//RE__ALLOW(00,01,10,11);
input s_74,s_75;//RE__ALLOW(00,01,10,11);
input s_76,s_77;//RE__ALLOW(00,01,10,11);
input s_78,s_79;//RE__ALLOW(00,01,10,11);
input s_80,s_81;//RE__ALLOW(00,01,10,11);
input s_82,s_83;//RE__ALLOW(00,01,10,11);
input s_84,s_85;//RE__ALLOW(00,01,10,11);
input s_86,s_87;//RE__ALLOW(00,01,10,11);
input s_88,s_89;//RE__ALLOW(00,01,10,11);
input s_90,s_91;//RE__ALLOW(00,01,10,11);
input s_92,s_93;//RE__ALLOW(00,01,10,11);
input s_94,s_95;//RE__ALLOW(00,01,10,11);
input s_96,s_97;//RE__ALLOW(00,01,10,11);
input s_98,s_99;//RE__ALLOW(00,01,10,11);
input s_100,s_101;//RE__ALLOW(00,01,10,11);
input s_102,s_103;//RE__ALLOW(00,01,10,11);
input s_104,s_105;//RE__ALLOW(00,01,10,11);
input s_106,s_107;//RE__ALLOW(00,01,10,11);
input s_108,s_109;//RE__ALLOW(00,01,10,11);
input s_110,s_111;//RE__ALLOW(00,01,10,11);
input s_112,s_113;//RE__ALLOW(00,01,10,11);
input s_114,s_115;//RE__ALLOW(00,01,10,11);
input s_116,s_117;//RE__ALLOW(00,01,10,11);
input s_118,s_119;//RE__ALLOW(00,01,10,11);
input s_120,s_121;//RE__ALLOW(00,01,10,11);
input s_122,s_123;//RE__ALLOW(00,01,10,11);
input s_124,s_125;//RE__ALLOW(00,01,10,11);
input s_126,s_127;//RE__ALLOW(00,01,10,11);
input s_128,s_129;//RE__ALLOW(00,01,10,11);
input s_130,s_131;//RE__ALLOW(00,01,10,11);
input s_132,s_133;//RE__ALLOW(00,01,10,11);
input s_134,s_135;//RE__ALLOW(00,01,10,11);
input s_136,s_137;//RE__ALLOW(00,01,10,11);
input s_138,s_139;//RE__ALLOW(00,01,10,11);
input s_140,s_141;//RE__ALLOW(00,01,10,11);
input s_142,s_143;//RE__ALLOW(00,01,10,11);
input s_144,s_145;//RE__ALLOW(00,01,10,11);
input s_146,s_147;//RE__ALLOW(00,01,10,11);
input s_148,s_149;//RE__ALLOW(00,01,10,11);
input s_150,s_151;//RE__ALLOW(00,01,10,11);
input s_152,s_153;//RE__ALLOW(00,01,10,11);
input s_154,s_155;//RE__ALLOW(00,01,10,11);
input s_156,s_157;//RE__ALLOW(00,01,10,11);
input s_158,s_159;//RE__ALLOW(00,01,10,11);
input s_160,s_161;//RE__ALLOW(00,01,10,11);
input s_162,s_163;//RE__ALLOW(00,01,10,11);
input s_164,s_165;//RE__ALLOW(00,01,10,11);
input s_166,s_167;//RE__ALLOW(00,01,10,11);
input s_168,s_169;//RE__ALLOW(00,01,10,11);
input s_170,s_171;//RE__ALLOW(00,01,10,11);
input s_172,s_173;//RE__ALLOW(00,01,10,11);
input s_174,s_175;//RE__ALLOW(00,01,10,11);
input s_176,s_177;//RE__ALLOW(00,01,10,11);
input s_178,s_179;//RE__ALLOW(00,01,10,11);
input s_180,s_181;//RE__ALLOW(00,01,10,11);
input s_182,s_183;//RE__ALLOW(00,01,10,11);
input s_184,s_185;//RE__ALLOW(00,01,10,11);
input s_186,s_187;//RE__ALLOW(00,01,10,11);
input s_188,s_189;//RE__ALLOW(00,01,10,11);
input s_190,s_191;//RE__ALLOW(00,01,10,11);
input s_192,s_193;//RE__ALLOW(00,01,10,11);
input s_194,s_195;//RE__ALLOW(00,01,10,11);
input s_196,s_197;//RE__ALLOW(00,01,10,11);
input s_198,s_199;//RE__ALLOW(00,01,10,11);
input s_200,s_201;//RE__ALLOW(00,01,10,11);
input s_202,s_203;//RE__ALLOW(00,01,10,11);
input s_204,s_205;//RE__ALLOW(00,01,10,11);
input s_206,s_207;//RE__ALLOW(00,01,10,11);
input s_208,s_209;//RE__ALLOW(00,01,10,11);
input s_210,s_211;//RE__ALLOW(00,01,10,11);
input s_212,s_213;//RE__ALLOW(00,01,10,11);
input s_214,s_215;//RE__ALLOW(00,01,10,11);
input s_216,s_217;//RE__ALLOW(00,01,10,11);
input s_218,s_219;//RE__ALLOW(00,01,10,11);
input s_220,s_221;//RE__ALLOW(00,01,10,11);
input s_222,s_223;//RE__ALLOW(00,01,10,11);
input s_224,s_225;//RE__ALLOW(00,01,10,11);
input s_226,s_227;//RE__ALLOW(00,01,10,11);
input s_228,s_229;//RE__ALLOW(00,01,10,11);
input s_230,s_231;//RE__ALLOW(00,01,10,11);
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;

  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate402inter0, gate402inter1, gate402inter2, gate402inter3, gate402inter4, gate402inter5, gate402inter6, gate402inter7, gate402inter8, gate402inter9, gate402inter10, gate402inter11, gate402inter12, gate65inter0, gate65inter1, gate65inter2, gate65inter3, gate65inter4, gate65inter5, gate65inter6, gate65inter7, gate65inter8, gate65inter9, gate65inter10, gate65inter11, gate65inter12, gate276inter0, gate276inter1, gate276inter2, gate276inter3, gate276inter4, gate276inter5, gate276inter6, gate276inter7, gate276inter8, gate276inter9, gate276inter10, gate276inter11, gate276inter12, gate428inter0, gate428inter1, gate428inter2, gate428inter3, gate428inter4, gate428inter5, gate428inter6, gate428inter7, gate428inter8, gate428inter9, gate428inter10, gate428inter11, gate428inter12, gate440inter0, gate440inter1, gate440inter2, gate440inter3, gate440inter4, gate440inter5, gate440inter6, gate440inter7, gate440inter8, gate440inter9, gate440inter10, gate440inter11, gate440inter12, gate434inter0, gate434inter1, gate434inter2, gate434inter3, gate434inter4, gate434inter5, gate434inter6, gate434inter7, gate434inter8, gate434inter9, gate434inter10, gate434inter11, gate434inter12, gate251inter0, gate251inter1, gate251inter2, gate251inter3, gate251inter4, gate251inter5, gate251inter6, gate251inter7, gate251inter8, gate251inter9, gate251inter10, gate251inter11, gate251inter12, gate225inter0, gate225inter1, gate225inter2, gate225inter3, gate225inter4, gate225inter5, gate225inter6, gate225inter7, gate225inter8, gate225inter9, gate225inter10, gate225inter11, gate225inter12, gate157inter0, gate157inter1, gate157inter2, gate157inter3, gate157inter4, gate157inter5, gate157inter6, gate157inter7, gate157inter8, gate157inter9, gate157inter10, gate157inter11, gate157inter12, gate92inter0, gate92inter1, gate92inter2, gate92inter3, gate92inter4, gate92inter5, gate92inter6, gate92inter7, gate92inter8, gate92inter9, gate92inter10, gate92inter11, gate92inter12, gate153inter0, gate153inter1, gate153inter2, gate153inter3, gate153inter4, gate153inter5, gate153inter6, gate153inter7, gate153inter8, gate153inter9, gate153inter10, gate153inter11, gate153inter12, gate469inter0, gate469inter1, gate469inter2, gate469inter3, gate469inter4, gate469inter5, gate469inter6, gate469inter7, gate469inter8, gate469inter9, gate469inter10, gate469inter11, gate469inter12, gate423inter0, gate423inter1, gate423inter2, gate423inter3, gate423inter4, gate423inter5, gate423inter6, gate423inter7, gate423inter8, gate423inter9, gate423inter10, gate423inter11, gate423inter12, gate421inter0, gate421inter1, gate421inter2, gate421inter3, gate421inter4, gate421inter5, gate421inter6, gate421inter7, gate421inter8, gate421inter9, gate421inter10, gate421inter11, gate421inter12, gate248inter0, gate248inter1, gate248inter2, gate248inter3, gate248inter4, gate248inter5, gate248inter6, gate248inter7, gate248inter8, gate248inter9, gate248inter10, gate248inter11, gate248inter12, gate261inter0, gate261inter1, gate261inter2, gate261inter3, gate261inter4, gate261inter5, gate261inter6, gate261inter7, gate261inter8, gate261inter9, gate261inter10, gate261inter11, gate261inter12, gate501inter0, gate501inter1, gate501inter2, gate501inter3, gate501inter4, gate501inter5, gate501inter6, gate501inter7, gate501inter8, gate501inter9, gate501inter10, gate501inter11, gate501inter12, gate74inter0, gate74inter1, gate74inter2, gate74inter3, gate74inter4, gate74inter5, gate74inter6, gate74inter7, gate74inter8, gate74inter9, gate74inter10, gate74inter11, gate74inter12, gate123inter0, gate123inter1, gate123inter2, gate123inter3, gate123inter4, gate123inter5, gate123inter6, gate123inter7, gate123inter8, gate123inter9, gate123inter10, gate123inter11, gate123inter12, gate513inter0, gate513inter1, gate513inter2, gate513inter3, gate513inter4, gate513inter5, gate513inter6, gate513inter7, gate513inter8, gate513inter9, gate513inter10, gate513inter11, gate513inter12, gate409inter0, gate409inter1, gate409inter2, gate409inter3, gate409inter4, gate409inter5, gate409inter6, gate409inter7, gate409inter8, gate409inter9, gate409inter10, gate409inter11, gate409inter12, gate97inter0, gate97inter1, gate97inter2, gate97inter3, gate97inter4, gate97inter5, gate97inter6, gate97inter7, gate97inter8, gate97inter9, gate97inter10, gate97inter11, gate97inter12, gate241inter0, gate241inter1, gate241inter2, gate241inter3, gate241inter4, gate241inter5, gate241inter6, gate241inter7, gate241inter8, gate241inter9, gate241inter10, gate241inter11, gate241inter12, gate128inter0, gate128inter1, gate128inter2, gate128inter3, gate128inter4, gate128inter5, gate128inter6, gate128inter7, gate128inter8, gate128inter9, gate128inter10, gate128inter11, gate128inter12, gate209inter0, gate209inter1, gate209inter2, gate209inter3, gate209inter4, gate209inter5, gate209inter6, gate209inter7, gate209inter8, gate209inter9, gate209inter10, gate209inter11, gate209inter12, gate63inter0, gate63inter1, gate63inter2, gate63inter3, gate63inter4, gate63inter5, gate63inter6, gate63inter7, gate63inter8, gate63inter9, gate63inter10, gate63inter11, gate63inter12, gate234inter0, gate234inter1, gate234inter2, gate234inter3, gate234inter4, gate234inter5, gate234inter6, gate234inter7, gate234inter8, gate234inter9, gate234inter10, gate234inter11, gate234inter12, gate258inter0, gate258inter1, gate258inter2, gate258inter3, gate258inter4, gate258inter5, gate258inter6, gate258inter7, gate258inter8, gate258inter9, gate258inter10, gate258inter11, gate258inter12, gate411inter0, gate411inter1, gate411inter2, gate411inter3, gate411inter4, gate411inter5, gate411inter6, gate411inter7, gate411inter8, gate411inter9, gate411inter10, gate411inter11, gate411inter12, gate275inter0, gate275inter1, gate275inter2, gate275inter3, gate275inter4, gate275inter5, gate275inter6, gate275inter7, gate275inter8, gate275inter9, gate275inter10, gate275inter11, gate275inter12, gate19inter0, gate19inter1, gate19inter2, gate19inter3, gate19inter4, gate19inter5, gate19inter6, gate19inter7, gate19inter8, gate19inter9, gate19inter10, gate19inter11, gate19inter12, gate29inter0, gate29inter1, gate29inter2, gate29inter3, gate29inter4, gate29inter5, gate29inter6, gate29inter7, gate29inter8, gate29inter9, gate29inter10, gate29inter11, gate29inter12, gate94inter0, gate94inter1, gate94inter2, gate94inter3, gate94inter4, gate94inter5, gate94inter6, gate94inter7, gate94inter8, gate94inter9, gate94inter10, gate94inter11, gate94inter12, gate193inter0, gate193inter1, gate193inter2, gate193inter3, gate193inter4, gate193inter5, gate193inter6, gate193inter7, gate193inter8, gate193inter9, gate193inter10, gate193inter11, gate193inter12, gate147inter0, gate147inter1, gate147inter2, gate147inter3, gate147inter4, gate147inter5, gate147inter6, gate147inter7, gate147inter8, gate147inter9, gate147inter10, gate147inter11, gate147inter12, gate250inter0, gate250inter1, gate250inter2, gate250inter3, gate250inter4, gate250inter5, gate250inter6, gate250inter7, gate250inter8, gate250inter9, gate250inter10, gate250inter11, gate250inter12, gate189inter0, gate189inter1, gate189inter2, gate189inter3, gate189inter4, gate189inter5, gate189inter6, gate189inter7, gate189inter8, gate189inter9, gate189inter10, gate189inter11, gate189inter12, gate77inter0, gate77inter1, gate77inter2, gate77inter3, gate77inter4, gate77inter5, gate77inter6, gate77inter7, gate77inter8, gate77inter9, gate77inter10, gate77inter11, gate77inter12, gate176inter0, gate176inter1, gate176inter2, gate176inter3, gate176inter4, gate176inter5, gate176inter6, gate176inter7, gate176inter8, gate176inter9, gate176inter10, gate176inter11, gate176inter12, gate262inter0, gate262inter1, gate262inter2, gate262inter3, gate262inter4, gate262inter5, gate262inter6, gate262inter7, gate262inter8, gate262inter9, gate262inter10, gate262inter11, gate262inter12, gate215inter0, gate215inter1, gate215inter2, gate215inter3, gate215inter4, gate215inter5, gate215inter6, gate215inter7, gate215inter8, gate215inter9, gate215inter10, gate215inter11, gate215inter12, gate108inter0, gate108inter1, gate108inter2, gate108inter3, gate108inter4, gate108inter5, gate108inter6, gate108inter7, gate108inter8, gate108inter9, gate108inter10, gate108inter11, gate108inter12, gate54inter0, gate54inter1, gate54inter2, gate54inter3, gate54inter4, gate54inter5, gate54inter6, gate54inter7, gate54inter8, gate54inter9, gate54inter10, gate54inter11, gate54inter12, gate266inter0, gate266inter1, gate266inter2, gate266inter3, gate266inter4, gate266inter5, gate266inter6, gate266inter7, gate266inter8, gate266inter9, gate266inter10, gate266inter11, gate266inter12, gate150inter0, gate150inter1, gate150inter2, gate150inter3, gate150inter4, gate150inter5, gate150inter6, gate150inter7, gate150inter8, gate150inter9, gate150inter10, gate150inter11, gate150inter12, gate198inter0, gate198inter1, gate198inter2, gate198inter3, gate198inter4, gate198inter5, gate198inter6, gate198inter7, gate198inter8, gate198inter9, gate198inter10, gate198inter11, gate198inter12, gate91inter0, gate91inter1, gate91inter2, gate91inter3, gate91inter4, gate91inter5, gate91inter6, gate91inter7, gate91inter8, gate91inter9, gate91inter10, gate91inter11, gate91inter12, gate486inter0, gate486inter1, gate486inter2, gate486inter3, gate486inter4, gate486inter5, gate486inter6, gate486inter7, gate486inter8, gate486inter9, gate486inter10, gate486inter11, gate486inter12, gate39inter0, gate39inter1, gate39inter2, gate39inter3, gate39inter4, gate39inter5, gate39inter6, gate39inter7, gate39inter8, gate39inter9, gate39inter10, gate39inter11, gate39inter12, gate67inter0, gate67inter1, gate67inter2, gate67inter3, gate67inter4, gate67inter5, gate67inter6, gate67inter7, gate67inter8, gate67inter9, gate67inter10, gate67inter11, gate67inter12, gate68inter0, gate68inter1, gate68inter2, gate68inter3, gate68inter4, gate68inter5, gate68inter6, gate68inter7, gate68inter8, gate68inter9, gate68inter10, gate68inter11, gate68inter12, gate511inter0, gate511inter1, gate511inter2, gate511inter3, gate511inter4, gate511inter5, gate511inter6, gate511inter7, gate511inter8, gate511inter9, gate511inter10, gate511inter11, gate511inter12, gate269inter0, gate269inter1, gate269inter2, gate269inter3, gate269inter4, gate269inter5, gate269inter6, gate269inter7, gate269inter8, gate269inter9, gate269inter10, gate269inter11, gate269inter12, gate59inter0, gate59inter1, gate59inter2, gate59inter3, gate59inter4, gate59inter5, gate59inter6, gate59inter7, gate59inter8, gate59inter9, gate59inter10, gate59inter11, gate59inter12, gate506inter0, gate506inter1, gate506inter2, gate506inter3, gate506inter4, gate506inter5, gate506inter6, gate506inter7, gate506inter8, gate506inter9, gate506inter10, gate506inter11, gate506inter12, gate51inter0, gate51inter1, gate51inter2, gate51inter3, gate51inter4, gate51inter5, gate51inter6, gate51inter7, gate51inter8, gate51inter9, gate51inter10, gate51inter11, gate51inter12, gate472inter0, gate472inter1, gate472inter2, gate472inter3, gate472inter4, gate472inter5, gate472inter6, gate472inter7, gate472inter8, gate472inter9, gate472inter10, gate472inter11, gate472inter12, gate439inter0, gate439inter1, gate439inter2, gate439inter3, gate439inter4, gate439inter5, gate439inter6, gate439inter7, gate439inter8, gate439inter9, gate439inter10, gate439inter11, gate439inter12, gate279inter0, gate279inter1, gate279inter2, gate279inter3, gate279inter4, gate279inter5, gate279inter6, gate279inter7, gate279inter8, gate279inter9, gate279inter10, gate279inter11, gate279inter12, gate72inter0, gate72inter1, gate72inter2, gate72inter3, gate72inter4, gate72inter5, gate72inter6, gate72inter7, gate72inter8, gate72inter9, gate72inter10, gate72inter11, gate72inter12, gate125inter0, gate125inter1, gate125inter2, gate125inter3, gate125inter4, gate125inter5, gate125inter6, gate125inter7, gate125inter8, gate125inter9, gate125inter10, gate125inter11, gate125inter12, gate149inter0, gate149inter1, gate149inter2, gate149inter3, gate149inter4, gate149inter5, gate149inter6, gate149inter7, gate149inter8, gate149inter9, gate149inter10, gate149inter11, gate149inter12, gate430inter0, gate430inter1, gate430inter2, gate430inter3, gate430inter4, gate430inter5, gate430inter6, gate430inter7, gate430inter8, gate430inter9, gate430inter10, gate430inter11, gate430inter12, gate413inter0, gate413inter1, gate413inter2, gate413inter3, gate413inter4, gate413inter5, gate413inter6, gate413inter7, gate413inter8, gate413inter9, gate413inter10, gate413inter11, gate413inter12, gate491inter0, gate491inter1, gate491inter2, gate491inter3, gate491inter4, gate491inter5, gate491inter6, gate491inter7, gate491inter8, gate491inter9, gate491inter10, gate491inter11, gate491inter12, gate246inter0, gate246inter1, gate246inter2, gate246inter3, gate246inter4, gate246inter5, gate246inter6, gate246inter7, gate246inter8, gate246inter9, gate246inter10, gate246inter11, gate246inter12, gate207inter0, gate207inter1, gate207inter2, gate207inter3, gate207inter4, gate207inter5, gate207inter6, gate207inter7, gate207inter8, gate207inter9, gate207inter10, gate207inter11, gate207inter12, gate408inter0, gate408inter1, gate408inter2, gate408inter3, gate408inter4, gate408inter5, gate408inter6, gate408inter7, gate408inter8, gate408inter9, gate408inter10, gate408inter11, gate408inter12, gate22inter0, gate22inter1, gate22inter2, gate22inter3, gate22inter4, gate22inter5, gate22inter6, gate22inter7, gate22inter8, gate22inter9, gate22inter10, gate22inter11, gate22inter12, gate400inter0, gate400inter1, gate400inter2, gate400inter3, gate400inter4, gate400inter5, gate400inter6, gate400inter7, gate400inter8, gate400inter9, gate400inter10, gate400inter11, gate400inter12, gate220inter0, gate220inter1, gate220inter2, gate220inter3, gate220inter4, gate220inter5, gate220inter6, gate220inter7, gate220inter8, gate220inter9, gate220inter10, gate220inter11, gate220inter12, gate493inter0, gate493inter1, gate493inter2, gate493inter3, gate493inter4, gate493inter5, gate493inter6, gate493inter7, gate493inter8, gate493inter9, gate493inter10, gate493inter11, gate493inter12, gate105inter0, gate105inter1, gate105inter2, gate105inter3, gate105inter4, gate105inter5, gate105inter6, gate105inter7, gate105inter8, gate105inter9, gate105inter10, gate105inter11, gate105inter12, gate514inter0, gate514inter1, gate514inter2, gate514inter3, gate514inter4, gate514inter5, gate514inter6, gate514inter7, gate514inter8, gate514inter9, gate514inter10, gate514inter11, gate514inter12, gate206inter0, gate206inter1, gate206inter2, gate206inter3, gate206inter4, gate206inter5, gate206inter6, gate206inter7, gate206inter8, gate206inter9, gate206inter10, gate206inter11, gate206inter12, gate505inter0, gate505inter1, gate505inter2, gate505inter3, gate505inter4, gate505inter5, gate505inter6, gate505inter7, gate505inter8, gate505inter9, gate505inter10, gate505inter11, gate505inter12, gate243inter0, gate243inter1, gate243inter2, gate243inter3, gate243inter4, gate243inter5, gate243inter6, gate243inter7, gate243inter8, gate243inter9, gate243inter10, gate243inter11, gate243inter12, gate34inter0, gate34inter1, gate34inter2, gate34inter3, gate34inter4, gate34inter5, gate34inter6, gate34inter7, gate34inter8, gate34inter9, gate34inter10, gate34inter11, gate34inter12, gate64inter0, gate64inter1, gate64inter2, gate64inter3, gate64inter4, gate64inter5, gate64inter6, gate64inter7, gate64inter8, gate64inter9, gate64inter10, gate64inter11, gate64inter12, gate277inter0, gate277inter1, gate277inter2, gate277inter3, gate277inter4, gate277inter5, gate277inter6, gate277inter7, gate277inter8, gate277inter9, gate277inter10, gate277inter11, gate277inter12, gate172inter0, gate172inter1, gate172inter2, gate172inter3, gate172inter4, gate172inter5, gate172inter6, gate172inter7, gate172inter8, gate172inter9, gate172inter10, gate172inter11, gate172inter12, gate294inter0, gate294inter1, gate294inter2, gate294inter3, gate294inter4, gate294inter5, gate294inter6, gate294inter7, gate294inter8, gate294inter9, gate294inter10, gate294inter11, gate294inter12, gate100inter0, gate100inter1, gate100inter2, gate100inter3, gate100inter4, gate100inter5, gate100inter6, gate100inter7, gate100inter8, gate100inter9, gate100inter10, gate100inter11, gate100inter12, gate255inter0, gate255inter1, gate255inter2, gate255inter3, gate255inter4, gate255inter5, gate255inter6, gate255inter7, gate255inter8, gate255inter9, gate255inter10, gate255inter11, gate255inter12, gate396inter0, gate396inter1, gate396inter2, gate396inter3, gate396inter4, gate396inter5, gate396inter6, gate396inter7, gate396inter8, gate396inter9, gate396inter10, gate396inter11, gate396inter12, gate159inter0, gate159inter1, gate159inter2, gate159inter3, gate159inter4, gate159inter5, gate159inter6, gate159inter7, gate159inter8, gate159inter9, gate159inter10, gate159inter11, gate159inter12, gate140inter0, gate140inter1, gate140inter2, gate140inter3, gate140inter4, gate140inter5, gate140inter6, gate140inter7, gate140inter8, gate140inter9, gate140inter10, gate140inter11, gate140inter12, gate476inter0, gate476inter1, gate476inter2, gate476inter3, gate476inter4, gate476inter5, gate476inter6, gate476inter7, gate476inter8, gate476inter9, gate476inter10, gate476inter11, gate476inter12, gate393inter0, gate393inter1, gate393inter2, gate393inter3, gate393inter4, gate393inter5, gate393inter6, gate393inter7, gate393inter8, gate393inter9, gate393inter10, gate393inter11, gate393inter12, gate40inter0, gate40inter1, gate40inter2, gate40inter3, gate40inter4, gate40inter5, gate40inter6, gate40inter7, gate40inter8, gate40inter9, gate40inter10, gate40inter11, gate40inter12, gate475inter0, gate475inter1, gate475inter2, gate475inter3, gate475inter4, gate475inter5, gate475inter6, gate475inter7, gate475inter8, gate475inter9, gate475inter10, gate475inter11, gate475inter12, gate422inter0, gate422inter1, gate422inter2, gate422inter3, gate422inter4, gate422inter5, gate422inter6, gate422inter7, gate422inter8, gate422inter9, gate422inter10, gate422inter11, gate422inter12, gate163inter0, gate163inter1, gate163inter2, gate163inter3, gate163inter4, gate163inter5, gate163inter6, gate163inter7, gate163inter8, gate163inter9, gate163inter10, gate163inter11, gate163inter12, gate10inter0, gate10inter1, gate10inter2, gate10inter3, gate10inter4, gate10inter5, gate10inter6, gate10inter7, gate10inter8, gate10inter9, gate10inter10, gate10inter11, gate10inter12, gate221inter0, gate221inter1, gate221inter2, gate221inter3, gate221inter4, gate221inter5, gate221inter6, gate221inter7, gate221inter8, gate221inter9, gate221inter10, gate221inter11, gate221inter12, gate82inter0, gate82inter1, gate82inter2, gate82inter3, gate82inter4, gate82inter5, gate82inter6, gate82inter7, gate82inter8, gate82inter9, gate82inter10, gate82inter11, gate82inter12, gate416inter0, gate416inter1, gate416inter2, gate416inter3, gate416inter4, gate416inter5, gate416inter6, gate416inter7, gate416inter8, gate416inter9, gate416inter10, gate416inter11, gate416inter12, gate496inter0, gate496inter1, gate496inter2, gate496inter3, gate496inter4, gate496inter5, gate496inter6, gate496inter7, gate496inter8, gate496inter9, gate496inter10, gate496inter11, gate496inter12, gate477inter0, gate477inter1, gate477inter2, gate477inter3, gate477inter4, gate477inter5, gate477inter6, gate477inter7, gate477inter8, gate477inter9, gate477inter10, gate477inter11, gate477inter12, gate109inter0, gate109inter1, gate109inter2, gate109inter3, gate109inter4, gate109inter5, gate109inter6, gate109inter7, gate109inter8, gate109inter9, gate109inter10, gate109inter11, gate109inter12, gate99inter0, gate99inter1, gate99inter2, gate99inter3, gate99inter4, gate99inter5, gate99inter6, gate99inter7, gate99inter8, gate99inter9, gate99inter10, gate99inter11, gate99inter12, gate455inter0, gate455inter1, gate455inter2, gate455inter3, gate455inter4, gate455inter5, gate455inter6, gate455inter7, gate455inter8, gate455inter9, gate455inter10, gate455inter11, gate455inter12, gate418inter0, gate418inter1, gate418inter2, gate418inter3, gate418inter4, gate418inter5, gate418inter6, gate418inter7, gate418inter8, gate418inter9, gate418inter10, gate418inter11, gate418inter12, gate252inter0, gate252inter1, gate252inter2, gate252inter3, gate252inter4, gate252inter5, gate252inter6, gate252inter7, gate252inter8, gate252inter9, gate252inter10, gate252inter11, gate252inter12, gate201inter0, gate201inter1, gate201inter2, gate201inter3, gate201inter4, gate201inter5, gate201inter6, gate201inter7, gate201inter8, gate201inter9, gate201inter10, gate201inter11, gate201inter12, gate504inter0, gate504inter1, gate504inter2, gate504inter3, gate504inter4, gate504inter5, gate504inter6, gate504inter7, gate504inter8, gate504inter9, gate504inter10, gate504inter11, gate504inter12, gate397inter0, gate397inter1, gate397inter2, gate397inter3, gate397inter4, gate397inter5, gate397inter6, gate397inter7, gate397inter8, gate397inter9, gate397inter10, gate397inter11, gate397inter12, gate208inter0, gate208inter1, gate208inter2, gate208inter3, gate208inter4, gate208inter5, gate208inter6, gate208inter7, gate208inter8, gate208inter9, gate208inter10, gate208inter11, gate208inter12, gate293inter0, gate293inter1, gate293inter2, gate293inter3, gate293inter4, gate293inter5, gate293inter6, gate293inter7, gate293inter8, gate293inter9, gate293inter10, gate293inter11, gate293inter12, gate412inter0, gate412inter1, gate412inter2, gate412inter3, gate412inter4, gate412inter5, gate412inter6, gate412inter7, gate412inter8, gate412inter9, gate412inter10, gate412inter11, gate412inter12, gate211inter0, gate211inter1, gate211inter2, gate211inter3, gate211inter4, gate211inter5, gate211inter6, gate211inter7, gate211inter8, gate211inter9, gate211inter10, gate211inter11, gate211inter12, gate175inter0, gate175inter1, gate175inter2, gate175inter3, gate175inter4, gate175inter5, gate175inter6, gate175inter7, gate175inter8, gate175inter9, gate175inter10, gate175inter11, gate175inter12, gate165inter0, gate165inter1, gate165inter2, gate165inter3, gate165inter4, gate165inter5, gate165inter6, gate165inter7, gate165inter8, gate165inter9, gate165inter10, gate165inter11, gate165inter12, gate427inter0, gate427inter1, gate427inter2, gate427inter3, gate427inter4, gate427inter5, gate427inter6, gate427inter7, gate427inter8, gate427inter9, gate427inter10, gate427inter11, gate427inter12, gate459inter0, gate459inter1, gate459inter2, gate459inter3, gate459inter4, gate459inter5, gate459inter6, gate459inter7, gate459inter8, gate459inter9, gate459inter10, gate459inter11, gate459inter12, gate14inter0, gate14inter1, gate14inter2, gate14inter3, gate14inter4, gate14inter5, gate14inter6, gate14inter7, gate14inter8, gate14inter9, gate14inter10, gate14inter11, gate14inter12;



and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );
nand2 gate9( .a(G1), .b(G2), .O(G266) );

  xor2  gate1849(.a(G4), .b(G3), .O(gate10inter0));
  nand2 gate1850(.a(gate10inter0), .b(s_186), .O(gate10inter1));
  and2  gate1851(.a(G4), .b(G3), .O(gate10inter2));
  inv1  gate1852(.a(s_186), .O(gate10inter3));
  inv1  gate1853(.a(s_187), .O(gate10inter4));
  nand2 gate1854(.a(gate10inter4), .b(gate10inter3), .O(gate10inter5));
  nor2  gate1855(.a(gate10inter5), .b(gate10inter2), .O(gate10inter6));
  inv1  gate1856(.a(G3), .O(gate10inter7));
  inv1  gate1857(.a(G4), .O(gate10inter8));
  nand2 gate1858(.a(gate10inter8), .b(gate10inter7), .O(gate10inter9));
  nand2 gate1859(.a(s_187), .b(gate10inter3), .O(gate10inter10));
  nor2  gate1860(.a(gate10inter10), .b(gate10inter9), .O(gate10inter11));
  nor2  gate1861(.a(gate10inter11), .b(gate10inter6), .O(gate10inter12));
  nand2 gate1862(.a(gate10inter12), .b(gate10inter1), .O(G269));
nand2 gate11( .a(G5), .b(G6), .O(G272) );
nand2 gate12( .a(G7), .b(G8), .O(G275) );
nand2 gate13( .a(G9), .b(G10), .O(G278) );

  xor2  gate2157(.a(G12), .b(G11), .O(gate14inter0));
  nand2 gate2158(.a(gate14inter0), .b(s_230), .O(gate14inter1));
  and2  gate2159(.a(G12), .b(G11), .O(gate14inter2));
  inv1  gate2160(.a(s_230), .O(gate14inter3));
  inv1  gate2161(.a(s_231), .O(gate14inter4));
  nand2 gate2162(.a(gate14inter4), .b(gate14inter3), .O(gate14inter5));
  nor2  gate2163(.a(gate14inter5), .b(gate14inter2), .O(gate14inter6));
  inv1  gate2164(.a(G11), .O(gate14inter7));
  inv1  gate2165(.a(G12), .O(gate14inter8));
  nand2 gate2166(.a(gate14inter8), .b(gate14inter7), .O(gate14inter9));
  nand2 gate2167(.a(s_231), .b(gate14inter3), .O(gate14inter10));
  nor2  gate2168(.a(gate14inter10), .b(gate14inter9), .O(gate14inter11));
  nor2  gate2169(.a(gate14inter11), .b(gate14inter6), .O(gate14inter12));
  nand2 gate2170(.a(gate14inter12), .b(gate14inter1), .O(G281));
nand2 gate15( .a(G13), .b(G14), .O(G284) );
nand2 gate16( .a(G15), .b(G16), .O(G287) );
nand2 gate17( .a(G17), .b(G18), .O(G290) );
nand2 gate18( .a(G19), .b(G20), .O(G293) );

  xor2  gate967(.a(G22), .b(G21), .O(gate19inter0));
  nand2 gate968(.a(gate19inter0), .b(s_60), .O(gate19inter1));
  and2  gate969(.a(G22), .b(G21), .O(gate19inter2));
  inv1  gate970(.a(s_60), .O(gate19inter3));
  inv1  gate971(.a(s_61), .O(gate19inter4));
  nand2 gate972(.a(gate19inter4), .b(gate19inter3), .O(gate19inter5));
  nor2  gate973(.a(gate19inter5), .b(gate19inter2), .O(gate19inter6));
  inv1  gate974(.a(G21), .O(gate19inter7));
  inv1  gate975(.a(G22), .O(gate19inter8));
  nand2 gate976(.a(gate19inter8), .b(gate19inter7), .O(gate19inter9));
  nand2 gate977(.a(s_61), .b(gate19inter3), .O(gate19inter10));
  nor2  gate978(.a(gate19inter10), .b(gate19inter9), .O(gate19inter11));
  nor2  gate979(.a(gate19inter11), .b(gate19inter6), .O(gate19inter12));
  nand2 gate980(.a(gate19inter12), .b(gate19inter1), .O(G296));
nand2 gate20( .a(G23), .b(G24), .O(G299) );
nand2 gate21( .a(G25), .b(G26), .O(G302) );

  xor2  gate1499(.a(G28), .b(G27), .O(gate22inter0));
  nand2 gate1500(.a(gate22inter0), .b(s_136), .O(gate22inter1));
  and2  gate1501(.a(G28), .b(G27), .O(gate22inter2));
  inv1  gate1502(.a(s_136), .O(gate22inter3));
  inv1  gate1503(.a(s_137), .O(gate22inter4));
  nand2 gate1504(.a(gate22inter4), .b(gate22inter3), .O(gate22inter5));
  nor2  gate1505(.a(gate22inter5), .b(gate22inter2), .O(gate22inter6));
  inv1  gate1506(.a(G27), .O(gate22inter7));
  inv1  gate1507(.a(G28), .O(gate22inter8));
  nand2 gate1508(.a(gate22inter8), .b(gate22inter7), .O(gate22inter9));
  nand2 gate1509(.a(s_137), .b(gate22inter3), .O(gate22inter10));
  nor2  gate1510(.a(gate22inter10), .b(gate22inter9), .O(gate22inter11));
  nor2  gate1511(.a(gate22inter11), .b(gate22inter6), .O(gate22inter12));
  nand2 gate1512(.a(gate22inter12), .b(gate22inter1), .O(G305));
nand2 gate23( .a(G29), .b(G30), .O(G308) );
nand2 gate24( .a(G31), .b(G32), .O(G311) );
nand2 gate25( .a(G1), .b(G5), .O(G314) );
nand2 gate26( .a(G9), .b(G13), .O(G317) );
nand2 gate27( .a(G2), .b(G6), .O(G320) );
nand2 gate28( .a(G10), .b(G14), .O(G323) );

  xor2  gate981(.a(G7), .b(G3), .O(gate29inter0));
  nand2 gate982(.a(gate29inter0), .b(s_62), .O(gate29inter1));
  and2  gate983(.a(G7), .b(G3), .O(gate29inter2));
  inv1  gate984(.a(s_62), .O(gate29inter3));
  inv1  gate985(.a(s_63), .O(gate29inter4));
  nand2 gate986(.a(gate29inter4), .b(gate29inter3), .O(gate29inter5));
  nor2  gate987(.a(gate29inter5), .b(gate29inter2), .O(gate29inter6));
  inv1  gate988(.a(G3), .O(gate29inter7));
  inv1  gate989(.a(G7), .O(gate29inter8));
  nand2 gate990(.a(gate29inter8), .b(gate29inter7), .O(gate29inter9));
  nand2 gate991(.a(s_63), .b(gate29inter3), .O(gate29inter10));
  nor2  gate992(.a(gate29inter10), .b(gate29inter9), .O(gate29inter11));
  nor2  gate993(.a(gate29inter11), .b(gate29inter6), .O(gate29inter12));
  nand2 gate994(.a(gate29inter12), .b(gate29inter1), .O(G326));
nand2 gate30( .a(G11), .b(G15), .O(G329) );
nand2 gate31( .a(G4), .b(G8), .O(G332) );
nand2 gate32( .a(G12), .b(G16), .O(G335) );
nand2 gate33( .a(G17), .b(G21), .O(G338) );

  xor2  gate1625(.a(G29), .b(G25), .O(gate34inter0));
  nand2 gate1626(.a(gate34inter0), .b(s_154), .O(gate34inter1));
  and2  gate1627(.a(G29), .b(G25), .O(gate34inter2));
  inv1  gate1628(.a(s_154), .O(gate34inter3));
  inv1  gate1629(.a(s_155), .O(gate34inter4));
  nand2 gate1630(.a(gate34inter4), .b(gate34inter3), .O(gate34inter5));
  nor2  gate1631(.a(gate34inter5), .b(gate34inter2), .O(gate34inter6));
  inv1  gate1632(.a(G25), .O(gate34inter7));
  inv1  gate1633(.a(G29), .O(gate34inter8));
  nand2 gate1634(.a(gate34inter8), .b(gate34inter7), .O(gate34inter9));
  nand2 gate1635(.a(s_155), .b(gate34inter3), .O(gate34inter10));
  nor2  gate1636(.a(gate34inter10), .b(gate34inter9), .O(gate34inter11));
  nor2  gate1637(.a(gate34inter11), .b(gate34inter6), .O(gate34inter12));
  nand2 gate1638(.a(gate34inter12), .b(gate34inter1), .O(G341));
nand2 gate35( .a(G18), .b(G22), .O(G344) );
nand2 gate36( .a(G26), .b(G30), .O(G347) );
nand2 gate37( .a(G19), .b(G23), .O(G350) );
nand2 gate38( .a(G27), .b(G31), .O(G353) );

  xor2  gate1219(.a(G24), .b(G20), .O(gate39inter0));
  nand2 gate1220(.a(gate39inter0), .b(s_96), .O(gate39inter1));
  and2  gate1221(.a(G24), .b(G20), .O(gate39inter2));
  inv1  gate1222(.a(s_96), .O(gate39inter3));
  inv1  gate1223(.a(s_97), .O(gate39inter4));
  nand2 gate1224(.a(gate39inter4), .b(gate39inter3), .O(gate39inter5));
  nor2  gate1225(.a(gate39inter5), .b(gate39inter2), .O(gate39inter6));
  inv1  gate1226(.a(G20), .O(gate39inter7));
  inv1  gate1227(.a(G24), .O(gate39inter8));
  nand2 gate1228(.a(gate39inter8), .b(gate39inter7), .O(gate39inter9));
  nand2 gate1229(.a(s_97), .b(gate39inter3), .O(gate39inter10));
  nor2  gate1230(.a(gate39inter10), .b(gate39inter9), .O(gate39inter11));
  nor2  gate1231(.a(gate39inter11), .b(gate39inter6), .O(gate39inter12));
  nand2 gate1232(.a(gate39inter12), .b(gate39inter1), .O(G356));

  xor2  gate1793(.a(G32), .b(G28), .O(gate40inter0));
  nand2 gate1794(.a(gate40inter0), .b(s_178), .O(gate40inter1));
  and2  gate1795(.a(G32), .b(G28), .O(gate40inter2));
  inv1  gate1796(.a(s_178), .O(gate40inter3));
  inv1  gate1797(.a(s_179), .O(gate40inter4));
  nand2 gate1798(.a(gate40inter4), .b(gate40inter3), .O(gate40inter5));
  nor2  gate1799(.a(gate40inter5), .b(gate40inter2), .O(gate40inter6));
  inv1  gate1800(.a(G28), .O(gate40inter7));
  inv1  gate1801(.a(G32), .O(gate40inter8));
  nand2 gate1802(.a(gate40inter8), .b(gate40inter7), .O(gate40inter9));
  nand2 gate1803(.a(s_179), .b(gate40inter3), .O(gate40inter10));
  nor2  gate1804(.a(gate40inter10), .b(gate40inter9), .O(gate40inter11));
  nor2  gate1805(.a(gate40inter11), .b(gate40inter6), .O(gate40inter12));
  nand2 gate1806(.a(gate40inter12), .b(gate40inter1), .O(G359));
nand2 gate41( .a(G1), .b(G266), .O(G362) );
nand2 gate42( .a(G2), .b(G266), .O(G363) );
nand2 gate43( .a(G3), .b(G269), .O(G364) );
nand2 gate44( .a(G4), .b(G269), .O(G365) );
nand2 gate45( .a(G5), .b(G272), .O(G366) );
nand2 gate46( .a(G6), .b(G272), .O(G367) );
nand2 gate47( .a(G7), .b(G275), .O(G368) );
nand2 gate48( .a(G8), .b(G275), .O(G369) );
nand2 gate49( .a(G9), .b(G278), .O(G370) );
nand2 gate50( .a(G10), .b(G278), .O(G371) );

  xor2  gate1317(.a(G281), .b(G11), .O(gate51inter0));
  nand2 gate1318(.a(gate51inter0), .b(s_110), .O(gate51inter1));
  and2  gate1319(.a(G281), .b(G11), .O(gate51inter2));
  inv1  gate1320(.a(s_110), .O(gate51inter3));
  inv1  gate1321(.a(s_111), .O(gate51inter4));
  nand2 gate1322(.a(gate51inter4), .b(gate51inter3), .O(gate51inter5));
  nor2  gate1323(.a(gate51inter5), .b(gate51inter2), .O(gate51inter6));
  inv1  gate1324(.a(G11), .O(gate51inter7));
  inv1  gate1325(.a(G281), .O(gate51inter8));
  nand2 gate1326(.a(gate51inter8), .b(gate51inter7), .O(gate51inter9));
  nand2 gate1327(.a(s_111), .b(gate51inter3), .O(gate51inter10));
  nor2  gate1328(.a(gate51inter10), .b(gate51inter9), .O(gate51inter11));
  nor2  gate1329(.a(gate51inter11), .b(gate51inter6), .O(gate51inter12));
  nand2 gate1330(.a(gate51inter12), .b(gate51inter1), .O(G372));
nand2 gate52( .a(G12), .b(G281), .O(G373) );
nand2 gate53( .a(G13), .b(G284), .O(G374) );

  xor2  gate1135(.a(G284), .b(G14), .O(gate54inter0));
  nand2 gate1136(.a(gate54inter0), .b(s_84), .O(gate54inter1));
  and2  gate1137(.a(G284), .b(G14), .O(gate54inter2));
  inv1  gate1138(.a(s_84), .O(gate54inter3));
  inv1  gate1139(.a(s_85), .O(gate54inter4));
  nand2 gate1140(.a(gate54inter4), .b(gate54inter3), .O(gate54inter5));
  nor2  gate1141(.a(gate54inter5), .b(gate54inter2), .O(gate54inter6));
  inv1  gate1142(.a(G14), .O(gate54inter7));
  inv1  gate1143(.a(G284), .O(gate54inter8));
  nand2 gate1144(.a(gate54inter8), .b(gate54inter7), .O(gate54inter9));
  nand2 gate1145(.a(s_85), .b(gate54inter3), .O(gate54inter10));
  nor2  gate1146(.a(gate54inter10), .b(gate54inter9), .O(gate54inter11));
  nor2  gate1147(.a(gate54inter11), .b(gate54inter6), .O(gate54inter12));
  nand2 gate1148(.a(gate54inter12), .b(gate54inter1), .O(G375));
nand2 gate55( .a(G15), .b(G287), .O(G376) );
nand2 gate56( .a(G16), .b(G287), .O(G377) );
nand2 gate57( .a(G17), .b(G290), .O(G378) );
nand2 gate58( .a(G18), .b(G290), .O(G379) );

  xor2  gate1289(.a(G293), .b(G19), .O(gate59inter0));
  nand2 gate1290(.a(gate59inter0), .b(s_106), .O(gate59inter1));
  and2  gate1291(.a(G293), .b(G19), .O(gate59inter2));
  inv1  gate1292(.a(s_106), .O(gate59inter3));
  inv1  gate1293(.a(s_107), .O(gate59inter4));
  nand2 gate1294(.a(gate59inter4), .b(gate59inter3), .O(gate59inter5));
  nor2  gate1295(.a(gate59inter5), .b(gate59inter2), .O(gate59inter6));
  inv1  gate1296(.a(G19), .O(gate59inter7));
  inv1  gate1297(.a(G293), .O(gate59inter8));
  nand2 gate1298(.a(gate59inter8), .b(gate59inter7), .O(gate59inter9));
  nand2 gate1299(.a(s_107), .b(gate59inter3), .O(gate59inter10));
  nor2  gate1300(.a(gate59inter10), .b(gate59inter9), .O(gate59inter11));
  nor2  gate1301(.a(gate59inter11), .b(gate59inter6), .O(gate59inter12));
  nand2 gate1302(.a(gate59inter12), .b(gate59inter1), .O(G380));
nand2 gate60( .a(G20), .b(G293), .O(G381) );
nand2 gate61( .a(G21), .b(G296), .O(G382) );
nand2 gate62( .a(G22), .b(G296), .O(G383) );

  xor2  gate897(.a(G299), .b(G23), .O(gate63inter0));
  nand2 gate898(.a(gate63inter0), .b(s_50), .O(gate63inter1));
  and2  gate899(.a(G299), .b(G23), .O(gate63inter2));
  inv1  gate900(.a(s_50), .O(gate63inter3));
  inv1  gate901(.a(s_51), .O(gate63inter4));
  nand2 gate902(.a(gate63inter4), .b(gate63inter3), .O(gate63inter5));
  nor2  gate903(.a(gate63inter5), .b(gate63inter2), .O(gate63inter6));
  inv1  gate904(.a(G23), .O(gate63inter7));
  inv1  gate905(.a(G299), .O(gate63inter8));
  nand2 gate906(.a(gate63inter8), .b(gate63inter7), .O(gate63inter9));
  nand2 gate907(.a(s_51), .b(gate63inter3), .O(gate63inter10));
  nor2  gate908(.a(gate63inter10), .b(gate63inter9), .O(gate63inter11));
  nor2  gate909(.a(gate63inter11), .b(gate63inter6), .O(gate63inter12));
  nand2 gate910(.a(gate63inter12), .b(gate63inter1), .O(G384));

  xor2  gate1639(.a(G299), .b(G24), .O(gate64inter0));
  nand2 gate1640(.a(gate64inter0), .b(s_156), .O(gate64inter1));
  and2  gate1641(.a(G299), .b(G24), .O(gate64inter2));
  inv1  gate1642(.a(s_156), .O(gate64inter3));
  inv1  gate1643(.a(s_157), .O(gate64inter4));
  nand2 gate1644(.a(gate64inter4), .b(gate64inter3), .O(gate64inter5));
  nor2  gate1645(.a(gate64inter5), .b(gate64inter2), .O(gate64inter6));
  inv1  gate1646(.a(G24), .O(gate64inter7));
  inv1  gate1647(.a(G299), .O(gate64inter8));
  nand2 gate1648(.a(gate64inter8), .b(gate64inter7), .O(gate64inter9));
  nand2 gate1649(.a(s_157), .b(gate64inter3), .O(gate64inter10));
  nor2  gate1650(.a(gate64inter10), .b(gate64inter9), .O(gate64inter11));
  nor2  gate1651(.a(gate64inter11), .b(gate64inter6), .O(gate64inter12));
  nand2 gate1652(.a(gate64inter12), .b(gate64inter1), .O(G385));

  xor2  gate561(.a(G302), .b(G25), .O(gate65inter0));
  nand2 gate562(.a(gate65inter0), .b(s_2), .O(gate65inter1));
  and2  gate563(.a(G302), .b(G25), .O(gate65inter2));
  inv1  gate564(.a(s_2), .O(gate65inter3));
  inv1  gate565(.a(s_3), .O(gate65inter4));
  nand2 gate566(.a(gate65inter4), .b(gate65inter3), .O(gate65inter5));
  nor2  gate567(.a(gate65inter5), .b(gate65inter2), .O(gate65inter6));
  inv1  gate568(.a(G25), .O(gate65inter7));
  inv1  gate569(.a(G302), .O(gate65inter8));
  nand2 gate570(.a(gate65inter8), .b(gate65inter7), .O(gate65inter9));
  nand2 gate571(.a(s_3), .b(gate65inter3), .O(gate65inter10));
  nor2  gate572(.a(gate65inter10), .b(gate65inter9), .O(gate65inter11));
  nor2  gate573(.a(gate65inter11), .b(gate65inter6), .O(gate65inter12));
  nand2 gate574(.a(gate65inter12), .b(gate65inter1), .O(G386));
nand2 gate66( .a(G26), .b(G302), .O(G387) );

  xor2  gate1233(.a(G305), .b(G27), .O(gate67inter0));
  nand2 gate1234(.a(gate67inter0), .b(s_98), .O(gate67inter1));
  and2  gate1235(.a(G305), .b(G27), .O(gate67inter2));
  inv1  gate1236(.a(s_98), .O(gate67inter3));
  inv1  gate1237(.a(s_99), .O(gate67inter4));
  nand2 gate1238(.a(gate67inter4), .b(gate67inter3), .O(gate67inter5));
  nor2  gate1239(.a(gate67inter5), .b(gate67inter2), .O(gate67inter6));
  inv1  gate1240(.a(G27), .O(gate67inter7));
  inv1  gate1241(.a(G305), .O(gate67inter8));
  nand2 gate1242(.a(gate67inter8), .b(gate67inter7), .O(gate67inter9));
  nand2 gate1243(.a(s_99), .b(gate67inter3), .O(gate67inter10));
  nor2  gate1244(.a(gate67inter10), .b(gate67inter9), .O(gate67inter11));
  nor2  gate1245(.a(gate67inter11), .b(gate67inter6), .O(gate67inter12));
  nand2 gate1246(.a(gate67inter12), .b(gate67inter1), .O(G388));

  xor2  gate1247(.a(G305), .b(G28), .O(gate68inter0));
  nand2 gate1248(.a(gate68inter0), .b(s_100), .O(gate68inter1));
  and2  gate1249(.a(G305), .b(G28), .O(gate68inter2));
  inv1  gate1250(.a(s_100), .O(gate68inter3));
  inv1  gate1251(.a(s_101), .O(gate68inter4));
  nand2 gate1252(.a(gate68inter4), .b(gate68inter3), .O(gate68inter5));
  nor2  gate1253(.a(gate68inter5), .b(gate68inter2), .O(gate68inter6));
  inv1  gate1254(.a(G28), .O(gate68inter7));
  inv1  gate1255(.a(G305), .O(gate68inter8));
  nand2 gate1256(.a(gate68inter8), .b(gate68inter7), .O(gate68inter9));
  nand2 gate1257(.a(s_101), .b(gate68inter3), .O(gate68inter10));
  nor2  gate1258(.a(gate68inter10), .b(gate68inter9), .O(gate68inter11));
  nor2  gate1259(.a(gate68inter11), .b(gate68inter6), .O(gate68inter12));
  nand2 gate1260(.a(gate68inter12), .b(gate68inter1), .O(G389));
nand2 gate69( .a(G29), .b(G308), .O(G390) );
nand2 gate70( .a(G30), .b(G308), .O(G391) );
nand2 gate71( .a(G31), .b(G311), .O(G392) );

  xor2  gate1373(.a(G311), .b(G32), .O(gate72inter0));
  nand2 gate1374(.a(gate72inter0), .b(s_118), .O(gate72inter1));
  and2  gate1375(.a(G311), .b(G32), .O(gate72inter2));
  inv1  gate1376(.a(s_118), .O(gate72inter3));
  inv1  gate1377(.a(s_119), .O(gate72inter4));
  nand2 gate1378(.a(gate72inter4), .b(gate72inter3), .O(gate72inter5));
  nor2  gate1379(.a(gate72inter5), .b(gate72inter2), .O(gate72inter6));
  inv1  gate1380(.a(G32), .O(gate72inter7));
  inv1  gate1381(.a(G311), .O(gate72inter8));
  nand2 gate1382(.a(gate72inter8), .b(gate72inter7), .O(gate72inter9));
  nand2 gate1383(.a(s_119), .b(gate72inter3), .O(gate72inter10));
  nor2  gate1384(.a(gate72inter10), .b(gate72inter9), .O(gate72inter11));
  nor2  gate1385(.a(gate72inter11), .b(gate72inter6), .O(gate72inter12));
  nand2 gate1386(.a(gate72inter12), .b(gate72inter1), .O(G393));
nand2 gate73( .a(G1), .b(G314), .O(G394) );

  xor2  gate785(.a(G314), .b(G5), .O(gate74inter0));
  nand2 gate786(.a(gate74inter0), .b(s_34), .O(gate74inter1));
  and2  gate787(.a(G314), .b(G5), .O(gate74inter2));
  inv1  gate788(.a(s_34), .O(gate74inter3));
  inv1  gate789(.a(s_35), .O(gate74inter4));
  nand2 gate790(.a(gate74inter4), .b(gate74inter3), .O(gate74inter5));
  nor2  gate791(.a(gate74inter5), .b(gate74inter2), .O(gate74inter6));
  inv1  gate792(.a(G5), .O(gate74inter7));
  inv1  gate793(.a(G314), .O(gate74inter8));
  nand2 gate794(.a(gate74inter8), .b(gate74inter7), .O(gate74inter9));
  nand2 gate795(.a(s_35), .b(gate74inter3), .O(gate74inter10));
  nor2  gate796(.a(gate74inter10), .b(gate74inter9), .O(gate74inter11));
  nor2  gate797(.a(gate74inter11), .b(gate74inter6), .O(gate74inter12));
  nand2 gate798(.a(gate74inter12), .b(gate74inter1), .O(G395));
nand2 gate75( .a(G9), .b(G317), .O(G396) );
nand2 gate76( .a(G13), .b(G317), .O(G397) );

  xor2  gate1065(.a(G320), .b(G2), .O(gate77inter0));
  nand2 gate1066(.a(gate77inter0), .b(s_74), .O(gate77inter1));
  and2  gate1067(.a(G320), .b(G2), .O(gate77inter2));
  inv1  gate1068(.a(s_74), .O(gate77inter3));
  inv1  gate1069(.a(s_75), .O(gate77inter4));
  nand2 gate1070(.a(gate77inter4), .b(gate77inter3), .O(gate77inter5));
  nor2  gate1071(.a(gate77inter5), .b(gate77inter2), .O(gate77inter6));
  inv1  gate1072(.a(G2), .O(gate77inter7));
  inv1  gate1073(.a(G320), .O(gate77inter8));
  nand2 gate1074(.a(gate77inter8), .b(gate77inter7), .O(gate77inter9));
  nand2 gate1075(.a(s_75), .b(gate77inter3), .O(gate77inter10));
  nor2  gate1076(.a(gate77inter10), .b(gate77inter9), .O(gate77inter11));
  nor2  gate1077(.a(gate77inter11), .b(gate77inter6), .O(gate77inter12));
  nand2 gate1078(.a(gate77inter12), .b(gate77inter1), .O(G398));
nand2 gate78( .a(G6), .b(G320), .O(G399) );
nand2 gate79( .a(G10), .b(G323), .O(G400) );
nand2 gate80( .a(G14), .b(G323), .O(G401) );
nand2 gate81( .a(G3), .b(G326), .O(G402) );

  xor2  gate1877(.a(G326), .b(G7), .O(gate82inter0));
  nand2 gate1878(.a(gate82inter0), .b(s_190), .O(gate82inter1));
  and2  gate1879(.a(G326), .b(G7), .O(gate82inter2));
  inv1  gate1880(.a(s_190), .O(gate82inter3));
  inv1  gate1881(.a(s_191), .O(gate82inter4));
  nand2 gate1882(.a(gate82inter4), .b(gate82inter3), .O(gate82inter5));
  nor2  gate1883(.a(gate82inter5), .b(gate82inter2), .O(gate82inter6));
  inv1  gate1884(.a(G7), .O(gate82inter7));
  inv1  gate1885(.a(G326), .O(gate82inter8));
  nand2 gate1886(.a(gate82inter8), .b(gate82inter7), .O(gate82inter9));
  nand2 gate1887(.a(s_191), .b(gate82inter3), .O(gate82inter10));
  nor2  gate1888(.a(gate82inter10), .b(gate82inter9), .O(gate82inter11));
  nor2  gate1889(.a(gate82inter11), .b(gate82inter6), .O(gate82inter12));
  nand2 gate1890(.a(gate82inter12), .b(gate82inter1), .O(G403));
nand2 gate83( .a(G11), .b(G329), .O(G404) );
nand2 gate84( .a(G15), .b(G329), .O(G405) );
nand2 gate85( .a(G4), .b(G332), .O(G406) );
nand2 gate86( .a(G8), .b(G332), .O(G407) );
nand2 gate87( .a(G12), .b(G335), .O(G408) );
nand2 gate88( .a(G16), .b(G335), .O(G409) );
nand2 gate89( .a(G17), .b(G338), .O(G410) );
nand2 gate90( .a(G21), .b(G338), .O(G411) );

  xor2  gate1191(.a(G341), .b(G25), .O(gate91inter0));
  nand2 gate1192(.a(gate91inter0), .b(s_92), .O(gate91inter1));
  and2  gate1193(.a(G341), .b(G25), .O(gate91inter2));
  inv1  gate1194(.a(s_92), .O(gate91inter3));
  inv1  gate1195(.a(s_93), .O(gate91inter4));
  nand2 gate1196(.a(gate91inter4), .b(gate91inter3), .O(gate91inter5));
  nor2  gate1197(.a(gate91inter5), .b(gate91inter2), .O(gate91inter6));
  inv1  gate1198(.a(G25), .O(gate91inter7));
  inv1  gate1199(.a(G341), .O(gate91inter8));
  nand2 gate1200(.a(gate91inter8), .b(gate91inter7), .O(gate91inter9));
  nand2 gate1201(.a(s_93), .b(gate91inter3), .O(gate91inter10));
  nor2  gate1202(.a(gate91inter10), .b(gate91inter9), .O(gate91inter11));
  nor2  gate1203(.a(gate91inter11), .b(gate91inter6), .O(gate91inter12));
  nand2 gate1204(.a(gate91inter12), .b(gate91inter1), .O(G412));

  xor2  gate673(.a(G341), .b(G29), .O(gate92inter0));
  nand2 gate674(.a(gate92inter0), .b(s_18), .O(gate92inter1));
  and2  gate675(.a(G341), .b(G29), .O(gate92inter2));
  inv1  gate676(.a(s_18), .O(gate92inter3));
  inv1  gate677(.a(s_19), .O(gate92inter4));
  nand2 gate678(.a(gate92inter4), .b(gate92inter3), .O(gate92inter5));
  nor2  gate679(.a(gate92inter5), .b(gate92inter2), .O(gate92inter6));
  inv1  gate680(.a(G29), .O(gate92inter7));
  inv1  gate681(.a(G341), .O(gate92inter8));
  nand2 gate682(.a(gate92inter8), .b(gate92inter7), .O(gate92inter9));
  nand2 gate683(.a(s_19), .b(gate92inter3), .O(gate92inter10));
  nor2  gate684(.a(gate92inter10), .b(gate92inter9), .O(gate92inter11));
  nor2  gate685(.a(gate92inter11), .b(gate92inter6), .O(gate92inter12));
  nand2 gate686(.a(gate92inter12), .b(gate92inter1), .O(G413));
nand2 gate93( .a(G18), .b(G344), .O(G414) );

  xor2  gate995(.a(G344), .b(G22), .O(gate94inter0));
  nand2 gate996(.a(gate94inter0), .b(s_64), .O(gate94inter1));
  and2  gate997(.a(G344), .b(G22), .O(gate94inter2));
  inv1  gate998(.a(s_64), .O(gate94inter3));
  inv1  gate999(.a(s_65), .O(gate94inter4));
  nand2 gate1000(.a(gate94inter4), .b(gate94inter3), .O(gate94inter5));
  nor2  gate1001(.a(gate94inter5), .b(gate94inter2), .O(gate94inter6));
  inv1  gate1002(.a(G22), .O(gate94inter7));
  inv1  gate1003(.a(G344), .O(gate94inter8));
  nand2 gate1004(.a(gate94inter8), .b(gate94inter7), .O(gate94inter9));
  nand2 gate1005(.a(s_65), .b(gate94inter3), .O(gate94inter10));
  nor2  gate1006(.a(gate94inter10), .b(gate94inter9), .O(gate94inter11));
  nor2  gate1007(.a(gate94inter11), .b(gate94inter6), .O(gate94inter12));
  nand2 gate1008(.a(gate94inter12), .b(gate94inter1), .O(G415));
nand2 gate95( .a(G26), .b(G347), .O(G416) );
nand2 gate96( .a(G30), .b(G347), .O(G417) );

  xor2  gate841(.a(G350), .b(G19), .O(gate97inter0));
  nand2 gate842(.a(gate97inter0), .b(s_42), .O(gate97inter1));
  and2  gate843(.a(G350), .b(G19), .O(gate97inter2));
  inv1  gate844(.a(s_42), .O(gate97inter3));
  inv1  gate845(.a(s_43), .O(gate97inter4));
  nand2 gate846(.a(gate97inter4), .b(gate97inter3), .O(gate97inter5));
  nor2  gate847(.a(gate97inter5), .b(gate97inter2), .O(gate97inter6));
  inv1  gate848(.a(G19), .O(gate97inter7));
  inv1  gate849(.a(G350), .O(gate97inter8));
  nand2 gate850(.a(gate97inter8), .b(gate97inter7), .O(gate97inter9));
  nand2 gate851(.a(s_43), .b(gate97inter3), .O(gate97inter10));
  nor2  gate852(.a(gate97inter10), .b(gate97inter9), .O(gate97inter11));
  nor2  gate853(.a(gate97inter11), .b(gate97inter6), .O(gate97inter12));
  nand2 gate854(.a(gate97inter12), .b(gate97inter1), .O(G418));
nand2 gate98( .a(G23), .b(G350), .O(G419) );

  xor2  gate1947(.a(G353), .b(G27), .O(gate99inter0));
  nand2 gate1948(.a(gate99inter0), .b(s_200), .O(gate99inter1));
  and2  gate1949(.a(G353), .b(G27), .O(gate99inter2));
  inv1  gate1950(.a(s_200), .O(gate99inter3));
  inv1  gate1951(.a(s_201), .O(gate99inter4));
  nand2 gate1952(.a(gate99inter4), .b(gate99inter3), .O(gate99inter5));
  nor2  gate1953(.a(gate99inter5), .b(gate99inter2), .O(gate99inter6));
  inv1  gate1954(.a(G27), .O(gate99inter7));
  inv1  gate1955(.a(G353), .O(gate99inter8));
  nand2 gate1956(.a(gate99inter8), .b(gate99inter7), .O(gate99inter9));
  nand2 gate1957(.a(s_201), .b(gate99inter3), .O(gate99inter10));
  nor2  gate1958(.a(gate99inter10), .b(gate99inter9), .O(gate99inter11));
  nor2  gate1959(.a(gate99inter11), .b(gate99inter6), .O(gate99inter12));
  nand2 gate1960(.a(gate99inter12), .b(gate99inter1), .O(G420));

  xor2  gate1695(.a(G353), .b(G31), .O(gate100inter0));
  nand2 gate1696(.a(gate100inter0), .b(s_164), .O(gate100inter1));
  and2  gate1697(.a(G353), .b(G31), .O(gate100inter2));
  inv1  gate1698(.a(s_164), .O(gate100inter3));
  inv1  gate1699(.a(s_165), .O(gate100inter4));
  nand2 gate1700(.a(gate100inter4), .b(gate100inter3), .O(gate100inter5));
  nor2  gate1701(.a(gate100inter5), .b(gate100inter2), .O(gate100inter6));
  inv1  gate1702(.a(G31), .O(gate100inter7));
  inv1  gate1703(.a(G353), .O(gate100inter8));
  nand2 gate1704(.a(gate100inter8), .b(gate100inter7), .O(gate100inter9));
  nand2 gate1705(.a(s_165), .b(gate100inter3), .O(gate100inter10));
  nor2  gate1706(.a(gate100inter10), .b(gate100inter9), .O(gate100inter11));
  nor2  gate1707(.a(gate100inter11), .b(gate100inter6), .O(gate100inter12));
  nand2 gate1708(.a(gate100inter12), .b(gate100inter1), .O(G421));
nand2 gate101( .a(G20), .b(G356), .O(G422) );
nand2 gate102( .a(G24), .b(G356), .O(G423) );
nand2 gate103( .a(G28), .b(G359), .O(G424) );
nand2 gate104( .a(G32), .b(G359), .O(G425) );

  xor2  gate1555(.a(G363), .b(G362), .O(gate105inter0));
  nand2 gate1556(.a(gate105inter0), .b(s_144), .O(gate105inter1));
  and2  gate1557(.a(G363), .b(G362), .O(gate105inter2));
  inv1  gate1558(.a(s_144), .O(gate105inter3));
  inv1  gate1559(.a(s_145), .O(gate105inter4));
  nand2 gate1560(.a(gate105inter4), .b(gate105inter3), .O(gate105inter5));
  nor2  gate1561(.a(gate105inter5), .b(gate105inter2), .O(gate105inter6));
  inv1  gate1562(.a(G362), .O(gate105inter7));
  inv1  gate1563(.a(G363), .O(gate105inter8));
  nand2 gate1564(.a(gate105inter8), .b(gate105inter7), .O(gate105inter9));
  nand2 gate1565(.a(s_145), .b(gate105inter3), .O(gate105inter10));
  nor2  gate1566(.a(gate105inter10), .b(gate105inter9), .O(gate105inter11));
  nor2  gate1567(.a(gate105inter11), .b(gate105inter6), .O(gate105inter12));
  nand2 gate1568(.a(gate105inter12), .b(gate105inter1), .O(G426));
nand2 gate106( .a(G364), .b(G365), .O(G429) );
nand2 gate107( .a(G366), .b(G367), .O(G432) );

  xor2  gate1121(.a(G369), .b(G368), .O(gate108inter0));
  nand2 gate1122(.a(gate108inter0), .b(s_82), .O(gate108inter1));
  and2  gate1123(.a(G369), .b(G368), .O(gate108inter2));
  inv1  gate1124(.a(s_82), .O(gate108inter3));
  inv1  gate1125(.a(s_83), .O(gate108inter4));
  nand2 gate1126(.a(gate108inter4), .b(gate108inter3), .O(gate108inter5));
  nor2  gate1127(.a(gate108inter5), .b(gate108inter2), .O(gate108inter6));
  inv1  gate1128(.a(G368), .O(gate108inter7));
  inv1  gate1129(.a(G369), .O(gate108inter8));
  nand2 gate1130(.a(gate108inter8), .b(gate108inter7), .O(gate108inter9));
  nand2 gate1131(.a(s_83), .b(gate108inter3), .O(gate108inter10));
  nor2  gate1132(.a(gate108inter10), .b(gate108inter9), .O(gate108inter11));
  nor2  gate1133(.a(gate108inter11), .b(gate108inter6), .O(gate108inter12));
  nand2 gate1134(.a(gate108inter12), .b(gate108inter1), .O(G435));

  xor2  gate1933(.a(G371), .b(G370), .O(gate109inter0));
  nand2 gate1934(.a(gate109inter0), .b(s_198), .O(gate109inter1));
  and2  gate1935(.a(G371), .b(G370), .O(gate109inter2));
  inv1  gate1936(.a(s_198), .O(gate109inter3));
  inv1  gate1937(.a(s_199), .O(gate109inter4));
  nand2 gate1938(.a(gate109inter4), .b(gate109inter3), .O(gate109inter5));
  nor2  gate1939(.a(gate109inter5), .b(gate109inter2), .O(gate109inter6));
  inv1  gate1940(.a(G370), .O(gate109inter7));
  inv1  gate1941(.a(G371), .O(gate109inter8));
  nand2 gate1942(.a(gate109inter8), .b(gate109inter7), .O(gate109inter9));
  nand2 gate1943(.a(s_199), .b(gate109inter3), .O(gate109inter10));
  nor2  gate1944(.a(gate109inter10), .b(gate109inter9), .O(gate109inter11));
  nor2  gate1945(.a(gate109inter11), .b(gate109inter6), .O(gate109inter12));
  nand2 gate1946(.a(gate109inter12), .b(gate109inter1), .O(G438));
nand2 gate110( .a(G372), .b(G373), .O(G441) );
nand2 gate111( .a(G374), .b(G375), .O(G444) );
nand2 gate112( .a(G376), .b(G377), .O(G447) );
nand2 gate113( .a(G378), .b(G379), .O(G450) );
nand2 gate114( .a(G380), .b(G381), .O(G453) );
nand2 gate115( .a(G382), .b(G383), .O(G456) );
nand2 gate116( .a(G384), .b(G385), .O(G459) );
nand2 gate117( .a(G386), .b(G387), .O(G462) );
nand2 gate118( .a(G388), .b(G389), .O(G465) );
nand2 gate119( .a(G390), .b(G391), .O(G468) );
nand2 gate120( .a(G392), .b(G393), .O(G471) );
nand2 gate121( .a(G394), .b(G395), .O(G474) );
nand2 gate122( .a(G396), .b(G397), .O(G477) );

  xor2  gate799(.a(G399), .b(G398), .O(gate123inter0));
  nand2 gate800(.a(gate123inter0), .b(s_36), .O(gate123inter1));
  and2  gate801(.a(G399), .b(G398), .O(gate123inter2));
  inv1  gate802(.a(s_36), .O(gate123inter3));
  inv1  gate803(.a(s_37), .O(gate123inter4));
  nand2 gate804(.a(gate123inter4), .b(gate123inter3), .O(gate123inter5));
  nor2  gate805(.a(gate123inter5), .b(gate123inter2), .O(gate123inter6));
  inv1  gate806(.a(G398), .O(gate123inter7));
  inv1  gate807(.a(G399), .O(gate123inter8));
  nand2 gate808(.a(gate123inter8), .b(gate123inter7), .O(gate123inter9));
  nand2 gate809(.a(s_37), .b(gate123inter3), .O(gate123inter10));
  nor2  gate810(.a(gate123inter10), .b(gate123inter9), .O(gate123inter11));
  nor2  gate811(.a(gate123inter11), .b(gate123inter6), .O(gate123inter12));
  nand2 gate812(.a(gate123inter12), .b(gate123inter1), .O(G480));
nand2 gate124( .a(G400), .b(G401), .O(G483) );

  xor2  gate1387(.a(G403), .b(G402), .O(gate125inter0));
  nand2 gate1388(.a(gate125inter0), .b(s_120), .O(gate125inter1));
  and2  gate1389(.a(G403), .b(G402), .O(gate125inter2));
  inv1  gate1390(.a(s_120), .O(gate125inter3));
  inv1  gate1391(.a(s_121), .O(gate125inter4));
  nand2 gate1392(.a(gate125inter4), .b(gate125inter3), .O(gate125inter5));
  nor2  gate1393(.a(gate125inter5), .b(gate125inter2), .O(gate125inter6));
  inv1  gate1394(.a(G402), .O(gate125inter7));
  inv1  gate1395(.a(G403), .O(gate125inter8));
  nand2 gate1396(.a(gate125inter8), .b(gate125inter7), .O(gate125inter9));
  nand2 gate1397(.a(s_121), .b(gate125inter3), .O(gate125inter10));
  nor2  gate1398(.a(gate125inter10), .b(gate125inter9), .O(gate125inter11));
  nor2  gate1399(.a(gate125inter11), .b(gate125inter6), .O(gate125inter12));
  nand2 gate1400(.a(gate125inter12), .b(gate125inter1), .O(G486));
nand2 gate126( .a(G404), .b(G405), .O(G489) );
nand2 gate127( .a(G406), .b(G407), .O(G492) );

  xor2  gate869(.a(G409), .b(G408), .O(gate128inter0));
  nand2 gate870(.a(gate128inter0), .b(s_46), .O(gate128inter1));
  and2  gate871(.a(G409), .b(G408), .O(gate128inter2));
  inv1  gate872(.a(s_46), .O(gate128inter3));
  inv1  gate873(.a(s_47), .O(gate128inter4));
  nand2 gate874(.a(gate128inter4), .b(gate128inter3), .O(gate128inter5));
  nor2  gate875(.a(gate128inter5), .b(gate128inter2), .O(gate128inter6));
  inv1  gate876(.a(G408), .O(gate128inter7));
  inv1  gate877(.a(G409), .O(gate128inter8));
  nand2 gate878(.a(gate128inter8), .b(gate128inter7), .O(gate128inter9));
  nand2 gate879(.a(s_47), .b(gate128inter3), .O(gate128inter10));
  nor2  gate880(.a(gate128inter10), .b(gate128inter9), .O(gate128inter11));
  nor2  gate881(.a(gate128inter11), .b(gate128inter6), .O(gate128inter12));
  nand2 gate882(.a(gate128inter12), .b(gate128inter1), .O(G495));
nand2 gate129( .a(G410), .b(G411), .O(G498) );
nand2 gate130( .a(G412), .b(G413), .O(G501) );
nand2 gate131( .a(G414), .b(G415), .O(G504) );
nand2 gate132( .a(G416), .b(G417), .O(G507) );
nand2 gate133( .a(G418), .b(G419), .O(G510) );
nand2 gate134( .a(G420), .b(G421), .O(G513) );
nand2 gate135( .a(G422), .b(G423), .O(G516) );
nand2 gate136( .a(G424), .b(G425), .O(G519) );
nand2 gate137( .a(G426), .b(G429), .O(G522) );
nand2 gate138( .a(G432), .b(G435), .O(G525) );
nand2 gate139( .a(G438), .b(G441), .O(G528) );

  xor2  gate1751(.a(G447), .b(G444), .O(gate140inter0));
  nand2 gate1752(.a(gate140inter0), .b(s_172), .O(gate140inter1));
  and2  gate1753(.a(G447), .b(G444), .O(gate140inter2));
  inv1  gate1754(.a(s_172), .O(gate140inter3));
  inv1  gate1755(.a(s_173), .O(gate140inter4));
  nand2 gate1756(.a(gate140inter4), .b(gate140inter3), .O(gate140inter5));
  nor2  gate1757(.a(gate140inter5), .b(gate140inter2), .O(gate140inter6));
  inv1  gate1758(.a(G444), .O(gate140inter7));
  inv1  gate1759(.a(G447), .O(gate140inter8));
  nand2 gate1760(.a(gate140inter8), .b(gate140inter7), .O(gate140inter9));
  nand2 gate1761(.a(s_173), .b(gate140inter3), .O(gate140inter10));
  nor2  gate1762(.a(gate140inter10), .b(gate140inter9), .O(gate140inter11));
  nor2  gate1763(.a(gate140inter11), .b(gate140inter6), .O(gate140inter12));
  nand2 gate1764(.a(gate140inter12), .b(gate140inter1), .O(G531));
nand2 gate141( .a(G450), .b(G453), .O(G534) );
nand2 gate142( .a(G456), .b(G459), .O(G537) );
nand2 gate143( .a(G462), .b(G465), .O(G540) );
nand2 gate144( .a(G468), .b(G471), .O(G543) );
nand2 gate145( .a(G474), .b(G477), .O(G546) );
nand2 gate146( .a(G480), .b(G483), .O(G549) );

  xor2  gate1023(.a(G489), .b(G486), .O(gate147inter0));
  nand2 gate1024(.a(gate147inter0), .b(s_68), .O(gate147inter1));
  and2  gate1025(.a(G489), .b(G486), .O(gate147inter2));
  inv1  gate1026(.a(s_68), .O(gate147inter3));
  inv1  gate1027(.a(s_69), .O(gate147inter4));
  nand2 gate1028(.a(gate147inter4), .b(gate147inter3), .O(gate147inter5));
  nor2  gate1029(.a(gate147inter5), .b(gate147inter2), .O(gate147inter6));
  inv1  gate1030(.a(G486), .O(gate147inter7));
  inv1  gate1031(.a(G489), .O(gate147inter8));
  nand2 gate1032(.a(gate147inter8), .b(gate147inter7), .O(gate147inter9));
  nand2 gate1033(.a(s_69), .b(gate147inter3), .O(gate147inter10));
  nor2  gate1034(.a(gate147inter10), .b(gate147inter9), .O(gate147inter11));
  nor2  gate1035(.a(gate147inter11), .b(gate147inter6), .O(gate147inter12));
  nand2 gate1036(.a(gate147inter12), .b(gate147inter1), .O(G552));
nand2 gate148( .a(G492), .b(G495), .O(G555) );

  xor2  gate1401(.a(G501), .b(G498), .O(gate149inter0));
  nand2 gate1402(.a(gate149inter0), .b(s_122), .O(gate149inter1));
  and2  gate1403(.a(G501), .b(G498), .O(gate149inter2));
  inv1  gate1404(.a(s_122), .O(gate149inter3));
  inv1  gate1405(.a(s_123), .O(gate149inter4));
  nand2 gate1406(.a(gate149inter4), .b(gate149inter3), .O(gate149inter5));
  nor2  gate1407(.a(gate149inter5), .b(gate149inter2), .O(gate149inter6));
  inv1  gate1408(.a(G498), .O(gate149inter7));
  inv1  gate1409(.a(G501), .O(gate149inter8));
  nand2 gate1410(.a(gate149inter8), .b(gate149inter7), .O(gate149inter9));
  nand2 gate1411(.a(s_123), .b(gate149inter3), .O(gate149inter10));
  nor2  gate1412(.a(gate149inter10), .b(gate149inter9), .O(gate149inter11));
  nor2  gate1413(.a(gate149inter11), .b(gate149inter6), .O(gate149inter12));
  nand2 gate1414(.a(gate149inter12), .b(gate149inter1), .O(G558));

  xor2  gate1163(.a(G507), .b(G504), .O(gate150inter0));
  nand2 gate1164(.a(gate150inter0), .b(s_88), .O(gate150inter1));
  and2  gate1165(.a(G507), .b(G504), .O(gate150inter2));
  inv1  gate1166(.a(s_88), .O(gate150inter3));
  inv1  gate1167(.a(s_89), .O(gate150inter4));
  nand2 gate1168(.a(gate150inter4), .b(gate150inter3), .O(gate150inter5));
  nor2  gate1169(.a(gate150inter5), .b(gate150inter2), .O(gate150inter6));
  inv1  gate1170(.a(G504), .O(gate150inter7));
  inv1  gate1171(.a(G507), .O(gate150inter8));
  nand2 gate1172(.a(gate150inter8), .b(gate150inter7), .O(gate150inter9));
  nand2 gate1173(.a(s_89), .b(gate150inter3), .O(gate150inter10));
  nor2  gate1174(.a(gate150inter10), .b(gate150inter9), .O(gate150inter11));
  nor2  gate1175(.a(gate150inter11), .b(gate150inter6), .O(gate150inter12));
  nand2 gate1176(.a(gate150inter12), .b(gate150inter1), .O(G561));
nand2 gate151( .a(G510), .b(G513), .O(G564) );
nand2 gate152( .a(G516), .b(G519), .O(G567) );

  xor2  gate687(.a(G522), .b(G426), .O(gate153inter0));
  nand2 gate688(.a(gate153inter0), .b(s_20), .O(gate153inter1));
  and2  gate689(.a(G522), .b(G426), .O(gate153inter2));
  inv1  gate690(.a(s_20), .O(gate153inter3));
  inv1  gate691(.a(s_21), .O(gate153inter4));
  nand2 gate692(.a(gate153inter4), .b(gate153inter3), .O(gate153inter5));
  nor2  gate693(.a(gate153inter5), .b(gate153inter2), .O(gate153inter6));
  inv1  gate694(.a(G426), .O(gate153inter7));
  inv1  gate695(.a(G522), .O(gate153inter8));
  nand2 gate696(.a(gate153inter8), .b(gate153inter7), .O(gate153inter9));
  nand2 gate697(.a(s_21), .b(gate153inter3), .O(gate153inter10));
  nor2  gate698(.a(gate153inter10), .b(gate153inter9), .O(gate153inter11));
  nor2  gate699(.a(gate153inter11), .b(gate153inter6), .O(gate153inter12));
  nand2 gate700(.a(gate153inter12), .b(gate153inter1), .O(G570));
nand2 gate154( .a(G429), .b(G522), .O(G571) );
nand2 gate155( .a(G432), .b(G525), .O(G572) );
nand2 gate156( .a(G435), .b(G525), .O(G573) );

  xor2  gate659(.a(G528), .b(G438), .O(gate157inter0));
  nand2 gate660(.a(gate157inter0), .b(s_16), .O(gate157inter1));
  and2  gate661(.a(G528), .b(G438), .O(gate157inter2));
  inv1  gate662(.a(s_16), .O(gate157inter3));
  inv1  gate663(.a(s_17), .O(gate157inter4));
  nand2 gate664(.a(gate157inter4), .b(gate157inter3), .O(gate157inter5));
  nor2  gate665(.a(gate157inter5), .b(gate157inter2), .O(gate157inter6));
  inv1  gate666(.a(G438), .O(gate157inter7));
  inv1  gate667(.a(G528), .O(gate157inter8));
  nand2 gate668(.a(gate157inter8), .b(gate157inter7), .O(gate157inter9));
  nand2 gate669(.a(s_17), .b(gate157inter3), .O(gate157inter10));
  nor2  gate670(.a(gate157inter10), .b(gate157inter9), .O(gate157inter11));
  nor2  gate671(.a(gate157inter11), .b(gate157inter6), .O(gate157inter12));
  nand2 gate672(.a(gate157inter12), .b(gate157inter1), .O(G574));
nand2 gate158( .a(G441), .b(G528), .O(G575) );

  xor2  gate1737(.a(G531), .b(G444), .O(gate159inter0));
  nand2 gate1738(.a(gate159inter0), .b(s_170), .O(gate159inter1));
  and2  gate1739(.a(G531), .b(G444), .O(gate159inter2));
  inv1  gate1740(.a(s_170), .O(gate159inter3));
  inv1  gate1741(.a(s_171), .O(gate159inter4));
  nand2 gate1742(.a(gate159inter4), .b(gate159inter3), .O(gate159inter5));
  nor2  gate1743(.a(gate159inter5), .b(gate159inter2), .O(gate159inter6));
  inv1  gate1744(.a(G444), .O(gate159inter7));
  inv1  gate1745(.a(G531), .O(gate159inter8));
  nand2 gate1746(.a(gate159inter8), .b(gate159inter7), .O(gate159inter9));
  nand2 gate1747(.a(s_171), .b(gate159inter3), .O(gate159inter10));
  nor2  gate1748(.a(gate159inter10), .b(gate159inter9), .O(gate159inter11));
  nor2  gate1749(.a(gate159inter11), .b(gate159inter6), .O(gate159inter12));
  nand2 gate1750(.a(gate159inter12), .b(gate159inter1), .O(G576));
nand2 gate160( .a(G447), .b(G531), .O(G577) );
nand2 gate161( .a(G450), .b(G534), .O(G578) );
nand2 gate162( .a(G453), .b(G534), .O(G579) );

  xor2  gate1835(.a(G537), .b(G456), .O(gate163inter0));
  nand2 gate1836(.a(gate163inter0), .b(s_184), .O(gate163inter1));
  and2  gate1837(.a(G537), .b(G456), .O(gate163inter2));
  inv1  gate1838(.a(s_184), .O(gate163inter3));
  inv1  gate1839(.a(s_185), .O(gate163inter4));
  nand2 gate1840(.a(gate163inter4), .b(gate163inter3), .O(gate163inter5));
  nor2  gate1841(.a(gate163inter5), .b(gate163inter2), .O(gate163inter6));
  inv1  gate1842(.a(G456), .O(gate163inter7));
  inv1  gate1843(.a(G537), .O(gate163inter8));
  nand2 gate1844(.a(gate163inter8), .b(gate163inter7), .O(gate163inter9));
  nand2 gate1845(.a(s_185), .b(gate163inter3), .O(gate163inter10));
  nor2  gate1846(.a(gate163inter10), .b(gate163inter9), .O(gate163inter11));
  nor2  gate1847(.a(gate163inter11), .b(gate163inter6), .O(gate163inter12));
  nand2 gate1848(.a(gate163inter12), .b(gate163inter1), .O(G580));
nand2 gate164( .a(G459), .b(G537), .O(G581) );

  xor2  gate2115(.a(G540), .b(G462), .O(gate165inter0));
  nand2 gate2116(.a(gate165inter0), .b(s_224), .O(gate165inter1));
  and2  gate2117(.a(G540), .b(G462), .O(gate165inter2));
  inv1  gate2118(.a(s_224), .O(gate165inter3));
  inv1  gate2119(.a(s_225), .O(gate165inter4));
  nand2 gate2120(.a(gate165inter4), .b(gate165inter3), .O(gate165inter5));
  nor2  gate2121(.a(gate165inter5), .b(gate165inter2), .O(gate165inter6));
  inv1  gate2122(.a(G462), .O(gate165inter7));
  inv1  gate2123(.a(G540), .O(gate165inter8));
  nand2 gate2124(.a(gate165inter8), .b(gate165inter7), .O(gate165inter9));
  nand2 gate2125(.a(s_225), .b(gate165inter3), .O(gate165inter10));
  nor2  gate2126(.a(gate165inter10), .b(gate165inter9), .O(gate165inter11));
  nor2  gate2127(.a(gate165inter11), .b(gate165inter6), .O(gate165inter12));
  nand2 gate2128(.a(gate165inter12), .b(gate165inter1), .O(G582));
nand2 gate166( .a(G465), .b(G540), .O(G583) );
nand2 gate167( .a(G468), .b(G543), .O(G584) );
nand2 gate168( .a(G471), .b(G543), .O(G585) );
nand2 gate169( .a(G474), .b(G546), .O(G586) );
nand2 gate170( .a(G477), .b(G546), .O(G587) );
nand2 gate171( .a(G480), .b(G549), .O(G588) );

  xor2  gate1667(.a(G549), .b(G483), .O(gate172inter0));
  nand2 gate1668(.a(gate172inter0), .b(s_160), .O(gate172inter1));
  and2  gate1669(.a(G549), .b(G483), .O(gate172inter2));
  inv1  gate1670(.a(s_160), .O(gate172inter3));
  inv1  gate1671(.a(s_161), .O(gate172inter4));
  nand2 gate1672(.a(gate172inter4), .b(gate172inter3), .O(gate172inter5));
  nor2  gate1673(.a(gate172inter5), .b(gate172inter2), .O(gate172inter6));
  inv1  gate1674(.a(G483), .O(gate172inter7));
  inv1  gate1675(.a(G549), .O(gate172inter8));
  nand2 gate1676(.a(gate172inter8), .b(gate172inter7), .O(gate172inter9));
  nand2 gate1677(.a(s_161), .b(gate172inter3), .O(gate172inter10));
  nor2  gate1678(.a(gate172inter10), .b(gate172inter9), .O(gate172inter11));
  nor2  gate1679(.a(gate172inter11), .b(gate172inter6), .O(gate172inter12));
  nand2 gate1680(.a(gate172inter12), .b(gate172inter1), .O(G589));
nand2 gate173( .a(G486), .b(G552), .O(G590) );
nand2 gate174( .a(G489), .b(G552), .O(G591) );

  xor2  gate2101(.a(G555), .b(G492), .O(gate175inter0));
  nand2 gate2102(.a(gate175inter0), .b(s_222), .O(gate175inter1));
  and2  gate2103(.a(G555), .b(G492), .O(gate175inter2));
  inv1  gate2104(.a(s_222), .O(gate175inter3));
  inv1  gate2105(.a(s_223), .O(gate175inter4));
  nand2 gate2106(.a(gate175inter4), .b(gate175inter3), .O(gate175inter5));
  nor2  gate2107(.a(gate175inter5), .b(gate175inter2), .O(gate175inter6));
  inv1  gate2108(.a(G492), .O(gate175inter7));
  inv1  gate2109(.a(G555), .O(gate175inter8));
  nand2 gate2110(.a(gate175inter8), .b(gate175inter7), .O(gate175inter9));
  nand2 gate2111(.a(s_223), .b(gate175inter3), .O(gate175inter10));
  nor2  gate2112(.a(gate175inter10), .b(gate175inter9), .O(gate175inter11));
  nor2  gate2113(.a(gate175inter11), .b(gate175inter6), .O(gate175inter12));
  nand2 gate2114(.a(gate175inter12), .b(gate175inter1), .O(G592));

  xor2  gate1079(.a(G555), .b(G495), .O(gate176inter0));
  nand2 gate1080(.a(gate176inter0), .b(s_76), .O(gate176inter1));
  and2  gate1081(.a(G555), .b(G495), .O(gate176inter2));
  inv1  gate1082(.a(s_76), .O(gate176inter3));
  inv1  gate1083(.a(s_77), .O(gate176inter4));
  nand2 gate1084(.a(gate176inter4), .b(gate176inter3), .O(gate176inter5));
  nor2  gate1085(.a(gate176inter5), .b(gate176inter2), .O(gate176inter6));
  inv1  gate1086(.a(G495), .O(gate176inter7));
  inv1  gate1087(.a(G555), .O(gate176inter8));
  nand2 gate1088(.a(gate176inter8), .b(gate176inter7), .O(gate176inter9));
  nand2 gate1089(.a(s_77), .b(gate176inter3), .O(gate176inter10));
  nor2  gate1090(.a(gate176inter10), .b(gate176inter9), .O(gate176inter11));
  nor2  gate1091(.a(gate176inter11), .b(gate176inter6), .O(gate176inter12));
  nand2 gate1092(.a(gate176inter12), .b(gate176inter1), .O(G593));
nand2 gate177( .a(G498), .b(G558), .O(G594) );
nand2 gate178( .a(G501), .b(G558), .O(G595) );
nand2 gate179( .a(G504), .b(G561), .O(G596) );
nand2 gate180( .a(G507), .b(G561), .O(G597) );
nand2 gate181( .a(G510), .b(G564), .O(G598) );
nand2 gate182( .a(G513), .b(G564), .O(G599) );
nand2 gate183( .a(G516), .b(G567), .O(G600) );
nand2 gate184( .a(G519), .b(G567), .O(G601) );
nand2 gate185( .a(G570), .b(G571), .O(G602) );
nand2 gate186( .a(G572), .b(G573), .O(G607) );
nand2 gate187( .a(G574), .b(G575), .O(G612) );
nand2 gate188( .a(G576), .b(G577), .O(G617) );

  xor2  gate1051(.a(G579), .b(G578), .O(gate189inter0));
  nand2 gate1052(.a(gate189inter0), .b(s_72), .O(gate189inter1));
  and2  gate1053(.a(G579), .b(G578), .O(gate189inter2));
  inv1  gate1054(.a(s_72), .O(gate189inter3));
  inv1  gate1055(.a(s_73), .O(gate189inter4));
  nand2 gate1056(.a(gate189inter4), .b(gate189inter3), .O(gate189inter5));
  nor2  gate1057(.a(gate189inter5), .b(gate189inter2), .O(gate189inter6));
  inv1  gate1058(.a(G578), .O(gate189inter7));
  inv1  gate1059(.a(G579), .O(gate189inter8));
  nand2 gate1060(.a(gate189inter8), .b(gate189inter7), .O(gate189inter9));
  nand2 gate1061(.a(s_73), .b(gate189inter3), .O(gate189inter10));
  nor2  gate1062(.a(gate189inter10), .b(gate189inter9), .O(gate189inter11));
  nor2  gate1063(.a(gate189inter11), .b(gate189inter6), .O(gate189inter12));
  nand2 gate1064(.a(gate189inter12), .b(gate189inter1), .O(G622));
nand2 gate190( .a(G580), .b(G581), .O(G627) );
nand2 gate191( .a(G582), .b(G583), .O(G632) );
nand2 gate192( .a(G584), .b(G585), .O(G637) );

  xor2  gate1009(.a(G587), .b(G586), .O(gate193inter0));
  nand2 gate1010(.a(gate193inter0), .b(s_66), .O(gate193inter1));
  and2  gate1011(.a(G587), .b(G586), .O(gate193inter2));
  inv1  gate1012(.a(s_66), .O(gate193inter3));
  inv1  gate1013(.a(s_67), .O(gate193inter4));
  nand2 gate1014(.a(gate193inter4), .b(gate193inter3), .O(gate193inter5));
  nor2  gate1015(.a(gate193inter5), .b(gate193inter2), .O(gate193inter6));
  inv1  gate1016(.a(G586), .O(gate193inter7));
  inv1  gate1017(.a(G587), .O(gate193inter8));
  nand2 gate1018(.a(gate193inter8), .b(gate193inter7), .O(gate193inter9));
  nand2 gate1019(.a(s_67), .b(gate193inter3), .O(gate193inter10));
  nor2  gate1020(.a(gate193inter10), .b(gate193inter9), .O(gate193inter11));
  nor2  gate1021(.a(gate193inter11), .b(gate193inter6), .O(gate193inter12));
  nand2 gate1022(.a(gate193inter12), .b(gate193inter1), .O(G642));
nand2 gate194( .a(G588), .b(G589), .O(G645) );
nand2 gate195( .a(G590), .b(G591), .O(G648) );
nand2 gate196( .a(G592), .b(G593), .O(G651) );
nand2 gate197( .a(G594), .b(G595), .O(G654) );

  xor2  gate1177(.a(G597), .b(G596), .O(gate198inter0));
  nand2 gate1178(.a(gate198inter0), .b(s_90), .O(gate198inter1));
  and2  gate1179(.a(G597), .b(G596), .O(gate198inter2));
  inv1  gate1180(.a(s_90), .O(gate198inter3));
  inv1  gate1181(.a(s_91), .O(gate198inter4));
  nand2 gate1182(.a(gate198inter4), .b(gate198inter3), .O(gate198inter5));
  nor2  gate1183(.a(gate198inter5), .b(gate198inter2), .O(gate198inter6));
  inv1  gate1184(.a(G596), .O(gate198inter7));
  inv1  gate1185(.a(G597), .O(gate198inter8));
  nand2 gate1186(.a(gate198inter8), .b(gate198inter7), .O(gate198inter9));
  nand2 gate1187(.a(s_91), .b(gate198inter3), .O(gate198inter10));
  nor2  gate1188(.a(gate198inter10), .b(gate198inter9), .O(gate198inter11));
  nor2  gate1189(.a(gate198inter11), .b(gate198inter6), .O(gate198inter12));
  nand2 gate1190(.a(gate198inter12), .b(gate198inter1), .O(G657));
nand2 gate199( .a(G598), .b(G599), .O(G660) );
nand2 gate200( .a(G600), .b(G601), .O(G663) );

  xor2  gate2003(.a(G607), .b(G602), .O(gate201inter0));
  nand2 gate2004(.a(gate201inter0), .b(s_208), .O(gate201inter1));
  and2  gate2005(.a(G607), .b(G602), .O(gate201inter2));
  inv1  gate2006(.a(s_208), .O(gate201inter3));
  inv1  gate2007(.a(s_209), .O(gate201inter4));
  nand2 gate2008(.a(gate201inter4), .b(gate201inter3), .O(gate201inter5));
  nor2  gate2009(.a(gate201inter5), .b(gate201inter2), .O(gate201inter6));
  inv1  gate2010(.a(G602), .O(gate201inter7));
  inv1  gate2011(.a(G607), .O(gate201inter8));
  nand2 gate2012(.a(gate201inter8), .b(gate201inter7), .O(gate201inter9));
  nand2 gate2013(.a(s_209), .b(gate201inter3), .O(gate201inter10));
  nor2  gate2014(.a(gate201inter10), .b(gate201inter9), .O(gate201inter11));
  nor2  gate2015(.a(gate201inter11), .b(gate201inter6), .O(gate201inter12));
  nand2 gate2016(.a(gate201inter12), .b(gate201inter1), .O(G666));
nand2 gate202( .a(G612), .b(G617), .O(G669) );
nand2 gate203( .a(G602), .b(G612), .O(G672) );
nand2 gate204( .a(G607), .b(G617), .O(G675) );
nand2 gate205( .a(G622), .b(G627), .O(G678) );

  xor2  gate1583(.a(G637), .b(G632), .O(gate206inter0));
  nand2 gate1584(.a(gate206inter0), .b(s_148), .O(gate206inter1));
  and2  gate1585(.a(G637), .b(G632), .O(gate206inter2));
  inv1  gate1586(.a(s_148), .O(gate206inter3));
  inv1  gate1587(.a(s_149), .O(gate206inter4));
  nand2 gate1588(.a(gate206inter4), .b(gate206inter3), .O(gate206inter5));
  nor2  gate1589(.a(gate206inter5), .b(gate206inter2), .O(gate206inter6));
  inv1  gate1590(.a(G632), .O(gate206inter7));
  inv1  gate1591(.a(G637), .O(gate206inter8));
  nand2 gate1592(.a(gate206inter8), .b(gate206inter7), .O(gate206inter9));
  nand2 gate1593(.a(s_149), .b(gate206inter3), .O(gate206inter10));
  nor2  gate1594(.a(gate206inter10), .b(gate206inter9), .O(gate206inter11));
  nor2  gate1595(.a(gate206inter11), .b(gate206inter6), .O(gate206inter12));
  nand2 gate1596(.a(gate206inter12), .b(gate206inter1), .O(G681));

  xor2  gate1471(.a(G632), .b(G622), .O(gate207inter0));
  nand2 gate1472(.a(gate207inter0), .b(s_132), .O(gate207inter1));
  and2  gate1473(.a(G632), .b(G622), .O(gate207inter2));
  inv1  gate1474(.a(s_132), .O(gate207inter3));
  inv1  gate1475(.a(s_133), .O(gate207inter4));
  nand2 gate1476(.a(gate207inter4), .b(gate207inter3), .O(gate207inter5));
  nor2  gate1477(.a(gate207inter5), .b(gate207inter2), .O(gate207inter6));
  inv1  gate1478(.a(G622), .O(gate207inter7));
  inv1  gate1479(.a(G632), .O(gate207inter8));
  nand2 gate1480(.a(gate207inter8), .b(gate207inter7), .O(gate207inter9));
  nand2 gate1481(.a(s_133), .b(gate207inter3), .O(gate207inter10));
  nor2  gate1482(.a(gate207inter10), .b(gate207inter9), .O(gate207inter11));
  nor2  gate1483(.a(gate207inter11), .b(gate207inter6), .O(gate207inter12));
  nand2 gate1484(.a(gate207inter12), .b(gate207inter1), .O(G684));

  xor2  gate2045(.a(G637), .b(G627), .O(gate208inter0));
  nand2 gate2046(.a(gate208inter0), .b(s_214), .O(gate208inter1));
  and2  gate2047(.a(G637), .b(G627), .O(gate208inter2));
  inv1  gate2048(.a(s_214), .O(gate208inter3));
  inv1  gate2049(.a(s_215), .O(gate208inter4));
  nand2 gate2050(.a(gate208inter4), .b(gate208inter3), .O(gate208inter5));
  nor2  gate2051(.a(gate208inter5), .b(gate208inter2), .O(gate208inter6));
  inv1  gate2052(.a(G627), .O(gate208inter7));
  inv1  gate2053(.a(G637), .O(gate208inter8));
  nand2 gate2054(.a(gate208inter8), .b(gate208inter7), .O(gate208inter9));
  nand2 gate2055(.a(s_215), .b(gate208inter3), .O(gate208inter10));
  nor2  gate2056(.a(gate208inter10), .b(gate208inter9), .O(gate208inter11));
  nor2  gate2057(.a(gate208inter11), .b(gate208inter6), .O(gate208inter12));
  nand2 gate2058(.a(gate208inter12), .b(gate208inter1), .O(G687));

  xor2  gate883(.a(G666), .b(G602), .O(gate209inter0));
  nand2 gate884(.a(gate209inter0), .b(s_48), .O(gate209inter1));
  and2  gate885(.a(G666), .b(G602), .O(gate209inter2));
  inv1  gate886(.a(s_48), .O(gate209inter3));
  inv1  gate887(.a(s_49), .O(gate209inter4));
  nand2 gate888(.a(gate209inter4), .b(gate209inter3), .O(gate209inter5));
  nor2  gate889(.a(gate209inter5), .b(gate209inter2), .O(gate209inter6));
  inv1  gate890(.a(G602), .O(gate209inter7));
  inv1  gate891(.a(G666), .O(gate209inter8));
  nand2 gate892(.a(gate209inter8), .b(gate209inter7), .O(gate209inter9));
  nand2 gate893(.a(s_49), .b(gate209inter3), .O(gate209inter10));
  nor2  gate894(.a(gate209inter10), .b(gate209inter9), .O(gate209inter11));
  nor2  gate895(.a(gate209inter11), .b(gate209inter6), .O(gate209inter12));
  nand2 gate896(.a(gate209inter12), .b(gate209inter1), .O(G690));
nand2 gate210( .a(G607), .b(G666), .O(G691) );

  xor2  gate2087(.a(G669), .b(G612), .O(gate211inter0));
  nand2 gate2088(.a(gate211inter0), .b(s_220), .O(gate211inter1));
  and2  gate2089(.a(G669), .b(G612), .O(gate211inter2));
  inv1  gate2090(.a(s_220), .O(gate211inter3));
  inv1  gate2091(.a(s_221), .O(gate211inter4));
  nand2 gate2092(.a(gate211inter4), .b(gate211inter3), .O(gate211inter5));
  nor2  gate2093(.a(gate211inter5), .b(gate211inter2), .O(gate211inter6));
  inv1  gate2094(.a(G612), .O(gate211inter7));
  inv1  gate2095(.a(G669), .O(gate211inter8));
  nand2 gate2096(.a(gate211inter8), .b(gate211inter7), .O(gate211inter9));
  nand2 gate2097(.a(s_221), .b(gate211inter3), .O(gate211inter10));
  nor2  gate2098(.a(gate211inter10), .b(gate211inter9), .O(gate211inter11));
  nor2  gate2099(.a(gate211inter11), .b(gate211inter6), .O(gate211inter12));
  nand2 gate2100(.a(gate211inter12), .b(gate211inter1), .O(G692));
nand2 gate212( .a(G617), .b(G669), .O(G693) );
nand2 gate213( .a(G602), .b(G672), .O(G694) );
nand2 gate214( .a(G612), .b(G672), .O(G695) );

  xor2  gate1107(.a(G675), .b(G607), .O(gate215inter0));
  nand2 gate1108(.a(gate215inter0), .b(s_80), .O(gate215inter1));
  and2  gate1109(.a(G675), .b(G607), .O(gate215inter2));
  inv1  gate1110(.a(s_80), .O(gate215inter3));
  inv1  gate1111(.a(s_81), .O(gate215inter4));
  nand2 gate1112(.a(gate215inter4), .b(gate215inter3), .O(gate215inter5));
  nor2  gate1113(.a(gate215inter5), .b(gate215inter2), .O(gate215inter6));
  inv1  gate1114(.a(G607), .O(gate215inter7));
  inv1  gate1115(.a(G675), .O(gate215inter8));
  nand2 gate1116(.a(gate215inter8), .b(gate215inter7), .O(gate215inter9));
  nand2 gate1117(.a(s_81), .b(gate215inter3), .O(gate215inter10));
  nor2  gate1118(.a(gate215inter10), .b(gate215inter9), .O(gate215inter11));
  nor2  gate1119(.a(gate215inter11), .b(gate215inter6), .O(gate215inter12));
  nand2 gate1120(.a(gate215inter12), .b(gate215inter1), .O(G696));
nand2 gate216( .a(G617), .b(G675), .O(G697) );
nand2 gate217( .a(G622), .b(G678), .O(G698) );
nand2 gate218( .a(G627), .b(G678), .O(G699) );
nand2 gate219( .a(G632), .b(G681), .O(G700) );

  xor2  gate1527(.a(G681), .b(G637), .O(gate220inter0));
  nand2 gate1528(.a(gate220inter0), .b(s_140), .O(gate220inter1));
  and2  gate1529(.a(G681), .b(G637), .O(gate220inter2));
  inv1  gate1530(.a(s_140), .O(gate220inter3));
  inv1  gate1531(.a(s_141), .O(gate220inter4));
  nand2 gate1532(.a(gate220inter4), .b(gate220inter3), .O(gate220inter5));
  nor2  gate1533(.a(gate220inter5), .b(gate220inter2), .O(gate220inter6));
  inv1  gate1534(.a(G637), .O(gate220inter7));
  inv1  gate1535(.a(G681), .O(gate220inter8));
  nand2 gate1536(.a(gate220inter8), .b(gate220inter7), .O(gate220inter9));
  nand2 gate1537(.a(s_141), .b(gate220inter3), .O(gate220inter10));
  nor2  gate1538(.a(gate220inter10), .b(gate220inter9), .O(gate220inter11));
  nor2  gate1539(.a(gate220inter11), .b(gate220inter6), .O(gate220inter12));
  nand2 gate1540(.a(gate220inter12), .b(gate220inter1), .O(G701));

  xor2  gate1863(.a(G684), .b(G622), .O(gate221inter0));
  nand2 gate1864(.a(gate221inter0), .b(s_188), .O(gate221inter1));
  and2  gate1865(.a(G684), .b(G622), .O(gate221inter2));
  inv1  gate1866(.a(s_188), .O(gate221inter3));
  inv1  gate1867(.a(s_189), .O(gate221inter4));
  nand2 gate1868(.a(gate221inter4), .b(gate221inter3), .O(gate221inter5));
  nor2  gate1869(.a(gate221inter5), .b(gate221inter2), .O(gate221inter6));
  inv1  gate1870(.a(G622), .O(gate221inter7));
  inv1  gate1871(.a(G684), .O(gate221inter8));
  nand2 gate1872(.a(gate221inter8), .b(gate221inter7), .O(gate221inter9));
  nand2 gate1873(.a(s_189), .b(gate221inter3), .O(gate221inter10));
  nor2  gate1874(.a(gate221inter10), .b(gate221inter9), .O(gate221inter11));
  nor2  gate1875(.a(gate221inter11), .b(gate221inter6), .O(gate221inter12));
  nand2 gate1876(.a(gate221inter12), .b(gate221inter1), .O(G702));
nand2 gate222( .a(G632), .b(G684), .O(G703) );
nand2 gate223( .a(G627), .b(G687), .O(G704) );
nand2 gate224( .a(G637), .b(G687), .O(G705) );

  xor2  gate645(.a(G691), .b(G690), .O(gate225inter0));
  nand2 gate646(.a(gate225inter0), .b(s_14), .O(gate225inter1));
  and2  gate647(.a(G691), .b(G690), .O(gate225inter2));
  inv1  gate648(.a(s_14), .O(gate225inter3));
  inv1  gate649(.a(s_15), .O(gate225inter4));
  nand2 gate650(.a(gate225inter4), .b(gate225inter3), .O(gate225inter5));
  nor2  gate651(.a(gate225inter5), .b(gate225inter2), .O(gate225inter6));
  inv1  gate652(.a(G690), .O(gate225inter7));
  inv1  gate653(.a(G691), .O(gate225inter8));
  nand2 gate654(.a(gate225inter8), .b(gate225inter7), .O(gate225inter9));
  nand2 gate655(.a(s_15), .b(gate225inter3), .O(gate225inter10));
  nor2  gate656(.a(gate225inter10), .b(gate225inter9), .O(gate225inter11));
  nor2  gate657(.a(gate225inter11), .b(gate225inter6), .O(gate225inter12));
  nand2 gate658(.a(gate225inter12), .b(gate225inter1), .O(G706));
nand2 gate226( .a(G692), .b(G693), .O(G709) );
nand2 gate227( .a(G694), .b(G695), .O(G712) );
nand2 gate228( .a(G696), .b(G697), .O(G715) );
nand2 gate229( .a(G698), .b(G699), .O(G718) );
nand2 gate230( .a(G700), .b(G701), .O(G721) );
nand2 gate231( .a(G702), .b(G703), .O(G724) );
nand2 gate232( .a(G704), .b(G705), .O(G727) );
nand2 gate233( .a(G242), .b(G718), .O(G730) );

  xor2  gate911(.a(G721), .b(G245), .O(gate234inter0));
  nand2 gate912(.a(gate234inter0), .b(s_52), .O(gate234inter1));
  and2  gate913(.a(G721), .b(G245), .O(gate234inter2));
  inv1  gate914(.a(s_52), .O(gate234inter3));
  inv1  gate915(.a(s_53), .O(gate234inter4));
  nand2 gate916(.a(gate234inter4), .b(gate234inter3), .O(gate234inter5));
  nor2  gate917(.a(gate234inter5), .b(gate234inter2), .O(gate234inter6));
  inv1  gate918(.a(G245), .O(gate234inter7));
  inv1  gate919(.a(G721), .O(gate234inter8));
  nand2 gate920(.a(gate234inter8), .b(gate234inter7), .O(gate234inter9));
  nand2 gate921(.a(s_53), .b(gate234inter3), .O(gate234inter10));
  nor2  gate922(.a(gate234inter10), .b(gate234inter9), .O(gate234inter11));
  nor2  gate923(.a(gate234inter11), .b(gate234inter6), .O(gate234inter12));
  nand2 gate924(.a(gate234inter12), .b(gate234inter1), .O(G733));
nand2 gate235( .a(G248), .b(G724), .O(G736) );
nand2 gate236( .a(G251), .b(G727), .O(G739) );
nand2 gate237( .a(G254), .b(G706), .O(G742) );
nand2 gate238( .a(G257), .b(G709), .O(G745) );
nand2 gate239( .a(G260), .b(G712), .O(G748) );
nand2 gate240( .a(G263), .b(G715), .O(G751) );

  xor2  gate855(.a(G730), .b(G242), .O(gate241inter0));
  nand2 gate856(.a(gate241inter0), .b(s_44), .O(gate241inter1));
  and2  gate857(.a(G730), .b(G242), .O(gate241inter2));
  inv1  gate858(.a(s_44), .O(gate241inter3));
  inv1  gate859(.a(s_45), .O(gate241inter4));
  nand2 gate860(.a(gate241inter4), .b(gate241inter3), .O(gate241inter5));
  nor2  gate861(.a(gate241inter5), .b(gate241inter2), .O(gate241inter6));
  inv1  gate862(.a(G242), .O(gate241inter7));
  inv1  gate863(.a(G730), .O(gate241inter8));
  nand2 gate864(.a(gate241inter8), .b(gate241inter7), .O(gate241inter9));
  nand2 gate865(.a(s_45), .b(gate241inter3), .O(gate241inter10));
  nor2  gate866(.a(gate241inter10), .b(gate241inter9), .O(gate241inter11));
  nor2  gate867(.a(gate241inter11), .b(gate241inter6), .O(gate241inter12));
  nand2 gate868(.a(gate241inter12), .b(gate241inter1), .O(G754));
nand2 gate242( .a(G718), .b(G730), .O(G755) );

  xor2  gate1611(.a(G733), .b(G245), .O(gate243inter0));
  nand2 gate1612(.a(gate243inter0), .b(s_152), .O(gate243inter1));
  and2  gate1613(.a(G733), .b(G245), .O(gate243inter2));
  inv1  gate1614(.a(s_152), .O(gate243inter3));
  inv1  gate1615(.a(s_153), .O(gate243inter4));
  nand2 gate1616(.a(gate243inter4), .b(gate243inter3), .O(gate243inter5));
  nor2  gate1617(.a(gate243inter5), .b(gate243inter2), .O(gate243inter6));
  inv1  gate1618(.a(G245), .O(gate243inter7));
  inv1  gate1619(.a(G733), .O(gate243inter8));
  nand2 gate1620(.a(gate243inter8), .b(gate243inter7), .O(gate243inter9));
  nand2 gate1621(.a(s_153), .b(gate243inter3), .O(gate243inter10));
  nor2  gate1622(.a(gate243inter10), .b(gate243inter9), .O(gate243inter11));
  nor2  gate1623(.a(gate243inter11), .b(gate243inter6), .O(gate243inter12));
  nand2 gate1624(.a(gate243inter12), .b(gate243inter1), .O(G756));
nand2 gate244( .a(G721), .b(G733), .O(G757) );
nand2 gate245( .a(G248), .b(G736), .O(G758) );

  xor2  gate1457(.a(G736), .b(G724), .O(gate246inter0));
  nand2 gate1458(.a(gate246inter0), .b(s_130), .O(gate246inter1));
  and2  gate1459(.a(G736), .b(G724), .O(gate246inter2));
  inv1  gate1460(.a(s_130), .O(gate246inter3));
  inv1  gate1461(.a(s_131), .O(gate246inter4));
  nand2 gate1462(.a(gate246inter4), .b(gate246inter3), .O(gate246inter5));
  nor2  gate1463(.a(gate246inter5), .b(gate246inter2), .O(gate246inter6));
  inv1  gate1464(.a(G724), .O(gate246inter7));
  inv1  gate1465(.a(G736), .O(gate246inter8));
  nand2 gate1466(.a(gate246inter8), .b(gate246inter7), .O(gate246inter9));
  nand2 gate1467(.a(s_131), .b(gate246inter3), .O(gate246inter10));
  nor2  gate1468(.a(gate246inter10), .b(gate246inter9), .O(gate246inter11));
  nor2  gate1469(.a(gate246inter11), .b(gate246inter6), .O(gate246inter12));
  nand2 gate1470(.a(gate246inter12), .b(gate246inter1), .O(G759));
nand2 gate247( .a(G251), .b(G739), .O(G760) );

  xor2  gate743(.a(G739), .b(G727), .O(gate248inter0));
  nand2 gate744(.a(gate248inter0), .b(s_28), .O(gate248inter1));
  and2  gate745(.a(G739), .b(G727), .O(gate248inter2));
  inv1  gate746(.a(s_28), .O(gate248inter3));
  inv1  gate747(.a(s_29), .O(gate248inter4));
  nand2 gate748(.a(gate248inter4), .b(gate248inter3), .O(gate248inter5));
  nor2  gate749(.a(gate248inter5), .b(gate248inter2), .O(gate248inter6));
  inv1  gate750(.a(G727), .O(gate248inter7));
  inv1  gate751(.a(G739), .O(gate248inter8));
  nand2 gate752(.a(gate248inter8), .b(gate248inter7), .O(gate248inter9));
  nand2 gate753(.a(s_29), .b(gate248inter3), .O(gate248inter10));
  nor2  gate754(.a(gate248inter10), .b(gate248inter9), .O(gate248inter11));
  nor2  gate755(.a(gate248inter11), .b(gate248inter6), .O(gate248inter12));
  nand2 gate756(.a(gate248inter12), .b(gate248inter1), .O(G761));
nand2 gate249( .a(G254), .b(G742), .O(G762) );

  xor2  gate1037(.a(G742), .b(G706), .O(gate250inter0));
  nand2 gate1038(.a(gate250inter0), .b(s_70), .O(gate250inter1));
  and2  gate1039(.a(G742), .b(G706), .O(gate250inter2));
  inv1  gate1040(.a(s_70), .O(gate250inter3));
  inv1  gate1041(.a(s_71), .O(gate250inter4));
  nand2 gate1042(.a(gate250inter4), .b(gate250inter3), .O(gate250inter5));
  nor2  gate1043(.a(gate250inter5), .b(gate250inter2), .O(gate250inter6));
  inv1  gate1044(.a(G706), .O(gate250inter7));
  inv1  gate1045(.a(G742), .O(gate250inter8));
  nand2 gate1046(.a(gate250inter8), .b(gate250inter7), .O(gate250inter9));
  nand2 gate1047(.a(s_71), .b(gate250inter3), .O(gate250inter10));
  nor2  gate1048(.a(gate250inter10), .b(gate250inter9), .O(gate250inter11));
  nor2  gate1049(.a(gate250inter11), .b(gate250inter6), .O(gate250inter12));
  nand2 gate1050(.a(gate250inter12), .b(gate250inter1), .O(G763));

  xor2  gate631(.a(G745), .b(G257), .O(gate251inter0));
  nand2 gate632(.a(gate251inter0), .b(s_12), .O(gate251inter1));
  and2  gate633(.a(G745), .b(G257), .O(gate251inter2));
  inv1  gate634(.a(s_12), .O(gate251inter3));
  inv1  gate635(.a(s_13), .O(gate251inter4));
  nand2 gate636(.a(gate251inter4), .b(gate251inter3), .O(gate251inter5));
  nor2  gate637(.a(gate251inter5), .b(gate251inter2), .O(gate251inter6));
  inv1  gate638(.a(G257), .O(gate251inter7));
  inv1  gate639(.a(G745), .O(gate251inter8));
  nand2 gate640(.a(gate251inter8), .b(gate251inter7), .O(gate251inter9));
  nand2 gate641(.a(s_13), .b(gate251inter3), .O(gate251inter10));
  nor2  gate642(.a(gate251inter10), .b(gate251inter9), .O(gate251inter11));
  nor2  gate643(.a(gate251inter11), .b(gate251inter6), .O(gate251inter12));
  nand2 gate644(.a(gate251inter12), .b(gate251inter1), .O(G764));

  xor2  gate1989(.a(G745), .b(G709), .O(gate252inter0));
  nand2 gate1990(.a(gate252inter0), .b(s_206), .O(gate252inter1));
  and2  gate1991(.a(G745), .b(G709), .O(gate252inter2));
  inv1  gate1992(.a(s_206), .O(gate252inter3));
  inv1  gate1993(.a(s_207), .O(gate252inter4));
  nand2 gate1994(.a(gate252inter4), .b(gate252inter3), .O(gate252inter5));
  nor2  gate1995(.a(gate252inter5), .b(gate252inter2), .O(gate252inter6));
  inv1  gate1996(.a(G709), .O(gate252inter7));
  inv1  gate1997(.a(G745), .O(gate252inter8));
  nand2 gate1998(.a(gate252inter8), .b(gate252inter7), .O(gate252inter9));
  nand2 gate1999(.a(s_207), .b(gate252inter3), .O(gate252inter10));
  nor2  gate2000(.a(gate252inter10), .b(gate252inter9), .O(gate252inter11));
  nor2  gate2001(.a(gate252inter11), .b(gate252inter6), .O(gate252inter12));
  nand2 gate2002(.a(gate252inter12), .b(gate252inter1), .O(G765));
nand2 gate253( .a(G260), .b(G748), .O(G766) );
nand2 gate254( .a(G712), .b(G748), .O(G767) );

  xor2  gate1709(.a(G751), .b(G263), .O(gate255inter0));
  nand2 gate1710(.a(gate255inter0), .b(s_166), .O(gate255inter1));
  and2  gate1711(.a(G751), .b(G263), .O(gate255inter2));
  inv1  gate1712(.a(s_166), .O(gate255inter3));
  inv1  gate1713(.a(s_167), .O(gate255inter4));
  nand2 gate1714(.a(gate255inter4), .b(gate255inter3), .O(gate255inter5));
  nor2  gate1715(.a(gate255inter5), .b(gate255inter2), .O(gate255inter6));
  inv1  gate1716(.a(G263), .O(gate255inter7));
  inv1  gate1717(.a(G751), .O(gate255inter8));
  nand2 gate1718(.a(gate255inter8), .b(gate255inter7), .O(gate255inter9));
  nand2 gate1719(.a(s_167), .b(gate255inter3), .O(gate255inter10));
  nor2  gate1720(.a(gate255inter10), .b(gate255inter9), .O(gate255inter11));
  nor2  gate1721(.a(gate255inter11), .b(gate255inter6), .O(gate255inter12));
  nand2 gate1722(.a(gate255inter12), .b(gate255inter1), .O(G768));
nand2 gate256( .a(G715), .b(G751), .O(G769) );
nand2 gate257( .a(G754), .b(G755), .O(G770) );

  xor2  gate925(.a(G757), .b(G756), .O(gate258inter0));
  nand2 gate926(.a(gate258inter0), .b(s_54), .O(gate258inter1));
  and2  gate927(.a(G757), .b(G756), .O(gate258inter2));
  inv1  gate928(.a(s_54), .O(gate258inter3));
  inv1  gate929(.a(s_55), .O(gate258inter4));
  nand2 gate930(.a(gate258inter4), .b(gate258inter3), .O(gate258inter5));
  nor2  gate931(.a(gate258inter5), .b(gate258inter2), .O(gate258inter6));
  inv1  gate932(.a(G756), .O(gate258inter7));
  inv1  gate933(.a(G757), .O(gate258inter8));
  nand2 gate934(.a(gate258inter8), .b(gate258inter7), .O(gate258inter9));
  nand2 gate935(.a(s_55), .b(gate258inter3), .O(gate258inter10));
  nor2  gate936(.a(gate258inter10), .b(gate258inter9), .O(gate258inter11));
  nor2  gate937(.a(gate258inter11), .b(gate258inter6), .O(gate258inter12));
  nand2 gate938(.a(gate258inter12), .b(gate258inter1), .O(G773));
nand2 gate259( .a(G758), .b(G759), .O(G776) );
nand2 gate260( .a(G760), .b(G761), .O(G779) );

  xor2  gate757(.a(G763), .b(G762), .O(gate261inter0));
  nand2 gate758(.a(gate261inter0), .b(s_30), .O(gate261inter1));
  and2  gate759(.a(G763), .b(G762), .O(gate261inter2));
  inv1  gate760(.a(s_30), .O(gate261inter3));
  inv1  gate761(.a(s_31), .O(gate261inter4));
  nand2 gate762(.a(gate261inter4), .b(gate261inter3), .O(gate261inter5));
  nor2  gate763(.a(gate261inter5), .b(gate261inter2), .O(gate261inter6));
  inv1  gate764(.a(G762), .O(gate261inter7));
  inv1  gate765(.a(G763), .O(gate261inter8));
  nand2 gate766(.a(gate261inter8), .b(gate261inter7), .O(gate261inter9));
  nand2 gate767(.a(s_31), .b(gate261inter3), .O(gate261inter10));
  nor2  gate768(.a(gate261inter10), .b(gate261inter9), .O(gate261inter11));
  nor2  gate769(.a(gate261inter11), .b(gate261inter6), .O(gate261inter12));
  nand2 gate770(.a(gate261inter12), .b(gate261inter1), .O(G782));

  xor2  gate1093(.a(G765), .b(G764), .O(gate262inter0));
  nand2 gate1094(.a(gate262inter0), .b(s_78), .O(gate262inter1));
  and2  gate1095(.a(G765), .b(G764), .O(gate262inter2));
  inv1  gate1096(.a(s_78), .O(gate262inter3));
  inv1  gate1097(.a(s_79), .O(gate262inter4));
  nand2 gate1098(.a(gate262inter4), .b(gate262inter3), .O(gate262inter5));
  nor2  gate1099(.a(gate262inter5), .b(gate262inter2), .O(gate262inter6));
  inv1  gate1100(.a(G764), .O(gate262inter7));
  inv1  gate1101(.a(G765), .O(gate262inter8));
  nand2 gate1102(.a(gate262inter8), .b(gate262inter7), .O(gate262inter9));
  nand2 gate1103(.a(s_79), .b(gate262inter3), .O(gate262inter10));
  nor2  gate1104(.a(gate262inter10), .b(gate262inter9), .O(gate262inter11));
  nor2  gate1105(.a(gate262inter11), .b(gate262inter6), .O(gate262inter12));
  nand2 gate1106(.a(gate262inter12), .b(gate262inter1), .O(G785));
nand2 gate263( .a(G766), .b(G767), .O(G788) );
nand2 gate264( .a(G768), .b(G769), .O(G791) );
nand2 gate265( .a(G642), .b(G770), .O(G794) );

  xor2  gate1149(.a(G773), .b(G645), .O(gate266inter0));
  nand2 gate1150(.a(gate266inter0), .b(s_86), .O(gate266inter1));
  and2  gate1151(.a(G773), .b(G645), .O(gate266inter2));
  inv1  gate1152(.a(s_86), .O(gate266inter3));
  inv1  gate1153(.a(s_87), .O(gate266inter4));
  nand2 gate1154(.a(gate266inter4), .b(gate266inter3), .O(gate266inter5));
  nor2  gate1155(.a(gate266inter5), .b(gate266inter2), .O(gate266inter6));
  inv1  gate1156(.a(G645), .O(gate266inter7));
  inv1  gate1157(.a(G773), .O(gate266inter8));
  nand2 gate1158(.a(gate266inter8), .b(gate266inter7), .O(gate266inter9));
  nand2 gate1159(.a(s_87), .b(gate266inter3), .O(gate266inter10));
  nor2  gate1160(.a(gate266inter10), .b(gate266inter9), .O(gate266inter11));
  nor2  gate1161(.a(gate266inter11), .b(gate266inter6), .O(gate266inter12));
  nand2 gate1162(.a(gate266inter12), .b(gate266inter1), .O(G797));
nand2 gate267( .a(G648), .b(G776), .O(G800) );
nand2 gate268( .a(G651), .b(G779), .O(G803) );

  xor2  gate1275(.a(G782), .b(G654), .O(gate269inter0));
  nand2 gate1276(.a(gate269inter0), .b(s_104), .O(gate269inter1));
  and2  gate1277(.a(G782), .b(G654), .O(gate269inter2));
  inv1  gate1278(.a(s_104), .O(gate269inter3));
  inv1  gate1279(.a(s_105), .O(gate269inter4));
  nand2 gate1280(.a(gate269inter4), .b(gate269inter3), .O(gate269inter5));
  nor2  gate1281(.a(gate269inter5), .b(gate269inter2), .O(gate269inter6));
  inv1  gate1282(.a(G654), .O(gate269inter7));
  inv1  gate1283(.a(G782), .O(gate269inter8));
  nand2 gate1284(.a(gate269inter8), .b(gate269inter7), .O(gate269inter9));
  nand2 gate1285(.a(s_105), .b(gate269inter3), .O(gate269inter10));
  nor2  gate1286(.a(gate269inter10), .b(gate269inter9), .O(gate269inter11));
  nor2  gate1287(.a(gate269inter11), .b(gate269inter6), .O(gate269inter12));
  nand2 gate1288(.a(gate269inter12), .b(gate269inter1), .O(G806));
nand2 gate270( .a(G657), .b(G785), .O(G809) );
nand2 gate271( .a(G660), .b(G788), .O(G812) );
nand2 gate272( .a(G663), .b(G791), .O(G815) );
nand2 gate273( .a(G642), .b(G794), .O(G818) );
nand2 gate274( .a(G770), .b(G794), .O(G819) );

  xor2  gate953(.a(G797), .b(G645), .O(gate275inter0));
  nand2 gate954(.a(gate275inter0), .b(s_58), .O(gate275inter1));
  and2  gate955(.a(G797), .b(G645), .O(gate275inter2));
  inv1  gate956(.a(s_58), .O(gate275inter3));
  inv1  gate957(.a(s_59), .O(gate275inter4));
  nand2 gate958(.a(gate275inter4), .b(gate275inter3), .O(gate275inter5));
  nor2  gate959(.a(gate275inter5), .b(gate275inter2), .O(gate275inter6));
  inv1  gate960(.a(G645), .O(gate275inter7));
  inv1  gate961(.a(G797), .O(gate275inter8));
  nand2 gate962(.a(gate275inter8), .b(gate275inter7), .O(gate275inter9));
  nand2 gate963(.a(s_59), .b(gate275inter3), .O(gate275inter10));
  nor2  gate964(.a(gate275inter10), .b(gate275inter9), .O(gate275inter11));
  nor2  gate965(.a(gate275inter11), .b(gate275inter6), .O(gate275inter12));
  nand2 gate966(.a(gate275inter12), .b(gate275inter1), .O(G820));

  xor2  gate575(.a(G797), .b(G773), .O(gate276inter0));
  nand2 gate576(.a(gate276inter0), .b(s_4), .O(gate276inter1));
  and2  gate577(.a(G797), .b(G773), .O(gate276inter2));
  inv1  gate578(.a(s_4), .O(gate276inter3));
  inv1  gate579(.a(s_5), .O(gate276inter4));
  nand2 gate580(.a(gate276inter4), .b(gate276inter3), .O(gate276inter5));
  nor2  gate581(.a(gate276inter5), .b(gate276inter2), .O(gate276inter6));
  inv1  gate582(.a(G773), .O(gate276inter7));
  inv1  gate583(.a(G797), .O(gate276inter8));
  nand2 gate584(.a(gate276inter8), .b(gate276inter7), .O(gate276inter9));
  nand2 gate585(.a(s_5), .b(gate276inter3), .O(gate276inter10));
  nor2  gate586(.a(gate276inter10), .b(gate276inter9), .O(gate276inter11));
  nor2  gate587(.a(gate276inter11), .b(gate276inter6), .O(gate276inter12));
  nand2 gate588(.a(gate276inter12), .b(gate276inter1), .O(G821));

  xor2  gate1653(.a(G800), .b(G648), .O(gate277inter0));
  nand2 gate1654(.a(gate277inter0), .b(s_158), .O(gate277inter1));
  and2  gate1655(.a(G800), .b(G648), .O(gate277inter2));
  inv1  gate1656(.a(s_158), .O(gate277inter3));
  inv1  gate1657(.a(s_159), .O(gate277inter4));
  nand2 gate1658(.a(gate277inter4), .b(gate277inter3), .O(gate277inter5));
  nor2  gate1659(.a(gate277inter5), .b(gate277inter2), .O(gate277inter6));
  inv1  gate1660(.a(G648), .O(gate277inter7));
  inv1  gate1661(.a(G800), .O(gate277inter8));
  nand2 gate1662(.a(gate277inter8), .b(gate277inter7), .O(gate277inter9));
  nand2 gate1663(.a(s_159), .b(gate277inter3), .O(gate277inter10));
  nor2  gate1664(.a(gate277inter10), .b(gate277inter9), .O(gate277inter11));
  nor2  gate1665(.a(gate277inter11), .b(gate277inter6), .O(gate277inter12));
  nand2 gate1666(.a(gate277inter12), .b(gate277inter1), .O(G822));
nand2 gate278( .a(G776), .b(G800), .O(G823) );

  xor2  gate1359(.a(G803), .b(G651), .O(gate279inter0));
  nand2 gate1360(.a(gate279inter0), .b(s_116), .O(gate279inter1));
  and2  gate1361(.a(G803), .b(G651), .O(gate279inter2));
  inv1  gate1362(.a(s_116), .O(gate279inter3));
  inv1  gate1363(.a(s_117), .O(gate279inter4));
  nand2 gate1364(.a(gate279inter4), .b(gate279inter3), .O(gate279inter5));
  nor2  gate1365(.a(gate279inter5), .b(gate279inter2), .O(gate279inter6));
  inv1  gate1366(.a(G651), .O(gate279inter7));
  inv1  gate1367(.a(G803), .O(gate279inter8));
  nand2 gate1368(.a(gate279inter8), .b(gate279inter7), .O(gate279inter9));
  nand2 gate1369(.a(s_117), .b(gate279inter3), .O(gate279inter10));
  nor2  gate1370(.a(gate279inter10), .b(gate279inter9), .O(gate279inter11));
  nor2  gate1371(.a(gate279inter11), .b(gate279inter6), .O(gate279inter12));
  nand2 gate1372(.a(gate279inter12), .b(gate279inter1), .O(G824));
nand2 gate280( .a(G779), .b(G803), .O(G825) );
nand2 gate281( .a(G654), .b(G806), .O(G826) );
nand2 gate282( .a(G782), .b(G806), .O(G827) );
nand2 gate283( .a(G657), .b(G809), .O(G828) );
nand2 gate284( .a(G785), .b(G809), .O(G829) );
nand2 gate285( .a(G660), .b(G812), .O(G830) );
nand2 gate286( .a(G788), .b(G812), .O(G831) );
nand2 gate287( .a(G663), .b(G815), .O(G832) );
nand2 gate288( .a(G791), .b(G815), .O(G833) );
nand2 gate289( .a(G818), .b(G819), .O(G834) );
nand2 gate290( .a(G820), .b(G821), .O(G847) );
nand2 gate291( .a(G822), .b(G823), .O(G860) );
nand2 gate292( .a(G824), .b(G825), .O(G873) );

  xor2  gate2059(.a(G829), .b(G828), .O(gate293inter0));
  nand2 gate2060(.a(gate293inter0), .b(s_216), .O(gate293inter1));
  and2  gate2061(.a(G829), .b(G828), .O(gate293inter2));
  inv1  gate2062(.a(s_216), .O(gate293inter3));
  inv1  gate2063(.a(s_217), .O(gate293inter4));
  nand2 gate2064(.a(gate293inter4), .b(gate293inter3), .O(gate293inter5));
  nor2  gate2065(.a(gate293inter5), .b(gate293inter2), .O(gate293inter6));
  inv1  gate2066(.a(G828), .O(gate293inter7));
  inv1  gate2067(.a(G829), .O(gate293inter8));
  nand2 gate2068(.a(gate293inter8), .b(gate293inter7), .O(gate293inter9));
  nand2 gate2069(.a(s_217), .b(gate293inter3), .O(gate293inter10));
  nor2  gate2070(.a(gate293inter10), .b(gate293inter9), .O(gate293inter11));
  nor2  gate2071(.a(gate293inter11), .b(gate293inter6), .O(gate293inter12));
  nand2 gate2072(.a(gate293inter12), .b(gate293inter1), .O(G886));

  xor2  gate1681(.a(G833), .b(G832), .O(gate294inter0));
  nand2 gate1682(.a(gate294inter0), .b(s_162), .O(gate294inter1));
  and2  gate1683(.a(G833), .b(G832), .O(gate294inter2));
  inv1  gate1684(.a(s_162), .O(gate294inter3));
  inv1  gate1685(.a(s_163), .O(gate294inter4));
  nand2 gate1686(.a(gate294inter4), .b(gate294inter3), .O(gate294inter5));
  nor2  gate1687(.a(gate294inter5), .b(gate294inter2), .O(gate294inter6));
  inv1  gate1688(.a(G832), .O(gate294inter7));
  inv1  gate1689(.a(G833), .O(gate294inter8));
  nand2 gate1690(.a(gate294inter8), .b(gate294inter7), .O(gate294inter9));
  nand2 gate1691(.a(s_163), .b(gate294inter3), .O(gate294inter10));
  nor2  gate1692(.a(gate294inter10), .b(gate294inter9), .O(gate294inter11));
  nor2  gate1693(.a(gate294inter11), .b(gate294inter6), .O(gate294inter12));
  nand2 gate1694(.a(gate294inter12), .b(gate294inter1), .O(G899));
nand2 gate295( .a(G830), .b(G831), .O(G912) );
nand2 gate296( .a(G826), .b(G827), .O(G925) );
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );
nand2 gate387( .a(G1), .b(G1036), .O(G1132) );
nand2 gate388( .a(G2), .b(G1039), .O(G1135) );
nand2 gate389( .a(G3), .b(G1042), .O(G1138) );
nand2 gate390( .a(G4), .b(G1045), .O(G1141) );
nand2 gate391( .a(G5), .b(G1048), .O(G1144) );
nand2 gate392( .a(G6), .b(G1051), .O(G1147) );

  xor2  gate1779(.a(G1054), .b(G7), .O(gate393inter0));
  nand2 gate1780(.a(gate393inter0), .b(s_176), .O(gate393inter1));
  and2  gate1781(.a(G1054), .b(G7), .O(gate393inter2));
  inv1  gate1782(.a(s_176), .O(gate393inter3));
  inv1  gate1783(.a(s_177), .O(gate393inter4));
  nand2 gate1784(.a(gate393inter4), .b(gate393inter3), .O(gate393inter5));
  nor2  gate1785(.a(gate393inter5), .b(gate393inter2), .O(gate393inter6));
  inv1  gate1786(.a(G7), .O(gate393inter7));
  inv1  gate1787(.a(G1054), .O(gate393inter8));
  nand2 gate1788(.a(gate393inter8), .b(gate393inter7), .O(gate393inter9));
  nand2 gate1789(.a(s_177), .b(gate393inter3), .O(gate393inter10));
  nor2  gate1790(.a(gate393inter10), .b(gate393inter9), .O(gate393inter11));
  nor2  gate1791(.a(gate393inter11), .b(gate393inter6), .O(gate393inter12));
  nand2 gate1792(.a(gate393inter12), .b(gate393inter1), .O(G1150));
nand2 gate394( .a(G8), .b(G1057), .O(G1153) );
nand2 gate395( .a(G9), .b(G1060), .O(G1156) );

  xor2  gate1723(.a(G1063), .b(G10), .O(gate396inter0));
  nand2 gate1724(.a(gate396inter0), .b(s_168), .O(gate396inter1));
  and2  gate1725(.a(G1063), .b(G10), .O(gate396inter2));
  inv1  gate1726(.a(s_168), .O(gate396inter3));
  inv1  gate1727(.a(s_169), .O(gate396inter4));
  nand2 gate1728(.a(gate396inter4), .b(gate396inter3), .O(gate396inter5));
  nor2  gate1729(.a(gate396inter5), .b(gate396inter2), .O(gate396inter6));
  inv1  gate1730(.a(G10), .O(gate396inter7));
  inv1  gate1731(.a(G1063), .O(gate396inter8));
  nand2 gate1732(.a(gate396inter8), .b(gate396inter7), .O(gate396inter9));
  nand2 gate1733(.a(s_169), .b(gate396inter3), .O(gate396inter10));
  nor2  gate1734(.a(gate396inter10), .b(gate396inter9), .O(gate396inter11));
  nor2  gate1735(.a(gate396inter11), .b(gate396inter6), .O(gate396inter12));
  nand2 gate1736(.a(gate396inter12), .b(gate396inter1), .O(G1159));

  xor2  gate2031(.a(G1066), .b(G11), .O(gate397inter0));
  nand2 gate2032(.a(gate397inter0), .b(s_212), .O(gate397inter1));
  and2  gate2033(.a(G1066), .b(G11), .O(gate397inter2));
  inv1  gate2034(.a(s_212), .O(gate397inter3));
  inv1  gate2035(.a(s_213), .O(gate397inter4));
  nand2 gate2036(.a(gate397inter4), .b(gate397inter3), .O(gate397inter5));
  nor2  gate2037(.a(gate397inter5), .b(gate397inter2), .O(gate397inter6));
  inv1  gate2038(.a(G11), .O(gate397inter7));
  inv1  gate2039(.a(G1066), .O(gate397inter8));
  nand2 gate2040(.a(gate397inter8), .b(gate397inter7), .O(gate397inter9));
  nand2 gate2041(.a(s_213), .b(gate397inter3), .O(gate397inter10));
  nor2  gate2042(.a(gate397inter10), .b(gate397inter9), .O(gate397inter11));
  nor2  gate2043(.a(gate397inter11), .b(gate397inter6), .O(gate397inter12));
  nand2 gate2044(.a(gate397inter12), .b(gate397inter1), .O(G1162));
nand2 gate398( .a(G12), .b(G1069), .O(G1165) );
nand2 gate399( .a(G13), .b(G1072), .O(G1168) );

  xor2  gate1513(.a(G1075), .b(G14), .O(gate400inter0));
  nand2 gate1514(.a(gate400inter0), .b(s_138), .O(gate400inter1));
  and2  gate1515(.a(G1075), .b(G14), .O(gate400inter2));
  inv1  gate1516(.a(s_138), .O(gate400inter3));
  inv1  gate1517(.a(s_139), .O(gate400inter4));
  nand2 gate1518(.a(gate400inter4), .b(gate400inter3), .O(gate400inter5));
  nor2  gate1519(.a(gate400inter5), .b(gate400inter2), .O(gate400inter6));
  inv1  gate1520(.a(G14), .O(gate400inter7));
  inv1  gate1521(.a(G1075), .O(gate400inter8));
  nand2 gate1522(.a(gate400inter8), .b(gate400inter7), .O(gate400inter9));
  nand2 gate1523(.a(s_139), .b(gate400inter3), .O(gate400inter10));
  nor2  gate1524(.a(gate400inter10), .b(gate400inter9), .O(gate400inter11));
  nor2  gate1525(.a(gate400inter11), .b(gate400inter6), .O(gate400inter12));
  nand2 gate1526(.a(gate400inter12), .b(gate400inter1), .O(G1171));
nand2 gate401( .a(G15), .b(G1078), .O(G1174) );

  xor2  gate547(.a(G1081), .b(G16), .O(gate402inter0));
  nand2 gate548(.a(gate402inter0), .b(s_0), .O(gate402inter1));
  and2  gate549(.a(G1081), .b(G16), .O(gate402inter2));
  inv1  gate550(.a(s_0), .O(gate402inter3));
  inv1  gate551(.a(s_1), .O(gate402inter4));
  nand2 gate552(.a(gate402inter4), .b(gate402inter3), .O(gate402inter5));
  nor2  gate553(.a(gate402inter5), .b(gate402inter2), .O(gate402inter6));
  inv1  gate554(.a(G16), .O(gate402inter7));
  inv1  gate555(.a(G1081), .O(gate402inter8));
  nand2 gate556(.a(gate402inter8), .b(gate402inter7), .O(gate402inter9));
  nand2 gate557(.a(s_1), .b(gate402inter3), .O(gate402inter10));
  nor2  gate558(.a(gate402inter10), .b(gate402inter9), .O(gate402inter11));
  nor2  gate559(.a(gate402inter11), .b(gate402inter6), .O(gate402inter12));
  nand2 gate560(.a(gate402inter12), .b(gate402inter1), .O(G1177));
nand2 gate403( .a(G17), .b(G1084), .O(G1180) );
nand2 gate404( .a(G18), .b(G1087), .O(G1183) );
nand2 gate405( .a(G19), .b(G1090), .O(G1186) );
nand2 gate406( .a(G20), .b(G1093), .O(G1189) );
nand2 gate407( .a(G21), .b(G1096), .O(G1192) );

  xor2  gate1485(.a(G1099), .b(G22), .O(gate408inter0));
  nand2 gate1486(.a(gate408inter0), .b(s_134), .O(gate408inter1));
  and2  gate1487(.a(G1099), .b(G22), .O(gate408inter2));
  inv1  gate1488(.a(s_134), .O(gate408inter3));
  inv1  gate1489(.a(s_135), .O(gate408inter4));
  nand2 gate1490(.a(gate408inter4), .b(gate408inter3), .O(gate408inter5));
  nor2  gate1491(.a(gate408inter5), .b(gate408inter2), .O(gate408inter6));
  inv1  gate1492(.a(G22), .O(gate408inter7));
  inv1  gate1493(.a(G1099), .O(gate408inter8));
  nand2 gate1494(.a(gate408inter8), .b(gate408inter7), .O(gate408inter9));
  nand2 gate1495(.a(s_135), .b(gate408inter3), .O(gate408inter10));
  nor2  gate1496(.a(gate408inter10), .b(gate408inter9), .O(gate408inter11));
  nor2  gate1497(.a(gate408inter11), .b(gate408inter6), .O(gate408inter12));
  nand2 gate1498(.a(gate408inter12), .b(gate408inter1), .O(G1195));

  xor2  gate827(.a(G1102), .b(G23), .O(gate409inter0));
  nand2 gate828(.a(gate409inter0), .b(s_40), .O(gate409inter1));
  and2  gate829(.a(G1102), .b(G23), .O(gate409inter2));
  inv1  gate830(.a(s_40), .O(gate409inter3));
  inv1  gate831(.a(s_41), .O(gate409inter4));
  nand2 gate832(.a(gate409inter4), .b(gate409inter3), .O(gate409inter5));
  nor2  gate833(.a(gate409inter5), .b(gate409inter2), .O(gate409inter6));
  inv1  gate834(.a(G23), .O(gate409inter7));
  inv1  gate835(.a(G1102), .O(gate409inter8));
  nand2 gate836(.a(gate409inter8), .b(gate409inter7), .O(gate409inter9));
  nand2 gate837(.a(s_41), .b(gate409inter3), .O(gate409inter10));
  nor2  gate838(.a(gate409inter10), .b(gate409inter9), .O(gate409inter11));
  nor2  gate839(.a(gate409inter11), .b(gate409inter6), .O(gate409inter12));
  nand2 gate840(.a(gate409inter12), .b(gate409inter1), .O(G1198));
nand2 gate410( .a(G24), .b(G1105), .O(G1201) );

  xor2  gate939(.a(G1108), .b(G25), .O(gate411inter0));
  nand2 gate940(.a(gate411inter0), .b(s_56), .O(gate411inter1));
  and2  gate941(.a(G1108), .b(G25), .O(gate411inter2));
  inv1  gate942(.a(s_56), .O(gate411inter3));
  inv1  gate943(.a(s_57), .O(gate411inter4));
  nand2 gate944(.a(gate411inter4), .b(gate411inter3), .O(gate411inter5));
  nor2  gate945(.a(gate411inter5), .b(gate411inter2), .O(gate411inter6));
  inv1  gate946(.a(G25), .O(gate411inter7));
  inv1  gate947(.a(G1108), .O(gate411inter8));
  nand2 gate948(.a(gate411inter8), .b(gate411inter7), .O(gate411inter9));
  nand2 gate949(.a(s_57), .b(gate411inter3), .O(gate411inter10));
  nor2  gate950(.a(gate411inter10), .b(gate411inter9), .O(gate411inter11));
  nor2  gate951(.a(gate411inter11), .b(gate411inter6), .O(gate411inter12));
  nand2 gate952(.a(gate411inter12), .b(gate411inter1), .O(G1204));

  xor2  gate2073(.a(G1111), .b(G26), .O(gate412inter0));
  nand2 gate2074(.a(gate412inter0), .b(s_218), .O(gate412inter1));
  and2  gate2075(.a(G1111), .b(G26), .O(gate412inter2));
  inv1  gate2076(.a(s_218), .O(gate412inter3));
  inv1  gate2077(.a(s_219), .O(gate412inter4));
  nand2 gate2078(.a(gate412inter4), .b(gate412inter3), .O(gate412inter5));
  nor2  gate2079(.a(gate412inter5), .b(gate412inter2), .O(gate412inter6));
  inv1  gate2080(.a(G26), .O(gate412inter7));
  inv1  gate2081(.a(G1111), .O(gate412inter8));
  nand2 gate2082(.a(gate412inter8), .b(gate412inter7), .O(gate412inter9));
  nand2 gate2083(.a(s_219), .b(gate412inter3), .O(gate412inter10));
  nor2  gate2084(.a(gate412inter10), .b(gate412inter9), .O(gate412inter11));
  nor2  gate2085(.a(gate412inter11), .b(gate412inter6), .O(gate412inter12));
  nand2 gate2086(.a(gate412inter12), .b(gate412inter1), .O(G1207));

  xor2  gate1429(.a(G1114), .b(G27), .O(gate413inter0));
  nand2 gate1430(.a(gate413inter0), .b(s_126), .O(gate413inter1));
  and2  gate1431(.a(G1114), .b(G27), .O(gate413inter2));
  inv1  gate1432(.a(s_126), .O(gate413inter3));
  inv1  gate1433(.a(s_127), .O(gate413inter4));
  nand2 gate1434(.a(gate413inter4), .b(gate413inter3), .O(gate413inter5));
  nor2  gate1435(.a(gate413inter5), .b(gate413inter2), .O(gate413inter6));
  inv1  gate1436(.a(G27), .O(gate413inter7));
  inv1  gate1437(.a(G1114), .O(gate413inter8));
  nand2 gate1438(.a(gate413inter8), .b(gate413inter7), .O(gate413inter9));
  nand2 gate1439(.a(s_127), .b(gate413inter3), .O(gate413inter10));
  nor2  gate1440(.a(gate413inter10), .b(gate413inter9), .O(gate413inter11));
  nor2  gate1441(.a(gate413inter11), .b(gate413inter6), .O(gate413inter12));
  nand2 gate1442(.a(gate413inter12), .b(gate413inter1), .O(G1210));
nand2 gate414( .a(G28), .b(G1117), .O(G1213) );
nand2 gate415( .a(G29), .b(G1120), .O(G1216) );

  xor2  gate1891(.a(G1123), .b(G30), .O(gate416inter0));
  nand2 gate1892(.a(gate416inter0), .b(s_192), .O(gate416inter1));
  and2  gate1893(.a(G1123), .b(G30), .O(gate416inter2));
  inv1  gate1894(.a(s_192), .O(gate416inter3));
  inv1  gate1895(.a(s_193), .O(gate416inter4));
  nand2 gate1896(.a(gate416inter4), .b(gate416inter3), .O(gate416inter5));
  nor2  gate1897(.a(gate416inter5), .b(gate416inter2), .O(gate416inter6));
  inv1  gate1898(.a(G30), .O(gate416inter7));
  inv1  gate1899(.a(G1123), .O(gate416inter8));
  nand2 gate1900(.a(gate416inter8), .b(gate416inter7), .O(gate416inter9));
  nand2 gate1901(.a(s_193), .b(gate416inter3), .O(gate416inter10));
  nor2  gate1902(.a(gate416inter10), .b(gate416inter9), .O(gate416inter11));
  nor2  gate1903(.a(gate416inter11), .b(gate416inter6), .O(gate416inter12));
  nand2 gate1904(.a(gate416inter12), .b(gate416inter1), .O(G1219));
nand2 gate417( .a(G31), .b(G1126), .O(G1222) );

  xor2  gate1975(.a(G1129), .b(G32), .O(gate418inter0));
  nand2 gate1976(.a(gate418inter0), .b(s_204), .O(gate418inter1));
  and2  gate1977(.a(G1129), .b(G32), .O(gate418inter2));
  inv1  gate1978(.a(s_204), .O(gate418inter3));
  inv1  gate1979(.a(s_205), .O(gate418inter4));
  nand2 gate1980(.a(gate418inter4), .b(gate418inter3), .O(gate418inter5));
  nor2  gate1981(.a(gate418inter5), .b(gate418inter2), .O(gate418inter6));
  inv1  gate1982(.a(G32), .O(gate418inter7));
  inv1  gate1983(.a(G1129), .O(gate418inter8));
  nand2 gate1984(.a(gate418inter8), .b(gate418inter7), .O(gate418inter9));
  nand2 gate1985(.a(s_205), .b(gate418inter3), .O(gate418inter10));
  nor2  gate1986(.a(gate418inter10), .b(gate418inter9), .O(gate418inter11));
  nor2  gate1987(.a(gate418inter11), .b(gate418inter6), .O(gate418inter12));
  nand2 gate1988(.a(gate418inter12), .b(gate418inter1), .O(G1225));
nand2 gate419( .a(G1), .b(G1132), .O(G1228) );
nand2 gate420( .a(G1036), .b(G1132), .O(G1229) );

  xor2  gate729(.a(G1135), .b(G2), .O(gate421inter0));
  nand2 gate730(.a(gate421inter0), .b(s_26), .O(gate421inter1));
  and2  gate731(.a(G1135), .b(G2), .O(gate421inter2));
  inv1  gate732(.a(s_26), .O(gate421inter3));
  inv1  gate733(.a(s_27), .O(gate421inter4));
  nand2 gate734(.a(gate421inter4), .b(gate421inter3), .O(gate421inter5));
  nor2  gate735(.a(gate421inter5), .b(gate421inter2), .O(gate421inter6));
  inv1  gate736(.a(G2), .O(gate421inter7));
  inv1  gate737(.a(G1135), .O(gate421inter8));
  nand2 gate738(.a(gate421inter8), .b(gate421inter7), .O(gate421inter9));
  nand2 gate739(.a(s_27), .b(gate421inter3), .O(gate421inter10));
  nor2  gate740(.a(gate421inter10), .b(gate421inter9), .O(gate421inter11));
  nor2  gate741(.a(gate421inter11), .b(gate421inter6), .O(gate421inter12));
  nand2 gate742(.a(gate421inter12), .b(gate421inter1), .O(G1230));

  xor2  gate1821(.a(G1135), .b(G1039), .O(gate422inter0));
  nand2 gate1822(.a(gate422inter0), .b(s_182), .O(gate422inter1));
  and2  gate1823(.a(G1135), .b(G1039), .O(gate422inter2));
  inv1  gate1824(.a(s_182), .O(gate422inter3));
  inv1  gate1825(.a(s_183), .O(gate422inter4));
  nand2 gate1826(.a(gate422inter4), .b(gate422inter3), .O(gate422inter5));
  nor2  gate1827(.a(gate422inter5), .b(gate422inter2), .O(gate422inter6));
  inv1  gate1828(.a(G1039), .O(gate422inter7));
  inv1  gate1829(.a(G1135), .O(gate422inter8));
  nand2 gate1830(.a(gate422inter8), .b(gate422inter7), .O(gate422inter9));
  nand2 gate1831(.a(s_183), .b(gate422inter3), .O(gate422inter10));
  nor2  gate1832(.a(gate422inter10), .b(gate422inter9), .O(gate422inter11));
  nor2  gate1833(.a(gate422inter11), .b(gate422inter6), .O(gate422inter12));
  nand2 gate1834(.a(gate422inter12), .b(gate422inter1), .O(G1231));

  xor2  gate715(.a(G1138), .b(G3), .O(gate423inter0));
  nand2 gate716(.a(gate423inter0), .b(s_24), .O(gate423inter1));
  and2  gate717(.a(G1138), .b(G3), .O(gate423inter2));
  inv1  gate718(.a(s_24), .O(gate423inter3));
  inv1  gate719(.a(s_25), .O(gate423inter4));
  nand2 gate720(.a(gate423inter4), .b(gate423inter3), .O(gate423inter5));
  nor2  gate721(.a(gate423inter5), .b(gate423inter2), .O(gate423inter6));
  inv1  gate722(.a(G3), .O(gate423inter7));
  inv1  gate723(.a(G1138), .O(gate423inter8));
  nand2 gate724(.a(gate423inter8), .b(gate423inter7), .O(gate423inter9));
  nand2 gate725(.a(s_25), .b(gate423inter3), .O(gate423inter10));
  nor2  gate726(.a(gate423inter10), .b(gate423inter9), .O(gate423inter11));
  nor2  gate727(.a(gate423inter11), .b(gate423inter6), .O(gate423inter12));
  nand2 gate728(.a(gate423inter12), .b(gate423inter1), .O(G1232));
nand2 gate424( .a(G1042), .b(G1138), .O(G1233) );
nand2 gate425( .a(G4), .b(G1141), .O(G1234) );
nand2 gate426( .a(G1045), .b(G1141), .O(G1235) );

  xor2  gate2129(.a(G1144), .b(G5), .O(gate427inter0));
  nand2 gate2130(.a(gate427inter0), .b(s_226), .O(gate427inter1));
  and2  gate2131(.a(G1144), .b(G5), .O(gate427inter2));
  inv1  gate2132(.a(s_226), .O(gate427inter3));
  inv1  gate2133(.a(s_227), .O(gate427inter4));
  nand2 gate2134(.a(gate427inter4), .b(gate427inter3), .O(gate427inter5));
  nor2  gate2135(.a(gate427inter5), .b(gate427inter2), .O(gate427inter6));
  inv1  gate2136(.a(G5), .O(gate427inter7));
  inv1  gate2137(.a(G1144), .O(gate427inter8));
  nand2 gate2138(.a(gate427inter8), .b(gate427inter7), .O(gate427inter9));
  nand2 gate2139(.a(s_227), .b(gate427inter3), .O(gate427inter10));
  nor2  gate2140(.a(gate427inter10), .b(gate427inter9), .O(gate427inter11));
  nor2  gate2141(.a(gate427inter11), .b(gate427inter6), .O(gate427inter12));
  nand2 gate2142(.a(gate427inter12), .b(gate427inter1), .O(G1236));

  xor2  gate589(.a(G1144), .b(G1048), .O(gate428inter0));
  nand2 gate590(.a(gate428inter0), .b(s_6), .O(gate428inter1));
  and2  gate591(.a(G1144), .b(G1048), .O(gate428inter2));
  inv1  gate592(.a(s_6), .O(gate428inter3));
  inv1  gate593(.a(s_7), .O(gate428inter4));
  nand2 gate594(.a(gate428inter4), .b(gate428inter3), .O(gate428inter5));
  nor2  gate595(.a(gate428inter5), .b(gate428inter2), .O(gate428inter6));
  inv1  gate596(.a(G1048), .O(gate428inter7));
  inv1  gate597(.a(G1144), .O(gate428inter8));
  nand2 gate598(.a(gate428inter8), .b(gate428inter7), .O(gate428inter9));
  nand2 gate599(.a(s_7), .b(gate428inter3), .O(gate428inter10));
  nor2  gate600(.a(gate428inter10), .b(gate428inter9), .O(gate428inter11));
  nor2  gate601(.a(gate428inter11), .b(gate428inter6), .O(gate428inter12));
  nand2 gate602(.a(gate428inter12), .b(gate428inter1), .O(G1237));
nand2 gate429( .a(G6), .b(G1147), .O(G1238) );

  xor2  gate1415(.a(G1147), .b(G1051), .O(gate430inter0));
  nand2 gate1416(.a(gate430inter0), .b(s_124), .O(gate430inter1));
  and2  gate1417(.a(G1147), .b(G1051), .O(gate430inter2));
  inv1  gate1418(.a(s_124), .O(gate430inter3));
  inv1  gate1419(.a(s_125), .O(gate430inter4));
  nand2 gate1420(.a(gate430inter4), .b(gate430inter3), .O(gate430inter5));
  nor2  gate1421(.a(gate430inter5), .b(gate430inter2), .O(gate430inter6));
  inv1  gate1422(.a(G1051), .O(gate430inter7));
  inv1  gate1423(.a(G1147), .O(gate430inter8));
  nand2 gate1424(.a(gate430inter8), .b(gate430inter7), .O(gate430inter9));
  nand2 gate1425(.a(s_125), .b(gate430inter3), .O(gate430inter10));
  nor2  gate1426(.a(gate430inter10), .b(gate430inter9), .O(gate430inter11));
  nor2  gate1427(.a(gate430inter11), .b(gate430inter6), .O(gate430inter12));
  nand2 gate1428(.a(gate430inter12), .b(gate430inter1), .O(G1239));
nand2 gate431( .a(G7), .b(G1150), .O(G1240) );
nand2 gate432( .a(G1054), .b(G1150), .O(G1241) );
nand2 gate433( .a(G8), .b(G1153), .O(G1242) );

  xor2  gate617(.a(G1153), .b(G1057), .O(gate434inter0));
  nand2 gate618(.a(gate434inter0), .b(s_10), .O(gate434inter1));
  and2  gate619(.a(G1153), .b(G1057), .O(gate434inter2));
  inv1  gate620(.a(s_10), .O(gate434inter3));
  inv1  gate621(.a(s_11), .O(gate434inter4));
  nand2 gate622(.a(gate434inter4), .b(gate434inter3), .O(gate434inter5));
  nor2  gate623(.a(gate434inter5), .b(gate434inter2), .O(gate434inter6));
  inv1  gate624(.a(G1057), .O(gate434inter7));
  inv1  gate625(.a(G1153), .O(gate434inter8));
  nand2 gate626(.a(gate434inter8), .b(gate434inter7), .O(gate434inter9));
  nand2 gate627(.a(s_11), .b(gate434inter3), .O(gate434inter10));
  nor2  gate628(.a(gate434inter10), .b(gate434inter9), .O(gate434inter11));
  nor2  gate629(.a(gate434inter11), .b(gate434inter6), .O(gate434inter12));
  nand2 gate630(.a(gate434inter12), .b(gate434inter1), .O(G1243));
nand2 gate435( .a(G9), .b(G1156), .O(G1244) );
nand2 gate436( .a(G1060), .b(G1156), .O(G1245) );
nand2 gate437( .a(G10), .b(G1159), .O(G1246) );
nand2 gate438( .a(G1063), .b(G1159), .O(G1247) );

  xor2  gate1345(.a(G1162), .b(G11), .O(gate439inter0));
  nand2 gate1346(.a(gate439inter0), .b(s_114), .O(gate439inter1));
  and2  gate1347(.a(G1162), .b(G11), .O(gate439inter2));
  inv1  gate1348(.a(s_114), .O(gate439inter3));
  inv1  gate1349(.a(s_115), .O(gate439inter4));
  nand2 gate1350(.a(gate439inter4), .b(gate439inter3), .O(gate439inter5));
  nor2  gate1351(.a(gate439inter5), .b(gate439inter2), .O(gate439inter6));
  inv1  gate1352(.a(G11), .O(gate439inter7));
  inv1  gate1353(.a(G1162), .O(gate439inter8));
  nand2 gate1354(.a(gate439inter8), .b(gate439inter7), .O(gate439inter9));
  nand2 gate1355(.a(s_115), .b(gate439inter3), .O(gate439inter10));
  nor2  gate1356(.a(gate439inter10), .b(gate439inter9), .O(gate439inter11));
  nor2  gate1357(.a(gate439inter11), .b(gate439inter6), .O(gate439inter12));
  nand2 gate1358(.a(gate439inter12), .b(gate439inter1), .O(G1248));

  xor2  gate603(.a(G1162), .b(G1066), .O(gate440inter0));
  nand2 gate604(.a(gate440inter0), .b(s_8), .O(gate440inter1));
  and2  gate605(.a(G1162), .b(G1066), .O(gate440inter2));
  inv1  gate606(.a(s_8), .O(gate440inter3));
  inv1  gate607(.a(s_9), .O(gate440inter4));
  nand2 gate608(.a(gate440inter4), .b(gate440inter3), .O(gate440inter5));
  nor2  gate609(.a(gate440inter5), .b(gate440inter2), .O(gate440inter6));
  inv1  gate610(.a(G1066), .O(gate440inter7));
  inv1  gate611(.a(G1162), .O(gate440inter8));
  nand2 gate612(.a(gate440inter8), .b(gate440inter7), .O(gate440inter9));
  nand2 gate613(.a(s_9), .b(gate440inter3), .O(gate440inter10));
  nor2  gate614(.a(gate440inter10), .b(gate440inter9), .O(gate440inter11));
  nor2  gate615(.a(gate440inter11), .b(gate440inter6), .O(gate440inter12));
  nand2 gate616(.a(gate440inter12), .b(gate440inter1), .O(G1249));
nand2 gate441( .a(G12), .b(G1165), .O(G1250) );
nand2 gate442( .a(G1069), .b(G1165), .O(G1251) );
nand2 gate443( .a(G13), .b(G1168), .O(G1252) );
nand2 gate444( .a(G1072), .b(G1168), .O(G1253) );
nand2 gate445( .a(G14), .b(G1171), .O(G1254) );
nand2 gate446( .a(G1075), .b(G1171), .O(G1255) );
nand2 gate447( .a(G15), .b(G1174), .O(G1256) );
nand2 gate448( .a(G1078), .b(G1174), .O(G1257) );
nand2 gate449( .a(G16), .b(G1177), .O(G1258) );
nand2 gate450( .a(G1081), .b(G1177), .O(G1259) );
nand2 gate451( .a(G17), .b(G1180), .O(G1260) );
nand2 gate452( .a(G1084), .b(G1180), .O(G1261) );
nand2 gate453( .a(G18), .b(G1183), .O(G1262) );
nand2 gate454( .a(G1087), .b(G1183), .O(G1263) );

  xor2  gate1961(.a(G1186), .b(G19), .O(gate455inter0));
  nand2 gate1962(.a(gate455inter0), .b(s_202), .O(gate455inter1));
  and2  gate1963(.a(G1186), .b(G19), .O(gate455inter2));
  inv1  gate1964(.a(s_202), .O(gate455inter3));
  inv1  gate1965(.a(s_203), .O(gate455inter4));
  nand2 gate1966(.a(gate455inter4), .b(gate455inter3), .O(gate455inter5));
  nor2  gate1967(.a(gate455inter5), .b(gate455inter2), .O(gate455inter6));
  inv1  gate1968(.a(G19), .O(gate455inter7));
  inv1  gate1969(.a(G1186), .O(gate455inter8));
  nand2 gate1970(.a(gate455inter8), .b(gate455inter7), .O(gate455inter9));
  nand2 gate1971(.a(s_203), .b(gate455inter3), .O(gate455inter10));
  nor2  gate1972(.a(gate455inter10), .b(gate455inter9), .O(gate455inter11));
  nor2  gate1973(.a(gate455inter11), .b(gate455inter6), .O(gate455inter12));
  nand2 gate1974(.a(gate455inter12), .b(gate455inter1), .O(G1264));
nand2 gate456( .a(G1090), .b(G1186), .O(G1265) );
nand2 gate457( .a(G20), .b(G1189), .O(G1266) );
nand2 gate458( .a(G1093), .b(G1189), .O(G1267) );

  xor2  gate2143(.a(G1192), .b(G21), .O(gate459inter0));
  nand2 gate2144(.a(gate459inter0), .b(s_228), .O(gate459inter1));
  and2  gate2145(.a(G1192), .b(G21), .O(gate459inter2));
  inv1  gate2146(.a(s_228), .O(gate459inter3));
  inv1  gate2147(.a(s_229), .O(gate459inter4));
  nand2 gate2148(.a(gate459inter4), .b(gate459inter3), .O(gate459inter5));
  nor2  gate2149(.a(gate459inter5), .b(gate459inter2), .O(gate459inter6));
  inv1  gate2150(.a(G21), .O(gate459inter7));
  inv1  gate2151(.a(G1192), .O(gate459inter8));
  nand2 gate2152(.a(gate459inter8), .b(gate459inter7), .O(gate459inter9));
  nand2 gate2153(.a(s_229), .b(gate459inter3), .O(gate459inter10));
  nor2  gate2154(.a(gate459inter10), .b(gate459inter9), .O(gate459inter11));
  nor2  gate2155(.a(gate459inter11), .b(gate459inter6), .O(gate459inter12));
  nand2 gate2156(.a(gate459inter12), .b(gate459inter1), .O(G1268));
nand2 gate460( .a(G1096), .b(G1192), .O(G1269) );
nand2 gate461( .a(G22), .b(G1195), .O(G1270) );
nand2 gate462( .a(G1099), .b(G1195), .O(G1271) );
nand2 gate463( .a(G23), .b(G1198), .O(G1272) );
nand2 gate464( .a(G1102), .b(G1198), .O(G1273) );
nand2 gate465( .a(G24), .b(G1201), .O(G1274) );
nand2 gate466( .a(G1105), .b(G1201), .O(G1275) );
nand2 gate467( .a(G25), .b(G1204), .O(G1276) );
nand2 gate468( .a(G1108), .b(G1204), .O(G1277) );

  xor2  gate701(.a(G1207), .b(G26), .O(gate469inter0));
  nand2 gate702(.a(gate469inter0), .b(s_22), .O(gate469inter1));
  and2  gate703(.a(G1207), .b(G26), .O(gate469inter2));
  inv1  gate704(.a(s_22), .O(gate469inter3));
  inv1  gate705(.a(s_23), .O(gate469inter4));
  nand2 gate706(.a(gate469inter4), .b(gate469inter3), .O(gate469inter5));
  nor2  gate707(.a(gate469inter5), .b(gate469inter2), .O(gate469inter6));
  inv1  gate708(.a(G26), .O(gate469inter7));
  inv1  gate709(.a(G1207), .O(gate469inter8));
  nand2 gate710(.a(gate469inter8), .b(gate469inter7), .O(gate469inter9));
  nand2 gate711(.a(s_23), .b(gate469inter3), .O(gate469inter10));
  nor2  gate712(.a(gate469inter10), .b(gate469inter9), .O(gate469inter11));
  nor2  gate713(.a(gate469inter11), .b(gate469inter6), .O(gate469inter12));
  nand2 gate714(.a(gate469inter12), .b(gate469inter1), .O(G1278));
nand2 gate470( .a(G1111), .b(G1207), .O(G1279) );
nand2 gate471( .a(G27), .b(G1210), .O(G1280) );

  xor2  gate1331(.a(G1210), .b(G1114), .O(gate472inter0));
  nand2 gate1332(.a(gate472inter0), .b(s_112), .O(gate472inter1));
  and2  gate1333(.a(G1210), .b(G1114), .O(gate472inter2));
  inv1  gate1334(.a(s_112), .O(gate472inter3));
  inv1  gate1335(.a(s_113), .O(gate472inter4));
  nand2 gate1336(.a(gate472inter4), .b(gate472inter3), .O(gate472inter5));
  nor2  gate1337(.a(gate472inter5), .b(gate472inter2), .O(gate472inter6));
  inv1  gate1338(.a(G1114), .O(gate472inter7));
  inv1  gate1339(.a(G1210), .O(gate472inter8));
  nand2 gate1340(.a(gate472inter8), .b(gate472inter7), .O(gate472inter9));
  nand2 gate1341(.a(s_113), .b(gate472inter3), .O(gate472inter10));
  nor2  gate1342(.a(gate472inter10), .b(gate472inter9), .O(gate472inter11));
  nor2  gate1343(.a(gate472inter11), .b(gate472inter6), .O(gate472inter12));
  nand2 gate1344(.a(gate472inter12), .b(gate472inter1), .O(G1281));
nand2 gate473( .a(G28), .b(G1213), .O(G1282) );
nand2 gate474( .a(G1117), .b(G1213), .O(G1283) );

  xor2  gate1807(.a(G1216), .b(G29), .O(gate475inter0));
  nand2 gate1808(.a(gate475inter0), .b(s_180), .O(gate475inter1));
  and2  gate1809(.a(G1216), .b(G29), .O(gate475inter2));
  inv1  gate1810(.a(s_180), .O(gate475inter3));
  inv1  gate1811(.a(s_181), .O(gate475inter4));
  nand2 gate1812(.a(gate475inter4), .b(gate475inter3), .O(gate475inter5));
  nor2  gate1813(.a(gate475inter5), .b(gate475inter2), .O(gate475inter6));
  inv1  gate1814(.a(G29), .O(gate475inter7));
  inv1  gate1815(.a(G1216), .O(gate475inter8));
  nand2 gate1816(.a(gate475inter8), .b(gate475inter7), .O(gate475inter9));
  nand2 gate1817(.a(s_181), .b(gate475inter3), .O(gate475inter10));
  nor2  gate1818(.a(gate475inter10), .b(gate475inter9), .O(gate475inter11));
  nor2  gate1819(.a(gate475inter11), .b(gate475inter6), .O(gate475inter12));
  nand2 gate1820(.a(gate475inter12), .b(gate475inter1), .O(G1284));

  xor2  gate1765(.a(G1216), .b(G1120), .O(gate476inter0));
  nand2 gate1766(.a(gate476inter0), .b(s_174), .O(gate476inter1));
  and2  gate1767(.a(G1216), .b(G1120), .O(gate476inter2));
  inv1  gate1768(.a(s_174), .O(gate476inter3));
  inv1  gate1769(.a(s_175), .O(gate476inter4));
  nand2 gate1770(.a(gate476inter4), .b(gate476inter3), .O(gate476inter5));
  nor2  gate1771(.a(gate476inter5), .b(gate476inter2), .O(gate476inter6));
  inv1  gate1772(.a(G1120), .O(gate476inter7));
  inv1  gate1773(.a(G1216), .O(gate476inter8));
  nand2 gate1774(.a(gate476inter8), .b(gate476inter7), .O(gate476inter9));
  nand2 gate1775(.a(s_175), .b(gate476inter3), .O(gate476inter10));
  nor2  gate1776(.a(gate476inter10), .b(gate476inter9), .O(gate476inter11));
  nor2  gate1777(.a(gate476inter11), .b(gate476inter6), .O(gate476inter12));
  nand2 gate1778(.a(gate476inter12), .b(gate476inter1), .O(G1285));

  xor2  gate1919(.a(G1219), .b(G30), .O(gate477inter0));
  nand2 gate1920(.a(gate477inter0), .b(s_196), .O(gate477inter1));
  and2  gate1921(.a(G1219), .b(G30), .O(gate477inter2));
  inv1  gate1922(.a(s_196), .O(gate477inter3));
  inv1  gate1923(.a(s_197), .O(gate477inter4));
  nand2 gate1924(.a(gate477inter4), .b(gate477inter3), .O(gate477inter5));
  nor2  gate1925(.a(gate477inter5), .b(gate477inter2), .O(gate477inter6));
  inv1  gate1926(.a(G30), .O(gate477inter7));
  inv1  gate1927(.a(G1219), .O(gate477inter8));
  nand2 gate1928(.a(gate477inter8), .b(gate477inter7), .O(gate477inter9));
  nand2 gate1929(.a(s_197), .b(gate477inter3), .O(gate477inter10));
  nor2  gate1930(.a(gate477inter10), .b(gate477inter9), .O(gate477inter11));
  nor2  gate1931(.a(gate477inter11), .b(gate477inter6), .O(gate477inter12));
  nand2 gate1932(.a(gate477inter12), .b(gate477inter1), .O(G1286));
nand2 gate478( .a(G1123), .b(G1219), .O(G1287) );
nand2 gate479( .a(G31), .b(G1222), .O(G1288) );
nand2 gate480( .a(G1126), .b(G1222), .O(G1289) );
nand2 gate481( .a(G32), .b(G1225), .O(G1290) );
nand2 gate482( .a(G1129), .b(G1225), .O(G1291) );
nand2 gate483( .a(G1228), .b(G1229), .O(G1292) );
nand2 gate484( .a(G1230), .b(G1231), .O(G1293) );
nand2 gate485( .a(G1232), .b(G1233), .O(G1294) );

  xor2  gate1205(.a(G1235), .b(G1234), .O(gate486inter0));
  nand2 gate1206(.a(gate486inter0), .b(s_94), .O(gate486inter1));
  and2  gate1207(.a(G1235), .b(G1234), .O(gate486inter2));
  inv1  gate1208(.a(s_94), .O(gate486inter3));
  inv1  gate1209(.a(s_95), .O(gate486inter4));
  nand2 gate1210(.a(gate486inter4), .b(gate486inter3), .O(gate486inter5));
  nor2  gate1211(.a(gate486inter5), .b(gate486inter2), .O(gate486inter6));
  inv1  gate1212(.a(G1234), .O(gate486inter7));
  inv1  gate1213(.a(G1235), .O(gate486inter8));
  nand2 gate1214(.a(gate486inter8), .b(gate486inter7), .O(gate486inter9));
  nand2 gate1215(.a(s_95), .b(gate486inter3), .O(gate486inter10));
  nor2  gate1216(.a(gate486inter10), .b(gate486inter9), .O(gate486inter11));
  nor2  gate1217(.a(gate486inter11), .b(gate486inter6), .O(gate486inter12));
  nand2 gate1218(.a(gate486inter12), .b(gate486inter1), .O(G1295));
nand2 gate487( .a(G1236), .b(G1237), .O(G1296) );
nand2 gate488( .a(G1238), .b(G1239), .O(G1297) );
nand2 gate489( .a(G1240), .b(G1241), .O(G1298) );
nand2 gate490( .a(G1242), .b(G1243), .O(G1299) );

  xor2  gate1443(.a(G1245), .b(G1244), .O(gate491inter0));
  nand2 gate1444(.a(gate491inter0), .b(s_128), .O(gate491inter1));
  and2  gate1445(.a(G1245), .b(G1244), .O(gate491inter2));
  inv1  gate1446(.a(s_128), .O(gate491inter3));
  inv1  gate1447(.a(s_129), .O(gate491inter4));
  nand2 gate1448(.a(gate491inter4), .b(gate491inter3), .O(gate491inter5));
  nor2  gate1449(.a(gate491inter5), .b(gate491inter2), .O(gate491inter6));
  inv1  gate1450(.a(G1244), .O(gate491inter7));
  inv1  gate1451(.a(G1245), .O(gate491inter8));
  nand2 gate1452(.a(gate491inter8), .b(gate491inter7), .O(gate491inter9));
  nand2 gate1453(.a(s_129), .b(gate491inter3), .O(gate491inter10));
  nor2  gate1454(.a(gate491inter10), .b(gate491inter9), .O(gate491inter11));
  nor2  gate1455(.a(gate491inter11), .b(gate491inter6), .O(gate491inter12));
  nand2 gate1456(.a(gate491inter12), .b(gate491inter1), .O(G1300));
nand2 gate492( .a(G1246), .b(G1247), .O(G1301) );

  xor2  gate1541(.a(G1249), .b(G1248), .O(gate493inter0));
  nand2 gate1542(.a(gate493inter0), .b(s_142), .O(gate493inter1));
  and2  gate1543(.a(G1249), .b(G1248), .O(gate493inter2));
  inv1  gate1544(.a(s_142), .O(gate493inter3));
  inv1  gate1545(.a(s_143), .O(gate493inter4));
  nand2 gate1546(.a(gate493inter4), .b(gate493inter3), .O(gate493inter5));
  nor2  gate1547(.a(gate493inter5), .b(gate493inter2), .O(gate493inter6));
  inv1  gate1548(.a(G1248), .O(gate493inter7));
  inv1  gate1549(.a(G1249), .O(gate493inter8));
  nand2 gate1550(.a(gate493inter8), .b(gate493inter7), .O(gate493inter9));
  nand2 gate1551(.a(s_143), .b(gate493inter3), .O(gate493inter10));
  nor2  gate1552(.a(gate493inter10), .b(gate493inter9), .O(gate493inter11));
  nor2  gate1553(.a(gate493inter11), .b(gate493inter6), .O(gate493inter12));
  nand2 gate1554(.a(gate493inter12), .b(gate493inter1), .O(G1302));
nand2 gate494( .a(G1250), .b(G1251), .O(G1303) );
nand2 gate495( .a(G1252), .b(G1253), .O(G1304) );

  xor2  gate1905(.a(G1255), .b(G1254), .O(gate496inter0));
  nand2 gate1906(.a(gate496inter0), .b(s_194), .O(gate496inter1));
  and2  gate1907(.a(G1255), .b(G1254), .O(gate496inter2));
  inv1  gate1908(.a(s_194), .O(gate496inter3));
  inv1  gate1909(.a(s_195), .O(gate496inter4));
  nand2 gate1910(.a(gate496inter4), .b(gate496inter3), .O(gate496inter5));
  nor2  gate1911(.a(gate496inter5), .b(gate496inter2), .O(gate496inter6));
  inv1  gate1912(.a(G1254), .O(gate496inter7));
  inv1  gate1913(.a(G1255), .O(gate496inter8));
  nand2 gate1914(.a(gate496inter8), .b(gate496inter7), .O(gate496inter9));
  nand2 gate1915(.a(s_195), .b(gate496inter3), .O(gate496inter10));
  nor2  gate1916(.a(gate496inter10), .b(gate496inter9), .O(gate496inter11));
  nor2  gate1917(.a(gate496inter11), .b(gate496inter6), .O(gate496inter12));
  nand2 gate1918(.a(gate496inter12), .b(gate496inter1), .O(G1305));
nand2 gate497( .a(G1256), .b(G1257), .O(G1306) );
nand2 gate498( .a(G1258), .b(G1259), .O(G1307) );
nand2 gate499( .a(G1260), .b(G1261), .O(G1308) );
nand2 gate500( .a(G1262), .b(G1263), .O(G1309) );

  xor2  gate771(.a(G1265), .b(G1264), .O(gate501inter0));
  nand2 gate772(.a(gate501inter0), .b(s_32), .O(gate501inter1));
  and2  gate773(.a(G1265), .b(G1264), .O(gate501inter2));
  inv1  gate774(.a(s_32), .O(gate501inter3));
  inv1  gate775(.a(s_33), .O(gate501inter4));
  nand2 gate776(.a(gate501inter4), .b(gate501inter3), .O(gate501inter5));
  nor2  gate777(.a(gate501inter5), .b(gate501inter2), .O(gate501inter6));
  inv1  gate778(.a(G1264), .O(gate501inter7));
  inv1  gate779(.a(G1265), .O(gate501inter8));
  nand2 gate780(.a(gate501inter8), .b(gate501inter7), .O(gate501inter9));
  nand2 gate781(.a(s_33), .b(gate501inter3), .O(gate501inter10));
  nor2  gate782(.a(gate501inter10), .b(gate501inter9), .O(gate501inter11));
  nor2  gate783(.a(gate501inter11), .b(gate501inter6), .O(gate501inter12));
  nand2 gate784(.a(gate501inter12), .b(gate501inter1), .O(G1310));
nand2 gate502( .a(G1266), .b(G1267), .O(G1311) );
nand2 gate503( .a(G1268), .b(G1269), .O(G1312) );

  xor2  gate2017(.a(G1271), .b(G1270), .O(gate504inter0));
  nand2 gate2018(.a(gate504inter0), .b(s_210), .O(gate504inter1));
  and2  gate2019(.a(G1271), .b(G1270), .O(gate504inter2));
  inv1  gate2020(.a(s_210), .O(gate504inter3));
  inv1  gate2021(.a(s_211), .O(gate504inter4));
  nand2 gate2022(.a(gate504inter4), .b(gate504inter3), .O(gate504inter5));
  nor2  gate2023(.a(gate504inter5), .b(gate504inter2), .O(gate504inter6));
  inv1  gate2024(.a(G1270), .O(gate504inter7));
  inv1  gate2025(.a(G1271), .O(gate504inter8));
  nand2 gate2026(.a(gate504inter8), .b(gate504inter7), .O(gate504inter9));
  nand2 gate2027(.a(s_211), .b(gate504inter3), .O(gate504inter10));
  nor2  gate2028(.a(gate504inter10), .b(gate504inter9), .O(gate504inter11));
  nor2  gate2029(.a(gate504inter11), .b(gate504inter6), .O(gate504inter12));
  nand2 gate2030(.a(gate504inter12), .b(gate504inter1), .O(G1313));

  xor2  gate1597(.a(G1273), .b(G1272), .O(gate505inter0));
  nand2 gate1598(.a(gate505inter0), .b(s_150), .O(gate505inter1));
  and2  gate1599(.a(G1273), .b(G1272), .O(gate505inter2));
  inv1  gate1600(.a(s_150), .O(gate505inter3));
  inv1  gate1601(.a(s_151), .O(gate505inter4));
  nand2 gate1602(.a(gate505inter4), .b(gate505inter3), .O(gate505inter5));
  nor2  gate1603(.a(gate505inter5), .b(gate505inter2), .O(gate505inter6));
  inv1  gate1604(.a(G1272), .O(gate505inter7));
  inv1  gate1605(.a(G1273), .O(gate505inter8));
  nand2 gate1606(.a(gate505inter8), .b(gate505inter7), .O(gate505inter9));
  nand2 gate1607(.a(s_151), .b(gate505inter3), .O(gate505inter10));
  nor2  gate1608(.a(gate505inter10), .b(gate505inter9), .O(gate505inter11));
  nor2  gate1609(.a(gate505inter11), .b(gate505inter6), .O(gate505inter12));
  nand2 gate1610(.a(gate505inter12), .b(gate505inter1), .O(G1314));

  xor2  gate1303(.a(G1275), .b(G1274), .O(gate506inter0));
  nand2 gate1304(.a(gate506inter0), .b(s_108), .O(gate506inter1));
  and2  gate1305(.a(G1275), .b(G1274), .O(gate506inter2));
  inv1  gate1306(.a(s_108), .O(gate506inter3));
  inv1  gate1307(.a(s_109), .O(gate506inter4));
  nand2 gate1308(.a(gate506inter4), .b(gate506inter3), .O(gate506inter5));
  nor2  gate1309(.a(gate506inter5), .b(gate506inter2), .O(gate506inter6));
  inv1  gate1310(.a(G1274), .O(gate506inter7));
  inv1  gate1311(.a(G1275), .O(gate506inter8));
  nand2 gate1312(.a(gate506inter8), .b(gate506inter7), .O(gate506inter9));
  nand2 gate1313(.a(s_109), .b(gate506inter3), .O(gate506inter10));
  nor2  gate1314(.a(gate506inter10), .b(gate506inter9), .O(gate506inter11));
  nor2  gate1315(.a(gate506inter11), .b(gate506inter6), .O(gate506inter12));
  nand2 gate1316(.a(gate506inter12), .b(gate506inter1), .O(G1315));
nand2 gate507( .a(G1276), .b(G1277), .O(G1316) );
nand2 gate508( .a(G1278), .b(G1279), .O(G1317) );
nand2 gate509( .a(G1280), .b(G1281), .O(G1318) );
nand2 gate510( .a(G1282), .b(G1283), .O(G1319) );

  xor2  gate1261(.a(G1285), .b(G1284), .O(gate511inter0));
  nand2 gate1262(.a(gate511inter0), .b(s_102), .O(gate511inter1));
  and2  gate1263(.a(G1285), .b(G1284), .O(gate511inter2));
  inv1  gate1264(.a(s_102), .O(gate511inter3));
  inv1  gate1265(.a(s_103), .O(gate511inter4));
  nand2 gate1266(.a(gate511inter4), .b(gate511inter3), .O(gate511inter5));
  nor2  gate1267(.a(gate511inter5), .b(gate511inter2), .O(gate511inter6));
  inv1  gate1268(.a(G1284), .O(gate511inter7));
  inv1  gate1269(.a(G1285), .O(gate511inter8));
  nand2 gate1270(.a(gate511inter8), .b(gate511inter7), .O(gate511inter9));
  nand2 gate1271(.a(s_103), .b(gate511inter3), .O(gate511inter10));
  nor2  gate1272(.a(gate511inter10), .b(gate511inter9), .O(gate511inter11));
  nor2  gate1273(.a(gate511inter11), .b(gate511inter6), .O(gate511inter12));
  nand2 gate1274(.a(gate511inter12), .b(gate511inter1), .O(G1320));
nand2 gate512( .a(G1286), .b(G1287), .O(G1321) );

  xor2  gate813(.a(G1289), .b(G1288), .O(gate513inter0));
  nand2 gate814(.a(gate513inter0), .b(s_38), .O(gate513inter1));
  and2  gate815(.a(G1289), .b(G1288), .O(gate513inter2));
  inv1  gate816(.a(s_38), .O(gate513inter3));
  inv1  gate817(.a(s_39), .O(gate513inter4));
  nand2 gate818(.a(gate513inter4), .b(gate513inter3), .O(gate513inter5));
  nor2  gate819(.a(gate513inter5), .b(gate513inter2), .O(gate513inter6));
  inv1  gate820(.a(G1288), .O(gate513inter7));
  inv1  gate821(.a(G1289), .O(gate513inter8));
  nand2 gate822(.a(gate513inter8), .b(gate513inter7), .O(gate513inter9));
  nand2 gate823(.a(s_39), .b(gate513inter3), .O(gate513inter10));
  nor2  gate824(.a(gate513inter10), .b(gate513inter9), .O(gate513inter11));
  nor2  gate825(.a(gate513inter11), .b(gate513inter6), .O(gate513inter12));
  nand2 gate826(.a(gate513inter12), .b(gate513inter1), .O(G1322));

  xor2  gate1569(.a(G1291), .b(G1290), .O(gate514inter0));
  nand2 gate1570(.a(gate514inter0), .b(s_146), .O(gate514inter1));
  and2  gate1571(.a(G1291), .b(G1290), .O(gate514inter2));
  inv1  gate1572(.a(s_146), .O(gate514inter3));
  inv1  gate1573(.a(s_147), .O(gate514inter4));
  nand2 gate1574(.a(gate514inter4), .b(gate514inter3), .O(gate514inter5));
  nor2  gate1575(.a(gate514inter5), .b(gate514inter2), .O(gate514inter6));
  inv1  gate1576(.a(G1290), .O(gate514inter7));
  inv1  gate1577(.a(G1291), .O(gate514inter8));
  nand2 gate1578(.a(gate514inter8), .b(gate514inter7), .O(gate514inter9));
  nand2 gate1579(.a(s_147), .b(gate514inter3), .O(gate514inter10));
  nor2  gate1580(.a(gate514inter10), .b(gate514inter9), .O(gate514inter11));
  nor2  gate1581(.a(gate514inter11), .b(gate514inter6), .O(gate514inter12));
  nand2 gate1582(.a(gate514inter12), .b(gate514inter1), .O(G1323));
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule