module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);

input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;//RE__PI;

input s_0,s_1;//RE__ALLOW(00,01,10,11);
input s_2,s_3;//RE__ALLOW(00,01,10,11);
input s_4,s_5;//RE__ALLOW(00,01,10,11);
input s_6,s_7;//RE__ALLOW(00,01,10,11);
input s_8,s_9;//RE__ALLOW(00,01,10,11);
input s_10,s_11;//RE__ALLOW(00,01,10,11);
input s_12,s_13;//RE__ALLOW(00,01,10,11);
input s_14,s_15;//RE__ALLOW(00,01,10,11);
input s_16,s_17;//RE__ALLOW(00,01,10,11);
input s_18,s_19;//RE__ALLOW(00,01,10,11);
input s_20,s_21;//RE__ALLOW(00,01,10,11);
input s_22,s_23;//RE__ALLOW(00,01,10,11);
input s_24,s_25;//RE__ALLOW(00,01,10,11);
input s_26,s_27;//RE__ALLOW(00,01,10,11);
input s_28,s_29;//RE__ALLOW(00,01,10,11);
input s_30,s_31;//RE__ALLOW(00,01,10,11);
input s_32,s_33;//RE__ALLOW(00,01,10,11);
input s_34,s_35;//RE__ALLOW(00,01,10,11);
input s_36,s_37;//RE__ALLOW(00,01,10,11);
input s_38,s_39;//RE__ALLOW(00,01,10,11);
input s_40,s_41;//RE__ALLOW(00,01,10,11);
input s_42,s_43;//RE__ALLOW(00,01,10,11);
input s_44,s_45;//RE__ALLOW(00,01,10,11);
input s_46,s_47;//RE__ALLOW(00,01,10,11);
input s_48,s_49;//RE__ALLOW(00,01,10,11);
input s_50,s_51;//RE__ALLOW(00,01,10,11);
input s_52,s_53;//RE__ALLOW(00,01,10,11);
input s_54,s_55;//RE__ALLOW(00,01,10,11);
input s_56,s_57;//RE__ALLOW(00,01,10,11);
input s_58,s_59;//RE__ALLOW(00,01,10,11);
input s_60,s_61;//RE__ALLOW(00,01,10,11);
input s_62,s_63;//RE__ALLOW(00,01,10,11);
input s_64,s_65;//RE__ALLOW(00,01,10,11);
input s_66,s_67;//RE__ALLOW(00,01,10,11);
input s_68,s_69;//RE__ALLOW(00,01,10,11);
input s_70,s_71;//RE__ALLOW(00,01,10,11);
input s_72,s_73;//RE__ALLOW(00,01,10,11);
input s_74,s_75;//RE__ALLOW(00,01,10,11);
input s_76,s_77;//RE__ALLOW(00,01,10,11);
input s_78,s_79;//RE__ALLOW(00,01,10,11);
input s_80,s_81;//RE__ALLOW(00,01,10,11);
input s_82,s_83;//RE__ALLOW(00,01,10,11);
input s_84,s_85;//RE__ALLOW(00,01,10,11);
input s_86,s_87;//RE__ALLOW(00,01,10,11);
input s_88,s_89;//RE__ALLOW(00,01,10,11);
input s_90,s_91;//RE__ALLOW(00,01,10,11);
input s_92,s_93;//RE__ALLOW(00,01,10,11);
input s_94,s_95;//RE__ALLOW(00,01,10,11);
input s_96,s_97;//RE__ALLOW(00,01,10,11);
input s_98,s_99;//RE__ALLOW(00,01,10,11);
input s_100,s_101;//RE__ALLOW(00,01,10,11);
input s_102,s_103;//RE__ALLOW(00,01,10,11);
input s_104,s_105;//RE__ALLOW(00,01,10,11);
input s_106,s_107;//RE__ALLOW(00,01,10,11);
input s_108,s_109;//RE__ALLOW(00,01,10,11);
input s_110,s_111;//RE__ALLOW(00,01,10,11);
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;

  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate207inter0, gate207inter1, gate207inter2, gate207inter3, gate207inter4, gate207inter5, gate207inter6, gate207inter7, gate207inter8, gate207inter9, gate207inter10, gate207inter11, gate207inter12, gate13inter0, gate13inter1, gate13inter2, gate13inter3, gate13inter4, gate13inter5, gate13inter6, gate13inter7, gate13inter8, gate13inter9, gate13inter10, gate13inter11, gate13inter12, gate422inter0, gate422inter1, gate422inter2, gate422inter3, gate422inter4, gate422inter5, gate422inter6, gate422inter7, gate422inter8, gate422inter9, gate422inter10, gate422inter11, gate422inter12, gate428inter0, gate428inter1, gate428inter2, gate428inter3, gate428inter4, gate428inter5, gate428inter6, gate428inter7, gate428inter8, gate428inter9, gate428inter10, gate428inter11, gate428inter12, gate256inter0, gate256inter1, gate256inter2, gate256inter3, gate256inter4, gate256inter5, gate256inter6, gate256inter7, gate256inter8, gate256inter9, gate256inter10, gate256inter11, gate256inter12, gate113inter0, gate113inter1, gate113inter2, gate113inter3, gate113inter4, gate113inter5, gate113inter6, gate113inter7, gate113inter8, gate113inter9, gate113inter10, gate113inter11, gate113inter12, gate477inter0, gate477inter1, gate477inter2, gate477inter3, gate477inter4, gate477inter5, gate477inter6, gate477inter7, gate477inter8, gate477inter9, gate477inter10, gate477inter11, gate477inter12, gate211inter0, gate211inter1, gate211inter2, gate211inter3, gate211inter4, gate211inter5, gate211inter6, gate211inter7, gate211inter8, gate211inter9, gate211inter10, gate211inter11, gate211inter12, gate210inter0, gate210inter1, gate210inter2, gate210inter3, gate210inter4, gate210inter5, gate210inter6, gate210inter7, gate210inter8, gate210inter9, gate210inter10, gate210inter11, gate210inter12, gate390inter0, gate390inter1, gate390inter2, gate390inter3, gate390inter4, gate390inter5, gate390inter6, gate390inter7, gate390inter8, gate390inter9, gate390inter10, gate390inter11, gate390inter12, gate107inter0, gate107inter1, gate107inter2, gate107inter3, gate107inter4, gate107inter5, gate107inter6, gate107inter7, gate107inter8, gate107inter9, gate107inter10, gate107inter11, gate107inter12, gate41inter0, gate41inter1, gate41inter2, gate41inter3, gate41inter4, gate41inter5, gate41inter6, gate41inter7, gate41inter8, gate41inter9, gate41inter10, gate41inter11, gate41inter12, gate432inter0, gate432inter1, gate432inter2, gate432inter3, gate432inter4, gate432inter5, gate432inter6, gate432inter7, gate432inter8, gate432inter9, gate432inter10, gate432inter11, gate432inter12, gate449inter0, gate449inter1, gate449inter2, gate449inter3, gate449inter4, gate449inter5, gate449inter6, gate449inter7, gate449inter8, gate449inter9, gate449inter10, gate449inter11, gate449inter12, gate158inter0, gate158inter1, gate158inter2, gate158inter3, gate158inter4, gate158inter5, gate158inter6, gate158inter7, gate158inter8, gate158inter9, gate158inter10, gate158inter11, gate158inter12, gate412inter0, gate412inter1, gate412inter2, gate412inter3, gate412inter4, gate412inter5, gate412inter6, gate412inter7, gate412inter8, gate412inter9, gate412inter10, gate412inter11, gate412inter12, gate244inter0, gate244inter1, gate244inter2, gate244inter3, gate244inter4, gate244inter5, gate244inter6, gate244inter7, gate244inter8, gate244inter9, gate244inter10, gate244inter11, gate244inter12, gate75inter0, gate75inter1, gate75inter2, gate75inter3, gate75inter4, gate75inter5, gate75inter6, gate75inter7, gate75inter8, gate75inter9, gate75inter10, gate75inter11, gate75inter12, gate254inter0, gate254inter1, gate254inter2, gate254inter3, gate254inter4, gate254inter5, gate254inter6, gate254inter7, gate254inter8, gate254inter9, gate254inter10, gate254inter11, gate254inter12, gate235inter0, gate235inter1, gate235inter2, gate235inter3, gate235inter4, gate235inter5, gate235inter6, gate235inter7, gate235inter8, gate235inter9, gate235inter10, gate235inter11, gate235inter12, gate218inter0, gate218inter1, gate218inter2, gate218inter3, gate218inter4, gate218inter5, gate218inter6, gate218inter7, gate218inter8, gate218inter9, gate218inter10, gate218inter11, gate218inter12, gate169inter0, gate169inter1, gate169inter2, gate169inter3, gate169inter4, gate169inter5, gate169inter6, gate169inter7, gate169inter8, gate169inter9, gate169inter10, gate169inter11, gate169inter12, gate200inter0, gate200inter1, gate200inter2, gate200inter3, gate200inter4, gate200inter5, gate200inter6, gate200inter7, gate200inter8, gate200inter9, gate200inter10, gate200inter11, gate200inter12, gate53inter0, gate53inter1, gate53inter2, gate53inter3, gate53inter4, gate53inter5, gate53inter6, gate53inter7, gate53inter8, gate53inter9, gate53inter10, gate53inter11, gate53inter12, gate141inter0, gate141inter1, gate141inter2, gate141inter3, gate141inter4, gate141inter5, gate141inter6, gate141inter7, gate141inter8, gate141inter9, gate141inter10, gate141inter11, gate141inter12, gate9inter0, gate9inter1, gate9inter2, gate9inter3, gate9inter4, gate9inter5, gate9inter6, gate9inter7, gate9inter8, gate9inter9, gate9inter10, gate9inter11, gate9inter12, gate223inter0, gate223inter1, gate223inter2, gate223inter3, gate223inter4, gate223inter5, gate223inter6, gate223inter7, gate223inter8, gate223inter9, gate223inter10, gate223inter11, gate223inter12, gate151inter0, gate151inter1, gate151inter2, gate151inter3, gate151inter4, gate151inter5, gate151inter6, gate151inter7, gate151inter8, gate151inter9, gate151inter10, gate151inter11, gate151inter12, gate406inter0, gate406inter1, gate406inter2, gate406inter3, gate406inter4, gate406inter5, gate406inter6, gate406inter7, gate406inter8, gate406inter9, gate406inter10, gate406inter11, gate406inter12, gate508inter0, gate508inter1, gate508inter2, gate508inter3, gate508inter4, gate508inter5, gate508inter6, gate508inter7, gate508inter8, gate508inter9, gate508inter10, gate508inter11, gate508inter12, gate179inter0, gate179inter1, gate179inter2, gate179inter3, gate179inter4, gate179inter5, gate179inter6, gate179inter7, gate179inter8, gate179inter9, gate179inter10, gate179inter11, gate179inter12, gate185inter0, gate185inter1, gate185inter2, gate185inter3, gate185inter4, gate185inter5, gate185inter6, gate185inter7, gate185inter8, gate185inter9, gate185inter10, gate185inter11, gate185inter12, gate276inter0, gate276inter1, gate276inter2, gate276inter3, gate276inter4, gate276inter5, gate276inter6, gate276inter7, gate276inter8, gate276inter9, gate276inter10, gate276inter11, gate276inter12, gate282inter0, gate282inter1, gate282inter2, gate282inter3, gate282inter4, gate282inter5, gate282inter6, gate282inter7, gate282inter8, gate282inter9, gate282inter10, gate282inter11, gate282inter12, gate499inter0, gate499inter1, gate499inter2, gate499inter3, gate499inter4, gate499inter5, gate499inter6, gate499inter7, gate499inter8, gate499inter9, gate499inter10, gate499inter11, gate499inter12, gate140inter0, gate140inter1, gate140inter2, gate140inter3, gate140inter4, gate140inter5, gate140inter6, gate140inter7, gate140inter8, gate140inter9, gate140inter10, gate140inter11, gate140inter12, gate64inter0, gate64inter1, gate64inter2, gate64inter3, gate64inter4, gate64inter5, gate64inter6, gate64inter7, gate64inter8, gate64inter9, gate64inter10, gate64inter11, gate64inter12, gate471inter0, gate471inter1, gate471inter2, gate471inter3, gate471inter4, gate471inter5, gate471inter6, gate471inter7, gate471inter8, gate471inter9, gate471inter10, gate471inter11, gate471inter12, gate504inter0, gate504inter1, gate504inter2, gate504inter3, gate504inter4, gate504inter5, gate504inter6, gate504inter7, gate504inter8, gate504inter9, gate504inter10, gate504inter11, gate504inter12, gate97inter0, gate97inter1, gate97inter2, gate97inter3, gate97inter4, gate97inter5, gate97inter6, gate97inter7, gate97inter8, gate97inter9, gate97inter10, gate97inter11, gate97inter12, gate51inter0, gate51inter1, gate51inter2, gate51inter3, gate51inter4, gate51inter5, gate51inter6, gate51inter7, gate51inter8, gate51inter9, gate51inter10, gate51inter11, gate51inter12, gate461inter0, gate461inter1, gate461inter2, gate461inter3, gate461inter4, gate461inter5, gate461inter6, gate461inter7, gate461inter8, gate461inter9, gate461inter10, gate461inter11, gate461inter12, gate415inter0, gate415inter1, gate415inter2, gate415inter3, gate415inter4, gate415inter5, gate415inter6, gate415inter7, gate415inter8, gate415inter9, gate415inter10, gate415inter11, gate415inter12, gate72inter0, gate72inter1, gate72inter2, gate72inter3, gate72inter4, gate72inter5, gate72inter6, gate72inter7, gate72inter8, gate72inter9, gate72inter10, gate72inter11, gate72inter12, gate396inter0, gate396inter1, gate396inter2, gate396inter3, gate396inter4, gate396inter5, gate396inter6, gate396inter7, gate396inter8, gate396inter9, gate396inter10, gate396inter11, gate396inter12, gate233inter0, gate233inter1, gate233inter2, gate233inter3, gate233inter4, gate233inter5, gate233inter6, gate233inter7, gate233inter8, gate233inter9, gate233inter10, gate233inter11, gate233inter12, gate234inter0, gate234inter1, gate234inter2, gate234inter3, gate234inter4, gate234inter5, gate234inter6, gate234inter7, gate234inter8, gate234inter9, gate234inter10, gate234inter11, gate234inter12, gate405inter0, gate405inter1, gate405inter2, gate405inter3, gate405inter4, gate405inter5, gate405inter6, gate405inter7, gate405inter8, gate405inter9, gate405inter10, gate405inter11, gate405inter12, gate201inter0, gate201inter1, gate201inter2, gate201inter3, gate201inter4, gate201inter5, gate201inter6, gate201inter7, gate201inter8, gate201inter9, gate201inter10, gate201inter11, gate201inter12, gate164inter0, gate164inter1, gate164inter2, gate164inter3, gate164inter4, gate164inter5, gate164inter6, gate164inter7, gate164inter8, gate164inter9, gate164inter10, gate164inter11, gate164inter12, gate170inter0, gate170inter1, gate170inter2, gate170inter3, gate170inter4, gate170inter5, gate170inter6, gate170inter7, gate170inter8, gate170inter9, gate170inter10, gate170inter11, gate170inter12, gate498inter0, gate498inter1, gate498inter2, gate498inter3, gate498inter4, gate498inter5, gate498inter6, gate498inter7, gate498inter8, gate498inter9, gate498inter10, gate498inter11, gate498inter12, gate274inter0, gate274inter1, gate274inter2, gate274inter3, gate274inter4, gate274inter5, gate274inter6, gate274inter7, gate274inter8, gate274inter9, gate274inter10, gate274inter11, gate274inter12, gate38inter0, gate38inter1, gate38inter2, gate38inter3, gate38inter4, gate38inter5, gate38inter6, gate38inter7, gate38inter8, gate38inter9, gate38inter10, gate38inter11, gate38inter12, gate33inter0, gate33inter1, gate33inter2, gate33inter3, gate33inter4, gate33inter5, gate33inter6, gate33inter7, gate33inter8, gate33inter9, gate33inter10, gate33inter11, gate33inter12, gate495inter0, gate495inter1, gate495inter2, gate495inter3, gate495inter4, gate495inter5, gate495inter6, gate495inter7, gate495inter8, gate495inter9, gate495inter10, gate495inter11, gate495inter12;



and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );

  xor2  gate897(.a(G2), .b(G1), .O(gate9inter0));
  nand2 gate898(.a(gate9inter0), .b(s_50), .O(gate9inter1));
  and2  gate899(.a(G2), .b(G1), .O(gate9inter2));
  inv1  gate900(.a(s_50), .O(gate9inter3));
  inv1  gate901(.a(s_51), .O(gate9inter4));
  nand2 gate902(.a(gate9inter4), .b(gate9inter3), .O(gate9inter5));
  nor2  gate903(.a(gate9inter5), .b(gate9inter2), .O(gate9inter6));
  inv1  gate904(.a(G1), .O(gate9inter7));
  inv1  gate905(.a(G2), .O(gate9inter8));
  nand2 gate906(.a(gate9inter8), .b(gate9inter7), .O(gate9inter9));
  nand2 gate907(.a(s_51), .b(gate9inter3), .O(gate9inter10));
  nor2  gate908(.a(gate9inter10), .b(gate9inter9), .O(gate9inter11));
  nor2  gate909(.a(gate9inter11), .b(gate9inter6), .O(gate9inter12));
  nand2 gate910(.a(gate9inter12), .b(gate9inter1), .O(G266));
nand2 gate10( .a(G3), .b(G4), .O(G269) );
nand2 gate11( .a(G5), .b(G6), .O(G272) );
nand2 gate12( .a(G7), .b(G8), .O(G275) );

  xor2  gate561(.a(G10), .b(G9), .O(gate13inter0));
  nand2 gate562(.a(gate13inter0), .b(s_2), .O(gate13inter1));
  and2  gate563(.a(G10), .b(G9), .O(gate13inter2));
  inv1  gate564(.a(s_2), .O(gate13inter3));
  inv1  gate565(.a(s_3), .O(gate13inter4));
  nand2 gate566(.a(gate13inter4), .b(gate13inter3), .O(gate13inter5));
  nor2  gate567(.a(gate13inter5), .b(gate13inter2), .O(gate13inter6));
  inv1  gate568(.a(G9), .O(gate13inter7));
  inv1  gate569(.a(G10), .O(gate13inter8));
  nand2 gate570(.a(gate13inter8), .b(gate13inter7), .O(gate13inter9));
  nand2 gate571(.a(s_3), .b(gate13inter3), .O(gate13inter10));
  nor2  gate572(.a(gate13inter10), .b(gate13inter9), .O(gate13inter11));
  nor2  gate573(.a(gate13inter11), .b(gate13inter6), .O(gate13inter12));
  nand2 gate574(.a(gate13inter12), .b(gate13inter1), .O(G278));
nand2 gate14( .a(G11), .b(G12), .O(G281) );
nand2 gate15( .a(G13), .b(G14), .O(G284) );
nand2 gate16( .a(G15), .b(G16), .O(G287) );
nand2 gate17( .a(G17), .b(G18), .O(G290) );
nand2 gate18( .a(G19), .b(G20), .O(G293) );
nand2 gate19( .a(G21), .b(G22), .O(G296) );
nand2 gate20( .a(G23), .b(G24), .O(G299) );
nand2 gate21( .a(G25), .b(G26), .O(G302) );
nand2 gate22( .a(G27), .b(G28), .O(G305) );
nand2 gate23( .a(G29), .b(G30), .O(G308) );
nand2 gate24( .a(G31), .b(G32), .O(G311) );
nand2 gate25( .a(G1), .b(G5), .O(G314) );
nand2 gate26( .a(G9), .b(G13), .O(G317) );
nand2 gate27( .a(G2), .b(G6), .O(G320) );
nand2 gate28( .a(G10), .b(G14), .O(G323) );
nand2 gate29( .a(G3), .b(G7), .O(G326) );
nand2 gate30( .a(G11), .b(G15), .O(G329) );
nand2 gate31( .a(G4), .b(G8), .O(G332) );
nand2 gate32( .a(G12), .b(G16), .O(G335) );

  xor2  gate1303(.a(G21), .b(G17), .O(gate33inter0));
  nand2 gate1304(.a(gate33inter0), .b(s_108), .O(gate33inter1));
  and2  gate1305(.a(G21), .b(G17), .O(gate33inter2));
  inv1  gate1306(.a(s_108), .O(gate33inter3));
  inv1  gate1307(.a(s_109), .O(gate33inter4));
  nand2 gate1308(.a(gate33inter4), .b(gate33inter3), .O(gate33inter5));
  nor2  gate1309(.a(gate33inter5), .b(gate33inter2), .O(gate33inter6));
  inv1  gate1310(.a(G17), .O(gate33inter7));
  inv1  gate1311(.a(G21), .O(gate33inter8));
  nand2 gate1312(.a(gate33inter8), .b(gate33inter7), .O(gate33inter9));
  nand2 gate1313(.a(s_109), .b(gate33inter3), .O(gate33inter10));
  nor2  gate1314(.a(gate33inter10), .b(gate33inter9), .O(gate33inter11));
  nor2  gate1315(.a(gate33inter11), .b(gate33inter6), .O(gate33inter12));
  nand2 gate1316(.a(gate33inter12), .b(gate33inter1), .O(G338));
nand2 gate34( .a(G25), .b(G29), .O(G341) );
nand2 gate35( .a(G18), .b(G22), .O(G344) );
nand2 gate36( .a(G26), .b(G30), .O(G347) );
nand2 gate37( .a(G19), .b(G23), .O(G350) );

  xor2  gate1289(.a(G31), .b(G27), .O(gate38inter0));
  nand2 gate1290(.a(gate38inter0), .b(s_106), .O(gate38inter1));
  and2  gate1291(.a(G31), .b(G27), .O(gate38inter2));
  inv1  gate1292(.a(s_106), .O(gate38inter3));
  inv1  gate1293(.a(s_107), .O(gate38inter4));
  nand2 gate1294(.a(gate38inter4), .b(gate38inter3), .O(gate38inter5));
  nor2  gate1295(.a(gate38inter5), .b(gate38inter2), .O(gate38inter6));
  inv1  gate1296(.a(G27), .O(gate38inter7));
  inv1  gate1297(.a(G31), .O(gate38inter8));
  nand2 gate1298(.a(gate38inter8), .b(gate38inter7), .O(gate38inter9));
  nand2 gate1299(.a(s_107), .b(gate38inter3), .O(gate38inter10));
  nor2  gate1300(.a(gate38inter10), .b(gate38inter9), .O(gate38inter11));
  nor2  gate1301(.a(gate38inter11), .b(gate38inter6), .O(gate38inter12));
  nand2 gate1302(.a(gate38inter12), .b(gate38inter1), .O(G353));
nand2 gate39( .a(G20), .b(G24), .O(G356) );
nand2 gate40( .a(G28), .b(G32), .O(G359) );

  xor2  gate701(.a(G266), .b(G1), .O(gate41inter0));
  nand2 gate702(.a(gate41inter0), .b(s_22), .O(gate41inter1));
  and2  gate703(.a(G266), .b(G1), .O(gate41inter2));
  inv1  gate704(.a(s_22), .O(gate41inter3));
  inv1  gate705(.a(s_23), .O(gate41inter4));
  nand2 gate706(.a(gate41inter4), .b(gate41inter3), .O(gate41inter5));
  nor2  gate707(.a(gate41inter5), .b(gate41inter2), .O(gate41inter6));
  inv1  gate708(.a(G1), .O(gate41inter7));
  inv1  gate709(.a(G266), .O(gate41inter8));
  nand2 gate710(.a(gate41inter8), .b(gate41inter7), .O(gate41inter9));
  nand2 gate711(.a(s_23), .b(gate41inter3), .O(gate41inter10));
  nor2  gate712(.a(gate41inter10), .b(gate41inter9), .O(gate41inter11));
  nor2  gate713(.a(gate41inter11), .b(gate41inter6), .O(gate41inter12));
  nand2 gate714(.a(gate41inter12), .b(gate41inter1), .O(G362));
nand2 gate42( .a(G2), .b(G266), .O(G363) );
nand2 gate43( .a(G3), .b(G269), .O(G364) );
nand2 gate44( .a(G4), .b(G269), .O(G365) );
nand2 gate45( .a(G5), .b(G272), .O(G366) );
nand2 gate46( .a(G6), .b(G272), .O(G367) );
nand2 gate47( .a(G7), .b(G275), .O(G368) );
nand2 gate48( .a(G8), .b(G275), .O(G369) );
nand2 gate49( .a(G9), .b(G278), .O(G370) );
nand2 gate50( .a(G10), .b(G278), .O(G371) );

  xor2  gate1107(.a(G281), .b(G11), .O(gate51inter0));
  nand2 gate1108(.a(gate51inter0), .b(s_80), .O(gate51inter1));
  and2  gate1109(.a(G281), .b(G11), .O(gate51inter2));
  inv1  gate1110(.a(s_80), .O(gate51inter3));
  inv1  gate1111(.a(s_81), .O(gate51inter4));
  nand2 gate1112(.a(gate51inter4), .b(gate51inter3), .O(gate51inter5));
  nor2  gate1113(.a(gate51inter5), .b(gate51inter2), .O(gate51inter6));
  inv1  gate1114(.a(G11), .O(gate51inter7));
  inv1  gate1115(.a(G281), .O(gate51inter8));
  nand2 gate1116(.a(gate51inter8), .b(gate51inter7), .O(gate51inter9));
  nand2 gate1117(.a(s_81), .b(gate51inter3), .O(gate51inter10));
  nor2  gate1118(.a(gate51inter10), .b(gate51inter9), .O(gate51inter11));
  nor2  gate1119(.a(gate51inter11), .b(gate51inter6), .O(gate51inter12));
  nand2 gate1120(.a(gate51inter12), .b(gate51inter1), .O(G372));
nand2 gate52( .a(G12), .b(G281), .O(G373) );

  xor2  gate869(.a(G284), .b(G13), .O(gate53inter0));
  nand2 gate870(.a(gate53inter0), .b(s_46), .O(gate53inter1));
  and2  gate871(.a(G284), .b(G13), .O(gate53inter2));
  inv1  gate872(.a(s_46), .O(gate53inter3));
  inv1  gate873(.a(s_47), .O(gate53inter4));
  nand2 gate874(.a(gate53inter4), .b(gate53inter3), .O(gate53inter5));
  nor2  gate875(.a(gate53inter5), .b(gate53inter2), .O(gate53inter6));
  inv1  gate876(.a(G13), .O(gate53inter7));
  inv1  gate877(.a(G284), .O(gate53inter8));
  nand2 gate878(.a(gate53inter8), .b(gate53inter7), .O(gate53inter9));
  nand2 gate879(.a(s_47), .b(gate53inter3), .O(gate53inter10));
  nor2  gate880(.a(gate53inter10), .b(gate53inter9), .O(gate53inter11));
  nor2  gate881(.a(gate53inter11), .b(gate53inter6), .O(gate53inter12));
  nand2 gate882(.a(gate53inter12), .b(gate53inter1), .O(G374));
nand2 gate54( .a(G14), .b(G284), .O(G375) );
nand2 gate55( .a(G15), .b(G287), .O(G376) );
nand2 gate56( .a(G16), .b(G287), .O(G377) );
nand2 gate57( .a(G17), .b(G290), .O(G378) );
nand2 gate58( .a(G18), .b(G290), .O(G379) );
nand2 gate59( .a(G19), .b(G293), .O(G380) );
nand2 gate60( .a(G20), .b(G293), .O(G381) );
nand2 gate61( .a(G21), .b(G296), .O(G382) );
nand2 gate62( .a(G22), .b(G296), .O(G383) );
nand2 gate63( .a(G23), .b(G299), .O(G384) );

  xor2  gate1051(.a(G299), .b(G24), .O(gate64inter0));
  nand2 gate1052(.a(gate64inter0), .b(s_72), .O(gate64inter1));
  and2  gate1053(.a(G299), .b(G24), .O(gate64inter2));
  inv1  gate1054(.a(s_72), .O(gate64inter3));
  inv1  gate1055(.a(s_73), .O(gate64inter4));
  nand2 gate1056(.a(gate64inter4), .b(gate64inter3), .O(gate64inter5));
  nor2  gate1057(.a(gate64inter5), .b(gate64inter2), .O(gate64inter6));
  inv1  gate1058(.a(G24), .O(gate64inter7));
  inv1  gate1059(.a(G299), .O(gate64inter8));
  nand2 gate1060(.a(gate64inter8), .b(gate64inter7), .O(gate64inter9));
  nand2 gate1061(.a(s_73), .b(gate64inter3), .O(gate64inter10));
  nor2  gate1062(.a(gate64inter10), .b(gate64inter9), .O(gate64inter11));
  nor2  gate1063(.a(gate64inter11), .b(gate64inter6), .O(gate64inter12));
  nand2 gate1064(.a(gate64inter12), .b(gate64inter1), .O(G385));
nand2 gate65( .a(G25), .b(G302), .O(G386) );
nand2 gate66( .a(G26), .b(G302), .O(G387) );
nand2 gate67( .a(G27), .b(G305), .O(G388) );
nand2 gate68( .a(G28), .b(G305), .O(G389) );
nand2 gate69( .a(G29), .b(G308), .O(G390) );
nand2 gate70( .a(G30), .b(G308), .O(G391) );
nand2 gate71( .a(G31), .b(G311), .O(G392) );

  xor2  gate1149(.a(G311), .b(G32), .O(gate72inter0));
  nand2 gate1150(.a(gate72inter0), .b(s_86), .O(gate72inter1));
  and2  gate1151(.a(G311), .b(G32), .O(gate72inter2));
  inv1  gate1152(.a(s_86), .O(gate72inter3));
  inv1  gate1153(.a(s_87), .O(gate72inter4));
  nand2 gate1154(.a(gate72inter4), .b(gate72inter3), .O(gate72inter5));
  nor2  gate1155(.a(gate72inter5), .b(gate72inter2), .O(gate72inter6));
  inv1  gate1156(.a(G32), .O(gate72inter7));
  inv1  gate1157(.a(G311), .O(gate72inter8));
  nand2 gate1158(.a(gate72inter8), .b(gate72inter7), .O(gate72inter9));
  nand2 gate1159(.a(s_87), .b(gate72inter3), .O(gate72inter10));
  nor2  gate1160(.a(gate72inter10), .b(gate72inter9), .O(gate72inter11));
  nor2  gate1161(.a(gate72inter11), .b(gate72inter6), .O(gate72inter12));
  nand2 gate1162(.a(gate72inter12), .b(gate72inter1), .O(G393));
nand2 gate73( .a(G1), .b(G314), .O(G394) );
nand2 gate74( .a(G5), .b(G314), .O(G395) );

  xor2  gate785(.a(G317), .b(G9), .O(gate75inter0));
  nand2 gate786(.a(gate75inter0), .b(s_34), .O(gate75inter1));
  and2  gate787(.a(G317), .b(G9), .O(gate75inter2));
  inv1  gate788(.a(s_34), .O(gate75inter3));
  inv1  gate789(.a(s_35), .O(gate75inter4));
  nand2 gate790(.a(gate75inter4), .b(gate75inter3), .O(gate75inter5));
  nor2  gate791(.a(gate75inter5), .b(gate75inter2), .O(gate75inter6));
  inv1  gate792(.a(G9), .O(gate75inter7));
  inv1  gate793(.a(G317), .O(gate75inter8));
  nand2 gate794(.a(gate75inter8), .b(gate75inter7), .O(gate75inter9));
  nand2 gate795(.a(s_35), .b(gate75inter3), .O(gate75inter10));
  nor2  gate796(.a(gate75inter10), .b(gate75inter9), .O(gate75inter11));
  nor2  gate797(.a(gate75inter11), .b(gate75inter6), .O(gate75inter12));
  nand2 gate798(.a(gate75inter12), .b(gate75inter1), .O(G396));
nand2 gate76( .a(G13), .b(G317), .O(G397) );
nand2 gate77( .a(G2), .b(G320), .O(G398) );
nand2 gate78( .a(G6), .b(G320), .O(G399) );
nand2 gate79( .a(G10), .b(G323), .O(G400) );
nand2 gate80( .a(G14), .b(G323), .O(G401) );
nand2 gate81( .a(G3), .b(G326), .O(G402) );
nand2 gate82( .a(G7), .b(G326), .O(G403) );
nand2 gate83( .a(G11), .b(G329), .O(G404) );
nand2 gate84( .a(G15), .b(G329), .O(G405) );
nand2 gate85( .a(G4), .b(G332), .O(G406) );
nand2 gate86( .a(G8), .b(G332), .O(G407) );
nand2 gate87( .a(G12), .b(G335), .O(G408) );
nand2 gate88( .a(G16), .b(G335), .O(G409) );
nand2 gate89( .a(G17), .b(G338), .O(G410) );
nand2 gate90( .a(G21), .b(G338), .O(G411) );
nand2 gate91( .a(G25), .b(G341), .O(G412) );
nand2 gate92( .a(G29), .b(G341), .O(G413) );
nand2 gate93( .a(G18), .b(G344), .O(G414) );
nand2 gate94( .a(G22), .b(G344), .O(G415) );
nand2 gate95( .a(G26), .b(G347), .O(G416) );
nand2 gate96( .a(G30), .b(G347), .O(G417) );

  xor2  gate1093(.a(G350), .b(G19), .O(gate97inter0));
  nand2 gate1094(.a(gate97inter0), .b(s_78), .O(gate97inter1));
  and2  gate1095(.a(G350), .b(G19), .O(gate97inter2));
  inv1  gate1096(.a(s_78), .O(gate97inter3));
  inv1  gate1097(.a(s_79), .O(gate97inter4));
  nand2 gate1098(.a(gate97inter4), .b(gate97inter3), .O(gate97inter5));
  nor2  gate1099(.a(gate97inter5), .b(gate97inter2), .O(gate97inter6));
  inv1  gate1100(.a(G19), .O(gate97inter7));
  inv1  gate1101(.a(G350), .O(gate97inter8));
  nand2 gate1102(.a(gate97inter8), .b(gate97inter7), .O(gate97inter9));
  nand2 gate1103(.a(s_79), .b(gate97inter3), .O(gate97inter10));
  nor2  gate1104(.a(gate97inter10), .b(gate97inter9), .O(gate97inter11));
  nor2  gate1105(.a(gate97inter11), .b(gate97inter6), .O(gate97inter12));
  nand2 gate1106(.a(gate97inter12), .b(gate97inter1), .O(G418));
nand2 gate98( .a(G23), .b(G350), .O(G419) );
nand2 gate99( .a(G27), .b(G353), .O(G420) );
nand2 gate100( .a(G31), .b(G353), .O(G421) );
nand2 gate101( .a(G20), .b(G356), .O(G422) );
nand2 gate102( .a(G24), .b(G356), .O(G423) );
nand2 gate103( .a(G28), .b(G359), .O(G424) );
nand2 gate104( .a(G32), .b(G359), .O(G425) );
nand2 gate105( .a(G362), .b(G363), .O(G426) );
nand2 gate106( .a(G364), .b(G365), .O(G429) );

  xor2  gate687(.a(G367), .b(G366), .O(gate107inter0));
  nand2 gate688(.a(gate107inter0), .b(s_20), .O(gate107inter1));
  and2  gate689(.a(G367), .b(G366), .O(gate107inter2));
  inv1  gate690(.a(s_20), .O(gate107inter3));
  inv1  gate691(.a(s_21), .O(gate107inter4));
  nand2 gate692(.a(gate107inter4), .b(gate107inter3), .O(gate107inter5));
  nor2  gate693(.a(gate107inter5), .b(gate107inter2), .O(gate107inter6));
  inv1  gate694(.a(G366), .O(gate107inter7));
  inv1  gate695(.a(G367), .O(gate107inter8));
  nand2 gate696(.a(gate107inter8), .b(gate107inter7), .O(gate107inter9));
  nand2 gate697(.a(s_21), .b(gate107inter3), .O(gate107inter10));
  nor2  gate698(.a(gate107inter10), .b(gate107inter9), .O(gate107inter11));
  nor2  gate699(.a(gate107inter11), .b(gate107inter6), .O(gate107inter12));
  nand2 gate700(.a(gate107inter12), .b(gate107inter1), .O(G432));
nand2 gate108( .a(G368), .b(G369), .O(G435) );
nand2 gate109( .a(G370), .b(G371), .O(G438) );
nand2 gate110( .a(G372), .b(G373), .O(G441) );
nand2 gate111( .a(G374), .b(G375), .O(G444) );
nand2 gate112( .a(G376), .b(G377), .O(G447) );

  xor2  gate617(.a(G379), .b(G378), .O(gate113inter0));
  nand2 gate618(.a(gate113inter0), .b(s_10), .O(gate113inter1));
  and2  gate619(.a(G379), .b(G378), .O(gate113inter2));
  inv1  gate620(.a(s_10), .O(gate113inter3));
  inv1  gate621(.a(s_11), .O(gate113inter4));
  nand2 gate622(.a(gate113inter4), .b(gate113inter3), .O(gate113inter5));
  nor2  gate623(.a(gate113inter5), .b(gate113inter2), .O(gate113inter6));
  inv1  gate624(.a(G378), .O(gate113inter7));
  inv1  gate625(.a(G379), .O(gate113inter8));
  nand2 gate626(.a(gate113inter8), .b(gate113inter7), .O(gate113inter9));
  nand2 gate627(.a(s_11), .b(gate113inter3), .O(gate113inter10));
  nor2  gate628(.a(gate113inter10), .b(gate113inter9), .O(gate113inter11));
  nor2  gate629(.a(gate113inter11), .b(gate113inter6), .O(gate113inter12));
  nand2 gate630(.a(gate113inter12), .b(gate113inter1), .O(G450));
nand2 gate114( .a(G380), .b(G381), .O(G453) );
nand2 gate115( .a(G382), .b(G383), .O(G456) );
nand2 gate116( .a(G384), .b(G385), .O(G459) );
nand2 gate117( .a(G386), .b(G387), .O(G462) );
nand2 gate118( .a(G388), .b(G389), .O(G465) );
nand2 gate119( .a(G390), .b(G391), .O(G468) );
nand2 gate120( .a(G392), .b(G393), .O(G471) );
nand2 gate121( .a(G394), .b(G395), .O(G474) );
nand2 gate122( .a(G396), .b(G397), .O(G477) );
nand2 gate123( .a(G398), .b(G399), .O(G480) );
nand2 gate124( .a(G400), .b(G401), .O(G483) );
nand2 gate125( .a(G402), .b(G403), .O(G486) );
nand2 gate126( .a(G404), .b(G405), .O(G489) );
nand2 gate127( .a(G406), .b(G407), .O(G492) );
nand2 gate128( .a(G408), .b(G409), .O(G495) );
nand2 gate129( .a(G410), .b(G411), .O(G498) );
nand2 gate130( .a(G412), .b(G413), .O(G501) );
nand2 gate131( .a(G414), .b(G415), .O(G504) );
nand2 gate132( .a(G416), .b(G417), .O(G507) );
nand2 gate133( .a(G418), .b(G419), .O(G510) );
nand2 gate134( .a(G420), .b(G421), .O(G513) );
nand2 gate135( .a(G422), .b(G423), .O(G516) );
nand2 gate136( .a(G424), .b(G425), .O(G519) );
nand2 gate137( .a(G426), .b(G429), .O(G522) );
nand2 gate138( .a(G432), .b(G435), .O(G525) );
nand2 gate139( .a(G438), .b(G441), .O(G528) );

  xor2  gate1037(.a(G447), .b(G444), .O(gate140inter0));
  nand2 gate1038(.a(gate140inter0), .b(s_70), .O(gate140inter1));
  and2  gate1039(.a(G447), .b(G444), .O(gate140inter2));
  inv1  gate1040(.a(s_70), .O(gate140inter3));
  inv1  gate1041(.a(s_71), .O(gate140inter4));
  nand2 gate1042(.a(gate140inter4), .b(gate140inter3), .O(gate140inter5));
  nor2  gate1043(.a(gate140inter5), .b(gate140inter2), .O(gate140inter6));
  inv1  gate1044(.a(G444), .O(gate140inter7));
  inv1  gate1045(.a(G447), .O(gate140inter8));
  nand2 gate1046(.a(gate140inter8), .b(gate140inter7), .O(gate140inter9));
  nand2 gate1047(.a(s_71), .b(gate140inter3), .O(gate140inter10));
  nor2  gate1048(.a(gate140inter10), .b(gate140inter9), .O(gate140inter11));
  nor2  gate1049(.a(gate140inter11), .b(gate140inter6), .O(gate140inter12));
  nand2 gate1050(.a(gate140inter12), .b(gate140inter1), .O(G531));

  xor2  gate883(.a(G453), .b(G450), .O(gate141inter0));
  nand2 gate884(.a(gate141inter0), .b(s_48), .O(gate141inter1));
  and2  gate885(.a(G453), .b(G450), .O(gate141inter2));
  inv1  gate886(.a(s_48), .O(gate141inter3));
  inv1  gate887(.a(s_49), .O(gate141inter4));
  nand2 gate888(.a(gate141inter4), .b(gate141inter3), .O(gate141inter5));
  nor2  gate889(.a(gate141inter5), .b(gate141inter2), .O(gate141inter6));
  inv1  gate890(.a(G450), .O(gate141inter7));
  inv1  gate891(.a(G453), .O(gate141inter8));
  nand2 gate892(.a(gate141inter8), .b(gate141inter7), .O(gate141inter9));
  nand2 gate893(.a(s_49), .b(gate141inter3), .O(gate141inter10));
  nor2  gate894(.a(gate141inter10), .b(gate141inter9), .O(gate141inter11));
  nor2  gate895(.a(gate141inter11), .b(gate141inter6), .O(gate141inter12));
  nand2 gate896(.a(gate141inter12), .b(gate141inter1), .O(G534));
nand2 gate142( .a(G456), .b(G459), .O(G537) );
nand2 gate143( .a(G462), .b(G465), .O(G540) );
nand2 gate144( .a(G468), .b(G471), .O(G543) );
nand2 gate145( .a(G474), .b(G477), .O(G546) );
nand2 gate146( .a(G480), .b(G483), .O(G549) );
nand2 gate147( .a(G486), .b(G489), .O(G552) );
nand2 gate148( .a(G492), .b(G495), .O(G555) );
nand2 gate149( .a(G498), .b(G501), .O(G558) );
nand2 gate150( .a(G504), .b(G507), .O(G561) );

  xor2  gate925(.a(G513), .b(G510), .O(gate151inter0));
  nand2 gate926(.a(gate151inter0), .b(s_54), .O(gate151inter1));
  and2  gate927(.a(G513), .b(G510), .O(gate151inter2));
  inv1  gate928(.a(s_54), .O(gate151inter3));
  inv1  gate929(.a(s_55), .O(gate151inter4));
  nand2 gate930(.a(gate151inter4), .b(gate151inter3), .O(gate151inter5));
  nor2  gate931(.a(gate151inter5), .b(gate151inter2), .O(gate151inter6));
  inv1  gate932(.a(G510), .O(gate151inter7));
  inv1  gate933(.a(G513), .O(gate151inter8));
  nand2 gate934(.a(gate151inter8), .b(gate151inter7), .O(gate151inter9));
  nand2 gate935(.a(s_55), .b(gate151inter3), .O(gate151inter10));
  nor2  gate936(.a(gate151inter10), .b(gate151inter9), .O(gate151inter11));
  nor2  gate937(.a(gate151inter11), .b(gate151inter6), .O(gate151inter12));
  nand2 gate938(.a(gate151inter12), .b(gate151inter1), .O(G564));
nand2 gate152( .a(G516), .b(G519), .O(G567) );
nand2 gate153( .a(G426), .b(G522), .O(G570) );
nand2 gate154( .a(G429), .b(G522), .O(G571) );
nand2 gate155( .a(G432), .b(G525), .O(G572) );
nand2 gate156( .a(G435), .b(G525), .O(G573) );
nand2 gate157( .a(G438), .b(G528), .O(G574) );

  xor2  gate743(.a(G528), .b(G441), .O(gate158inter0));
  nand2 gate744(.a(gate158inter0), .b(s_28), .O(gate158inter1));
  and2  gate745(.a(G528), .b(G441), .O(gate158inter2));
  inv1  gate746(.a(s_28), .O(gate158inter3));
  inv1  gate747(.a(s_29), .O(gate158inter4));
  nand2 gate748(.a(gate158inter4), .b(gate158inter3), .O(gate158inter5));
  nor2  gate749(.a(gate158inter5), .b(gate158inter2), .O(gate158inter6));
  inv1  gate750(.a(G441), .O(gate158inter7));
  inv1  gate751(.a(G528), .O(gate158inter8));
  nand2 gate752(.a(gate158inter8), .b(gate158inter7), .O(gate158inter9));
  nand2 gate753(.a(s_29), .b(gate158inter3), .O(gate158inter10));
  nor2  gate754(.a(gate158inter10), .b(gate158inter9), .O(gate158inter11));
  nor2  gate755(.a(gate158inter11), .b(gate158inter6), .O(gate158inter12));
  nand2 gate756(.a(gate158inter12), .b(gate158inter1), .O(G575));
nand2 gate159( .a(G444), .b(G531), .O(G576) );
nand2 gate160( .a(G447), .b(G531), .O(G577) );
nand2 gate161( .a(G450), .b(G534), .O(G578) );
nand2 gate162( .a(G453), .b(G534), .O(G579) );
nand2 gate163( .a(G456), .b(G537), .O(G580) );

  xor2  gate1233(.a(G537), .b(G459), .O(gate164inter0));
  nand2 gate1234(.a(gate164inter0), .b(s_98), .O(gate164inter1));
  and2  gate1235(.a(G537), .b(G459), .O(gate164inter2));
  inv1  gate1236(.a(s_98), .O(gate164inter3));
  inv1  gate1237(.a(s_99), .O(gate164inter4));
  nand2 gate1238(.a(gate164inter4), .b(gate164inter3), .O(gate164inter5));
  nor2  gate1239(.a(gate164inter5), .b(gate164inter2), .O(gate164inter6));
  inv1  gate1240(.a(G459), .O(gate164inter7));
  inv1  gate1241(.a(G537), .O(gate164inter8));
  nand2 gate1242(.a(gate164inter8), .b(gate164inter7), .O(gate164inter9));
  nand2 gate1243(.a(s_99), .b(gate164inter3), .O(gate164inter10));
  nor2  gate1244(.a(gate164inter10), .b(gate164inter9), .O(gate164inter11));
  nor2  gate1245(.a(gate164inter11), .b(gate164inter6), .O(gate164inter12));
  nand2 gate1246(.a(gate164inter12), .b(gate164inter1), .O(G581));
nand2 gate165( .a(G462), .b(G540), .O(G582) );
nand2 gate166( .a(G465), .b(G540), .O(G583) );
nand2 gate167( .a(G468), .b(G543), .O(G584) );
nand2 gate168( .a(G471), .b(G543), .O(G585) );

  xor2  gate841(.a(G546), .b(G474), .O(gate169inter0));
  nand2 gate842(.a(gate169inter0), .b(s_42), .O(gate169inter1));
  and2  gate843(.a(G546), .b(G474), .O(gate169inter2));
  inv1  gate844(.a(s_42), .O(gate169inter3));
  inv1  gate845(.a(s_43), .O(gate169inter4));
  nand2 gate846(.a(gate169inter4), .b(gate169inter3), .O(gate169inter5));
  nor2  gate847(.a(gate169inter5), .b(gate169inter2), .O(gate169inter6));
  inv1  gate848(.a(G474), .O(gate169inter7));
  inv1  gate849(.a(G546), .O(gate169inter8));
  nand2 gate850(.a(gate169inter8), .b(gate169inter7), .O(gate169inter9));
  nand2 gate851(.a(s_43), .b(gate169inter3), .O(gate169inter10));
  nor2  gate852(.a(gate169inter10), .b(gate169inter9), .O(gate169inter11));
  nor2  gate853(.a(gate169inter11), .b(gate169inter6), .O(gate169inter12));
  nand2 gate854(.a(gate169inter12), .b(gate169inter1), .O(G586));

  xor2  gate1247(.a(G546), .b(G477), .O(gate170inter0));
  nand2 gate1248(.a(gate170inter0), .b(s_100), .O(gate170inter1));
  and2  gate1249(.a(G546), .b(G477), .O(gate170inter2));
  inv1  gate1250(.a(s_100), .O(gate170inter3));
  inv1  gate1251(.a(s_101), .O(gate170inter4));
  nand2 gate1252(.a(gate170inter4), .b(gate170inter3), .O(gate170inter5));
  nor2  gate1253(.a(gate170inter5), .b(gate170inter2), .O(gate170inter6));
  inv1  gate1254(.a(G477), .O(gate170inter7));
  inv1  gate1255(.a(G546), .O(gate170inter8));
  nand2 gate1256(.a(gate170inter8), .b(gate170inter7), .O(gate170inter9));
  nand2 gate1257(.a(s_101), .b(gate170inter3), .O(gate170inter10));
  nor2  gate1258(.a(gate170inter10), .b(gate170inter9), .O(gate170inter11));
  nor2  gate1259(.a(gate170inter11), .b(gate170inter6), .O(gate170inter12));
  nand2 gate1260(.a(gate170inter12), .b(gate170inter1), .O(G587));
nand2 gate171( .a(G480), .b(G549), .O(G588) );
nand2 gate172( .a(G483), .b(G549), .O(G589) );
nand2 gate173( .a(G486), .b(G552), .O(G590) );
nand2 gate174( .a(G489), .b(G552), .O(G591) );
nand2 gate175( .a(G492), .b(G555), .O(G592) );
nand2 gate176( .a(G495), .b(G555), .O(G593) );
nand2 gate177( .a(G498), .b(G558), .O(G594) );
nand2 gate178( .a(G501), .b(G558), .O(G595) );

  xor2  gate967(.a(G561), .b(G504), .O(gate179inter0));
  nand2 gate968(.a(gate179inter0), .b(s_60), .O(gate179inter1));
  and2  gate969(.a(G561), .b(G504), .O(gate179inter2));
  inv1  gate970(.a(s_60), .O(gate179inter3));
  inv1  gate971(.a(s_61), .O(gate179inter4));
  nand2 gate972(.a(gate179inter4), .b(gate179inter3), .O(gate179inter5));
  nor2  gate973(.a(gate179inter5), .b(gate179inter2), .O(gate179inter6));
  inv1  gate974(.a(G504), .O(gate179inter7));
  inv1  gate975(.a(G561), .O(gate179inter8));
  nand2 gate976(.a(gate179inter8), .b(gate179inter7), .O(gate179inter9));
  nand2 gate977(.a(s_61), .b(gate179inter3), .O(gate179inter10));
  nor2  gate978(.a(gate179inter10), .b(gate179inter9), .O(gate179inter11));
  nor2  gate979(.a(gate179inter11), .b(gate179inter6), .O(gate179inter12));
  nand2 gate980(.a(gate179inter12), .b(gate179inter1), .O(G596));
nand2 gate180( .a(G507), .b(G561), .O(G597) );
nand2 gate181( .a(G510), .b(G564), .O(G598) );
nand2 gate182( .a(G513), .b(G564), .O(G599) );
nand2 gate183( .a(G516), .b(G567), .O(G600) );
nand2 gate184( .a(G519), .b(G567), .O(G601) );

  xor2  gate981(.a(G571), .b(G570), .O(gate185inter0));
  nand2 gate982(.a(gate185inter0), .b(s_62), .O(gate185inter1));
  and2  gate983(.a(G571), .b(G570), .O(gate185inter2));
  inv1  gate984(.a(s_62), .O(gate185inter3));
  inv1  gate985(.a(s_63), .O(gate185inter4));
  nand2 gate986(.a(gate185inter4), .b(gate185inter3), .O(gate185inter5));
  nor2  gate987(.a(gate185inter5), .b(gate185inter2), .O(gate185inter6));
  inv1  gate988(.a(G570), .O(gate185inter7));
  inv1  gate989(.a(G571), .O(gate185inter8));
  nand2 gate990(.a(gate185inter8), .b(gate185inter7), .O(gate185inter9));
  nand2 gate991(.a(s_63), .b(gate185inter3), .O(gate185inter10));
  nor2  gate992(.a(gate185inter10), .b(gate185inter9), .O(gate185inter11));
  nor2  gate993(.a(gate185inter11), .b(gate185inter6), .O(gate185inter12));
  nand2 gate994(.a(gate185inter12), .b(gate185inter1), .O(G602));
nand2 gate186( .a(G572), .b(G573), .O(G607) );
nand2 gate187( .a(G574), .b(G575), .O(G612) );
nand2 gate188( .a(G576), .b(G577), .O(G617) );
nand2 gate189( .a(G578), .b(G579), .O(G622) );
nand2 gate190( .a(G580), .b(G581), .O(G627) );
nand2 gate191( .a(G582), .b(G583), .O(G632) );
nand2 gate192( .a(G584), .b(G585), .O(G637) );
nand2 gate193( .a(G586), .b(G587), .O(G642) );
nand2 gate194( .a(G588), .b(G589), .O(G645) );
nand2 gate195( .a(G590), .b(G591), .O(G648) );
nand2 gate196( .a(G592), .b(G593), .O(G651) );
nand2 gate197( .a(G594), .b(G595), .O(G654) );
nand2 gate198( .a(G596), .b(G597), .O(G657) );
nand2 gate199( .a(G598), .b(G599), .O(G660) );

  xor2  gate855(.a(G601), .b(G600), .O(gate200inter0));
  nand2 gate856(.a(gate200inter0), .b(s_44), .O(gate200inter1));
  and2  gate857(.a(G601), .b(G600), .O(gate200inter2));
  inv1  gate858(.a(s_44), .O(gate200inter3));
  inv1  gate859(.a(s_45), .O(gate200inter4));
  nand2 gate860(.a(gate200inter4), .b(gate200inter3), .O(gate200inter5));
  nor2  gate861(.a(gate200inter5), .b(gate200inter2), .O(gate200inter6));
  inv1  gate862(.a(G600), .O(gate200inter7));
  inv1  gate863(.a(G601), .O(gate200inter8));
  nand2 gate864(.a(gate200inter8), .b(gate200inter7), .O(gate200inter9));
  nand2 gate865(.a(s_45), .b(gate200inter3), .O(gate200inter10));
  nor2  gate866(.a(gate200inter10), .b(gate200inter9), .O(gate200inter11));
  nor2  gate867(.a(gate200inter11), .b(gate200inter6), .O(gate200inter12));
  nand2 gate868(.a(gate200inter12), .b(gate200inter1), .O(G663));

  xor2  gate1219(.a(G607), .b(G602), .O(gate201inter0));
  nand2 gate1220(.a(gate201inter0), .b(s_96), .O(gate201inter1));
  and2  gate1221(.a(G607), .b(G602), .O(gate201inter2));
  inv1  gate1222(.a(s_96), .O(gate201inter3));
  inv1  gate1223(.a(s_97), .O(gate201inter4));
  nand2 gate1224(.a(gate201inter4), .b(gate201inter3), .O(gate201inter5));
  nor2  gate1225(.a(gate201inter5), .b(gate201inter2), .O(gate201inter6));
  inv1  gate1226(.a(G602), .O(gate201inter7));
  inv1  gate1227(.a(G607), .O(gate201inter8));
  nand2 gate1228(.a(gate201inter8), .b(gate201inter7), .O(gate201inter9));
  nand2 gate1229(.a(s_97), .b(gate201inter3), .O(gate201inter10));
  nor2  gate1230(.a(gate201inter10), .b(gate201inter9), .O(gate201inter11));
  nor2  gate1231(.a(gate201inter11), .b(gate201inter6), .O(gate201inter12));
  nand2 gate1232(.a(gate201inter12), .b(gate201inter1), .O(G666));
nand2 gate202( .a(G612), .b(G617), .O(G669) );
nand2 gate203( .a(G602), .b(G612), .O(G672) );
nand2 gate204( .a(G607), .b(G617), .O(G675) );
nand2 gate205( .a(G622), .b(G627), .O(G678) );
nand2 gate206( .a(G632), .b(G637), .O(G681) );

  xor2  gate547(.a(G632), .b(G622), .O(gate207inter0));
  nand2 gate548(.a(gate207inter0), .b(s_0), .O(gate207inter1));
  and2  gate549(.a(G632), .b(G622), .O(gate207inter2));
  inv1  gate550(.a(s_0), .O(gate207inter3));
  inv1  gate551(.a(s_1), .O(gate207inter4));
  nand2 gate552(.a(gate207inter4), .b(gate207inter3), .O(gate207inter5));
  nor2  gate553(.a(gate207inter5), .b(gate207inter2), .O(gate207inter6));
  inv1  gate554(.a(G622), .O(gate207inter7));
  inv1  gate555(.a(G632), .O(gate207inter8));
  nand2 gate556(.a(gate207inter8), .b(gate207inter7), .O(gate207inter9));
  nand2 gate557(.a(s_1), .b(gate207inter3), .O(gate207inter10));
  nor2  gate558(.a(gate207inter10), .b(gate207inter9), .O(gate207inter11));
  nor2  gate559(.a(gate207inter11), .b(gate207inter6), .O(gate207inter12));
  nand2 gate560(.a(gate207inter12), .b(gate207inter1), .O(G684));
nand2 gate208( .a(G627), .b(G637), .O(G687) );
nand2 gate209( .a(G602), .b(G666), .O(G690) );

  xor2  gate659(.a(G666), .b(G607), .O(gate210inter0));
  nand2 gate660(.a(gate210inter0), .b(s_16), .O(gate210inter1));
  and2  gate661(.a(G666), .b(G607), .O(gate210inter2));
  inv1  gate662(.a(s_16), .O(gate210inter3));
  inv1  gate663(.a(s_17), .O(gate210inter4));
  nand2 gate664(.a(gate210inter4), .b(gate210inter3), .O(gate210inter5));
  nor2  gate665(.a(gate210inter5), .b(gate210inter2), .O(gate210inter6));
  inv1  gate666(.a(G607), .O(gate210inter7));
  inv1  gate667(.a(G666), .O(gate210inter8));
  nand2 gate668(.a(gate210inter8), .b(gate210inter7), .O(gate210inter9));
  nand2 gate669(.a(s_17), .b(gate210inter3), .O(gate210inter10));
  nor2  gate670(.a(gate210inter10), .b(gate210inter9), .O(gate210inter11));
  nor2  gate671(.a(gate210inter11), .b(gate210inter6), .O(gate210inter12));
  nand2 gate672(.a(gate210inter12), .b(gate210inter1), .O(G691));

  xor2  gate645(.a(G669), .b(G612), .O(gate211inter0));
  nand2 gate646(.a(gate211inter0), .b(s_14), .O(gate211inter1));
  and2  gate647(.a(G669), .b(G612), .O(gate211inter2));
  inv1  gate648(.a(s_14), .O(gate211inter3));
  inv1  gate649(.a(s_15), .O(gate211inter4));
  nand2 gate650(.a(gate211inter4), .b(gate211inter3), .O(gate211inter5));
  nor2  gate651(.a(gate211inter5), .b(gate211inter2), .O(gate211inter6));
  inv1  gate652(.a(G612), .O(gate211inter7));
  inv1  gate653(.a(G669), .O(gate211inter8));
  nand2 gate654(.a(gate211inter8), .b(gate211inter7), .O(gate211inter9));
  nand2 gate655(.a(s_15), .b(gate211inter3), .O(gate211inter10));
  nor2  gate656(.a(gate211inter10), .b(gate211inter9), .O(gate211inter11));
  nor2  gate657(.a(gate211inter11), .b(gate211inter6), .O(gate211inter12));
  nand2 gate658(.a(gate211inter12), .b(gate211inter1), .O(G692));
nand2 gate212( .a(G617), .b(G669), .O(G693) );
nand2 gate213( .a(G602), .b(G672), .O(G694) );
nand2 gate214( .a(G612), .b(G672), .O(G695) );
nand2 gate215( .a(G607), .b(G675), .O(G696) );
nand2 gate216( .a(G617), .b(G675), .O(G697) );
nand2 gate217( .a(G622), .b(G678), .O(G698) );

  xor2  gate827(.a(G678), .b(G627), .O(gate218inter0));
  nand2 gate828(.a(gate218inter0), .b(s_40), .O(gate218inter1));
  and2  gate829(.a(G678), .b(G627), .O(gate218inter2));
  inv1  gate830(.a(s_40), .O(gate218inter3));
  inv1  gate831(.a(s_41), .O(gate218inter4));
  nand2 gate832(.a(gate218inter4), .b(gate218inter3), .O(gate218inter5));
  nor2  gate833(.a(gate218inter5), .b(gate218inter2), .O(gate218inter6));
  inv1  gate834(.a(G627), .O(gate218inter7));
  inv1  gate835(.a(G678), .O(gate218inter8));
  nand2 gate836(.a(gate218inter8), .b(gate218inter7), .O(gate218inter9));
  nand2 gate837(.a(s_41), .b(gate218inter3), .O(gate218inter10));
  nor2  gate838(.a(gate218inter10), .b(gate218inter9), .O(gate218inter11));
  nor2  gate839(.a(gate218inter11), .b(gate218inter6), .O(gate218inter12));
  nand2 gate840(.a(gate218inter12), .b(gate218inter1), .O(G699));
nand2 gate219( .a(G632), .b(G681), .O(G700) );
nand2 gate220( .a(G637), .b(G681), .O(G701) );
nand2 gate221( .a(G622), .b(G684), .O(G702) );
nand2 gate222( .a(G632), .b(G684), .O(G703) );

  xor2  gate911(.a(G687), .b(G627), .O(gate223inter0));
  nand2 gate912(.a(gate223inter0), .b(s_52), .O(gate223inter1));
  and2  gate913(.a(G687), .b(G627), .O(gate223inter2));
  inv1  gate914(.a(s_52), .O(gate223inter3));
  inv1  gate915(.a(s_53), .O(gate223inter4));
  nand2 gate916(.a(gate223inter4), .b(gate223inter3), .O(gate223inter5));
  nor2  gate917(.a(gate223inter5), .b(gate223inter2), .O(gate223inter6));
  inv1  gate918(.a(G627), .O(gate223inter7));
  inv1  gate919(.a(G687), .O(gate223inter8));
  nand2 gate920(.a(gate223inter8), .b(gate223inter7), .O(gate223inter9));
  nand2 gate921(.a(s_53), .b(gate223inter3), .O(gate223inter10));
  nor2  gate922(.a(gate223inter10), .b(gate223inter9), .O(gate223inter11));
  nor2  gate923(.a(gate223inter11), .b(gate223inter6), .O(gate223inter12));
  nand2 gate924(.a(gate223inter12), .b(gate223inter1), .O(G704));
nand2 gate224( .a(G637), .b(G687), .O(G705) );
nand2 gate225( .a(G690), .b(G691), .O(G706) );
nand2 gate226( .a(G692), .b(G693), .O(G709) );
nand2 gate227( .a(G694), .b(G695), .O(G712) );
nand2 gate228( .a(G696), .b(G697), .O(G715) );
nand2 gate229( .a(G698), .b(G699), .O(G718) );
nand2 gate230( .a(G700), .b(G701), .O(G721) );
nand2 gate231( .a(G702), .b(G703), .O(G724) );
nand2 gate232( .a(G704), .b(G705), .O(G727) );

  xor2  gate1177(.a(G718), .b(G242), .O(gate233inter0));
  nand2 gate1178(.a(gate233inter0), .b(s_90), .O(gate233inter1));
  and2  gate1179(.a(G718), .b(G242), .O(gate233inter2));
  inv1  gate1180(.a(s_90), .O(gate233inter3));
  inv1  gate1181(.a(s_91), .O(gate233inter4));
  nand2 gate1182(.a(gate233inter4), .b(gate233inter3), .O(gate233inter5));
  nor2  gate1183(.a(gate233inter5), .b(gate233inter2), .O(gate233inter6));
  inv1  gate1184(.a(G242), .O(gate233inter7));
  inv1  gate1185(.a(G718), .O(gate233inter8));
  nand2 gate1186(.a(gate233inter8), .b(gate233inter7), .O(gate233inter9));
  nand2 gate1187(.a(s_91), .b(gate233inter3), .O(gate233inter10));
  nor2  gate1188(.a(gate233inter10), .b(gate233inter9), .O(gate233inter11));
  nor2  gate1189(.a(gate233inter11), .b(gate233inter6), .O(gate233inter12));
  nand2 gate1190(.a(gate233inter12), .b(gate233inter1), .O(G730));

  xor2  gate1191(.a(G721), .b(G245), .O(gate234inter0));
  nand2 gate1192(.a(gate234inter0), .b(s_92), .O(gate234inter1));
  and2  gate1193(.a(G721), .b(G245), .O(gate234inter2));
  inv1  gate1194(.a(s_92), .O(gate234inter3));
  inv1  gate1195(.a(s_93), .O(gate234inter4));
  nand2 gate1196(.a(gate234inter4), .b(gate234inter3), .O(gate234inter5));
  nor2  gate1197(.a(gate234inter5), .b(gate234inter2), .O(gate234inter6));
  inv1  gate1198(.a(G245), .O(gate234inter7));
  inv1  gate1199(.a(G721), .O(gate234inter8));
  nand2 gate1200(.a(gate234inter8), .b(gate234inter7), .O(gate234inter9));
  nand2 gate1201(.a(s_93), .b(gate234inter3), .O(gate234inter10));
  nor2  gate1202(.a(gate234inter10), .b(gate234inter9), .O(gate234inter11));
  nor2  gate1203(.a(gate234inter11), .b(gate234inter6), .O(gate234inter12));
  nand2 gate1204(.a(gate234inter12), .b(gate234inter1), .O(G733));

  xor2  gate813(.a(G724), .b(G248), .O(gate235inter0));
  nand2 gate814(.a(gate235inter0), .b(s_38), .O(gate235inter1));
  and2  gate815(.a(G724), .b(G248), .O(gate235inter2));
  inv1  gate816(.a(s_38), .O(gate235inter3));
  inv1  gate817(.a(s_39), .O(gate235inter4));
  nand2 gate818(.a(gate235inter4), .b(gate235inter3), .O(gate235inter5));
  nor2  gate819(.a(gate235inter5), .b(gate235inter2), .O(gate235inter6));
  inv1  gate820(.a(G248), .O(gate235inter7));
  inv1  gate821(.a(G724), .O(gate235inter8));
  nand2 gate822(.a(gate235inter8), .b(gate235inter7), .O(gate235inter9));
  nand2 gate823(.a(s_39), .b(gate235inter3), .O(gate235inter10));
  nor2  gate824(.a(gate235inter10), .b(gate235inter9), .O(gate235inter11));
  nor2  gate825(.a(gate235inter11), .b(gate235inter6), .O(gate235inter12));
  nand2 gate826(.a(gate235inter12), .b(gate235inter1), .O(G736));
nand2 gate236( .a(G251), .b(G727), .O(G739) );
nand2 gate237( .a(G254), .b(G706), .O(G742) );
nand2 gate238( .a(G257), .b(G709), .O(G745) );
nand2 gate239( .a(G260), .b(G712), .O(G748) );
nand2 gate240( .a(G263), .b(G715), .O(G751) );
nand2 gate241( .a(G242), .b(G730), .O(G754) );
nand2 gate242( .a(G718), .b(G730), .O(G755) );
nand2 gate243( .a(G245), .b(G733), .O(G756) );

  xor2  gate771(.a(G733), .b(G721), .O(gate244inter0));
  nand2 gate772(.a(gate244inter0), .b(s_32), .O(gate244inter1));
  and2  gate773(.a(G733), .b(G721), .O(gate244inter2));
  inv1  gate774(.a(s_32), .O(gate244inter3));
  inv1  gate775(.a(s_33), .O(gate244inter4));
  nand2 gate776(.a(gate244inter4), .b(gate244inter3), .O(gate244inter5));
  nor2  gate777(.a(gate244inter5), .b(gate244inter2), .O(gate244inter6));
  inv1  gate778(.a(G721), .O(gate244inter7));
  inv1  gate779(.a(G733), .O(gate244inter8));
  nand2 gate780(.a(gate244inter8), .b(gate244inter7), .O(gate244inter9));
  nand2 gate781(.a(s_33), .b(gate244inter3), .O(gate244inter10));
  nor2  gate782(.a(gate244inter10), .b(gate244inter9), .O(gate244inter11));
  nor2  gate783(.a(gate244inter11), .b(gate244inter6), .O(gate244inter12));
  nand2 gate784(.a(gate244inter12), .b(gate244inter1), .O(G757));
nand2 gate245( .a(G248), .b(G736), .O(G758) );
nand2 gate246( .a(G724), .b(G736), .O(G759) );
nand2 gate247( .a(G251), .b(G739), .O(G760) );
nand2 gate248( .a(G727), .b(G739), .O(G761) );
nand2 gate249( .a(G254), .b(G742), .O(G762) );
nand2 gate250( .a(G706), .b(G742), .O(G763) );
nand2 gate251( .a(G257), .b(G745), .O(G764) );
nand2 gate252( .a(G709), .b(G745), .O(G765) );
nand2 gate253( .a(G260), .b(G748), .O(G766) );

  xor2  gate799(.a(G748), .b(G712), .O(gate254inter0));
  nand2 gate800(.a(gate254inter0), .b(s_36), .O(gate254inter1));
  and2  gate801(.a(G748), .b(G712), .O(gate254inter2));
  inv1  gate802(.a(s_36), .O(gate254inter3));
  inv1  gate803(.a(s_37), .O(gate254inter4));
  nand2 gate804(.a(gate254inter4), .b(gate254inter3), .O(gate254inter5));
  nor2  gate805(.a(gate254inter5), .b(gate254inter2), .O(gate254inter6));
  inv1  gate806(.a(G712), .O(gate254inter7));
  inv1  gate807(.a(G748), .O(gate254inter8));
  nand2 gate808(.a(gate254inter8), .b(gate254inter7), .O(gate254inter9));
  nand2 gate809(.a(s_37), .b(gate254inter3), .O(gate254inter10));
  nor2  gate810(.a(gate254inter10), .b(gate254inter9), .O(gate254inter11));
  nor2  gate811(.a(gate254inter11), .b(gate254inter6), .O(gate254inter12));
  nand2 gate812(.a(gate254inter12), .b(gate254inter1), .O(G767));
nand2 gate255( .a(G263), .b(G751), .O(G768) );

  xor2  gate603(.a(G751), .b(G715), .O(gate256inter0));
  nand2 gate604(.a(gate256inter0), .b(s_8), .O(gate256inter1));
  and2  gate605(.a(G751), .b(G715), .O(gate256inter2));
  inv1  gate606(.a(s_8), .O(gate256inter3));
  inv1  gate607(.a(s_9), .O(gate256inter4));
  nand2 gate608(.a(gate256inter4), .b(gate256inter3), .O(gate256inter5));
  nor2  gate609(.a(gate256inter5), .b(gate256inter2), .O(gate256inter6));
  inv1  gate610(.a(G715), .O(gate256inter7));
  inv1  gate611(.a(G751), .O(gate256inter8));
  nand2 gate612(.a(gate256inter8), .b(gate256inter7), .O(gate256inter9));
  nand2 gate613(.a(s_9), .b(gate256inter3), .O(gate256inter10));
  nor2  gate614(.a(gate256inter10), .b(gate256inter9), .O(gate256inter11));
  nor2  gate615(.a(gate256inter11), .b(gate256inter6), .O(gate256inter12));
  nand2 gate616(.a(gate256inter12), .b(gate256inter1), .O(G769));
nand2 gate257( .a(G754), .b(G755), .O(G770) );
nand2 gate258( .a(G756), .b(G757), .O(G773) );
nand2 gate259( .a(G758), .b(G759), .O(G776) );
nand2 gate260( .a(G760), .b(G761), .O(G779) );
nand2 gate261( .a(G762), .b(G763), .O(G782) );
nand2 gate262( .a(G764), .b(G765), .O(G785) );
nand2 gate263( .a(G766), .b(G767), .O(G788) );
nand2 gate264( .a(G768), .b(G769), .O(G791) );
nand2 gate265( .a(G642), .b(G770), .O(G794) );
nand2 gate266( .a(G645), .b(G773), .O(G797) );
nand2 gate267( .a(G648), .b(G776), .O(G800) );
nand2 gate268( .a(G651), .b(G779), .O(G803) );
nand2 gate269( .a(G654), .b(G782), .O(G806) );
nand2 gate270( .a(G657), .b(G785), .O(G809) );
nand2 gate271( .a(G660), .b(G788), .O(G812) );
nand2 gate272( .a(G663), .b(G791), .O(G815) );
nand2 gate273( .a(G642), .b(G794), .O(G818) );

  xor2  gate1275(.a(G794), .b(G770), .O(gate274inter0));
  nand2 gate1276(.a(gate274inter0), .b(s_104), .O(gate274inter1));
  and2  gate1277(.a(G794), .b(G770), .O(gate274inter2));
  inv1  gate1278(.a(s_104), .O(gate274inter3));
  inv1  gate1279(.a(s_105), .O(gate274inter4));
  nand2 gate1280(.a(gate274inter4), .b(gate274inter3), .O(gate274inter5));
  nor2  gate1281(.a(gate274inter5), .b(gate274inter2), .O(gate274inter6));
  inv1  gate1282(.a(G770), .O(gate274inter7));
  inv1  gate1283(.a(G794), .O(gate274inter8));
  nand2 gate1284(.a(gate274inter8), .b(gate274inter7), .O(gate274inter9));
  nand2 gate1285(.a(s_105), .b(gate274inter3), .O(gate274inter10));
  nor2  gate1286(.a(gate274inter10), .b(gate274inter9), .O(gate274inter11));
  nor2  gate1287(.a(gate274inter11), .b(gate274inter6), .O(gate274inter12));
  nand2 gate1288(.a(gate274inter12), .b(gate274inter1), .O(G819));
nand2 gate275( .a(G645), .b(G797), .O(G820) );

  xor2  gate995(.a(G797), .b(G773), .O(gate276inter0));
  nand2 gate996(.a(gate276inter0), .b(s_64), .O(gate276inter1));
  and2  gate997(.a(G797), .b(G773), .O(gate276inter2));
  inv1  gate998(.a(s_64), .O(gate276inter3));
  inv1  gate999(.a(s_65), .O(gate276inter4));
  nand2 gate1000(.a(gate276inter4), .b(gate276inter3), .O(gate276inter5));
  nor2  gate1001(.a(gate276inter5), .b(gate276inter2), .O(gate276inter6));
  inv1  gate1002(.a(G773), .O(gate276inter7));
  inv1  gate1003(.a(G797), .O(gate276inter8));
  nand2 gate1004(.a(gate276inter8), .b(gate276inter7), .O(gate276inter9));
  nand2 gate1005(.a(s_65), .b(gate276inter3), .O(gate276inter10));
  nor2  gate1006(.a(gate276inter10), .b(gate276inter9), .O(gate276inter11));
  nor2  gate1007(.a(gate276inter11), .b(gate276inter6), .O(gate276inter12));
  nand2 gate1008(.a(gate276inter12), .b(gate276inter1), .O(G821));
nand2 gate277( .a(G648), .b(G800), .O(G822) );
nand2 gate278( .a(G776), .b(G800), .O(G823) );
nand2 gate279( .a(G651), .b(G803), .O(G824) );
nand2 gate280( .a(G779), .b(G803), .O(G825) );
nand2 gate281( .a(G654), .b(G806), .O(G826) );

  xor2  gate1009(.a(G806), .b(G782), .O(gate282inter0));
  nand2 gate1010(.a(gate282inter0), .b(s_66), .O(gate282inter1));
  and2  gate1011(.a(G806), .b(G782), .O(gate282inter2));
  inv1  gate1012(.a(s_66), .O(gate282inter3));
  inv1  gate1013(.a(s_67), .O(gate282inter4));
  nand2 gate1014(.a(gate282inter4), .b(gate282inter3), .O(gate282inter5));
  nor2  gate1015(.a(gate282inter5), .b(gate282inter2), .O(gate282inter6));
  inv1  gate1016(.a(G782), .O(gate282inter7));
  inv1  gate1017(.a(G806), .O(gate282inter8));
  nand2 gate1018(.a(gate282inter8), .b(gate282inter7), .O(gate282inter9));
  nand2 gate1019(.a(s_67), .b(gate282inter3), .O(gate282inter10));
  nor2  gate1020(.a(gate282inter10), .b(gate282inter9), .O(gate282inter11));
  nor2  gate1021(.a(gate282inter11), .b(gate282inter6), .O(gate282inter12));
  nand2 gate1022(.a(gate282inter12), .b(gate282inter1), .O(G827));
nand2 gate283( .a(G657), .b(G809), .O(G828) );
nand2 gate284( .a(G785), .b(G809), .O(G829) );
nand2 gate285( .a(G660), .b(G812), .O(G830) );
nand2 gate286( .a(G788), .b(G812), .O(G831) );
nand2 gate287( .a(G663), .b(G815), .O(G832) );
nand2 gate288( .a(G791), .b(G815), .O(G833) );
nand2 gate289( .a(G818), .b(G819), .O(G834) );
nand2 gate290( .a(G820), .b(G821), .O(G847) );
nand2 gate291( .a(G822), .b(G823), .O(G860) );
nand2 gate292( .a(G824), .b(G825), .O(G873) );
nand2 gate293( .a(G828), .b(G829), .O(G886) );
nand2 gate294( .a(G832), .b(G833), .O(G899) );
nand2 gate295( .a(G830), .b(G831), .O(G912) );
nand2 gate296( .a(G826), .b(G827), .O(G925) );
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );
nand2 gate387( .a(G1), .b(G1036), .O(G1132) );
nand2 gate388( .a(G2), .b(G1039), .O(G1135) );
nand2 gate389( .a(G3), .b(G1042), .O(G1138) );

  xor2  gate673(.a(G1045), .b(G4), .O(gate390inter0));
  nand2 gate674(.a(gate390inter0), .b(s_18), .O(gate390inter1));
  and2  gate675(.a(G1045), .b(G4), .O(gate390inter2));
  inv1  gate676(.a(s_18), .O(gate390inter3));
  inv1  gate677(.a(s_19), .O(gate390inter4));
  nand2 gate678(.a(gate390inter4), .b(gate390inter3), .O(gate390inter5));
  nor2  gate679(.a(gate390inter5), .b(gate390inter2), .O(gate390inter6));
  inv1  gate680(.a(G4), .O(gate390inter7));
  inv1  gate681(.a(G1045), .O(gate390inter8));
  nand2 gate682(.a(gate390inter8), .b(gate390inter7), .O(gate390inter9));
  nand2 gate683(.a(s_19), .b(gate390inter3), .O(gate390inter10));
  nor2  gate684(.a(gate390inter10), .b(gate390inter9), .O(gate390inter11));
  nor2  gate685(.a(gate390inter11), .b(gate390inter6), .O(gate390inter12));
  nand2 gate686(.a(gate390inter12), .b(gate390inter1), .O(G1141));
nand2 gate391( .a(G5), .b(G1048), .O(G1144) );
nand2 gate392( .a(G6), .b(G1051), .O(G1147) );
nand2 gate393( .a(G7), .b(G1054), .O(G1150) );
nand2 gate394( .a(G8), .b(G1057), .O(G1153) );
nand2 gate395( .a(G9), .b(G1060), .O(G1156) );

  xor2  gate1163(.a(G1063), .b(G10), .O(gate396inter0));
  nand2 gate1164(.a(gate396inter0), .b(s_88), .O(gate396inter1));
  and2  gate1165(.a(G1063), .b(G10), .O(gate396inter2));
  inv1  gate1166(.a(s_88), .O(gate396inter3));
  inv1  gate1167(.a(s_89), .O(gate396inter4));
  nand2 gate1168(.a(gate396inter4), .b(gate396inter3), .O(gate396inter5));
  nor2  gate1169(.a(gate396inter5), .b(gate396inter2), .O(gate396inter6));
  inv1  gate1170(.a(G10), .O(gate396inter7));
  inv1  gate1171(.a(G1063), .O(gate396inter8));
  nand2 gate1172(.a(gate396inter8), .b(gate396inter7), .O(gate396inter9));
  nand2 gate1173(.a(s_89), .b(gate396inter3), .O(gate396inter10));
  nor2  gate1174(.a(gate396inter10), .b(gate396inter9), .O(gate396inter11));
  nor2  gate1175(.a(gate396inter11), .b(gate396inter6), .O(gate396inter12));
  nand2 gate1176(.a(gate396inter12), .b(gate396inter1), .O(G1159));
nand2 gate397( .a(G11), .b(G1066), .O(G1162) );
nand2 gate398( .a(G12), .b(G1069), .O(G1165) );
nand2 gate399( .a(G13), .b(G1072), .O(G1168) );
nand2 gate400( .a(G14), .b(G1075), .O(G1171) );
nand2 gate401( .a(G15), .b(G1078), .O(G1174) );
nand2 gate402( .a(G16), .b(G1081), .O(G1177) );
nand2 gate403( .a(G17), .b(G1084), .O(G1180) );
nand2 gate404( .a(G18), .b(G1087), .O(G1183) );

  xor2  gate1205(.a(G1090), .b(G19), .O(gate405inter0));
  nand2 gate1206(.a(gate405inter0), .b(s_94), .O(gate405inter1));
  and2  gate1207(.a(G1090), .b(G19), .O(gate405inter2));
  inv1  gate1208(.a(s_94), .O(gate405inter3));
  inv1  gate1209(.a(s_95), .O(gate405inter4));
  nand2 gate1210(.a(gate405inter4), .b(gate405inter3), .O(gate405inter5));
  nor2  gate1211(.a(gate405inter5), .b(gate405inter2), .O(gate405inter6));
  inv1  gate1212(.a(G19), .O(gate405inter7));
  inv1  gate1213(.a(G1090), .O(gate405inter8));
  nand2 gate1214(.a(gate405inter8), .b(gate405inter7), .O(gate405inter9));
  nand2 gate1215(.a(s_95), .b(gate405inter3), .O(gate405inter10));
  nor2  gate1216(.a(gate405inter10), .b(gate405inter9), .O(gate405inter11));
  nor2  gate1217(.a(gate405inter11), .b(gate405inter6), .O(gate405inter12));
  nand2 gate1218(.a(gate405inter12), .b(gate405inter1), .O(G1186));

  xor2  gate939(.a(G1093), .b(G20), .O(gate406inter0));
  nand2 gate940(.a(gate406inter0), .b(s_56), .O(gate406inter1));
  and2  gate941(.a(G1093), .b(G20), .O(gate406inter2));
  inv1  gate942(.a(s_56), .O(gate406inter3));
  inv1  gate943(.a(s_57), .O(gate406inter4));
  nand2 gate944(.a(gate406inter4), .b(gate406inter3), .O(gate406inter5));
  nor2  gate945(.a(gate406inter5), .b(gate406inter2), .O(gate406inter6));
  inv1  gate946(.a(G20), .O(gate406inter7));
  inv1  gate947(.a(G1093), .O(gate406inter8));
  nand2 gate948(.a(gate406inter8), .b(gate406inter7), .O(gate406inter9));
  nand2 gate949(.a(s_57), .b(gate406inter3), .O(gate406inter10));
  nor2  gate950(.a(gate406inter10), .b(gate406inter9), .O(gate406inter11));
  nor2  gate951(.a(gate406inter11), .b(gate406inter6), .O(gate406inter12));
  nand2 gate952(.a(gate406inter12), .b(gate406inter1), .O(G1189));
nand2 gate407( .a(G21), .b(G1096), .O(G1192) );
nand2 gate408( .a(G22), .b(G1099), .O(G1195) );
nand2 gate409( .a(G23), .b(G1102), .O(G1198) );
nand2 gate410( .a(G24), .b(G1105), .O(G1201) );
nand2 gate411( .a(G25), .b(G1108), .O(G1204) );

  xor2  gate757(.a(G1111), .b(G26), .O(gate412inter0));
  nand2 gate758(.a(gate412inter0), .b(s_30), .O(gate412inter1));
  and2  gate759(.a(G1111), .b(G26), .O(gate412inter2));
  inv1  gate760(.a(s_30), .O(gate412inter3));
  inv1  gate761(.a(s_31), .O(gate412inter4));
  nand2 gate762(.a(gate412inter4), .b(gate412inter3), .O(gate412inter5));
  nor2  gate763(.a(gate412inter5), .b(gate412inter2), .O(gate412inter6));
  inv1  gate764(.a(G26), .O(gate412inter7));
  inv1  gate765(.a(G1111), .O(gate412inter8));
  nand2 gate766(.a(gate412inter8), .b(gate412inter7), .O(gate412inter9));
  nand2 gate767(.a(s_31), .b(gate412inter3), .O(gate412inter10));
  nor2  gate768(.a(gate412inter10), .b(gate412inter9), .O(gate412inter11));
  nor2  gate769(.a(gate412inter11), .b(gate412inter6), .O(gate412inter12));
  nand2 gate770(.a(gate412inter12), .b(gate412inter1), .O(G1207));
nand2 gate413( .a(G27), .b(G1114), .O(G1210) );
nand2 gate414( .a(G28), .b(G1117), .O(G1213) );

  xor2  gate1135(.a(G1120), .b(G29), .O(gate415inter0));
  nand2 gate1136(.a(gate415inter0), .b(s_84), .O(gate415inter1));
  and2  gate1137(.a(G1120), .b(G29), .O(gate415inter2));
  inv1  gate1138(.a(s_84), .O(gate415inter3));
  inv1  gate1139(.a(s_85), .O(gate415inter4));
  nand2 gate1140(.a(gate415inter4), .b(gate415inter3), .O(gate415inter5));
  nor2  gate1141(.a(gate415inter5), .b(gate415inter2), .O(gate415inter6));
  inv1  gate1142(.a(G29), .O(gate415inter7));
  inv1  gate1143(.a(G1120), .O(gate415inter8));
  nand2 gate1144(.a(gate415inter8), .b(gate415inter7), .O(gate415inter9));
  nand2 gate1145(.a(s_85), .b(gate415inter3), .O(gate415inter10));
  nor2  gate1146(.a(gate415inter10), .b(gate415inter9), .O(gate415inter11));
  nor2  gate1147(.a(gate415inter11), .b(gate415inter6), .O(gate415inter12));
  nand2 gate1148(.a(gate415inter12), .b(gate415inter1), .O(G1216));
nand2 gate416( .a(G30), .b(G1123), .O(G1219) );
nand2 gate417( .a(G31), .b(G1126), .O(G1222) );
nand2 gate418( .a(G32), .b(G1129), .O(G1225) );
nand2 gate419( .a(G1), .b(G1132), .O(G1228) );
nand2 gate420( .a(G1036), .b(G1132), .O(G1229) );
nand2 gate421( .a(G2), .b(G1135), .O(G1230) );

  xor2  gate575(.a(G1135), .b(G1039), .O(gate422inter0));
  nand2 gate576(.a(gate422inter0), .b(s_4), .O(gate422inter1));
  and2  gate577(.a(G1135), .b(G1039), .O(gate422inter2));
  inv1  gate578(.a(s_4), .O(gate422inter3));
  inv1  gate579(.a(s_5), .O(gate422inter4));
  nand2 gate580(.a(gate422inter4), .b(gate422inter3), .O(gate422inter5));
  nor2  gate581(.a(gate422inter5), .b(gate422inter2), .O(gate422inter6));
  inv1  gate582(.a(G1039), .O(gate422inter7));
  inv1  gate583(.a(G1135), .O(gate422inter8));
  nand2 gate584(.a(gate422inter8), .b(gate422inter7), .O(gate422inter9));
  nand2 gate585(.a(s_5), .b(gate422inter3), .O(gate422inter10));
  nor2  gate586(.a(gate422inter10), .b(gate422inter9), .O(gate422inter11));
  nor2  gate587(.a(gate422inter11), .b(gate422inter6), .O(gate422inter12));
  nand2 gate588(.a(gate422inter12), .b(gate422inter1), .O(G1231));
nand2 gate423( .a(G3), .b(G1138), .O(G1232) );
nand2 gate424( .a(G1042), .b(G1138), .O(G1233) );
nand2 gate425( .a(G4), .b(G1141), .O(G1234) );
nand2 gate426( .a(G1045), .b(G1141), .O(G1235) );
nand2 gate427( .a(G5), .b(G1144), .O(G1236) );

  xor2  gate589(.a(G1144), .b(G1048), .O(gate428inter0));
  nand2 gate590(.a(gate428inter0), .b(s_6), .O(gate428inter1));
  and2  gate591(.a(G1144), .b(G1048), .O(gate428inter2));
  inv1  gate592(.a(s_6), .O(gate428inter3));
  inv1  gate593(.a(s_7), .O(gate428inter4));
  nand2 gate594(.a(gate428inter4), .b(gate428inter3), .O(gate428inter5));
  nor2  gate595(.a(gate428inter5), .b(gate428inter2), .O(gate428inter6));
  inv1  gate596(.a(G1048), .O(gate428inter7));
  inv1  gate597(.a(G1144), .O(gate428inter8));
  nand2 gate598(.a(gate428inter8), .b(gate428inter7), .O(gate428inter9));
  nand2 gate599(.a(s_7), .b(gate428inter3), .O(gate428inter10));
  nor2  gate600(.a(gate428inter10), .b(gate428inter9), .O(gate428inter11));
  nor2  gate601(.a(gate428inter11), .b(gate428inter6), .O(gate428inter12));
  nand2 gate602(.a(gate428inter12), .b(gate428inter1), .O(G1237));
nand2 gate429( .a(G6), .b(G1147), .O(G1238) );
nand2 gate430( .a(G1051), .b(G1147), .O(G1239) );
nand2 gate431( .a(G7), .b(G1150), .O(G1240) );

  xor2  gate715(.a(G1150), .b(G1054), .O(gate432inter0));
  nand2 gate716(.a(gate432inter0), .b(s_24), .O(gate432inter1));
  and2  gate717(.a(G1150), .b(G1054), .O(gate432inter2));
  inv1  gate718(.a(s_24), .O(gate432inter3));
  inv1  gate719(.a(s_25), .O(gate432inter4));
  nand2 gate720(.a(gate432inter4), .b(gate432inter3), .O(gate432inter5));
  nor2  gate721(.a(gate432inter5), .b(gate432inter2), .O(gate432inter6));
  inv1  gate722(.a(G1054), .O(gate432inter7));
  inv1  gate723(.a(G1150), .O(gate432inter8));
  nand2 gate724(.a(gate432inter8), .b(gate432inter7), .O(gate432inter9));
  nand2 gate725(.a(s_25), .b(gate432inter3), .O(gate432inter10));
  nor2  gate726(.a(gate432inter10), .b(gate432inter9), .O(gate432inter11));
  nor2  gate727(.a(gate432inter11), .b(gate432inter6), .O(gate432inter12));
  nand2 gate728(.a(gate432inter12), .b(gate432inter1), .O(G1241));
nand2 gate433( .a(G8), .b(G1153), .O(G1242) );
nand2 gate434( .a(G1057), .b(G1153), .O(G1243) );
nand2 gate435( .a(G9), .b(G1156), .O(G1244) );
nand2 gate436( .a(G1060), .b(G1156), .O(G1245) );
nand2 gate437( .a(G10), .b(G1159), .O(G1246) );
nand2 gate438( .a(G1063), .b(G1159), .O(G1247) );
nand2 gate439( .a(G11), .b(G1162), .O(G1248) );
nand2 gate440( .a(G1066), .b(G1162), .O(G1249) );
nand2 gate441( .a(G12), .b(G1165), .O(G1250) );
nand2 gate442( .a(G1069), .b(G1165), .O(G1251) );
nand2 gate443( .a(G13), .b(G1168), .O(G1252) );
nand2 gate444( .a(G1072), .b(G1168), .O(G1253) );
nand2 gate445( .a(G14), .b(G1171), .O(G1254) );
nand2 gate446( .a(G1075), .b(G1171), .O(G1255) );
nand2 gate447( .a(G15), .b(G1174), .O(G1256) );
nand2 gate448( .a(G1078), .b(G1174), .O(G1257) );

  xor2  gate729(.a(G1177), .b(G16), .O(gate449inter0));
  nand2 gate730(.a(gate449inter0), .b(s_26), .O(gate449inter1));
  and2  gate731(.a(G1177), .b(G16), .O(gate449inter2));
  inv1  gate732(.a(s_26), .O(gate449inter3));
  inv1  gate733(.a(s_27), .O(gate449inter4));
  nand2 gate734(.a(gate449inter4), .b(gate449inter3), .O(gate449inter5));
  nor2  gate735(.a(gate449inter5), .b(gate449inter2), .O(gate449inter6));
  inv1  gate736(.a(G16), .O(gate449inter7));
  inv1  gate737(.a(G1177), .O(gate449inter8));
  nand2 gate738(.a(gate449inter8), .b(gate449inter7), .O(gate449inter9));
  nand2 gate739(.a(s_27), .b(gate449inter3), .O(gate449inter10));
  nor2  gate740(.a(gate449inter10), .b(gate449inter9), .O(gate449inter11));
  nor2  gate741(.a(gate449inter11), .b(gate449inter6), .O(gate449inter12));
  nand2 gate742(.a(gate449inter12), .b(gate449inter1), .O(G1258));
nand2 gate450( .a(G1081), .b(G1177), .O(G1259) );
nand2 gate451( .a(G17), .b(G1180), .O(G1260) );
nand2 gate452( .a(G1084), .b(G1180), .O(G1261) );
nand2 gate453( .a(G18), .b(G1183), .O(G1262) );
nand2 gate454( .a(G1087), .b(G1183), .O(G1263) );
nand2 gate455( .a(G19), .b(G1186), .O(G1264) );
nand2 gate456( .a(G1090), .b(G1186), .O(G1265) );
nand2 gate457( .a(G20), .b(G1189), .O(G1266) );
nand2 gate458( .a(G1093), .b(G1189), .O(G1267) );
nand2 gate459( .a(G21), .b(G1192), .O(G1268) );
nand2 gate460( .a(G1096), .b(G1192), .O(G1269) );

  xor2  gate1121(.a(G1195), .b(G22), .O(gate461inter0));
  nand2 gate1122(.a(gate461inter0), .b(s_82), .O(gate461inter1));
  and2  gate1123(.a(G1195), .b(G22), .O(gate461inter2));
  inv1  gate1124(.a(s_82), .O(gate461inter3));
  inv1  gate1125(.a(s_83), .O(gate461inter4));
  nand2 gate1126(.a(gate461inter4), .b(gate461inter3), .O(gate461inter5));
  nor2  gate1127(.a(gate461inter5), .b(gate461inter2), .O(gate461inter6));
  inv1  gate1128(.a(G22), .O(gate461inter7));
  inv1  gate1129(.a(G1195), .O(gate461inter8));
  nand2 gate1130(.a(gate461inter8), .b(gate461inter7), .O(gate461inter9));
  nand2 gate1131(.a(s_83), .b(gate461inter3), .O(gate461inter10));
  nor2  gate1132(.a(gate461inter10), .b(gate461inter9), .O(gate461inter11));
  nor2  gate1133(.a(gate461inter11), .b(gate461inter6), .O(gate461inter12));
  nand2 gate1134(.a(gate461inter12), .b(gate461inter1), .O(G1270));
nand2 gate462( .a(G1099), .b(G1195), .O(G1271) );
nand2 gate463( .a(G23), .b(G1198), .O(G1272) );
nand2 gate464( .a(G1102), .b(G1198), .O(G1273) );
nand2 gate465( .a(G24), .b(G1201), .O(G1274) );
nand2 gate466( .a(G1105), .b(G1201), .O(G1275) );
nand2 gate467( .a(G25), .b(G1204), .O(G1276) );
nand2 gate468( .a(G1108), .b(G1204), .O(G1277) );
nand2 gate469( .a(G26), .b(G1207), .O(G1278) );
nand2 gate470( .a(G1111), .b(G1207), .O(G1279) );

  xor2  gate1065(.a(G1210), .b(G27), .O(gate471inter0));
  nand2 gate1066(.a(gate471inter0), .b(s_74), .O(gate471inter1));
  and2  gate1067(.a(G1210), .b(G27), .O(gate471inter2));
  inv1  gate1068(.a(s_74), .O(gate471inter3));
  inv1  gate1069(.a(s_75), .O(gate471inter4));
  nand2 gate1070(.a(gate471inter4), .b(gate471inter3), .O(gate471inter5));
  nor2  gate1071(.a(gate471inter5), .b(gate471inter2), .O(gate471inter6));
  inv1  gate1072(.a(G27), .O(gate471inter7));
  inv1  gate1073(.a(G1210), .O(gate471inter8));
  nand2 gate1074(.a(gate471inter8), .b(gate471inter7), .O(gate471inter9));
  nand2 gate1075(.a(s_75), .b(gate471inter3), .O(gate471inter10));
  nor2  gate1076(.a(gate471inter10), .b(gate471inter9), .O(gate471inter11));
  nor2  gate1077(.a(gate471inter11), .b(gate471inter6), .O(gate471inter12));
  nand2 gate1078(.a(gate471inter12), .b(gate471inter1), .O(G1280));
nand2 gate472( .a(G1114), .b(G1210), .O(G1281) );
nand2 gate473( .a(G28), .b(G1213), .O(G1282) );
nand2 gate474( .a(G1117), .b(G1213), .O(G1283) );
nand2 gate475( .a(G29), .b(G1216), .O(G1284) );
nand2 gate476( .a(G1120), .b(G1216), .O(G1285) );

  xor2  gate631(.a(G1219), .b(G30), .O(gate477inter0));
  nand2 gate632(.a(gate477inter0), .b(s_12), .O(gate477inter1));
  and2  gate633(.a(G1219), .b(G30), .O(gate477inter2));
  inv1  gate634(.a(s_12), .O(gate477inter3));
  inv1  gate635(.a(s_13), .O(gate477inter4));
  nand2 gate636(.a(gate477inter4), .b(gate477inter3), .O(gate477inter5));
  nor2  gate637(.a(gate477inter5), .b(gate477inter2), .O(gate477inter6));
  inv1  gate638(.a(G30), .O(gate477inter7));
  inv1  gate639(.a(G1219), .O(gate477inter8));
  nand2 gate640(.a(gate477inter8), .b(gate477inter7), .O(gate477inter9));
  nand2 gate641(.a(s_13), .b(gate477inter3), .O(gate477inter10));
  nor2  gate642(.a(gate477inter10), .b(gate477inter9), .O(gate477inter11));
  nor2  gate643(.a(gate477inter11), .b(gate477inter6), .O(gate477inter12));
  nand2 gate644(.a(gate477inter12), .b(gate477inter1), .O(G1286));
nand2 gate478( .a(G1123), .b(G1219), .O(G1287) );
nand2 gate479( .a(G31), .b(G1222), .O(G1288) );
nand2 gate480( .a(G1126), .b(G1222), .O(G1289) );
nand2 gate481( .a(G32), .b(G1225), .O(G1290) );
nand2 gate482( .a(G1129), .b(G1225), .O(G1291) );
nand2 gate483( .a(G1228), .b(G1229), .O(G1292) );
nand2 gate484( .a(G1230), .b(G1231), .O(G1293) );
nand2 gate485( .a(G1232), .b(G1233), .O(G1294) );
nand2 gate486( .a(G1234), .b(G1235), .O(G1295) );
nand2 gate487( .a(G1236), .b(G1237), .O(G1296) );
nand2 gate488( .a(G1238), .b(G1239), .O(G1297) );
nand2 gate489( .a(G1240), .b(G1241), .O(G1298) );
nand2 gate490( .a(G1242), .b(G1243), .O(G1299) );
nand2 gate491( .a(G1244), .b(G1245), .O(G1300) );
nand2 gate492( .a(G1246), .b(G1247), .O(G1301) );
nand2 gate493( .a(G1248), .b(G1249), .O(G1302) );
nand2 gate494( .a(G1250), .b(G1251), .O(G1303) );

  xor2  gate1317(.a(G1253), .b(G1252), .O(gate495inter0));
  nand2 gate1318(.a(gate495inter0), .b(s_110), .O(gate495inter1));
  and2  gate1319(.a(G1253), .b(G1252), .O(gate495inter2));
  inv1  gate1320(.a(s_110), .O(gate495inter3));
  inv1  gate1321(.a(s_111), .O(gate495inter4));
  nand2 gate1322(.a(gate495inter4), .b(gate495inter3), .O(gate495inter5));
  nor2  gate1323(.a(gate495inter5), .b(gate495inter2), .O(gate495inter6));
  inv1  gate1324(.a(G1252), .O(gate495inter7));
  inv1  gate1325(.a(G1253), .O(gate495inter8));
  nand2 gate1326(.a(gate495inter8), .b(gate495inter7), .O(gate495inter9));
  nand2 gate1327(.a(s_111), .b(gate495inter3), .O(gate495inter10));
  nor2  gate1328(.a(gate495inter10), .b(gate495inter9), .O(gate495inter11));
  nor2  gate1329(.a(gate495inter11), .b(gate495inter6), .O(gate495inter12));
  nand2 gate1330(.a(gate495inter12), .b(gate495inter1), .O(G1304));
nand2 gate496( .a(G1254), .b(G1255), .O(G1305) );
nand2 gate497( .a(G1256), .b(G1257), .O(G1306) );

  xor2  gate1261(.a(G1259), .b(G1258), .O(gate498inter0));
  nand2 gate1262(.a(gate498inter0), .b(s_102), .O(gate498inter1));
  and2  gate1263(.a(G1259), .b(G1258), .O(gate498inter2));
  inv1  gate1264(.a(s_102), .O(gate498inter3));
  inv1  gate1265(.a(s_103), .O(gate498inter4));
  nand2 gate1266(.a(gate498inter4), .b(gate498inter3), .O(gate498inter5));
  nor2  gate1267(.a(gate498inter5), .b(gate498inter2), .O(gate498inter6));
  inv1  gate1268(.a(G1258), .O(gate498inter7));
  inv1  gate1269(.a(G1259), .O(gate498inter8));
  nand2 gate1270(.a(gate498inter8), .b(gate498inter7), .O(gate498inter9));
  nand2 gate1271(.a(s_103), .b(gate498inter3), .O(gate498inter10));
  nor2  gate1272(.a(gate498inter10), .b(gate498inter9), .O(gate498inter11));
  nor2  gate1273(.a(gate498inter11), .b(gate498inter6), .O(gate498inter12));
  nand2 gate1274(.a(gate498inter12), .b(gate498inter1), .O(G1307));

  xor2  gate1023(.a(G1261), .b(G1260), .O(gate499inter0));
  nand2 gate1024(.a(gate499inter0), .b(s_68), .O(gate499inter1));
  and2  gate1025(.a(G1261), .b(G1260), .O(gate499inter2));
  inv1  gate1026(.a(s_68), .O(gate499inter3));
  inv1  gate1027(.a(s_69), .O(gate499inter4));
  nand2 gate1028(.a(gate499inter4), .b(gate499inter3), .O(gate499inter5));
  nor2  gate1029(.a(gate499inter5), .b(gate499inter2), .O(gate499inter6));
  inv1  gate1030(.a(G1260), .O(gate499inter7));
  inv1  gate1031(.a(G1261), .O(gate499inter8));
  nand2 gate1032(.a(gate499inter8), .b(gate499inter7), .O(gate499inter9));
  nand2 gate1033(.a(s_69), .b(gate499inter3), .O(gate499inter10));
  nor2  gate1034(.a(gate499inter10), .b(gate499inter9), .O(gate499inter11));
  nor2  gate1035(.a(gate499inter11), .b(gate499inter6), .O(gate499inter12));
  nand2 gate1036(.a(gate499inter12), .b(gate499inter1), .O(G1308));
nand2 gate500( .a(G1262), .b(G1263), .O(G1309) );
nand2 gate501( .a(G1264), .b(G1265), .O(G1310) );
nand2 gate502( .a(G1266), .b(G1267), .O(G1311) );
nand2 gate503( .a(G1268), .b(G1269), .O(G1312) );

  xor2  gate1079(.a(G1271), .b(G1270), .O(gate504inter0));
  nand2 gate1080(.a(gate504inter0), .b(s_76), .O(gate504inter1));
  and2  gate1081(.a(G1271), .b(G1270), .O(gate504inter2));
  inv1  gate1082(.a(s_76), .O(gate504inter3));
  inv1  gate1083(.a(s_77), .O(gate504inter4));
  nand2 gate1084(.a(gate504inter4), .b(gate504inter3), .O(gate504inter5));
  nor2  gate1085(.a(gate504inter5), .b(gate504inter2), .O(gate504inter6));
  inv1  gate1086(.a(G1270), .O(gate504inter7));
  inv1  gate1087(.a(G1271), .O(gate504inter8));
  nand2 gate1088(.a(gate504inter8), .b(gate504inter7), .O(gate504inter9));
  nand2 gate1089(.a(s_77), .b(gate504inter3), .O(gate504inter10));
  nor2  gate1090(.a(gate504inter10), .b(gate504inter9), .O(gate504inter11));
  nor2  gate1091(.a(gate504inter11), .b(gate504inter6), .O(gate504inter12));
  nand2 gate1092(.a(gate504inter12), .b(gate504inter1), .O(G1313));
nand2 gate505( .a(G1272), .b(G1273), .O(G1314) );
nand2 gate506( .a(G1274), .b(G1275), .O(G1315) );
nand2 gate507( .a(G1276), .b(G1277), .O(G1316) );

  xor2  gate953(.a(G1279), .b(G1278), .O(gate508inter0));
  nand2 gate954(.a(gate508inter0), .b(s_58), .O(gate508inter1));
  and2  gate955(.a(G1279), .b(G1278), .O(gate508inter2));
  inv1  gate956(.a(s_58), .O(gate508inter3));
  inv1  gate957(.a(s_59), .O(gate508inter4));
  nand2 gate958(.a(gate508inter4), .b(gate508inter3), .O(gate508inter5));
  nor2  gate959(.a(gate508inter5), .b(gate508inter2), .O(gate508inter6));
  inv1  gate960(.a(G1278), .O(gate508inter7));
  inv1  gate961(.a(G1279), .O(gate508inter8));
  nand2 gate962(.a(gate508inter8), .b(gate508inter7), .O(gate508inter9));
  nand2 gate963(.a(s_59), .b(gate508inter3), .O(gate508inter10));
  nor2  gate964(.a(gate508inter10), .b(gate508inter9), .O(gate508inter11));
  nor2  gate965(.a(gate508inter11), .b(gate508inter6), .O(gate508inter12));
  nand2 gate966(.a(gate508inter12), .b(gate508inter1), .O(G1317));
nand2 gate509( .a(G1280), .b(G1281), .O(G1318) );
nand2 gate510( .a(G1282), .b(G1283), .O(G1319) );
nand2 gate511( .a(G1284), .b(G1285), .O(G1320) );
nand2 gate512( .a(G1286), .b(G1287), .O(G1321) );
nand2 gate513( .a(G1288), .b(G1289), .O(G1322) );
nand2 gate514( .a(G1290), .b(G1291), .O(G1323) );
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule