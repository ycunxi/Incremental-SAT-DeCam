module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);

input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;//RE__PI;

input s_0,s_1;//RE__ALLOW(00,01,10,11);
input s_2,s_3;//RE__ALLOW(00,01,10,11);
input s_4,s_5;//RE__ALLOW(00,01,10,11);
input s_6,s_7;//RE__ALLOW(00,01,10,11);
input s_8,s_9;//RE__ALLOW(00,01,10,11);
input s_10,s_11;//RE__ALLOW(00,01,10,11);
input s_12,s_13;//RE__ALLOW(00,01,10,11);
input s_14,s_15;//RE__ALLOW(00,01,10,11);
input s_16,s_17;//RE__ALLOW(00,01,10,11);
input s_18,s_19;//RE__ALLOW(00,01,10,11);
input s_20,s_21;//RE__ALLOW(00,01,10,11);
input s_22,s_23;//RE__ALLOW(00,01,10,11);
input s_24,s_25;//RE__ALLOW(00,01,10,11);
input s_26,s_27;//RE__ALLOW(00,01,10,11);
input s_28,s_29;//RE__ALLOW(00,01,10,11);
input s_30,s_31;//RE__ALLOW(00,01,10,11);
input s_32,s_33;//RE__ALLOW(00,01,10,11);
input s_34,s_35;//RE__ALLOW(00,01,10,11);
input s_36,s_37;//RE__ALLOW(00,01,10,11);
input s_38,s_39;//RE__ALLOW(00,01,10,11);
input s_40,s_41;//RE__ALLOW(00,01,10,11);
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;

  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate27inter0, gate27inter1, gate27inter2, gate27inter3, gate27inter4, gate27inter5, gate27inter6, gate27inter7, gate27inter8, gate27inter9, gate27inter10, gate27inter11, gate27inter12, gate212inter0, gate212inter1, gate212inter2, gate212inter3, gate212inter4, gate212inter5, gate212inter6, gate212inter7, gate212inter8, gate212inter9, gate212inter10, gate212inter11, gate212inter12, gate61inter0, gate61inter1, gate61inter2, gate61inter3, gate61inter4, gate61inter5, gate61inter6, gate61inter7, gate61inter8, gate61inter9, gate61inter10, gate61inter11, gate61inter12, gate246inter0, gate246inter1, gate246inter2, gate246inter3, gate246inter4, gate246inter5, gate246inter6, gate246inter7, gate246inter8, gate246inter9, gate246inter10, gate246inter11, gate246inter12, gate456inter0, gate456inter1, gate456inter2, gate456inter3, gate456inter4, gate456inter5, gate456inter6, gate456inter7, gate456inter8, gate456inter9, gate456inter10, gate456inter11, gate456inter12, gate106inter0, gate106inter1, gate106inter2, gate106inter3, gate106inter4, gate106inter5, gate106inter6, gate106inter7, gate106inter8, gate106inter9, gate106inter10, gate106inter11, gate106inter12, gate110inter0, gate110inter1, gate110inter2, gate110inter3, gate110inter4, gate110inter5, gate110inter6, gate110inter7, gate110inter8, gate110inter9, gate110inter10, gate110inter11, gate110inter12, gate40inter0, gate40inter1, gate40inter2, gate40inter3, gate40inter4, gate40inter5, gate40inter6, gate40inter7, gate40inter8, gate40inter9, gate40inter10, gate40inter11, gate40inter12, gate434inter0, gate434inter1, gate434inter2, gate434inter3, gate434inter4, gate434inter5, gate434inter6, gate434inter7, gate434inter8, gate434inter9, gate434inter10, gate434inter11, gate434inter12, gate149inter0, gate149inter1, gate149inter2, gate149inter3, gate149inter4, gate149inter5, gate149inter6, gate149inter7, gate149inter8, gate149inter9, gate149inter10, gate149inter11, gate149inter12, gate152inter0, gate152inter1, gate152inter2, gate152inter3, gate152inter4, gate152inter5, gate152inter6, gate152inter7, gate152inter8, gate152inter9, gate152inter10, gate152inter11, gate152inter12, gate111inter0, gate111inter1, gate111inter2, gate111inter3, gate111inter4, gate111inter5, gate111inter6, gate111inter7, gate111inter8, gate111inter9, gate111inter10, gate111inter11, gate111inter12, gate435inter0, gate435inter1, gate435inter2, gate435inter3, gate435inter4, gate435inter5, gate435inter6, gate435inter7, gate435inter8, gate435inter9, gate435inter10, gate435inter11, gate435inter12, gate183inter0, gate183inter1, gate183inter2, gate183inter3, gate183inter4, gate183inter5, gate183inter6, gate183inter7, gate183inter8, gate183inter9, gate183inter10, gate183inter11, gate183inter12, gate156inter0, gate156inter1, gate156inter2, gate156inter3, gate156inter4, gate156inter5, gate156inter6, gate156inter7, gate156inter8, gate156inter9, gate156inter10, gate156inter11, gate156inter12, gate251inter0, gate251inter1, gate251inter2, gate251inter3, gate251inter4, gate251inter5, gate251inter6, gate251inter7, gate251inter8, gate251inter9, gate251inter10, gate251inter11, gate251inter12, gate49inter0, gate49inter1, gate49inter2, gate49inter3, gate49inter4, gate49inter5, gate49inter6, gate49inter7, gate49inter8, gate49inter9, gate49inter10, gate49inter11, gate49inter12, gate128inter0, gate128inter1, gate128inter2, gate128inter3, gate128inter4, gate128inter5, gate128inter6, gate128inter7, gate128inter8, gate128inter9, gate128inter10, gate128inter11, gate128inter12, gate420inter0, gate420inter1, gate420inter2, gate420inter3, gate420inter4, gate420inter5, gate420inter6, gate420inter7, gate420inter8, gate420inter9, gate420inter10, gate420inter11, gate420inter12, gate215inter0, gate215inter1, gate215inter2, gate215inter3, gate215inter4, gate215inter5, gate215inter6, gate215inter7, gate215inter8, gate215inter9, gate215inter10, gate215inter11, gate215inter12, gate476inter0, gate476inter1, gate476inter2, gate476inter3, gate476inter4, gate476inter5, gate476inter6, gate476inter7, gate476inter8, gate476inter9, gate476inter10, gate476inter11, gate476inter12;



and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );
nand2 gate9( .a(G1), .b(G2), .O(G266) );
nand2 gate10( .a(G3), .b(G4), .O(G269) );
nand2 gate11( .a(G5), .b(G6), .O(G272) );
nand2 gate12( .a(G7), .b(G8), .O(G275) );
nand2 gate13( .a(G9), .b(G10), .O(G278) );
nand2 gate14( .a(G11), .b(G12), .O(G281) );
nand2 gate15( .a(G13), .b(G14), .O(G284) );
nand2 gate16( .a(G15), .b(G16), .O(G287) );
nand2 gate17( .a(G17), .b(G18), .O(G290) );
nand2 gate18( .a(G19), .b(G20), .O(G293) );
nand2 gate19( .a(G21), .b(G22), .O(G296) );
nand2 gate20( .a(G23), .b(G24), .O(G299) );
nand2 gate21( .a(G25), .b(G26), .O(G302) );
nand2 gate22( .a(G27), .b(G28), .O(G305) );
nand2 gate23( .a(G29), .b(G30), .O(G308) );
nand2 gate24( .a(G31), .b(G32), .O(G311) );
nand2 gate25( .a(G1), .b(G5), .O(G314) );
nand2 gate26( .a(G9), .b(G13), .O(G317) );

  xor2  gate547(.a(G6), .b(G2), .O(gate27inter0));
  nand2 gate548(.a(gate27inter0), .b(s_0), .O(gate27inter1));
  and2  gate549(.a(G6), .b(G2), .O(gate27inter2));
  inv1  gate550(.a(s_0), .O(gate27inter3));
  inv1  gate551(.a(s_1), .O(gate27inter4));
  nand2 gate552(.a(gate27inter4), .b(gate27inter3), .O(gate27inter5));
  nor2  gate553(.a(gate27inter5), .b(gate27inter2), .O(gate27inter6));
  inv1  gate554(.a(G2), .O(gate27inter7));
  inv1  gate555(.a(G6), .O(gate27inter8));
  nand2 gate556(.a(gate27inter8), .b(gate27inter7), .O(gate27inter9));
  nand2 gate557(.a(s_1), .b(gate27inter3), .O(gate27inter10));
  nor2  gate558(.a(gate27inter10), .b(gate27inter9), .O(gate27inter11));
  nor2  gate559(.a(gate27inter11), .b(gate27inter6), .O(gate27inter12));
  nand2 gate560(.a(gate27inter12), .b(gate27inter1), .O(G320));
nand2 gate28( .a(G10), .b(G14), .O(G323) );
nand2 gate29( .a(G3), .b(G7), .O(G326) );
nand2 gate30( .a(G11), .b(G15), .O(G329) );
nand2 gate31( .a(G4), .b(G8), .O(G332) );
nand2 gate32( .a(G12), .b(G16), .O(G335) );
nand2 gate33( .a(G17), .b(G21), .O(G338) );
nand2 gate34( .a(G25), .b(G29), .O(G341) );
nand2 gate35( .a(G18), .b(G22), .O(G344) );
nand2 gate36( .a(G26), .b(G30), .O(G347) );
nand2 gate37( .a(G19), .b(G23), .O(G350) );
nand2 gate38( .a(G27), .b(G31), .O(G353) );
nand2 gate39( .a(G20), .b(G24), .O(G356) );

  xor2  gate645(.a(G32), .b(G28), .O(gate40inter0));
  nand2 gate646(.a(gate40inter0), .b(s_14), .O(gate40inter1));
  and2  gate647(.a(G32), .b(G28), .O(gate40inter2));
  inv1  gate648(.a(s_14), .O(gate40inter3));
  inv1  gate649(.a(s_15), .O(gate40inter4));
  nand2 gate650(.a(gate40inter4), .b(gate40inter3), .O(gate40inter5));
  nor2  gate651(.a(gate40inter5), .b(gate40inter2), .O(gate40inter6));
  inv1  gate652(.a(G28), .O(gate40inter7));
  inv1  gate653(.a(G32), .O(gate40inter8));
  nand2 gate654(.a(gate40inter8), .b(gate40inter7), .O(gate40inter9));
  nand2 gate655(.a(s_15), .b(gate40inter3), .O(gate40inter10));
  nor2  gate656(.a(gate40inter10), .b(gate40inter9), .O(gate40inter11));
  nor2  gate657(.a(gate40inter11), .b(gate40inter6), .O(gate40inter12));
  nand2 gate658(.a(gate40inter12), .b(gate40inter1), .O(G359));
nand2 gate41( .a(G1), .b(G266), .O(G362) );
nand2 gate42( .a(G2), .b(G266), .O(G363) );
nand2 gate43( .a(G3), .b(G269), .O(G364) );
nand2 gate44( .a(G4), .b(G269), .O(G365) );
nand2 gate45( .a(G5), .b(G272), .O(G366) );
nand2 gate46( .a(G6), .b(G272), .O(G367) );
nand2 gate47( .a(G7), .b(G275), .O(G368) );
nand2 gate48( .a(G8), .b(G275), .O(G369) );

  xor2  gate771(.a(G278), .b(G9), .O(gate49inter0));
  nand2 gate772(.a(gate49inter0), .b(s_32), .O(gate49inter1));
  and2  gate773(.a(G278), .b(G9), .O(gate49inter2));
  inv1  gate774(.a(s_32), .O(gate49inter3));
  inv1  gate775(.a(s_33), .O(gate49inter4));
  nand2 gate776(.a(gate49inter4), .b(gate49inter3), .O(gate49inter5));
  nor2  gate777(.a(gate49inter5), .b(gate49inter2), .O(gate49inter6));
  inv1  gate778(.a(G9), .O(gate49inter7));
  inv1  gate779(.a(G278), .O(gate49inter8));
  nand2 gate780(.a(gate49inter8), .b(gate49inter7), .O(gate49inter9));
  nand2 gate781(.a(s_33), .b(gate49inter3), .O(gate49inter10));
  nor2  gate782(.a(gate49inter10), .b(gate49inter9), .O(gate49inter11));
  nor2  gate783(.a(gate49inter11), .b(gate49inter6), .O(gate49inter12));
  nand2 gate784(.a(gate49inter12), .b(gate49inter1), .O(G370));
nand2 gate50( .a(G10), .b(G278), .O(G371) );
nand2 gate51( .a(G11), .b(G281), .O(G372) );
nand2 gate52( .a(G12), .b(G281), .O(G373) );
nand2 gate53( .a(G13), .b(G284), .O(G374) );
nand2 gate54( .a(G14), .b(G284), .O(G375) );
nand2 gate55( .a(G15), .b(G287), .O(G376) );
nand2 gate56( .a(G16), .b(G287), .O(G377) );
nand2 gate57( .a(G17), .b(G290), .O(G378) );
nand2 gate58( .a(G18), .b(G290), .O(G379) );
nand2 gate59( .a(G19), .b(G293), .O(G380) );
nand2 gate60( .a(G20), .b(G293), .O(G381) );

  xor2  gate575(.a(G296), .b(G21), .O(gate61inter0));
  nand2 gate576(.a(gate61inter0), .b(s_4), .O(gate61inter1));
  and2  gate577(.a(G296), .b(G21), .O(gate61inter2));
  inv1  gate578(.a(s_4), .O(gate61inter3));
  inv1  gate579(.a(s_5), .O(gate61inter4));
  nand2 gate580(.a(gate61inter4), .b(gate61inter3), .O(gate61inter5));
  nor2  gate581(.a(gate61inter5), .b(gate61inter2), .O(gate61inter6));
  inv1  gate582(.a(G21), .O(gate61inter7));
  inv1  gate583(.a(G296), .O(gate61inter8));
  nand2 gate584(.a(gate61inter8), .b(gate61inter7), .O(gate61inter9));
  nand2 gate585(.a(s_5), .b(gate61inter3), .O(gate61inter10));
  nor2  gate586(.a(gate61inter10), .b(gate61inter9), .O(gate61inter11));
  nor2  gate587(.a(gate61inter11), .b(gate61inter6), .O(gate61inter12));
  nand2 gate588(.a(gate61inter12), .b(gate61inter1), .O(G382));
nand2 gate62( .a(G22), .b(G296), .O(G383) );
nand2 gate63( .a(G23), .b(G299), .O(G384) );
nand2 gate64( .a(G24), .b(G299), .O(G385) );
nand2 gate65( .a(G25), .b(G302), .O(G386) );
nand2 gate66( .a(G26), .b(G302), .O(G387) );
nand2 gate67( .a(G27), .b(G305), .O(G388) );
nand2 gate68( .a(G28), .b(G305), .O(G389) );
nand2 gate69( .a(G29), .b(G308), .O(G390) );
nand2 gate70( .a(G30), .b(G308), .O(G391) );
nand2 gate71( .a(G31), .b(G311), .O(G392) );
nand2 gate72( .a(G32), .b(G311), .O(G393) );
nand2 gate73( .a(G1), .b(G314), .O(G394) );
nand2 gate74( .a(G5), .b(G314), .O(G395) );
nand2 gate75( .a(G9), .b(G317), .O(G396) );
nand2 gate76( .a(G13), .b(G317), .O(G397) );
nand2 gate77( .a(G2), .b(G320), .O(G398) );
nand2 gate78( .a(G6), .b(G320), .O(G399) );
nand2 gate79( .a(G10), .b(G323), .O(G400) );
nand2 gate80( .a(G14), .b(G323), .O(G401) );
nand2 gate81( .a(G3), .b(G326), .O(G402) );
nand2 gate82( .a(G7), .b(G326), .O(G403) );
nand2 gate83( .a(G11), .b(G329), .O(G404) );
nand2 gate84( .a(G15), .b(G329), .O(G405) );
nand2 gate85( .a(G4), .b(G332), .O(G406) );
nand2 gate86( .a(G8), .b(G332), .O(G407) );
nand2 gate87( .a(G12), .b(G335), .O(G408) );
nand2 gate88( .a(G16), .b(G335), .O(G409) );
nand2 gate89( .a(G17), .b(G338), .O(G410) );
nand2 gate90( .a(G21), .b(G338), .O(G411) );
nand2 gate91( .a(G25), .b(G341), .O(G412) );
nand2 gate92( .a(G29), .b(G341), .O(G413) );
nand2 gate93( .a(G18), .b(G344), .O(G414) );
nand2 gate94( .a(G22), .b(G344), .O(G415) );
nand2 gate95( .a(G26), .b(G347), .O(G416) );
nand2 gate96( .a(G30), .b(G347), .O(G417) );
nand2 gate97( .a(G19), .b(G350), .O(G418) );
nand2 gate98( .a(G23), .b(G350), .O(G419) );
nand2 gate99( .a(G27), .b(G353), .O(G420) );
nand2 gate100( .a(G31), .b(G353), .O(G421) );
nand2 gate101( .a(G20), .b(G356), .O(G422) );
nand2 gate102( .a(G24), .b(G356), .O(G423) );
nand2 gate103( .a(G28), .b(G359), .O(G424) );
nand2 gate104( .a(G32), .b(G359), .O(G425) );
nand2 gate105( .a(G362), .b(G363), .O(G426) );

  xor2  gate617(.a(G365), .b(G364), .O(gate106inter0));
  nand2 gate618(.a(gate106inter0), .b(s_10), .O(gate106inter1));
  and2  gate619(.a(G365), .b(G364), .O(gate106inter2));
  inv1  gate620(.a(s_10), .O(gate106inter3));
  inv1  gate621(.a(s_11), .O(gate106inter4));
  nand2 gate622(.a(gate106inter4), .b(gate106inter3), .O(gate106inter5));
  nor2  gate623(.a(gate106inter5), .b(gate106inter2), .O(gate106inter6));
  inv1  gate624(.a(G364), .O(gate106inter7));
  inv1  gate625(.a(G365), .O(gate106inter8));
  nand2 gate626(.a(gate106inter8), .b(gate106inter7), .O(gate106inter9));
  nand2 gate627(.a(s_11), .b(gate106inter3), .O(gate106inter10));
  nor2  gate628(.a(gate106inter10), .b(gate106inter9), .O(gate106inter11));
  nor2  gate629(.a(gate106inter11), .b(gate106inter6), .O(gate106inter12));
  nand2 gate630(.a(gate106inter12), .b(gate106inter1), .O(G429));
nand2 gate107( .a(G366), .b(G367), .O(G432) );
nand2 gate108( .a(G368), .b(G369), .O(G435) );
nand2 gate109( .a(G370), .b(G371), .O(G438) );

  xor2  gate631(.a(G373), .b(G372), .O(gate110inter0));
  nand2 gate632(.a(gate110inter0), .b(s_12), .O(gate110inter1));
  and2  gate633(.a(G373), .b(G372), .O(gate110inter2));
  inv1  gate634(.a(s_12), .O(gate110inter3));
  inv1  gate635(.a(s_13), .O(gate110inter4));
  nand2 gate636(.a(gate110inter4), .b(gate110inter3), .O(gate110inter5));
  nor2  gate637(.a(gate110inter5), .b(gate110inter2), .O(gate110inter6));
  inv1  gate638(.a(G372), .O(gate110inter7));
  inv1  gate639(.a(G373), .O(gate110inter8));
  nand2 gate640(.a(gate110inter8), .b(gate110inter7), .O(gate110inter9));
  nand2 gate641(.a(s_13), .b(gate110inter3), .O(gate110inter10));
  nor2  gate642(.a(gate110inter10), .b(gate110inter9), .O(gate110inter11));
  nor2  gate643(.a(gate110inter11), .b(gate110inter6), .O(gate110inter12));
  nand2 gate644(.a(gate110inter12), .b(gate110inter1), .O(G441));

  xor2  gate701(.a(G375), .b(G374), .O(gate111inter0));
  nand2 gate702(.a(gate111inter0), .b(s_22), .O(gate111inter1));
  and2  gate703(.a(G375), .b(G374), .O(gate111inter2));
  inv1  gate704(.a(s_22), .O(gate111inter3));
  inv1  gate705(.a(s_23), .O(gate111inter4));
  nand2 gate706(.a(gate111inter4), .b(gate111inter3), .O(gate111inter5));
  nor2  gate707(.a(gate111inter5), .b(gate111inter2), .O(gate111inter6));
  inv1  gate708(.a(G374), .O(gate111inter7));
  inv1  gate709(.a(G375), .O(gate111inter8));
  nand2 gate710(.a(gate111inter8), .b(gate111inter7), .O(gate111inter9));
  nand2 gate711(.a(s_23), .b(gate111inter3), .O(gate111inter10));
  nor2  gate712(.a(gate111inter10), .b(gate111inter9), .O(gate111inter11));
  nor2  gate713(.a(gate111inter11), .b(gate111inter6), .O(gate111inter12));
  nand2 gate714(.a(gate111inter12), .b(gate111inter1), .O(G444));
nand2 gate112( .a(G376), .b(G377), .O(G447) );
nand2 gate113( .a(G378), .b(G379), .O(G450) );
nand2 gate114( .a(G380), .b(G381), .O(G453) );
nand2 gate115( .a(G382), .b(G383), .O(G456) );
nand2 gate116( .a(G384), .b(G385), .O(G459) );
nand2 gate117( .a(G386), .b(G387), .O(G462) );
nand2 gate118( .a(G388), .b(G389), .O(G465) );
nand2 gate119( .a(G390), .b(G391), .O(G468) );
nand2 gate120( .a(G392), .b(G393), .O(G471) );
nand2 gate121( .a(G394), .b(G395), .O(G474) );
nand2 gate122( .a(G396), .b(G397), .O(G477) );
nand2 gate123( .a(G398), .b(G399), .O(G480) );
nand2 gate124( .a(G400), .b(G401), .O(G483) );
nand2 gate125( .a(G402), .b(G403), .O(G486) );
nand2 gate126( .a(G404), .b(G405), .O(G489) );
nand2 gate127( .a(G406), .b(G407), .O(G492) );

  xor2  gate785(.a(G409), .b(G408), .O(gate128inter0));
  nand2 gate786(.a(gate128inter0), .b(s_34), .O(gate128inter1));
  and2  gate787(.a(G409), .b(G408), .O(gate128inter2));
  inv1  gate788(.a(s_34), .O(gate128inter3));
  inv1  gate789(.a(s_35), .O(gate128inter4));
  nand2 gate790(.a(gate128inter4), .b(gate128inter3), .O(gate128inter5));
  nor2  gate791(.a(gate128inter5), .b(gate128inter2), .O(gate128inter6));
  inv1  gate792(.a(G408), .O(gate128inter7));
  inv1  gate793(.a(G409), .O(gate128inter8));
  nand2 gate794(.a(gate128inter8), .b(gate128inter7), .O(gate128inter9));
  nand2 gate795(.a(s_35), .b(gate128inter3), .O(gate128inter10));
  nor2  gate796(.a(gate128inter10), .b(gate128inter9), .O(gate128inter11));
  nor2  gate797(.a(gate128inter11), .b(gate128inter6), .O(gate128inter12));
  nand2 gate798(.a(gate128inter12), .b(gate128inter1), .O(G495));
nand2 gate129( .a(G410), .b(G411), .O(G498) );
nand2 gate130( .a(G412), .b(G413), .O(G501) );
nand2 gate131( .a(G414), .b(G415), .O(G504) );
nand2 gate132( .a(G416), .b(G417), .O(G507) );
nand2 gate133( .a(G418), .b(G419), .O(G510) );
nand2 gate134( .a(G420), .b(G421), .O(G513) );
nand2 gate135( .a(G422), .b(G423), .O(G516) );
nand2 gate136( .a(G424), .b(G425), .O(G519) );
nand2 gate137( .a(G426), .b(G429), .O(G522) );
nand2 gate138( .a(G432), .b(G435), .O(G525) );
nand2 gate139( .a(G438), .b(G441), .O(G528) );
nand2 gate140( .a(G444), .b(G447), .O(G531) );
nand2 gate141( .a(G450), .b(G453), .O(G534) );
nand2 gate142( .a(G456), .b(G459), .O(G537) );
nand2 gate143( .a(G462), .b(G465), .O(G540) );
nand2 gate144( .a(G468), .b(G471), .O(G543) );
nand2 gate145( .a(G474), .b(G477), .O(G546) );
nand2 gate146( .a(G480), .b(G483), .O(G549) );
nand2 gate147( .a(G486), .b(G489), .O(G552) );
nand2 gate148( .a(G492), .b(G495), .O(G555) );

  xor2  gate673(.a(G501), .b(G498), .O(gate149inter0));
  nand2 gate674(.a(gate149inter0), .b(s_18), .O(gate149inter1));
  and2  gate675(.a(G501), .b(G498), .O(gate149inter2));
  inv1  gate676(.a(s_18), .O(gate149inter3));
  inv1  gate677(.a(s_19), .O(gate149inter4));
  nand2 gate678(.a(gate149inter4), .b(gate149inter3), .O(gate149inter5));
  nor2  gate679(.a(gate149inter5), .b(gate149inter2), .O(gate149inter6));
  inv1  gate680(.a(G498), .O(gate149inter7));
  inv1  gate681(.a(G501), .O(gate149inter8));
  nand2 gate682(.a(gate149inter8), .b(gate149inter7), .O(gate149inter9));
  nand2 gate683(.a(s_19), .b(gate149inter3), .O(gate149inter10));
  nor2  gate684(.a(gate149inter10), .b(gate149inter9), .O(gate149inter11));
  nor2  gate685(.a(gate149inter11), .b(gate149inter6), .O(gate149inter12));
  nand2 gate686(.a(gate149inter12), .b(gate149inter1), .O(G558));
nand2 gate150( .a(G504), .b(G507), .O(G561) );
nand2 gate151( .a(G510), .b(G513), .O(G564) );

  xor2  gate687(.a(G519), .b(G516), .O(gate152inter0));
  nand2 gate688(.a(gate152inter0), .b(s_20), .O(gate152inter1));
  and2  gate689(.a(G519), .b(G516), .O(gate152inter2));
  inv1  gate690(.a(s_20), .O(gate152inter3));
  inv1  gate691(.a(s_21), .O(gate152inter4));
  nand2 gate692(.a(gate152inter4), .b(gate152inter3), .O(gate152inter5));
  nor2  gate693(.a(gate152inter5), .b(gate152inter2), .O(gate152inter6));
  inv1  gate694(.a(G516), .O(gate152inter7));
  inv1  gate695(.a(G519), .O(gate152inter8));
  nand2 gate696(.a(gate152inter8), .b(gate152inter7), .O(gate152inter9));
  nand2 gate697(.a(s_21), .b(gate152inter3), .O(gate152inter10));
  nor2  gate698(.a(gate152inter10), .b(gate152inter9), .O(gate152inter11));
  nor2  gate699(.a(gate152inter11), .b(gate152inter6), .O(gate152inter12));
  nand2 gate700(.a(gate152inter12), .b(gate152inter1), .O(G567));
nand2 gate153( .a(G426), .b(G522), .O(G570) );
nand2 gate154( .a(G429), .b(G522), .O(G571) );
nand2 gate155( .a(G432), .b(G525), .O(G572) );

  xor2  gate743(.a(G525), .b(G435), .O(gate156inter0));
  nand2 gate744(.a(gate156inter0), .b(s_28), .O(gate156inter1));
  and2  gate745(.a(G525), .b(G435), .O(gate156inter2));
  inv1  gate746(.a(s_28), .O(gate156inter3));
  inv1  gate747(.a(s_29), .O(gate156inter4));
  nand2 gate748(.a(gate156inter4), .b(gate156inter3), .O(gate156inter5));
  nor2  gate749(.a(gate156inter5), .b(gate156inter2), .O(gate156inter6));
  inv1  gate750(.a(G435), .O(gate156inter7));
  inv1  gate751(.a(G525), .O(gate156inter8));
  nand2 gate752(.a(gate156inter8), .b(gate156inter7), .O(gate156inter9));
  nand2 gate753(.a(s_29), .b(gate156inter3), .O(gate156inter10));
  nor2  gate754(.a(gate156inter10), .b(gate156inter9), .O(gate156inter11));
  nor2  gate755(.a(gate156inter11), .b(gate156inter6), .O(gate156inter12));
  nand2 gate756(.a(gate156inter12), .b(gate156inter1), .O(G573));
nand2 gate157( .a(G438), .b(G528), .O(G574) );
nand2 gate158( .a(G441), .b(G528), .O(G575) );
nand2 gate159( .a(G444), .b(G531), .O(G576) );
nand2 gate160( .a(G447), .b(G531), .O(G577) );
nand2 gate161( .a(G450), .b(G534), .O(G578) );
nand2 gate162( .a(G453), .b(G534), .O(G579) );
nand2 gate163( .a(G456), .b(G537), .O(G580) );
nand2 gate164( .a(G459), .b(G537), .O(G581) );
nand2 gate165( .a(G462), .b(G540), .O(G582) );
nand2 gate166( .a(G465), .b(G540), .O(G583) );
nand2 gate167( .a(G468), .b(G543), .O(G584) );
nand2 gate168( .a(G471), .b(G543), .O(G585) );
nand2 gate169( .a(G474), .b(G546), .O(G586) );
nand2 gate170( .a(G477), .b(G546), .O(G587) );
nand2 gate171( .a(G480), .b(G549), .O(G588) );
nand2 gate172( .a(G483), .b(G549), .O(G589) );
nand2 gate173( .a(G486), .b(G552), .O(G590) );
nand2 gate174( .a(G489), .b(G552), .O(G591) );
nand2 gate175( .a(G492), .b(G555), .O(G592) );
nand2 gate176( .a(G495), .b(G555), .O(G593) );
nand2 gate177( .a(G498), .b(G558), .O(G594) );
nand2 gate178( .a(G501), .b(G558), .O(G595) );
nand2 gate179( .a(G504), .b(G561), .O(G596) );
nand2 gate180( .a(G507), .b(G561), .O(G597) );
nand2 gate181( .a(G510), .b(G564), .O(G598) );
nand2 gate182( .a(G513), .b(G564), .O(G599) );

  xor2  gate729(.a(G567), .b(G516), .O(gate183inter0));
  nand2 gate730(.a(gate183inter0), .b(s_26), .O(gate183inter1));
  and2  gate731(.a(G567), .b(G516), .O(gate183inter2));
  inv1  gate732(.a(s_26), .O(gate183inter3));
  inv1  gate733(.a(s_27), .O(gate183inter4));
  nand2 gate734(.a(gate183inter4), .b(gate183inter3), .O(gate183inter5));
  nor2  gate735(.a(gate183inter5), .b(gate183inter2), .O(gate183inter6));
  inv1  gate736(.a(G516), .O(gate183inter7));
  inv1  gate737(.a(G567), .O(gate183inter8));
  nand2 gate738(.a(gate183inter8), .b(gate183inter7), .O(gate183inter9));
  nand2 gate739(.a(s_27), .b(gate183inter3), .O(gate183inter10));
  nor2  gate740(.a(gate183inter10), .b(gate183inter9), .O(gate183inter11));
  nor2  gate741(.a(gate183inter11), .b(gate183inter6), .O(gate183inter12));
  nand2 gate742(.a(gate183inter12), .b(gate183inter1), .O(G600));
nand2 gate184( .a(G519), .b(G567), .O(G601) );
nand2 gate185( .a(G570), .b(G571), .O(G602) );
nand2 gate186( .a(G572), .b(G573), .O(G607) );
nand2 gate187( .a(G574), .b(G575), .O(G612) );
nand2 gate188( .a(G576), .b(G577), .O(G617) );
nand2 gate189( .a(G578), .b(G579), .O(G622) );
nand2 gate190( .a(G580), .b(G581), .O(G627) );
nand2 gate191( .a(G582), .b(G583), .O(G632) );
nand2 gate192( .a(G584), .b(G585), .O(G637) );
nand2 gate193( .a(G586), .b(G587), .O(G642) );
nand2 gate194( .a(G588), .b(G589), .O(G645) );
nand2 gate195( .a(G590), .b(G591), .O(G648) );
nand2 gate196( .a(G592), .b(G593), .O(G651) );
nand2 gate197( .a(G594), .b(G595), .O(G654) );
nand2 gate198( .a(G596), .b(G597), .O(G657) );
nand2 gate199( .a(G598), .b(G599), .O(G660) );
nand2 gate200( .a(G600), .b(G601), .O(G663) );
nand2 gate201( .a(G602), .b(G607), .O(G666) );
nand2 gate202( .a(G612), .b(G617), .O(G669) );
nand2 gate203( .a(G602), .b(G612), .O(G672) );
nand2 gate204( .a(G607), .b(G617), .O(G675) );
nand2 gate205( .a(G622), .b(G627), .O(G678) );
nand2 gate206( .a(G632), .b(G637), .O(G681) );
nand2 gate207( .a(G622), .b(G632), .O(G684) );
nand2 gate208( .a(G627), .b(G637), .O(G687) );
nand2 gate209( .a(G602), .b(G666), .O(G690) );
nand2 gate210( .a(G607), .b(G666), .O(G691) );
nand2 gate211( .a(G612), .b(G669), .O(G692) );

  xor2  gate561(.a(G669), .b(G617), .O(gate212inter0));
  nand2 gate562(.a(gate212inter0), .b(s_2), .O(gate212inter1));
  and2  gate563(.a(G669), .b(G617), .O(gate212inter2));
  inv1  gate564(.a(s_2), .O(gate212inter3));
  inv1  gate565(.a(s_3), .O(gate212inter4));
  nand2 gate566(.a(gate212inter4), .b(gate212inter3), .O(gate212inter5));
  nor2  gate567(.a(gate212inter5), .b(gate212inter2), .O(gate212inter6));
  inv1  gate568(.a(G617), .O(gate212inter7));
  inv1  gate569(.a(G669), .O(gate212inter8));
  nand2 gate570(.a(gate212inter8), .b(gate212inter7), .O(gate212inter9));
  nand2 gate571(.a(s_3), .b(gate212inter3), .O(gate212inter10));
  nor2  gate572(.a(gate212inter10), .b(gate212inter9), .O(gate212inter11));
  nor2  gate573(.a(gate212inter11), .b(gate212inter6), .O(gate212inter12));
  nand2 gate574(.a(gate212inter12), .b(gate212inter1), .O(G693));
nand2 gate213( .a(G602), .b(G672), .O(G694) );
nand2 gate214( .a(G612), .b(G672), .O(G695) );

  xor2  gate813(.a(G675), .b(G607), .O(gate215inter0));
  nand2 gate814(.a(gate215inter0), .b(s_38), .O(gate215inter1));
  and2  gate815(.a(G675), .b(G607), .O(gate215inter2));
  inv1  gate816(.a(s_38), .O(gate215inter3));
  inv1  gate817(.a(s_39), .O(gate215inter4));
  nand2 gate818(.a(gate215inter4), .b(gate215inter3), .O(gate215inter5));
  nor2  gate819(.a(gate215inter5), .b(gate215inter2), .O(gate215inter6));
  inv1  gate820(.a(G607), .O(gate215inter7));
  inv1  gate821(.a(G675), .O(gate215inter8));
  nand2 gate822(.a(gate215inter8), .b(gate215inter7), .O(gate215inter9));
  nand2 gate823(.a(s_39), .b(gate215inter3), .O(gate215inter10));
  nor2  gate824(.a(gate215inter10), .b(gate215inter9), .O(gate215inter11));
  nor2  gate825(.a(gate215inter11), .b(gate215inter6), .O(gate215inter12));
  nand2 gate826(.a(gate215inter12), .b(gate215inter1), .O(G696));
nand2 gate216( .a(G617), .b(G675), .O(G697) );
nand2 gate217( .a(G622), .b(G678), .O(G698) );
nand2 gate218( .a(G627), .b(G678), .O(G699) );
nand2 gate219( .a(G632), .b(G681), .O(G700) );
nand2 gate220( .a(G637), .b(G681), .O(G701) );
nand2 gate221( .a(G622), .b(G684), .O(G702) );
nand2 gate222( .a(G632), .b(G684), .O(G703) );
nand2 gate223( .a(G627), .b(G687), .O(G704) );
nand2 gate224( .a(G637), .b(G687), .O(G705) );
nand2 gate225( .a(G690), .b(G691), .O(G706) );
nand2 gate226( .a(G692), .b(G693), .O(G709) );
nand2 gate227( .a(G694), .b(G695), .O(G712) );
nand2 gate228( .a(G696), .b(G697), .O(G715) );
nand2 gate229( .a(G698), .b(G699), .O(G718) );
nand2 gate230( .a(G700), .b(G701), .O(G721) );
nand2 gate231( .a(G702), .b(G703), .O(G724) );
nand2 gate232( .a(G704), .b(G705), .O(G727) );
nand2 gate233( .a(G242), .b(G718), .O(G730) );
nand2 gate234( .a(G245), .b(G721), .O(G733) );
nand2 gate235( .a(G248), .b(G724), .O(G736) );
nand2 gate236( .a(G251), .b(G727), .O(G739) );
nand2 gate237( .a(G254), .b(G706), .O(G742) );
nand2 gate238( .a(G257), .b(G709), .O(G745) );
nand2 gate239( .a(G260), .b(G712), .O(G748) );
nand2 gate240( .a(G263), .b(G715), .O(G751) );
nand2 gate241( .a(G242), .b(G730), .O(G754) );
nand2 gate242( .a(G718), .b(G730), .O(G755) );
nand2 gate243( .a(G245), .b(G733), .O(G756) );
nand2 gate244( .a(G721), .b(G733), .O(G757) );
nand2 gate245( .a(G248), .b(G736), .O(G758) );

  xor2  gate589(.a(G736), .b(G724), .O(gate246inter0));
  nand2 gate590(.a(gate246inter0), .b(s_6), .O(gate246inter1));
  and2  gate591(.a(G736), .b(G724), .O(gate246inter2));
  inv1  gate592(.a(s_6), .O(gate246inter3));
  inv1  gate593(.a(s_7), .O(gate246inter4));
  nand2 gate594(.a(gate246inter4), .b(gate246inter3), .O(gate246inter5));
  nor2  gate595(.a(gate246inter5), .b(gate246inter2), .O(gate246inter6));
  inv1  gate596(.a(G724), .O(gate246inter7));
  inv1  gate597(.a(G736), .O(gate246inter8));
  nand2 gate598(.a(gate246inter8), .b(gate246inter7), .O(gate246inter9));
  nand2 gate599(.a(s_7), .b(gate246inter3), .O(gate246inter10));
  nor2  gate600(.a(gate246inter10), .b(gate246inter9), .O(gate246inter11));
  nor2  gate601(.a(gate246inter11), .b(gate246inter6), .O(gate246inter12));
  nand2 gate602(.a(gate246inter12), .b(gate246inter1), .O(G759));
nand2 gate247( .a(G251), .b(G739), .O(G760) );
nand2 gate248( .a(G727), .b(G739), .O(G761) );
nand2 gate249( .a(G254), .b(G742), .O(G762) );
nand2 gate250( .a(G706), .b(G742), .O(G763) );

  xor2  gate757(.a(G745), .b(G257), .O(gate251inter0));
  nand2 gate758(.a(gate251inter0), .b(s_30), .O(gate251inter1));
  and2  gate759(.a(G745), .b(G257), .O(gate251inter2));
  inv1  gate760(.a(s_30), .O(gate251inter3));
  inv1  gate761(.a(s_31), .O(gate251inter4));
  nand2 gate762(.a(gate251inter4), .b(gate251inter3), .O(gate251inter5));
  nor2  gate763(.a(gate251inter5), .b(gate251inter2), .O(gate251inter6));
  inv1  gate764(.a(G257), .O(gate251inter7));
  inv1  gate765(.a(G745), .O(gate251inter8));
  nand2 gate766(.a(gate251inter8), .b(gate251inter7), .O(gate251inter9));
  nand2 gate767(.a(s_31), .b(gate251inter3), .O(gate251inter10));
  nor2  gate768(.a(gate251inter10), .b(gate251inter9), .O(gate251inter11));
  nor2  gate769(.a(gate251inter11), .b(gate251inter6), .O(gate251inter12));
  nand2 gate770(.a(gate251inter12), .b(gate251inter1), .O(G764));
nand2 gate252( .a(G709), .b(G745), .O(G765) );
nand2 gate253( .a(G260), .b(G748), .O(G766) );
nand2 gate254( .a(G712), .b(G748), .O(G767) );
nand2 gate255( .a(G263), .b(G751), .O(G768) );
nand2 gate256( .a(G715), .b(G751), .O(G769) );
nand2 gate257( .a(G754), .b(G755), .O(G770) );
nand2 gate258( .a(G756), .b(G757), .O(G773) );
nand2 gate259( .a(G758), .b(G759), .O(G776) );
nand2 gate260( .a(G760), .b(G761), .O(G779) );
nand2 gate261( .a(G762), .b(G763), .O(G782) );
nand2 gate262( .a(G764), .b(G765), .O(G785) );
nand2 gate263( .a(G766), .b(G767), .O(G788) );
nand2 gate264( .a(G768), .b(G769), .O(G791) );
nand2 gate265( .a(G642), .b(G770), .O(G794) );
nand2 gate266( .a(G645), .b(G773), .O(G797) );
nand2 gate267( .a(G648), .b(G776), .O(G800) );
nand2 gate268( .a(G651), .b(G779), .O(G803) );
nand2 gate269( .a(G654), .b(G782), .O(G806) );
nand2 gate270( .a(G657), .b(G785), .O(G809) );
nand2 gate271( .a(G660), .b(G788), .O(G812) );
nand2 gate272( .a(G663), .b(G791), .O(G815) );
nand2 gate273( .a(G642), .b(G794), .O(G818) );
nand2 gate274( .a(G770), .b(G794), .O(G819) );
nand2 gate275( .a(G645), .b(G797), .O(G820) );
nand2 gate276( .a(G773), .b(G797), .O(G821) );
nand2 gate277( .a(G648), .b(G800), .O(G822) );
nand2 gate278( .a(G776), .b(G800), .O(G823) );
nand2 gate279( .a(G651), .b(G803), .O(G824) );
nand2 gate280( .a(G779), .b(G803), .O(G825) );
nand2 gate281( .a(G654), .b(G806), .O(G826) );
nand2 gate282( .a(G782), .b(G806), .O(G827) );
nand2 gate283( .a(G657), .b(G809), .O(G828) );
nand2 gate284( .a(G785), .b(G809), .O(G829) );
nand2 gate285( .a(G660), .b(G812), .O(G830) );
nand2 gate286( .a(G788), .b(G812), .O(G831) );
nand2 gate287( .a(G663), .b(G815), .O(G832) );
nand2 gate288( .a(G791), .b(G815), .O(G833) );
nand2 gate289( .a(G818), .b(G819), .O(G834) );
nand2 gate290( .a(G820), .b(G821), .O(G847) );
nand2 gate291( .a(G822), .b(G823), .O(G860) );
nand2 gate292( .a(G824), .b(G825), .O(G873) );
nand2 gate293( .a(G828), .b(G829), .O(G886) );
nand2 gate294( .a(G832), .b(G833), .O(G899) );
nand2 gate295( .a(G830), .b(G831), .O(G912) );
nand2 gate296( .a(G826), .b(G827), .O(G925) );
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );
nand2 gate387( .a(G1), .b(G1036), .O(G1132) );
nand2 gate388( .a(G2), .b(G1039), .O(G1135) );
nand2 gate389( .a(G3), .b(G1042), .O(G1138) );
nand2 gate390( .a(G4), .b(G1045), .O(G1141) );
nand2 gate391( .a(G5), .b(G1048), .O(G1144) );
nand2 gate392( .a(G6), .b(G1051), .O(G1147) );
nand2 gate393( .a(G7), .b(G1054), .O(G1150) );
nand2 gate394( .a(G8), .b(G1057), .O(G1153) );
nand2 gate395( .a(G9), .b(G1060), .O(G1156) );
nand2 gate396( .a(G10), .b(G1063), .O(G1159) );
nand2 gate397( .a(G11), .b(G1066), .O(G1162) );
nand2 gate398( .a(G12), .b(G1069), .O(G1165) );
nand2 gate399( .a(G13), .b(G1072), .O(G1168) );
nand2 gate400( .a(G14), .b(G1075), .O(G1171) );
nand2 gate401( .a(G15), .b(G1078), .O(G1174) );
nand2 gate402( .a(G16), .b(G1081), .O(G1177) );
nand2 gate403( .a(G17), .b(G1084), .O(G1180) );
nand2 gate404( .a(G18), .b(G1087), .O(G1183) );
nand2 gate405( .a(G19), .b(G1090), .O(G1186) );
nand2 gate406( .a(G20), .b(G1093), .O(G1189) );
nand2 gate407( .a(G21), .b(G1096), .O(G1192) );
nand2 gate408( .a(G22), .b(G1099), .O(G1195) );
nand2 gate409( .a(G23), .b(G1102), .O(G1198) );
nand2 gate410( .a(G24), .b(G1105), .O(G1201) );
nand2 gate411( .a(G25), .b(G1108), .O(G1204) );
nand2 gate412( .a(G26), .b(G1111), .O(G1207) );
nand2 gate413( .a(G27), .b(G1114), .O(G1210) );
nand2 gate414( .a(G28), .b(G1117), .O(G1213) );
nand2 gate415( .a(G29), .b(G1120), .O(G1216) );
nand2 gate416( .a(G30), .b(G1123), .O(G1219) );
nand2 gate417( .a(G31), .b(G1126), .O(G1222) );
nand2 gate418( .a(G32), .b(G1129), .O(G1225) );
nand2 gate419( .a(G1), .b(G1132), .O(G1228) );

  xor2  gate799(.a(G1132), .b(G1036), .O(gate420inter0));
  nand2 gate800(.a(gate420inter0), .b(s_36), .O(gate420inter1));
  and2  gate801(.a(G1132), .b(G1036), .O(gate420inter2));
  inv1  gate802(.a(s_36), .O(gate420inter3));
  inv1  gate803(.a(s_37), .O(gate420inter4));
  nand2 gate804(.a(gate420inter4), .b(gate420inter3), .O(gate420inter5));
  nor2  gate805(.a(gate420inter5), .b(gate420inter2), .O(gate420inter6));
  inv1  gate806(.a(G1036), .O(gate420inter7));
  inv1  gate807(.a(G1132), .O(gate420inter8));
  nand2 gate808(.a(gate420inter8), .b(gate420inter7), .O(gate420inter9));
  nand2 gate809(.a(s_37), .b(gate420inter3), .O(gate420inter10));
  nor2  gate810(.a(gate420inter10), .b(gate420inter9), .O(gate420inter11));
  nor2  gate811(.a(gate420inter11), .b(gate420inter6), .O(gate420inter12));
  nand2 gate812(.a(gate420inter12), .b(gate420inter1), .O(G1229));
nand2 gate421( .a(G2), .b(G1135), .O(G1230) );
nand2 gate422( .a(G1039), .b(G1135), .O(G1231) );
nand2 gate423( .a(G3), .b(G1138), .O(G1232) );
nand2 gate424( .a(G1042), .b(G1138), .O(G1233) );
nand2 gate425( .a(G4), .b(G1141), .O(G1234) );
nand2 gate426( .a(G1045), .b(G1141), .O(G1235) );
nand2 gate427( .a(G5), .b(G1144), .O(G1236) );
nand2 gate428( .a(G1048), .b(G1144), .O(G1237) );
nand2 gate429( .a(G6), .b(G1147), .O(G1238) );
nand2 gate430( .a(G1051), .b(G1147), .O(G1239) );
nand2 gate431( .a(G7), .b(G1150), .O(G1240) );
nand2 gate432( .a(G1054), .b(G1150), .O(G1241) );
nand2 gate433( .a(G8), .b(G1153), .O(G1242) );

  xor2  gate659(.a(G1153), .b(G1057), .O(gate434inter0));
  nand2 gate660(.a(gate434inter0), .b(s_16), .O(gate434inter1));
  and2  gate661(.a(G1153), .b(G1057), .O(gate434inter2));
  inv1  gate662(.a(s_16), .O(gate434inter3));
  inv1  gate663(.a(s_17), .O(gate434inter4));
  nand2 gate664(.a(gate434inter4), .b(gate434inter3), .O(gate434inter5));
  nor2  gate665(.a(gate434inter5), .b(gate434inter2), .O(gate434inter6));
  inv1  gate666(.a(G1057), .O(gate434inter7));
  inv1  gate667(.a(G1153), .O(gate434inter8));
  nand2 gate668(.a(gate434inter8), .b(gate434inter7), .O(gate434inter9));
  nand2 gate669(.a(s_17), .b(gate434inter3), .O(gate434inter10));
  nor2  gate670(.a(gate434inter10), .b(gate434inter9), .O(gate434inter11));
  nor2  gate671(.a(gate434inter11), .b(gate434inter6), .O(gate434inter12));
  nand2 gate672(.a(gate434inter12), .b(gate434inter1), .O(G1243));

  xor2  gate715(.a(G1156), .b(G9), .O(gate435inter0));
  nand2 gate716(.a(gate435inter0), .b(s_24), .O(gate435inter1));
  and2  gate717(.a(G1156), .b(G9), .O(gate435inter2));
  inv1  gate718(.a(s_24), .O(gate435inter3));
  inv1  gate719(.a(s_25), .O(gate435inter4));
  nand2 gate720(.a(gate435inter4), .b(gate435inter3), .O(gate435inter5));
  nor2  gate721(.a(gate435inter5), .b(gate435inter2), .O(gate435inter6));
  inv1  gate722(.a(G9), .O(gate435inter7));
  inv1  gate723(.a(G1156), .O(gate435inter8));
  nand2 gate724(.a(gate435inter8), .b(gate435inter7), .O(gate435inter9));
  nand2 gate725(.a(s_25), .b(gate435inter3), .O(gate435inter10));
  nor2  gate726(.a(gate435inter10), .b(gate435inter9), .O(gate435inter11));
  nor2  gate727(.a(gate435inter11), .b(gate435inter6), .O(gate435inter12));
  nand2 gate728(.a(gate435inter12), .b(gate435inter1), .O(G1244));
nand2 gate436( .a(G1060), .b(G1156), .O(G1245) );
nand2 gate437( .a(G10), .b(G1159), .O(G1246) );
nand2 gate438( .a(G1063), .b(G1159), .O(G1247) );
nand2 gate439( .a(G11), .b(G1162), .O(G1248) );
nand2 gate440( .a(G1066), .b(G1162), .O(G1249) );
nand2 gate441( .a(G12), .b(G1165), .O(G1250) );
nand2 gate442( .a(G1069), .b(G1165), .O(G1251) );
nand2 gate443( .a(G13), .b(G1168), .O(G1252) );
nand2 gate444( .a(G1072), .b(G1168), .O(G1253) );
nand2 gate445( .a(G14), .b(G1171), .O(G1254) );
nand2 gate446( .a(G1075), .b(G1171), .O(G1255) );
nand2 gate447( .a(G15), .b(G1174), .O(G1256) );
nand2 gate448( .a(G1078), .b(G1174), .O(G1257) );
nand2 gate449( .a(G16), .b(G1177), .O(G1258) );
nand2 gate450( .a(G1081), .b(G1177), .O(G1259) );
nand2 gate451( .a(G17), .b(G1180), .O(G1260) );
nand2 gate452( .a(G1084), .b(G1180), .O(G1261) );
nand2 gate453( .a(G18), .b(G1183), .O(G1262) );
nand2 gate454( .a(G1087), .b(G1183), .O(G1263) );
nand2 gate455( .a(G19), .b(G1186), .O(G1264) );

  xor2  gate603(.a(G1186), .b(G1090), .O(gate456inter0));
  nand2 gate604(.a(gate456inter0), .b(s_8), .O(gate456inter1));
  and2  gate605(.a(G1186), .b(G1090), .O(gate456inter2));
  inv1  gate606(.a(s_8), .O(gate456inter3));
  inv1  gate607(.a(s_9), .O(gate456inter4));
  nand2 gate608(.a(gate456inter4), .b(gate456inter3), .O(gate456inter5));
  nor2  gate609(.a(gate456inter5), .b(gate456inter2), .O(gate456inter6));
  inv1  gate610(.a(G1090), .O(gate456inter7));
  inv1  gate611(.a(G1186), .O(gate456inter8));
  nand2 gate612(.a(gate456inter8), .b(gate456inter7), .O(gate456inter9));
  nand2 gate613(.a(s_9), .b(gate456inter3), .O(gate456inter10));
  nor2  gate614(.a(gate456inter10), .b(gate456inter9), .O(gate456inter11));
  nor2  gate615(.a(gate456inter11), .b(gate456inter6), .O(gate456inter12));
  nand2 gate616(.a(gate456inter12), .b(gate456inter1), .O(G1265));
nand2 gate457( .a(G20), .b(G1189), .O(G1266) );
nand2 gate458( .a(G1093), .b(G1189), .O(G1267) );
nand2 gate459( .a(G21), .b(G1192), .O(G1268) );
nand2 gate460( .a(G1096), .b(G1192), .O(G1269) );
nand2 gate461( .a(G22), .b(G1195), .O(G1270) );
nand2 gate462( .a(G1099), .b(G1195), .O(G1271) );
nand2 gate463( .a(G23), .b(G1198), .O(G1272) );
nand2 gate464( .a(G1102), .b(G1198), .O(G1273) );
nand2 gate465( .a(G24), .b(G1201), .O(G1274) );
nand2 gate466( .a(G1105), .b(G1201), .O(G1275) );
nand2 gate467( .a(G25), .b(G1204), .O(G1276) );
nand2 gate468( .a(G1108), .b(G1204), .O(G1277) );
nand2 gate469( .a(G26), .b(G1207), .O(G1278) );
nand2 gate470( .a(G1111), .b(G1207), .O(G1279) );
nand2 gate471( .a(G27), .b(G1210), .O(G1280) );
nand2 gate472( .a(G1114), .b(G1210), .O(G1281) );
nand2 gate473( .a(G28), .b(G1213), .O(G1282) );
nand2 gate474( .a(G1117), .b(G1213), .O(G1283) );
nand2 gate475( .a(G29), .b(G1216), .O(G1284) );

  xor2  gate827(.a(G1216), .b(G1120), .O(gate476inter0));
  nand2 gate828(.a(gate476inter0), .b(s_40), .O(gate476inter1));
  and2  gate829(.a(G1216), .b(G1120), .O(gate476inter2));
  inv1  gate830(.a(s_40), .O(gate476inter3));
  inv1  gate831(.a(s_41), .O(gate476inter4));
  nand2 gate832(.a(gate476inter4), .b(gate476inter3), .O(gate476inter5));
  nor2  gate833(.a(gate476inter5), .b(gate476inter2), .O(gate476inter6));
  inv1  gate834(.a(G1120), .O(gate476inter7));
  inv1  gate835(.a(G1216), .O(gate476inter8));
  nand2 gate836(.a(gate476inter8), .b(gate476inter7), .O(gate476inter9));
  nand2 gate837(.a(s_41), .b(gate476inter3), .O(gate476inter10));
  nor2  gate838(.a(gate476inter10), .b(gate476inter9), .O(gate476inter11));
  nor2  gate839(.a(gate476inter11), .b(gate476inter6), .O(gate476inter12));
  nand2 gate840(.a(gate476inter12), .b(gate476inter1), .O(G1285));
nand2 gate477( .a(G30), .b(G1219), .O(G1286) );
nand2 gate478( .a(G1123), .b(G1219), .O(G1287) );
nand2 gate479( .a(G31), .b(G1222), .O(G1288) );
nand2 gate480( .a(G1126), .b(G1222), .O(G1289) );
nand2 gate481( .a(G32), .b(G1225), .O(G1290) );
nand2 gate482( .a(G1129), .b(G1225), .O(G1291) );
nand2 gate483( .a(G1228), .b(G1229), .O(G1292) );
nand2 gate484( .a(G1230), .b(G1231), .O(G1293) );
nand2 gate485( .a(G1232), .b(G1233), .O(G1294) );
nand2 gate486( .a(G1234), .b(G1235), .O(G1295) );
nand2 gate487( .a(G1236), .b(G1237), .O(G1296) );
nand2 gate488( .a(G1238), .b(G1239), .O(G1297) );
nand2 gate489( .a(G1240), .b(G1241), .O(G1298) );
nand2 gate490( .a(G1242), .b(G1243), .O(G1299) );
nand2 gate491( .a(G1244), .b(G1245), .O(G1300) );
nand2 gate492( .a(G1246), .b(G1247), .O(G1301) );
nand2 gate493( .a(G1248), .b(G1249), .O(G1302) );
nand2 gate494( .a(G1250), .b(G1251), .O(G1303) );
nand2 gate495( .a(G1252), .b(G1253), .O(G1304) );
nand2 gate496( .a(G1254), .b(G1255), .O(G1305) );
nand2 gate497( .a(G1256), .b(G1257), .O(G1306) );
nand2 gate498( .a(G1258), .b(G1259), .O(G1307) );
nand2 gate499( .a(G1260), .b(G1261), .O(G1308) );
nand2 gate500( .a(G1262), .b(G1263), .O(G1309) );
nand2 gate501( .a(G1264), .b(G1265), .O(G1310) );
nand2 gate502( .a(G1266), .b(G1267), .O(G1311) );
nand2 gate503( .a(G1268), .b(G1269), .O(G1312) );
nand2 gate504( .a(G1270), .b(G1271), .O(G1313) );
nand2 gate505( .a(G1272), .b(G1273), .O(G1314) );
nand2 gate506( .a(G1274), .b(G1275), .O(G1315) );
nand2 gate507( .a(G1276), .b(G1277), .O(G1316) );
nand2 gate508( .a(G1278), .b(G1279), .O(G1317) );
nand2 gate509( .a(G1280), .b(G1281), .O(G1318) );
nand2 gate510( .a(G1282), .b(G1283), .O(G1319) );
nand2 gate511( .a(G1284), .b(G1285), .O(G1320) );
nand2 gate512( .a(G1286), .b(G1287), .O(G1321) );
nand2 gate513( .a(G1288), .b(G1289), .O(G1322) );
nand2 gate514( .a(G1290), .b(G1291), .O(G1323) );
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule