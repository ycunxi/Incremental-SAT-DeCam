module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);

input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;//RE__PI;

input s_0,s_1;//RE__ALLOW(00,01,10,11);
input s_2,s_3;//RE__ALLOW(00,01,10,11);
input s_4,s_5;//RE__ALLOW(00,01,10,11);
input s_6,s_7;//RE__ALLOW(00,01,10,11);
input s_8,s_9;//RE__ALLOW(00,01,10,11);
input s_10,s_11;//RE__ALLOW(00,01,10,11);
input s_12,s_13;//RE__ALLOW(00,01,10,11);
input s_14,s_15;//RE__ALLOW(00,01,10,11);
input s_16,s_17;//RE__ALLOW(00,01,10,11);
input s_18,s_19;//RE__ALLOW(00,01,10,11);
input s_20,s_21;//RE__ALLOW(00,01,10,11);
input s_22,s_23;//RE__ALLOW(00,01,10,11);
input s_24,s_25;//RE__ALLOW(00,01,10,11);
input s_26,s_27;//RE__ALLOW(00,01,10,11);
input s_28,s_29;//RE__ALLOW(00,01,10,11);
input s_30,s_31;//RE__ALLOW(00,01,10,11);
input s_32,s_33;//RE__ALLOW(00,01,10,11);
input s_34,s_35;//RE__ALLOW(00,01,10,11);
input s_36,s_37;//RE__ALLOW(00,01,10,11);
input s_38,s_39;//RE__ALLOW(00,01,10,11);
input s_40,s_41;//RE__ALLOW(00,01,10,11);
input s_42,s_43;//RE__ALLOW(00,01,10,11);
input s_44,s_45;//RE__ALLOW(00,01,10,11);
input s_46,s_47;//RE__ALLOW(00,01,10,11);
input s_48,s_49;//RE__ALLOW(00,01,10,11);
input s_50,s_51;//RE__ALLOW(00,01,10,11);
input s_52,s_53;//RE__ALLOW(00,01,10,11);
input s_54,s_55;//RE__ALLOW(00,01,10,11);
input s_56,s_57;//RE__ALLOW(00,01,10,11);
input s_58,s_59;//RE__ALLOW(00,01,10,11);
input s_60,s_61;//RE__ALLOW(00,01,10,11);
input s_62,s_63;//RE__ALLOW(00,01,10,11);
input s_64,s_65;//RE__ALLOW(00,01,10,11);
input s_66,s_67;//RE__ALLOW(00,01,10,11);
input s_68,s_69;//RE__ALLOW(00,01,10,11);
input s_70,s_71;//RE__ALLOW(00,01,10,11);
input s_72,s_73;//RE__ALLOW(00,01,10,11);
input s_74,s_75;//RE__ALLOW(00,01,10,11);
input s_76,s_77;//RE__ALLOW(00,01,10,11);
input s_78,s_79;//RE__ALLOW(00,01,10,11);
input s_80,s_81;//RE__ALLOW(00,01,10,11);
input s_82,s_83;//RE__ALLOW(00,01,10,11);
input s_84,s_85;//RE__ALLOW(00,01,10,11);
input s_86,s_87;//RE__ALLOW(00,01,10,11);
input s_88,s_89;//RE__ALLOW(00,01,10,11);
input s_90,s_91;//RE__ALLOW(00,01,10,11);
input s_92,s_93;//RE__ALLOW(00,01,10,11);
input s_94,s_95;//RE__ALLOW(00,01,10,11);
input s_96,s_97;//RE__ALLOW(00,01,10,11);
input s_98,s_99;//RE__ALLOW(00,01,10,11);
input s_100,s_101;//RE__ALLOW(00,01,10,11);
input s_102,s_103;//RE__ALLOW(00,01,10,11);
input s_104,s_105;//RE__ALLOW(00,01,10,11);
input s_106,s_107;//RE__ALLOW(00,01,10,11);
input s_108,s_109;//RE__ALLOW(00,01,10,11);
input s_110,s_111;//RE__ALLOW(00,01,10,11);
input s_112,s_113;//RE__ALLOW(00,01,10,11);
input s_114,s_115;//RE__ALLOW(00,01,10,11);
input s_116,s_117;//RE__ALLOW(00,01,10,11);
input s_118,s_119;//RE__ALLOW(00,01,10,11);
input s_120,s_121;//RE__ALLOW(00,01,10,11);
input s_122,s_123;//RE__ALLOW(00,01,10,11);
input s_124,s_125;//RE__ALLOW(00,01,10,11);
input s_126,s_127;//RE__ALLOW(00,01,10,11);
input s_128,s_129;//RE__ALLOW(00,01,10,11);
input s_130,s_131;//RE__ALLOW(00,01,10,11);
input s_132,s_133;//RE__ALLOW(00,01,10,11);
input s_134,s_135;//RE__ALLOW(00,01,10,11);
input s_136,s_137;//RE__ALLOW(00,01,10,11);
input s_138,s_139;//RE__ALLOW(00,01,10,11);
input s_140,s_141;//RE__ALLOW(00,01,10,11);
input s_142,s_143;//RE__ALLOW(00,01,10,11);
input s_144,s_145;//RE__ALLOW(00,01,10,11);
input s_146,s_147;//RE__ALLOW(00,01,10,11);
input s_148,s_149;//RE__ALLOW(00,01,10,11);
input s_150,s_151;//RE__ALLOW(00,01,10,11);
input s_152,s_153;//RE__ALLOW(00,01,10,11);
input s_154,s_155;//RE__ALLOW(00,01,10,11);
input s_156,s_157;//RE__ALLOW(00,01,10,11);
input s_158,s_159;//RE__ALLOW(00,01,10,11);
input s_160,s_161;//RE__ALLOW(00,01,10,11);
input s_162,s_163;//RE__ALLOW(00,01,10,11);
input s_164,s_165;//RE__ALLOW(00,01,10,11);
input s_166,s_167;//RE__ALLOW(00,01,10,11);
input s_168,s_169;//RE__ALLOW(00,01,10,11);
input s_170,s_171;//RE__ALLOW(00,01,10,11);
input s_172,s_173;//RE__ALLOW(00,01,10,11);
input s_174,s_175;//RE__ALLOW(00,01,10,11);
input s_176,s_177;//RE__ALLOW(00,01,10,11);
input s_178,s_179;//RE__ALLOW(00,01,10,11);
input s_180,s_181;//RE__ALLOW(00,01,10,11);
input s_182,s_183;//RE__ALLOW(00,01,10,11);
input s_184,s_185;//RE__ALLOW(00,01,10,11);
input s_186,s_187;//RE__ALLOW(00,01,10,11);
input s_188,s_189;//RE__ALLOW(00,01,10,11);
input s_190,s_191;//RE__ALLOW(00,01,10,11);
input s_192,s_193;//RE__ALLOW(00,01,10,11);
input s_194,s_195;//RE__ALLOW(00,01,10,11);
input s_196,s_197;//RE__ALLOW(00,01,10,11);
input s_198,s_199;//RE__ALLOW(00,01,10,11);
input s_200,s_201;//RE__ALLOW(00,01,10,11);
input s_202,s_203;//RE__ALLOW(00,01,10,11);
input s_204,s_205;//RE__ALLOW(00,01,10,11);
input s_206,s_207;//RE__ALLOW(00,01,10,11);
input s_208,s_209;//RE__ALLOW(00,01,10,11);
input s_210,s_211;//RE__ALLOW(00,01,10,11);
input s_212,s_213;//RE__ALLOW(00,01,10,11);
input s_214,s_215;//RE__ALLOW(00,01,10,11);
input s_216,s_217;//RE__ALLOW(00,01,10,11);
input s_218,s_219;//RE__ALLOW(00,01,10,11);
input s_220,s_221;//RE__ALLOW(00,01,10,11);
input s_222,s_223;//RE__ALLOW(00,01,10,11);
input s_224,s_225;//RE__ALLOW(00,01,10,11);
input s_226,s_227;//RE__ALLOW(00,01,10,11);
input s_228,s_229;//RE__ALLOW(00,01,10,11);
input s_230,s_231;//RE__ALLOW(00,01,10,11);
input s_232,s_233;//RE__ALLOW(00,01,10,11);
input s_234,s_235;//RE__ALLOW(00,01,10,11);
input s_236,s_237;//RE__ALLOW(00,01,10,11);
input s_238,s_239;//RE__ALLOW(00,01,10,11);
input s_240,s_241;//RE__ALLOW(00,01,10,11);
input s_242,s_243;//RE__ALLOW(00,01,10,11);
input s_244,s_245;//RE__ALLOW(00,01,10,11);
input s_246,s_247;//RE__ALLOW(00,01,10,11);
input s_248,s_249;//RE__ALLOW(00,01,10,11);
input s_250,s_251;//RE__ALLOW(00,01,10,11);
input s_252,s_253;//RE__ALLOW(00,01,10,11);
input s_254,s_255;//RE__ALLOW(00,01,10,11);
input s_256,s_257;//RE__ALLOW(00,01,10,11);
input s_258,s_259;//RE__ALLOW(00,01,10,11);
input s_260,s_261;//RE__ALLOW(00,01,10,11);
input s_262,s_263;//RE__ALLOW(00,01,10,11);
input s_264,s_265;//RE__ALLOW(00,01,10,11);
input s_266,s_267;//RE__ALLOW(00,01,10,11);
input s_268,s_269;//RE__ALLOW(00,01,10,11);
input s_270,s_271;//RE__ALLOW(00,01,10,11);
input s_272,s_273;//RE__ALLOW(00,01,10,11);
input s_274,s_275;//RE__ALLOW(00,01,10,11);
input s_276,s_277;//RE__ALLOW(00,01,10,11);
input s_278,s_279;//RE__ALLOW(00,01,10,11);
input s_280,s_281;//RE__ALLOW(00,01,10,11);
input s_282,s_283;//RE__ALLOW(00,01,10,11);
input s_284,s_285;//RE__ALLOW(00,01,10,11);
input s_286,s_287;//RE__ALLOW(00,01,10,11);
input s_288,s_289;//RE__ALLOW(00,01,10,11);
input s_290,s_291;//RE__ALLOW(00,01,10,11);
input s_292,s_293;//RE__ALLOW(00,01,10,11);
input s_294,s_295;//RE__ALLOW(00,01,10,11);
input s_296,s_297;//RE__ALLOW(00,01,10,11);
input s_298,s_299;//RE__ALLOW(00,01,10,11);
input s_300,s_301;//RE__ALLOW(00,01,10,11);
input s_302,s_303;//RE__ALLOW(00,01,10,11);
input s_304,s_305;//RE__ALLOW(00,01,10,11);
input s_306,s_307;//RE__ALLOW(00,01,10,11);
input s_308,s_309;//RE__ALLOW(00,01,10,11);
input s_310,s_311;//RE__ALLOW(00,01,10,11);
input s_312,s_313;//RE__ALLOW(00,01,10,11);
input s_314,s_315;//RE__ALLOW(00,01,10,11);
input s_316,s_317;//RE__ALLOW(00,01,10,11);
input s_318,s_319;//RE__ALLOW(00,01,10,11);
input s_320,s_321;//RE__ALLOW(00,01,10,11);
input s_322,s_323;//RE__ALLOW(00,01,10,11);
input s_324,s_325;//RE__ALLOW(00,01,10,11);
input s_326,s_327;//RE__ALLOW(00,01,10,11);
input s_328,s_329;//RE__ALLOW(00,01,10,11);
input s_330,s_331;//RE__ALLOW(00,01,10,11);
input s_332,s_333;//RE__ALLOW(00,01,10,11);
input s_334,s_335;//RE__ALLOW(00,01,10,11);
input s_336,s_337;//RE__ALLOW(00,01,10,11);
input s_338,s_339;//RE__ALLOW(00,01,10,11);
input s_340,s_341;//RE__ALLOW(00,01,10,11);
input s_342,s_343;//RE__ALLOW(00,01,10,11);
input s_344,s_345;//RE__ALLOW(00,01,10,11);
input s_346,s_347;//RE__ALLOW(00,01,10,11);
input s_348,s_349;//RE__ALLOW(00,01,10,11);
input s_350,s_351;//RE__ALLOW(00,01,10,11);
input s_352,s_353;//RE__ALLOW(00,01,10,11);
input s_354,s_355;//RE__ALLOW(00,01,10,11);
input s_356,s_357;//RE__ALLOW(00,01,10,11);
input s_358,s_359;//RE__ALLOW(00,01,10,11);
input s_360,s_361;//RE__ALLOW(00,01,10,11);
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;

  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate157inter0, gate157inter1, gate157inter2, gate157inter3, gate157inter4, gate157inter5, gate157inter6, gate157inter7, gate157inter8, gate157inter9, gate157inter10, gate157inter11, gate157inter12, gate440inter0, gate440inter1, gate440inter2, gate440inter3, gate440inter4, gate440inter5, gate440inter6, gate440inter7, gate440inter8, gate440inter9, gate440inter10, gate440inter11, gate440inter12, gate489inter0, gate489inter1, gate489inter2, gate489inter3, gate489inter4, gate489inter5, gate489inter6, gate489inter7, gate489inter8, gate489inter9, gate489inter10, gate489inter11, gate489inter12, gate469inter0, gate469inter1, gate469inter2, gate469inter3, gate469inter4, gate469inter5, gate469inter6, gate469inter7, gate469inter8, gate469inter9, gate469inter10, gate469inter11, gate469inter12, gate160inter0, gate160inter1, gate160inter2, gate160inter3, gate160inter4, gate160inter5, gate160inter6, gate160inter7, gate160inter8, gate160inter9, gate160inter10, gate160inter11, gate160inter12, gate80inter0, gate80inter1, gate80inter2, gate80inter3, gate80inter4, gate80inter5, gate80inter6, gate80inter7, gate80inter8, gate80inter9, gate80inter10, gate80inter11, gate80inter12, gate75inter0, gate75inter1, gate75inter2, gate75inter3, gate75inter4, gate75inter5, gate75inter6, gate75inter7, gate75inter8, gate75inter9, gate75inter10, gate75inter11, gate75inter12, gate226inter0, gate226inter1, gate226inter2, gate226inter3, gate226inter4, gate226inter5, gate226inter6, gate226inter7, gate226inter8, gate226inter9, gate226inter10, gate226inter11, gate226inter12, gate250inter0, gate250inter1, gate250inter2, gate250inter3, gate250inter4, gate250inter5, gate250inter6, gate250inter7, gate250inter8, gate250inter9, gate250inter10, gate250inter11, gate250inter12, gate239inter0, gate239inter1, gate239inter2, gate239inter3, gate239inter4, gate239inter5, gate239inter6, gate239inter7, gate239inter8, gate239inter9, gate239inter10, gate239inter11, gate239inter12, gate451inter0, gate451inter1, gate451inter2, gate451inter3, gate451inter4, gate451inter5, gate451inter6, gate451inter7, gate451inter8, gate451inter9, gate451inter10, gate451inter11, gate451inter12, gate56inter0, gate56inter1, gate56inter2, gate56inter3, gate56inter4, gate56inter5, gate56inter6, gate56inter7, gate56inter8, gate56inter9, gate56inter10, gate56inter11, gate56inter12, gate413inter0, gate413inter1, gate413inter2, gate413inter3, gate413inter4, gate413inter5, gate413inter6, gate413inter7, gate413inter8, gate413inter9, gate413inter10, gate413inter11, gate413inter12, gate153inter0, gate153inter1, gate153inter2, gate153inter3, gate153inter4, gate153inter5, gate153inter6, gate153inter7, gate153inter8, gate153inter9, gate153inter10, gate153inter11, gate153inter12, gate39inter0, gate39inter1, gate39inter2, gate39inter3, gate39inter4, gate39inter5, gate39inter6, gate39inter7, gate39inter8, gate39inter9, gate39inter10, gate39inter11, gate39inter12, gate152inter0, gate152inter1, gate152inter2, gate152inter3, gate152inter4, gate152inter5, gate152inter6, gate152inter7, gate152inter8, gate152inter9, gate152inter10, gate152inter11, gate152inter12, gate389inter0, gate389inter1, gate389inter2, gate389inter3, gate389inter4, gate389inter5, gate389inter6, gate389inter7, gate389inter8, gate389inter9, gate389inter10, gate389inter11, gate389inter12, gate411inter0, gate411inter1, gate411inter2, gate411inter3, gate411inter4, gate411inter5, gate411inter6, gate411inter7, gate411inter8, gate411inter9, gate411inter10, gate411inter11, gate411inter12, gate443inter0, gate443inter1, gate443inter2, gate443inter3, gate443inter4, gate443inter5, gate443inter6, gate443inter7, gate443inter8, gate443inter9, gate443inter10, gate443inter11, gate443inter12, gate252inter0, gate252inter1, gate252inter2, gate252inter3, gate252inter4, gate252inter5, gate252inter6, gate252inter7, gate252inter8, gate252inter9, gate252inter10, gate252inter11, gate252inter12, gate82inter0, gate82inter1, gate82inter2, gate82inter3, gate82inter4, gate82inter5, gate82inter6, gate82inter7, gate82inter8, gate82inter9, gate82inter10, gate82inter11, gate82inter12, gate91inter0, gate91inter1, gate91inter2, gate91inter3, gate91inter4, gate91inter5, gate91inter6, gate91inter7, gate91inter8, gate91inter9, gate91inter10, gate91inter11, gate91inter12, gate207inter0, gate207inter1, gate207inter2, gate207inter3, gate207inter4, gate207inter5, gate207inter6, gate207inter7, gate207inter8, gate207inter9, gate207inter10, gate207inter11, gate207inter12, gate125inter0, gate125inter1, gate125inter2, gate125inter3, gate125inter4, gate125inter5, gate125inter6, gate125inter7, gate125inter8, gate125inter9, gate125inter10, gate125inter11, gate125inter12, gate434inter0, gate434inter1, gate434inter2, gate434inter3, gate434inter4, gate434inter5, gate434inter6, gate434inter7, gate434inter8, gate434inter9, gate434inter10, gate434inter11, gate434inter12, gate289inter0, gate289inter1, gate289inter2, gate289inter3, gate289inter4, gate289inter5, gate289inter6, gate289inter7, gate289inter8, gate289inter9, gate289inter10, gate289inter11, gate289inter12, gate111inter0, gate111inter1, gate111inter2, gate111inter3, gate111inter4, gate111inter5, gate111inter6, gate111inter7, gate111inter8, gate111inter9, gate111inter10, gate111inter11, gate111inter12, gate436inter0, gate436inter1, gate436inter2, gate436inter3, gate436inter4, gate436inter5, gate436inter6, gate436inter7, gate436inter8, gate436inter9, gate436inter10, gate436inter11, gate436inter12, gate70inter0, gate70inter1, gate70inter2, gate70inter3, gate70inter4, gate70inter5, gate70inter6, gate70inter7, gate70inter8, gate70inter9, gate70inter10, gate70inter11, gate70inter12, gate282inter0, gate282inter1, gate282inter2, gate282inter3, gate282inter4, gate282inter5, gate282inter6, gate282inter7, gate282inter8, gate282inter9, gate282inter10, gate282inter11, gate282inter12, gate280inter0, gate280inter1, gate280inter2, gate280inter3, gate280inter4, gate280inter5, gate280inter6, gate280inter7, gate280inter8, gate280inter9, gate280inter10, gate280inter11, gate280inter12, gate24inter0, gate24inter1, gate24inter2, gate24inter3, gate24inter4, gate24inter5, gate24inter6, gate24inter7, gate24inter8, gate24inter9, gate24inter10, gate24inter11, gate24inter12, gate9inter0, gate9inter1, gate9inter2, gate9inter3, gate9inter4, gate9inter5, gate9inter6, gate9inter7, gate9inter8, gate9inter9, gate9inter10, gate9inter11, gate9inter12, gate199inter0, gate199inter1, gate199inter2, gate199inter3, gate199inter4, gate199inter5, gate199inter6, gate199inter7, gate199inter8, gate199inter9, gate199inter10, gate199inter11, gate199inter12, gate67inter0, gate67inter1, gate67inter2, gate67inter3, gate67inter4, gate67inter5, gate67inter6, gate67inter7, gate67inter8, gate67inter9, gate67inter10, gate67inter11, gate67inter12, gate185inter0, gate185inter1, gate185inter2, gate185inter3, gate185inter4, gate185inter5, gate185inter6, gate185inter7, gate185inter8, gate185inter9, gate185inter10, gate185inter11, gate185inter12, gate400inter0, gate400inter1, gate400inter2, gate400inter3, gate400inter4, gate400inter5, gate400inter6, gate400inter7, gate400inter8, gate400inter9, gate400inter10, gate400inter11, gate400inter12, gate223inter0, gate223inter1, gate223inter2, gate223inter3, gate223inter4, gate223inter5, gate223inter6, gate223inter7, gate223inter8, gate223inter9, gate223inter10, gate223inter11, gate223inter12, gate161inter0, gate161inter1, gate161inter2, gate161inter3, gate161inter4, gate161inter5, gate161inter6, gate161inter7, gate161inter8, gate161inter9, gate161inter10, gate161inter11, gate161inter12, gate265inter0, gate265inter1, gate265inter2, gate265inter3, gate265inter4, gate265inter5, gate265inter6, gate265inter7, gate265inter8, gate265inter9, gate265inter10, gate265inter11, gate265inter12, gate86inter0, gate86inter1, gate86inter2, gate86inter3, gate86inter4, gate86inter5, gate86inter6, gate86inter7, gate86inter8, gate86inter9, gate86inter10, gate86inter11, gate86inter12, gate15inter0, gate15inter1, gate15inter2, gate15inter3, gate15inter4, gate15inter5, gate15inter6, gate15inter7, gate15inter8, gate15inter9, gate15inter10, gate15inter11, gate15inter12, gate134inter0, gate134inter1, gate134inter2, gate134inter3, gate134inter4, gate134inter5, gate134inter6, gate134inter7, gate134inter8, gate134inter9, gate134inter10, gate134inter11, gate134inter12, gate145inter0, gate145inter1, gate145inter2, gate145inter3, gate145inter4, gate145inter5, gate145inter6, gate145inter7, gate145inter8, gate145inter9, gate145inter10, gate145inter11, gate145inter12, gate512inter0, gate512inter1, gate512inter2, gate512inter3, gate512inter4, gate512inter5, gate512inter6, gate512inter7, gate512inter8, gate512inter9, gate512inter10, gate512inter11, gate512inter12, gate391inter0, gate391inter1, gate391inter2, gate391inter3, gate391inter4, gate391inter5, gate391inter6, gate391inter7, gate391inter8, gate391inter9, gate391inter10, gate391inter11, gate391inter12, gate191inter0, gate191inter1, gate191inter2, gate191inter3, gate191inter4, gate191inter5, gate191inter6, gate191inter7, gate191inter8, gate191inter9, gate191inter10, gate191inter11, gate191inter12, gate500inter0, gate500inter1, gate500inter2, gate500inter3, gate500inter4, gate500inter5, gate500inter6, gate500inter7, gate500inter8, gate500inter9, gate500inter10, gate500inter11, gate500inter12, gate419inter0, gate419inter1, gate419inter2, gate419inter3, gate419inter4, gate419inter5, gate419inter6, gate419inter7, gate419inter8, gate419inter9, gate419inter10, gate419inter11, gate419inter12, gate248inter0, gate248inter1, gate248inter2, gate248inter3, gate248inter4, gate248inter5, gate248inter6, gate248inter7, gate248inter8, gate248inter9, gate248inter10, gate248inter11, gate248inter12, gate18inter0, gate18inter1, gate18inter2, gate18inter3, gate18inter4, gate18inter5, gate18inter6, gate18inter7, gate18inter8, gate18inter9, gate18inter10, gate18inter11, gate18inter12, gate225inter0, gate225inter1, gate225inter2, gate225inter3, gate225inter4, gate225inter5, gate225inter6, gate225inter7, gate225inter8, gate225inter9, gate225inter10, gate225inter11, gate225inter12, gate427inter0, gate427inter1, gate427inter2, gate427inter3, gate427inter4, gate427inter5, gate427inter6, gate427inter7, gate427inter8, gate427inter9, gate427inter10, gate427inter11, gate427inter12, gate42inter0, gate42inter1, gate42inter2, gate42inter3, gate42inter4, gate42inter5, gate42inter6, gate42inter7, gate42inter8, gate42inter9, gate42inter10, gate42inter11, gate42inter12, gate21inter0, gate21inter1, gate21inter2, gate21inter3, gate21inter4, gate21inter5, gate21inter6, gate21inter7, gate21inter8, gate21inter9, gate21inter10, gate21inter11, gate21inter12, gate409inter0, gate409inter1, gate409inter2, gate409inter3, gate409inter4, gate409inter5, gate409inter6, gate409inter7, gate409inter8, gate409inter9, gate409inter10, gate409inter11, gate409inter12, gate188inter0, gate188inter1, gate188inter2, gate188inter3, gate188inter4, gate188inter5, gate188inter6, gate188inter7, gate188inter8, gate188inter9, gate188inter10, gate188inter11, gate188inter12, gate420inter0, gate420inter1, gate420inter2, gate420inter3, gate420inter4, gate420inter5, gate420inter6, gate420inter7, gate420inter8, gate420inter9, gate420inter10, gate420inter11, gate420inter12, gate429inter0, gate429inter1, gate429inter2, gate429inter3, gate429inter4, gate429inter5, gate429inter6, gate429inter7, gate429inter8, gate429inter9, gate429inter10, gate429inter11, gate429inter12, gate168inter0, gate168inter1, gate168inter2, gate168inter3, gate168inter4, gate168inter5, gate168inter6, gate168inter7, gate168inter8, gate168inter9, gate168inter10, gate168inter11, gate168inter12, gate399inter0, gate399inter1, gate399inter2, gate399inter3, gate399inter4, gate399inter5, gate399inter6, gate399inter7, gate399inter8, gate399inter9, gate399inter10, gate399inter11, gate399inter12, gate69inter0, gate69inter1, gate69inter2, gate69inter3, gate69inter4, gate69inter5, gate69inter6, gate69inter7, gate69inter8, gate69inter9, gate69inter10, gate69inter11, gate69inter12, gate163inter0, gate163inter1, gate163inter2, gate163inter3, gate163inter4, gate163inter5, gate163inter6, gate163inter7, gate163inter8, gate163inter9, gate163inter10, gate163inter11, gate163inter12, gate267inter0, gate267inter1, gate267inter2, gate267inter3, gate267inter4, gate267inter5, gate267inter6, gate267inter7, gate267inter8, gate267inter9, gate267inter10, gate267inter11, gate267inter12, gate27inter0, gate27inter1, gate27inter2, gate27inter3, gate27inter4, gate27inter5, gate27inter6, gate27inter7, gate27inter8, gate27inter9, gate27inter10, gate27inter11, gate27inter12, gate460inter0, gate460inter1, gate460inter2, gate460inter3, gate460inter4, gate460inter5, gate460inter6, gate460inter7, gate460inter8, gate460inter9, gate460inter10, gate460inter11, gate460inter12, gate240inter0, gate240inter1, gate240inter2, gate240inter3, gate240inter4, gate240inter5, gate240inter6, gate240inter7, gate240inter8, gate240inter9, gate240inter10, gate240inter11, gate240inter12, gate116inter0, gate116inter1, gate116inter2, gate116inter3, gate116inter4, gate116inter5, gate116inter6, gate116inter7, gate116inter8, gate116inter9, gate116inter10, gate116inter11, gate116inter12, gate259inter0, gate259inter1, gate259inter2, gate259inter3, gate259inter4, gate259inter5, gate259inter6, gate259inter7, gate259inter8, gate259inter9, gate259inter10, gate259inter11, gate259inter12, gate46inter0, gate46inter1, gate46inter2, gate46inter3, gate46inter4, gate46inter5, gate46inter6, gate46inter7, gate46inter8, gate46inter9, gate46inter10, gate46inter11, gate46inter12, gate484inter0, gate484inter1, gate484inter2, gate484inter3, gate484inter4, gate484inter5, gate484inter6, gate484inter7, gate484inter8, gate484inter9, gate484inter10, gate484inter11, gate484inter12, gate20inter0, gate20inter1, gate20inter2, gate20inter3, gate20inter4, gate20inter5, gate20inter6, gate20inter7, gate20inter8, gate20inter9, gate20inter10, gate20inter11, gate20inter12, gate40inter0, gate40inter1, gate40inter2, gate40inter3, gate40inter4, gate40inter5, gate40inter6, gate40inter7, gate40inter8, gate40inter9, gate40inter10, gate40inter11, gate40inter12, gate97inter0, gate97inter1, gate97inter2, gate97inter3, gate97inter4, gate97inter5, gate97inter6, gate97inter7, gate97inter8, gate97inter9, gate97inter10, gate97inter11, gate97inter12, gate506inter0, gate506inter1, gate506inter2, gate506inter3, gate506inter4, gate506inter5, gate506inter6, gate506inter7, gate506inter8, gate506inter9, gate506inter10, gate506inter11, gate506inter12, gate118inter0, gate118inter1, gate118inter2, gate118inter3, gate118inter4, gate118inter5, gate118inter6, gate118inter7, gate118inter8, gate118inter9, gate118inter10, gate118inter11, gate118inter12, gate10inter0, gate10inter1, gate10inter2, gate10inter3, gate10inter4, gate10inter5, gate10inter6, gate10inter7, gate10inter8, gate10inter9, gate10inter10, gate10inter11, gate10inter12, gate261inter0, gate261inter1, gate261inter2, gate261inter3, gate261inter4, gate261inter5, gate261inter6, gate261inter7, gate261inter8, gate261inter9, gate261inter10, gate261inter11, gate261inter12, gate35inter0, gate35inter1, gate35inter2, gate35inter3, gate35inter4, gate35inter5, gate35inter6, gate35inter7, gate35inter8, gate35inter9, gate35inter10, gate35inter11, gate35inter12, gate109inter0, gate109inter1, gate109inter2, gate109inter3, gate109inter4, gate109inter5, gate109inter6, gate109inter7, gate109inter8, gate109inter9, gate109inter10, gate109inter11, gate109inter12, gate423inter0, gate423inter1, gate423inter2, gate423inter3, gate423inter4, gate423inter5, gate423inter6, gate423inter7, gate423inter8, gate423inter9, gate423inter10, gate423inter11, gate423inter12, gate497inter0, gate497inter1, gate497inter2, gate497inter3, gate497inter4, gate497inter5, gate497inter6, gate497inter7, gate497inter8, gate497inter9, gate497inter10, gate497inter11, gate497inter12, gate96inter0, gate96inter1, gate96inter2, gate96inter3, gate96inter4, gate96inter5, gate96inter6, gate96inter7, gate96inter8, gate96inter9, gate96inter10, gate96inter11, gate96inter12, gate88inter0, gate88inter1, gate88inter2, gate88inter3, gate88inter4, gate88inter5, gate88inter6, gate88inter7, gate88inter8, gate88inter9, gate88inter10, gate88inter11, gate88inter12, gate238inter0, gate238inter1, gate238inter2, gate238inter3, gate238inter4, gate238inter5, gate238inter6, gate238inter7, gate238inter8, gate238inter9, gate238inter10, gate238inter11, gate238inter12, gate235inter0, gate235inter1, gate235inter2, gate235inter3, gate235inter4, gate235inter5, gate235inter6, gate235inter7, gate235inter8, gate235inter9, gate235inter10, gate235inter11, gate235inter12, gate251inter0, gate251inter1, gate251inter2, gate251inter3, gate251inter4, gate251inter5, gate251inter6, gate251inter7, gate251inter8, gate251inter9, gate251inter10, gate251inter11, gate251inter12, gate147inter0, gate147inter1, gate147inter2, gate147inter3, gate147inter4, gate147inter5, gate147inter6, gate147inter7, gate147inter8, gate147inter9, gate147inter10, gate147inter11, gate147inter12, gate465inter0, gate465inter1, gate465inter2, gate465inter3, gate465inter4, gate465inter5, gate465inter6, gate465inter7, gate465inter8, gate465inter9, gate465inter10, gate465inter11, gate465inter12, gate22inter0, gate22inter1, gate22inter2, gate22inter3, gate22inter4, gate22inter5, gate22inter6, gate22inter7, gate22inter8, gate22inter9, gate22inter10, gate22inter11, gate22inter12, gate61inter0, gate61inter1, gate61inter2, gate61inter3, gate61inter4, gate61inter5, gate61inter6, gate61inter7, gate61inter8, gate61inter9, gate61inter10, gate61inter11, gate61inter12, gate276inter0, gate276inter1, gate276inter2, gate276inter3, gate276inter4, gate276inter5, gate276inter6, gate276inter7, gate276inter8, gate276inter9, gate276inter10, gate276inter11, gate276inter12, gate43inter0, gate43inter1, gate43inter2, gate43inter3, gate43inter4, gate43inter5, gate43inter6, gate43inter7, gate43inter8, gate43inter9, gate43inter10, gate43inter11, gate43inter12, gate230inter0, gate230inter1, gate230inter2, gate230inter3, gate230inter4, gate230inter5, gate230inter6, gate230inter7, gate230inter8, gate230inter9, gate230inter10, gate230inter11, gate230inter12, gate492inter0, gate492inter1, gate492inter2, gate492inter3, gate492inter4, gate492inter5, gate492inter6, gate492inter7, gate492inter8, gate492inter9, gate492inter10, gate492inter11, gate492inter12, gate452inter0, gate452inter1, gate452inter2, gate452inter3, gate452inter4, gate452inter5, gate452inter6, gate452inter7, gate452inter8, gate452inter9, gate452inter10, gate452inter11, gate452inter12, gate285inter0, gate285inter1, gate285inter2, gate285inter3, gate285inter4, gate285inter5, gate285inter6, gate285inter7, gate285inter8, gate285inter9, gate285inter10, gate285inter11, gate285inter12, gate120inter0, gate120inter1, gate120inter2, gate120inter3, gate120inter4, gate120inter5, gate120inter6, gate120inter7, gate120inter8, gate120inter9, gate120inter10, gate120inter11, gate120inter12, gate455inter0, gate455inter1, gate455inter2, gate455inter3, gate455inter4, gate455inter5, gate455inter6, gate455inter7, gate455inter8, gate455inter9, gate455inter10, gate455inter11, gate455inter12, gate425inter0, gate425inter1, gate425inter2, gate425inter3, gate425inter4, gate425inter5, gate425inter6, gate425inter7, gate425inter8, gate425inter9, gate425inter10, gate425inter11, gate425inter12, gate117inter0, gate117inter1, gate117inter2, gate117inter3, gate117inter4, gate117inter5, gate117inter6, gate117inter7, gate117inter8, gate117inter9, gate117inter10, gate117inter11, gate117inter12, gate467inter0, gate467inter1, gate467inter2, gate467inter3, gate467inter4, gate467inter5, gate467inter6, gate467inter7, gate467inter8, gate467inter9, gate467inter10, gate467inter11, gate467inter12, gate28inter0, gate28inter1, gate28inter2, gate28inter3, gate28inter4, gate28inter5, gate28inter6, gate28inter7, gate28inter8, gate28inter9, gate28inter10, gate28inter11, gate28inter12, gate139inter0, gate139inter1, gate139inter2, gate139inter3, gate139inter4, gate139inter5, gate139inter6, gate139inter7, gate139inter8, gate139inter9, gate139inter10, gate139inter11, gate139inter12, gate93inter0, gate93inter1, gate93inter2, gate93inter3, gate93inter4, gate93inter5, gate93inter6, gate93inter7, gate93inter8, gate93inter9, gate93inter10, gate93inter11, gate93inter12, gate213inter0, gate213inter1, gate213inter2, gate213inter3, gate213inter4, gate213inter5, gate213inter6, gate213inter7, gate213inter8, gate213inter9, gate213inter10, gate213inter11, gate213inter12, gate217inter0, gate217inter1, gate217inter2, gate217inter3, gate217inter4, gate217inter5, gate217inter6, gate217inter7, gate217inter8, gate217inter9, gate217inter10, gate217inter11, gate217inter12, gate23inter0, gate23inter1, gate23inter2, gate23inter3, gate23inter4, gate23inter5, gate23inter6, gate23inter7, gate23inter8, gate23inter9, gate23inter10, gate23inter11, gate23inter12, gate143inter0, gate143inter1, gate143inter2, gate143inter3, gate143inter4, gate143inter5, gate143inter6, gate143inter7, gate143inter8, gate143inter9, gate143inter10, gate143inter11, gate143inter12, gate73inter0, gate73inter1, gate73inter2, gate73inter3, gate73inter4, gate73inter5, gate73inter6, gate73inter7, gate73inter8, gate73inter9, gate73inter10, gate73inter11, gate73inter12, gate479inter0, gate479inter1, gate479inter2, gate479inter3, gate479inter4, gate479inter5, gate479inter6, gate479inter7, gate479inter8, gate479inter9, gate479inter10, gate479inter11, gate479inter12, gate504inter0, gate504inter1, gate504inter2, gate504inter3, gate504inter4, gate504inter5, gate504inter6, gate504inter7, gate504inter8, gate504inter9, gate504inter10, gate504inter11, gate504inter12, gate128inter0, gate128inter1, gate128inter2, gate128inter3, gate128inter4, gate128inter5, gate128inter6, gate128inter7, gate128inter8, gate128inter9, gate128inter10, gate128inter11, gate128inter12, gate137inter0, gate137inter1, gate137inter2, gate137inter3, gate137inter4, gate137inter5, gate137inter6, gate137inter7, gate137inter8, gate137inter9, gate137inter10, gate137inter11, gate137inter12, gate16inter0, gate16inter1, gate16inter2, gate16inter3, gate16inter4, gate16inter5, gate16inter6, gate16inter7, gate16inter8, gate16inter9, gate16inter10, gate16inter11, gate16inter12, gate214inter0, gate214inter1, gate214inter2, gate214inter3, gate214inter4, gate214inter5, gate214inter6, gate214inter7, gate214inter8, gate214inter9, gate214inter10, gate214inter11, gate214inter12, gate174inter0, gate174inter1, gate174inter2, gate174inter3, gate174inter4, gate174inter5, gate174inter6, gate174inter7, gate174inter8, gate174inter9, gate174inter10, gate174inter11, gate174inter12, gate189inter0, gate189inter1, gate189inter2, gate189inter3, gate189inter4, gate189inter5, gate189inter6, gate189inter7, gate189inter8, gate189inter9, gate189inter10, gate189inter11, gate189inter12, gate167inter0, gate167inter1, gate167inter2, gate167inter3, gate167inter4, gate167inter5, gate167inter6, gate167inter7, gate167inter8, gate167inter9, gate167inter10, gate167inter11, gate167inter12, gate84inter0, gate84inter1, gate84inter2, gate84inter3, gate84inter4, gate84inter5, gate84inter6, gate84inter7, gate84inter8, gate84inter9, gate84inter10, gate84inter11, gate84inter12, gate509inter0, gate509inter1, gate509inter2, gate509inter3, gate509inter4, gate509inter5, gate509inter6, gate509inter7, gate509inter8, gate509inter9, gate509inter10, gate509inter11, gate509inter12, gate154inter0, gate154inter1, gate154inter2, gate154inter3, gate154inter4, gate154inter5, gate154inter6, gate154inter7, gate154inter8, gate154inter9, gate154inter10, gate154inter11, gate154inter12, gate229inter0, gate229inter1, gate229inter2, gate229inter3, gate229inter4, gate229inter5, gate229inter6, gate229inter7, gate229inter8, gate229inter9, gate229inter10, gate229inter11, gate229inter12, gate74inter0, gate74inter1, gate74inter2, gate74inter3, gate74inter4, gate74inter5, gate74inter6, gate74inter7, gate74inter8, gate74inter9, gate74inter10, gate74inter11, gate74inter12, gate41inter0, gate41inter1, gate41inter2, gate41inter3, gate41inter4, gate41inter5, gate41inter6, gate41inter7, gate41inter8, gate41inter9, gate41inter10, gate41inter11, gate41inter12, gate186inter0, gate186inter1, gate186inter2, gate186inter3, gate186inter4, gate186inter5, gate186inter6, gate186inter7, gate186inter8, gate186inter9, gate186inter10, gate186inter11, gate186inter12, gate11inter0, gate11inter1, gate11inter2, gate11inter3, gate11inter4, gate11inter5, gate11inter6, gate11inter7, gate11inter8, gate11inter9, gate11inter10, gate11inter11, gate11inter12, gate262inter0, gate262inter1, gate262inter2, gate262inter3, gate262inter4, gate262inter5, gate262inter6, gate262inter7, gate262inter8, gate262inter9, gate262inter10, gate262inter11, gate262inter12, gate433inter0, gate433inter1, gate433inter2, gate433inter3, gate433inter4, gate433inter5, gate433inter6, gate433inter7, gate433inter8, gate433inter9, gate433inter10, gate433inter11, gate433inter12, gate114inter0, gate114inter1, gate114inter2, gate114inter3, gate114inter4, gate114inter5, gate114inter6, gate114inter7, gate114inter8, gate114inter9, gate114inter10, gate114inter11, gate114inter12, gate477inter0, gate477inter1, gate477inter2, gate477inter3, gate477inter4, gate477inter5, gate477inter6, gate477inter7, gate477inter8, gate477inter9, gate477inter10, gate477inter11, gate477inter12, gate64inter0, gate64inter1, gate64inter2, gate64inter3, gate64inter4, gate64inter5, gate64inter6, gate64inter7, gate64inter8, gate64inter9, gate64inter10, gate64inter11, gate64inter12, gate119inter0, gate119inter1, gate119inter2, gate119inter3, gate119inter4, gate119inter5, gate119inter6, gate119inter7, gate119inter8, gate119inter9, gate119inter10, gate119inter11, gate119inter12, gate87inter0, gate87inter1, gate87inter2, gate87inter3, gate87inter4, gate87inter5, gate87inter6, gate87inter7, gate87inter8, gate87inter9, gate87inter10, gate87inter11, gate87inter12, gate454inter0, gate454inter1, gate454inter2, gate454inter3, gate454inter4, gate454inter5, gate454inter6, gate454inter7, gate454inter8, gate454inter9, gate454inter10, gate454inter11, gate454inter12, gate236inter0, gate236inter1, gate236inter2, gate236inter3, gate236inter4, gate236inter5, gate236inter6, gate236inter7, gate236inter8, gate236inter9, gate236inter10, gate236inter11, gate236inter12, gate209inter0, gate209inter1, gate209inter2, gate209inter3, gate209inter4, gate209inter5, gate209inter6, gate209inter7, gate209inter8, gate209inter9, gate209inter10, gate209inter11, gate209inter12, gate244inter0, gate244inter1, gate244inter2, gate244inter3, gate244inter4, gate244inter5, gate244inter6, gate244inter7, gate244inter8, gate244inter9, gate244inter10, gate244inter11, gate244inter12, gate107inter0, gate107inter1, gate107inter2, gate107inter3, gate107inter4, gate107inter5, gate107inter6, gate107inter7, gate107inter8, gate107inter9, gate107inter10, gate107inter11, gate107inter12, gate216inter0, gate216inter1, gate216inter2, gate216inter3, gate216inter4, gate216inter5, gate216inter6, gate216inter7, gate216inter8, gate216inter9, gate216inter10, gate216inter11, gate216inter12, gate275inter0, gate275inter1, gate275inter2, gate275inter3, gate275inter4, gate275inter5, gate275inter6, gate275inter7, gate275inter8, gate275inter9, gate275inter10, gate275inter11, gate275inter12, gate164inter0, gate164inter1, gate164inter2, gate164inter3, gate164inter4, gate164inter5, gate164inter6, gate164inter7, gate164inter8, gate164inter9, gate164inter10, gate164inter11, gate164inter12, gate392inter0, gate392inter1, gate392inter2, gate392inter3, gate392inter4, gate392inter5, gate392inter6, gate392inter7, gate392inter8, gate392inter9, gate392inter10, gate392inter11, gate392inter12, gate482inter0, gate482inter1, gate482inter2, gate482inter3, gate482inter4, gate482inter5, gate482inter6, gate482inter7, gate482inter8, gate482inter9, gate482inter10, gate482inter11, gate482inter12, gate181inter0, gate181inter1, gate181inter2, gate181inter3, gate181inter4, gate181inter5, gate181inter6, gate181inter7, gate181inter8, gate181inter9, gate181inter10, gate181inter11, gate181inter12, gate410inter0, gate410inter1, gate410inter2, gate410inter3, gate410inter4, gate410inter5, gate410inter6, gate410inter7, gate410inter8, gate410inter9, gate410inter10, gate410inter11, gate410inter12, gate58inter0, gate58inter1, gate58inter2, gate58inter3, gate58inter4, gate58inter5, gate58inter6, gate58inter7, gate58inter8, gate58inter9, gate58inter10, gate58inter11, gate58inter12, gate278inter0, gate278inter1, gate278inter2, gate278inter3, gate278inter4, gate278inter5, gate278inter6, gate278inter7, gate278inter8, gate278inter9, gate278inter10, gate278inter11, gate278inter12, gate100inter0, gate100inter1, gate100inter2, gate100inter3, gate100inter4, gate100inter5, gate100inter6, gate100inter7, gate100inter8, gate100inter9, gate100inter10, gate100inter11, gate100inter12, gate461inter0, gate461inter1, gate461inter2, gate461inter3, gate461inter4, gate461inter5, gate461inter6, gate461inter7, gate461inter8, gate461inter9, gate461inter10, gate461inter11, gate461inter12, gate192inter0, gate192inter1, gate192inter2, gate192inter3, gate192inter4, gate192inter5, gate192inter6, gate192inter7, gate192inter8, gate192inter9, gate192inter10, gate192inter11, gate192inter12, gate173inter0, gate173inter1, gate173inter2, gate173inter3, gate173inter4, gate173inter5, gate173inter6, gate173inter7, gate173inter8, gate173inter9, gate173inter10, gate173inter11, gate173inter12, gate98inter0, gate98inter1, gate98inter2, gate98inter3, gate98inter4, gate98inter5, gate98inter6, gate98inter7, gate98inter8, gate98inter9, gate98inter10, gate98inter11, gate98inter12, gate444inter0, gate444inter1, gate444inter2, gate444inter3, gate444inter4, gate444inter5, gate444inter6, gate444inter7, gate444inter8, gate444inter9, gate444inter10, gate444inter11, gate444inter12, gate150inter0, gate150inter1, gate150inter2, gate150inter3, gate150inter4, gate150inter5, gate150inter6, gate150inter7, gate150inter8, gate150inter9, gate150inter10, gate150inter11, gate150inter12, gate151inter0, gate151inter1, gate151inter2, gate151inter3, gate151inter4, gate151inter5, gate151inter6, gate151inter7, gate151inter8, gate151inter9, gate151inter10, gate151inter11, gate151inter12, gate94inter0, gate94inter1, gate94inter2, gate94inter3, gate94inter4, gate94inter5, gate94inter6, gate94inter7, gate94inter8, gate94inter9, gate94inter10, gate94inter11, gate94inter12, gate14inter0, gate14inter1, gate14inter2, gate14inter3, gate14inter4, gate14inter5, gate14inter6, gate14inter7, gate14inter8, gate14inter9, gate14inter10, gate14inter11, gate14inter12, gate201inter0, gate201inter1, gate201inter2, gate201inter3, gate201inter4, gate201inter5, gate201inter6, gate201inter7, gate201inter8, gate201inter9, gate201inter10, gate201inter11, gate201inter12, gate503inter0, gate503inter1, gate503inter2, gate503inter3, gate503inter4, gate503inter5, gate503inter6, gate503inter7, gate503inter8, gate503inter9, gate503inter10, gate503inter11, gate503inter12, gate408inter0, gate408inter1, gate408inter2, gate408inter3, gate408inter4, gate408inter5, gate408inter6, gate408inter7, gate408inter8, gate408inter9, gate408inter10, gate408inter11, gate408inter12, gate256inter0, gate256inter1, gate256inter2, gate256inter3, gate256inter4, gate256inter5, gate256inter6, gate256inter7, gate256inter8, gate256inter9, gate256inter10, gate256inter11, gate256inter12, gate193inter0, gate193inter1, gate193inter2, gate193inter3, gate193inter4, gate193inter5, gate193inter6, gate193inter7, gate193inter8, gate193inter9, gate193inter10, gate193inter11, gate193inter12, gate133inter0, gate133inter1, gate133inter2, gate133inter3, gate133inter4, gate133inter5, gate133inter6, gate133inter7, gate133inter8, gate133inter9, gate133inter10, gate133inter11, gate133inter12, gate60inter0, gate60inter1, gate60inter2, gate60inter3, gate60inter4, gate60inter5, gate60inter6, gate60inter7, gate60inter8, gate60inter9, gate60inter10, gate60inter11, gate60inter12, gate85inter0, gate85inter1, gate85inter2, gate85inter3, gate85inter4, gate85inter5, gate85inter6, gate85inter7, gate85inter8, gate85inter9, gate85inter10, gate85inter11, gate85inter12, gate462inter0, gate462inter1, gate462inter2, gate462inter3, gate462inter4, gate462inter5, gate462inter6, gate462inter7, gate462inter8, gate462inter9, gate462inter10, gate462inter11, gate462inter12, gate89inter0, gate89inter1, gate89inter2, gate89inter3, gate89inter4, gate89inter5, gate89inter6, gate89inter7, gate89inter8, gate89inter9, gate89inter10, gate89inter11, gate89inter12, gate387inter0, gate387inter1, gate387inter2, gate387inter3, gate387inter4, gate387inter5, gate387inter6, gate387inter7, gate387inter8, gate387inter9, gate387inter10, gate387inter11, gate387inter12, gate233inter0, gate233inter1, gate233inter2, gate233inter3, gate233inter4, gate233inter5, gate233inter6, gate233inter7, gate233inter8, gate233inter9, gate233inter10, gate233inter11, gate233inter12, gate513inter0, gate513inter1, gate513inter2, gate513inter3, gate513inter4, gate513inter5, gate513inter6, gate513inter7, gate513inter8, gate513inter9, gate513inter10, gate513inter11, gate513inter12, gate426inter0, gate426inter1, gate426inter2, gate426inter3, gate426inter4, gate426inter5, gate426inter6, gate426inter7, gate426inter8, gate426inter9, gate426inter10, gate426inter11, gate426inter12, gate480inter0, gate480inter1, gate480inter2, gate480inter3, gate480inter4, gate480inter5, gate480inter6, gate480inter7, gate480inter8, gate480inter9, gate480inter10, gate480inter11, gate480inter12, gate115inter0, gate115inter1, gate115inter2, gate115inter3, gate115inter4, gate115inter5, gate115inter6, gate115inter7, gate115inter8, gate115inter9, gate115inter10, gate115inter11, gate115inter12, gate388inter0, gate388inter1, gate388inter2, gate388inter3, gate388inter4, gate388inter5, gate388inter6, gate388inter7, gate388inter8, gate388inter9, gate388inter10, gate388inter11, gate388inter12, gate76inter0, gate76inter1, gate76inter2, gate76inter3, gate76inter4, gate76inter5, gate76inter6, gate76inter7, gate76inter8, gate76inter9, gate76inter10, gate76inter11, gate76inter12, gate54inter0, gate54inter1, gate54inter2, gate54inter3, gate54inter4, gate54inter5, gate54inter6, gate54inter7, gate54inter8, gate54inter9, gate54inter10, gate54inter11, gate54inter12, gate149inter0, gate149inter1, gate149inter2, gate149inter3, gate149inter4, gate149inter5, gate149inter6, gate149inter7, gate149inter8, gate149inter9, gate149inter10, gate149inter11, gate149inter12, gate247inter0, gate247inter1, gate247inter2, gate247inter3, gate247inter4, gate247inter5, gate247inter6, gate247inter7, gate247inter8, gate247inter9, gate247inter10, gate247inter11, gate247inter12, gate292inter0, gate292inter1, gate292inter2, gate292inter3, gate292inter4, gate292inter5, gate292inter6, gate292inter7, gate292inter8, gate292inter9, gate292inter10, gate292inter11, gate292inter12, gate123inter0, gate123inter1, gate123inter2, gate123inter3, gate123inter4, gate123inter5, gate123inter6, gate123inter7, gate123inter8, gate123inter9, gate123inter10, gate123inter11, gate123inter12;



and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );

  xor2  gate995(.a(G2), .b(G1), .O(gate9inter0));
  nand2 gate996(.a(gate9inter0), .b(s_64), .O(gate9inter1));
  and2  gate997(.a(G2), .b(G1), .O(gate9inter2));
  inv1  gate998(.a(s_64), .O(gate9inter3));
  inv1  gate999(.a(s_65), .O(gate9inter4));
  nand2 gate1000(.a(gate9inter4), .b(gate9inter3), .O(gate9inter5));
  nor2  gate1001(.a(gate9inter5), .b(gate9inter2), .O(gate9inter6));
  inv1  gate1002(.a(G1), .O(gate9inter7));
  inv1  gate1003(.a(G2), .O(gate9inter8));
  nand2 gate1004(.a(gate9inter8), .b(gate9inter7), .O(gate9inter9));
  nand2 gate1005(.a(s_65), .b(gate9inter3), .O(gate9inter10));
  nor2  gate1006(.a(gate9inter10), .b(gate9inter9), .O(gate9inter11));
  nor2  gate1007(.a(gate9inter11), .b(gate9inter6), .O(gate9inter12));
  nand2 gate1008(.a(gate9inter12), .b(gate9inter1), .O(G266));

  xor2  gate1611(.a(G4), .b(G3), .O(gate10inter0));
  nand2 gate1612(.a(gate10inter0), .b(s_152), .O(gate10inter1));
  and2  gate1613(.a(G4), .b(G3), .O(gate10inter2));
  inv1  gate1614(.a(s_152), .O(gate10inter3));
  inv1  gate1615(.a(s_153), .O(gate10inter4));
  nand2 gate1616(.a(gate10inter4), .b(gate10inter3), .O(gate10inter5));
  nor2  gate1617(.a(gate10inter5), .b(gate10inter2), .O(gate10inter6));
  inv1  gate1618(.a(G3), .O(gate10inter7));
  inv1  gate1619(.a(G4), .O(gate10inter8));
  nand2 gate1620(.a(gate10inter8), .b(gate10inter7), .O(gate10inter9));
  nand2 gate1621(.a(s_153), .b(gate10inter3), .O(gate10inter10));
  nor2  gate1622(.a(gate10inter10), .b(gate10inter9), .O(gate10inter11));
  nor2  gate1623(.a(gate10inter11), .b(gate10inter6), .O(gate10inter12));
  nand2 gate1624(.a(gate10inter12), .b(gate10inter1), .O(G269));

  xor2  gate2311(.a(G6), .b(G5), .O(gate11inter0));
  nand2 gate2312(.a(gate11inter0), .b(s_252), .O(gate11inter1));
  and2  gate2313(.a(G6), .b(G5), .O(gate11inter2));
  inv1  gate2314(.a(s_252), .O(gate11inter3));
  inv1  gate2315(.a(s_253), .O(gate11inter4));
  nand2 gate2316(.a(gate11inter4), .b(gate11inter3), .O(gate11inter5));
  nor2  gate2317(.a(gate11inter5), .b(gate11inter2), .O(gate11inter6));
  inv1  gate2318(.a(G5), .O(gate11inter7));
  inv1  gate2319(.a(G6), .O(gate11inter8));
  nand2 gate2320(.a(gate11inter8), .b(gate11inter7), .O(gate11inter9));
  nand2 gate2321(.a(s_253), .b(gate11inter3), .O(gate11inter10));
  nor2  gate2322(.a(gate11inter10), .b(gate11inter9), .O(gate11inter11));
  nor2  gate2323(.a(gate11inter11), .b(gate11inter6), .O(gate11inter12));
  nand2 gate2324(.a(gate11inter12), .b(gate11inter1), .O(G272));
nand2 gate12( .a(G7), .b(G8), .O(G275) );
nand2 gate13( .a(G9), .b(G10), .O(G278) );

  xor2  gate2745(.a(G12), .b(G11), .O(gate14inter0));
  nand2 gate2746(.a(gate14inter0), .b(s_314), .O(gate14inter1));
  and2  gate2747(.a(G12), .b(G11), .O(gate14inter2));
  inv1  gate2748(.a(s_314), .O(gate14inter3));
  inv1  gate2749(.a(s_315), .O(gate14inter4));
  nand2 gate2750(.a(gate14inter4), .b(gate14inter3), .O(gate14inter5));
  nor2  gate2751(.a(gate14inter5), .b(gate14inter2), .O(gate14inter6));
  inv1  gate2752(.a(G11), .O(gate14inter7));
  inv1  gate2753(.a(G12), .O(gate14inter8));
  nand2 gate2754(.a(gate14inter8), .b(gate14inter7), .O(gate14inter9));
  nand2 gate2755(.a(s_315), .b(gate14inter3), .O(gate14inter10));
  nor2  gate2756(.a(gate14inter10), .b(gate14inter9), .O(gate14inter11));
  nor2  gate2757(.a(gate14inter11), .b(gate14inter6), .O(gate14inter12));
  nand2 gate2758(.a(gate14inter12), .b(gate14inter1), .O(G281));

  xor2  gate1121(.a(G14), .b(G13), .O(gate15inter0));
  nand2 gate1122(.a(gate15inter0), .b(s_82), .O(gate15inter1));
  and2  gate1123(.a(G14), .b(G13), .O(gate15inter2));
  inv1  gate1124(.a(s_82), .O(gate15inter3));
  inv1  gate1125(.a(s_83), .O(gate15inter4));
  nand2 gate1126(.a(gate15inter4), .b(gate15inter3), .O(gate15inter5));
  nor2  gate1127(.a(gate15inter5), .b(gate15inter2), .O(gate15inter6));
  inv1  gate1128(.a(G13), .O(gate15inter7));
  inv1  gate1129(.a(G14), .O(gate15inter8));
  nand2 gate1130(.a(gate15inter8), .b(gate15inter7), .O(gate15inter9));
  nand2 gate1131(.a(s_83), .b(gate15inter3), .O(gate15inter10));
  nor2  gate1132(.a(gate15inter10), .b(gate15inter9), .O(gate15inter11));
  nor2  gate1133(.a(gate15inter11), .b(gate15inter6), .O(gate15inter12));
  nand2 gate1134(.a(gate15inter12), .b(gate15inter1), .O(G284));

  xor2  gate2143(.a(G16), .b(G15), .O(gate16inter0));
  nand2 gate2144(.a(gate16inter0), .b(s_228), .O(gate16inter1));
  and2  gate2145(.a(G16), .b(G15), .O(gate16inter2));
  inv1  gate2146(.a(s_228), .O(gate16inter3));
  inv1  gate2147(.a(s_229), .O(gate16inter4));
  nand2 gate2148(.a(gate16inter4), .b(gate16inter3), .O(gate16inter5));
  nor2  gate2149(.a(gate16inter5), .b(gate16inter2), .O(gate16inter6));
  inv1  gate2150(.a(G15), .O(gate16inter7));
  inv1  gate2151(.a(G16), .O(gate16inter8));
  nand2 gate2152(.a(gate16inter8), .b(gate16inter7), .O(gate16inter9));
  nand2 gate2153(.a(s_229), .b(gate16inter3), .O(gate16inter10));
  nor2  gate2154(.a(gate16inter10), .b(gate16inter9), .O(gate16inter11));
  nor2  gate2155(.a(gate16inter11), .b(gate16inter6), .O(gate16inter12));
  nand2 gate2156(.a(gate16inter12), .b(gate16inter1), .O(G287));
nand2 gate17( .a(G17), .b(G18), .O(G290) );

  xor2  gate1247(.a(G20), .b(G19), .O(gate18inter0));
  nand2 gate1248(.a(gate18inter0), .b(s_100), .O(gate18inter1));
  and2  gate1249(.a(G20), .b(G19), .O(gate18inter2));
  inv1  gate1250(.a(s_100), .O(gate18inter3));
  inv1  gate1251(.a(s_101), .O(gate18inter4));
  nand2 gate1252(.a(gate18inter4), .b(gate18inter3), .O(gate18inter5));
  nor2  gate1253(.a(gate18inter5), .b(gate18inter2), .O(gate18inter6));
  inv1  gate1254(.a(G19), .O(gate18inter7));
  inv1  gate1255(.a(G20), .O(gate18inter8));
  nand2 gate1256(.a(gate18inter8), .b(gate18inter7), .O(gate18inter9));
  nand2 gate1257(.a(s_101), .b(gate18inter3), .O(gate18inter10));
  nor2  gate1258(.a(gate18inter10), .b(gate18inter9), .O(gate18inter11));
  nor2  gate1259(.a(gate18inter11), .b(gate18inter6), .O(gate18inter12));
  nand2 gate1260(.a(gate18inter12), .b(gate18inter1), .O(G293));
nand2 gate19( .a(G21), .b(G22), .O(G296) );

  xor2  gate1541(.a(G24), .b(G23), .O(gate20inter0));
  nand2 gate1542(.a(gate20inter0), .b(s_142), .O(gate20inter1));
  and2  gate1543(.a(G24), .b(G23), .O(gate20inter2));
  inv1  gate1544(.a(s_142), .O(gate20inter3));
  inv1  gate1545(.a(s_143), .O(gate20inter4));
  nand2 gate1546(.a(gate20inter4), .b(gate20inter3), .O(gate20inter5));
  nor2  gate1547(.a(gate20inter5), .b(gate20inter2), .O(gate20inter6));
  inv1  gate1548(.a(G23), .O(gate20inter7));
  inv1  gate1549(.a(G24), .O(gate20inter8));
  nand2 gate1550(.a(gate20inter8), .b(gate20inter7), .O(gate20inter9));
  nand2 gate1551(.a(s_143), .b(gate20inter3), .O(gate20inter10));
  nor2  gate1552(.a(gate20inter10), .b(gate20inter9), .O(gate20inter11));
  nor2  gate1553(.a(gate20inter11), .b(gate20inter6), .O(gate20inter12));
  nand2 gate1554(.a(gate20inter12), .b(gate20inter1), .O(G299));

  xor2  gate1303(.a(G26), .b(G25), .O(gate21inter0));
  nand2 gate1304(.a(gate21inter0), .b(s_108), .O(gate21inter1));
  and2  gate1305(.a(G26), .b(G25), .O(gate21inter2));
  inv1  gate1306(.a(s_108), .O(gate21inter3));
  inv1  gate1307(.a(s_109), .O(gate21inter4));
  nand2 gate1308(.a(gate21inter4), .b(gate21inter3), .O(gate21inter5));
  nor2  gate1309(.a(gate21inter5), .b(gate21inter2), .O(gate21inter6));
  inv1  gate1310(.a(G25), .O(gate21inter7));
  inv1  gate1311(.a(G26), .O(gate21inter8));
  nand2 gate1312(.a(gate21inter8), .b(gate21inter7), .O(gate21inter9));
  nand2 gate1313(.a(s_109), .b(gate21inter3), .O(gate21inter10));
  nor2  gate1314(.a(gate21inter10), .b(gate21inter9), .O(gate21inter11));
  nor2  gate1315(.a(gate21inter11), .b(gate21inter6), .O(gate21inter12));
  nand2 gate1316(.a(gate21inter12), .b(gate21inter1), .O(G302));

  xor2  gate1793(.a(G28), .b(G27), .O(gate22inter0));
  nand2 gate1794(.a(gate22inter0), .b(s_178), .O(gate22inter1));
  and2  gate1795(.a(G28), .b(G27), .O(gate22inter2));
  inv1  gate1796(.a(s_178), .O(gate22inter3));
  inv1  gate1797(.a(s_179), .O(gate22inter4));
  nand2 gate1798(.a(gate22inter4), .b(gate22inter3), .O(gate22inter5));
  nor2  gate1799(.a(gate22inter5), .b(gate22inter2), .O(gate22inter6));
  inv1  gate1800(.a(G27), .O(gate22inter7));
  inv1  gate1801(.a(G28), .O(gate22inter8));
  nand2 gate1802(.a(gate22inter8), .b(gate22inter7), .O(gate22inter9));
  nand2 gate1803(.a(s_179), .b(gate22inter3), .O(gate22inter10));
  nor2  gate1804(.a(gate22inter10), .b(gate22inter9), .O(gate22inter11));
  nor2  gate1805(.a(gate22inter11), .b(gate22inter6), .O(gate22inter12));
  nand2 gate1806(.a(gate22inter12), .b(gate22inter1), .O(G305));

  xor2  gate2045(.a(G30), .b(G29), .O(gate23inter0));
  nand2 gate2046(.a(gate23inter0), .b(s_214), .O(gate23inter1));
  and2  gate2047(.a(G30), .b(G29), .O(gate23inter2));
  inv1  gate2048(.a(s_214), .O(gate23inter3));
  inv1  gate2049(.a(s_215), .O(gate23inter4));
  nand2 gate2050(.a(gate23inter4), .b(gate23inter3), .O(gate23inter5));
  nor2  gate2051(.a(gate23inter5), .b(gate23inter2), .O(gate23inter6));
  inv1  gate2052(.a(G29), .O(gate23inter7));
  inv1  gate2053(.a(G30), .O(gate23inter8));
  nand2 gate2054(.a(gate23inter8), .b(gate23inter7), .O(gate23inter9));
  nand2 gate2055(.a(s_215), .b(gate23inter3), .O(gate23inter10));
  nor2  gate2056(.a(gate23inter10), .b(gate23inter9), .O(gate23inter11));
  nor2  gate2057(.a(gate23inter11), .b(gate23inter6), .O(gate23inter12));
  nand2 gate2058(.a(gate23inter12), .b(gate23inter1), .O(G308));

  xor2  gate981(.a(G32), .b(G31), .O(gate24inter0));
  nand2 gate982(.a(gate24inter0), .b(s_62), .O(gate24inter1));
  and2  gate983(.a(G32), .b(G31), .O(gate24inter2));
  inv1  gate984(.a(s_62), .O(gate24inter3));
  inv1  gate985(.a(s_63), .O(gate24inter4));
  nand2 gate986(.a(gate24inter4), .b(gate24inter3), .O(gate24inter5));
  nor2  gate987(.a(gate24inter5), .b(gate24inter2), .O(gate24inter6));
  inv1  gate988(.a(G31), .O(gate24inter7));
  inv1  gate989(.a(G32), .O(gate24inter8));
  nand2 gate990(.a(gate24inter8), .b(gate24inter7), .O(gate24inter9));
  nand2 gate991(.a(s_63), .b(gate24inter3), .O(gate24inter10));
  nor2  gate992(.a(gate24inter10), .b(gate24inter9), .O(gate24inter11));
  nor2  gate993(.a(gate24inter11), .b(gate24inter6), .O(gate24inter12));
  nand2 gate994(.a(gate24inter12), .b(gate24inter1), .O(G311));
nand2 gate25( .a(G1), .b(G5), .O(G314) );
nand2 gate26( .a(G9), .b(G13), .O(G317) );

  xor2  gate1443(.a(G6), .b(G2), .O(gate27inter0));
  nand2 gate1444(.a(gate27inter0), .b(s_128), .O(gate27inter1));
  and2  gate1445(.a(G6), .b(G2), .O(gate27inter2));
  inv1  gate1446(.a(s_128), .O(gate27inter3));
  inv1  gate1447(.a(s_129), .O(gate27inter4));
  nand2 gate1448(.a(gate27inter4), .b(gate27inter3), .O(gate27inter5));
  nor2  gate1449(.a(gate27inter5), .b(gate27inter2), .O(gate27inter6));
  inv1  gate1450(.a(G2), .O(gate27inter7));
  inv1  gate1451(.a(G6), .O(gate27inter8));
  nand2 gate1452(.a(gate27inter8), .b(gate27inter7), .O(gate27inter9));
  nand2 gate1453(.a(s_129), .b(gate27inter3), .O(gate27inter10));
  nor2  gate1454(.a(gate27inter10), .b(gate27inter9), .O(gate27inter11));
  nor2  gate1455(.a(gate27inter11), .b(gate27inter6), .O(gate27inter12));
  nand2 gate1456(.a(gate27inter12), .b(gate27inter1), .O(G320));

  xor2  gate1975(.a(G14), .b(G10), .O(gate28inter0));
  nand2 gate1976(.a(gate28inter0), .b(s_204), .O(gate28inter1));
  and2  gate1977(.a(G14), .b(G10), .O(gate28inter2));
  inv1  gate1978(.a(s_204), .O(gate28inter3));
  inv1  gate1979(.a(s_205), .O(gate28inter4));
  nand2 gate1980(.a(gate28inter4), .b(gate28inter3), .O(gate28inter5));
  nor2  gate1981(.a(gate28inter5), .b(gate28inter2), .O(gate28inter6));
  inv1  gate1982(.a(G10), .O(gate28inter7));
  inv1  gate1983(.a(G14), .O(gate28inter8));
  nand2 gate1984(.a(gate28inter8), .b(gate28inter7), .O(gate28inter9));
  nand2 gate1985(.a(s_205), .b(gate28inter3), .O(gate28inter10));
  nor2  gate1986(.a(gate28inter10), .b(gate28inter9), .O(gate28inter11));
  nor2  gate1987(.a(gate28inter11), .b(gate28inter6), .O(gate28inter12));
  nand2 gate1988(.a(gate28inter12), .b(gate28inter1), .O(G323));
nand2 gate29( .a(G3), .b(G7), .O(G326) );
nand2 gate30( .a(G11), .b(G15), .O(G329) );
nand2 gate31( .a(G4), .b(G8), .O(G332) );
nand2 gate32( .a(G12), .b(G16), .O(G335) );
nand2 gate33( .a(G17), .b(G21), .O(G338) );
nand2 gate34( .a(G25), .b(G29), .O(G341) );

  xor2  gate1639(.a(G22), .b(G18), .O(gate35inter0));
  nand2 gate1640(.a(gate35inter0), .b(s_156), .O(gate35inter1));
  and2  gate1641(.a(G22), .b(G18), .O(gate35inter2));
  inv1  gate1642(.a(s_156), .O(gate35inter3));
  inv1  gate1643(.a(s_157), .O(gate35inter4));
  nand2 gate1644(.a(gate35inter4), .b(gate35inter3), .O(gate35inter5));
  nor2  gate1645(.a(gate35inter5), .b(gate35inter2), .O(gate35inter6));
  inv1  gate1646(.a(G18), .O(gate35inter7));
  inv1  gate1647(.a(G22), .O(gate35inter8));
  nand2 gate1648(.a(gate35inter8), .b(gate35inter7), .O(gate35inter9));
  nand2 gate1649(.a(s_157), .b(gate35inter3), .O(gate35inter10));
  nor2  gate1650(.a(gate35inter10), .b(gate35inter9), .O(gate35inter11));
  nor2  gate1651(.a(gate35inter11), .b(gate35inter6), .O(gate35inter12));
  nand2 gate1652(.a(gate35inter12), .b(gate35inter1), .O(G344));
nand2 gate36( .a(G26), .b(G30), .O(G347) );
nand2 gate37( .a(G19), .b(G23), .O(G350) );
nand2 gate38( .a(G27), .b(G31), .O(G353) );

  xor2  gate743(.a(G24), .b(G20), .O(gate39inter0));
  nand2 gate744(.a(gate39inter0), .b(s_28), .O(gate39inter1));
  and2  gate745(.a(G24), .b(G20), .O(gate39inter2));
  inv1  gate746(.a(s_28), .O(gate39inter3));
  inv1  gate747(.a(s_29), .O(gate39inter4));
  nand2 gate748(.a(gate39inter4), .b(gate39inter3), .O(gate39inter5));
  nor2  gate749(.a(gate39inter5), .b(gate39inter2), .O(gate39inter6));
  inv1  gate750(.a(G20), .O(gate39inter7));
  inv1  gate751(.a(G24), .O(gate39inter8));
  nand2 gate752(.a(gate39inter8), .b(gate39inter7), .O(gate39inter9));
  nand2 gate753(.a(s_29), .b(gate39inter3), .O(gate39inter10));
  nor2  gate754(.a(gate39inter10), .b(gate39inter9), .O(gate39inter11));
  nor2  gate755(.a(gate39inter11), .b(gate39inter6), .O(gate39inter12));
  nand2 gate756(.a(gate39inter12), .b(gate39inter1), .O(G356));

  xor2  gate1555(.a(G32), .b(G28), .O(gate40inter0));
  nand2 gate1556(.a(gate40inter0), .b(s_144), .O(gate40inter1));
  and2  gate1557(.a(G32), .b(G28), .O(gate40inter2));
  inv1  gate1558(.a(s_144), .O(gate40inter3));
  inv1  gate1559(.a(s_145), .O(gate40inter4));
  nand2 gate1560(.a(gate40inter4), .b(gate40inter3), .O(gate40inter5));
  nor2  gate1561(.a(gate40inter5), .b(gate40inter2), .O(gate40inter6));
  inv1  gate1562(.a(G28), .O(gate40inter7));
  inv1  gate1563(.a(G32), .O(gate40inter8));
  nand2 gate1564(.a(gate40inter8), .b(gate40inter7), .O(gate40inter9));
  nand2 gate1565(.a(s_145), .b(gate40inter3), .O(gate40inter10));
  nor2  gate1566(.a(gate40inter10), .b(gate40inter9), .O(gate40inter11));
  nor2  gate1567(.a(gate40inter11), .b(gate40inter6), .O(gate40inter12));
  nand2 gate1568(.a(gate40inter12), .b(gate40inter1), .O(G359));

  xor2  gate2283(.a(G266), .b(G1), .O(gate41inter0));
  nand2 gate2284(.a(gate41inter0), .b(s_248), .O(gate41inter1));
  and2  gate2285(.a(G266), .b(G1), .O(gate41inter2));
  inv1  gate2286(.a(s_248), .O(gate41inter3));
  inv1  gate2287(.a(s_249), .O(gate41inter4));
  nand2 gate2288(.a(gate41inter4), .b(gate41inter3), .O(gate41inter5));
  nor2  gate2289(.a(gate41inter5), .b(gate41inter2), .O(gate41inter6));
  inv1  gate2290(.a(G1), .O(gate41inter7));
  inv1  gate2291(.a(G266), .O(gate41inter8));
  nand2 gate2292(.a(gate41inter8), .b(gate41inter7), .O(gate41inter9));
  nand2 gate2293(.a(s_249), .b(gate41inter3), .O(gate41inter10));
  nor2  gate2294(.a(gate41inter10), .b(gate41inter9), .O(gate41inter11));
  nor2  gate2295(.a(gate41inter11), .b(gate41inter6), .O(gate41inter12));
  nand2 gate2296(.a(gate41inter12), .b(gate41inter1), .O(G362));

  xor2  gate1289(.a(G266), .b(G2), .O(gate42inter0));
  nand2 gate1290(.a(gate42inter0), .b(s_106), .O(gate42inter1));
  and2  gate1291(.a(G266), .b(G2), .O(gate42inter2));
  inv1  gate1292(.a(s_106), .O(gate42inter3));
  inv1  gate1293(.a(s_107), .O(gate42inter4));
  nand2 gate1294(.a(gate42inter4), .b(gate42inter3), .O(gate42inter5));
  nor2  gate1295(.a(gate42inter5), .b(gate42inter2), .O(gate42inter6));
  inv1  gate1296(.a(G2), .O(gate42inter7));
  inv1  gate1297(.a(G266), .O(gate42inter8));
  nand2 gate1298(.a(gate42inter8), .b(gate42inter7), .O(gate42inter9));
  nand2 gate1299(.a(s_107), .b(gate42inter3), .O(gate42inter10));
  nor2  gate1300(.a(gate42inter10), .b(gate42inter9), .O(gate42inter11));
  nor2  gate1301(.a(gate42inter11), .b(gate42inter6), .O(gate42inter12));
  nand2 gate1302(.a(gate42inter12), .b(gate42inter1), .O(G363));

  xor2  gate1835(.a(G269), .b(G3), .O(gate43inter0));
  nand2 gate1836(.a(gate43inter0), .b(s_184), .O(gate43inter1));
  and2  gate1837(.a(G269), .b(G3), .O(gate43inter2));
  inv1  gate1838(.a(s_184), .O(gate43inter3));
  inv1  gate1839(.a(s_185), .O(gate43inter4));
  nand2 gate1840(.a(gate43inter4), .b(gate43inter3), .O(gate43inter5));
  nor2  gate1841(.a(gate43inter5), .b(gate43inter2), .O(gate43inter6));
  inv1  gate1842(.a(G3), .O(gate43inter7));
  inv1  gate1843(.a(G269), .O(gate43inter8));
  nand2 gate1844(.a(gate43inter8), .b(gate43inter7), .O(gate43inter9));
  nand2 gate1845(.a(s_185), .b(gate43inter3), .O(gate43inter10));
  nor2  gate1846(.a(gate43inter10), .b(gate43inter9), .O(gate43inter11));
  nor2  gate1847(.a(gate43inter11), .b(gate43inter6), .O(gate43inter12));
  nand2 gate1848(.a(gate43inter12), .b(gate43inter1), .O(G364));
nand2 gate44( .a(G4), .b(G269), .O(G365) );
nand2 gate45( .a(G5), .b(G272), .O(G366) );

  xor2  gate1513(.a(G272), .b(G6), .O(gate46inter0));
  nand2 gate1514(.a(gate46inter0), .b(s_138), .O(gate46inter1));
  and2  gate1515(.a(G272), .b(G6), .O(gate46inter2));
  inv1  gate1516(.a(s_138), .O(gate46inter3));
  inv1  gate1517(.a(s_139), .O(gate46inter4));
  nand2 gate1518(.a(gate46inter4), .b(gate46inter3), .O(gate46inter5));
  nor2  gate1519(.a(gate46inter5), .b(gate46inter2), .O(gate46inter6));
  inv1  gate1520(.a(G6), .O(gate46inter7));
  inv1  gate1521(.a(G272), .O(gate46inter8));
  nand2 gate1522(.a(gate46inter8), .b(gate46inter7), .O(gate46inter9));
  nand2 gate1523(.a(s_139), .b(gate46inter3), .O(gate46inter10));
  nor2  gate1524(.a(gate46inter10), .b(gate46inter9), .O(gate46inter11));
  nor2  gate1525(.a(gate46inter11), .b(gate46inter6), .O(gate46inter12));
  nand2 gate1526(.a(gate46inter12), .b(gate46inter1), .O(G367));
nand2 gate47( .a(G7), .b(G275), .O(G368) );
nand2 gate48( .a(G8), .b(G275), .O(G369) );
nand2 gate49( .a(G9), .b(G278), .O(G370) );
nand2 gate50( .a(G10), .b(G278), .O(G371) );
nand2 gate51( .a(G11), .b(G281), .O(G372) );
nand2 gate52( .a(G12), .b(G281), .O(G373) );
nand2 gate53( .a(G13), .b(G284), .O(G374) );

  xor2  gate3011(.a(G284), .b(G14), .O(gate54inter0));
  nand2 gate3012(.a(gate54inter0), .b(s_352), .O(gate54inter1));
  and2  gate3013(.a(G284), .b(G14), .O(gate54inter2));
  inv1  gate3014(.a(s_352), .O(gate54inter3));
  inv1  gate3015(.a(s_353), .O(gate54inter4));
  nand2 gate3016(.a(gate54inter4), .b(gate54inter3), .O(gate54inter5));
  nor2  gate3017(.a(gate54inter5), .b(gate54inter2), .O(gate54inter6));
  inv1  gate3018(.a(G14), .O(gate54inter7));
  inv1  gate3019(.a(G284), .O(gate54inter8));
  nand2 gate3020(.a(gate54inter8), .b(gate54inter7), .O(gate54inter9));
  nand2 gate3021(.a(s_353), .b(gate54inter3), .O(gate54inter10));
  nor2  gate3022(.a(gate54inter10), .b(gate54inter9), .O(gate54inter11));
  nor2  gate3023(.a(gate54inter11), .b(gate54inter6), .O(gate54inter12));
  nand2 gate3024(.a(gate54inter12), .b(gate54inter1), .O(G375));
nand2 gate55( .a(G15), .b(G287), .O(G376) );

  xor2  gate701(.a(G287), .b(G16), .O(gate56inter0));
  nand2 gate702(.a(gate56inter0), .b(s_22), .O(gate56inter1));
  and2  gate703(.a(G287), .b(G16), .O(gate56inter2));
  inv1  gate704(.a(s_22), .O(gate56inter3));
  inv1  gate705(.a(s_23), .O(gate56inter4));
  nand2 gate706(.a(gate56inter4), .b(gate56inter3), .O(gate56inter5));
  nor2  gate707(.a(gate56inter5), .b(gate56inter2), .O(gate56inter6));
  inv1  gate708(.a(G16), .O(gate56inter7));
  inv1  gate709(.a(G287), .O(gate56inter8));
  nand2 gate710(.a(gate56inter8), .b(gate56inter7), .O(gate56inter9));
  nand2 gate711(.a(s_23), .b(gate56inter3), .O(gate56inter10));
  nor2  gate712(.a(gate56inter10), .b(gate56inter9), .O(gate56inter11));
  nor2  gate713(.a(gate56inter11), .b(gate56inter6), .O(gate56inter12));
  nand2 gate714(.a(gate56inter12), .b(gate56inter1), .O(G377));
nand2 gate57( .a(G17), .b(G290), .O(G378) );

  xor2  gate2591(.a(G290), .b(G18), .O(gate58inter0));
  nand2 gate2592(.a(gate58inter0), .b(s_292), .O(gate58inter1));
  and2  gate2593(.a(G290), .b(G18), .O(gate58inter2));
  inv1  gate2594(.a(s_292), .O(gate58inter3));
  inv1  gate2595(.a(s_293), .O(gate58inter4));
  nand2 gate2596(.a(gate58inter4), .b(gate58inter3), .O(gate58inter5));
  nor2  gate2597(.a(gate58inter5), .b(gate58inter2), .O(gate58inter6));
  inv1  gate2598(.a(G18), .O(gate58inter7));
  inv1  gate2599(.a(G290), .O(gate58inter8));
  nand2 gate2600(.a(gate58inter8), .b(gate58inter7), .O(gate58inter9));
  nand2 gate2601(.a(s_293), .b(gate58inter3), .O(gate58inter10));
  nor2  gate2602(.a(gate58inter10), .b(gate58inter9), .O(gate58inter11));
  nor2  gate2603(.a(gate58inter11), .b(gate58inter6), .O(gate58inter12));
  nand2 gate2604(.a(gate58inter12), .b(gate58inter1), .O(G379));
nand2 gate59( .a(G19), .b(G293), .O(G380) );

  xor2  gate2843(.a(G293), .b(G20), .O(gate60inter0));
  nand2 gate2844(.a(gate60inter0), .b(s_328), .O(gate60inter1));
  and2  gate2845(.a(G293), .b(G20), .O(gate60inter2));
  inv1  gate2846(.a(s_328), .O(gate60inter3));
  inv1  gate2847(.a(s_329), .O(gate60inter4));
  nand2 gate2848(.a(gate60inter4), .b(gate60inter3), .O(gate60inter5));
  nor2  gate2849(.a(gate60inter5), .b(gate60inter2), .O(gate60inter6));
  inv1  gate2850(.a(G20), .O(gate60inter7));
  inv1  gate2851(.a(G293), .O(gate60inter8));
  nand2 gate2852(.a(gate60inter8), .b(gate60inter7), .O(gate60inter9));
  nand2 gate2853(.a(s_329), .b(gate60inter3), .O(gate60inter10));
  nor2  gate2854(.a(gate60inter10), .b(gate60inter9), .O(gate60inter11));
  nor2  gate2855(.a(gate60inter11), .b(gate60inter6), .O(gate60inter12));
  nand2 gate2856(.a(gate60inter12), .b(gate60inter1), .O(G381));

  xor2  gate1807(.a(G296), .b(G21), .O(gate61inter0));
  nand2 gate1808(.a(gate61inter0), .b(s_180), .O(gate61inter1));
  and2  gate1809(.a(G296), .b(G21), .O(gate61inter2));
  inv1  gate1810(.a(s_180), .O(gate61inter3));
  inv1  gate1811(.a(s_181), .O(gate61inter4));
  nand2 gate1812(.a(gate61inter4), .b(gate61inter3), .O(gate61inter5));
  nor2  gate1813(.a(gate61inter5), .b(gate61inter2), .O(gate61inter6));
  inv1  gate1814(.a(G21), .O(gate61inter7));
  inv1  gate1815(.a(G296), .O(gate61inter8));
  nand2 gate1816(.a(gate61inter8), .b(gate61inter7), .O(gate61inter9));
  nand2 gate1817(.a(s_181), .b(gate61inter3), .O(gate61inter10));
  nor2  gate1818(.a(gate61inter10), .b(gate61inter9), .O(gate61inter11));
  nor2  gate1819(.a(gate61inter11), .b(gate61inter6), .O(gate61inter12));
  nand2 gate1820(.a(gate61inter12), .b(gate61inter1), .O(G382));
nand2 gate62( .a(G22), .b(G296), .O(G383) );
nand2 gate63( .a(G23), .b(G299), .O(G384) );

  xor2  gate2381(.a(G299), .b(G24), .O(gate64inter0));
  nand2 gate2382(.a(gate64inter0), .b(s_262), .O(gate64inter1));
  and2  gate2383(.a(G299), .b(G24), .O(gate64inter2));
  inv1  gate2384(.a(s_262), .O(gate64inter3));
  inv1  gate2385(.a(s_263), .O(gate64inter4));
  nand2 gate2386(.a(gate64inter4), .b(gate64inter3), .O(gate64inter5));
  nor2  gate2387(.a(gate64inter5), .b(gate64inter2), .O(gate64inter6));
  inv1  gate2388(.a(G24), .O(gate64inter7));
  inv1  gate2389(.a(G299), .O(gate64inter8));
  nand2 gate2390(.a(gate64inter8), .b(gate64inter7), .O(gate64inter9));
  nand2 gate2391(.a(s_263), .b(gate64inter3), .O(gate64inter10));
  nor2  gate2392(.a(gate64inter10), .b(gate64inter9), .O(gate64inter11));
  nor2  gate2393(.a(gate64inter11), .b(gate64inter6), .O(gate64inter12));
  nand2 gate2394(.a(gate64inter12), .b(gate64inter1), .O(G385));
nand2 gate65( .a(G25), .b(G302), .O(G386) );
nand2 gate66( .a(G26), .b(G302), .O(G387) );

  xor2  gate1023(.a(G305), .b(G27), .O(gate67inter0));
  nand2 gate1024(.a(gate67inter0), .b(s_68), .O(gate67inter1));
  and2  gate1025(.a(G305), .b(G27), .O(gate67inter2));
  inv1  gate1026(.a(s_68), .O(gate67inter3));
  inv1  gate1027(.a(s_69), .O(gate67inter4));
  nand2 gate1028(.a(gate67inter4), .b(gate67inter3), .O(gate67inter5));
  nor2  gate1029(.a(gate67inter5), .b(gate67inter2), .O(gate67inter6));
  inv1  gate1030(.a(G27), .O(gate67inter7));
  inv1  gate1031(.a(G305), .O(gate67inter8));
  nand2 gate1032(.a(gate67inter8), .b(gate67inter7), .O(gate67inter9));
  nand2 gate1033(.a(s_69), .b(gate67inter3), .O(gate67inter10));
  nor2  gate1034(.a(gate67inter10), .b(gate67inter9), .O(gate67inter11));
  nor2  gate1035(.a(gate67inter11), .b(gate67inter6), .O(gate67inter12));
  nand2 gate1036(.a(gate67inter12), .b(gate67inter1), .O(G388));
nand2 gate68( .a(G28), .b(G305), .O(G389) );

  xor2  gate1401(.a(G308), .b(G29), .O(gate69inter0));
  nand2 gate1402(.a(gate69inter0), .b(s_122), .O(gate69inter1));
  and2  gate1403(.a(G308), .b(G29), .O(gate69inter2));
  inv1  gate1404(.a(s_122), .O(gate69inter3));
  inv1  gate1405(.a(s_123), .O(gate69inter4));
  nand2 gate1406(.a(gate69inter4), .b(gate69inter3), .O(gate69inter5));
  nor2  gate1407(.a(gate69inter5), .b(gate69inter2), .O(gate69inter6));
  inv1  gate1408(.a(G29), .O(gate69inter7));
  inv1  gate1409(.a(G308), .O(gate69inter8));
  nand2 gate1410(.a(gate69inter8), .b(gate69inter7), .O(gate69inter9));
  nand2 gate1411(.a(s_123), .b(gate69inter3), .O(gate69inter10));
  nor2  gate1412(.a(gate69inter10), .b(gate69inter9), .O(gate69inter11));
  nor2  gate1413(.a(gate69inter11), .b(gate69inter6), .O(gate69inter12));
  nand2 gate1414(.a(gate69inter12), .b(gate69inter1), .O(G390));

  xor2  gate939(.a(G308), .b(G30), .O(gate70inter0));
  nand2 gate940(.a(gate70inter0), .b(s_56), .O(gate70inter1));
  and2  gate941(.a(G308), .b(G30), .O(gate70inter2));
  inv1  gate942(.a(s_56), .O(gate70inter3));
  inv1  gate943(.a(s_57), .O(gate70inter4));
  nand2 gate944(.a(gate70inter4), .b(gate70inter3), .O(gate70inter5));
  nor2  gate945(.a(gate70inter5), .b(gate70inter2), .O(gate70inter6));
  inv1  gate946(.a(G30), .O(gate70inter7));
  inv1  gate947(.a(G308), .O(gate70inter8));
  nand2 gate948(.a(gate70inter8), .b(gate70inter7), .O(gate70inter9));
  nand2 gate949(.a(s_57), .b(gate70inter3), .O(gate70inter10));
  nor2  gate950(.a(gate70inter10), .b(gate70inter9), .O(gate70inter11));
  nor2  gate951(.a(gate70inter11), .b(gate70inter6), .O(gate70inter12));
  nand2 gate952(.a(gate70inter12), .b(gate70inter1), .O(G391));
nand2 gate71( .a(G31), .b(G311), .O(G392) );
nand2 gate72( .a(G32), .b(G311), .O(G393) );

  xor2  gate2073(.a(G314), .b(G1), .O(gate73inter0));
  nand2 gate2074(.a(gate73inter0), .b(s_218), .O(gate73inter1));
  and2  gate2075(.a(G314), .b(G1), .O(gate73inter2));
  inv1  gate2076(.a(s_218), .O(gate73inter3));
  inv1  gate2077(.a(s_219), .O(gate73inter4));
  nand2 gate2078(.a(gate73inter4), .b(gate73inter3), .O(gate73inter5));
  nor2  gate2079(.a(gate73inter5), .b(gate73inter2), .O(gate73inter6));
  inv1  gate2080(.a(G1), .O(gate73inter7));
  inv1  gate2081(.a(G314), .O(gate73inter8));
  nand2 gate2082(.a(gate73inter8), .b(gate73inter7), .O(gate73inter9));
  nand2 gate2083(.a(s_219), .b(gate73inter3), .O(gate73inter10));
  nor2  gate2084(.a(gate73inter10), .b(gate73inter9), .O(gate73inter11));
  nor2  gate2085(.a(gate73inter11), .b(gate73inter6), .O(gate73inter12));
  nand2 gate2086(.a(gate73inter12), .b(gate73inter1), .O(G394));

  xor2  gate2269(.a(G314), .b(G5), .O(gate74inter0));
  nand2 gate2270(.a(gate74inter0), .b(s_246), .O(gate74inter1));
  and2  gate2271(.a(G314), .b(G5), .O(gate74inter2));
  inv1  gate2272(.a(s_246), .O(gate74inter3));
  inv1  gate2273(.a(s_247), .O(gate74inter4));
  nand2 gate2274(.a(gate74inter4), .b(gate74inter3), .O(gate74inter5));
  nor2  gate2275(.a(gate74inter5), .b(gate74inter2), .O(gate74inter6));
  inv1  gate2276(.a(G5), .O(gate74inter7));
  inv1  gate2277(.a(G314), .O(gate74inter8));
  nand2 gate2278(.a(gate74inter8), .b(gate74inter7), .O(gate74inter9));
  nand2 gate2279(.a(s_247), .b(gate74inter3), .O(gate74inter10));
  nor2  gate2280(.a(gate74inter10), .b(gate74inter9), .O(gate74inter11));
  nor2  gate2281(.a(gate74inter11), .b(gate74inter6), .O(gate74inter12));
  nand2 gate2282(.a(gate74inter12), .b(gate74inter1), .O(G395));

  xor2  gate631(.a(G317), .b(G9), .O(gate75inter0));
  nand2 gate632(.a(gate75inter0), .b(s_12), .O(gate75inter1));
  and2  gate633(.a(G317), .b(G9), .O(gate75inter2));
  inv1  gate634(.a(s_12), .O(gate75inter3));
  inv1  gate635(.a(s_13), .O(gate75inter4));
  nand2 gate636(.a(gate75inter4), .b(gate75inter3), .O(gate75inter5));
  nor2  gate637(.a(gate75inter5), .b(gate75inter2), .O(gate75inter6));
  inv1  gate638(.a(G9), .O(gate75inter7));
  inv1  gate639(.a(G317), .O(gate75inter8));
  nand2 gate640(.a(gate75inter8), .b(gate75inter7), .O(gate75inter9));
  nand2 gate641(.a(s_13), .b(gate75inter3), .O(gate75inter10));
  nor2  gate642(.a(gate75inter10), .b(gate75inter9), .O(gate75inter11));
  nor2  gate643(.a(gate75inter11), .b(gate75inter6), .O(gate75inter12));
  nand2 gate644(.a(gate75inter12), .b(gate75inter1), .O(G396));

  xor2  gate2997(.a(G317), .b(G13), .O(gate76inter0));
  nand2 gate2998(.a(gate76inter0), .b(s_350), .O(gate76inter1));
  and2  gate2999(.a(G317), .b(G13), .O(gate76inter2));
  inv1  gate3000(.a(s_350), .O(gate76inter3));
  inv1  gate3001(.a(s_351), .O(gate76inter4));
  nand2 gate3002(.a(gate76inter4), .b(gate76inter3), .O(gate76inter5));
  nor2  gate3003(.a(gate76inter5), .b(gate76inter2), .O(gate76inter6));
  inv1  gate3004(.a(G13), .O(gate76inter7));
  inv1  gate3005(.a(G317), .O(gate76inter8));
  nand2 gate3006(.a(gate76inter8), .b(gate76inter7), .O(gate76inter9));
  nand2 gate3007(.a(s_351), .b(gate76inter3), .O(gate76inter10));
  nor2  gate3008(.a(gate76inter10), .b(gate76inter9), .O(gate76inter11));
  nor2  gate3009(.a(gate76inter11), .b(gate76inter6), .O(gate76inter12));
  nand2 gate3010(.a(gate76inter12), .b(gate76inter1), .O(G397));
nand2 gate77( .a(G2), .b(G320), .O(G398) );
nand2 gate78( .a(G6), .b(G320), .O(G399) );
nand2 gate79( .a(G10), .b(G323), .O(G400) );

  xor2  gate617(.a(G323), .b(G14), .O(gate80inter0));
  nand2 gate618(.a(gate80inter0), .b(s_10), .O(gate80inter1));
  and2  gate619(.a(G323), .b(G14), .O(gate80inter2));
  inv1  gate620(.a(s_10), .O(gate80inter3));
  inv1  gate621(.a(s_11), .O(gate80inter4));
  nand2 gate622(.a(gate80inter4), .b(gate80inter3), .O(gate80inter5));
  nor2  gate623(.a(gate80inter5), .b(gate80inter2), .O(gate80inter6));
  inv1  gate624(.a(G14), .O(gate80inter7));
  inv1  gate625(.a(G323), .O(gate80inter8));
  nand2 gate626(.a(gate80inter8), .b(gate80inter7), .O(gate80inter9));
  nand2 gate627(.a(s_11), .b(gate80inter3), .O(gate80inter10));
  nor2  gate628(.a(gate80inter10), .b(gate80inter9), .O(gate80inter11));
  nor2  gate629(.a(gate80inter11), .b(gate80inter6), .O(gate80inter12));
  nand2 gate630(.a(gate80inter12), .b(gate80inter1), .O(G401));
nand2 gate81( .a(G3), .b(G326), .O(G402) );

  xor2  gate827(.a(G326), .b(G7), .O(gate82inter0));
  nand2 gate828(.a(gate82inter0), .b(s_40), .O(gate82inter1));
  and2  gate829(.a(G326), .b(G7), .O(gate82inter2));
  inv1  gate830(.a(s_40), .O(gate82inter3));
  inv1  gate831(.a(s_41), .O(gate82inter4));
  nand2 gate832(.a(gate82inter4), .b(gate82inter3), .O(gate82inter5));
  nor2  gate833(.a(gate82inter5), .b(gate82inter2), .O(gate82inter6));
  inv1  gate834(.a(G7), .O(gate82inter7));
  inv1  gate835(.a(G326), .O(gate82inter8));
  nand2 gate836(.a(gate82inter8), .b(gate82inter7), .O(gate82inter9));
  nand2 gate837(.a(s_41), .b(gate82inter3), .O(gate82inter10));
  nor2  gate838(.a(gate82inter10), .b(gate82inter9), .O(gate82inter11));
  nor2  gate839(.a(gate82inter11), .b(gate82inter6), .O(gate82inter12));
  nand2 gate840(.a(gate82inter12), .b(gate82inter1), .O(G403));
nand2 gate83( .a(G11), .b(G329), .O(G404) );

  xor2  gate2213(.a(G329), .b(G15), .O(gate84inter0));
  nand2 gate2214(.a(gate84inter0), .b(s_238), .O(gate84inter1));
  and2  gate2215(.a(G329), .b(G15), .O(gate84inter2));
  inv1  gate2216(.a(s_238), .O(gate84inter3));
  inv1  gate2217(.a(s_239), .O(gate84inter4));
  nand2 gate2218(.a(gate84inter4), .b(gate84inter3), .O(gate84inter5));
  nor2  gate2219(.a(gate84inter5), .b(gate84inter2), .O(gate84inter6));
  inv1  gate2220(.a(G15), .O(gate84inter7));
  inv1  gate2221(.a(G329), .O(gate84inter8));
  nand2 gate2222(.a(gate84inter8), .b(gate84inter7), .O(gate84inter9));
  nand2 gate2223(.a(s_239), .b(gate84inter3), .O(gate84inter10));
  nor2  gate2224(.a(gate84inter10), .b(gate84inter9), .O(gate84inter11));
  nor2  gate2225(.a(gate84inter11), .b(gate84inter6), .O(gate84inter12));
  nand2 gate2226(.a(gate84inter12), .b(gate84inter1), .O(G405));

  xor2  gate2857(.a(G332), .b(G4), .O(gate85inter0));
  nand2 gate2858(.a(gate85inter0), .b(s_330), .O(gate85inter1));
  and2  gate2859(.a(G332), .b(G4), .O(gate85inter2));
  inv1  gate2860(.a(s_330), .O(gate85inter3));
  inv1  gate2861(.a(s_331), .O(gate85inter4));
  nand2 gate2862(.a(gate85inter4), .b(gate85inter3), .O(gate85inter5));
  nor2  gate2863(.a(gate85inter5), .b(gate85inter2), .O(gate85inter6));
  inv1  gate2864(.a(G4), .O(gate85inter7));
  inv1  gate2865(.a(G332), .O(gate85inter8));
  nand2 gate2866(.a(gate85inter8), .b(gate85inter7), .O(gate85inter9));
  nand2 gate2867(.a(s_331), .b(gate85inter3), .O(gate85inter10));
  nor2  gate2868(.a(gate85inter10), .b(gate85inter9), .O(gate85inter11));
  nor2  gate2869(.a(gate85inter11), .b(gate85inter6), .O(gate85inter12));
  nand2 gate2870(.a(gate85inter12), .b(gate85inter1), .O(G406));

  xor2  gate1107(.a(G332), .b(G8), .O(gate86inter0));
  nand2 gate1108(.a(gate86inter0), .b(s_80), .O(gate86inter1));
  and2  gate1109(.a(G332), .b(G8), .O(gate86inter2));
  inv1  gate1110(.a(s_80), .O(gate86inter3));
  inv1  gate1111(.a(s_81), .O(gate86inter4));
  nand2 gate1112(.a(gate86inter4), .b(gate86inter3), .O(gate86inter5));
  nor2  gate1113(.a(gate86inter5), .b(gate86inter2), .O(gate86inter6));
  inv1  gate1114(.a(G8), .O(gate86inter7));
  inv1  gate1115(.a(G332), .O(gate86inter8));
  nand2 gate1116(.a(gate86inter8), .b(gate86inter7), .O(gate86inter9));
  nand2 gate1117(.a(s_81), .b(gate86inter3), .O(gate86inter10));
  nor2  gate1118(.a(gate86inter10), .b(gate86inter9), .O(gate86inter11));
  nor2  gate1119(.a(gate86inter11), .b(gate86inter6), .O(gate86inter12));
  nand2 gate1120(.a(gate86inter12), .b(gate86inter1), .O(G407));

  xor2  gate2409(.a(G335), .b(G12), .O(gate87inter0));
  nand2 gate2410(.a(gate87inter0), .b(s_266), .O(gate87inter1));
  and2  gate2411(.a(G335), .b(G12), .O(gate87inter2));
  inv1  gate2412(.a(s_266), .O(gate87inter3));
  inv1  gate2413(.a(s_267), .O(gate87inter4));
  nand2 gate2414(.a(gate87inter4), .b(gate87inter3), .O(gate87inter5));
  nor2  gate2415(.a(gate87inter5), .b(gate87inter2), .O(gate87inter6));
  inv1  gate2416(.a(G12), .O(gate87inter7));
  inv1  gate2417(.a(G335), .O(gate87inter8));
  nand2 gate2418(.a(gate87inter8), .b(gate87inter7), .O(gate87inter9));
  nand2 gate2419(.a(s_267), .b(gate87inter3), .O(gate87inter10));
  nor2  gate2420(.a(gate87inter10), .b(gate87inter9), .O(gate87inter11));
  nor2  gate2421(.a(gate87inter11), .b(gate87inter6), .O(gate87inter12));
  nand2 gate2422(.a(gate87inter12), .b(gate87inter1), .O(G408));

  xor2  gate1709(.a(G335), .b(G16), .O(gate88inter0));
  nand2 gate1710(.a(gate88inter0), .b(s_166), .O(gate88inter1));
  and2  gate1711(.a(G335), .b(G16), .O(gate88inter2));
  inv1  gate1712(.a(s_166), .O(gate88inter3));
  inv1  gate1713(.a(s_167), .O(gate88inter4));
  nand2 gate1714(.a(gate88inter4), .b(gate88inter3), .O(gate88inter5));
  nor2  gate1715(.a(gate88inter5), .b(gate88inter2), .O(gate88inter6));
  inv1  gate1716(.a(G16), .O(gate88inter7));
  inv1  gate1717(.a(G335), .O(gate88inter8));
  nand2 gate1718(.a(gate88inter8), .b(gate88inter7), .O(gate88inter9));
  nand2 gate1719(.a(s_167), .b(gate88inter3), .O(gate88inter10));
  nor2  gate1720(.a(gate88inter10), .b(gate88inter9), .O(gate88inter11));
  nor2  gate1721(.a(gate88inter11), .b(gate88inter6), .O(gate88inter12));
  nand2 gate1722(.a(gate88inter12), .b(gate88inter1), .O(G409));

  xor2  gate2885(.a(G338), .b(G17), .O(gate89inter0));
  nand2 gate2886(.a(gate89inter0), .b(s_334), .O(gate89inter1));
  and2  gate2887(.a(G338), .b(G17), .O(gate89inter2));
  inv1  gate2888(.a(s_334), .O(gate89inter3));
  inv1  gate2889(.a(s_335), .O(gate89inter4));
  nand2 gate2890(.a(gate89inter4), .b(gate89inter3), .O(gate89inter5));
  nor2  gate2891(.a(gate89inter5), .b(gate89inter2), .O(gate89inter6));
  inv1  gate2892(.a(G17), .O(gate89inter7));
  inv1  gate2893(.a(G338), .O(gate89inter8));
  nand2 gate2894(.a(gate89inter8), .b(gate89inter7), .O(gate89inter9));
  nand2 gate2895(.a(s_335), .b(gate89inter3), .O(gate89inter10));
  nor2  gate2896(.a(gate89inter10), .b(gate89inter9), .O(gate89inter11));
  nor2  gate2897(.a(gate89inter11), .b(gate89inter6), .O(gate89inter12));
  nand2 gate2898(.a(gate89inter12), .b(gate89inter1), .O(G410));
nand2 gate90( .a(G21), .b(G338), .O(G411) );

  xor2  gate841(.a(G341), .b(G25), .O(gate91inter0));
  nand2 gate842(.a(gate91inter0), .b(s_42), .O(gate91inter1));
  and2  gate843(.a(G341), .b(G25), .O(gate91inter2));
  inv1  gate844(.a(s_42), .O(gate91inter3));
  inv1  gate845(.a(s_43), .O(gate91inter4));
  nand2 gate846(.a(gate91inter4), .b(gate91inter3), .O(gate91inter5));
  nor2  gate847(.a(gate91inter5), .b(gate91inter2), .O(gate91inter6));
  inv1  gate848(.a(G25), .O(gate91inter7));
  inv1  gate849(.a(G341), .O(gate91inter8));
  nand2 gate850(.a(gate91inter8), .b(gate91inter7), .O(gate91inter9));
  nand2 gate851(.a(s_43), .b(gate91inter3), .O(gate91inter10));
  nor2  gate852(.a(gate91inter10), .b(gate91inter9), .O(gate91inter11));
  nor2  gate853(.a(gate91inter11), .b(gate91inter6), .O(gate91inter12));
  nand2 gate854(.a(gate91inter12), .b(gate91inter1), .O(G412));
nand2 gate92( .a(G29), .b(G341), .O(G413) );

  xor2  gate2003(.a(G344), .b(G18), .O(gate93inter0));
  nand2 gate2004(.a(gate93inter0), .b(s_208), .O(gate93inter1));
  and2  gate2005(.a(G344), .b(G18), .O(gate93inter2));
  inv1  gate2006(.a(s_208), .O(gate93inter3));
  inv1  gate2007(.a(s_209), .O(gate93inter4));
  nand2 gate2008(.a(gate93inter4), .b(gate93inter3), .O(gate93inter5));
  nor2  gate2009(.a(gate93inter5), .b(gate93inter2), .O(gate93inter6));
  inv1  gate2010(.a(G18), .O(gate93inter7));
  inv1  gate2011(.a(G344), .O(gate93inter8));
  nand2 gate2012(.a(gate93inter8), .b(gate93inter7), .O(gate93inter9));
  nand2 gate2013(.a(s_209), .b(gate93inter3), .O(gate93inter10));
  nor2  gate2014(.a(gate93inter10), .b(gate93inter9), .O(gate93inter11));
  nor2  gate2015(.a(gate93inter11), .b(gate93inter6), .O(gate93inter12));
  nand2 gate2016(.a(gate93inter12), .b(gate93inter1), .O(G414));

  xor2  gate2731(.a(G344), .b(G22), .O(gate94inter0));
  nand2 gate2732(.a(gate94inter0), .b(s_312), .O(gate94inter1));
  and2  gate2733(.a(G344), .b(G22), .O(gate94inter2));
  inv1  gate2734(.a(s_312), .O(gate94inter3));
  inv1  gate2735(.a(s_313), .O(gate94inter4));
  nand2 gate2736(.a(gate94inter4), .b(gate94inter3), .O(gate94inter5));
  nor2  gate2737(.a(gate94inter5), .b(gate94inter2), .O(gate94inter6));
  inv1  gate2738(.a(G22), .O(gate94inter7));
  inv1  gate2739(.a(G344), .O(gate94inter8));
  nand2 gate2740(.a(gate94inter8), .b(gate94inter7), .O(gate94inter9));
  nand2 gate2741(.a(s_313), .b(gate94inter3), .O(gate94inter10));
  nor2  gate2742(.a(gate94inter10), .b(gate94inter9), .O(gate94inter11));
  nor2  gate2743(.a(gate94inter11), .b(gate94inter6), .O(gate94inter12));
  nand2 gate2744(.a(gate94inter12), .b(gate94inter1), .O(G415));
nand2 gate95( .a(G26), .b(G347), .O(G416) );

  xor2  gate1695(.a(G347), .b(G30), .O(gate96inter0));
  nand2 gate1696(.a(gate96inter0), .b(s_164), .O(gate96inter1));
  and2  gate1697(.a(G347), .b(G30), .O(gate96inter2));
  inv1  gate1698(.a(s_164), .O(gate96inter3));
  inv1  gate1699(.a(s_165), .O(gate96inter4));
  nand2 gate1700(.a(gate96inter4), .b(gate96inter3), .O(gate96inter5));
  nor2  gate1701(.a(gate96inter5), .b(gate96inter2), .O(gate96inter6));
  inv1  gate1702(.a(G30), .O(gate96inter7));
  inv1  gate1703(.a(G347), .O(gate96inter8));
  nand2 gate1704(.a(gate96inter8), .b(gate96inter7), .O(gate96inter9));
  nand2 gate1705(.a(s_165), .b(gate96inter3), .O(gate96inter10));
  nor2  gate1706(.a(gate96inter10), .b(gate96inter9), .O(gate96inter11));
  nor2  gate1707(.a(gate96inter11), .b(gate96inter6), .O(gate96inter12));
  nand2 gate1708(.a(gate96inter12), .b(gate96inter1), .O(G417));

  xor2  gate1569(.a(G350), .b(G19), .O(gate97inter0));
  nand2 gate1570(.a(gate97inter0), .b(s_146), .O(gate97inter1));
  and2  gate1571(.a(G350), .b(G19), .O(gate97inter2));
  inv1  gate1572(.a(s_146), .O(gate97inter3));
  inv1  gate1573(.a(s_147), .O(gate97inter4));
  nand2 gate1574(.a(gate97inter4), .b(gate97inter3), .O(gate97inter5));
  nor2  gate1575(.a(gate97inter5), .b(gate97inter2), .O(gate97inter6));
  inv1  gate1576(.a(G19), .O(gate97inter7));
  inv1  gate1577(.a(G350), .O(gate97inter8));
  nand2 gate1578(.a(gate97inter8), .b(gate97inter7), .O(gate97inter9));
  nand2 gate1579(.a(s_147), .b(gate97inter3), .O(gate97inter10));
  nor2  gate1580(.a(gate97inter10), .b(gate97inter9), .O(gate97inter11));
  nor2  gate1581(.a(gate97inter11), .b(gate97inter6), .O(gate97inter12));
  nand2 gate1582(.a(gate97inter12), .b(gate97inter1), .O(G418));

  xor2  gate2675(.a(G350), .b(G23), .O(gate98inter0));
  nand2 gate2676(.a(gate98inter0), .b(s_304), .O(gate98inter1));
  and2  gate2677(.a(G350), .b(G23), .O(gate98inter2));
  inv1  gate2678(.a(s_304), .O(gate98inter3));
  inv1  gate2679(.a(s_305), .O(gate98inter4));
  nand2 gate2680(.a(gate98inter4), .b(gate98inter3), .O(gate98inter5));
  nor2  gate2681(.a(gate98inter5), .b(gate98inter2), .O(gate98inter6));
  inv1  gate2682(.a(G23), .O(gate98inter7));
  inv1  gate2683(.a(G350), .O(gate98inter8));
  nand2 gate2684(.a(gate98inter8), .b(gate98inter7), .O(gate98inter9));
  nand2 gate2685(.a(s_305), .b(gate98inter3), .O(gate98inter10));
  nor2  gate2686(.a(gate98inter10), .b(gate98inter9), .O(gate98inter11));
  nor2  gate2687(.a(gate98inter11), .b(gate98inter6), .O(gate98inter12));
  nand2 gate2688(.a(gate98inter12), .b(gate98inter1), .O(G419));
nand2 gate99( .a(G27), .b(G353), .O(G420) );

  xor2  gate2619(.a(G353), .b(G31), .O(gate100inter0));
  nand2 gate2620(.a(gate100inter0), .b(s_296), .O(gate100inter1));
  and2  gate2621(.a(G353), .b(G31), .O(gate100inter2));
  inv1  gate2622(.a(s_296), .O(gate100inter3));
  inv1  gate2623(.a(s_297), .O(gate100inter4));
  nand2 gate2624(.a(gate100inter4), .b(gate100inter3), .O(gate100inter5));
  nor2  gate2625(.a(gate100inter5), .b(gate100inter2), .O(gate100inter6));
  inv1  gate2626(.a(G31), .O(gate100inter7));
  inv1  gate2627(.a(G353), .O(gate100inter8));
  nand2 gate2628(.a(gate100inter8), .b(gate100inter7), .O(gate100inter9));
  nand2 gate2629(.a(s_297), .b(gate100inter3), .O(gate100inter10));
  nor2  gate2630(.a(gate100inter10), .b(gate100inter9), .O(gate100inter11));
  nor2  gate2631(.a(gate100inter11), .b(gate100inter6), .O(gate100inter12));
  nand2 gate2632(.a(gate100inter12), .b(gate100inter1), .O(G421));
nand2 gate101( .a(G20), .b(G356), .O(G422) );
nand2 gate102( .a(G24), .b(G356), .O(G423) );
nand2 gate103( .a(G28), .b(G359), .O(G424) );
nand2 gate104( .a(G32), .b(G359), .O(G425) );
nand2 gate105( .a(G362), .b(G363), .O(G426) );
nand2 gate106( .a(G364), .b(G365), .O(G429) );

  xor2  gate2479(.a(G367), .b(G366), .O(gate107inter0));
  nand2 gate2480(.a(gate107inter0), .b(s_276), .O(gate107inter1));
  and2  gate2481(.a(G367), .b(G366), .O(gate107inter2));
  inv1  gate2482(.a(s_276), .O(gate107inter3));
  inv1  gate2483(.a(s_277), .O(gate107inter4));
  nand2 gate2484(.a(gate107inter4), .b(gate107inter3), .O(gate107inter5));
  nor2  gate2485(.a(gate107inter5), .b(gate107inter2), .O(gate107inter6));
  inv1  gate2486(.a(G366), .O(gate107inter7));
  inv1  gate2487(.a(G367), .O(gate107inter8));
  nand2 gate2488(.a(gate107inter8), .b(gate107inter7), .O(gate107inter9));
  nand2 gate2489(.a(s_277), .b(gate107inter3), .O(gate107inter10));
  nor2  gate2490(.a(gate107inter10), .b(gate107inter9), .O(gate107inter11));
  nor2  gate2491(.a(gate107inter11), .b(gate107inter6), .O(gate107inter12));
  nand2 gate2492(.a(gate107inter12), .b(gate107inter1), .O(G432));
nand2 gate108( .a(G368), .b(G369), .O(G435) );

  xor2  gate1653(.a(G371), .b(G370), .O(gate109inter0));
  nand2 gate1654(.a(gate109inter0), .b(s_158), .O(gate109inter1));
  and2  gate1655(.a(G371), .b(G370), .O(gate109inter2));
  inv1  gate1656(.a(s_158), .O(gate109inter3));
  inv1  gate1657(.a(s_159), .O(gate109inter4));
  nand2 gate1658(.a(gate109inter4), .b(gate109inter3), .O(gate109inter5));
  nor2  gate1659(.a(gate109inter5), .b(gate109inter2), .O(gate109inter6));
  inv1  gate1660(.a(G370), .O(gate109inter7));
  inv1  gate1661(.a(G371), .O(gate109inter8));
  nand2 gate1662(.a(gate109inter8), .b(gate109inter7), .O(gate109inter9));
  nand2 gate1663(.a(s_159), .b(gate109inter3), .O(gate109inter10));
  nor2  gate1664(.a(gate109inter10), .b(gate109inter9), .O(gate109inter11));
  nor2  gate1665(.a(gate109inter11), .b(gate109inter6), .O(gate109inter12));
  nand2 gate1666(.a(gate109inter12), .b(gate109inter1), .O(G438));
nand2 gate110( .a(G372), .b(G373), .O(G441) );

  xor2  gate911(.a(G375), .b(G374), .O(gate111inter0));
  nand2 gate912(.a(gate111inter0), .b(s_52), .O(gate111inter1));
  and2  gate913(.a(G375), .b(G374), .O(gate111inter2));
  inv1  gate914(.a(s_52), .O(gate111inter3));
  inv1  gate915(.a(s_53), .O(gate111inter4));
  nand2 gate916(.a(gate111inter4), .b(gate111inter3), .O(gate111inter5));
  nor2  gate917(.a(gate111inter5), .b(gate111inter2), .O(gate111inter6));
  inv1  gate918(.a(G374), .O(gate111inter7));
  inv1  gate919(.a(G375), .O(gate111inter8));
  nand2 gate920(.a(gate111inter8), .b(gate111inter7), .O(gate111inter9));
  nand2 gate921(.a(s_53), .b(gate111inter3), .O(gate111inter10));
  nor2  gate922(.a(gate111inter10), .b(gate111inter9), .O(gate111inter11));
  nor2  gate923(.a(gate111inter11), .b(gate111inter6), .O(gate111inter12));
  nand2 gate924(.a(gate111inter12), .b(gate111inter1), .O(G444));
nand2 gate112( .a(G376), .b(G377), .O(G447) );
nand2 gate113( .a(G378), .b(G379), .O(G450) );

  xor2  gate2353(.a(G381), .b(G380), .O(gate114inter0));
  nand2 gate2354(.a(gate114inter0), .b(s_258), .O(gate114inter1));
  and2  gate2355(.a(G381), .b(G380), .O(gate114inter2));
  inv1  gate2356(.a(s_258), .O(gate114inter3));
  inv1  gate2357(.a(s_259), .O(gate114inter4));
  nand2 gate2358(.a(gate114inter4), .b(gate114inter3), .O(gate114inter5));
  nor2  gate2359(.a(gate114inter5), .b(gate114inter2), .O(gate114inter6));
  inv1  gate2360(.a(G380), .O(gate114inter7));
  inv1  gate2361(.a(G381), .O(gate114inter8));
  nand2 gate2362(.a(gate114inter8), .b(gate114inter7), .O(gate114inter9));
  nand2 gate2363(.a(s_259), .b(gate114inter3), .O(gate114inter10));
  nor2  gate2364(.a(gate114inter10), .b(gate114inter9), .O(gate114inter11));
  nor2  gate2365(.a(gate114inter11), .b(gate114inter6), .O(gate114inter12));
  nand2 gate2366(.a(gate114inter12), .b(gate114inter1), .O(G453));

  xor2  gate2969(.a(G383), .b(G382), .O(gate115inter0));
  nand2 gate2970(.a(gate115inter0), .b(s_346), .O(gate115inter1));
  and2  gate2971(.a(G383), .b(G382), .O(gate115inter2));
  inv1  gate2972(.a(s_346), .O(gate115inter3));
  inv1  gate2973(.a(s_347), .O(gate115inter4));
  nand2 gate2974(.a(gate115inter4), .b(gate115inter3), .O(gate115inter5));
  nor2  gate2975(.a(gate115inter5), .b(gate115inter2), .O(gate115inter6));
  inv1  gate2976(.a(G382), .O(gate115inter7));
  inv1  gate2977(.a(G383), .O(gate115inter8));
  nand2 gate2978(.a(gate115inter8), .b(gate115inter7), .O(gate115inter9));
  nand2 gate2979(.a(s_347), .b(gate115inter3), .O(gate115inter10));
  nor2  gate2980(.a(gate115inter10), .b(gate115inter9), .O(gate115inter11));
  nor2  gate2981(.a(gate115inter11), .b(gate115inter6), .O(gate115inter12));
  nand2 gate2982(.a(gate115inter12), .b(gate115inter1), .O(G456));

  xor2  gate1485(.a(G385), .b(G384), .O(gate116inter0));
  nand2 gate1486(.a(gate116inter0), .b(s_134), .O(gate116inter1));
  and2  gate1487(.a(G385), .b(G384), .O(gate116inter2));
  inv1  gate1488(.a(s_134), .O(gate116inter3));
  inv1  gate1489(.a(s_135), .O(gate116inter4));
  nand2 gate1490(.a(gate116inter4), .b(gate116inter3), .O(gate116inter5));
  nor2  gate1491(.a(gate116inter5), .b(gate116inter2), .O(gate116inter6));
  inv1  gate1492(.a(G384), .O(gate116inter7));
  inv1  gate1493(.a(G385), .O(gate116inter8));
  nand2 gate1494(.a(gate116inter8), .b(gate116inter7), .O(gate116inter9));
  nand2 gate1495(.a(s_135), .b(gate116inter3), .O(gate116inter10));
  nor2  gate1496(.a(gate116inter10), .b(gate116inter9), .O(gate116inter11));
  nor2  gate1497(.a(gate116inter11), .b(gate116inter6), .O(gate116inter12));
  nand2 gate1498(.a(gate116inter12), .b(gate116inter1), .O(G459));

  xor2  gate1947(.a(G387), .b(G386), .O(gate117inter0));
  nand2 gate1948(.a(gate117inter0), .b(s_200), .O(gate117inter1));
  and2  gate1949(.a(G387), .b(G386), .O(gate117inter2));
  inv1  gate1950(.a(s_200), .O(gate117inter3));
  inv1  gate1951(.a(s_201), .O(gate117inter4));
  nand2 gate1952(.a(gate117inter4), .b(gate117inter3), .O(gate117inter5));
  nor2  gate1953(.a(gate117inter5), .b(gate117inter2), .O(gate117inter6));
  inv1  gate1954(.a(G386), .O(gate117inter7));
  inv1  gate1955(.a(G387), .O(gate117inter8));
  nand2 gate1956(.a(gate117inter8), .b(gate117inter7), .O(gate117inter9));
  nand2 gate1957(.a(s_201), .b(gate117inter3), .O(gate117inter10));
  nor2  gate1958(.a(gate117inter10), .b(gate117inter9), .O(gate117inter11));
  nor2  gate1959(.a(gate117inter11), .b(gate117inter6), .O(gate117inter12));
  nand2 gate1960(.a(gate117inter12), .b(gate117inter1), .O(G462));

  xor2  gate1597(.a(G389), .b(G388), .O(gate118inter0));
  nand2 gate1598(.a(gate118inter0), .b(s_150), .O(gate118inter1));
  and2  gate1599(.a(G389), .b(G388), .O(gate118inter2));
  inv1  gate1600(.a(s_150), .O(gate118inter3));
  inv1  gate1601(.a(s_151), .O(gate118inter4));
  nand2 gate1602(.a(gate118inter4), .b(gate118inter3), .O(gate118inter5));
  nor2  gate1603(.a(gate118inter5), .b(gate118inter2), .O(gate118inter6));
  inv1  gate1604(.a(G388), .O(gate118inter7));
  inv1  gate1605(.a(G389), .O(gate118inter8));
  nand2 gate1606(.a(gate118inter8), .b(gate118inter7), .O(gate118inter9));
  nand2 gate1607(.a(s_151), .b(gate118inter3), .O(gate118inter10));
  nor2  gate1608(.a(gate118inter10), .b(gate118inter9), .O(gate118inter11));
  nor2  gate1609(.a(gate118inter11), .b(gate118inter6), .O(gate118inter12));
  nand2 gate1610(.a(gate118inter12), .b(gate118inter1), .O(G465));

  xor2  gate2395(.a(G391), .b(G390), .O(gate119inter0));
  nand2 gate2396(.a(gate119inter0), .b(s_264), .O(gate119inter1));
  and2  gate2397(.a(G391), .b(G390), .O(gate119inter2));
  inv1  gate2398(.a(s_264), .O(gate119inter3));
  inv1  gate2399(.a(s_265), .O(gate119inter4));
  nand2 gate2400(.a(gate119inter4), .b(gate119inter3), .O(gate119inter5));
  nor2  gate2401(.a(gate119inter5), .b(gate119inter2), .O(gate119inter6));
  inv1  gate2402(.a(G390), .O(gate119inter7));
  inv1  gate2403(.a(G391), .O(gate119inter8));
  nand2 gate2404(.a(gate119inter8), .b(gate119inter7), .O(gate119inter9));
  nand2 gate2405(.a(s_265), .b(gate119inter3), .O(gate119inter10));
  nor2  gate2406(.a(gate119inter10), .b(gate119inter9), .O(gate119inter11));
  nor2  gate2407(.a(gate119inter11), .b(gate119inter6), .O(gate119inter12));
  nand2 gate2408(.a(gate119inter12), .b(gate119inter1), .O(G468));

  xor2  gate1905(.a(G393), .b(G392), .O(gate120inter0));
  nand2 gate1906(.a(gate120inter0), .b(s_194), .O(gate120inter1));
  and2  gate1907(.a(G393), .b(G392), .O(gate120inter2));
  inv1  gate1908(.a(s_194), .O(gate120inter3));
  inv1  gate1909(.a(s_195), .O(gate120inter4));
  nand2 gate1910(.a(gate120inter4), .b(gate120inter3), .O(gate120inter5));
  nor2  gate1911(.a(gate120inter5), .b(gate120inter2), .O(gate120inter6));
  inv1  gate1912(.a(G392), .O(gate120inter7));
  inv1  gate1913(.a(G393), .O(gate120inter8));
  nand2 gate1914(.a(gate120inter8), .b(gate120inter7), .O(gate120inter9));
  nand2 gate1915(.a(s_195), .b(gate120inter3), .O(gate120inter10));
  nor2  gate1916(.a(gate120inter10), .b(gate120inter9), .O(gate120inter11));
  nor2  gate1917(.a(gate120inter11), .b(gate120inter6), .O(gate120inter12));
  nand2 gate1918(.a(gate120inter12), .b(gate120inter1), .O(G471));
nand2 gate121( .a(G394), .b(G395), .O(G474) );
nand2 gate122( .a(G396), .b(G397), .O(G477) );

  xor2  gate3067(.a(G399), .b(G398), .O(gate123inter0));
  nand2 gate3068(.a(gate123inter0), .b(s_360), .O(gate123inter1));
  and2  gate3069(.a(G399), .b(G398), .O(gate123inter2));
  inv1  gate3070(.a(s_360), .O(gate123inter3));
  inv1  gate3071(.a(s_361), .O(gate123inter4));
  nand2 gate3072(.a(gate123inter4), .b(gate123inter3), .O(gate123inter5));
  nor2  gate3073(.a(gate123inter5), .b(gate123inter2), .O(gate123inter6));
  inv1  gate3074(.a(G398), .O(gate123inter7));
  inv1  gate3075(.a(G399), .O(gate123inter8));
  nand2 gate3076(.a(gate123inter8), .b(gate123inter7), .O(gate123inter9));
  nand2 gate3077(.a(s_361), .b(gate123inter3), .O(gate123inter10));
  nor2  gate3078(.a(gate123inter10), .b(gate123inter9), .O(gate123inter11));
  nor2  gate3079(.a(gate123inter11), .b(gate123inter6), .O(gate123inter12));
  nand2 gate3080(.a(gate123inter12), .b(gate123inter1), .O(G480));
nand2 gate124( .a(G400), .b(G401), .O(G483) );

  xor2  gate869(.a(G403), .b(G402), .O(gate125inter0));
  nand2 gate870(.a(gate125inter0), .b(s_46), .O(gate125inter1));
  and2  gate871(.a(G403), .b(G402), .O(gate125inter2));
  inv1  gate872(.a(s_46), .O(gate125inter3));
  inv1  gate873(.a(s_47), .O(gate125inter4));
  nand2 gate874(.a(gate125inter4), .b(gate125inter3), .O(gate125inter5));
  nor2  gate875(.a(gate125inter5), .b(gate125inter2), .O(gate125inter6));
  inv1  gate876(.a(G402), .O(gate125inter7));
  inv1  gate877(.a(G403), .O(gate125inter8));
  nand2 gate878(.a(gate125inter8), .b(gate125inter7), .O(gate125inter9));
  nand2 gate879(.a(s_47), .b(gate125inter3), .O(gate125inter10));
  nor2  gate880(.a(gate125inter10), .b(gate125inter9), .O(gate125inter11));
  nor2  gate881(.a(gate125inter11), .b(gate125inter6), .O(gate125inter12));
  nand2 gate882(.a(gate125inter12), .b(gate125inter1), .O(G486));
nand2 gate126( .a(G404), .b(G405), .O(G489) );
nand2 gate127( .a(G406), .b(G407), .O(G492) );

  xor2  gate2115(.a(G409), .b(G408), .O(gate128inter0));
  nand2 gate2116(.a(gate128inter0), .b(s_224), .O(gate128inter1));
  and2  gate2117(.a(G409), .b(G408), .O(gate128inter2));
  inv1  gate2118(.a(s_224), .O(gate128inter3));
  inv1  gate2119(.a(s_225), .O(gate128inter4));
  nand2 gate2120(.a(gate128inter4), .b(gate128inter3), .O(gate128inter5));
  nor2  gate2121(.a(gate128inter5), .b(gate128inter2), .O(gate128inter6));
  inv1  gate2122(.a(G408), .O(gate128inter7));
  inv1  gate2123(.a(G409), .O(gate128inter8));
  nand2 gate2124(.a(gate128inter8), .b(gate128inter7), .O(gate128inter9));
  nand2 gate2125(.a(s_225), .b(gate128inter3), .O(gate128inter10));
  nor2  gate2126(.a(gate128inter10), .b(gate128inter9), .O(gate128inter11));
  nor2  gate2127(.a(gate128inter11), .b(gate128inter6), .O(gate128inter12));
  nand2 gate2128(.a(gate128inter12), .b(gate128inter1), .O(G495));
nand2 gate129( .a(G410), .b(G411), .O(G498) );
nand2 gate130( .a(G412), .b(G413), .O(G501) );
nand2 gate131( .a(G414), .b(G415), .O(G504) );
nand2 gate132( .a(G416), .b(G417), .O(G507) );

  xor2  gate2829(.a(G419), .b(G418), .O(gate133inter0));
  nand2 gate2830(.a(gate133inter0), .b(s_326), .O(gate133inter1));
  and2  gate2831(.a(G419), .b(G418), .O(gate133inter2));
  inv1  gate2832(.a(s_326), .O(gate133inter3));
  inv1  gate2833(.a(s_327), .O(gate133inter4));
  nand2 gate2834(.a(gate133inter4), .b(gate133inter3), .O(gate133inter5));
  nor2  gate2835(.a(gate133inter5), .b(gate133inter2), .O(gate133inter6));
  inv1  gate2836(.a(G418), .O(gate133inter7));
  inv1  gate2837(.a(G419), .O(gate133inter8));
  nand2 gate2838(.a(gate133inter8), .b(gate133inter7), .O(gate133inter9));
  nand2 gate2839(.a(s_327), .b(gate133inter3), .O(gate133inter10));
  nor2  gate2840(.a(gate133inter10), .b(gate133inter9), .O(gate133inter11));
  nor2  gate2841(.a(gate133inter11), .b(gate133inter6), .O(gate133inter12));
  nand2 gate2842(.a(gate133inter12), .b(gate133inter1), .O(G510));

  xor2  gate1135(.a(G421), .b(G420), .O(gate134inter0));
  nand2 gate1136(.a(gate134inter0), .b(s_84), .O(gate134inter1));
  and2  gate1137(.a(G421), .b(G420), .O(gate134inter2));
  inv1  gate1138(.a(s_84), .O(gate134inter3));
  inv1  gate1139(.a(s_85), .O(gate134inter4));
  nand2 gate1140(.a(gate134inter4), .b(gate134inter3), .O(gate134inter5));
  nor2  gate1141(.a(gate134inter5), .b(gate134inter2), .O(gate134inter6));
  inv1  gate1142(.a(G420), .O(gate134inter7));
  inv1  gate1143(.a(G421), .O(gate134inter8));
  nand2 gate1144(.a(gate134inter8), .b(gate134inter7), .O(gate134inter9));
  nand2 gate1145(.a(s_85), .b(gate134inter3), .O(gate134inter10));
  nor2  gate1146(.a(gate134inter10), .b(gate134inter9), .O(gate134inter11));
  nor2  gate1147(.a(gate134inter11), .b(gate134inter6), .O(gate134inter12));
  nand2 gate1148(.a(gate134inter12), .b(gate134inter1), .O(G513));
nand2 gate135( .a(G422), .b(G423), .O(G516) );
nand2 gate136( .a(G424), .b(G425), .O(G519) );

  xor2  gate2129(.a(G429), .b(G426), .O(gate137inter0));
  nand2 gate2130(.a(gate137inter0), .b(s_226), .O(gate137inter1));
  and2  gate2131(.a(G429), .b(G426), .O(gate137inter2));
  inv1  gate2132(.a(s_226), .O(gate137inter3));
  inv1  gate2133(.a(s_227), .O(gate137inter4));
  nand2 gate2134(.a(gate137inter4), .b(gate137inter3), .O(gate137inter5));
  nor2  gate2135(.a(gate137inter5), .b(gate137inter2), .O(gate137inter6));
  inv1  gate2136(.a(G426), .O(gate137inter7));
  inv1  gate2137(.a(G429), .O(gate137inter8));
  nand2 gate2138(.a(gate137inter8), .b(gate137inter7), .O(gate137inter9));
  nand2 gate2139(.a(s_227), .b(gate137inter3), .O(gate137inter10));
  nor2  gate2140(.a(gate137inter10), .b(gate137inter9), .O(gate137inter11));
  nor2  gate2141(.a(gate137inter11), .b(gate137inter6), .O(gate137inter12));
  nand2 gate2142(.a(gate137inter12), .b(gate137inter1), .O(G522));
nand2 gate138( .a(G432), .b(G435), .O(G525) );

  xor2  gate1989(.a(G441), .b(G438), .O(gate139inter0));
  nand2 gate1990(.a(gate139inter0), .b(s_206), .O(gate139inter1));
  and2  gate1991(.a(G441), .b(G438), .O(gate139inter2));
  inv1  gate1992(.a(s_206), .O(gate139inter3));
  inv1  gate1993(.a(s_207), .O(gate139inter4));
  nand2 gate1994(.a(gate139inter4), .b(gate139inter3), .O(gate139inter5));
  nor2  gate1995(.a(gate139inter5), .b(gate139inter2), .O(gate139inter6));
  inv1  gate1996(.a(G438), .O(gate139inter7));
  inv1  gate1997(.a(G441), .O(gate139inter8));
  nand2 gate1998(.a(gate139inter8), .b(gate139inter7), .O(gate139inter9));
  nand2 gate1999(.a(s_207), .b(gate139inter3), .O(gate139inter10));
  nor2  gate2000(.a(gate139inter10), .b(gate139inter9), .O(gate139inter11));
  nor2  gate2001(.a(gate139inter11), .b(gate139inter6), .O(gate139inter12));
  nand2 gate2002(.a(gate139inter12), .b(gate139inter1), .O(G528));
nand2 gate140( .a(G444), .b(G447), .O(G531) );
nand2 gate141( .a(G450), .b(G453), .O(G534) );
nand2 gate142( .a(G456), .b(G459), .O(G537) );

  xor2  gate2059(.a(G465), .b(G462), .O(gate143inter0));
  nand2 gate2060(.a(gate143inter0), .b(s_216), .O(gate143inter1));
  and2  gate2061(.a(G465), .b(G462), .O(gate143inter2));
  inv1  gate2062(.a(s_216), .O(gate143inter3));
  inv1  gate2063(.a(s_217), .O(gate143inter4));
  nand2 gate2064(.a(gate143inter4), .b(gate143inter3), .O(gate143inter5));
  nor2  gate2065(.a(gate143inter5), .b(gate143inter2), .O(gate143inter6));
  inv1  gate2066(.a(G462), .O(gate143inter7));
  inv1  gate2067(.a(G465), .O(gate143inter8));
  nand2 gate2068(.a(gate143inter8), .b(gate143inter7), .O(gate143inter9));
  nand2 gate2069(.a(s_217), .b(gate143inter3), .O(gate143inter10));
  nor2  gate2070(.a(gate143inter10), .b(gate143inter9), .O(gate143inter11));
  nor2  gate2071(.a(gate143inter11), .b(gate143inter6), .O(gate143inter12));
  nand2 gate2072(.a(gate143inter12), .b(gate143inter1), .O(G540));
nand2 gate144( .a(G468), .b(G471), .O(G543) );

  xor2  gate1149(.a(G477), .b(G474), .O(gate145inter0));
  nand2 gate1150(.a(gate145inter0), .b(s_86), .O(gate145inter1));
  and2  gate1151(.a(G477), .b(G474), .O(gate145inter2));
  inv1  gate1152(.a(s_86), .O(gate145inter3));
  inv1  gate1153(.a(s_87), .O(gate145inter4));
  nand2 gate1154(.a(gate145inter4), .b(gate145inter3), .O(gate145inter5));
  nor2  gate1155(.a(gate145inter5), .b(gate145inter2), .O(gate145inter6));
  inv1  gate1156(.a(G474), .O(gate145inter7));
  inv1  gate1157(.a(G477), .O(gate145inter8));
  nand2 gate1158(.a(gate145inter8), .b(gate145inter7), .O(gate145inter9));
  nand2 gate1159(.a(s_87), .b(gate145inter3), .O(gate145inter10));
  nor2  gate1160(.a(gate145inter10), .b(gate145inter9), .O(gate145inter11));
  nor2  gate1161(.a(gate145inter11), .b(gate145inter6), .O(gate145inter12));
  nand2 gate1162(.a(gate145inter12), .b(gate145inter1), .O(G546));
nand2 gate146( .a(G480), .b(G483), .O(G549) );

  xor2  gate1765(.a(G489), .b(G486), .O(gate147inter0));
  nand2 gate1766(.a(gate147inter0), .b(s_174), .O(gate147inter1));
  and2  gate1767(.a(G489), .b(G486), .O(gate147inter2));
  inv1  gate1768(.a(s_174), .O(gate147inter3));
  inv1  gate1769(.a(s_175), .O(gate147inter4));
  nand2 gate1770(.a(gate147inter4), .b(gate147inter3), .O(gate147inter5));
  nor2  gate1771(.a(gate147inter5), .b(gate147inter2), .O(gate147inter6));
  inv1  gate1772(.a(G486), .O(gate147inter7));
  inv1  gate1773(.a(G489), .O(gate147inter8));
  nand2 gate1774(.a(gate147inter8), .b(gate147inter7), .O(gate147inter9));
  nand2 gate1775(.a(s_175), .b(gate147inter3), .O(gate147inter10));
  nor2  gate1776(.a(gate147inter10), .b(gate147inter9), .O(gate147inter11));
  nor2  gate1777(.a(gate147inter11), .b(gate147inter6), .O(gate147inter12));
  nand2 gate1778(.a(gate147inter12), .b(gate147inter1), .O(G552));
nand2 gate148( .a(G492), .b(G495), .O(G555) );

  xor2  gate3025(.a(G501), .b(G498), .O(gate149inter0));
  nand2 gate3026(.a(gate149inter0), .b(s_354), .O(gate149inter1));
  and2  gate3027(.a(G501), .b(G498), .O(gate149inter2));
  inv1  gate3028(.a(s_354), .O(gate149inter3));
  inv1  gate3029(.a(s_355), .O(gate149inter4));
  nand2 gate3030(.a(gate149inter4), .b(gate149inter3), .O(gate149inter5));
  nor2  gate3031(.a(gate149inter5), .b(gate149inter2), .O(gate149inter6));
  inv1  gate3032(.a(G498), .O(gate149inter7));
  inv1  gate3033(.a(G501), .O(gate149inter8));
  nand2 gate3034(.a(gate149inter8), .b(gate149inter7), .O(gate149inter9));
  nand2 gate3035(.a(s_355), .b(gate149inter3), .O(gate149inter10));
  nor2  gate3036(.a(gate149inter10), .b(gate149inter9), .O(gate149inter11));
  nor2  gate3037(.a(gate149inter11), .b(gate149inter6), .O(gate149inter12));
  nand2 gate3038(.a(gate149inter12), .b(gate149inter1), .O(G558));

  xor2  gate2703(.a(G507), .b(G504), .O(gate150inter0));
  nand2 gate2704(.a(gate150inter0), .b(s_308), .O(gate150inter1));
  and2  gate2705(.a(G507), .b(G504), .O(gate150inter2));
  inv1  gate2706(.a(s_308), .O(gate150inter3));
  inv1  gate2707(.a(s_309), .O(gate150inter4));
  nand2 gate2708(.a(gate150inter4), .b(gate150inter3), .O(gate150inter5));
  nor2  gate2709(.a(gate150inter5), .b(gate150inter2), .O(gate150inter6));
  inv1  gate2710(.a(G504), .O(gate150inter7));
  inv1  gate2711(.a(G507), .O(gate150inter8));
  nand2 gate2712(.a(gate150inter8), .b(gate150inter7), .O(gate150inter9));
  nand2 gate2713(.a(s_309), .b(gate150inter3), .O(gate150inter10));
  nor2  gate2714(.a(gate150inter10), .b(gate150inter9), .O(gate150inter11));
  nor2  gate2715(.a(gate150inter11), .b(gate150inter6), .O(gate150inter12));
  nand2 gate2716(.a(gate150inter12), .b(gate150inter1), .O(G561));

  xor2  gate2717(.a(G513), .b(G510), .O(gate151inter0));
  nand2 gate2718(.a(gate151inter0), .b(s_310), .O(gate151inter1));
  and2  gate2719(.a(G513), .b(G510), .O(gate151inter2));
  inv1  gate2720(.a(s_310), .O(gate151inter3));
  inv1  gate2721(.a(s_311), .O(gate151inter4));
  nand2 gate2722(.a(gate151inter4), .b(gate151inter3), .O(gate151inter5));
  nor2  gate2723(.a(gate151inter5), .b(gate151inter2), .O(gate151inter6));
  inv1  gate2724(.a(G510), .O(gate151inter7));
  inv1  gate2725(.a(G513), .O(gate151inter8));
  nand2 gate2726(.a(gate151inter8), .b(gate151inter7), .O(gate151inter9));
  nand2 gate2727(.a(s_311), .b(gate151inter3), .O(gate151inter10));
  nor2  gate2728(.a(gate151inter10), .b(gate151inter9), .O(gate151inter11));
  nor2  gate2729(.a(gate151inter11), .b(gate151inter6), .O(gate151inter12));
  nand2 gate2730(.a(gate151inter12), .b(gate151inter1), .O(G564));

  xor2  gate757(.a(G519), .b(G516), .O(gate152inter0));
  nand2 gate758(.a(gate152inter0), .b(s_30), .O(gate152inter1));
  and2  gate759(.a(G519), .b(G516), .O(gate152inter2));
  inv1  gate760(.a(s_30), .O(gate152inter3));
  inv1  gate761(.a(s_31), .O(gate152inter4));
  nand2 gate762(.a(gate152inter4), .b(gate152inter3), .O(gate152inter5));
  nor2  gate763(.a(gate152inter5), .b(gate152inter2), .O(gate152inter6));
  inv1  gate764(.a(G516), .O(gate152inter7));
  inv1  gate765(.a(G519), .O(gate152inter8));
  nand2 gate766(.a(gate152inter8), .b(gate152inter7), .O(gate152inter9));
  nand2 gate767(.a(s_31), .b(gate152inter3), .O(gate152inter10));
  nor2  gate768(.a(gate152inter10), .b(gate152inter9), .O(gate152inter11));
  nor2  gate769(.a(gate152inter11), .b(gate152inter6), .O(gate152inter12));
  nand2 gate770(.a(gate152inter12), .b(gate152inter1), .O(G567));

  xor2  gate729(.a(G522), .b(G426), .O(gate153inter0));
  nand2 gate730(.a(gate153inter0), .b(s_26), .O(gate153inter1));
  and2  gate731(.a(G522), .b(G426), .O(gate153inter2));
  inv1  gate732(.a(s_26), .O(gate153inter3));
  inv1  gate733(.a(s_27), .O(gate153inter4));
  nand2 gate734(.a(gate153inter4), .b(gate153inter3), .O(gate153inter5));
  nor2  gate735(.a(gate153inter5), .b(gate153inter2), .O(gate153inter6));
  inv1  gate736(.a(G426), .O(gate153inter7));
  inv1  gate737(.a(G522), .O(gate153inter8));
  nand2 gate738(.a(gate153inter8), .b(gate153inter7), .O(gate153inter9));
  nand2 gate739(.a(s_27), .b(gate153inter3), .O(gate153inter10));
  nor2  gate740(.a(gate153inter10), .b(gate153inter9), .O(gate153inter11));
  nor2  gate741(.a(gate153inter11), .b(gate153inter6), .O(gate153inter12));
  nand2 gate742(.a(gate153inter12), .b(gate153inter1), .O(G570));

  xor2  gate2241(.a(G522), .b(G429), .O(gate154inter0));
  nand2 gate2242(.a(gate154inter0), .b(s_242), .O(gate154inter1));
  and2  gate2243(.a(G522), .b(G429), .O(gate154inter2));
  inv1  gate2244(.a(s_242), .O(gate154inter3));
  inv1  gate2245(.a(s_243), .O(gate154inter4));
  nand2 gate2246(.a(gate154inter4), .b(gate154inter3), .O(gate154inter5));
  nor2  gate2247(.a(gate154inter5), .b(gate154inter2), .O(gate154inter6));
  inv1  gate2248(.a(G429), .O(gate154inter7));
  inv1  gate2249(.a(G522), .O(gate154inter8));
  nand2 gate2250(.a(gate154inter8), .b(gate154inter7), .O(gate154inter9));
  nand2 gate2251(.a(s_243), .b(gate154inter3), .O(gate154inter10));
  nor2  gate2252(.a(gate154inter10), .b(gate154inter9), .O(gate154inter11));
  nor2  gate2253(.a(gate154inter11), .b(gate154inter6), .O(gate154inter12));
  nand2 gate2254(.a(gate154inter12), .b(gate154inter1), .O(G571));
nand2 gate155( .a(G432), .b(G525), .O(G572) );
nand2 gate156( .a(G435), .b(G525), .O(G573) );

  xor2  gate547(.a(G528), .b(G438), .O(gate157inter0));
  nand2 gate548(.a(gate157inter0), .b(s_0), .O(gate157inter1));
  and2  gate549(.a(G528), .b(G438), .O(gate157inter2));
  inv1  gate550(.a(s_0), .O(gate157inter3));
  inv1  gate551(.a(s_1), .O(gate157inter4));
  nand2 gate552(.a(gate157inter4), .b(gate157inter3), .O(gate157inter5));
  nor2  gate553(.a(gate157inter5), .b(gate157inter2), .O(gate157inter6));
  inv1  gate554(.a(G438), .O(gate157inter7));
  inv1  gate555(.a(G528), .O(gate157inter8));
  nand2 gate556(.a(gate157inter8), .b(gate157inter7), .O(gate157inter9));
  nand2 gate557(.a(s_1), .b(gate157inter3), .O(gate157inter10));
  nor2  gate558(.a(gate157inter10), .b(gate157inter9), .O(gate157inter11));
  nor2  gate559(.a(gate157inter11), .b(gate157inter6), .O(gate157inter12));
  nand2 gate560(.a(gate157inter12), .b(gate157inter1), .O(G574));
nand2 gate158( .a(G441), .b(G528), .O(G575) );
nand2 gate159( .a(G444), .b(G531), .O(G576) );

  xor2  gate603(.a(G531), .b(G447), .O(gate160inter0));
  nand2 gate604(.a(gate160inter0), .b(s_8), .O(gate160inter1));
  and2  gate605(.a(G531), .b(G447), .O(gate160inter2));
  inv1  gate606(.a(s_8), .O(gate160inter3));
  inv1  gate607(.a(s_9), .O(gate160inter4));
  nand2 gate608(.a(gate160inter4), .b(gate160inter3), .O(gate160inter5));
  nor2  gate609(.a(gate160inter5), .b(gate160inter2), .O(gate160inter6));
  inv1  gate610(.a(G447), .O(gate160inter7));
  inv1  gate611(.a(G531), .O(gate160inter8));
  nand2 gate612(.a(gate160inter8), .b(gate160inter7), .O(gate160inter9));
  nand2 gate613(.a(s_9), .b(gate160inter3), .O(gate160inter10));
  nor2  gate614(.a(gate160inter10), .b(gate160inter9), .O(gate160inter11));
  nor2  gate615(.a(gate160inter11), .b(gate160inter6), .O(gate160inter12));
  nand2 gate616(.a(gate160inter12), .b(gate160inter1), .O(G577));

  xor2  gate1079(.a(G534), .b(G450), .O(gate161inter0));
  nand2 gate1080(.a(gate161inter0), .b(s_76), .O(gate161inter1));
  and2  gate1081(.a(G534), .b(G450), .O(gate161inter2));
  inv1  gate1082(.a(s_76), .O(gate161inter3));
  inv1  gate1083(.a(s_77), .O(gate161inter4));
  nand2 gate1084(.a(gate161inter4), .b(gate161inter3), .O(gate161inter5));
  nor2  gate1085(.a(gate161inter5), .b(gate161inter2), .O(gate161inter6));
  inv1  gate1086(.a(G450), .O(gate161inter7));
  inv1  gate1087(.a(G534), .O(gate161inter8));
  nand2 gate1088(.a(gate161inter8), .b(gate161inter7), .O(gate161inter9));
  nand2 gate1089(.a(s_77), .b(gate161inter3), .O(gate161inter10));
  nor2  gate1090(.a(gate161inter10), .b(gate161inter9), .O(gate161inter11));
  nor2  gate1091(.a(gate161inter11), .b(gate161inter6), .O(gate161inter12));
  nand2 gate1092(.a(gate161inter12), .b(gate161inter1), .O(G578));
nand2 gate162( .a(G453), .b(G534), .O(G579) );

  xor2  gate1415(.a(G537), .b(G456), .O(gate163inter0));
  nand2 gate1416(.a(gate163inter0), .b(s_124), .O(gate163inter1));
  and2  gate1417(.a(G537), .b(G456), .O(gate163inter2));
  inv1  gate1418(.a(s_124), .O(gate163inter3));
  inv1  gate1419(.a(s_125), .O(gate163inter4));
  nand2 gate1420(.a(gate163inter4), .b(gate163inter3), .O(gate163inter5));
  nor2  gate1421(.a(gate163inter5), .b(gate163inter2), .O(gate163inter6));
  inv1  gate1422(.a(G456), .O(gate163inter7));
  inv1  gate1423(.a(G537), .O(gate163inter8));
  nand2 gate1424(.a(gate163inter8), .b(gate163inter7), .O(gate163inter9));
  nand2 gate1425(.a(s_125), .b(gate163inter3), .O(gate163inter10));
  nor2  gate1426(.a(gate163inter10), .b(gate163inter9), .O(gate163inter11));
  nor2  gate1427(.a(gate163inter11), .b(gate163inter6), .O(gate163inter12));
  nand2 gate1428(.a(gate163inter12), .b(gate163inter1), .O(G580));

  xor2  gate2521(.a(G537), .b(G459), .O(gate164inter0));
  nand2 gate2522(.a(gate164inter0), .b(s_282), .O(gate164inter1));
  and2  gate2523(.a(G537), .b(G459), .O(gate164inter2));
  inv1  gate2524(.a(s_282), .O(gate164inter3));
  inv1  gate2525(.a(s_283), .O(gate164inter4));
  nand2 gate2526(.a(gate164inter4), .b(gate164inter3), .O(gate164inter5));
  nor2  gate2527(.a(gate164inter5), .b(gate164inter2), .O(gate164inter6));
  inv1  gate2528(.a(G459), .O(gate164inter7));
  inv1  gate2529(.a(G537), .O(gate164inter8));
  nand2 gate2530(.a(gate164inter8), .b(gate164inter7), .O(gate164inter9));
  nand2 gate2531(.a(s_283), .b(gate164inter3), .O(gate164inter10));
  nor2  gate2532(.a(gate164inter10), .b(gate164inter9), .O(gate164inter11));
  nor2  gate2533(.a(gate164inter11), .b(gate164inter6), .O(gate164inter12));
  nand2 gate2534(.a(gate164inter12), .b(gate164inter1), .O(G581));
nand2 gate165( .a(G462), .b(G540), .O(G582) );
nand2 gate166( .a(G465), .b(G540), .O(G583) );

  xor2  gate2199(.a(G543), .b(G468), .O(gate167inter0));
  nand2 gate2200(.a(gate167inter0), .b(s_236), .O(gate167inter1));
  and2  gate2201(.a(G543), .b(G468), .O(gate167inter2));
  inv1  gate2202(.a(s_236), .O(gate167inter3));
  inv1  gate2203(.a(s_237), .O(gate167inter4));
  nand2 gate2204(.a(gate167inter4), .b(gate167inter3), .O(gate167inter5));
  nor2  gate2205(.a(gate167inter5), .b(gate167inter2), .O(gate167inter6));
  inv1  gate2206(.a(G468), .O(gate167inter7));
  inv1  gate2207(.a(G543), .O(gate167inter8));
  nand2 gate2208(.a(gate167inter8), .b(gate167inter7), .O(gate167inter9));
  nand2 gate2209(.a(s_237), .b(gate167inter3), .O(gate167inter10));
  nor2  gate2210(.a(gate167inter10), .b(gate167inter9), .O(gate167inter11));
  nor2  gate2211(.a(gate167inter11), .b(gate167inter6), .O(gate167inter12));
  nand2 gate2212(.a(gate167inter12), .b(gate167inter1), .O(G584));

  xor2  gate1373(.a(G543), .b(G471), .O(gate168inter0));
  nand2 gate1374(.a(gate168inter0), .b(s_118), .O(gate168inter1));
  and2  gate1375(.a(G543), .b(G471), .O(gate168inter2));
  inv1  gate1376(.a(s_118), .O(gate168inter3));
  inv1  gate1377(.a(s_119), .O(gate168inter4));
  nand2 gate1378(.a(gate168inter4), .b(gate168inter3), .O(gate168inter5));
  nor2  gate1379(.a(gate168inter5), .b(gate168inter2), .O(gate168inter6));
  inv1  gate1380(.a(G471), .O(gate168inter7));
  inv1  gate1381(.a(G543), .O(gate168inter8));
  nand2 gate1382(.a(gate168inter8), .b(gate168inter7), .O(gate168inter9));
  nand2 gate1383(.a(s_119), .b(gate168inter3), .O(gate168inter10));
  nor2  gate1384(.a(gate168inter10), .b(gate168inter9), .O(gate168inter11));
  nor2  gate1385(.a(gate168inter11), .b(gate168inter6), .O(gate168inter12));
  nand2 gate1386(.a(gate168inter12), .b(gate168inter1), .O(G585));
nand2 gate169( .a(G474), .b(G546), .O(G586) );
nand2 gate170( .a(G477), .b(G546), .O(G587) );
nand2 gate171( .a(G480), .b(G549), .O(G588) );
nand2 gate172( .a(G483), .b(G549), .O(G589) );

  xor2  gate2661(.a(G552), .b(G486), .O(gate173inter0));
  nand2 gate2662(.a(gate173inter0), .b(s_302), .O(gate173inter1));
  and2  gate2663(.a(G552), .b(G486), .O(gate173inter2));
  inv1  gate2664(.a(s_302), .O(gate173inter3));
  inv1  gate2665(.a(s_303), .O(gate173inter4));
  nand2 gate2666(.a(gate173inter4), .b(gate173inter3), .O(gate173inter5));
  nor2  gate2667(.a(gate173inter5), .b(gate173inter2), .O(gate173inter6));
  inv1  gate2668(.a(G486), .O(gate173inter7));
  inv1  gate2669(.a(G552), .O(gate173inter8));
  nand2 gate2670(.a(gate173inter8), .b(gate173inter7), .O(gate173inter9));
  nand2 gate2671(.a(s_303), .b(gate173inter3), .O(gate173inter10));
  nor2  gate2672(.a(gate173inter10), .b(gate173inter9), .O(gate173inter11));
  nor2  gate2673(.a(gate173inter11), .b(gate173inter6), .O(gate173inter12));
  nand2 gate2674(.a(gate173inter12), .b(gate173inter1), .O(G590));

  xor2  gate2171(.a(G552), .b(G489), .O(gate174inter0));
  nand2 gate2172(.a(gate174inter0), .b(s_232), .O(gate174inter1));
  and2  gate2173(.a(G552), .b(G489), .O(gate174inter2));
  inv1  gate2174(.a(s_232), .O(gate174inter3));
  inv1  gate2175(.a(s_233), .O(gate174inter4));
  nand2 gate2176(.a(gate174inter4), .b(gate174inter3), .O(gate174inter5));
  nor2  gate2177(.a(gate174inter5), .b(gate174inter2), .O(gate174inter6));
  inv1  gate2178(.a(G489), .O(gate174inter7));
  inv1  gate2179(.a(G552), .O(gate174inter8));
  nand2 gate2180(.a(gate174inter8), .b(gate174inter7), .O(gate174inter9));
  nand2 gate2181(.a(s_233), .b(gate174inter3), .O(gate174inter10));
  nor2  gate2182(.a(gate174inter10), .b(gate174inter9), .O(gate174inter11));
  nor2  gate2183(.a(gate174inter11), .b(gate174inter6), .O(gate174inter12));
  nand2 gate2184(.a(gate174inter12), .b(gate174inter1), .O(G591));
nand2 gate175( .a(G492), .b(G555), .O(G592) );
nand2 gate176( .a(G495), .b(G555), .O(G593) );
nand2 gate177( .a(G498), .b(G558), .O(G594) );
nand2 gate178( .a(G501), .b(G558), .O(G595) );
nand2 gate179( .a(G504), .b(G561), .O(G596) );
nand2 gate180( .a(G507), .b(G561), .O(G597) );

  xor2  gate2563(.a(G564), .b(G510), .O(gate181inter0));
  nand2 gate2564(.a(gate181inter0), .b(s_288), .O(gate181inter1));
  and2  gate2565(.a(G564), .b(G510), .O(gate181inter2));
  inv1  gate2566(.a(s_288), .O(gate181inter3));
  inv1  gate2567(.a(s_289), .O(gate181inter4));
  nand2 gate2568(.a(gate181inter4), .b(gate181inter3), .O(gate181inter5));
  nor2  gate2569(.a(gate181inter5), .b(gate181inter2), .O(gate181inter6));
  inv1  gate2570(.a(G510), .O(gate181inter7));
  inv1  gate2571(.a(G564), .O(gate181inter8));
  nand2 gate2572(.a(gate181inter8), .b(gate181inter7), .O(gate181inter9));
  nand2 gate2573(.a(s_289), .b(gate181inter3), .O(gate181inter10));
  nor2  gate2574(.a(gate181inter10), .b(gate181inter9), .O(gate181inter11));
  nor2  gate2575(.a(gate181inter11), .b(gate181inter6), .O(gate181inter12));
  nand2 gate2576(.a(gate181inter12), .b(gate181inter1), .O(G598));
nand2 gate182( .a(G513), .b(G564), .O(G599) );
nand2 gate183( .a(G516), .b(G567), .O(G600) );
nand2 gate184( .a(G519), .b(G567), .O(G601) );

  xor2  gate1037(.a(G571), .b(G570), .O(gate185inter0));
  nand2 gate1038(.a(gate185inter0), .b(s_70), .O(gate185inter1));
  and2  gate1039(.a(G571), .b(G570), .O(gate185inter2));
  inv1  gate1040(.a(s_70), .O(gate185inter3));
  inv1  gate1041(.a(s_71), .O(gate185inter4));
  nand2 gate1042(.a(gate185inter4), .b(gate185inter3), .O(gate185inter5));
  nor2  gate1043(.a(gate185inter5), .b(gate185inter2), .O(gate185inter6));
  inv1  gate1044(.a(G570), .O(gate185inter7));
  inv1  gate1045(.a(G571), .O(gate185inter8));
  nand2 gate1046(.a(gate185inter8), .b(gate185inter7), .O(gate185inter9));
  nand2 gate1047(.a(s_71), .b(gate185inter3), .O(gate185inter10));
  nor2  gate1048(.a(gate185inter10), .b(gate185inter9), .O(gate185inter11));
  nor2  gate1049(.a(gate185inter11), .b(gate185inter6), .O(gate185inter12));
  nand2 gate1050(.a(gate185inter12), .b(gate185inter1), .O(G602));

  xor2  gate2297(.a(G573), .b(G572), .O(gate186inter0));
  nand2 gate2298(.a(gate186inter0), .b(s_250), .O(gate186inter1));
  and2  gate2299(.a(G573), .b(G572), .O(gate186inter2));
  inv1  gate2300(.a(s_250), .O(gate186inter3));
  inv1  gate2301(.a(s_251), .O(gate186inter4));
  nand2 gate2302(.a(gate186inter4), .b(gate186inter3), .O(gate186inter5));
  nor2  gate2303(.a(gate186inter5), .b(gate186inter2), .O(gate186inter6));
  inv1  gate2304(.a(G572), .O(gate186inter7));
  inv1  gate2305(.a(G573), .O(gate186inter8));
  nand2 gate2306(.a(gate186inter8), .b(gate186inter7), .O(gate186inter9));
  nand2 gate2307(.a(s_251), .b(gate186inter3), .O(gate186inter10));
  nor2  gate2308(.a(gate186inter10), .b(gate186inter9), .O(gate186inter11));
  nor2  gate2309(.a(gate186inter11), .b(gate186inter6), .O(gate186inter12));
  nand2 gate2310(.a(gate186inter12), .b(gate186inter1), .O(G607));
nand2 gate187( .a(G574), .b(G575), .O(G612) );

  xor2  gate1331(.a(G577), .b(G576), .O(gate188inter0));
  nand2 gate1332(.a(gate188inter0), .b(s_112), .O(gate188inter1));
  and2  gate1333(.a(G577), .b(G576), .O(gate188inter2));
  inv1  gate1334(.a(s_112), .O(gate188inter3));
  inv1  gate1335(.a(s_113), .O(gate188inter4));
  nand2 gate1336(.a(gate188inter4), .b(gate188inter3), .O(gate188inter5));
  nor2  gate1337(.a(gate188inter5), .b(gate188inter2), .O(gate188inter6));
  inv1  gate1338(.a(G576), .O(gate188inter7));
  inv1  gate1339(.a(G577), .O(gate188inter8));
  nand2 gate1340(.a(gate188inter8), .b(gate188inter7), .O(gate188inter9));
  nand2 gate1341(.a(s_113), .b(gate188inter3), .O(gate188inter10));
  nor2  gate1342(.a(gate188inter10), .b(gate188inter9), .O(gate188inter11));
  nor2  gate1343(.a(gate188inter11), .b(gate188inter6), .O(gate188inter12));
  nand2 gate1344(.a(gate188inter12), .b(gate188inter1), .O(G617));

  xor2  gate2185(.a(G579), .b(G578), .O(gate189inter0));
  nand2 gate2186(.a(gate189inter0), .b(s_234), .O(gate189inter1));
  and2  gate2187(.a(G579), .b(G578), .O(gate189inter2));
  inv1  gate2188(.a(s_234), .O(gate189inter3));
  inv1  gate2189(.a(s_235), .O(gate189inter4));
  nand2 gate2190(.a(gate189inter4), .b(gate189inter3), .O(gate189inter5));
  nor2  gate2191(.a(gate189inter5), .b(gate189inter2), .O(gate189inter6));
  inv1  gate2192(.a(G578), .O(gate189inter7));
  inv1  gate2193(.a(G579), .O(gate189inter8));
  nand2 gate2194(.a(gate189inter8), .b(gate189inter7), .O(gate189inter9));
  nand2 gate2195(.a(s_235), .b(gate189inter3), .O(gate189inter10));
  nor2  gate2196(.a(gate189inter10), .b(gate189inter9), .O(gate189inter11));
  nor2  gate2197(.a(gate189inter11), .b(gate189inter6), .O(gate189inter12));
  nand2 gate2198(.a(gate189inter12), .b(gate189inter1), .O(G622));
nand2 gate190( .a(G580), .b(G581), .O(G627) );

  xor2  gate1191(.a(G583), .b(G582), .O(gate191inter0));
  nand2 gate1192(.a(gate191inter0), .b(s_92), .O(gate191inter1));
  and2  gate1193(.a(G583), .b(G582), .O(gate191inter2));
  inv1  gate1194(.a(s_92), .O(gate191inter3));
  inv1  gate1195(.a(s_93), .O(gate191inter4));
  nand2 gate1196(.a(gate191inter4), .b(gate191inter3), .O(gate191inter5));
  nor2  gate1197(.a(gate191inter5), .b(gate191inter2), .O(gate191inter6));
  inv1  gate1198(.a(G582), .O(gate191inter7));
  inv1  gate1199(.a(G583), .O(gate191inter8));
  nand2 gate1200(.a(gate191inter8), .b(gate191inter7), .O(gate191inter9));
  nand2 gate1201(.a(s_93), .b(gate191inter3), .O(gate191inter10));
  nor2  gate1202(.a(gate191inter10), .b(gate191inter9), .O(gate191inter11));
  nor2  gate1203(.a(gate191inter11), .b(gate191inter6), .O(gate191inter12));
  nand2 gate1204(.a(gate191inter12), .b(gate191inter1), .O(G632));

  xor2  gate2647(.a(G585), .b(G584), .O(gate192inter0));
  nand2 gate2648(.a(gate192inter0), .b(s_300), .O(gate192inter1));
  and2  gate2649(.a(G585), .b(G584), .O(gate192inter2));
  inv1  gate2650(.a(s_300), .O(gate192inter3));
  inv1  gate2651(.a(s_301), .O(gate192inter4));
  nand2 gate2652(.a(gate192inter4), .b(gate192inter3), .O(gate192inter5));
  nor2  gate2653(.a(gate192inter5), .b(gate192inter2), .O(gate192inter6));
  inv1  gate2654(.a(G584), .O(gate192inter7));
  inv1  gate2655(.a(G585), .O(gate192inter8));
  nand2 gate2656(.a(gate192inter8), .b(gate192inter7), .O(gate192inter9));
  nand2 gate2657(.a(s_301), .b(gate192inter3), .O(gate192inter10));
  nor2  gate2658(.a(gate192inter10), .b(gate192inter9), .O(gate192inter11));
  nor2  gate2659(.a(gate192inter11), .b(gate192inter6), .O(gate192inter12));
  nand2 gate2660(.a(gate192inter12), .b(gate192inter1), .O(G637));

  xor2  gate2815(.a(G587), .b(G586), .O(gate193inter0));
  nand2 gate2816(.a(gate193inter0), .b(s_324), .O(gate193inter1));
  and2  gate2817(.a(G587), .b(G586), .O(gate193inter2));
  inv1  gate2818(.a(s_324), .O(gate193inter3));
  inv1  gate2819(.a(s_325), .O(gate193inter4));
  nand2 gate2820(.a(gate193inter4), .b(gate193inter3), .O(gate193inter5));
  nor2  gate2821(.a(gate193inter5), .b(gate193inter2), .O(gate193inter6));
  inv1  gate2822(.a(G586), .O(gate193inter7));
  inv1  gate2823(.a(G587), .O(gate193inter8));
  nand2 gate2824(.a(gate193inter8), .b(gate193inter7), .O(gate193inter9));
  nand2 gate2825(.a(s_325), .b(gate193inter3), .O(gate193inter10));
  nor2  gate2826(.a(gate193inter10), .b(gate193inter9), .O(gate193inter11));
  nor2  gate2827(.a(gate193inter11), .b(gate193inter6), .O(gate193inter12));
  nand2 gate2828(.a(gate193inter12), .b(gate193inter1), .O(G642));
nand2 gate194( .a(G588), .b(G589), .O(G645) );
nand2 gate195( .a(G590), .b(G591), .O(G648) );
nand2 gate196( .a(G592), .b(G593), .O(G651) );
nand2 gate197( .a(G594), .b(G595), .O(G654) );
nand2 gate198( .a(G596), .b(G597), .O(G657) );

  xor2  gate1009(.a(G599), .b(G598), .O(gate199inter0));
  nand2 gate1010(.a(gate199inter0), .b(s_66), .O(gate199inter1));
  and2  gate1011(.a(G599), .b(G598), .O(gate199inter2));
  inv1  gate1012(.a(s_66), .O(gate199inter3));
  inv1  gate1013(.a(s_67), .O(gate199inter4));
  nand2 gate1014(.a(gate199inter4), .b(gate199inter3), .O(gate199inter5));
  nor2  gate1015(.a(gate199inter5), .b(gate199inter2), .O(gate199inter6));
  inv1  gate1016(.a(G598), .O(gate199inter7));
  inv1  gate1017(.a(G599), .O(gate199inter8));
  nand2 gate1018(.a(gate199inter8), .b(gate199inter7), .O(gate199inter9));
  nand2 gate1019(.a(s_67), .b(gate199inter3), .O(gate199inter10));
  nor2  gate1020(.a(gate199inter10), .b(gate199inter9), .O(gate199inter11));
  nor2  gate1021(.a(gate199inter11), .b(gate199inter6), .O(gate199inter12));
  nand2 gate1022(.a(gate199inter12), .b(gate199inter1), .O(G660));
nand2 gate200( .a(G600), .b(G601), .O(G663) );

  xor2  gate2759(.a(G607), .b(G602), .O(gate201inter0));
  nand2 gate2760(.a(gate201inter0), .b(s_316), .O(gate201inter1));
  and2  gate2761(.a(G607), .b(G602), .O(gate201inter2));
  inv1  gate2762(.a(s_316), .O(gate201inter3));
  inv1  gate2763(.a(s_317), .O(gate201inter4));
  nand2 gate2764(.a(gate201inter4), .b(gate201inter3), .O(gate201inter5));
  nor2  gate2765(.a(gate201inter5), .b(gate201inter2), .O(gate201inter6));
  inv1  gate2766(.a(G602), .O(gate201inter7));
  inv1  gate2767(.a(G607), .O(gate201inter8));
  nand2 gate2768(.a(gate201inter8), .b(gate201inter7), .O(gate201inter9));
  nand2 gate2769(.a(s_317), .b(gate201inter3), .O(gate201inter10));
  nor2  gate2770(.a(gate201inter10), .b(gate201inter9), .O(gate201inter11));
  nor2  gate2771(.a(gate201inter11), .b(gate201inter6), .O(gate201inter12));
  nand2 gate2772(.a(gate201inter12), .b(gate201inter1), .O(G666));
nand2 gate202( .a(G612), .b(G617), .O(G669) );
nand2 gate203( .a(G602), .b(G612), .O(G672) );
nand2 gate204( .a(G607), .b(G617), .O(G675) );
nand2 gate205( .a(G622), .b(G627), .O(G678) );
nand2 gate206( .a(G632), .b(G637), .O(G681) );

  xor2  gate855(.a(G632), .b(G622), .O(gate207inter0));
  nand2 gate856(.a(gate207inter0), .b(s_44), .O(gate207inter1));
  and2  gate857(.a(G632), .b(G622), .O(gate207inter2));
  inv1  gate858(.a(s_44), .O(gate207inter3));
  inv1  gate859(.a(s_45), .O(gate207inter4));
  nand2 gate860(.a(gate207inter4), .b(gate207inter3), .O(gate207inter5));
  nor2  gate861(.a(gate207inter5), .b(gate207inter2), .O(gate207inter6));
  inv1  gate862(.a(G622), .O(gate207inter7));
  inv1  gate863(.a(G632), .O(gate207inter8));
  nand2 gate864(.a(gate207inter8), .b(gate207inter7), .O(gate207inter9));
  nand2 gate865(.a(s_45), .b(gate207inter3), .O(gate207inter10));
  nor2  gate866(.a(gate207inter10), .b(gate207inter9), .O(gate207inter11));
  nor2  gate867(.a(gate207inter11), .b(gate207inter6), .O(gate207inter12));
  nand2 gate868(.a(gate207inter12), .b(gate207inter1), .O(G684));
nand2 gate208( .a(G627), .b(G637), .O(G687) );

  xor2  gate2451(.a(G666), .b(G602), .O(gate209inter0));
  nand2 gate2452(.a(gate209inter0), .b(s_272), .O(gate209inter1));
  and2  gate2453(.a(G666), .b(G602), .O(gate209inter2));
  inv1  gate2454(.a(s_272), .O(gate209inter3));
  inv1  gate2455(.a(s_273), .O(gate209inter4));
  nand2 gate2456(.a(gate209inter4), .b(gate209inter3), .O(gate209inter5));
  nor2  gate2457(.a(gate209inter5), .b(gate209inter2), .O(gate209inter6));
  inv1  gate2458(.a(G602), .O(gate209inter7));
  inv1  gate2459(.a(G666), .O(gate209inter8));
  nand2 gate2460(.a(gate209inter8), .b(gate209inter7), .O(gate209inter9));
  nand2 gate2461(.a(s_273), .b(gate209inter3), .O(gate209inter10));
  nor2  gate2462(.a(gate209inter10), .b(gate209inter9), .O(gate209inter11));
  nor2  gate2463(.a(gate209inter11), .b(gate209inter6), .O(gate209inter12));
  nand2 gate2464(.a(gate209inter12), .b(gate209inter1), .O(G690));
nand2 gate210( .a(G607), .b(G666), .O(G691) );
nand2 gate211( .a(G612), .b(G669), .O(G692) );
nand2 gate212( .a(G617), .b(G669), .O(G693) );

  xor2  gate2017(.a(G672), .b(G602), .O(gate213inter0));
  nand2 gate2018(.a(gate213inter0), .b(s_210), .O(gate213inter1));
  and2  gate2019(.a(G672), .b(G602), .O(gate213inter2));
  inv1  gate2020(.a(s_210), .O(gate213inter3));
  inv1  gate2021(.a(s_211), .O(gate213inter4));
  nand2 gate2022(.a(gate213inter4), .b(gate213inter3), .O(gate213inter5));
  nor2  gate2023(.a(gate213inter5), .b(gate213inter2), .O(gate213inter6));
  inv1  gate2024(.a(G602), .O(gate213inter7));
  inv1  gate2025(.a(G672), .O(gate213inter8));
  nand2 gate2026(.a(gate213inter8), .b(gate213inter7), .O(gate213inter9));
  nand2 gate2027(.a(s_211), .b(gate213inter3), .O(gate213inter10));
  nor2  gate2028(.a(gate213inter10), .b(gate213inter9), .O(gate213inter11));
  nor2  gate2029(.a(gate213inter11), .b(gate213inter6), .O(gate213inter12));
  nand2 gate2030(.a(gate213inter12), .b(gate213inter1), .O(G694));

  xor2  gate2157(.a(G672), .b(G612), .O(gate214inter0));
  nand2 gate2158(.a(gate214inter0), .b(s_230), .O(gate214inter1));
  and2  gate2159(.a(G672), .b(G612), .O(gate214inter2));
  inv1  gate2160(.a(s_230), .O(gate214inter3));
  inv1  gate2161(.a(s_231), .O(gate214inter4));
  nand2 gate2162(.a(gate214inter4), .b(gate214inter3), .O(gate214inter5));
  nor2  gate2163(.a(gate214inter5), .b(gate214inter2), .O(gate214inter6));
  inv1  gate2164(.a(G612), .O(gate214inter7));
  inv1  gate2165(.a(G672), .O(gate214inter8));
  nand2 gate2166(.a(gate214inter8), .b(gate214inter7), .O(gate214inter9));
  nand2 gate2167(.a(s_231), .b(gate214inter3), .O(gate214inter10));
  nor2  gate2168(.a(gate214inter10), .b(gate214inter9), .O(gate214inter11));
  nor2  gate2169(.a(gate214inter11), .b(gate214inter6), .O(gate214inter12));
  nand2 gate2170(.a(gate214inter12), .b(gate214inter1), .O(G695));
nand2 gate215( .a(G607), .b(G675), .O(G696) );

  xor2  gate2493(.a(G675), .b(G617), .O(gate216inter0));
  nand2 gate2494(.a(gate216inter0), .b(s_278), .O(gate216inter1));
  and2  gate2495(.a(G675), .b(G617), .O(gate216inter2));
  inv1  gate2496(.a(s_278), .O(gate216inter3));
  inv1  gate2497(.a(s_279), .O(gate216inter4));
  nand2 gate2498(.a(gate216inter4), .b(gate216inter3), .O(gate216inter5));
  nor2  gate2499(.a(gate216inter5), .b(gate216inter2), .O(gate216inter6));
  inv1  gate2500(.a(G617), .O(gate216inter7));
  inv1  gate2501(.a(G675), .O(gate216inter8));
  nand2 gate2502(.a(gate216inter8), .b(gate216inter7), .O(gate216inter9));
  nand2 gate2503(.a(s_279), .b(gate216inter3), .O(gate216inter10));
  nor2  gate2504(.a(gate216inter10), .b(gate216inter9), .O(gate216inter11));
  nor2  gate2505(.a(gate216inter11), .b(gate216inter6), .O(gate216inter12));
  nand2 gate2506(.a(gate216inter12), .b(gate216inter1), .O(G697));

  xor2  gate2031(.a(G678), .b(G622), .O(gate217inter0));
  nand2 gate2032(.a(gate217inter0), .b(s_212), .O(gate217inter1));
  and2  gate2033(.a(G678), .b(G622), .O(gate217inter2));
  inv1  gate2034(.a(s_212), .O(gate217inter3));
  inv1  gate2035(.a(s_213), .O(gate217inter4));
  nand2 gate2036(.a(gate217inter4), .b(gate217inter3), .O(gate217inter5));
  nor2  gate2037(.a(gate217inter5), .b(gate217inter2), .O(gate217inter6));
  inv1  gate2038(.a(G622), .O(gate217inter7));
  inv1  gate2039(.a(G678), .O(gate217inter8));
  nand2 gate2040(.a(gate217inter8), .b(gate217inter7), .O(gate217inter9));
  nand2 gate2041(.a(s_213), .b(gate217inter3), .O(gate217inter10));
  nor2  gate2042(.a(gate217inter10), .b(gate217inter9), .O(gate217inter11));
  nor2  gate2043(.a(gate217inter11), .b(gate217inter6), .O(gate217inter12));
  nand2 gate2044(.a(gate217inter12), .b(gate217inter1), .O(G698));
nand2 gate218( .a(G627), .b(G678), .O(G699) );
nand2 gate219( .a(G632), .b(G681), .O(G700) );
nand2 gate220( .a(G637), .b(G681), .O(G701) );
nand2 gate221( .a(G622), .b(G684), .O(G702) );
nand2 gate222( .a(G632), .b(G684), .O(G703) );

  xor2  gate1065(.a(G687), .b(G627), .O(gate223inter0));
  nand2 gate1066(.a(gate223inter0), .b(s_74), .O(gate223inter1));
  and2  gate1067(.a(G687), .b(G627), .O(gate223inter2));
  inv1  gate1068(.a(s_74), .O(gate223inter3));
  inv1  gate1069(.a(s_75), .O(gate223inter4));
  nand2 gate1070(.a(gate223inter4), .b(gate223inter3), .O(gate223inter5));
  nor2  gate1071(.a(gate223inter5), .b(gate223inter2), .O(gate223inter6));
  inv1  gate1072(.a(G627), .O(gate223inter7));
  inv1  gate1073(.a(G687), .O(gate223inter8));
  nand2 gate1074(.a(gate223inter8), .b(gate223inter7), .O(gate223inter9));
  nand2 gate1075(.a(s_75), .b(gate223inter3), .O(gate223inter10));
  nor2  gate1076(.a(gate223inter10), .b(gate223inter9), .O(gate223inter11));
  nor2  gate1077(.a(gate223inter11), .b(gate223inter6), .O(gate223inter12));
  nand2 gate1078(.a(gate223inter12), .b(gate223inter1), .O(G704));
nand2 gate224( .a(G637), .b(G687), .O(G705) );

  xor2  gate1261(.a(G691), .b(G690), .O(gate225inter0));
  nand2 gate1262(.a(gate225inter0), .b(s_102), .O(gate225inter1));
  and2  gate1263(.a(G691), .b(G690), .O(gate225inter2));
  inv1  gate1264(.a(s_102), .O(gate225inter3));
  inv1  gate1265(.a(s_103), .O(gate225inter4));
  nand2 gate1266(.a(gate225inter4), .b(gate225inter3), .O(gate225inter5));
  nor2  gate1267(.a(gate225inter5), .b(gate225inter2), .O(gate225inter6));
  inv1  gate1268(.a(G690), .O(gate225inter7));
  inv1  gate1269(.a(G691), .O(gate225inter8));
  nand2 gate1270(.a(gate225inter8), .b(gate225inter7), .O(gate225inter9));
  nand2 gate1271(.a(s_103), .b(gate225inter3), .O(gate225inter10));
  nor2  gate1272(.a(gate225inter10), .b(gate225inter9), .O(gate225inter11));
  nor2  gate1273(.a(gate225inter11), .b(gate225inter6), .O(gate225inter12));
  nand2 gate1274(.a(gate225inter12), .b(gate225inter1), .O(G706));

  xor2  gate645(.a(G693), .b(G692), .O(gate226inter0));
  nand2 gate646(.a(gate226inter0), .b(s_14), .O(gate226inter1));
  and2  gate647(.a(G693), .b(G692), .O(gate226inter2));
  inv1  gate648(.a(s_14), .O(gate226inter3));
  inv1  gate649(.a(s_15), .O(gate226inter4));
  nand2 gate650(.a(gate226inter4), .b(gate226inter3), .O(gate226inter5));
  nor2  gate651(.a(gate226inter5), .b(gate226inter2), .O(gate226inter6));
  inv1  gate652(.a(G692), .O(gate226inter7));
  inv1  gate653(.a(G693), .O(gate226inter8));
  nand2 gate654(.a(gate226inter8), .b(gate226inter7), .O(gate226inter9));
  nand2 gate655(.a(s_15), .b(gate226inter3), .O(gate226inter10));
  nor2  gate656(.a(gate226inter10), .b(gate226inter9), .O(gate226inter11));
  nor2  gate657(.a(gate226inter11), .b(gate226inter6), .O(gate226inter12));
  nand2 gate658(.a(gate226inter12), .b(gate226inter1), .O(G709));
nand2 gate227( .a(G694), .b(G695), .O(G712) );
nand2 gate228( .a(G696), .b(G697), .O(G715) );

  xor2  gate2255(.a(G699), .b(G698), .O(gate229inter0));
  nand2 gate2256(.a(gate229inter0), .b(s_244), .O(gate229inter1));
  and2  gate2257(.a(G699), .b(G698), .O(gate229inter2));
  inv1  gate2258(.a(s_244), .O(gate229inter3));
  inv1  gate2259(.a(s_245), .O(gate229inter4));
  nand2 gate2260(.a(gate229inter4), .b(gate229inter3), .O(gate229inter5));
  nor2  gate2261(.a(gate229inter5), .b(gate229inter2), .O(gate229inter6));
  inv1  gate2262(.a(G698), .O(gate229inter7));
  inv1  gate2263(.a(G699), .O(gate229inter8));
  nand2 gate2264(.a(gate229inter8), .b(gate229inter7), .O(gate229inter9));
  nand2 gate2265(.a(s_245), .b(gate229inter3), .O(gate229inter10));
  nor2  gate2266(.a(gate229inter10), .b(gate229inter9), .O(gate229inter11));
  nor2  gate2267(.a(gate229inter11), .b(gate229inter6), .O(gate229inter12));
  nand2 gate2268(.a(gate229inter12), .b(gate229inter1), .O(G718));

  xor2  gate1849(.a(G701), .b(G700), .O(gate230inter0));
  nand2 gate1850(.a(gate230inter0), .b(s_186), .O(gate230inter1));
  and2  gate1851(.a(G701), .b(G700), .O(gate230inter2));
  inv1  gate1852(.a(s_186), .O(gate230inter3));
  inv1  gate1853(.a(s_187), .O(gate230inter4));
  nand2 gate1854(.a(gate230inter4), .b(gate230inter3), .O(gate230inter5));
  nor2  gate1855(.a(gate230inter5), .b(gate230inter2), .O(gate230inter6));
  inv1  gate1856(.a(G700), .O(gate230inter7));
  inv1  gate1857(.a(G701), .O(gate230inter8));
  nand2 gate1858(.a(gate230inter8), .b(gate230inter7), .O(gate230inter9));
  nand2 gate1859(.a(s_187), .b(gate230inter3), .O(gate230inter10));
  nor2  gate1860(.a(gate230inter10), .b(gate230inter9), .O(gate230inter11));
  nor2  gate1861(.a(gate230inter11), .b(gate230inter6), .O(gate230inter12));
  nand2 gate1862(.a(gate230inter12), .b(gate230inter1), .O(G721));
nand2 gate231( .a(G702), .b(G703), .O(G724) );
nand2 gate232( .a(G704), .b(G705), .O(G727) );

  xor2  gate2913(.a(G718), .b(G242), .O(gate233inter0));
  nand2 gate2914(.a(gate233inter0), .b(s_338), .O(gate233inter1));
  and2  gate2915(.a(G718), .b(G242), .O(gate233inter2));
  inv1  gate2916(.a(s_338), .O(gate233inter3));
  inv1  gate2917(.a(s_339), .O(gate233inter4));
  nand2 gate2918(.a(gate233inter4), .b(gate233inter3), .O(gate233inter5));
  nor2  gate2919(.a(gate233inter5), .b(gate233inter2), .O(gate233inter6));
  inv1  gate2920(.a(G242), .O(gate233inter7));
  inv1  gate2921(.a(G718), .O(gate233inter8));
  nand2 gate2922(.a(gate233inter8), .b(gate233inter7), .O(gate233inter9));
  nand2 gate2923(.a(s_339), .b(gate233inter3), .O(gate233inter10));
  nor2  gate2924(.a(gate233inter10), .b(gate233inter9), .O(gate233inter11));
  nor2  gate2925(.a(gate233inter11), .b(gate233inter6), .O(gate233inter12));
  nand2 gate2926(.a(gate233inter12), .b(gate233inter1), .O(G730));
nand2 gate234( .a(G245), .b(G721), .O(G733) );

  xor2  gate1737(.a(G724), .b(G248), .O(gate235inter0));
  nand2 gate1738(.a(gate235inter0), .b(s_170), .O(gate235inter1));
  and2  gate1739(.a(G724), .b(G248), .O(gate235inter2));
  inv1  gate1740(.a(s_170), .O(gate235inter3));
  inv1  gate1741(.a(s_171), .O(gate235inter4));
  nand2 gate1742(.a(gate235inter4), .b(gate235inter3), .O(gate235inter5));
  nor2  gate1743(.a(gate235inter5), .b(gate235inter2), .O(gate235inter6));
  inv1  gate1744(.a(G248), .O(gate235inter7));
  inv1  gate1745(.a(G724), .O(gate235inter8));
  nand2 gate1746(.a(gate235inter8), .b(gate235inter7), .O(gate235inter9));
  nand2 gate1747(.a(s_171), .b(gate235inter3), .O(gate235inter10));
  nor2  gate1748(.a(gate235inter10), .b(gate235inter9), .O(gate235inter11));
  nor2  gate1749(.a(gate235inter11), .b(gate235inter6), .O(gate235inter12));
  nand2 gate1750(.a(gate235inter12), .b(gate235inter1), .O(G736));

  xor2  gate2437(.a(G727), .b(G251), .O(gate236inter0));
  nand2 gate2438(.a(gate236inter0), .b(s_270), .O(gate236inter1));
  and2  gate2439(.a(G727), .b(G251), .O(gate236inter2));
  inv1  gate2440(.a(s_270), .O(gate236inter3));
  inv1  gate2441(.a(s_271), .O(gate236inter4));
  nand2 gate2442(.a(gate236inter4), .b(gate236inter3), .O(gate236inter5));
  nor2  gate2443(.a(gate236inter5), .b(gate236inter2), .O(gate236inter6));
  inv1  gate2444(.a(G251), .O(gate236inter7));
  inv1  gate2445(.a(G727), .O(gate236inter8));
  nand2 gate2446(.a(gate236inter8), .b(gate236inter7), .O(gate236inter9));
  nand2 gate2447(.a(s_271), .b(gate236inter3), .O(gate236inter10));
  nor2  gate2448(.a(gate236inter10), .b(gate236inter9), .O(gate236inter11));
  nor2  gate2449(.a(gate236inter11), .b(gate236inter6), .O(gate236inter12));
  nand2 gate2450(.a(gate236inter12), .b(gate236inter1), .O(G739));
nand2 gate237( .a(G254), .b(G706), .O(G742) );

  xor2  gate1723(.a(G709), .b(G257), .O(gate238inter0));
  nand2 gate1724(.a(gate238inter0), .b(s_168), .O(gate238inter1));
  and2  gate1725(.a(G709), .b(G257), .O(gate238inter2));
  inv1  gate1726(.a(s_168), .O(gate238inter3));
  inv1  gate1727(.a(s_169), .O(gate238inter4));
  nand2 gate1728(.a(gate238inter4), .b(gate238inter3), .O(gate238inter5));
  nor2  gate1729(.a(gate238inter5), .b(gate238inter2), .O(gate238inter6));
  inv1  gate1730(.a(G257), .O(gate238inter7));
  inv1  gate1731(.a(G709), .O(gate238inter8));
  nand2 gate1732(.a(gate238inter8), .b(gate238inter7), .O(gate238inter9));
  nand2 gate1733(.a(s_169), .b(gate238inter3), .O(gate238inter10));
  nor2  gate1734(.a(gate238inter10), .b(gate238inter9), .O(gate238inter11));
  nor2  gate1735(.a(gate238inter11), .b(gate238inter6), .O(gate238inter12));
  nand2 gate1736(.a(gate238inter12), .b(gate238inter1), .O(G745));

  xor2  gate673(.a(G712), .b(G260), .O(gate239inter0));
  nand2 gate674(.a(gate239inter0), .b(s_18), .O(gate239inter1));
  and2  gate675(.a(G712), .b(G260), .O(gate239inter2));
  inv1  gate676(.a(s_18), .O(gate239inter3));
  inv1  gate677(.a(s_19), .O(gate239inter4));
  nand2 gate678(.a(gate239inter4), .b(gate239inter3), .O(gate239inter5));
  nor2  gate679(.a(gate239inter5), .b(gate239inter2), .O(gate239inter6));
  inv1  gate680(.a(G260), .O(gate239inter7));
  inv1  gate681(.a(G712), .O(gate239inter8));
  nand2 gate682(.a(gate239inter8), .b(gate239inter7), .O(gate239inter9));
  nand2 gate683(.a(s_19), .b(gate239inter3), .O(gate239inter10));
  nor2  gate684(.a(gate239inter10), .b(gate239inter9), .O(gate239inter11));
  nor2  gate685(.a(gate239inter11), .b(gate239inter6), .O(gate239inter12));
  nand2 gate686(.a(gate239inter12), .b(gate239inter1), .O(G748));

  xor2  gate1471(.a(G715), .b(G263), .O(gate240inter0));
  nand2 gate1472(.a(gate240inter0), .b(s_132), .O(gate240inter1));
  and2  gate1473(.a(G715), .b(G263), .O(gate240inter2));
  inv1  gate1474(.a(s_132), .O(gate240inter3));
  inv1  gate1475(.a(s_133), .O(gate240inter4));
  nand2 gate1476(.a(gate240inter4), .b(gate240inter3), .O(gate240inter5));
  nor2  gate1477(.a(gate240inter5), .b(gate240inter2), .O(gate240inter6));
  inv1  gate1478(.a(G263), .O(gate240inter7));
  inv1  gate1479(.a(G715), .O(gate240inter8));
  nand2 gate1480(.a(gate240inter8), .b(gate240inter7), .O(gate240inter9));
  nand2 gate1481(.a(s_133), .b(gate240inter3), .O(gate240inter10));
  nor2  gate1482(.a(gate240inter10), .b(gate240inter9), .O(gate240inter11));
  nor2  gate1483(.a(gate240inter11), .b(gate240inter6), .O(gate240inter12));
  nand2 gate1484(.a(gate240inter12), .b(gate240inter1), .O(G751));
nand2 gate241( .a(G242), .b(G730), .O(G754) );
nand2 gate242( .a(G718), .b(G730), .O(G755) );
nand2 gate243( .a(G245), .b(G733), .O(G756) );

  xor2  gate2465(.a(G733), .b(G721), .O(gate244inter0));
  nand2 gate2466(.a(gate244inter0), .b(s_274), .O(gate244inter1));
  and2  gate2467(.a(G733), .b(G721), .O(gate244inter2));
  inv1  gate2468(.a(s_274), .O(gate244inter3));
  inv1  gate2469(.a(s_275), .O(gate244inter4));
  nand2 gate2470(.a(gate244inter4), .b(gate244inter3), .O(gate244inter5));
  nor2  gate2471(.a(gate244inter5), .b(gate244inter2), .O(gate244inter6));
  inv1  gate2472(.a(G721), .O(gate244inter7));
  inv1  gate2473(.a(G733), .O(gate244inter8));
  nand2 gate2474(.a(gate244inter8), .b(gate244inter7), .O(gate244inter9));
  nand2 gate2475(.a(s_275), .b(gate244inter3), .O(gate244inter10));
  nor2  gate2476(.a(gate244inter10), .b(gate244inter9), .O(gate244inter11));
  nor2  gate2477(.a(gate244inter11), .b(gate244inter6), .O(gate244inter12));
  nand2 gate2478(.a(gate244inter12), .b(gate244inter1), .O(G757));
nand2 gate245( .a(G248), .b(G736), .O(G758) );
nand2 gate246( .a(G724), .b(G736), .O(G759) );

  xor2  gate3039(.a(G739), .b(G251), .O(gate247inter0));
  nand2 gate3040(.a(gate247inter0), .b(s_356), .O(gate247inter1));
  and2  gate3041(.a(G739), .b(G251), .O(gate247inter2));
  inv1  gate3042(.a(s_356), .O(gate247inter3));
  inv1  gate3043(.a(s_357), .O(gate247inter4));
  nand2 gate3044(.a(gate247inter4), .b(gate247inter3), .O(gate247inter5));
  nor2  gate3045(.a(gate247inter5), .b(gate247inter2), .O(gate247inter6));
  inv1  gate3046(.a(G251), .O(gate247inter7));
  inv1  gate3047(.a(G739), .O(gate247inter8));
  nand2 gate3048(.a(gate247inter8), .b(gate247inter7), .O(gate247inter9));
  nand2 gate3049(.a(s_357), .b(gate247inter3), .O(gate247inter10));
  nor2  gate3050(.a(gate247inter10), .b(gate247inter9), .O(gate247inter11));
  nor2  gate3051(.a(gate247inter11), .b(gate247inter6), .O(gate247inter12));
  nand2 gate3052(.a(gate247inter12), .b(gate247inter1), .O(G760));

  xor2  gate1233(.a(G739), .b(G727), .O(gate248inter0));
  nand2 gate1234(.a(gate248inter0), .b(s_98), .O(gate248inter1));
  and2  gate1235(.a(G739), .b(G727), .O(gate248inter2));
  inv1  gate1236(.a(s_98), .O(gate248inter3));
  inv1  gate1237(.a(s_99), .O(gate248inter4));
  nand2 gate1238(.a(gate248inter4), .b(gate248inter3), .O(gate248inter5));
  nor2  gate1239(.a(gate248inter5), .b(gate248inter2), .O(gate248inter6));
  inv1  gate1240(.a(G727), .O(gate248inter7));
  inv1  gate1241(.a(G739), .O(gate248inter8));
  nand2 gate1242(.a(gate248inter8), .b(gate248inter7), .O(gate248inter9));
  nand2 gate1243(.a(s_99), .b(gate248inter3), .O(gate248inter10));
  nor2  gate1244(.a(gate248inter10), .b(gate248inter9), .O(gate248inter11));
  nor2  gate1245(.a(gate248inter11), .b(gate248inter6), .O(gate248inter12));
  nand2 gate1246(.a(gate248inter12), .b(gate248inter1), .O(G761));
nand2 gate249( .a(G254), .b(G742), .O(G762) );

  xor2  gate659(.a(G742), .b(G706), .O(gate250inter0));
  nand2 gate660(.a(gate250inter0), .b(s_16), .O(gate250inter1));
  and2  gate661(.a(G742), .b(G706), .O(gate250inter2));
  inv1  gate662(.a(s_16), .O(gate250inter3));
  inv1  gate663(.a(s_17), .O(gate250inter4));
  nand2 gate664(.a(gate250inter4), .b(gate250inter3), .O(gate250inter5));
  nor2  gate665(.a(gate250inter5), .b(gate250inter2), .O(gate250inter6));
  inv1  gate666(.a(G706), .O(gate250inter7));
  inv1  gate667(.a(G742), .O(gate250inter8));
  nand2 gate668(.a(gate250inter8), .b(gate250inter7), .O(gate250inter9));
  nand2 gate669(.a(s_17), .b(gate250inter3), .O(gate250inter10));
  nor2  gate670(.a(gate250inter10), .b(gate250inter9), .O(gate250inter11));
  nor2  gate671(.a(gate250inter11), .b(gate250inter6), .O(gate250inter12));
  nand2 gate672(.a(gate250inter12), .b(gate250inter1), .O(G763));

  xor2  gate1751(.a(G745), .b(G257), .O(gate251inter0));
  nand2 gate1752(.a(gate251inter0), .b(s_172), .O(gate251inter1));
  and2  gate1753(.a(G745), .b(G257), .O(gate251inter2));
  inv1  gate1754(.a(s_172), .O(gate251inter3));
  inv1  gate1755(.a(s_173), .O(gate251inter4));
  nand2 gate1756(.a(gate251inter4), .b(gate251inter3), .O(gate251inter5));
  nor2  gate1757(.a(gate251inter5), .b(gate251inter2), .O(gate251inter6));
  inv1  gate1758(.a(G257), .O(gate251inter7));
  inv1  gate1759(.a(G745), .O(gate251inter8));
  nand2 gate1760(.a(gate251inter8), .b(gate251inter7), .O(gate251inter9));
  nand2 gate1761(.a(s_173), .b(gate251inter3), .O(gate251inter10));
  nor2  gate1762(.a(gate251inter10), .b(gate251inter9), .O(gate251inter11));
  nor2  gate1763(.a(gate251inter11), .b(gate251inter6), .O(gate251inter12));
  nand2 gate1764(.a(gate251inter12), .b(gate251inter1), .O(G764));

  xor2  gate813(.a(G745), .b(G709), .O(gate252inter0));
  nand2 gate814(.a(gate252inter0), .b(s_38), .O(gate252inter1));
  and2  gate815(.a(G745), .b(G709), .O(gate252inter2));
  inv1  gate816(.a(s_38), .O(gate252inter3));
  inv1  gate817(.a(s_39), .O(gate252inter4));
  nand2 gate818(.a(gate252inter4), .b(gate252inter3), .O(gate252inter5));
  nor2  gate819(.a(gate252inter5), .b(gate252inter2), .O(gate252inter6));
  inv1  gate820(.a(G709), .O(gate252inter7));
  inv1  gate821(.a(G745), .O(gate252inter8));
  nand2 gate822(.a(gate252inter8), .b(gate252inter7), .O(gate252inter9));
  nand2 gate823(.a(s_39), .b(gate252inter3), .O(gate252inter10));
  nor2  gate824(.a(gate252inter10), .b(gate252inter9), .O(gate252inter11));
  nor2  gate825(.a(gate252inter11), .b(gate252inter6), .O(gate252inter12));
  nand2 gate826(.a(gate252inter12), .b(gate252inter1), .O(G765));
nand2 gate253( .a(G260), .b(G748), .O(G766) );
nand2 gate254( .a(G712), .b(G748), .O(G767) );
nand2 gate255( .a(G263), .b(G751), .O(G768) );

  xor2  gate2801(.a(G751), .b(G715), .O(gate256inter0));
  nand2 gate2802(.a(gate256inter0), .b(s_322), .O(gate256inter1));
  and2  gate2803(.a(G751), .b(G715), .O(gate256inter2));
  inv1  gate2804(.a(s_322), .O(gate256inter3));
  inv1  gate2805(.a(s_323), .O(gate256inter4));
  nand2 gate2806(.a(gate256inter4), .b(gate256inter3), .O(gate256inter5));
  nor2  gate2807(.a(gate256inter5), .b(gate256inter2), .O(gate256inter6));
  inv1  gate2808(.a(G715), .O(gate256inter7));
  inv1  gate2809(.a(G751), .O(gate256inter8));
  nand2 gate2810(.a(gate256inter8), .b(gate256inter7), .O(gate256inter9));
  nand2 gate2811(.a(s_323), .b(gate256inter3), .O(gate256inter10));
  nor2  gate2812(.a(gate256inter10), .b(gate256inter9), .O(gate256inter11));
  nor2  gate2813(.a(gate256inter11), .b(gate256inter6), .O(gate256inter12));
  nand2 gate2814(.a(gate256inter12), .b(gate256inter1), .O(G769));
nand2 gate257( .a(G754), .b(G755), .O(G770) );
nand2 gate258( .a(G756), .b(G757), .O(G773) );

  xor2  gate1499(.a(G759), .b(G758), .O(gate259inter0));
  nand2 gate1500(.a(gate259inter0), .b(s_136), .O(gate259inter1));
  and2  gate1501(.a(G759), .b(G758), .O(gate259inter2));
  inv1  gate1502(.a(s_136), .O(gate259inter3));
  inv1  gate1503(.a(s_137), .O(gate259inter4));
  nand2 gate1504(.a(gate259inter4), .b(gate259inter3), .O(gate259inter5));
  nor2  gate1505(.a(gate259inter5), .b(gate259inter2), .O(gate259inter6));
  inv1  gate1506(.a(G758), .O(gate259inter7));
  inv1  gate1507(.a(G759), .O(gate259inter8));
  nand2 gate1508(.a(gate259inter8), .b(gate259inter7), .O(gate259inter9));
  nand2 gate1509(.a(s_137), .b(gate259inter3), .O(gate259inter10));
  nor2  gate1510(.a(gate259inter10), .b(gate259inter9), .O(gate259inter11));
  nor2  gate1511(.a(gate259inter11), .b(gate259inter6), .O(gate259inter12));
  nand2 gate1512(.a(gate259inter12), .b(gate259inter1), .O(G776));
nand2 gate260( .a(G760), .b(G761), .O(G779) );

  xor2  gate1625(.a(G763), .b(G762), .O(gate261inter0));
  nand2 gate1626(.a(gate261inter0), .b(s_154), .O(gate261inter1));
  and2  gate1627(.a(G763), .b(G762), .O(gate261inter2));
  inv1  gate1628(.a(s_154), .O(gate261inter3));
  inv1  gate1629(.a(s_155), .O(gate261inter4));
  nand2 gate1630(.a(gate261inter4), .b(gate261inter3), .O(gate261inter5));
  nor2  gate1631(.a(gate261inter5), .b(gate261inter2), .O(gate261inter6));
  inv1  gate1632(.a(G762), .O(gate261inter7));
  inv1  gate1633(.a(G763), .O(gate261inter8));
  nand2 gate1634(.a(gate261inter8), .b(gate261inter7), .O(gate261inter9));
  nand2 gate1635(.a(s_155), .b(gate261inter3), .O(gate261inter10));
  nor2  gate1636(.a(gate261inter10), .b(gate261inter9), .O(gate261inter11));
  nor2  gate1637(.a(gate261inter11), .b(gate261inter6), .O(gate261inter12));
  nand2 gate1638(.a(gate261inter12), .b(gate261inter1), .O(G782));

  xor2  gate2325(.a(G765), .b(G764), .O(gate262inter0));
  nand2 gate2326(.a(gate262inter0), .b(s_254), .O(gate262inter1));
  and2  gate2327(.a(G765), .b(G764), .O(gate262inter2));
  inv1  gate2328(.a(s_254), .O(gate262inter3));
  inv1  gate2329(.a(s_255), .O(gate262inter4));
  nand2 gate2330(.a(gate262inter4), .b(gate262inter3), .O(gate262inter5));
  nor2  gate2331(.a(gate262inter5), .b(gate262inter2), .O(gate262inter6));
  inv1  gate2332(.a(G764), .O(gate262inter7));
  inv1  gate2333(.a(G765), .O(gate262inter8));
  nand2 gate2334(.a(gate262inter8), .b(gate262inter7), .O(gate262inter9));
  nand2 gate2335(.a(s_255), .b(gate262inter3), .O(gate262inter10));
  nor2  gate2336(.a(gate262inter10), .b(gate262inter9), .O(gate262inter11));
  nor2  gate2337(.a(gate262inter11), .b(gate262inter6), .O(gate262inter12));
  nand2 gate2338(.a(gate262inter12), .b(gate262inter1), .O(G785));
nand2 gate263( .a(G766), .b(G767), .O(G788) );
nand2 gate264( .a(G768), .b(G769), .O(G791) );

  xor2  gate1093(.a(G770), .b(G642), .O(gate265inter0));
  nand2 gate1094(.a(gate265inter0), .b(s_78), .O(gate265inter1));
  and2  gate1095(.a(G770), .b(G642), .O(gate265inter2));
  inv1  gate1096(.a(s_78), .O(gate265inter3));
  inv1  gate1097(.a(s_79), .O(gate265inter4));
  nand2 gate1098(.a(gate265inter4), .b(gate265inter3), .O(gate265inter5));
  nor2  gate1099(.a(gate265inter5), .b(gate265inter2), .O(gate265inter6));
  inv1  gate1100(.a(G642), .O(gate265inter7));
  inv1  gate1101(.a(G770), .O(gate265inter8));
  nand2 gate1102(.a(gate265inter8), .b(gate265inter7), .O(gate265inter9));
  nand2 gate1103(.a(s_79), .b(gate265inter3), .O(gate265inter10));
  nor2  gate1104(.a(gate265inter10), .b(gate265inter9), .O(gate265inter11));
  nor2  gate1105(.a(gate265inter11), .b(gate265inter6), .O(gate265inter12));
  nand2 gate1106(.a(gate265inter12), .b(gate265inter1), .O(G794));
nand2 gate266( .a(G645), .b(G773), .O(G797) );

  xor2  gate1429(.a(G776), .b(G648), .O(gate267inter0));
  nand2 gate1430(.a(gate267inter0), .b(s_126), .O(gate267inter1));
  and2  gate1431(.a(G776), .b(G648), .O(gate267inter2));
  inv1  gate1432(.a(s_126), .O(gate267inter3));
  inv1  gate1433(.a(s_127), .O(gate267inter4));
  nand2 gate1434(.a(gate267inter4), .b(gate267inter3), .O(gate267inter5));
  nor2  gate1435(.a(gate267inter5), .b(gate267inter2), .O(gate267inter6));
  inv1  gate1436(.a(G648), .O(gate267inter7));
  inv1  gate1437(.a(G776), .O(gate267inter8));
  nand2 gate1438(.a(gate267inter8), .b(gate267inter7), .O(gate267inter9));
  nand2 gate1439(.a(s_127), .b(gate267inter3), .O(gate267inter10));
  nor2  gate1440(.a(gate267inter10), .b(gate267inter9), .O(gate267inter11));
  nor2  gate1441(.a(gate267inter11), .b(gate267inter6), .O(gate267inter12));
  nand2 gate1442(.a(gate267inter12), .b(gate267inter1), .O(G800));
nand2 gate268( .a(G651), .b(G779), .O(G803) );
nand2 gate269( .a(G654), .b(G782), .O(G806) );
nand2 gate270( .a(G657), .b(G785), .O(G809) );
nand2 gate271( .a(G660), .b(G788), .O(G812) );
nand2 gate272( .a(G663), .b(G791), .O(G815) );
nand2 gate273( .a(G642), .b(G794), .O(G818) );
nand2 gate274( .a(G770), .b(G794), .O(G819) );

  xor2  gate2507(.a(G797), .b(G645), .O(gate275inter0));
  nand2 gate2508(.a(gate275inter0), .b(s_280), .O(gate275inter1));
  and2  gate2509(.a(G797), .b(G645), .O(gate275inter2));
  inv1  gate2510(.a(s_280), .O(gate275inter3));
  inv1  gate2511(.a(s_281), .O(gate275inter4));
  nand2 gate2512(.a(gate275inter4), .b(gate275inter3), .O(gate275inter5));
  nor2  gate2513(.a(gate275inter5), .b(gate275inter2), .O(gate275inter6));
  inv1  gate2514(.a(G645), .O(gate275inter7));
  inv1  gate2515(.a(G797), .O(gate275inter8));
  nand2 gate2516(.a(gate275inter8), .b(gate275inter7), .O(gate275inter9));
  nand2 gate2517(.a(s_281), .b(gate275inter3), .O(gate275inter10));
  nor2  gate2518(.a(gate275inter10), .b(gate275inter9), .O(gate275inter11));
  nor2  gate2519(.a(gate275inter11), .b(gate275inter6), .O(gate275inter12));
  nand2 gate2520(.a(gate275inter12), .b(gate275inter1), .O(G820));

  xor2  gate1821(.a(G797), .b(G773), .O(gate276inter0));
  nand2 gate1822(.a(gate276inter0), .b(s_182), .O(gate276inter1));
  and2  gate1823(.a(G797), .b(G773), .O(gate276inter2));
  inv1  gate1824(.a(s_182), .O(gate276inter3));
  inv1  gate1825(.a(s_183), .O(gate276inter4));
  nand2 gate1826(.a(gate276inter4), .b(gate276inter3), .O(gate276inter5));
  nor2  gate1827(.a(gate276inter5), .b(gate276inter2), .O(gate276inter6));
  inv1  gate1828(.a(G773), .O(gate276inter7));
  inv1  gate1829(.a(G797), .O(gate276inter8));
  nand2 gate1830(.a(gate276inter8), .b(gate276inter7), .O(gate276inter9));
  nand2 gate1831(.a(s_183), .b(gate276inter3), .O(gate276inter10));
  nor2  gate1832(.a(gate276inter10), .b(gate276inter9), .O(gate276inter11));
  nor2  gate1833(.a(gate276inter11), .b(gate276inter6), .O(gate276inter12));
  nand2 gate1834(.a(gate276inter12), .b(gate276inter1), .O(G821));
nand2 gate277( .a(G648), .b(G800), .O(G822) );

  xor2  gate2605(.a(G800), .b(G776), .O(gate278inter0));
  nand2 gate2606(.a(gate278inter0), .b(s_294), .O(gate278inter1));
  and2  gate2607(.a(G800), .b(G776), .O(gate278inter2));
  inv1  gate2608(.a(s_294), .O(gate278inter3));
  inv1  gate2609(.a(s_295), .O(gate278inter4));
  nand2 gate2610(.a(gate278inter4), .b(gate278inter3), .O(gate278inter5));
  nor2  gate2611(.a(gate278inter5), .b(gate278inter2), .O(gate278inter6));
  inv1  gate2612(.a(G776), .O(gate278inter7));
  inv1  gate2613(.a(G800), .O(gate278inter8));
  nand2 gate2614(.a(gate278inter8), .b(gate278inter7), .O(gate278inter9));
  nand2 gate2615(.a(s_295), .b(gate278inter3), .O(gate278inter10));
  nor2  gate2616(.a(gate278inter10), .b(gate278inter9), .O(gate278inter11));
  nor2  gate2617(.a(gate278inter11), .b(gate278inter6), .O(gate278inter12));
  nand2 gate2618(.a(gate278inter12), .b(gate278inter1), .O(G823));
nand2 gate279( .a(G651), .b(G803), .O(G824) );

  xor2  gate967(.a(G803), .b(G779), .O(gate280inter0));
  nand2 gate968(.a(gate280inter0), .b(s_60), .O(gate280inter1));
  and2  gate969(.a(G803), .b(G779), .O(gate280inter2));
  inv1  gate970(.a(s_60), .O(gate280inter3));
  inv1  gate971(.a(s_61), .O(gate280inter4));
  nand2 gate972(.a(gate280inter4), .b(gate280inter3), .O(gate280inter5));
  nor2  gate973(.a(gate280inter5), .b(gate280inter2), .O(gate280inter6));
  inv1  gate974(.a(G779), .O(gate280inter7));
  inv1  gate975(.a(G803), .O(gate280inter8));
  nand2 gate976(.a(gate280inter8), .b(gate280inter7), .O(gate280inter9));
  nand2 gate977(.a(s_61), .b(gate280inter3), .O(gate280inter10));
  nor2  gate978(.a(gate280inter10), .b(gate280inter9), .O(gate280inter11));
  nor2  gate979(.a(gate280inter11), .b(gate280inter6), .O(gate280inter12));
  nand2 gate980(.a(gate280inter12), .b(gate280inter1), .O(G825));
nand2 gate281( .a(G654), .b(G806), .O(G826) );

  xor2  gate953(.a(G806), .b(G782), .O(gate282inter0));
  nand2 gate954(.a(gate282inter0), .b(s_58), .O(gate282inter1));
  and2  gate955(.a(G806), .b(G782), .O(gate282inter2));
  inv1  gate956(.a(s_58), .O(gate282inter3));
  inv1  gate957(.a(s_59), .O(gate282inter4));
  nand2 gate958(.a(gate282inter4), .b(gate282inter3), .O(gate282inter5));
  nor2  gate959(.a(gate282inter5), .b(gate282inter2), .O(gate282inter6));
  inv1  gate960(.a(G782), .O(gate282inter7));
  inv1  gate961(.a(G806), .O(gate282inter8));
  nand2 gate962(.a(gate282inter8), .b(gate282inter7), .O(gate282inter9));
  nand2 gate963(.a(s_59), .b(gate282inter3), .O(gate282inter10));
  nor2  gate964(.a(gate282inter10), .b(gate282inter9), .O(gate282inter11));
  nor2  gate965(.a(gate282inter11), .b(gate282inter6), .O(gate282inter12));
  nand2 gate966(.a(gate282inter12), .b(gate282inter1), .O(G827));
nand2 gate283( .a(G657), .b(G809), .O(G828) );
nand2 gate284( .a(G785), .b(G809), .O(G829) );

  xor2  gate1891(.a(G812), .b(G660), .O(gate285inter0));
  nand2 gate1892(.a(gate285inter0), .b(s_192), .O(gate285inter1));
  and2  gate1893(.a(G812), .b(G660), .O(gate285inter2));
  inv1  gate1894(.a(s_192), .O(gate285inter3));
  inv1  gate1895(.a(s_193), .O(gate285inter4));
  nand2 gate1896(.a(gate285inter4), .b(gate285inter3), .O(gate285inter5));
  nor2  gate1897(.a(gate285inter5), .b(gate285inter2), .O(gate285inter6));
  inv1  gate1898(.a(G660), .O(gate285inter7));
  inv1  gate1899(.a(G812), .O(gate285inter8));
  nand2 gate1900(.a(gate285inter8), .b(gate285inter7), .O(gate285inter9));
  nand2 gate1901(.a(s_193), .b(gate285inter3), .O(gate285inter10));
  nor2  gate1902(.a(gate285inter10), .b(gate285inter9), .O(gate285inter11));
  nor2  gate1903(.a(gate285inter11), .b(gate285inter6), .O(gate285inter12));
  nand2 gate1904(.a(gate285inter12), .b(gate285inter1), .O(G830));
nand2 gate286( .a(G788), .b(G812), .O(G831) );
nand2 gate287( .a(G663), .b(G815), .O(G832) );
nand2 gate288( .a(G791), .b(G815), .O(G833) );

  xor2  gate897(.a(G819), .b(G818), .O(gate289inter0));
  nand2 gate898(.a(gate289inter0), .b(s_50), .O(gate289inter1));
  and2  gate899(.a(G819), .b(G818), .O(gate289inter2));
  inv1  gate900(.a(s_50), .O(gate289inter3));
  inv1  gate901(.a(s_51), .O(gate289inter4));
  nand2 gate902(.a(gate289inter4), .b(gate289inter3), .O(gate289inter5));
  nor2  gate903(.a(gate289inter5), .b(gate289inter2), .O(gate289inter6));
  inv1  gate904(.a(G818), .O(gate289inter7));
  inv1  gate905(.a(G819), .O(gate289inter8));
  nand2 gate906(.a(gate289inter8), .b(gate289inter7), .O(gate289inter9));
  nand2 gate907(.a(s_51), .b(gate289inter3), .O(gate289inter10));
  nor2  gate908(.a(gate289inter10), .b(gate289inter9), .O(gate289inter11));
  nor2  gate909(.a(gate289inter11), .b(gate289inter6), .O(gate289inter12));
  nand2 gate910(.a(gate289inter12), .b(gate289inter1), .O(G834));
nand2 gate290( .a(G820), .b(G821), .O(G847) );
nand2 gate291( .a(G822), .b(G823), .O(G860) );

  xor2  gate3053(.a(G825), .b(G824), .O(gate292inter0));
  nand2 gate3054(.a(gate292inter0), .b(s_358), .O(gate292inter1));
  and2  gate3055(.a(G825), .b(G824), .O(gate292inter2));
  inv1  gate3056(.a(s_358), .O(gate292inter3));
  inv1  gate3057(.a(s_359), .O(gate292inter4));
  nand2 gate3058(.a(gate292inter4), .b(gate292inter3), .O(gate292inter5));
  nor2  gate3059(.a(gate292inter5), .b(gate292inter2), .O(gate292inter6));
  inv1  gate3060(.a(G824), .O(gate292inter7));
  inv1  gate3061(.a(G825), .O(gate292inter8));
  nand2 gate3062(.a(gate292inter8), .b(gate292inter7), .O(gate292inter9));
  nand2 gate3063(.a(s_359), .b(gate292inter3), .O(gate292inter10));
  nor2  gate3064(.a(gate292inter10), .b(gate292inter9), .O(gate292inter11));
  nor2  gate3065(.a(gate292inter11), .b(gate292inter6), .O(gate292inter12));
  nand2 gate3066(.a(gate292inter12), .b(gate292inter1), .O(G873));
nand2 gate293( .a(G828), .b(G829), .O(G886) );
nand2 gate294( .a(G832), .b(G833), .O(G899) );
nand2 gate295( .a(G830), .b(G831), .O(G912) );
nand2 gate296( .a(G826), .b(G827), .O(G925) );
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );

  xor2  gate2899(.a(G1036), .b(G1), .O(gate387inter0));
  nand2 gate2900(.a(gate387inter0), .b(s_336), .O(gate387inter1));
  and2  gate2901(.a(G1036), .b(G1), .O(gate387inter2));
  inv1  gate2902(.a(s_336), .O(gate387inter3));
  inv1  gate2903(.a(s_337), .O(gate387inter4));
  nand2 gate2904(.a(gate387inter4), .b(gate387inter3), .O(gate387inter5));
  nor2  gate2905(.a(gate387inter5), .b(gate387inter2), .O(gate387inter6));
  inv1  gate2906(.a(G1), .O(gate387inter7));
  inv1  gate2907(.a(G1036), .O(gate387inter8));
  nand2 gate2908(.a(gate387inter8), .b(gate387inter7), .O(gate387inter9));
  nand2 gate2909(.a(s_337), .b(gate387inter3), .O(gate387inter10));
  nor2  gate2910(.a(gate387inter10), .b(gate387inter9), .O(gate387inter11));
  nor2  gate2911(.a(gate387inter11), .b(gate387inter6), .O(gate387inter12));
  nand2 gate2912(.a(gate387inter12), .b(gate387inter1), .O(G1132));

  xor2  gate2983(.a(G1039), .b(G2), .O(gate388inter0));
  nand2 gate2984(.a(gate388inter0), .b(s_348), .O(gate388inter1));
  and2  gate2985(.a(G1039), .b(G2), .O(gate388inter2));
  inv1  gate2986(.a(s_348), .O(gate388inter3));
  inv1  gate2987(.a(s_349), .O(gate388inter4));
  nand2 gate2988(.a(gate388inter4), .b(gate388inter3), .O(gate388inter5));
  nor2  gate2989(.a(gate388inter5), .b(gate388inter2), .O(gate388inter6));
  inv1  gate2990(.a(G2), .O(gate388inter7));
  inv1  gate2991(.a(G1039), .O(gate388inter8));
  nand2 gate2992(.a(gate388inter8), .b(gate388inter7), .O(gate388inter9));
  nand2 gate2993(.a(s_349), .b(gate388inter3), .O(gate388inter10));
  nor2  gate2994(.a(gate388inter10), .b(gate388inter9), .O(gate388inter11));
  nor2  gate2995(.a(gate388inter11), .b(gate388inter6), .O(gate388inter12));
  nand2 gate2996(.a(gate388inter12), .b(gate388inter1), .O(G1135));

  xor2  gate771(.a(G1042), .b(G3), .O(gate389inter0));
  nand2 gate772(.a(gate389inter0), .b(s_32), .O(gate389inter1));
  and2  gate773(.a(G1042), .b(G3), .O(gate389inter2));
  inv1  gate774(.a(s_32), .O(gate389inter3));
  inv1  gate775(.a(s_33), .O(gate389inter4));
  nand2 gate776(.a(gate389inter4), .b(gate389inter3), .O(gate389inter5));
  nor2  gate777(.a(gate389inter5), .b(gate389inter2), .O(gate389inter6));
  inv1  gate778(.a(G3), .O(gate389inter7));
  inv1  gate779(.a(G1042), .O(gate389inter8));
  nand2 gate780(.a(gate389inter8), .b(gate389inter7), .O(gate389inter9));
  nand2 gate781(.a(s_33), .b(gate389inter3), .O(gate389inter10));
  nor2  gate782(.a(gate389inter10), .b(gate389inter9), .O(gate389inter11));
  nor2  gate783(.a(gate389inter11), .b(gate389inter6), .O(gate389inter12));
  nand2 gate784(.a(gate389inter12), .b(gate389inter1), .O(G1138));
nand2 gate390( .a(G4), .b(G1045), .O(G1141) );

  xor2  gate1177(.a(G1048), .b(G5), .O(gate391inter0));
  nand2 gate1178(.a(gate391inter0), .b(s_90), .O(gate391inter1));
  and2  gate1179(.a(G1048), .b(G5), .O(gate391inter2));
  inv1  gate1180(.a(s_90), .O(gate391inter3));
  inv1  gate1181(.a(s_91), .O(gate391inter4));
  nand2 gate1182(.a(gate391inter4), .b(gate391inter3), .O(gate391inter5));
  nor2  gate1183(.a(gate391inter5), .b(gate391inter2), .O(gate391inter6));
  inv1  gate1184(.a(G5), .O(gate391inter7));
  inv1  gate1185(.a(G1048), .O(gate391inter8));
  nand2 gate1186(.a(gate391inter8), .b(gate391inter7), .O(gate391inter9));
  nand2 gate1187(.a(s_91), .b(gate391inter3), .O(gate391inter10));
  nor2  gate1188(.a(gate391inter10), .b(gate391inter9), .O(gate391inter11));
  nor2  gate1189(.a(gate391inter11), .b(gate391inter6), .O(gate391inter12));
  nand2 gate1190(.a(gate391inter12), .b(gate391inter1), .O(G1144));

  xor2  gate2535(.a(G1051), .b(G6), .O(gate392inter0));
  nand2 gate2536(.a(gate392inter0), .b(s_284), .O(gate392inter1));
  and2  gate2537(.a(G1051), .b(G6), .O(gate392inter2));
  inv1  gate2538(.a(s_284), .O(gate392inter3));
  inv1  gate2539(.a(s_285), .O(gate392inter4));
  nand2 gate2540(.a(gate392inter4), .b(gate392inter3), .O(gate392inter5));
  nor2  gate2541(.a(gate392inter5), .b(gate392inter2), .O(gate392inter6));
  inv1  gate2542(.a(G6), .O(gate392inter7));
  inv1  gate2543(.a(G1051), .O(gate392inter8));
  nand2 gate2544(.a(gate392inter8), .b(gate392inter7), .O(gate392inter9));
  nand2 gate2545(.a(s_285), .b(gate392inter3), .O(gate392inter10));
  nor2  gate2546(.a(gate392inter10), .b(gate392inter9), .O(gate392inter11));
  nor2  gate2547(.a(gate392inter11), .b(gate392inter6), .O(gate392inter12));
  nand2 gate2548(.a(gate392inter12), .b(gate392inter1), .O(G1147));
nand2 gate393( .a(G7), .b(G1054), .O(G1150) );
nand2 gate394( .a(G8), .b(G1057), .O(G1153) );
nand2 gate395( .a(G9), .b(G1060), .O(G1156) );
nand2 gate396( .a(G10), .b(G1063), .O(G1159) );
nand2 gate397( .a(G11), .b(G1066), .O(G1162) );
nand2 gate398( .a(G12), .b(G1069), .O(G1165) );

  xor2  gate1387(.a(G1072), .b(G13), .O(gate399inter0));
  nand2 gate1388(.a(gate399inter0), .b(s_120), .O(gate399inter1));
  and2  gate1389(.a(G1072), .b(G13), .O(gate399inter2));
  inv1  gate1390(.a(s_120), .O(gate399inter3));
  inv1  gate1391(.a(s_121), .O(gate399inter4));
  nand2 gate1392(.a(gate399inter4), .b(gate399inter3), .O(gate399inter5));
  nor2  gate1393(.a(gate399inter5), .b(gate399inter2), .O(gate399inter6));
  inv1  gate1394(.a(G13), .O(gate399inter7));
  inv1  gate1395(.a(G1072), .O(gate399inter8));
  nand2 gate1396(.a(gate399inter8), .b(gate399inter7), .O(gate399inter9));
  nand2 gate1397(.a(s_121), .b(gate399inter3), .O(gate399inter10));
  nor2  gate1398(.a(gate399inter10), .b(gate399inter9), .O(gate399inter11));
  nor2  gate1399(.a(gate399inter11), .b(gate399inter6), .O(gate399inter12));
  nand2 gate1400(.a(gate399inter12), .b(gate399inter1), .O(G1168));

  xor2  gate1051(.a(G1075), .b(G14), .O(gate400inter0));
  nand2 gate1052(.a(gate400inter0), .b(s_72), .O(gate400inter1));
  and2  gate1053(.a(G1075), .b(G14), .O(gate400inter2));
  inv1  gate1054(.a(s_72), .O(gate400inter3));
  inv1  gate1055(.a(s_73), .O(gate400inter4));
  nand2 gate1056(.a(gate400inter4), .b(gate400inter3), .O(gate400inter5));
  nor2  gate1057(.a(gate400inter5), .b(gate400inter2), .O(gate400inter6));
  inv1  gate1058(.a(G14), .O(gate400inter7));
  inv1  gate1059(.a(G1075), .O(gate400inter8));
  nand2 gate1060(.a(gate400inter8), .b(gate400inter7), .O(gate400inter9));
  nand2 gate1061(.a(s_73), .b(gate400inter3), .O(gate400inter10));
  nor2  gate1062(.a(gate400inter10), .b(gate400inter9), .O(gate400inter11));
  nor2  gate1063(.a(gate400inter11), .b(gate400inter6), .O(gate400inter12));
  nand2 gate1064(.a(gate400inter12), .b(gate400inter1), .O(G1171));
nand2 gate401( .a(G15), .b(G1078), .O(G1174) );
nand2 gate402( .a(G16), .b(G1081), .O(G1177) );
nand2 gate403( .a(G17), .b(G1084), .O(G1180) );
nand2 gate404( .a(G18), .b(G1087), .O(G1183) );
nand2 gate405( .a(G19), .b(G1090), .O(G1186) );
nand2 gate406( .a(G20), .b(G1093), .O(G1189) );
nand2 gate407( .a(G21), .b(G1096), .O(G1192) );

  xor2  gate2787(.a(G1099), .b(G22), .O(gate408inter0));
  nand2 gate2788(.a(gate408inter0), .b(s_320), .O(gate408inter1));
  and2  gate2789(.a(G1099), .b(G22), .O(gate408inter2));
  inv1  gate2790(.a(s_320), .O(gate408inter3));
  inv1  gate2791(.a(s_321), .O(gate408inter4));
  nand2 gate2792(.a(gate408inter4), .b(gate408inter3), .O(gate408inter5));
  nor2  gate2793(.a(gate408inter5), .b(gate408inter2), .O(gate408inter6));
  inv1  gate2794(.a(G22), .O(gate408inter7));
  inv1  gate2795(.a(G1099), .O(gate408inter8));
  nand2 gate2796(.a(gate408inter8), .b(gate408inter7), .O(gate408inter9));
  nand2 gate2797(.a(s_321), .b(gate408inter3), .O(gate408inter10));
  nor2  gate2798(.a(gate408inter10), .b(gate408inter9), .O(gate408inter11));
  nor2  gate2799(.a(gate408inter11), .b(gate408inter6), .O(gate408inter12));
  nand2 gate2800(.a(gate408inter12), .b(gate408inter1), .O(G1195));

  xor2  gate1317(.a(G1102), .b(G23), .O(gate409inter0));
  nand2 gate1318(.a(gate409inter0), .b(s_110), .O(gate409inter1));
  and2  gate1319(.a(G1102), .b(G23), .O(gate409inter2));
  inv1  gate1320(.a(s_110), .O(gate409inter3));
  inv1  gate1321(.a(s_111), .O(gate409inter4));
  nand2 gate1322(.a(gate409inter4), .b(gate409inter3), .O(gate409inter5));
  nor2  gate1323(.a(gate409inter5), .b(gate409inter2), .O(gate409inter6));
  inv1  gate1324(.a(G23), .O(gate409inter7));
  inv1  gate1325(.a(G1102), .O(gate409inter8));
  nand2 gate1326(.a(gate409inter8), .b(gate409inter7), .O(gate409inter9));
  nand2 gate1327(.a(s_111), .b(gate409inter3), .O(gate409inter10));
  nor2  gate1328(.a(gate409inter10), .b(gate409inter9), .O(gate409inter11));
  nor2  gate1329(.a(gate409inter11), .b(gate409inter6), .O(gate409inter12));
  nand2 gate1330(.a(gate409inter12), .b(gate409inter1), .O(G1198));

  xor2  gate2577(.a(G1105), .b(G24), .O(gate410inter0));
  nand2 gate2578(.a(gate410inter0), .b(s_290), .O(gate410inter1));
  and2  gate2579(.a(G1105), .b(G24), .O(gate410inter2));
  inv1  gate2580(.a(s_290), .O(gate410inter3));
  inv1  gate2581(.a(s_291), .O(gate410inter4));
  nand2 gate2582(.a(gate410inter4), .b(gate410inter3), .O(gate410inter5));
  nor2  gate2583(.a(gate410inter5), .b(gate410inter2), .O(gate410inter6));
  inv1  gate2584(.a(G24), .O(gate410inter7));
  inv1  gate2585(.a(G1105), .O(gate410inter8));
  nand2 gate2586(.a(gate410inter8), .b(gate410inter7), .O(gate410inter9));
  nand2 gate2587(.a(s_291), .b(gate410inter3), .O(gate410inter10));
  nor2  gate2588(.a(gate410inter10), .b(gate410inter9), .O(gate410inter11));
  nor2  gate2589(.a(gate410inter11), .b(gate410inter6), .O(gate410inter12));
  nand2 gate2590(.a(gate410inter12), .b(gate410inter1), .O(G1201));

  xor2  gate785(.a(G1108), .b(G25), .O(gate411inter0));
  nand2 gate786(.a(gate411inter0), .b(s_34), .O(gate411inter1));
  and2  gate787(.a(G1108), .b(G25), .O(gate411inter2));
  inv1  gate788(.a(s_34), .O(gate411inter3));
  inv1  gate789(.a(s_35), .O(gate411inter4));
  nand2 gate790(.a(gate411inter4), .b(gate411inter3), .O(gate411inter5));
  nor2  gate791(.a(gate411inter5), .b(gate411inter2), .O(gate411inter6));
  inv1  gate792(.a(G25), .O(gate411inter7));
  inv1  gate793(.a(G1108), .O(gate411inter8));
  nand2 gate794(.a(gate411inter8), .b(gate411inter7), .O(gate411inter9));
  nand2 gate795(.a(s_35), .b(gate411inter3), .O(gate411inter10));
  nor2  gate796(.a(gate411inter10), .b(gate411inter9), .O(gate411inter11));
  nor2  gate797(.a(gate411inter11), .b(gate411inter6), .O(gate411inter12));
  nand2 gate798(.a(gate411inter12), .b(gate411inter1), .O(G1204));
nand2 gate412( .a(G26), .b(G1111), .O(G1207) );

  xor2  gate715(.a(G1114), .b(G27), .O(gate413inter0));
  nand2 gate716(.a(gate413inter0), .b(s_24), .O(gate413inter1));
  and2  gate717(.a(G1114), .b(G27), .O(gate413inter2));
  inv1  gate718(.a(s_24), .O(gate413inter3));
  inv1  gate719(.a(s_25), .O(gate413inter4));
  nand2 gate720(.a(gate413inter4), .b(gate413inter3), .O(gate413inter5));
  nor2  gate721(.a(gate413inter5), .b(gate413inter2), .O(gate413inter6));
  inv1  gate722(.a(G27), .O(gate413inter7));
  inv1  gate723(.a(G1114), .O(gate413inter8));
  nand2 gate724(.a(gate413inter8), .b(gate413inter7), .O(gate413inter9));
  nand2 gate725(.a(s_25), .b(gate413inter3), .O(gate413inter10));
  nor2  gate726(.a(gate413inter10), .b(gate413inter9), .O(gate413inter11));
  nor2  gate727(.a(gate413inter11), .b(gate413inter6), .O(gate413inter12));
  nand2 gate728(.a(gate413inter12), .b(gate413inter1), .O(G1210));
nand2 gate414( .a(G28), .b(G1117), .O(G1213) );
nand2 gate415( .a(G29), .b(G1120), .O(G1216) );
nand2 gate416( .a(G30), .b(G1123), .O(G1219) );
nand2 gate417( .a(G31), .b(G1126), .O(G1222) );
nand2 gate418( .a(G32), .b(G1129), .O(G1225) );

  xor2  gate1219(.a(G1132), .b(G1), .O(gate419inter0));
  nand2 gate1220(.a(gate419inter0), .b(s_96), .O(gate419inter1));
  and2  gate1221(.a(G1132), .b(G1), .O(gate419inter2));
  inv1  gate1222(.a(s_96), .O(gate419inter3));
  inv1  gate1223(.a(s_97), .O(gate419inter4));
  nand2 gate1224(.a(gate419inter4), .b(gate419inter3), .O(gate419inter5));
  nor2  gate1225(.a(gate419inter5), .b(gate419inter2), .O(gate419inter6));
  inv1  gate1226(.a(G1), .O(gate419inter7));
  inv1  gate1227(.a(G1132), .O(gate419inter8));
  nand2 gate1228(.a(gate419inter8), .b(gate419inter7), .O(gate419inter9));
  nand2 gate1229(.a(s_97), .b(gate419inter3), .O(gate419inter10));
  nor2  gate1230(.a(gate419inter10), .b(gate419inter9), .O(gate419inter11));
  nor2  gate1231(.a(gate419inter11), .b(gate419inter6), .O(gate419inter12));
  nand2 gate1232(.a(gate419inter12), .b(gate419inter1), .O(G1228));

  xor2  gate1345(.a(G1132), .b(G1036), .O(gate420inter0));
  nand2 gate1346(.a(gate420inter0), .b(s_114), .O(gate420inter1));
  and2  gate1347(.a(G1132), .b(G1036), .O(gate420inter2));
  inv1  gate1348(.a(s_114), .O(gate420inter3));
  inv1  gate1349(.a(s_115), .O(gate420inter4));
  nand2 gate1350(.a(gate420inter4), .b(gate420inter3), .O(gate420inter5));
  nor2  gate1351(.a(gate420inter5), .b(gate420inter2), .O(gate420inter6));
  inv1  gate1352(.a(G1036), .O(gate420inter7));
  inv1  gate1353(.a(G1132), .O(gate420inter8));
  nand2 gate1354(.a(gate420inter8), .b(gate420inter7), .O(gate420inter9));
  nand2 gate1355(.a(s_115), .b(gate420inter3), .O(gate420inter10));
  nor2  gate1356(.a(gate420inter10), .b(gate420inter9), .O(gate420inter11));
  nor2  gate1357(.a(gate420inter11), .b(gate420inter6), .O(gate420inter12));
  nand2 gate1358(.a(gate420inter12), .b(gate420inter1), .O(G1229));
nand2 gate421( .a(G2), .b(G1135), .O(G1230) );
nand2 gate422( .a(G1039), .b(G1135), .O(G1231) );

  xor2  gate1667(.a(G1138), .b(G3), .O(gate423inter0));
  nand2 gate1668(.a(gate423inter0), .b(s_160), .O(gate423inter1));
  and2  gate1669(.a(G1138), .b(G3), .O(gate423inter2));
  inv1  gate1670(.a(s_160), .O(gate423inter3));
  inv1  gate1671(.a(s_161), .O(gate423inter4));
  nand2 gate1672(.a(gate423inter4), .b(gate423inter3), .O(gate423inter5));
  nor2  gate1673(.a(gate423inter5), .b(gate423inter2), .O(gate423inter6));
  inv1  gate1674(.a(G3), .O(gate423inter7));
  inv1  gate1675(.a(G1138), .O(gate423inter8));
  nand2 gate1676(.a(gate423inter8), .b(gate423inter7), .O(gate423inter9));
  nand2 gate1677(.a(s_161), .b(gate423inter3), .O(gate423inter10));
  nor2  gate1678(.a(gate423inter10), .b(gate423inter9), .O(gate423inter11));
  nor2  gate1679(.a(gate423inter11), .b(gate423inter6), .O(gate423inter12));
  nand2 gate1680(.a(gate423inter12), .b(gate423inter1), .O(G1232));
nand2 gate424( .a(G1042), .b(G1138), .O(G1233) );

  xor2  gate1933(.a(G1141), .b(G4), .O(gate425inter0));
  nand2 gate1934(.a(gate425inter0), .b(s_198), .O(gate425inter1));
  and2  gate1935(.a(G1141), .b(G4), .O(gate425inter2));
  inv1  gate1936(.a(s_198), .O(gate425inter3));
  inv1  gate1937(.a(s_199), .O(gate425inter4));
  nand2 gate1938(.a(gate425inter4), .b(gate425inter3), .O(gate425inter5));
  nor2  gate1939(.a(gate425inter5), .b(gate425inter2), .O(gate425inter6));
  inv1  gate1940(.a(G4), .O(gate425inter7));
  inv1  gate1941(.a(G1141), .O(gate425inter8));
  nand2 gate1942(.a(gate425inter8), .b(gate425inter7), .O(gate425inter9));
  nand2 gate1943(.a(s_199), .b(gate425inter3), .O(gate425inter10));
  nor2  gate1944(.a(gate425inter10), .b(gate425inter9), .O(gate425inter11));
  nor2  gate1945(.a(gate425inter11), .b(gate425inter6), .O(gate425inter12));
  nand2 gate1946(.a(gate425inter12), .b(gate425inter1), .O(G1234));

  xor2  gate2941(.a(G1141), .b(G1045), .O(gate426inter0));
  nand2 gate2942(.a(gate426inter0), .b(s_342), .O(gate426inter1));
  and2  gate2943(.a(G1141), .b(G1045), .O(gate426inter2));
  inv1  gate2944(.a(s_342), .O(gate426inter3));
  inv1  gate2945(.a(s_343), .O(gate426inter4));
  nand2 gate2946(.a(gate426inter4), .b(gate426inter3), .O(gate426inter5));
  nor2  gate2947(.a(gate426inter5), .b(gate426inter2), .O(gate426inter6));
  inv1  gate2948(.a(G1045), .O(gate426inter7));
  inv1  gate2949(.a(G1141), .O(gate426inter8));
  nand2 gate2950(.a(gate426inter8), .b(gate426inter7), .O(gate426inter9));
  nand2 gate2951(.a(s_343), .b(gate426inter3), .O(gate426inter10));
  nor2  gate2952(.a(gate426inter10), .b(gate426inter9), .O(gate426inter11));
  nor2  gate2953(.a(gate426inter11), .b(gate426inter6), .O(gate426inter12));
  nand2 gate2954(.a(gate426inter12), .b(gate426inter1), .O(G1235));

  xor2  gate1275(.a(G1144), .b(G5), .O(gate427inter0));
  nand2 gate1276(.a(gate427inter0), .b(s_104), .O(gate427inter1));
  and2  gate1277(.a(G1144), .b(G5), .O(gate427inter2));
  inv1  gate1278(.a(s_104), .O(gate427inter3));
  inv1  gate1279(.a(s_105), .O(gate427inter4));
  nand2 gate1280(.a(gate427inter4), .b(gate427inter3), .O(gate427inter5));
  nor2  gate1281(.a(gate427inter5), .b(gate427inter2), .O(gate427inter6));
  inv1  gate1282(.a(G5), .O(gate427inter7));
  inv1  gate1283(.a(G1144), .O(gate427inter8));
  nand2 gate1284(.a(gate427inter8), .b(gate427inter7), .O(gate427inter9));
  nand2 gate1285(.a(s_105), .b(gate427inter3), .O(gate427inter10));
  nor2  gate1286(.a(gate427inter10), .b(gate427inter9), .O(gate427inter11));
  nor2  gate1287(.a(gate427inter11), .b(gate427inter6), .O(gate427inter12));
  nand2 gate1288(.a(gate427inter12), .b(gate427inter1), .O(G1236));
nand2 gate428( .a(G1048), .b(G1144), .O(G1237) );

  xor2  gate1359(.a(G1147), .b(G6), .O(gate429inter0));
  nand2 gate1360(.a(gate429inter0), .b(s_116), .O(gate429inter1));
  and2  gate1361(.a(G1147), .b(G6), .O(gate429inter2));
  inv1  gate1362(.a(s_116), .O(gate429inter3));
  inv1  gate1363(.a(s_117), .O(gate429inter4));
  nand2 gate1364(.a(gate429inter4), .b(gate429inter3), .O(gate429inter5));
  nor2  gate1365(.a(gate429inter5), .b(gate429inter2), .O(gate429inter6));
  inv1  gate1366(.a(G6), .O(gate429inter7));
  inv1  gate1367(.a(G1147), .O(gate429inter8));
  nand2 gate1368(.a(gate429inter8), .b(gate429inter7), .O(gate429inter9));
  nand2 gate1369(.a(s_117), .b(gate429inter3), .O(gate429inter10));
  nor2  gate1370(.a(gate429inter10), .b(gate429inter9), .O(gate429inter11));
  nor2  gate1371(.a(gate429inter11), .b(gate429inter6), .O(gate429inter12));
  nand2 gate1372(.a(gate429inter12), .b(gate429inter1), .O(G1238));
nand2 gate430( .a(G1051), .b(G1147), .O(G1239) );
nand2 gate431( .a(G7), .b(G1150), .O(G1240) );
nand2 gate432( .a(G1054), .b(G1150), .O(G1241) );

  xor2  gate2339(.a(G1153), .b(G8), .O(gate433inter0));
  nand2 gate2340(.a(gate433inter0), .b(s_256), .O(gate433inter1));
  and2  gate2341(.a(G1153), .b(G8), .O(gate433inter2));
  inv1  gate2342(.a(s_256), .O(gate433inter3));
  inv1  gate2343(.a(s_257), .O(gate433inter4));
  nand2 gate2344(.a(gate433inter4), .b(gate433inter3), .O(gate433inter5));
  nor2  gate2345(.a(gate433inter5), .b(gate433inter2), .O(gate433inter6));
  inv1  gate2346(.a(G8), .O(gate433inter7));
  inv1  gate2347(.a(G1153), .O(gate433inter8));
  nand2 gate2348(.a(gate433inter8), .b(gate433inter7), .O(gate433inter9));
  nand2 gate2349(.a(s_257), .b(gate433inter3), .O(gate433inter10));
  nor2  gate2350(.a(gate433inter10), .b(gate433inter9), .O(gate433inter11));
  nor2  gate2351(.a(gate433inter11), .b(gate433inter6), .O(gate433inter12));
  nand2 gate2352(.a(gate433inter12), .b(gate433inter1), .O(G1242));

  xor2  gate883(.a(G1153), .b(G1057), .O(gate434inter0));
  nand2 gate884(.a(gate434inter0), .b(s_48), .O(gate434inter1));
  and2  gate885(.a(G1153), .b(G1057), .O(gate434inter2));
  inv1  gate886(.a(s_48), .O(gate434inter3));
  inv1  gate887(.a(s_49), .O(gate434inter4));
  nand2 gate888(.a(gate434inter4), .b(gate434inter3), .O(gate434inter5));
  nor2  gate889(.a(gate434inter5), .b(gate434inter2), .O(gate434inter6));
  inv1  gate890(.a(G1057), .O(gate434inter7));
  inv1  gate891(.a(G1153), .O(gate434inter8));
  nand2 gate892(.a(gate434inter8), .b(gate434inter7), .O(gate434inter9));
  nand2 gate893(.a(s_49), .b(gate434inter3), .O(gate434inter10));
  nor2  gate894(.a(gate434inter10), .b(gate434inter9), .O(gate434inter11));
  nor2  gate895(.a(gate434inter11), .b(gate434inter6), .O(gate434inter12));
  nand2 gate896(.a(gate434inter12), .b(gate434inter1), .O(G1243));
nand2 gate435( .a(G9), .b(G1156), .O(G1244) );

  xor2  gate925(.a(G1156), .b(G1060), .O(gate436inter0));
  nand2 gate926(.a(gate436inter0), .b(s_54), .O(gate436inter1));
  and2  gate927(.a(G1156), .b(G1060), .O(gate436inter2));
  inv1  gate928(.a(s_54), .O(gate436inter3));
  inv1  gate929(.a(s_55), .O(gate436inter4));
  nand2 gate930(.a(gate436inter4), .b(gate436inter3), .O(gate436inter5));
  nor2  gate931(.a(gate436inter5), .b(gate436inter2), .O(gate436inter6));
  inv1  gate932(.a(G1060), .O(gate436inter7));
  inv1  gate933(.a(G1156), .O(gate436inter8));
  nand2 gate934(.a(gate436inter8), .b(gate436inter7), .O(gate436inter9));
  nand2 gate935(.a(s_55), .b(gate436inter3), .O(gate436inter10));
  nor2  gate936(.a(gate436inter10), .b(gate436inter9), .O(gate436inter11));
  nor2  gate937(.a(gate436inter11), .b(gate436inter6), .O(gate436inter12));
  nand2 gate938(.a(gate436inter12), .b(gate436inter1), .O(G1245));
nand2 gate437( .a(G10), .b(G1159), .O(G1246) );
nand2 gate438( .a(G1063), .b(G1159), .O(G1247) );
nand2 gate439( .a(G11), .b(G1162), .O(G1248) );

  xor2  gate561(.a(G1162), .b(G1066), .O(gate440inter0));
  nand2 gate562(.a(gate440inter0), .b(s_2), .O(gate440inter1));
  and2  gate563(.a(G1162), .b(G1066), .O(gate440inter2));
  inv1  gate564(.a(s_2), .O(gate440inter3));
  inv1  gate565(.a(s_3), .O(gate440inter4));
  nand2 gate566(.a(gate440inter4), .b(gate440inter3), .O(gate440inter5));
  nor2  gate567(.a(gate440inter5), .b(gate440inter2), .O(gate440inter6));
  inv1  gate568(.a(G1066), .O(gate440inter7));
  inv1  gate569(.a(G1162), .O(gate440inter8));
  nand2 gate570(.a(gate440inter8), .b(gate440inter7), .O(gate440inter9));
  nand2 gate571(.a(s_3), .b(gate440inter3), .O(gate440inter10));
  nor2  gate572(.a(gate440inter10), .b(gate440inter9), .O(gate440inter11));
  nor2  gate573(.a(gate440inter11), .b(gate440inter6), .O(gate440inter12));
  nand2 gate574(.a(gate440inter12), .b(gate440inter1), .O(G1249));
nand2 gate441( .a(G12), .b(G1165), .O(G1250) );
nand2 gate442( .a(G1069), .b(G1165), .O(G1251) );

  xor2  gate799(.a(G1168), .b(G13), .O(gate443inter0));
  nand2 gate800(.a(gate443inter0), .b(s_36), .O(gate443inter1));
  and2  gate801(.a(G1168), .b(G13), .O(gate443inter2));
  inv1  gate802(.a(s_36), .O(gate443inter3));
  inv1  gate803(.a(s_37), .O(gate443inter4));
  nand2 gate804(.a(gate443inter4), .b(gate443inter3), .O(gate443inter5));
  nor2  gate805(.a(gate443inter5), .b(gate443inter2), .O(gate443inter6));
  inv1  gate806(.a(G13), .O(gate443inter7));
  inv1  gate807(.a(G1168), .O(gate443inter8));
  nand2 gate808(.a(gate443inter8), .b(gate443inter7), .O(gate443inter9));
  nand2 gate809(.a(s_37), .b(gate443inter3), .O(gate443inter10));
  nor2  gate810(.a(gate443inter10), .b(gate443inter9), .O(gate443inter11));
  nor2  gate811(.a(gate443inter11), .b(gate443inter6), .O(gate443inter12));
  nand2 gate812(.a(gate443inter12), .b(gate443inter1), .O(G1252));

  xor2  gate2689(.a(G1168), .b(G1072), .O(gate444inter0));
  nand2 gate2690(.a(gate444inter0), .b(s_306), .O(gate444inter1));
  and2  gate2691(.a(G1168), .b(G1072), .O(gate444inter2));
  inv1  gate2692(.a(s_306), .O(gate444inter3));
  inv1  gate2693(.a(s_307), .O(gate444inter4));
  nand2 gate2694(.a(gate444inter4), .b(gate444inter3), .O(gate444inter5));
  nor2  gate2695(.a(gate444inter5), .b(gate444inter2), .O(gate444inter6));
  inv1  gate2696(.a(G1072), .O(gate444inter7));
  inv1  gate2697(.a(G1168), .O(gate444inter8));
  nand2 gate2698(.a(gate444inter8), .b(gate444inter7), .O(gate444inter9));
  nand2 gate2699(.a(s_307), .b(gate444inter3), .O(gate444inter10));
  nor2  gate2700(.a(gate444inter10), .b(gate444inter9), .O(gate444inter11));
  nor2  gate2701(.a(gate444inter11), .b(gate444inter6), .O(gate444inter12));
  nand2 gate2702(.a(gate444inter12), .b(gate444inter1), .O(G1253));
nand2 gate445( .a(G14), .b(G1171), .O(G1254) );
nand2 gate446( .a(G1075), .b(G1171), .O(G1255) );
nand2 gate447( .a(G15), .b(G1174), .O(G1256) );
nand2 gate448( .a(G1078), .b(G1174), .O(G1257) );
nand2 gate449( .a(G16), .b(G1177), .O(G1258) );
nand2 gate450( .a(G1081), .b(G1177), .O(G1259) );

  xor2  gate687(.a(G1180), .b(G17), .O(gate451inter0));
  nand2 gate688(.a(gate451inter0), .b(s_20), .O(gate451inter1));
  and2  gate689(.a(G1180), .b(G17), .O(gate451inter2));
  inv1  gate690(.a(s_20), .O(gate451inter3));
  inv1  gate691(.a(s_21), .O(gate451inter4));
  nand2 gate692(.a(gate451inter4), .b(gate451inter3), .O(gate451inter5));
  nor2  gate693(.a(gate451inter5), .b(gate451inter2), .O(gate451inter6));
  inv1  gate694(.a(G17), .O(gate451inter7));
  inv1  gate695(.a(G1180), .O(gate451inter8));
  nand2 gate696(.a(gate451inter8), .b(gate451inter7), .O(gate451inter9));
  nand2 gate697(.a(s_21), .b(gate451inter3), .O(gate451inter10));
  nor2  gate698(.a(gate451inter10), .b(gate451inter9), .O(gate451inter11));
  nor2  gate699(.a(gate451inter11), .b(gate451inter6), .O(gate451inter12));
  nand2 gate700(.a(gate451inter12), .b(gate451inter1), .O(G1260));

  xor2  gate1877(.a(G1180), .b(G1084), .O(gate452inter0));
  nand2 gate1878(.a(gate452inter0), .b(s_190), .O(gate452inter1));
  and2  gate1879(.a(G1180), .b(G1084), .O(gate452inter2));
  inv1  gate1880(.a(s_190), .O(gate452inter3));
  inv1  gate1881(.a(s_191), .O(gate452inter4));
  nand2 gate1882(.a(gate452inter4), .b(gate452inter3), .O(gate452inter5));
  nor2  gate1883(.a(gate452inter5), .b(gate452inter2), .O(gate452inter6));
  inv1  gate1884(.a(G1084), .O(gate452inter7));
  inv1  gate1885(.a(G1180), .O(gate452inter8));
  nand2 gate1886(.a(gate452inter8), .b(gate452inter7), .O(gate452inter9));
  nand2 gate1887(.a(s_191), .b(gate452inter3), .O(gate452inter10));
  nor2  gate1888(.a(gate452inter10), .b(gate452inter9), .O(gate452inter11));
  nor2  gate1889(.a(gate452inter11), .b(gate452inter6), .O(gate452inter12));
  nand2 gate1890(.a(gate452inter12), .b(gate452inter1), .O(G1261));
nand2 gate453( .a(G18), .b(G1183), .O(G1262) );

  xor2  gate2423(.a(G1183), .b(G1087), .O(gate454inter0));
  nand2 gate2424(.a(gate454inter0), .b(s_268), .O(gate454inter1));
  and2  gate2425(.a(G1183), .b(G1087), .O(gate454inter2));
  inv1  gate2426(.a(s_268), .O(gate454inter3));
  inv1  gate2427(.a(s_269), .O(gate454inter4));
  nand2 gate2428(.a(gate454inter4), .b(gate454inter3), .O(gate454inter5));
  nor2  gate2429(.a(gate454inter5), .b(gate454inter2), .O(gate454inter6));
  inv1  gate2430(.a(G1087), .O(gate454inter7));
  inv1  gate2431(.a(G1183), .O(gate454inter8));
  nand2 gate2432(.a(gate454inter8), .b(gate454inter7), .O(gate454inter9));
  nand2 gate2433(.a(s_269), .b(gate454inter3), .O(gate454inter10));
  nor2  gate2434(.a(gate454inter10), .b(gate454inter9), .O(gate454inter11));
  nor2  gate2435(.a(gate454inter11), .b(gate454inter6), .O(gate454inter12));
  nand2 gate2436(.a(gate454inter12), .b(gate454inter1), .O(G1263));

  xor2  gate1919(.a(G1186), .b(G19), .O(gate455inter0));
  nand2 gate1920(.a(gate455inter0), .b(s_196), .O(gate455inter1));
  and2  gate1921(.a(G1186), .b(G19), .O(gate455inter2));
  inv1  gate1922(.a(s_196), .O(gate455inter3));
  inv1  gate1923(.a(s_197), .O(gate455inter4));
  nand2 gate1924(.a(gate455inter4), .b(gate455inter3), .O(gate455inter5));
  nor2  gate1925(.a(gate455inter5), .b(gate455inter2), .O(gate455inter6));
  inv1  gate1926(.a(G19), .O(gate455inter7));
  inv1  gate1927(.a(G1186), .O(gate455inter8));
  nand2 gate1928(.a(gate455inter8), .b(gate455inter7), .O(gate455inter9));
  nand2 gate1929(.a(s_197), .b(gate455inter3), .O(gate455inter10));
  nor2  gate1930(.a(gate455inter10), .b(gate455inter9), .O(gate455inter11));
  nor2  gate1931(.a(gate455inter11), .b(gate455inter6), .O(gate455inter12));
  nand2 gate1932(.a(gate455inter12), .b(gate455inter1), .O(G1264));
nand2 gate456( .a(G1090), .b(G1186), .O(G1265) );
nand2 gate457( .a(G20), .b(G1189), .O(G1266) );
nand2 gate458( .a(G1093), .b(G1189), .O(G1267) );
nand2 gate459( .a(G21), .b(G1192), .O(G1268) );

  xor2  gate1457(.a(G1192), .b(G1096), .O(gate460inter0));
  nand2 gate1458(.a(gate460inter0), .b(s_130), .O(gate460inter1));
  and2  gate1459(.a(G1192), .b(G1096), .O(gate460inter2));
  inv1  gate1460(.a(s_130), .O(gate460inter3));
  inv1  gate1461(.a(s_131), .O(gate460inter4));
  nand2 gate1462(.a(gate460inter4), .b(gate460inter3), .O(gate460inter5));
  nor2  gate1463(.a(gate460inter5), .b(gate460inter2), .O(gate460inter6));
  inv1  gate1464(.a(G1096), .O(gate460inter7));
  inv1  gate1465(.a(G1192), .O(gate460inter8));
  nand2 gate1466(.a(gate460inter8), .b(gate460inter7), .O(gate460inter9));
  nand2 gate1467(.a(s_131), .b(gate460inter3), .O(gate460inter10));
  nor2  gate1468(.a(gate460inter10), .b(gate460inter9), .O(gate460inter11));
  nor2  gate1469(.a(gate460inter11), .b(gate460inter6), .O(gate460inter12));
  nand2 gate1470(.a(gate460inter12), .b(gate460inter1), .O(G1269));

  xor2  gate2633(.a(G1195), .b(G22), .O(gate461inter0));
  nand2 gate2634(.a(gate461inter0), .b(s_298), .O(gate461inter1));
  and2  gate2635(.a(G1195), .b(G22), .O(gate461inter2));
  inv1  gate2636(.a(s_298), .O(gate461inter3));
  inv1  gate2637(.a(s_299), .O(gate461inter4));
  nand2 gate2638(.a(gate461inter4), .b(gate461inter3), .O(gate461inter5));
  nor2  gate2639(.a(gate461inter5), .b(gate461inter2), .O(gate461inter6));
  inv1  gate2640(.a(G22), .O(gate461inter7));
  inv1  gate2641(.a(G1195), .O(gate461inter8));
  nand2 gate2642(.a(gate461inter8), .b(gate461inter7), .O(gate461inter9));
  nand2 gate2643(.a(s_299), .b(gate461inter3), .O(gate461inter10));
  nor2  gate2644(.a(gate461inter10), .b(gate461inter9), .O(gate461inter11));
  nor2  gate2645(.a(gate461inter11), .b(gate461inter6), .O(gate461inter12));
  nand2 gate2646(.a(gate461inter12), .b(gate461inter1), .O(G1270));

  xor2  gate2871(.a(G1195), .b(G1099), .O(gate462inter0));
  nand2 gate2872(.a(gate462inter0), .b(s_332), .O(gate462inter1));
  and2  gate2873(.a(G1195), .b(G1099), .O(gate462inter2));
  inv1  gate2874(.a(s_332), .O(gate462inter3));
  inv1  gate2875(.a(s_333), .O(gate462inter4));
  nand2 gate2876(.a(gate462inter4), .b(gate462inter3), .O(gate462inter5));
  nor2  gate2877(.a(gate462inter5), .b(gate462inter2), .O(gate462inter6));
  inv1  gate2878(.a(G1099), .O(gate462inter7));
  inv1  gate2879(.a(G1195), .O(gate462inter8));
  nand2 gate2880(.a(gate462inter8), .b(gate462inter7), .O(gate462inter9));
  nand2 gate2881(.a(s_333), .b(gate462inter3), .O(gate462inter10));
  nor2  gate2882(.a(gate462inter10), .b(gate462inter9), .O(gate462inter11));
  nor2  gate2883(.a(gate462inter11), .b(gate462inter6), .O(gate462inter12));
  nand2 gate2884(.a(gate462inter12), .b(gate462inter1), .O(G1271));
nand2 gate463( .a(G23), .b(G1198), .O(G1272) );
nand2 gate464( .a(G1102), .b(G1198), .O(G1273) );

  xor2  gate1779(.a(G1201), .b(G24), .O(gate465inter0));
  nand2 gate1780(.a(gate465inter0), .b(s_176), .O(gate465inter1));
  and2  gate1781(.a(G1201), .b(G24), .O(gate465inter2));
  inv1  gate1782(.a(s_176), .O(gate465inter3));
  inv1  gate1783(.a(s_177), .O(gate465inter4));
  nand2 gate1784(.a(gate465inter4), .b(gate465inter3), .O(gate465inter5));
  nor2  gate1785(.a(gate465inter5), .b(gate465inter2), .O(gate465inter6));
  inv1  gate1786(.a(G24), .O(gate465inter7));
  inv1  gate1787(.a(G1201), .O(gate465inter8));
  nand2 gate1788(.a(gate465inter8), .b(gate465inter7), .O(gate465inter9));
  nand2 gate1789(.a(s_177), .b(gate465inter3), .O(gate465inter10));
  nor2  gate1790(.a(gate465inter10), .b(gate465inter9), .O(gate465inter11));
  nor2  gate1791(.a(gate465inter11), .b(gate465inter6), .O(gate465inter12));
  nand2 gate1792(.a(gate465inter12), .b(gate465inter1), .O(G1274));
nand2 gate466( .a(G1105), .b(G1201), .O(G1275) );

  xor2  gate1961(.a(G1204), .b(G25), .O(gate467inter0));
  nand2 gate1962(.a(gate467inter0), .b(s_202), .O(gate467inter1));
  and2  gate1963(.a(G1204), .b(G25), .O(gate467inter2));
  inv1  gate1964(.a(s_202), .O(gate467inter3));
  inv1  gate1965(.a(s_203), .O(gate467inter4));
  nand2 gate1966(.a(gate467inter4), .b(gate467inter3), .O(gate467inter5));
  nor2  gate1967(.a(gate467inter5), .b(gate467inter2), .O(gate467inter6));
  inv1  gate1968(.a(G25), .O(gate467inter7));
  inv1  gate1969(.a(G1204), .O(gate467inter8));
  nand2 gate1970(.a(gate467inter8), .b(gate467inter7), .O(gate467inter9));
  nand2 gate1971(.a(s_203), .b(gate467inter3), .O(gate467inter10));
  nor2  gate1972(.a(gate467inter10), .b(gate467inter9), .O(gate467inter11));
  nor2  gate1973(.a(gate467inter11), .b(gate467inter6), .O(gate467inter12));
  nand2 gate1974(.a(gate467inter12), .b(gate467inter1), .O(G1276));
nand2 gate468( .a(G1108), .b(G1204), .O(G1277) );

  xor2  gate589(.a(G1207), .b(G26), .O(gate469inter0));
  nand2 gate590(.a(gate469inter0), .b(s_6), .O(gate469inter1));
  and2  gate591(.a(G1207), .b(G26), .O(gate469inter2));
  inv1  gate592(.a(s_6), .O(gate469inter3));
  inv1  gate593(.a(s_7), .O(gate469inter4));
  nand2 gate594(.a(gate469inter4), .b(gate469inter3), .O(gate469inter5));
  nor2  gate595(.a(gate469inter5), .b(gate469inter2), .O(gate469inter6));
  inv1  gate596(.a(G26), .O(gate469inter7));
  inv1  gate597(.a(G1207), .O(gate469inter8));
  nand2 gate598(.a(gate469inter8), .b(gate469inter7), .O(gate469inter9));
  nand2 gate599(.a(s_7), .b(gate469inter3), .O(gate469inter10));
  nor2  gate600(.a(gate469inter10), .b(gate469inter9), .O(gate469inter11));
  nor2  gate601(.a(gate469inter11), .b(gate469inter6), .O(gate469inter12));
  nand2 gate602(.a(gate469inter12), .b(gate469inter1), .O(G1278));
nand2 gate470( .a(G1111), .b(G1207), .O(G1279) );
nand2 gate471( .a(G27), .b(G1210), .O(G1280) );
nand2 gate472( .a(G1114), .b(G1210), .O(G1281) );
nand2 gate473( .a(G28), .b(G1213), .O(G1282) );
nand2 gate474( .a(G1117), .b(G1213), .O(G1283) );
nand2 gate475( .a(G29), .b(G1216), .O(G1284) );
nand2 gate476( .a(G1120), .b(G1216), .O(G1285) );

  xor2  gate2367(.a(G1219), .b(G30), .O(gate477inter0));
  nand2 gate2368(.a(gate477inter0), .b(s_260), .O(gate477inter1));
  and2  gate2369(.a(G1219), .b(G30), .O(gate477inter2));
  inv1  gate2370(.a(s_260), .O(gate477inter3));
  inv1  gate2371(.a(s_261), .O(gate477inter4));
  nand2 gate2372(.a(gate477inter4), .b(gate477inter3), .O(gate477inter5));
  nor2  gate2373(.a(gate477inter5), .b(gate477inter2), .O(gate477inter6));
  inv1  gate2374(.a(G30), .O(gate477inter7));
  inv1  gate2375(.a(G1219), .O(gate477inter8));
  nand2 gate2376(.a(gate477inter8), .b(gate477inter7), .O(gate477inter9));
  nand2 gate2377(.a(s_261), .b(gate477inter3), .O(gate477inter10));
  nor2  gate2378(.a(gate477inter10), .b(gate477inter9), .O(gate477inter11));
  nor2  gate2379(.a(gate477inter11), .b(gate477inter6), .O(gate477inter12));
  nand2 gate2380(.a(gate477inter12), .b(gate477inter1), .O(G1286));
nand2 gate478( .a(G1123), .b(G1219), .O(G1287) );

  xor2  gate2087(.a(G1222), .b(G31), .O(gate479inter0));
  nand2 gate2088(.a(gate479inter0), .b(s_220), .O(gate479inter1));
  and2  gate2089(.a(G1222), .b(G31), .O(gate479inter2));
  inv1  gate2090(.a(s_220), .O(gate479inter3));
  inv1  gate2091(.a(s_221), .O(gate479inter4));
  nand2 gate2092(.a(gate479inter4), .b(gate479inter3), .O(gate479inter5));
  nor2  gate2093(.a(gate479inter5), .b(gate479inter2), .O(gate479inter6));
  inv1  gate2094(.a(G31), .O(gate479inter7));
  inv1  gate2095(.a(G1222), .O(gate479inter8));
  nand2 gate2096(.a(gate479inter8), .b(gate479inter7), .O(gate479inter9));
  nand2 gate2097(.a(s_221), .b(gate479inter3), .O(gate479inter10));
  nor2  gate2098(.a(gate479inter10), .b(gate479inter9), .O(gate479inter11));
  nor2  gate2099(.a(gate479inter11), .b(gate479inter6), .O(gate479inter12));
  nand2 gate2100(.a(gate479inter12), .b(gate479inter1), .O(G1288));

  xor2  gate2955(.a(G1222), .b(G1126), .O(gate480inter0));
  nand2 gate2956(.a(gate480inter0), .b(s_344), .O(gate480inter1));
  and2  gate2957(.a(G1222), .b(G1126), .O(gate480inter2));
  inv1  gate2958(.a(s_344), .O(gate480inter3));
  inv1  gate2959(.a(s_345), .O(gate480inter4));
  nand2 gate2960(.a(gate480inter4), .b(gate480inter3), .O(gate480inter5));
  nor2  gate2961(.a(gate480inter5), .b(gate480inter2), .O(gate480inter6));
  inv1  gate2962(.a(G1126), .O(gate480inter7));
  inv1  gate2963(.a(G1222), .O(gate480inter8));
  nand2 gate2964(.a(gate480inter8), .b(gate480inter7), .O(gate480inter9));
  nand2 gate2965(.a(s_345), .b(gate480inter3), .O(gate480inter10));
  nor2  gate2966(.a(gate480inter10), .b(gate480inter9), .O(gate480inter11));
  nor2  gate2967(.a(gate480inter11), .b(gate480inter6), .O(gate480inter12));
  nand2 gate2968(.a(gate480inter12), .b(gate480inter1), .O(G1289));
nand2 gate481( .a(G32), .b(G1225), .O(G1290) );

  xor2  gate2549(.a(G1225), .b(G1129), .O(gate482inter0));
  nand2 gate2550(.a(gate482inter0), .b(s_286), .O(gate482inter1));
  and2  gate2551(.a(G1225), .b(G1129), .O(gate482inter2));
  inv1  gate2552(.a(s_286), .O(gate482inter3));
  inv1  gate2553(.a(s_287), .O(gate482inter4));
  nand2 gate2554(.a(gate482inter4), .b(gate482inter3), .O(gate482inter5));
  nor2  gate2555(.a(gate482inter5), .b(gate482inter2), .O(gate482inter6));
  inv1  gate2556(.a(G1129), .O(gate482inter7));
  inv1  gate2557(.a(G1225), .O(gate482inter8));
  nand2 gate2558(.a(gate482inter8), .b(gate482inter7), .O(gate482inter9));
  nand2 gate2559(.a(s_287), .b(gate482inter3), .O(gate482inter10));
  nor2  gate2560(.a(gate482inter10), .b(gate482inter9), .O(gate482inter11));
  nor2  gate2561(.a(gate482inter11), .b(gate482inter6), .O(gate482inter12));
  nand2 gate2562(.a(gate482inter12), .b(gate482inter1), .O(G1291));
nand2 gate483( .a(G1228), .b(G1229), .O(G1292) );

  xor2  gate1527(.a(G1231), .b(G1230), .O(gate484inter0));
  nand2 gate1528(.a(gate484inter0), .b(s_140), .O(gate484inter1));
  and2  gate1529(.a(G1231), .b(G1230), .O(gate484inter2));
  inv1  gate1530(.a(s_140), .O(gate484inter3));
  inv1  gate1531(.a(s_141), .O(gate484inter4));
  nand2 gate1532(.a(gate484inter4), .b(gate484inter3), .O(gate484inter5));
  nor2  gate1533(.a(gate484inter5), .b(gate484inter2), .O(gate484inter6));
  inv1  gate1534(.a(G1230), .O(gate484inter7));
  inv1  gate1535(.a(G1231), .O(gate484inter8));
  nand2 gate1536(.a(gate484inter8), .b(gate484inter7), .O(gate484inter9));
  nand2 gate1537(.a(s_141), .b(gate484inter3), .O(gate484inter10));
  nor2  gate1538(.a(gate484inter10), .b(gate484inter9), .O(gate484inter11));
  nor2  gate1539(.a(gate484inter11), .b(gate484inter6), .O(gate484inter12));
  nand2 gate1540(.a(gate484inter12), .b(gate484inter1), .O(G1293));
nand2 gate485( .a(G1232), .b(G1233), .O(G1294) );
nand2 gate486( .a(G1234), .b(G1235), .O(G1295) );
nand2 gate487( .a(G1236), .b(G1237), .O(G1296) );
nand2 gate488( .a(G1238), .b(G1239), .O(G1297) );

  xor2  gate575(.a(G1241), .b(G1240), .O(gate489inter0));
  nand2 gate576(.a(gate489inter0), .b(s_4), .O(gate489inter1));
  and2  gate577(.a(G1241), .b(G1240), .O(gate489inter2));
  inv1  gate578(.a(s_4), .O(gate489inter3));
  inv1  gate579(.a(s_5), .O(gate489inter4));
  nand2 gate580(.a(gate489inter4), .b(gate489inter3), .O(gate489inter5));
  nor2  gate581(.a(gate489inter5), .b(gate489inter2), .O(gate489inter6));
  inv1  gate582(.a(G1240), .O(gate489inter7));
  inv1  gate583(.a(G1241), .O(gate489inter8));
  nand2 gate584(.a(gate489inter8), .b(gate489inter7), .O(gate489inter9));
  nand2 gate585(.a(s_5), .b(gate489inter3), .O(gate489inter10));
  nor2  gate586(.a(gate489inter10), .b(gate489inter9), .O(gate489inter11));
  nor2  gate587(.a(gate489inter11), .b(gate489inter6), .O(gate489inter12));
  nand2 gate588(.a(gate489inter12), .b(gate489inter1), .O(G1298));
nand2 gate490( .a(G1242), .b(G1243), .O(G1299) );
nand2 gate491( .a(G1244), .b(G1245), .O(G1300) );

  xor2  gate1863(.a(G1247), .b(G1246), .O(gate492inter0));
  nand2 gate1864(.a(gate492inter0), .b(s_188), .O(gate492inter1));
  and2  gate1865(.a(G1247), .b(G1246), .O(gate492inter2));
  inv1  gate1866(.a(s_188), .O(gate492inter3));
  inv1  gate1867(.a(s_189), .O(gate492inter4));
  nand2 gate1868(.a(gate492inter4), .b(gate492inter3), .O(gate492inter5));
  nor2  gate1869(.a(gate492inter5), .b(gate492inter2), .O(gate492inter6));
  inv1  gate1870(.a(G1246), .O(gate492inter7));
  inv1  gate1871(.a(G1247), .O(gate492inter8));
  nand2 gate1872(.a(gate492inter8), .b(gate492inter7), .O(gate492inter9));
  nand2 gate1873(.a(s_189), .b(gate492inter3), .O(gate492inter10));
  nor2  gate1874(.a(gate492inter10), .b(gate492inter9), .O(gate492inter11));
  nor2  gate1875(.a(gate492inter11), .b(gate492inter6), .O(gate492inter12));
  nand2 gate1876(.a(gate492inter12), .b(gate492inter1), .O(G1301));
nand2 gate493( .a(G1248), .b(G1249), .O(G1302) );
nand2 gate494( .a(G1250), .b(G1251), .O(G1303) );
nand2 gate495( .a(G1252), .b(G1253), .O(G1304) );
nand2 gate496( .a(G1254), .b(G1255), .O(G1305) );

  xor2  gate1681(.a(G1257), .b(G1256), .O(gate497inter0));
  nand2 gate1682(.a(gate497inter0), .b(s_162), .O(gate497inter1));
  and2  gate1683(.a(G1257), .b(G1256), .O(gate497inter2));
  inv1  gate1684(.a(s_162), .O(gate497inter3));
  inv1  gate1685(.a(s_163), .O(gate497inter4));
  nand2 gate1686(.a(gate497inter4), .b(gate497inter3), .O(gate497inter5));
  nor2  gate1687(.a(gate497inter5), .b(gate497inter2), .O(gate497inter6));
  inv1  gate1688(.a(G1256), .O(gate497inter7));
  inv1  gate1689(.a(G1257), .O(gate497inter8));
  nand2 gate1690(.a(gate497inter8), .b(gate497inter7), .O(gate497inter9));
  nand2 gate1691(.a(s_163), .b(gate497inter3), .O(gate497inter10));
  nor2  gate1692(.a(gate497inter10), .b(gate497inter9), .O(gate497inter11));
  nor2  gate1693(.a(gate497inter11), .b(gate497inter6), .O(gate497inter12));
  nand2 gate1694(.a(gate497inter12), .b(gate497inter1), .O(G1306));
nand2 gate498( .a(G1258), .b(G1259), .O(G1307) );
nand2 gate499( .a(G1260), .b(G1261), .O(G1308) );

  xor2  gate1205(.a(G1263), .b(G1262), .O(gate500inter0));
  nand2 gate1206(.a(gate500inter0), .b(s_94), .O(gate500inter1));
  and2  gate1207(.a(G1263), .b(G1262), .O(gate500inter2));
  inv1  gate1208(.a(s_94), .O(gate500inter3));
  inv1  gate1209(.a(s_95), .O(gate500inter4));
  nand2 gate1210(.a(gate500inter4), .b(gate500inter3), .O(gate500inter5));
  nor2  gate1211(.a(gate500inter5), .b(gate500inter2), .O(gate500inter6));
  inv1  gate1212(.a(G1262), .O(gate500inter7));
  inv1  gate1213(.a(G1263), .O(gate500inter8));
  nand2 gate1214(.a(gate500inter8), .b(gate500inter7), .O(gate500inter9));
  nand2 gate1215(.a(s_95), .b(gate500inter3), .O(gate500inter10));
  nor2  gate1216(.a(gate500inter10), .b(gate500inter9), .O(gate500inter11));
  nor2  gate1217(.a(gate500inter11), .b(gate500inter6), .O(gate500inter12));
  nand2 gate1218(.a(gate500inter12), .b(gate500inter1), .O(G1309));
nand2 gate501( .a(G1264), .b(G1265), .O(G1310) );
nand2 gate502( .a(G1266), .b(G1267), .O(G1311) );

  xor2  gate2773(.a(G1269), .b(G1268), .O(gate503inter0));
  nand2 gate2774(.a(gate503inter0), .b(s_318), .O(gate503inter1));
  and2  gate2775(.a(G1269), .b(G1268), .O(gate503inter2));
  inv1  gate2776(.a(s_318), .O(gate503inter3));
  inv1  gate2777(.a(s_319), .O(gate503inter4));
  nand2 gate2778(.a(gate503inter4), .b(gate503inter3), .O(gate503inter5));
  nor2  gate2779(.a(gate503inter5), .b(gate503inter2), .O(gate503inter6));
  inv1  gate2780(.a(G1268), .O(gate503inter7));
  inv1  gate2781(.a(G1269), .O(gate503inter8));
  nand2 gate2782(.a(gate503inter8), .b(gate503inter7), .O(gate503inter9));
  nand2 gate2783(.a(s_319), .b(gate503inter3), .O(gate503inter10));
  nor2  gate2784(.a(gate503inter10), .b(gate503inter9), .O(gate503inter11));
  nor2  gate2785(.a(gate503inter11), .b(gate503inter6), .O(gate503inter12));
  nand2 gate2786(.a(gate503inter12), .b(gate503inter1), .O(G1312));

  xor2  gate2101(.a(G1271), .b(G1270), .O(gate504inter0));
  nand2 gate2102(.a(gate504inter0), .b(s_222), .O(gate504inter1));
  and2  gate2103(.a(G1271), .b(G1270), .O(gate504inter2));
  inv1  gate2104(.a(s_222), .O(gate504inter3));
  inv1  gate2105(.a(s_223), .O(gate504inter4));
  nand2 gate2106(.a(gate504inter4), .b(gate504inter3), .O(gate504inter5));
  nor2  gate2107(.a(gate504inter5), .b(gate504inter2), .O(gate504inter6));
  inv1  gate2108(.a(G1270), .O(gate504inter7));
  inv1  gate2109(.a(G1271), .O(gate504inter8));
  nand2 gate2110(.a(gate504inter8), .b(gate504inter7), .O(gate504inter9));
  nand2 gate2111(.a(s_223), .b(gate504inter3), .O(gate504inter10));
  nor2  gate2112(.a(gate504inter10), .b(gate504inter9), .O(gate504inter11));
  nor2  gate2113(.a(gate504inter11), .b(gate504inter6), .O(gate504inter12));
  nand2 gate2114(.a(gate504inter12), .b(gate504inter1), .O(G1313));
nand2 gate505( .a(G1272), .b(G1273), .O(G1314) );

  xor2  gate1583(.a(G1275), .b(G1274), .O(gate506inter0));
  nand2 gate1584(.a(gate506inter0), .b(s_148), .O(gate506inter1));
  and2  gate1585(.a(G1275), .b(G1274), .O(gate506inter2));
  inv1  gate1586(.a(s_148), .O(gate506inter3));
  inv1  gate1587(.a(s_149), .O(gate506inter4));
  nand2 gate1588(.a(gate506inter4), .b(gate506inter3), .O(gate506inter5));
  nor2  gate1589(.a(gate506inter5), .b(gate506inter2), .O(gate506inter6));
  inv1  gate1590(.a(G1274), .O(gate506inter7));
  inv1  gate1591(.a(G1275), .O(gate506inter8));
  nand2 gate1592(.a(gate506inter8), .b(gate506inter7), .O(gate506inter9));
  nand2 gate1593(.a(s_149), .b(gate506inter3), .O(gate506inter10));
  nor2  gate1594(.a(gate506inter10), .b(gate506inter9), .O(gate506inter11));
  nor2  gate1595(.a(gate506inter11), .b(gate506inter6), .O(gate506inter12));
  nand2 gate1596(.a(gate506inter12), .b(gate506inter1), .O(G1315));
nand2 gate507( .a(G1276), .b(G1277), .O(G1316) );
nand2 gate508( .a(G1278), .b(G1279), .O(G1317) );

  xor2  gate2227(.a(G1281), .b(G1280), .O(gate509inter0));
  nand2 gate2228(.a(gate509inter0), .b(s_240), .O(gate509inter1));
  and2  gate2229(.a(G1281), .b(G1280), .O(gate509inter2));
  inv1  gate2230(.a(s_240), .O(gate509inter3));
  inv1  gate2231(.a(s_241), .O(gate509inter4));
  nand2 gate2232(.a(gate509inter4), .b(gate509inter3), .O(gate509inter5));
  nor2  gate2233(.a(gate509inter5), .b(gate509inter2), .O(gate509inter6));
  inv1  gate2234(.a(G1280), .O(gate509inter7));
  inv1  gate2235(.a(G1281), .O(gate509inter8));
  nand2 gate2236(.a(gate509inter8), .b(gate509inter7), .O(gate509inter9));
  nand2 gate2237(.a(s_241), .b(gate509inter3), .O(gate509inter10));
  nor2  gate2238(.a(gate509inter10), .b(gate509inter9), .O(gate509inter11));
  nor2  gate2239(.a(gate509inter11), .b(gate509inter6), .O(gate509inter12));
  nand2 gate2240(.a(gate509inter12), .b(gate509inter1), .O(G1318));
nand2 gate510( .a(G1282), .b(G1283), .O(G1319) );
nand2 gate511( .a(G1284), .b(G1285), .O(G1320) );

  xor2  gate1163(.a(G1287), .b(G1286), .O(gate512inter0));
  nand2 gate1164(.a(gate512inter0), .b(s_88), .O(gate512inter1));
  and2  gate1165(.a(G1287), .b(G1286), .O(gate512inter2));
  inv1  gate1166(.a(s_88), .O(gate512inter3));
  inv1  gate1167(.a(s_89), .O(gate512inter4));
  nand2 gate1168(.a(gate512inter4), .b(gate512inter3), .O(gate512inter5));
  nor2  gate1169(.a(gate512inter5), .b(gate512inter2), .O(gate512inter6));
  inv1  gate1170(.a(G1286), .O(gate512inter7));
  inv1  gate1171(.a(G1287), .O(gate512inter8));
  nand2 gate1172(.a(gate512inter8), .b(gate512inter7), .O(gate512inter9));
  nand2 gate1173(.a(s_89), .b(gate512inter3), .O(gate512inter10));
  nor2  gate1174(.a(gate512inter10), .b(gate512inter9), .O(gate512inter11));
  nor2  gate1175(.a(gate512inter11), .b(gate512inter6), .O(gate512inter12));
  nand2 gate1176(.a(gate512inter12), .b(gate512inter1), .O(G1321));

  xor2  gate2927(.a(G1289), .b(G1288), .O(gate513inter0));
  nand2 gate2928(.a(gate513inter0), .b(s_340), .O(gate513inter1));
  and2  gate2929(.a(G1289), .b(G1288), .O(gate513inter2));
  inv1  gate2930(.a(s_340), .O(gate513inter3));
  inv1  gate2931(.a(s_341), .O(gate513inter4));
  nand2 gate2932(.a(gate513inter4), .b(gate513inter3), .O(gate513inter5));
  nor2  gate2933(.a(gate513inter5), .b(gate513inter2), .O(gate513inter6));
  inv1  gate2934(.a(G1288), .O(gate513inter7));
  inv1  gate2935(.a(G1289), .O(gate513inter8));
  nand2 gate2936(.a(gate513inter8), .b(gate513inter7), .O(gate513inter9));
  nand2 gate2937(.a(s_341), .b(gate513inter3), .O(gate513inter10));
  nor2  gate2938(.a(gate513inter10), .b(gate513inter9), .O(gate513inter11));
  nor2  gate2939(.a(gate513inter11), .b(gate513inter6), .O(gate513inter12));
  nand2 gate2940(.a(gate513inter12), .b(gate513inter1), .O(G1322));
nand2 gate514( .a(G1290), .b(G1291), .O(G1323) );
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule