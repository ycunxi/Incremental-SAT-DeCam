module c499 (N1,N5,N9,N13,N17,N21,N25,N29,N33,N37,
             N41,N45,N49,N53,N57,N61,N65,N69,N73,N77,
             N81,N85,N89,N93,N97,N101,N105,N109,N113,N117,
             N121,N125,N129,N130,N131,N132,N133,N134,N135,N136,
             N137,N724,N725,N726,N727,N728,N729,N730,N731,N732,
             N733,N734,N735,N736,N737,N738,N739,N740,N741,N742,
             N743,N744,N745,N746,N747,N748,N749,N750,N751,N752,
             N753,N754,N755);

input N1,N5,N9,N13,N17,N21,N25,N29,N33,N37,
      N41,N45,N49,N53,N57,N61,N65,N69,N73,N77,
      N81,N85,N89,N93,N97,N101,N105,N109,N113,N117,
      N121,N125,N129,N130,N131,N132,N133,N134,N135,N136,
      N137;//RE__PI;

input s_0,s_1;//RE__ALLOW(00,01,10,11);
input s_2,s_3;//RE__ALLOW(00,01,10,11);
input s_4,s_5;//RE__ALLOW(00,01,10,11);
input s_6,s_7;//RE__ALLOW(00,01,10,11);
input s_8,s_9;//RE__ALLOW(00,01,10,11);
input s_10,s_11;//RE__ALLOW(00,01,10,11);
input s_12,s_13;//RE__ALLOW(00,01,10,11);
input s_14,s_15;//RE__ALLOW(00,01,10,11);
input s_16,s_17;//RE__ALLOW(00,01,10,11);
input s_18,s_19;//RE__ALLOW(00,01,10,11);
input s_20,s_21;//RE__ALLOW(00,01,10,11);
input s_22,s_23;//RE__ALLOW(00,01,10,11);
input s_24,s_25;//RE__ALLOW(00,01,10,11);
input s_26,s_27;//RE__ALLOW(00,01,10,11);
input s_28,s_29;//RE__ALLOW(00,01,10,11);
input s_30,s_31;//RE__ALLOW(00,01,10,11);
input s_32,s_33;//RE__ALLOW(00,01,10,11);
input s_34,s_35;//RE__ALLOW(00,01,10,11);
input s_36,s_37;//RE__ALLOW(00,01,10,11);
input s_38,s_39;//RE__ALLOW(00,01,10,11);
input s_40,s_41;//RE__ALLOW(00,01,10,11);
output N724,N725,N726,N727,N728,N729,N730,N731,N732,N733,
       N734,N735,N736,N737,N738,N739,N740,N741,N742,N743,
       N744,N745,N746,N747,N748,N749,N750,N751,N752,N753,
       N754,N755;

wire N250,N251,N252,N253,N254,N255,N256,N257,N258,N259,
     N260,N261,N262,N263,N264,N265,N266,N267,N268,N269,
     N270,N271,N272,N273,N274,N275,N276,N277,N278,N279,
     N280,N281,N282,N283,N284,N285,N286,N287,N288,N289,
     N290,N293,N296,N299,N302,N305,N308,N311,N314,N315,
     N316,N317,N318,N319,N320,N321,N338,N339,N340,N341,
     N342,N343,N344,N345,N346,N347,N348,N349,N350,N351,
     N352,N353,N354,N367,N380,N393,N406,N419,N432,N445,
     N554,N555,N556,N557,N558,N559,N560,N561,N562,N563,
     N564,N565,N566,N567,N568,N569,N570,N571,N572,N573,
     N574,N575,N576,N577,N578,N579,N580,N581,N582,N583,
     N584,N585,N586,N587,N588,N589,N590,N591,N592,N593,
     N594,N595,N596,N597,N598,N599,N600,N601,N602,N607,
     N620,N625,N630,N635,N640,N645,N650,N655,N692,N693,
     N694,N695,N696,N697,N698,N699,N700,N701,N702,N703,
     N704,N705,N706,N707,N708,N709,N710,N711,N712,N713,
     N714,N715,N716,N717,N718,N719,N720,N721,N722,N723, gate188inter0, gate188inter1, gate188inter2, gate188inter3, gate188inter4, gate188inter5, gate188inter6, gate188inter7, gate188inter8, gate188inter9, gate188inter10, gate188inter11, gate188inter12, gate187inter0, gate187inter1, gate187inter2, gate187inter3, gate187inter4, gate187inter5, gate187inter6, gate187inter7, gate187inter8, gate187inter9, gate187inter10, gate187inter11, gate187inter12, gate196inter0, gate196inter1, gate196inter2, gate196inter3, gate196inter4, gate196inter5, gate196inter6, gate196inter7, gate196inter8, gate196inter9, gate196inter10, gate196inter11, gate196inter12, gate64inter0, gate64inter1, gate64inter2, gate64inter3, gate64inter4, gate64inter5, gate64inter6, gate64inter7, gate64inter8, gate64inter9, gate64inter10, gate64inter11, gate64inter12, gate36inter0, gate36inter1, gate36inter2, gate36inter3, gate36inter4, gate36inter5, gate36inter6, gate36inter7, gate36inter8, gate36inter9, gate36inter10, gate36inter11, gate36inter12, gate172inter0, gate172inter1, gate172inter2, gate172inter3, gate172inter4, gate172inter5, gate172inter6, gate172inter7, gate172inter8, gate172inter9, gate172inter10, gate172inter11, gate172inter12, gate26inter0, gate26inter1, gate26inter2, gate26inter3, gate26inter4, gate26inter5, gate26inter6, gate26inter7, gate26inter8, gate26inter9, gate26inter10, gate26inter11, gate26inter12, gate10inter0, gate10inter1, gate10inter2, gate10inter3, gate10inter4, gate10inter5, gate10inter6, gate10inter7, gate10inter8, gate10inter9, gate10inter10, gate10inter11, gate10inter12, gate201inter0, gate201inter1, gate201inter2, gate201inter3, gate201inter4, gate201inter5, gate201inter6, gate201inter7, gate201inter8, gate201inter9, gate201inter10, gate201inter11, gate201inter12, gate190inter0, gate190inter1, gate190inter2, gate190inter3, gate190inter4, gate190inter5, gate190inter6, gate190inter7, gate190inter8, gate190inter9, gate190inter10, gate190inter11, gate190inter12, gate70inter0, gate70inter1, gate70inter2, gate70inter3, gate70inter4, gate70inter5, gate70inter6, gate70inter7, gate70inter8, gate70inter9, gate70inter10, gate70inter11, gate70inter12, gate25inter0, gate25inter1, gate25inter2, gate25inter3, gate25inter4, gate25inter5, gate25inter6, gate25inter7, gate25inter8, gate25inter9, gate25inter10, gate25inter11, gate25inter12, gate42inter0, gate42inter1, gate42inter2, gate42inter3, gate42inter4, gate42inter5, gate42inter6, gate42inter7, gate42inter8, gate42inter9, gate42inter10, gate42inter11, gate42inter12, gate198inter0, gate198inter1, gate198inter2, gate198inter3, gate198inter4, gate198inter5, gate198inter6, gate198inter7, gate198inter8, gate198inter9, gate198inter10, gate198inter11, gate198inter12, gate69inter0, gate69inter1, gate69inter2, gate69inter3, gate69inter4, gate69inter5, gate69inter6, gate69inter7, gate69inter8, gate69inter9, gate69inter10, gate69inter11, gate69inter12, gate71inter0, gate71inter1, gate71inter2, gate71inter3, gate71inter4, gate71inter5, gate71inter6, gate71inter7, gate71inter8, gate71inter9, gate71inter10, gate71inter11, gate71inter12, gate58inter0, gate58inter1, gate58inter2, gate58inter3, gate58inter4, gate58inter5, gate58inter6, gate58inter7, gate58inter8, gate58inter9, gate58inter10, gate58inter11, gate58inter12, gate54inter0, gate54inter1, gate54inter2, gate54inter3, gate54inter4, gate54inter5, gate54inter6, gate54inter7, gate54inter8, gate54inter9, gate54inter10, gate54inter11, gate54inter12, gate61inter0, gate61inter1, gate61inter2, gate61inter3, gate61inter4, gate61inter5, gate61inter6, gate61inter7, gate61inter8, gate61inter9, gate61inter10, gate61inter11, gate61inter12, gate33inter0, gate33inter1, gate33inter2, gate33inter3, gate33inter4, gate33inter5, gate33inter6, gate33inter7, gate33inter8, gate33inter9, gate33inter10, gate33inter11, gate33inter12, gate80inter0, gate80inter1, gate80inter2, gate80inter3, gate80inter4, gate80inter5, gate80inter6, gate80inter7, gate80inter8, gate80inter9, gate80inter10, gate80inter11, gate80inter12;



xor2 gate1( .a(N1), .b(N5), .O(N250) );
xor2 gate2( .a(N9), .b(N13), .O(N251) );
xor2 gate3( .a(N17), .b(N21), .O(N252) );
xor2 gate4( .a(N25), .b(N29), .O(N253) );
xor2 gate5( .a(N33), .b(N37), .O(N254) );
xor2 gate6( .a(N41), .b(N45), .O(N255) );
xor2 gate7( .a(N49), .b(N53), .O(N256) );
xor2 gate8( .a(N57), .b(N61), .O(N257) );
xor2 gate9( .a(N65), .b(N69), .O(N258) );

  xor2  gate301(.a(N77), .b(N73), .O(gate10inter0));
  nand2 gate302(.a(gate10inter0), .b(s_14), .O(gate10inter1));
  and2  gate303(.a(N77), .b(N73), .O(gate10inter2));
  inv1  gate304(.a(s_14), .O(gate10inter3));
  inv1  gate305(.a(s_15), .O(gate10inter4));
  nand2 gate306(.a(gate10inter4), .b(gate10inter3), .O(gate10inter5));
  nor2  gate307(.a(gate10inter5), .b(gate10inter2), .O(gate10inter6));
  inv1  gate308(.a(N73), .O(gate10inter7));
  inv1  gate309(.a(N77), .O(gate10inter8));
  nand2 gate310(.a(gate10inter8), .b(gate10inter7), .O(gate10inter9));
  nand2 gate311(.a(s_15), .b(gate10inter3), .O(gate10inter10));
  nor2  gate312(.a(gate10inter10), .b(gate10inter9), .O(gate10inter11));
  nor2  gate313(.a(gate10inter11), .b(gate10inter6), .O(gate10inter12));
  nand2 gate314(.a(gate10inter12), .b(gate10inter1), .O(N259));
xor2 gate11( .a(N81), .b(N85), .O(N260) );
xor2 gate12( .a(N89), .b(N93), .O(N261) );
xor2 gate13( .a(N97), .b(N101), .O(N262) );
xor2 gate14( .a(N105), .b(N109), .O(N263) );
xor2 gate15( .a(N113), .b(N117), .O(N264) );
xor2 gate16( .a(N121), .b(N125), .O(N265) );
and2 gate17( .a(N129), .b(N137), .O(N266) );
and2 gate18( .a(N130), .b(N137), .O(N267) );
and2 gate19( .a(N131), .b(N137), .O(N268) );
and2 gate20( .a(N132), .b(N137), .O(N269) );
and2 gate21( .a(N133), .b(N137), .O(N270) );
and2 gate22( .a(N134), .b(N137), .O(N271) );
and2 gate23( .a(N135), .b(N137), .O(N272) );
and2 gate24( .a(N136), .b(N137), .O(N273) );

  xor2  gate357(.a(N17), .b(N1), .O(gate25inter0));
  nand2 gate358(.a(gate25inter0), .b(s_22), .O(gate25inter1));
  and2  gate359(.a(N17), .b(N1), .O(gate25inter2));
  inv1  gate360(.a(s_22), .O(gate25inter3));
  inv1  gate361(.a(s_23), .O(gate25inter4));
  nand2 gate362(.a(gate25inter4), .b(gate25inter3), .O(gate25inter5));
  nor2  gate363(.a(gate25inter5), .b(gate25inter2), .O(gate25inter6));
  inv1  gate364(.a(N1), .O(gate25inter7));
  inv1  gate365(.a(N17), .O(gate25inter8));
  nand2 gate366(.a(gate25inter8), .b(gate25inter7), .O(gate25inter9));
  nand2 gate367(.a(s_23), .b(gate25inter3), .O(gate25inter10));
  nor2  gate368(.a(gate25inter10), .b(gate25inter9), .O(gate25inter11));
  nor2  gate369(.a(gate25inter11), .b(gate25inter6), .O(gate25inter12));
  nand2 gate370(.a(gate25inter12), .b(gate25inter1), .O(N274));

  xor2  gate287(.a(N49), .b(N33), .O(gate26inter0));
  nand2 gate288(.a(gate26inter0), .b(s_12), .O(gate26inter1));
  and2  gate289(.a(N49), .b(N33), .O(gate26inter2));
  inv1  gate290(.a(s_12), .O(gate26inter3));
  inv1  gate291(.a(s_13), .O(gate26inter4));
  nand2 gate292(.a(gate26inter4), .b(gate26inter3), .O(gate26inter5));
  nor2  gate293(.a(gate26inter5), .b(gate26inter2), .O(gate26inter6));
  inv1  gate294(.a(N33), .O(gate26inter7));
  inv1  gate295(.a(N49), .O(gate26inter8));
  nand2 gate296(.a(gate26inter8), .b(gate26inter7), .O(gate26inter9));
  nand2 gate297(.a(s_13), .b(gate26inter3), .O(gate26inter10));
  nor2  gate298(.a(gate26inter10), .b(gate26inter9), .O(gate26inter11));
  nor2  gate299(.a(gate26inter11), .b(gate26inter6), .O(gate26inter12));
  nand2 gate300(.a(gate26inter12), .b(gate26inter1), .O(N275));
xor2 gate27( .a(N5), .b(N21), .O(N276) );
xor2 gate28( .a(N37), .b(N53), .O(N277) );
xor2 gate29( .a(N9), .b(N25), .O(N278) );
xor2 gate30( .a(N41), .b(N57), .O(N279) );
xor2 gate31( .a(N13), .b(N29), .O(N280) );
xor2 gate32( .a(N45), .b(N61), .O(N281) );

  xor2  gate469(.a(N81), .b(N65), .O(gate33inter0));
  nand2 gate470(.a(gate33inter0), .b(s_38), .O(gate33inter1));
  and2  gate471(.a(N81), .b(N65), .O(gate33inter2));
  inv1  gate472(.a(s_38), .O(gate33inter3));
  inv1  gate473(.a(s_39), .O(gate33inter4));
  nand2 gate474(.a(gate33inter4), .b(gate33inter3), .O(gate33inter5));
  nor2  gate475(.a(gate33inter5), .b(gate33inter2), .O(gate33inter6));
  inv1  gate476(.a(N65), .O(gate33inter7));
  inv1  gate477(.a(N81), .O(gate33inter8));
  nand2 gate478(.a(gate33inter8), .b(gate33inter7), .O(gate33inter9));
  nand2 gate479(.a(s_39), .b(gate33inter3), .O(gate33inter10));
  nor2  gate480(.a(gate33inter10), .b(gate33inter9), .O(gate33inter11));
  nor2  gate481(.a(gate33inter11), .b(gate33inter6), .O(gate33inter12));
  nand2 gate482(.a(gate33inter12), .b(gate33inter1), .O(N282));
xor2 gate34( .a(N97), .b(N113), .O(N283) );
xor2 gate35( .a(N69), .b(N85), .O(N284) );

  xor2  gate259(.a(N117), .b(N101), .O(gate36inter0));
  nand2 gate260(.a(gate36inter0), .b(s_8), .O(gate36inter1));
  and2  gate261(.a(N117), .b(N101), .O(gate36inter2));
  inv1  gate262(.a(s_8), .O(gate36inter3));
  inv1  gate263(.a(s_9), .O(gate36inter4));
  nand2 gate264(.a(gate36inter4), .b(gate36inter3), .O(gate36inter5));
  nor2  gate265(.a(gate36inter5), .b(gate36inter2), .O(gate36inter6));
  inv1  gate266(.a(N101), .O(gate36inter7));
  inv1  gate267(.a(N117), .O(gate36inter8));
  nand2 gate268(.a(gate36inter8), .b(gate36inter7), .O(gate36inter9));
  nand2 gate269(.a(s_9), .b(gate36inter3), .O(gate36inter10));
  nor2  gate270(.a(gate36inter10), .b(gate36inter9), .O(gate36inter11));
  nor2  gate271(.a(gate36inter11), .b(gate36inter6), .O(gate36inter12));
  nand2 gate272(.a(gate36inter12), .b(gate36inter1), .O(N285));
xor2 gate37( .a(N73), .b(N89), .O(N286) );
xor2 gate38( .a(N105), .b(N121), .O(N287) );
xor2 gate39( .a(N77), .b(N93), .O(N288) );
xor2 gate40( .a(N109), .b(N125), .O(N289) );
xor2 gate41( .a(N250), .b(N251), .O(N290) );

  xor2  gate371(.a(N253), .b(N252), .O(gate42inter0));
  nand2 gate372(.a(gate42inter0), .b(s_24), .O(gate42inter1));
  and2  gate373(.a(N253), .b(N252), .O(gate42inter2));
  inv1  gate374(.a(s_24), .O(gate42inter3));
  inv1  gate375(.a(s_25), .O(gate42inter4));
  nand2 gate376(.a(gate42inter4), .b(gate42inter3), .O(gate42inter5));
  nor2  gate377(.a(gate42inter5), .b(gate42inter2), .O(gate42inter6));
  inv1  gate378(.a(N252), .O(gate42inter7));
  inv1  gate379(.a(N253), .O(gate42inter8));
  nand2 gate380(.a(gate42inter8), .b(gate42inter7), .O(gate42inter9));
  nand2 gate381(.a(s_25), .b(gate42inter3), .O(gate42inter10));
  nor2  gate382(.a(gate42inter10), .b(gate42inter9), .O(gate42inter11));
  nor2  gate383(.a(gate42inter11), .b(gate42inter6), .O(gate42inter12));
  nand2 gate384(.a(gate42inter12), .b(gate42inter1), .O(N293));
xor2 gate43( .a(N254), .b(N255), .O(N296) );
xor2 gate44( .a(N256), .b(N257), .O(N299) );
xor2 gate45( .a(N258), .b(N259), .O(N302) );
xor2 gate46( .a(N260), .b(N261), .O(N305) );
xor2 gate47( .a(N262), .b(N263), .O(N308) );
xor2 gate48( .a(N264), .b(N265), .O(N311) );
xor2 gate49( .a(N274), .b(N275), .O(N314) );
xor2 gate50( .a(N276), .b(N277), .O(N315) );
xor2 gate51( .a(N278), .b(N279), .O(N316) );
xor2 gate52( .a(N280), .b(N281), .O(N317) );
xor2 gate53( .a(N282), .b(N283), .O(N318) );

  xor2  gate441(.a(N285), .b(N284), .O(gate54inter0));
  nand2 gate442(.a(gate54inter0), .b(s_34), .O(gate54inter1));
  and2  gate443(.a(N285), .b(N284), .O(gate54inter2));
  inv1  gate444(.a(s_34), .O(gate54inter3));
  inv1  gate445(.a(s_35), .O(gate54inter4));
  nand2 gate446(.a(gate54inter4), .b(gate54inter3), .O(gate54inter5));
  nor2  gate447(.a(gate54inter5), .b(gate54inter2), .O(gate54inter6));
  inv1  gate448(.a(N284), .O(gate54inter7));
  inv1  gate449(.a(N285), .O(gate54inter8));
  nand2 gate450(.a(gate54inter8), .b(gate54inter7), .O(gate54inter9));
  nand2 gate451(.a(s_35), .b(gate54inter3), .O(gate54inter10));
  nor2  gate452(.a(gate54inter10), .b(gate54inter9), .O(gate54inter11));
  nor2  gate453(.a(gate54inter11), .b(gate54inter6), .O(gate54inter12));
  nand2 gate454(.a(gate54inter12), .b(gate54inter1), .O(N319));
xor2 gate55( .a(N286), .b(N287), .O(N320) );
xor2 gate56( .a(N288), .b(N289), .O(N321) );
xor2 gate57( .a(N290), .b(N293), .O(N338) );

  xor2  gate427(.a(N299), .b(N296), .O(gate58inter0));
  nand2 gate428(.a(gate58inter0), .b(s_32), .O(gate58inter1));
  and2  gate429(.a(N299), .b(N296), .O(gate58inter2));
  inv1  gate430(.a(s_32), .O(gate58inter3));
  inv1  gate431(.a(s_33), .O(gate58inter4));
  nand2 gate432(.a(gate58inter4), .b(gate58inter3), .O(gate58inter5));
  nor2  gate433(.a(gate58inter5), .b(gate58inter2), .O(gate58inter6));
  inv1  gate434(.a(N296), .O(gate58inter7));
  inv1  gate435(.a(N299), .O(gate58inter8));
  nand2 gate436(.a(gate58inter8), .b(gate58inter7), .O(gate58inter9));
  nand2 gate437(.a(s_33), .b(gate58inter3), .O(gate58inter10));
  nor2  gate438(.a(gate58inter10), .b(gate58inter9), .O(gate58inter11));
  nor2  gate439(.a(gate58inter11), .b(gate58inter6), .O(gate58inter12));
  nand2 gate440(.a(gate58inter12), .b(gate58inter1), .O(N339));
xor2 gate59( .a(N290), .b(N296), .O(N340) );
xor2 gate60( .a(N293), .b(N299), .O(N341) );

  xor2  gate455(.a(N305), .b(N302), .O(gate61inter0));
  nand2 gate456(.a(gate61inter0), .b(s_36), .O(gate61inter1));
  and2  gate457(.a(N305), .b(N302), .O(gate61inter2));
  inv1  gate458(.a(s_36), .O(gate61inter3));
  inv1  gate459(.a(s_37), .O(gate61inter4));
  nand2 gate460(.a(gate61inter4), .b(gate61inter3), .O(gate61inter5));
  nor2  gate461(.a(gate61inter5), .b(gate61inter2), .O(gate61inter6));
  inv1  gate462(.a(N302), .O(gate61inter7));
  inv1  gate463(.a(N305), .O(gate61inter8));
  nand2 gate464(.a(gate61inter8), .b(gate61inter7), .O(gate61inter9));
  nand2 gate465(.a(s_37), .b(gate61inter3), .O(gate61inter10));
  nor2  gate466(.a(gate61inter10), .b(gate61inter9), .O(gate61inter11));
  nor2  gate467(.a(gate61inter11), .b(gate61inter6), .O(gate61inter12));
  nand2 gate468(.a(gate61inter12), .b(gate61inter1), .O(N342));
xor2 gate62( .a(N308), .b(N311), .O(N343) );
xor2 gate63( .a(N302), .b(N308), .O(N344) );

  xor2  gate245(.a(N311), .b(N305), .O(gate64inter0));
  nand2 gate246(.a(gate64inter0), .b(s_6), .O(gate64inter1));
  and2  gate247(.a(N311), .b(N305), .O(gate64inter2));
  inv1  gate248(.a(s_6), .O(gate64inter3));
  inv1  gate249(.a(s_7), .O(gate64inter4));
  nand2 gate250(.a(gate64inter4), .b(gate64inter3), .O(gate64inter5));
  nor2  gate251(.a(gate64inter5), .b(gate64inter2), .O(gate64inter6));
  inv1  gate252(.a(N305), .O(gate64inter7));
  inv1  gate253(.a(N311), .O(gate64inter8));
  nand2 gate254(.a(gate64inter8), .b(gate64inter7), .O(gate64inter9));
  nand2 gate255(.a(s_7), .b(gate64inter3), .O(gate64inter10));
  nor2  gate256(.a(gate64inter10), .b(gate64inter9), .O(gate64inter11));
  nor2  gate257(.a(gate64inter11), .b(gate64inter6), .O(gate64inter12));
  nand2 gate258(.a(gate64inter12), .b(gate64inter1), .O(N345));
xor2 gate65( .a(N266), .b(N342), .O(N346) );
xor2 gate66( .a(N267), .b(N343), .O(N347) );
xor2 gate67( .a(N268), .b(N344), .O(N348) );
xor2 gate68( .a(N269), .b(N345), .O(N349) );

  xor2  gate399(.a(N338), .b(N270), .O(gate69inter0));
  nand2 gate400(.a(gate69inter0), .b(s_28), .O(gate69inter1));
  and2  gate401(.a(N338), .b(N270), .O(gate69inter2));
  inv1  gate402(.a(s_28), .O(gate69inter3));
  inv1  gate403(.a(s_29), .O(gate69inter4));
  nand2 gate404(.a(gate69inter4), .b(gate69inter3), .O(gate69inter5));
  nor2  gate405(.a(gate69inter5), .b(gate69inter2), .O(gate69inter6));
  inv1  gate406(.a(N270), .O(gate69inter7));
  inv1  gate407(.a(N338), .O(gate69inter8));
  nand2 gate408(.a(gate69inter8), .b(gate69inter7), .O(gate69inter9));
  nand2 gate409(.a(s_29), .b(gate69inter3), .O(gate69inter10));
  nor2  gate410(.a(gate69inter10), .b(gate69inter9), .O(gate69inter11));
  nor2  gate411(.a(gate69inter11), .b(gate69inter6), .O(gate69inter12));
  nand2 gate412(.a(gate69inter12), .b(gate69inter1), .O(N350));

  xor2  gate343(.a(N339), .b(N271), .O(gate70inter0));
  nand2 gate344(.a(gate70inter0), .b(s_20), .O(gate70inter1));
  and2  gate345(.a(N339), .b(N271), .O(gate70inter2));
  inv1  gate346(.a(s_20), .O(gate70inter3));
  inv1  gate347(.a(s_21), .O(gate70inter4));
  nand2 gate348(.a(gate70inter4), .b(gate70inter3), .O(gate70inter5));
  nor2  gate349(.a(gate70inter5), .b(gate70inter2), .O(gate70inter6));
  inv1  gate350(.a(N271), .O(gate70inter7));
  inv1  gate351(.a(N339), .O(gate70inter8));
  nand2 gate352(.a(gate70inter8), .b(gate70inter7), .O(gate70inter9));
  nand2 gate353(.a(s_21), .b(gate70inter3), .O(gate70inter10));
  nor2  gate354(.a(gate70inter10), .b(gate70inter9), .O(gate70inter11));
  nor2  gate355(.a(gate70inter11), .b(gate70inter6), .O(gate70inter12));
  nand2 gate356(.a(gate70inter12), .b(gate70inter1), .O(N351));

  xor2  gate413(.a(N340), .b(N272), .O(gate71inter0));
  nand2 gate414(.a(gate71inter0), .b(s_30), .O(gate71inter1));
  and2  gate415(.a(N340), .b(N272), .O(gate71inter2));
  inv1  gate416(.a(s_30), .O(gate71inter3));
  inv1  gate417(.a(s_31), .O(gate71inter4));
  nand2 gate418(.a(gate71inter4), .b(gate71inter3), .O(gate71inter5));
  nor2  gate419(.a(gate71inter5), .b(gate71inter2), .O(gate71inter6));
  inv1  gate420(.a(N272), .O(gate71inter7));
  inv1  gate421(.a(N340), .O(gate71inter8));
  nand2 gate422(.a(gate71inter8), .b(gate71inter7), .O(gate71inter9));
  nand2 gate423(.a(s_31), .b(gate71inter3), .O(gate71inter10));
  nor2  gate424(.a(gate71inter10), .b(gate71inter9), .O(gate71inter11));
  nor2  gate425(.a(gate71inter11), .b(gate71inter6), .O(gate71inter12));
  nand2 gate426(.a(gate71inter12), .b(gate71inter1), .O(N352));
xor2 gate72( .a(N273), .b(N341), .O(N353) );
xor2 gate73( .a(N314), .b(N346), .O(N354) );
xor2 gate74( .a(N315), .b(N347), .O(N367) );
xor2 gate75( .a(N316), .b(N348), .O(N380) );
xor2 gate76( .a(N317), .b(N349), .O(N393) );
xor2 gate77( .a(N318), .b(N350), .O(N406) );
xor2 gate78( .a(N319), .b(N351), .O(N419) );
xor2 gate79( .a(N320), .b(N352), .O(N432) );

  xor2  gate483(.a(N353), .b(N321), .O(gate80inter0));
  nand2 gate484(.a(gate80inter0), .b(s_40), .O(gate80inter1));
  and2  gate485(.a(N353), .b(N321), .O(gate80inter2));
  inv1  gate486(.a(s_40), .O(gate80inter3));
  inv1  gate487(.a(s_41), .O(gate80inter4));
  nand2 gate488(.a(gate80inter4), .b(gate80inter3), .O(gate80inter5));
  nor2  gate489(.a(gate80inter5), .b(gate80inter2), .O(gate80inter6));
  inv1  gate490(.a(N321), .O(gate80inter7));
  inv1  gate491(.a(N353), .O(gate80inter8));
  nand2 gate492(.a(gate80inter8), .b(gate80inter7), .O(gate80inter9));
  nand2 gate493(.a(s_41), .b(gate80inter3), .O(gate80inter10));
  nor2  gate494(.a(gate80inter10), .b(gate80inter9), .O(gate80inter11));
  nor2  gate495(.a(gate80inter11), .b(gate80inter6), .O(gate80inter12));
  nand2 gate496(.a(gate80inter12), .b(gate80inter1), .O(N445));
inv1 gate81( .a(N354), .O(N554) );
inv1 gate82( .a(N367), .O(N555) );
inv1 gate83( .a(N380), .O(N556) );
inv1 gate84( .a(N354), .O(N557) );
inv1 gate85( .a(N367), .O(N558) );
inv1 gate86( .a(N393), .O(N559) );
inv1 gate87( .a(N354), .O(N560) );
inv1 gate88( .a(N380), .O(N561) );
inv1 gate89( .a(N393), .O(N562) );
inv1 gate90( .a(N367), .O(N563) );
inv1 gate91( .a(N380), .O(N564) );
inv1 gate92( .a(N393), .O(N565) );
inv1 gate93( .a(N419), .O(N566) );
inv1 gate94( .a(N445), .O(N567) );
inv1 gate95( .a(N419), .O(N568) );
inv1 gate96( .a(N432), .O(N569) );
inv1 gate97( .a(N406), .O(N570) );
inv1 gate98( .a(N445), .O(N571) );
inv1 gate99( .a(N406), .O(N572) );
inv1 gate100( .a(N432), .O(N573) );
inv1 gate101( .a(N406), .O(N574) );
inv1 gate102( .a(N419), .O(N575) );
inv1 gate103( .a(N432), .O(N576) );
inv1 gate104( .a(N406), .O(N577) );
inv1 gate105( .a(N419), .O(N578) );
inv1 gate106( .a(N445), .O(N579) );
inv1 gate107( .a(N406), .O(N580) );
inv1 gate108( .a(N432), .O(N581) );
inv1 gate109( .a(N445), .O(N582) );
inv1 gate110( .a(N419), .O(N583) );
inv1 gate111( .a(N432), .O(N584) );
inv1 gate112( .a(N445), .O(N585) );
inv1 gate113( .a(N367), .O(N586) );
inv1 gate114( .a(N393), .O(N587) );
inv1 gate115( .a(N367), .O(N588) );
inv1 gate116( .a(N380), .O(N589) );
inv1 gate117( .a(N354), .O(N590) );
inv1 gate118( .a(N393), .O(N591) );
inv1 gate119( .a(N354), .O(N592) );
inv1 gate120( .a(N380), .O(N593) );
and4 gate121( .a(N554), .b(N555), .c(N556), .d(N393), .O(N594) );
and4 gate122( .a(N557), .b(N558), .c(N380), .d(N559), .O(N595) );
and4 gate123( .a(N560), .b(N367), .c(N561), .d(N562), .O(N596) );
and4 gate124( .a(N354), .b(N563), .c(N564), .d(N565), .O(N597) );
and4 gate125( .a(N574), .b(N575), .c(N576), .d(N445), .O(N598) );
and4 gate126( .a(N577), .b(N578), .c(N432), .d(N579), .O(N599) );
and4 gate127( .a(N580), .b(N419), .c(N581), .d(N582), .O(N600) );
and4 gate128( .a(N406), .b(N583), .c(N584), .d(N585), .O(N601) );
or4 gate129( .a(N594), .b(N595), .c(N596), .d(N597), .O(N602) );
or4 gate130( .a(N598), .b(N599), .c(N600), .d(N601), .O(N607) );
and5 gate131( .a(N406), .b(N566), .c(N432), .d(N567), .e(N602), .O(N620) );
and5 gate132( .a(N406), .b(N568), .c(N569), .d(N445), .e(N602), .O(N625) );
and5 gate133( .a(N570), .b(N419), .c(N432), .d(N571), .e(N602), .O(N630) );
and5 gate134( .a(N572), .b(N419), .c(N573), .d(N445), .e(N602), .O(N635) );
and5 gate135( .a(N354), .b(N586), .c(N380), .d(N587), .e(N607), .O(N640) );
and5 gate136( .a(N354), .b(N588), .c(N589), .d(N393), .e(N607), .O(N645) );
and5 gate137( .a(N590), .b(N367), .c(N380), .d(N591), .e(N607), .O(N650) );
and5 gate138( .a(N592), .b(N367), .c(N593), .d(N393), .e(N607), .O(N655) );
and2 gate139( .a(N354), .b(N620), .O(N692) );
and2 gate140( .a(N367), .b(N620), .O(N693) );
and2 gate141( .a(N380), .b(N620), .O(N694) );
and2 gate142( .a(N393), .b(N620), .O(N695) );
and2 gate143( .a(N354), .b(N625), .O(N696) );
and2 gate144( .a(N367), .b(N625), .O(N697) );
and2 gate145( .a(N380), .b(N625), .O(N698) );
and2 gate146( .a(N393), .b(N625), .O(N699) );
and2 gate147( .a(N354), .b(N630), .O(N700) );
and2 gate148( .a(N367), .b(N630), .O(N701) );
and2 gate149( .a(N380), .b(N630), .O(N702) );
and2 gate150( .a(N393), .b(N630), .O(N703) );
and2 gate151( .a(N354), .b(N635), .O(N704) );
and2 gate152( .a(N367), .b(N635), .O(N705) );
and2 gate153( .a(N380), .b(N635), .O(N706) );
and2 gate154( .a(N393), .b(N635), .O(N707) );
and2 gate155( .a(N406), .b(N640), .O(N708) );
and2 gate156( .a(N419), .b(N640), .O(N709) );
and2 gate157( .a(N432), .b(N640), .O(N710) );
and2 gate158( .a(N445), .b(N640), .O(N711) );
and2 gate159( .a(N406), .b(N645), .O(N712) );
and2 gate160( .a(N419), .b(N645), .O(N713) );
and2 gate161( .a(N432), .b(N645), .O(N714) );
and2 gate162( .a(N445), .b(N645), .O(N715) );
and2 gate163( .a(N406), .b(N650), .O(N716) );
and2 gate164( .a(N419), .b(N650), .O(N717) );
and2 gate165( .a(N432), .b(N650), .O(N718) );
and2 gate166( .a(N445), .b(N650), .O(N719) );
and2 gate167( .a(N406), .b(N655), .O(N720) );
and2 gate168( .a(N419), .b(N655), .O(N721) );
and2 gate169( .a(N432), .b(N655), .O(N722) );
and2 gate170( .a(N445), .b(N655), .O(N723) );
xor2 gate171( .a(N1), .b(N692), .O(N724) );

  xor2  gate273(.a(N693), .b(N5), .O(gate172inter0));
  nand2 gate274(.a(gate172inter0), .b(s_10), .O(gate172inter1));
  and2  gate275(.a(N693), .b(N5), .O(gate172inter2));
  inv1  gate276(.a(s_10), .O(gate172inter3));
  inv1  gate277(.a(s_11), .O(gate172inter4));
  nand2 gate278(.a(gate172inter4), .b(gate172inter3), .O(gate172inter5));
  nor2  gate279(.a(gate172inter5), .b(gate172inter2), .O(gate172inter6));
  inv1  gate280(.a(N5), .O(gate172inter7));
  inv1  gate281(.a(N693), .O(gate172inter8));
  nand2 gate282(.a(gate172inter8), .b(gate172inter7), .O(gate172inter9));
  nand2 gate283(.a(s_11), .b(gate172inter3), .O(gate172inter10));
  nor2  gate284(.a(gate172inter10), .b(gate172inter9), .O(gate172inter11));
  nor2  gate285(.a(gate172inter11), .b(gate172inter6), .O(gate172inter12));
  nand2 gate286(.a(gate172inter12), .b(gate172inter1), .O(N725));
xor2 gate173( .a(N9), .b(N694), .O(N726) );
xor2 gate174( .a(N13), .b(N695), .O(N727) );
xor2 gate175( .a(N17), .b(N696), .O(N728) );
xor2 gate176( .a(N21), .b(N697), .O(N729) );
xor2 gate177( .a(N25), .b(N698), .O(N730) );
xor2 gate178( .a(N29), .b(N699), .O(N731) );
xor2 gate179( .a(N33), .b(N700), .O(N732) );
xor2 gate180( .a(N37), .b(N701), .O(N733) );
xor2 gate181( .a(N41), .b(N702), .O(N734) );
xor2 gate182( .a(N45), .b(N703), .O(N735) );
xor2 gate183( .a(N49), .b(N704), .O(N736) );
xor2 gate184( .a(N53), .b(N705), .O(N737) );
xor2 gate185( .a(N57), .b(N706), .O(N738) );
xor2 gate186( .a(N61), .b(N707), .O(N739) );

  xor2  gate217(.a(N708), .b(N65), .O(gate187inter0));
  nand2 gate218(.a(gate187inter0), .b(s_2), .O(gate187inter1));
  and2  gate219(.a(N708), .b(N65), .O(gate187inter2));
  inv1  gate220(.a(s_2), .O(gate187inter3));
  inv1  gate221(.a(s_3), .O(gate187inter4));
  nand2 gate222(.a(gate187inter4), .b(gate187inter3), .O(gate187inter5));
  nor2  gate223(.a(gate187inter5), .b(gate187inter2), .O(gate187inter6));
  inv1  gate224(.a(N65), .O(gate187inter7));
  inv1  gate225(.a(N708), .O(gate187inter8));
  nand2 gate226(.a(gate187inter8), .b(gate187inter7), .O(gate187inter9));
  nand2 gate227(.a(s_3), .b(gate187inter3), .O(gate187inter10));
  nor2  gate228(.a(gate187inter10), .b(gate187inter9), .O(gate187inter11));
  nor2  gate229(.a(gate187inter11), .b(gate187inter6), .O(gate187inter12));
  nand2 gate230(.a(gate187inter12), .b(gate187inter1), .O(N740));

  xor2  gate203(.a(N709), .b(N69), .O(gate188inter0));
  nand2 gate204(.a(gate188inter0), .b(s_0), .O(gate188inter1));
  and2  gate205(.a(N709), .b(N69), .O(gate188inter2));
  inv1  gate206(.a(s_0), .O(gate188inter3));
  inv1  gate207(.a(s_1), .O(gate188inter4));
  nand2 gate208(.a(gate188inter4), .b(gate188inter3), .O(gate188inter5));
  nor2  gate209(.a(gate188inter5), .b(gate188inter2), .O(gate188inter6));
  inv1  gate210(.a(N69), .O(gate188inter7));
  inv1  gate211(.a(N709), .O(gate188inter8));
  nand2 gate212(.a(gate188inter8), .b(gate188inter7), .O(gate188inter9));
  nand2 gate213(.a(s_1), .b(gate188inter3), .O(gate188inter10));
  nor2  gate214(.a(gate188inter10), .b(gate188inter9), .O(gate188inter11));
  nor2  gate215(.a(gate188inter11), .b(gate188inter6), .O(gate188inter12));
  nand2 gate216(.a(gate188inter12), .b(gate188inter1), .O(N741));
xor2 gate189( .a(N73), .b(N710), .O(N742) );

  xor2  gate329(.a(N711), .b(N77), .O(gate190inter0));
  nand2 gate330(.a(gate190inter0), .b(s_18), .O(gate190inter1));
  and2  gate331(.a(N711), .b(N77), .O(gate190inter2));
  inv1  gate332(.a(s_18), .O(gate190inter3));
  inv1  gate333(.a(s_19), .O(gate190inter4));
  nand2 gate334(.a(gate190inter4), .b(gate190inter3), .O(gate190inter5));
  nor2  gate335(.a(gate190inter5), .b(gate190inter2), .O(gate190inter6));
  inv1  gate336(.a(N77), .O(gate190inter7));
  inv1  gate337(.a(N711), .O(gate190inter8));
  nand2 gate338(.a(gate190inter8), .b(gate190inter7), .O(gate190inter9));
  nand2 gate339(.a(s_19), .b(gate190inter3), .O(gate190inter10));
  nor2  gate340(.a(gate190inter10), .b(gate190inter9), .O(gate190inter11));
  nor2  gate341(.a(gate190inter11), .b(gate190inter6), .O(gate190inter12));
  nand2 gate342(.a(gate190inter12), .b(gate190inter1), .O(N743));
xor2 gate191( .a(N81), .b(N712), .O(N744) );
xor2 gate192( .a(N85), .b(N713), .O(N745) );
xor2 gate193( .a(N89), .b(N714), .O(N746) );
xor2 gate194( .a(N93), .b(N715), .O(N747) );
xor2 gate195( .a(N97), .b(N716), .O(N748) );

  xor2  gate231(.a(N717), .b(N101), .O(gate196inter0));
  nand2 gate232(.a(gate196inter0), .b(s_4), .O(gate196inter1));
  and2  gate233(.a(N717), .b(N101), .O(gate196inter2));
  inv1  gate234(.a(s_4), .O(gate196inter3));
  inv1  gate235(.a(s_5), .O(gate196inter4));
  nand2 gate236(.a(gate196inter4), .b(gate196inter3), .O(gate196inter5));
  nor2  gate237(.a(gate196inter5), .b(gate196inter2), .O(gate196inter6));
  inv1  gate238(.a(N101), .O(gate196inter7));
  inv1  gate239(.a(N717), .O(gate196inter8));
  nand2 gate240(.a(gate196inter8), .b(gate196inter7), .O(gate196inter9));
  nand2 gate241(.a(s_5), .b(gate196inter3), .O(gate196inter10));
  nor2  gate242(.a(gate196inter10), .b(gate196inter9), .O(gate196inter11));
  nor2  gate243(.a(gate196inter11), .b(gate196inter6), .O(gate196inter12));
  nand2 gate244(.a(gate196inter12), .b(gate196inter1), .O(N749));
xor2 gate197( .a(N105), .b(N718), .O(N750) );

  xor2  gate385(.a(N719), .b(N109), .O(gate198inter0));
  nand2 gate386(.a(gate198inter0), .b(s_26), .O(gate198inter1));
  and2  gate387(.a(N719), .b(N109), .O(gate198inter2));
  inv1  gate388(.a(s_26), .O(gate198inter3));
  inv1  gate389(.a(s_27), .O(gate198inter4));
  nand2 gate390(.a(gate198inter4), .b(gate198inter3), .O(gate198inter5));
  nor2  gate391(.a(gate198inter5), .b(gate198inter2), .O(gate198inter6));
  inv1  gate392(.a(N109), .O(gate198inter7));
  inv1  gate393(.a(N719), .O(gate198inter8));
  nand2 gate394(.a(gate198inter8), .b(gate198inter7), .O(gate198inter9));
  nand2 gate395(.a(s_27), .b(gate198inter3), .O(gate198inter10));
  nor2  gate396(.a(gate198inter10), .b(gate198inter9), .O(gate198inter11));
  nor2  gate397(.a(gate198inter11), .b(gate198inter6), .O(gate198inter12));
  nand2 gate398(.a(gate198inter12), .b(gate198inter1), .O(N751));
xor2 gate199( .a(N113), .b(N720), .O(N752) );
xor2 gate200( .a(N117), .b(N721), .O(N753) );

  xor2  gate315(.a(N722), .b(N121), .O(gate201inter0));
  nand2 gate316(.a(gate201inter0), .b(s_16), .O(gate201inter1));
  and2  gate317(.a(N722), .b(N121), .O(gate201inter2));
  inv1  gate318(.a(s_16), .O(gate201inter3));
  inv1  gate319(.a(s_17), .O(gate201inter4));
  nand2 gate320(.a(gate201inter4), .b(gate201inter3), .O(gate201inter5));
  nor2  gate321(.a(gate201inter5), .b(gate201inter2), .O(gate201inter6));
  inv1  gate322(.a(N121), .O(gate201inter7));
  inv1  gate323(.a(N722), .O(gate201inter8));
  nand2 gate324(.a(gate201inter8), .b(gate201inter7), .O(gate201inter9));
  nand2 gate325(.a(s_17), .b(gate201inter3), .O(gate201inter10));
  nor2  gate326(.a(gate201inter10), .b(gate201inter9), .O(gate201inter11));
  nor2  gate327(.a(gate201inter11), .b(gate201inter6), .O(gate201inter12));
  nand2 gate328(.a(gate201inter12), .b(gate201inter1), .O(N754));
xor2 gate202( .a(N125), .b(N723), .O(N755) );

endmodule