module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);

input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;//RE__PI;

input s_0,s_1;//RE__ALLOW(00,01,10,11);
input s_2,s_3;//RE__ALLOW(00,01,10,11);
input s_4,s_5;//RE__ALLOW(00,01,10,11);
input s_6,s_7;//RE__ALLOW(00,01,10,11);
input s_8,s_9;//RE__ALLOW(00,01,10,11);
input s_10,s_11;//RE__ALLOW(00,01,10,11);
input s_12,s_13;//RE__ALLOW(00,01,10,11);
input s_14,s_15;//RE__ALLOW(00,01,10,11);
input s_16,s_17;//RE__ALLOW(00,01,10,11);
input s_18,s_19;//RE__ALLOW(00,01,10,11);
input s_20,s_21;//RE__ALLOW(00,01,10,11);
input s_22,s_23;//RE__ALLOW(00,01,10,11);
input s_24,s_25;//RE__ALLOW(00,01,10,11);
input s_26,s_27;//RE__ALLOW(00,01,10,11);
input s_28,s_29;//RE__ALLOW(00,01,10,11);
input s_30,s_31;//RE__ALLOW(00,01,10,11);
input s_32,s_33;//RE__ALLOW(00,01,10,11);
input s_34,s_35;//RE__ALLOW(00,01,10,11);
input s_36,s_37;//RE__ALLOW(00,01,10,11);
input s_38,s_39;//RE__ALLOW(00,01,10,11);
input s_40,s_41;//RE__ALLOW(00,01,10,11);
input s_42,s_43;//RE__ALLOW(00,01,10,11);
input s_44,s_45;//RE__ALLOW(00,01,10,11);
input s_46,s_47;//RE__ALLOW(00,01,10,11);
input s_48,s_49;//RE__ALLOW(00,01,10,11);
input s_50,s_51;//RE__ALLOW(00,01,10,11);
input s_52,s_53;//RE__ALLOW(00,01,10,11);
input s_54,s_55;//RE__ALLOW(00,01,10,11);
input s_56,s_57;//RE__ALLOW(00,01,10,11);
input s_58,s_59;//RE__ALLOW(00,01,10,11);
input s_60,s_61;//RE__ALLOW(00,01,10,11);
input s_62,s_63;//RE__ALLOW(00,01,10,11);
input s_64,s_65;//RE__ALLOW(00,01,10,11);
input s_66,s_67;//RE__ALLOW(00,01,10,11);
input s_68,s_69;//RE__ALLOW(00,01,10,11);
input s_70,s_71;//RE__ALLOW(00,01,10,11);
input s_72,s_73;//RE__ALLOW(00,01,10,11);
input s_74,s_75;//RE__ALLOW(00,01,10,11);
input s_76,s_77;//RE__ALLOW(00,01,10,11);
input s_78,s_79;//RE__ALLOW(00,01,10,11);
input s_80,s_81;//RE__ALLOW(00,01,10,11);
input s_82,s_83;//RE__ALLOW(00,01,10,11);
input s_84,s_85;//RE__ALLOW(00,01,10,11);
input s_86,s_87;//RE__ALLOW(00,01,10,11);
input s_88,s_89;//RE__ALLOW(00,01,10,11);
input s_90,s_91;//RE__ALLOW(00,01,10,11);
input s_92,s_93;//RE__ALLOW(00,01,10,11);
input s_94,s_95;//RE__ALLOW(00,01,10,11);
input s_96,s_97;//RE__ALLOW(00,01,10,11);
input s_98,s_99;//RE__ALLOW(00,01,10,11);
input s_100,s_101;//RE__ALLOW(00,01,10,11);
input s_102,s_103;//RE__ALLOW(00,01,10,11);
input s_104,s_105;//RE__ALLOW(00,01,10,11);
input s_106,s_107;//RE__ALLOW(00,01,10,11);
input s_108,s_109;//RE__ALLOW(00,01,10,11);
input s_110,s_111;//RE__ALLOW(00,01,10,11);
input s_112,s_113;//RE__ALLOW(00,01,10,11);
input s_114,s_115;//RE__ALLOW(00,01,10,11);
input s_116,s_117;//RE__ALLOW(00,01,10,11);
input s_118,s_119;//RE__ALLOW(00,01,10,11);
input s_120,s_121;//RE__ALLOW(00,01,10,11);
input s_122,s_123;//RE__ALLOW(00,01,10,11);
input s_124,s_125;//RE__ALLOW(00,01,10,11);
input s_126,s_127;//RE__ALLOW(00,01,10,11);
input s_128,s_129;//RE__ALLOW(00,01,10,11);
input s_130,s_131;//RE__ALLOW(00,01,10,11);
input s_132,s_133;//RE__ALLOW(00,01,10,11);
input s_134,s_135;//RE__ALLOW(00,01,10,11);
input s_136,s_137;//RE__ALLOW(00,01,10,11);
input s_138,s_139;//RE__ALLOW(00,01,10,11);
input s_140,s_141;//RE__ALLOW(00,01,10,11);
input s_142,s_143;//RE__ALLOW(00,01,10,11);
input s_144,s_145;//RE__ALLOW(00,01,10,11);
input s_146,s_147;//RE__ALLOW(00,01,10,11);
input s_148,s_149;//RE__ALLOW(00,01,10,11);
input s_150,s_151;//RE__ALLOW(00,01,10,11);
input s_152,s_153;//RE__ALLOW(00,01,10,11);
input s_154,s_155;//RE__ALLOW(00,01,10,11);
input s_156,s_157;//RE__ALLOW(00,01,10,11);
input s_158,s_159;//RE__ALLOW(00,01,10,11);
input s_160,s_161;//RE__ALLOW(00,01,10,11);
input s_162,s_163;//RE__ALLOW(00,01,10,11);
input s_164,s_165;//RE__ALLOW(00,01,10,11);
input s_166,s_167;//RE__ALLOW(00,01,10,11);
input s_168,s_169;//RE__ALLOW(00,01,10,11);
input s_170,s_171;//RE__ALLOW(00,01,10,11);
input s_172,s_173;//RE__ALLOW(00,01,10,11);
input s_174,s_175;//RE__ALLOW(00,01,10,11);
input s_176,s_177;//RE__ALLOW(00,01,10,11);
input s_178,s_179;//RE__ALLOW(00,01,10,11);
input s_180,s_181;//RE__ALLOW(00,01,10,11);
input s_182,s_183;//RE__ALLOW(00,01,10,11);
input s_184,s_185;//RE__ALLOW(00,01,10,11);
input s_186,s_187;//RE__ALLOW(00,01,10,11);
input s_188,s_189;//RE__ALLOW(00,01,10,11);
input s_190,s_191;//RE__ALLOW(00,01,10,11);
input s_192,s_193;//RE__ALLOW(00,01,10,11);
input s_194,s_195;//RE__ALLOW(00,01,10,11);
input s_196,s_197;//RE__ALLOW(00,01,10,11);
input s_198,s_199;//RE__ALLOW(00,01,10,11);
input s_200,s_201;//RE__ALLOW(00,01,10,11);
input s_202,s_203;//RE__ALLOW(00,01,10,11);
input s_204,s_205;//RE__ALLOW(00,01,10,11);
input s_206,s_207;//RE__ALLOW(00,01,10,11);
input s_208,s_209;//RE__ALLOW(00,01,10,11);
input s_210,s_211;//RE__ALLOW(00,01,10,11);
input s_212,s_213;//RE__ALLOW(00,01,10,11);
input s_214,s_215;//RE__ALLOW(00,01,10,11);
input s_216,s_217;//RE__ALLOW(00,01,10,11);
input s_218,s_219;//RE__ALLOW(00,01,10,11);
input s_220,s_221;//RE__ALLOW(00,01,10,11);
input s_222,s_223;//RE__ALLOW(00,01,10,11);
input s_224,s_225;//RE__ALLOW(00,01,10,11);
input s_226,s_227;//RE__ALLOW(00,01,10,11);
input s_228,s_229;//RE__ALLOW(00,01,10,11);
input s_230,s_231;//RE__ALLOW(00,01,10,11);
input s_232,s_233;//RE__ALLOW(00,01,10,11);
input s_234,s_235;//RE__ALLOW(00,01,10,11);
input s_236,s_237;//RE__ALLOW(00,01,10,11);
input s_238,s_239;//RE__ALLOW(00,01,10,11);
input s_240,s_241;//RE__ALLOW(00,01,10,11);
input s_242,s_243;//RE__ALLOW(00,01,10,11);
input s_244,s_245;//RE__ALLOW(00,01,10,11);
input s_246,s_247;//RE__ALLOW(00,01,10,11);
input s_248,s_249;//RE__ALLOW(00,01,10,11);
input s_250,s_251;//RE__ALLOW(00,01,10,11);
input s_252,s_253;//RE__ALLOW(00,01,10,11);
input s_254,s_255;//RE__ALLOW(00,01,10,11);
input s_256,s_257;//RE__ALLOW(00,01,10,11);
input s_258,s_259;//RE__ALLOW(00,01,10,11);
input s_260,s_261;//RE__ALLOW(00,01,10,11);
input s_262,s_263;//RE__ALLOW(00,01,10,11);
input s_264,s_265;//RE__ALLOW(00,01,10,11);
input s_266,s_267;//RE__ALLOW(00,01,10,11);
input s_268,s_269;//RE__ALLOW(00,01,10,11);
input s_270,s_271;//RE__ALLOW(00,01,10,11);
input s_272,s_273;//RE__ALLOW(00,01,10,11);
input s_274,s_275;//RE__ALLOW(00,01,10,11);
input s_276,s_277;//RE__ALLOW(00,01,10,11);
input s_278,s_279;//RE__ALLOW(00,01,10,11);
input s_280,s_281;//RE__ALLOW(00,01,10,11);
input s_282,s_283;//RE__ALLOW(00,01,10,11);
input s_284,s_285;//RE__ALLOW(00,01,10,11);
input s_286,s_287;//RE__ALLOW(00,01,10,11);
input s_288,s_289;//RE__ALLOW(00,01,10,11);
input s_290,s_291;//RE__ALLOW(00,01,10,11);
input s_292,s_293;//RE__ALLOW(00,01,10,11);
input s_294,s_295;//RE__ALLOW(00,01,10,11);
input s_296,s_297;//RE__ALLOW(00,01,10,11);
input s_298,s_299;//RE__ALLOW(00,01,10,11);
input s_300,s_301;//RE__ALLOW(00,01,10,11);
input s_302,s_303;//RE__ALLOW(00,01,10,11);
input s_304,s_305;//RE__ALLOW(00,01,10,11);
input s_306,s_307;//RE__ALLOW(00,01,10,11);
input s_308,s_309;//RE__ALLOW(00,01,10,11);
input s_310,s_311;//RE__ALLOW(00,01,10,11);
input s_312,s_313;//RE__ALLOW(00,01,10,11);
input s_314,s_315;//RE__ALLOW(00,01,10,11);
input s_316,s_317;//RE__ALLOW(00,01,10,11);
input s_318,s_319;//RE__ALLOW(00,01,10,11);
input s_320,s_321;//RE__ALLOW(00,01,10,11);
input s_322,s_323;//RE__ALLOW(00,01,10,11);
input s_324,s_325;//RE__ALLOW(00,01,10,11);
input s_326,s_327;//RE__ALLOW(00,01,10,11);
input s_328,s_329;//RE__ALLOW(00,01,10,11);
input s_330,s_331;//RE__ALLOW(00,01,10,11);
input s_332,s_333;//RE__ALLOW(00,01,10,11);
input s_334,s_335;//RE__ALLOW(00,01,10,11);
input s_336,s_337;//RE__ALLOW(00,01,10,11);
input s_338,s_339;//RE__ALLOW(00,01,10,11);
input s_340,s_341;//RE__ALLOW(00,01,10,11);
input s_342,s_343;//RE__ALLOW(00,01,10,11);
input s_344,s_345;//RE__ALLOW(00,01,10,11);
input s_346,s_347;//RE__ALLOW(00,01,10,11);
input s_348,s_349;//RE__ALLOW(00,01,10,11);
input s_350,s_351;//RE__ALLOW(00,01,10,11);
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;

  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate445inter0, gate445inter1, gate445inter2, gate445inter3, gate445inter4, gate445inter5, gate445inter6, gate445inter7, gate445inter8, gate445inter9, gate445inter10, gate445inter11, gate445inter12, gate510inter0, gate510inter1, gate510inter2, gate510inter3, gate510inter4, gate510inter5, gate510inter6, gate510inter7, gate510inter8, gate510inter9, gate510inter10, gate510inter11, gate510inter12, gate273inter0, gate273inter1, gate273inter2, gate273inter3, gate273inter4, gate273inter5, gate273inter6, gate273inter7, gate273inter8, gate273inter9, gate273inter10, gate273inter11, gate273inter12, gate256inter0, gate256inter1, gate256inter2, gate256inter3, gate256inter4, gate256inter5, gate256inter6, gate256inter7, gate256inter8, gate256inter9, gate256inter10, gate256inter11, gate256inter12, gate155inter0, gate155inter1, gate155inter2, gate155inter3, gate155inter4, gate155inter5, gate155inter6, gate155inter7, gate155inter8, gate155inter9, gate155inter10, gate155inter11, gate155inter12, gate460inter0, gate460inter1, gate460inter2, gate460inter3, gate460inter4, gate460inter5, gate460inter6, gate460inter7, gate460inter8, gate460inter9, gate460inter10, gate460inter11, gate460inter12, gate509inter0, gate509inter1, gate509inter2, gate509inter3, gate509inter4, gate509inter5, gate509inter6, gate509inter7, gate509inter8, gate509inter9, gate509inter10, gate509inter11, gate509inter12, gate433inter0, gate433inter1, gate433inter2, gate433inter3, gate433inter4, gate433inter5, gate433inter6, gate433inter7, gate433inter8, gate433inter9, gate433inter10, gate433inter11, gate433inter12, gate109inter0, gate109inter1, gate109inter2, gate109inter3, gate109inter4, gate109inter5, gate109inter6, gate109inter7, gate109inter8, gate109inter9, gate109inter10, gate109inter11, gate109inter12, gate62inter0, gate62inter1, gate62inter2, gate62inter3, gate62inter4, gate62inter5, gate62inter6, gate62inter7, gate62inter8, gate62inter9, gate62inter10, gate62inter11, gate62inter12, gate247inter0, gate247inter1, gate247inter2, gate247inter3, gate247inter4, gate247inter5, gate247inter6, gate247inter7, gate247inter8, gate247inter9, gate247inter10, gate247inter11, gate247inter12, gate453inter0, gate453inter1, gate453inter2, gate453inter3, gate453inter4, gate453inter5, gate453inter6, gate453inter7, gate453inter8, gate453inter9, gate453inter10, gate453inter11, gate453inter12, gate467inter0, gate467inter1, gate467inter2, gate467inter3, gate467inter4, gate467inter5, gate467inter6, gate467inter7, gate467inter8, gate467inter9, gate467inter10, gate467inter11, gate467inter12, gate281inter0, gate281inter1, gate281inter2, gate281inter3, gate281inter4, gate281inter5, gate281inter6, gate281inter7, gate281inter8, gate281inter9, gate281inter10, gate281inter11, gate281inter12, gate208inter0, gate208inter1, gate208inter2, gate208inter3, gate208inter4, gate208inter5, gate208inter6, gate208inter7, gate208inter8, gate208inter9, gate208inter10, gate208inter11, gate208inter12, gate65inter0, gate65inter1, gate65inter2, gate65inter3, gate65inter4, gate65inter5, gate65inter6, gate65inter7, gate65inter8, gate65inter9, gate65inter10, gate65inter11, gate65inter12, gate263inter0, gate263inter1, gate263inter2, gate263inter3, gate263inter4, gate263inter5, gate263inter6, gate263inter7, gate263inter8, gate263inter9, gate263inter10, gate263inter11, gate263inter12, gate85inter0, gate85inter1, gate85inter2, gate85inter3, gate85inter4, gate85inter5, gate85inter6, gate85inter7, gate85inter8, gate85inter9, gate85inter10, gate85inter11, gate85inter12, gate224inter0, gate224inter1, gate224inter2, gate224inter3, gate224inter4, gate224inter5, gate224inter6, gate224inter7, gate224inter8, gate224inter9, gate224inter10, gate224inter11, gate224inter12, gate161inter0, gate161inter1, gate161inter2, gate161inter3, gate161inter4, gate161inter5, gate161inter6, gate161inter7, gate161inter8, gate161inter9, gate161inter10, gate161inter11, gate161inter12, gate59inter0, gate59inter1, gate59inter2, gate59inter3, gate59inter4, gate59inter5, gate59inter6, gate59inter7, gate59inter8, gate59inter9, gate59inter10, gate59inter11, gate59inter12, gate29inter0, gate29inter1, gate29inter2, gate29inter3, gate29inter4, gate29inter5, gate29inter6, gate29inter7, gate29inter8, gate29inter9, gate29inter10, gate29inter11, gate29inter12, gate153inter0, gate153inter1, gate153inter2, gate153inter3, gate153inter4, gate153inter5, gate153inter6, gate153inter7, gate153inter8, gate153inter9, gate153inter10, gate153inter11, gate153inter12, gate16inter0, gate16inter1, gate16inter2, gate16inter3, gate16inter4, gate16inter5, gate16inter6, gate16inter7, gate16inter8, gate16inter9, gate16inter10, gate16inter11, gate16inter12, gate205inter0, gate205inter1, gate205inter2, gate205inter3, gate205inter4, gate205inter5, gate205inter6, gate205inter7, gate205inter8, gate205inter9, gate205inter10, gate205inter11, gate205inter12, gate254inter0, gate254inter1, gate254inter2, gate254inter3, gate254inter4, gate254inter5, gate254inter6, gate254inter7, gate254inter8, gate254inter9, gate254inter10, gate254inter11, gate254inter12, gate43inter0, gate43inter1, gate43inter2, gate43inter3, gate43inter4, gate43inter5, gate43inter6, gate43inter7, gate43inter8, gate43inter9, gate43inter10, gate43inter11, gate43inter12, gate37inter0, gate37inter1, gate37inter2, gate37inter3, gate37inter4, gate37inter5, gate37inter6, gate37inter7, gate37inter8, gate37inter9, gate37inter10, gate37inter11, gate37inter12, gate240inter0, gate240inter1, gate240inter2, gate240inter3, gate240inter4, gate240inter5, gate240inter6, gate240inter7, gate240inter8, gate240inter9, gate240inter10, gate240inter11, gate240inter12, gate216inter0, gate216inter1, gate216inter2, gate216inter3, gate216inter4, gate216inter5, gate216inter6, gate216inter7, gate216inter8, gate216inter9, gate216inter10, gate216inter11, gate216inter12, gate54inter0, gate54inter1, gate54inter2, gate54inter3, gate54inter4, gate54inter5, gate54inter6, gate54inter7, gate54inter8, gate54inter9, gate54inter10, gate54inter11, gate54inter12, gate506inter0, gate506inter1, gate506inter2, gate506inter3, gate506inter4, gate506inter5, gate506inter6, gate506inter7, gate506inter8, gate506inter9, gate506inter10, gate506inter11, gate506inter12, gate296inter0, gate296inter1, gate296inter2, gate296inter3, gate296inter4, gate296inter5, gate296inter6, gate296inter7, gate296inter8, gate296inter9, gate296inter10, gate296inter11, gate296inter12, gate128inter0, gate128inter1, gate128inter2, gate128inter3, gate128inter4, gate128inter5, gate128inter6, gate128inter7, gate128inter8, gate128inter9, gate128inter10, gate128inter11, gate128inter12, gate38inter0, gate38inter1, gate38inter2, gate38inter3, gate38inter4, gate38inter5, gate38inter6, gate38inter7, gate38inter8, gate38inter9, gate38inter10, gate38inter11, gate38inter12, gate105inter0, gate105inter1, gate105inter2, gate105inter3, gate105inter4, gate105inter5, gate105inter6, gate105inter7, gate105inter8, gate105inter9, gate105inter10, gate105inter11, gate105inter12, gate10inter0, gate10inter1, gate10inter2, gate10inter3, gate10inter4, gate10inter5, gate10inter6, gate10inter7, gate10inter8, gate10inter9, gate10inter10, gate10inter11, gate10inter12, gate145inter0, gate145inter1, gate145inter2, gate145inter3, gate145inter4, gate145inter5, gate145inter6, gate145inter7, gate145inter8, gate145inter9, gate145inter10, gate145inter11, gate145inter12, gate99inter0, gate99inter1, gate99inter2, gate99inter3, gate99inter4, gate99inter5, gate99inter6, gate99inter7, gate99inter8, gate99inter9, gate99inter10, gate99inter11, gate99inter12, gate462inter0, gate462inter1, gate462inter2, gate462inter3, gate462inter4, gate462inter5, gate462inter6, gate462inter7, gate462inter8, gate462inter9, gate462inter10, gate462inter11, gate462inter12, gate57inter0, gate57inter1, gate57inter2, gate57inter3, gate57inter4, gate57inter5, gate57inter6, gate57inter7, gate57inter8, gate57inter9, gate57inter10, gate57inter11, gate57inter12, gate36inter0, gate36inter1, gate36inter2, gate36inter3, gate36inter4, gate36inter5, gate36inter6, gate36inter7, gate36inter8, gate36inter9, gate36inter10, gate36inter11, gate36inter12, gate110inter0, gate110inter1, gate110inter2, gate110inter3, gate110inter4, gate110inter5, gate110inter6, gate110inter7, gate110inter8, gate110inter9, gate110inter10, gate110inter11, gate110inter12, gate75inter0, gate75inter1, gate75inter2, gate75inter3, gate75inter4, gate75inter5, gate75inter6, gate75inter7, gate75inter8, gate75inter9, gate75inter10, gate75inter11, gate75inter12, gate146inter0, gate146inter1, gate146inter2, gate146inter3, gate146inter4, gate146inter5, gate146inter6, gate146inter7, gate146inter8, gate146inter9, gate146inter10, gate146inter11, gate146inter12, gate96inter0, gate96inter1, gate96inter2, gate96inter3, gate96inter4, gate96inter5, gate96inter6, gate96inter7, gate96inter8, gate96inter9, gate96inter10, gate96inter11, gate96inter12, gate53inter0, gate53inter1, gate53inter2, gate53inter3, gate53inter4, gate53inter5, gate53inter6, gate53inter7, gate53inter8, gate53inter9, gate53inter10, gate53inter11, gate53inter12, gate84inter0, gate84inter1, gate84inter2, gate84inter3, gate84inter4, gate84inter5, gate84inter6, gate84inter7, gate84inter8, gate84inter9, gate84inter10, gate84inter11, gate84inter12, gate295inter0, gate295inter1, gate295inter2, gate295inter3, gate295inter4, gate295inter5, gate295inter6, gate295inter7, gate295inter8, gate295inter9, gate295inter10, gate295inter11, gate295inter12, gate292inter0, gate292inter1, gate292inter2, gate292inter3, gate292inter4, gate292inter5, gate292inter6, gate292inter7, gate292inter8, gate292inter9, gate292inter10, gate292inter11, gate292inter12, gate413inter0, gate413inter1, gate413inter2, gate413inter3, gate413inter4, gate413inter5, gate413inter6, gate413inter7, gate413inter8, gate413inter9, gate413inter10, gate413inter11, gate413inter12, gate428inter0, gate428inter1, gate428inter2, gate428inter3, gate428inter4, gate428inter5, gate428inter6, gate428inter7, gate428inter8, gate428inter9, gate428inter10, gate428inter11, gate428inter12, gate103inter0, gate103inter1, gate103inter2, gate103inter3, gate103inter4, gate103inter5, gate103inter6, gate103inter7, gate103inter8, gate103inter9, gate103inter10, gate103inter11, gate103inter12, gate136inter0, gate136inter1, gate136inter2, gate136inter3, gate136inter4, gate136inter5, gate136inter6, gate136inter7, gate136inter8, gate136inter9, gate136inter10, gate136inter11, gate136inter12, gate238inter0, gate238inter1, gate238inter2, gate238inter3, gate238inter4, gate238inter5, gate238inter6, gate238inter7, gate238inter8, gate238inter9, gate238inter10, gate238inter11, gate238inter12, gate58inter0, gate58inter1, gate58inter2, gate58inter3, gate58inter4, gate58inter5, gate58inter6, gate58inter7, gate58inter8, gate58inter9, gate58inter10, gate58inter11, gate58inter12, gate288inter0, gate288inter1, gate288inter2, gate288inter3, gate288inter4, gate288inter5, gate288inter6, gate288inter7, gate288inter8, gate288inter9, gate288inter10, gate288inter11, gate288inter12, gate15inter0, gate15inter1, gate15inter2, gate15inter3, gate15inter4, gate15inter5, gate15inter6, gate15inter7, gate15inter8, gate15inter9, gate15inter10, gate15inter11, gate15inter12, gate246inter0, gate246inter1, gate246inter2, gate246inter3, gate246inter4, gate246inter5, gate246inter6, gate246inter7, gate246inter8, gate246inter9, gate246inter10, gate246inter11, gate246inter12, gate139inter0, gate139inter1, gate139inter2, gate139inter3, gate139inter4, gate139inter5, gate139inter6, gate139inter7, gate139inter8, gate139inter9, gate139inter10, gate139inter11, gate139inter12, gate63inter0, gate63inter1, gate63inter2, gate63inter3, gate63inter4, gate63inter5, gate63inter6, gate63inter7, gate63inter8, gate63inter9, gate63inter10, gate63inter11, gate63inter12, gate264inter0, gate264inter1, gate264inter2, gate264inter3, gate264inter4, gate264inter5, gate264inter6, gate264inter7, gate264inter8, gate264inter9, gate264inter10, gate264inter11, gate264inter12, gate27inter0, gate27inter1, gate27inter2, gate27inter3, gate27inter4, gate27inter5, gate27inter6, gate27inter7, gate27inter8, gate27inter9, gate27inter10, gate27inter11, gate27inter12, gate480inter0, gate480inter1, gate480inter2, gate480inter3, gate480inter4, gate480inter5, gate480inter6, gate480inter7, gate480inter8, gate480inter9, gate480inter10, gate480inter11, gate480inter12, gate260inter0, gate260inter1, gate260inter2, gate260inter3, gate260inter4, gate260inter5, gate260inter6, gate260inter7, gate260inter8, gate260inter9, gate260inter10, gate260inter11, gate260inter12, gate507inter0, gate507inter1, gate507inter2, gate507inter3, gate507inter4, gate507inter5, gate507inter6, gate507inter7, gate507inter8, gate507inter9, gate507inter10, gate507inter11, gate507inter12, gate459inter0, gate459inter1, gate459inter2, gate459inter3, gate459inter4, gate459inter5, gate459inter6, gate459inter7, gate459inter8, gate459inter9, gate459inter10, gate459inter11, gate459inter12, gate122inter0, gate122inter1, gate122inter2, gate122inter3, gate122inter4, gate122inter5, gate122inter6, gate122inter7, gate122inter8, gate122inter9, gate122inter10, gate122inter11, gate122inter12, gate83inter0, gate83inter1, gate83inter2, gate83inter3, gate83inter4, gate83inter5, gate83inter6, gate83inter7, gate83inter8, gate83inter9, gate83inter10, gate83inter11, gate83inter12, gate167inter0, gate167inter1, gate167inter2, gate167inter3, gate167inter4, gate167inter5, gate167inter6, gate167inter7, gate167inter8, gate167inter9, gate167inter10, gate167inter11, gate167inter12, gate135inter0, gate135inter1, gate135inter2, gate135inter3, gate135inter4, gate135inter5, gate135inter6, gate135inter7, gate135inter8, gate135inter9, gate135inter10, gate135inter11, gate135inter12, gate293inter0, gate293inter1, gate293inter2, gate293inter3, gate293inter4, gate293inter5, gate293inter6, gate293inter7, gate293inter8, gate293inter9, gate293inter10, gate293inter11, gate293inter12, gate392inter0, gate392inter1, gate392inter2, gate392inter3, gate392inter4, gate392inter5, gate392inter6, gate392inter7, gate392inter8, gate392inter9, gate392inter10, gate392inter11, gate392inter12, gate22inter0, gate22inter1, gate22inter2, gate22inter3, gate22inter4, gate22inter5, gate22inter6, gate22inter7, gate22inter8, gate22inter9, gate22inter10, gate22inter11, gate22inter12, gate421inter0, gate421inter1, gate421inter2, gate421inter3, gate421inter4, gate421inter5, gate421inter6, gate421inter7, gate421inter8, gate421inter9, gate421inter10, gate421inter11, gate421inter12, gate132inter0, gate132inter1, gate132inter2, gate132inter3, gate132inter4, gate132inter5, gate132inter6, gate132inter7, gate132inter8, gate132inter9, gate132inter10, gate132inter11, gate132inter12, gate405inter0, gate405inter1, gate405inter2, gate405inter3, gate405inter4, gate405inter5, gate405inter6, gate405inter7, gate405inter8, gate405inter9, gate405inter10, gate405inter11, gate405inter12, gate446inter0, gate446inter1, gate446inter2, gate446inter3, gate446inter4, gate446inter5, gate446inter6, gate446inter7, gate446inter8, gate446inter9, gate446inter10, gate446inter11, gate446inter12, gate21inter0, gate21inter1, gate21inter2, gate21inter3, gate21inter4, gate21inter5, gate21inter6, gate21inter7, gate21inter8, gate21inter9, gate21inter10, gate21inter11, gate21inter12, gate201inter0, gate201inter1, gate201inter2, gate201inter3, gate201inter4, gate201inter5, gate201inter6, gate201inter7, gate201inter8, gate201inter9, gate201inter10, gate201inter11, gate201inter12, gate206inter0, gate206inter1, gate206inter2, gate206inter3, gate206inter4, gate206inter5, gate206inter6, gate206inter7, gate206inter8, gate206inter9, gate206inter10, gate206inter11, gate206inter12, gate118inter0, gate118inter1, gate118inter2, gate118inter3, gate118inter4, gate118inter5, gate118inter6, gate118inter7, gate118inter8, gate118inter9, gate118inter10, gate118inter11, gate118inter12, gate66inter0, gate66inter1, gate66inter2, gate66inter3, gate66inter4, gate66inter5, gate66inter6, gate66inter7, gate66inter8, gate66inter9, gate66inter10, gate66inter11, gate66inter12, gate394inter0, gate394inter1, gate394inter2, gate394inter3, gate394inter4, gate394inter5, gate394inter6, gate394inter7, gate394inter8, gate394inter9, gate394inter10, gate394inter11, gate394inter12, gate236inter0, gate236inter1, gate236inter2, gate236inter3, gate236inter4, gate236inter5, gate236inter6, gate236inter7, gate236inter8, gate236inter9, gate236inter10, gate236inter11, gate236inter12, gate481inter0, gate481inter1, gate481inter2, gate481inter3, gate481inter4, gate481inter5, gate481inter6, gate481inter7, gate481inter8, gate481inter9, gate481inter10, gate481inter11, gate481inter12, gate389inter0, gate389inter1, gate389inter2, gate389inter3, gate389inter4, gate389inter5, gate389inter6, gate389inter7, gate389inter8, gate389inter9, gate389inter10, gate389inter11, gate389inter12, gate49inter0, gate49inter1, gate49inter2, gate49inter3, gate49inter4, gate49inter5, gate49inter6, gate49inter7, gate49inter8, gate49inter9, gate49inter10, gate49inter11, gate49inter12, gate162inter0, gate162inter1, gate162inter2, gate162inter3, gate162inter4, gate162inter5, gate162inter6, gate162inter7, gate162inter8, gate162inter9, gate162inter10, gate162inter11, gate162inter12, gate239inter0, gate239inter1, gate239inter2, gate239inter3, gate239inter4, gate239inter5, gate239inter6, gate239inter7, gate239inter8, gate239inter9, gate239inter10, gate239inter11, gate239inter12, gate218inter0, gate218inter1, gate218inter2, gate218inter3, gate218inter4, gate218inter5, gate218inter6, gate218inter7, gate218inter8, gate218inter9, gate218inter10, gate218inter11, gate218inter12, gate207inter0, gate207inter1, gate207inter2, gate207inter3, gate207inter4, gate207inter5, gate207inter6, gate207inter7, gate207inter8, gate207inter9, gate207inter10, gate207inter11, gate207inter12, gate466inter0, gate466inter1, gate466inter2, gate466inter3, gate466inter4, gate466inter5, gate466inter6, gate466inter7, gate466inter8, gate466inter9, gate466inter10, gate466inter11, gate466inter12, gate489inter0, gate489inter1, gate489inter2, gate489inter3, gate489inter4, gate489inter5, gate489inter6, gate489inter7, gate489inter8, gate489inter9, gate489inter10, gate489inter11, gate489inter12, gate469inter0, gate469inter1, gate469inter2, gate469inter3, gate469inter4, gate469inter5, gate469inter6, gate469inter7, gate469inter8, gate469inter9, gate469inter10, gate469inter11, gate469inter12, gate60inter0, gate60inter1, gate60inter2, gate60inter3, gate60inter4, gate60inter5, gate60inter6, gate60inter7, gate60inter8, gate60inter9, gate60inter10, gate60inter11, gate60inter12, gate18inter0, gate18inter1, gate18inter2, gate18inter3, gate18inter4, gate18inter5, gate18inter6, gate18inter7, gate18inter8, gate18inter9, gate18inter10, gate18inter11, gate18inter12, gate439inter0, gate439inter1, gate439inter2, gate439inter3, gate439inter4, gate439inter5, gate439inter6, gate439inter7, gate439inter8, gate439inter9, gate439inter10, gate439inter11, gate439inter12, gate280inter0, gate280inter1, gate280inter2, gate280inter3, gate280inter4, gate280inter5, gate280inter6, gate280inter7, gate280inter8, gate280inter9, gate280inter10, gate280inter11, gate280inter12, gate101inter0, gate101inter1, gate101inter2, gate101inter3, gate101inter4, gate101inter5, gate101inter6, gate101inter7, gate101inter8, gate101inter9, gate101inter10, gate101inter11, gate101inter12, gate159inter0, gate159inter1, gate159inter2, gate159inter3, gate159inter4, gate159inter5, gate159inter6, gate159inter7, gate159inter8, gate159inter9, gate159inter10, gate159inter11, gate159inter12, gate409inter0, gate409inter1, gate409inter2, gate409inter3, gate409inter4, gate409inter5, gate409inter6, gate409inter7, gate409inter8, gate409inter9, gate409inter10, gate409inter11, gate409inter12, gate448inter0, gate448inter1, gate448inter2, gate448inter3, gate448inter4, gate448inter5, gate448inter6, gate448inter7, gate448inter8, gate448inter9, gate448inter10, gate448inter11, gate448inter12, gate187inter0, gate187inter1, gate187inter2, gate187inter3, gate187inter4, gate187inter5, gate187inter6, gate187inter7, gate187inter8, gate187inter9, gate187inter10, gate187inter11, gate187inter12, gate194inter0, gate194inter1, gate194inter2, gate194inter3, gate194inter4, gate194inter5, gate194inter6, gate194inter7, gate194inter8, gate194inter9, gate194inter10, gate194inter11, gate194inter12, gate410inter0, gate410inter1, gate410inter2, gate410inter3, gate410inter4, gate410inter5, gate410inter6, gate410inter7, gate410inter8, gate410inter9, gate410inter10, gate410inter11, gate410inter12, gate147inter0, gate147inter1, gate147inter2, gate147inter3, gate147inter4, gate147inter5, gate147inter6, gate147inter7, gate147inter8, gate147inter9, gate147inter10, gate147inter11, gate147inter12, gate129inter0, gate129inter1, gate129inter2, gate129inter3, gate129inter4, gate129inter5, gate129inter6, gate129inter7, gate129inter8, gate129inter9, gate129inter10, gate129inter11, gate129inter12, gate277inter0, gate277inter1, gate277inter2, gate277inter3, gate277inter4, gate277inter5, gate277inter6, gate277inter7, gate277inter8, gate277inter9, gate277inter10, gate277inter11, gate277inter12, gate486inter0, gate486inter1, gate486inter2, gate486inter3, gate486inter4, gate486inter5, gate486inter6, gate486inter7, gate486inter8, gate486inter9, gate486inter10, gate486inter11, gate486inter12, gate74inter0, gate74inter1, gate74inter2, gate74inter3, gate74inter4, gate74inter5, gate74inter6, gate74inter7, gate74inter8, gate74inter9, gate74inter10, gate74inter11, gate74inter12, gate470inter0, gate470inter1, gate470inter2, gate470inter3, gate470inter4, gate470inter5, gate470inter6, gate470inter7, gate470inter8, gate470inter9, gate470inter10, gate470inter11, gate470inter12, gate396inter0, gate396inter1, gate396inter2, gate396inter3, gate396inter4, gate396inter5, gate396inter6, gate396inter7, gate396inter8, gate396inter9, gate396inter10, gate396inter11, gate396inter12, gate144inter0, gate144inter1, gate144inter2, gate144inter3, gate144inter4, gate144inter5, gate144inter6, gate144inter7, gate144inter8, gate144inter9, gate144inter10, gate144inter11, gate144inter12, gate412inter0, gate412inter1, gate412inter2, gate412inter3, gate412inter4, gate412inter5, gate412inter6, gate412inter7, gate412inter8, gate412inter9, gate412inter10, gate412inter11, gate412inter12, gate427inter0, gate427inter1, gate427inter2, gate427inter3, gate427inter4, gate427inter5, gate427inter6, gate427inter7, gate427inter8, gate427inter9, gate427inter10, gate427inter11, gate427inter12, gate126inter0, gate126inter1, gate126inter2, gate126inter3, gate126inter4, gate126inter5, gate126inter6, gate126inter7, gate126inter8, gate126inter9, gate126inter10, gate126inter11, gate126inter12, gate514inter0, gate514inter1, gate514inter2, gate514inter3, gate514inter4, gate514inter5, gate514inter6, gate514inter7, gate514inter8, gate514inter9, gate514inter10, gate514inter11, gate514inter12, gate11inter0, gate11inter1, gate11inter2, gate11inter3, gate11inter4, gate11inter5, gate11inter6, gate11inter7, gate11inter8, gate11inter9, gate11inter10, gate11inter11, gate11inter12, gate48inter0, gate48inter1, gate48inter2, gate48inter3, gate48inter4, gate48inter5, gate48inter6, gate48inter7, gate48inter8, gate48inter9, gate48inter10, gate48inter11, gate48inter12, gate141inter0, gate141inter1, gate141inter2, gate141inter3, gate141inter4, gate141inter5, gate141inter6, gate141inter7, gate141inter8, gate141inter9, gate141inter10, gate141inter11, gate141inter12, gate495inter0, gate495inter1, gate495inter2, gate495inter3, gate495inter4, gate495inter5, gate495inter6, gate495inter7, gate495inter8, gate495inter9, gate495inter10, gate495inter11, gate495inter12, gate9inter0, gate9inter1, gate9inter2, gate9inter3, gate9inter4, gate9inter5, gate9inter6, gate9inter7, gate9inter8, gate9inter9, gate9inter10, gate9inter11, gate9inter12, gate102inter0, gate102inter1, gate102inter2, gate102inter3, gate102inter4, gate102inter5, gate102inter6, gate102inter7, gate102inter8, gate102inter9, gate102inter10, gate102inter11, gate102inter12, gate69inter0, gate69inter1, gate69inter2, gate69inter3, gate69inter4, gate69inter5, gate69inter6, gate69inter7, gate69inter8, gate69inter9, gate69inter10, gate69inter11, gate69inter12, gate45inter0, gate45inter1, gate45inter2, gate45inter3, gate45inter4, gate45inter5, gate45inter6, gate45inter7, gate45inter8, gate45inter9, gate45inter10, gate45inter11, gate45inter12, gate71inter0, gate71inter1, gate71inter2, gate71inter3, gate71inter4, gate71inter5, gate71inter6, gate71inter7, gate71inter8, gate71inter9, gate71inter10, gate71inter11, gate71inter12, gate24inter0, gate24inter1, gate24inter2, gate24inter3, gate24inter4, gate24inter5, gate24inter6, gate24inter7, gate24inter8, gate24inter9, gate24inter10, gate24inter11, gate24inter12, gate221inter0, gate221inter1, gate221inter2, gate221inter3, gate221inter4, gate221inter5, gate221inter6, gate221inter7, gate221inter8, gate221inter9, gate221inter10, gate221inter11, gate221inter12, gate39inter0, gate39inter1, gate39inter2, gate39inter3, gate39inter4, gate39inter5, gate39inter6, gate39inter7, gate39inter8, gate39inter9, gate39inter10, gate39inter11, gate39inter12, gate494inter0, gate494inter1, gate494inter2, gate494inter3, gate494inter4, gate494inter5, gate494inter6, gate494inter7, gate494inter8, gate494inter9, gate494inter10, gate494inter11, gate494inter12, gate511inter0, gate511inter1, gate511inter2, gate511inter3, gate511inter4, gate511inter5, gate511inter6, gate511inter7, gate511inter8, gate511inter9, gate511inter10, gate511inter11, gate511inter12, gate443inter0, gate443inter1, gate443inter2, gate443inter3, gate443inter4, gate443inter5, gate443inter6, gate443inter7, gate443inter8, gate443inter9, gate443inter10, gate443inter11, gate443inter12, gate286inter0, gate286inter1, gate286inter2, gate286inter3, gate286inter4, gate286inter5, gate286inter6, gate286inter7, gate286inter8, gate286inter9, gate286inter10, gate286inter11, gate286inter12, gate426inter0, gate426inter1, gate426inter2, gate426inter3, gate426inter4, gate426inter5, gate426inter6, gate426inter7, gate426inter8, gate426inter9, gate426inter10, gate426inter11, gate426inter12, gate497inter0, gate497inter1, gate497inter2, gate497inter3, gate497inter4, gate497inter5, gate497inter6, gate497inter7, gate497inter8, gate497inter9, gate497inter10, gate497inter11, gate497inter12, gate425inter0, gate425inter1, gate425inter2, gate425inter3, gate425inter4, gate425inter5, gate425inter6, gate425inter7, gate425inter8, gate425inter9, gate425inter10, gate425inter11, gate425inter12, gate416inter0, gate416inter1, gate416inter2, gate416inter3, gate416inter4, gate416inter5, gate416inter6, gate416inter7, gate416inter8, gate416inter9, gate416inter10, gate416inter11, gate416inter12, gate262inter0, gate262inter1, gate262inter2, gate262inter3, gate262inter4, gate262inter5, gate262inter6, gate262inter7, gate262inter8, gate262inter9, gate262inter10, gate262inter11, gate262inter12, gate252inter0, gate252inter1, gate252inter2, gate252inter3, gate252inter4, gate252inter5, gate252inter6, gate252inter7, gate252inter8, gate252inter9, gate252inter10, gate252inter11, gate252inter12, gate498inter0, gate498inter1, gate498inter2, gate498inter3, gate498inter4, gate498inter5, gate498inter6, gate498inter7, gate498inter8, gate498inter9, gate498inter10, gate498inter11, gate498inter12, gate93inter0, gate93inter1, gate93inter2, gate93inter3, gate93inter4, gate93inter5, gate93inter6, gate93inter7, gate93inter8, gate93inter9, gate93inter10, gate93inter11, gate93inter12, gate278inter0, gate278inter1, gate278inter2, gate278inter3, gate278inter4, gate278inter5, gate278inter6, gate278inter7, gate278inter8, gate278inter9, gate278inter10, gate278inter11, gate278inter12, gate415inter0, gate415inter1, gate415inter2, gate415inter3, gate415inter4, gate415inter5, gate415inter6, gate415inter7, gate415inter8, gate415inter9, gate415inter10, gate415inter11, gate415inter12, gate88inter0, gate88inter1, gate88inter2, gate88inter3, gate88inter4, gate88inter5, gate88inter6, gate88inter7, gate88inter8, gate88inter9, gate88inter10, gate88inter11, gate88inter12, gate251inter0, gate251inter1, gate251inter2, gate251inter3, gate251inter4, gate251inter5, gate251inter6, gate251inter7, gate251inter8, gate251inter9, gate251inter10, gate251inter11, gate251inter12, gate270inter0, gate270inter1, gate270inter2, gate270inter3, gate270inter4, gate270inter5, gate270inter6, gate270inter7, gate270inter8, gate270inter9, gate270inter10, gate270inter11, gate270inter12, gate13inter0, gate13inter1, gate13inter2, gate13inter3, gate13inter4, gate13inter5, gate13inter6, gate13inter7, gate13inter8, gate13inter9, gate13inter10, gate13inter11, gate13inter12, gate438inter0, gate438inter1, gate438inter2, gate438inter3, gate438inter4, gate438inter5, gate438inter6, gate438inter7, gate438inter8, gate438inter9, gate438inter10, gate438inter11, gate438inter12, gate98inter0, gate98inter1, gate98inter2, gate98inter3, gate98inter4, gate98inter5, gate98inter6, gate98inter7, gate98inter8, gate98inter9, gate98inter10, gate98inter11, gate98inter12, gate505inter0, gate505inter1, gate505inter2, gate505inter3, gate505inter4, gate505inter5, gate505inter6, gate505inter7, gate505inter8, gate505inter9, gate505inter10, gate505inter11, gate505inter12, gate164inter0, gate164inter1, gate164inter2, gate164inter3, gate164inter4, gate164inter5, gate164inter6, gate164inter7, gate164inter8, gate164inter9, gate164inter10, gate164inter11, gate164inter12, gate493inter0, gate493inter1, gate493inter2, gate493inter3, gate493inter4, gate493inter5, gate493inter6, gate493inter7, gate493inter8, gate493inter9, gate493inter10, gate493inter11, gate493inter12, gate166inter0, gate166inter1, gate166inter2, gate166inter3, gate166inter4, gate166inter5, gate166inter6, gate166inter7, gate166inter8, gate166inter9, gate166inter10, gate166inter11, gate166inter12, gate154inter0, gate154inter1, gate154inter2, gate154inter3, gate154inter4, gate154inter5, gate154inter6, gate154inter7, gate154inter8, gate154inter9, gate154inter10, gate154inter11, gate154inter12, gate152inter0, gate152inter1, gate152inter2, gate152inter3, gate152inter4, gate152inter5, gate152inter6, gate152inter7, gate152inter8, gate152inter9, gate152inter10, gate152inter11, gate152inter12, gate492inter0, gate492inter1, gate492inter2, gate492inter3, gate492inter4, gate492inter5, gate492inter6, gate492inter7, gate492inter8, gate492inter9, gate492inter10, gate492inter11, gate492inter12, gate192inter0, gate192inter1, gate192inter2, gate192inter3, gate192inter4, gate192inter5, gate192inter6, gate192inter7, gate192inter8, gate192inter9, gate192inter10, gate192inter11, gate192inter12, gate117inter0, gate117inter1, gate117inter2, gate117inter3, gate117inter4, gate117inter5, gate117inter6, gate117inter7, gate117inter8, gate117inter9, gate117inter10, gate117inter11, gate117inter12, gate138inter0, gate138inter1, gate138inter2, gate138inter3, gate138inter4, gate138inter5, gate138inter6, gate138inter7, gate138inter8, gate138inter9, gate138inter10, gate138inter11, gate138inter12, gate231inter0, gate231inter1, gate231inter2, gate231inter3, gate231inter4, gate231inter5, gate231inter6, gate231inter7, gate231inter8, gate231inter9, gate231inter10, gate231inter11, gate231inter12, gate393inter0, gate393inter1, gate393inter2, gate393inter3, gate393inter4, gate393inter5, gate393inter6, gate393inter7, gate393inter8, gate393inter9, gate393inter10, gate393inter11, gate393inter12, gate33inter0, gate33inter1, gate33inter2, gate33inter3, gate33inter4, gate33inter5, gate33inter6, gate33inter7, gate33inter8, gate33inter9, gate33inter10, gate33inter11, gate33inter12, gate485inter0, gate485inter1, gate485inter2, gate485inter3, gate485inter4, gate485inter5, gate485inter6, gate485inter7, gate485inter8, gate485inter9, gate485inter10, gate485inter11, gate485inter12, gate290inter0, gate290inter1, gate290inter2, gate290inter3, gate290inter4, gate290inter5, gate290inter6, gate290inter7, gate290inter8, gate290inter9, gate290inter10, gate290inter11, gate290inter12, gate230inter0, gate230inter1, gate230inter2, gate230inter3, gate230inter4, gate230inter5, gate230inter6, gate230inter7, gate230inter8, gate230inter9, gate230inter10, gate230inter11, gate230inter12, gate211inter0, gate211inter1, gate211inter2, gate211inter3, gate211inter4, gate211inter5, gate211inter6, gate211inter7, gate211inter8, gate211inter9, gate211inter10, gate211inter11, gate211inter12, gate483inter0, gate483inter1, gate483inter2, gate483inter3, gate483inter4, gate483inter5, gate483inter6, gate483inter7, gate483inter8, gate483inter9, gate483inter10, gate483inter11, gate483inter12, gate131inter0, gate131inter1, gate131inter2, gate131inter3, gate131inter4, gate131inter5, gate131inter6, gate131inter7, gate131inter8, gate131inter9, gate131inter10, gate131inter11, gate131inter12, gate488inter0, gate488inter1, gate488inter2, gate488inter3, gate488inter4, gate488inter5, gate488inter6, gate488inter7, gate488inter8, gate488inter9, gate488inter10, gate488inter11, gate488inter12, gate30inter0, gate30inter1, gate30inter2, gate30inter3, gate30inter4, gate30inter5, gate30inter6, gate30inter7, gate30inter8, gate30inter9, gate30inter10, gate30inter11, gate30inter12, gate268inter0, gate268inter1, gate268inter2, gate268inter3, gate268inter4, gate268inter5, gate268inter6, gate268inter7, gate268inter8, gate268inter9, gate268inter10, gate268inter11, gate268inter12, gate112inter0, gate112inter1, gate112inter2, gate112inter3, gate112inter4, gate112inter5, gate112inter6, gate112inter7, gate112inter8, gate112inter9, gate112inter10, gate112inter11, gate112inter12, gate168inter0, gate168inter1, gate168inter2, gate168inter3, gate168inter4, gate168inter5, gate168inter6, gate168inter7, gate168inter8, gate168inter9, gate168inter10, gate168inter11, gate168inter12, gate55inter0, gate55inter1, gate55inter2, gate55inter3, gate55inter4, gate55inter5, gate55inter6, gate55inter7, gate55inter8, gate55inter9, gate55inter10, gate55inter11, gate55inter12, gate78inter0, gate78inter1, gate78inter2, gate78inter3, gate78inter4, gate78inter5, gate78inter6, gate78inter7, gate78inter8, gate78inter9, gate78inter10, gate78inter11, gate78inter12;



and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );

  xor2  gate2255(.a(G2), .b(G1), .O(gate9inter0));
  nand2 gate2256(.a(gate9inter0), .b(s_244), .O(gate9inter1));
  and2  gate2257(.a(G2), .b(G1), .O(gate9inter2));
  inv1  gate2258(.a(s_244), .O(gate9inter3));
  inv1  gate2259(.a(s_245), .O(gate9inter4));
  nand2 gate2260(.a(gate9inter4), .b(gate9inter3), .O(gate9inter5));
  nor2  gate2261(.a(gate9inter5), .b(gate9inter2), .O(gate9inter6));
  inv1  gate2262(.a(G1), .O(gate9inter7));
  inv1  gate2263(.a(G2), .O(gate9inter8));
  nand2 gate2264(.a(gate9inter8), .b(gate9inter7), .O(gate9inter9));
  nand2 gate2265(.a(s_245), .b(gate9inter3), .O(gate9inter10));
  nor2  gate2266(.a(gate9inter10), .b(gate9inter9), .O(gate9inter11));
  nor2  gate2267(.a(gate9inter11), .b(gate9inter6), .O(gate9inter12));
  nand2 gate2268(.a(gate9inter12), .b(gate9inter1), .O(G266));

  xor2  gate1051(.a(G4), .b(G3), .O(gate10inter0));
  nand2 gate1052(.a(gate10inter0), .b(s_72), .O(gate10inter1));
  and2  gate1053(.a(G4), .b(G3), .O(gate10inter2));
  inv1  gate1054(.a(s_72), .O(gate10inter3));
  inv1  gate1055(.a(s_73), .O(gate10inter4));
  nand2 gate1056(.a(gate10inter4), .b(gate10inter3), .O(gate10inter5));
  nor2  gate1057(.a(gate10inter5), .b(gate10inter2), .O(gate10inter6));
  inv1  gate1058(.a(G3), .O(gate10inter7));
  inv1  gate1059(.a(G4), .O(gate10inter8));
  nand2 gate1060(.a(gate10inter8), .b(gate10inter7), .O(gate10inter9));
  nand2 gate1061(.a(s_73), .b(gate10inter3), .O(gate10inter10));
  nor2  gate1062(.a(gate10inter10), .b(gate10inter9), .O(gate10inter11));
  nor2  gate1063(.a(gate10inter11), .b(gate10inter6), .O(gate10inter12));
  nand2 gate1064(.a(gate10inter12), .b(gate10inter1), .O(G269));

  xor2  gate2199(.a(G6), .b(G5), .O(gate11inter0));
  nand2 gate2200(.a(gate11inter0), .b(s_236), .O(gate11inter1));
  and2  gate2201(.a(G6), .b(G5), .O(gate11inter2));
  inv1  gate2202(.a(s_236), .O(gate11inter3));
  inv1  gate2203(.a(s_237), .O(gate11inter4));
  nand2 gate2204(.a(gate11inter4), .b(gate11inter3), .O(gate11inter5));
  nor2  gate2205(.a(gate11inter5), .b(gate11inter2), .O(gate11inter6));
  inv1  gate2206(.a(G5), .O(gate11inter7));
  inv1  gate2207(.a(G6), .O(gate11inter8));
  nand2 gate2208(.a(gate11inter8), .b(gate11inter7), .O(gate11inter9));
  nand2 gate2209(.a(s_237), .b(gate11inter3), .O(gate11inter10));
  nor2  gate2210(.a(gate11inter10), .b(gate11inter9), .O(gate11inter11));
  nor2  gate2211(.a(gate11inter11), .b(gate11inter6), .O(gate11inter12));
  nand2 gate2212(.a(gate11inter12), .b(gate11inter1), .O(G272));
nand2 gate12( .a(G7), .b(G8), .O(G275) );

  xor2  gate2605(.a(G10), .b(G9), .O(gate13inter0));
  nand2 gate2606(.a(gate13inter0), .b(s_294), .O(gate13inter1));
  and2  gate2607(.a(G10), .b(G9), .O(gate13inter2));
  inv1  gate2608(.a(s_294), .O(gate13inter3));
  inv1  gate2609(.a(s_295), .O(gate13inter4));
  nand2 gate2610(.a(gate13inter4), .b(gate13inter3), .O(gate13inter5));
  nor2  gate2611(.a(gate13inter5), .b(gate13inter2), .O(gate13inter6));
  inv1  gate2612(.a(G9), .O(gate13inter7));
  inv1  gate2613(.a(G10), .O(gate13inter8));
  nand2 gate2614(.a(gate13inter8), .b(gate13inter7), .O(gate13inter9));
  nand2 gate2615(.a(s_295), .b(gate13inter3), .O(gate13inter10));
  nor2  gate2616(.a(gate13inter10), .b(gate13inter9), .O(gate13inter11));
  nor2  gate2617(.a(gate13inter11), .b(gate13inter6), .O(gate13inter12));
  nand2 gate2618(.a(gate13inter12), .b(gate13inter1), .O(G278));
nand2 gate14( .a(G11), .b(G12), .O(G281) );

  xor2  gate1345(.a(G14), .b(G13), .O(gate15inter0));
  nand2 gate1346(.a(gate15inter0), .b(s_114), .O(gate15inter1));
  and2  gate1347(.a(G14), .b(G13), .O(gate15inter2));
  inv1  gate1348(.a(s_114), .O(gate15inter3));
  inv1  gate1349(.a(s_115), .O(gate15inter4));
  nand2 gate1350(.a(gate15inter4), .b(gate15inter3), .O(gate15inter5));
  nor2  gate1351(.a(gate15inter5), .b(gate15inter2), .O(gate15inter6));
  inv1  gate1352(.a(G13), .O(gate15inter7));
  inv1  gate1353(.a(G14), .O(gate15inter8));
  nand2 gate1354(.a(gate15inter8), .b(gate15inter7), .O(gate15inter9));
  nand2 gate1355(.a(s_115), .b(gate15inter3), .O(gate15inter10));
  nor2  gate1356(.a(gate15inter10), .b(gate15inter9), .O(gate15inter11));
  nor2  gate1357(.a(gate15inter11), .b(gate15inter6), .O(gate15inter12));
  nand2 gate1358(.a(gate15inter12), .b(gate15inter1), .O(G284));

  xor2  gate869(.a(G16), .b(G15), .O(gate16inter0));
  nand2 gate870(.a(gate16inter0), .b(s_46), .O(gate16inter1));
  and2  gate871(.a(G16), .b(G15), .O(gate16inter2));
  inv1  gate872(.a(s_46), .O(gate16inter3));
  inv1  gate873(.a(s_47), .O(gate16inter4));
  nand2 gate874(.a(gate16inter4), .b(gate16inter3), .O(gate16inter5));
  nor2  gate875(.a(gate16inter5), .b(gate16inter2), .O(gate16inter6));
  inv1  gate876(.a(G15), .O(gate16inter7));
  inv1  gate877(.a(G16), .O(gate16inter8));
  nand2 gate878(.a(gate16inter8), .b(gate16inter7), .O(gate16inter9));
  nand2 gate879(.a(s_47), .b(gate16inter3), .O(gate16inter10));
  nor2  gate880(.a(gate16inter10), .b(gate16inter9), .O(gate16inter11));
  nor2  gate881(.a(gate16inter11), .b(gate16inter6), .O(gate16inter12));
  nand2 gate882(.a(gate16inter12), .b(gate16inter1), .O(G287));
nand2 gate17( .a(G17), .b(G18), .O(G290) );

  xor2  gate1891(.a(G20), .b(G19), .O(gate18inter0));
  nand2 gate1892(.a(gate18inter0), .b(s_192), .O(gate18inter1));
  and2  gate1893(.a(G20), .b(G19), .O(gate18inter2));
  inv1  gate1894(.a(s_192), .O(gate18inter3));
  inv1  gate1895(.a(s_193), .O(gate18inter4));
  nand2 gate1896(.a(gate18inter4), .b(gate18inter3), .O(gate18inter5));
  nor2  gate1897(.a(gate18inter5), .b(gate18inter2), .O(gate18inter6));
  inv1  gate1898(.a(G19), .O(gate18inter7));
  inv1  gate1899(.a(G20), .O(gate18inter8));
  nand2 gate1900(.a(gate18inter8), .b(gate18inter7), .O(gate18inter9));
  nand2 gate1901(.a(s_193), .b(gate18inter3), .O(gate18inter10));
  nor2  gate1902(.a(gate18inter10), .b(gate18inter9), .O(gate18inter11));
  nor2  gate1903(.a(gate18inter11), .b(gate18inter6), .O(gate18inter12));
  nand2 gate1904(.a(gate18inter12), .b(gate18inter1), .O(G293));
nand2 gate19( .a(G21), .b(G22), .O(G296) );
nand2 gate20( .a(G23), .b(G24), .O(G299) );

  xor2  gate1639(.a(G26), .b(G25), .O(gate21inter0));
  nand2 gate1640(.a(gate21inter0), .b(s_156), .O(gate21inter1));
  and2  gate1641(.a(G26), .b(G25), .O(gate21inter2));
  inv1  gate1642(.a(s_156), .O(gate21inter3));
  inv1  gate1643(.a(s_157), .O(gate21inter4));
  nand2 gate1644(.a(gate21inter4), .b(gate21inter3), .O(gate21inter5));
  nor2  gate1645(.a(gate21inter5), .b(gate21inter2), .O(gate21inter6));
  inv1  gate1646(.a(G25), .O(gate21inter7));
  inv1  gate1647(.a(G26), .O(gate21inter8));
  nand2 gate1648(.a(gate21inter8), .b(gate21inter7), .O(gate21inter9));
  nand2 gate1649(.a(s_157), .b(gate21inter3), .O(gate21inter10));
  nor2  gate1650(.a(gate21inter10), .b(gate21inter9), .O(gate21inter11));
  nor2  gate1651(.a(gate21inter11), .b(gate21inter6), .O(gate21inter12));
  nand2 gate1652(.a(gate21inter12), .b(gate21inter1), .O(G302));

  xor2  gate1569(.a(G28), .b(G27), .O(gate22inter0));
  nand2 gate1570(.a(gate22inter0), .b(s_146), .O(gate22inter1));
  and2  gate1571(.a(G28), .b(G27), .O(gate22inter2));
  inv1  gate1572(.a(s_146), .O(gate22inter3));
  inv1  gate1573(.a(s_147), .O(gate22inter4));
  nand2 gate1574(.a(gate22inter4), .b(gate22inter3), .O(gate22inter5));
  nor2  gate1575(.a(gate22inter5), .b(gate22inter2), .O(gate22inter6));
  inv1  gate1576(.a(G27), .O(gate22inter7));
  inv1  gate1577(.a(G28), .O(gate22inter8));
  nand2 gate1578(.a(gate22inter8), .b(gate22inter7), .O(gate22inter9));
  nand2 gate1579(.a(s_147), .b(gate22inter3), .O(gate22inter10));
  nor2  gate1580(.a(gate22inter10), .b(gate22inter9), .O(gate22inter11));
  nor2  gate1581(.a(gate22inter11), .b(gate22inter6), .O(gate22inter12));
  nand2 gate1582(.a(gate22inter12), .b(gate22inter1), .O(G305));
nand2 gate23( .a(G29), .b(G30), .O(G308) );

  xor2  gate2325(.a(G32), .b(G31), .O(gate24inter0));
  nand2 gate2326(.a(gate24inter0), .b(s_254), .O(gate24inter1));
  and2  gate2327(.a(G32), .b(G31), .O(gate24inter2));
  inv1  gate2328(.a(s_254), .O(gate24inter3));
  inv1  gate2329(.a(s_255), .O(gate24inter4));
  nand2 gate2330(.a(gate24inter4), .b(gate24inter3), .O(gate24inter5));
  nor2  gate2331(.a(gate24inter5), .b(gate24inter2), .O(gate24inter6));
  inv1  gate2332(.a(G31), .O(gate24inter7));
  inv1  gate2333(.a(G32), .O(gate24inter8));
  nand2 gate2334(.a(gate24inter8), .b(gate24inter7), .O(gate24inter9));
  nand2 gate2335(.a(s_255), .b(gate24inter3), .O(gate24inter10));
  nor2  gate2336(.a(gate24inter10), .b(gate24inter9), .O(gate24inter11));
  nor2  gate2337(.a(gate24inter11), .b(gate24inter6), .O(gate24inter12));
  nand2 gate2338(.a(gate24inter12), .b(gate24inter1), .O(G311));
nand2 gate25( .a(G1), .b(G5), .O(G314) );
nand2 gate26( .a(G9), .b(G13), .O(G317) );

  xor2  gate1415(.a(G6), .b(G2), .O(gate27inter0));
  nand2 gate1416(.a(gate27inter0), .b(s_124), .O(gate27inter1));
  and2  gate1417(.a(G6), .b(G2), .O(gate27inter2));
  inv1  gate1418(.a(s_124), .O(gate27inter3));
  inv1  gate1419(.a(s_125), .O(gate27inter4));
  nand2 gate1420(.a(gate27inter4), .b(gate27inter3), .O(gate27inter5));
  nor2  gate1421(.a(gate27inter5), .b(gate27inter2), .O(gate27inter6));
  inv1  gate1422(.a(G2), .O(gate27inter7));
  inv1  gate1423(.a(G6), .O(gate27inter8));
  nand2 gate1424(.a(gate27inter8), .b(gate27inter7), .O(gate27inter9));
  nand2 gate1425(.a(s_125), .b(gate27inter3), .O(gate27inter10));
  nor2  gate1426(.a(gate27inter10), .b(gate27inter9), .O(gate27inter11));
  nor2  gate1427(.a(gate27inter11), .b(gate27inter6), .O(gate27inter12));
  nand2 gate1428(.a(gate27inter12), .b(gate27inter1), .O(G320));
nand2 gate28( .a(G10), .b(G14), .O(G323) );

  xor2  gate841(.a(G7), .b(G3), .O(gate29inter0));
  nand2 gate842(.a(gate29inter0), .b(s_42), .O(gate29inter1));
  and2  gate843(.a(G7), .b(G3), .O(gate29inter2));
  inv1  gate844(.a(s_42), .O(gate29inter3));
  inv1  gate845(.a(s_43), .O(gate29inter4));
  nand2 gate846(.a(gate29inter4), .b(gate29inter3), .O(gate29inter5));
  nor2  gate847(.a(gate29inter5), .b(gate29inter2), .O(gate29inter6));
  inv1  gate848(.a(G3), .O(gate29inter7));
  inv1  gate849(.a(G7), .O(gate29inter8));
  nand2 gate850(.a(gate29inter8), .b(gate29inter7), .O(gate29inter9));
  nand2 gate851(.a(s_43), .b(gate29inter3), .O(gate29inter10));
  nor2  gate852(.a(gate29inter10), .b(gate29inter9), .O(gate29inter11));
  nor2  gate853(.a(gate29inter11), .b(gate29inter6), .O(gate29inter12));
  nand2 gate854(.a(gate29inter12), .b(gate29inter1), .O(G326));

  xor2  gate2927(.a(G15), .b(G11), .O(gate30inter0));
  nand2 gate2928(.a(gate30inter0), .b(s_340), .O(gate30inter1));
  and2  gate2929(.a(G15), .b(G11), .O(gate30inter2));
  inv1  gate2930(.a(s_340), .O(gate30inter3));
  inv1  gate2931(.a(s_341), .O(gate30inter4));
  nand2 gate2932(.a(gate30inter4), .b(gate30inter3), .O(gate30inter5));
  nor2  gate2933(.a(gate30inter5), .b(gate30inter2), .O(gate30inter6));
  inv1  gate2934(.a(G11), .O(gate30inter7));
  inv1  gate2935(.a(G15), .O(gate30inter8));
  nand2 gate2936(.a(gate30inter8), .b(gate30inter7), .O(gate30inter9));
  nand2 gate2937(.a(s_341), .b(gate30inter3), .O(gate30inter10));
  nor2  gate2938(.a(gate30inter10), .b(gate30inter9), .O(gate30inter11));
  nor2  gate2939(.a(gate30inter11), .b(gate30inter6), .O(gate30inter12));
  nand2 gate2940(.a(gate30inter12), .b(gate30inter1), .O(G329));
nand2 gate31( .a(G4), .b(G8), .O(G332) );
nand2 gate32( .a(G12), .b(G16), .O(G335) );

  xor2  gate2815(.a(G21), .b(G17), .O(gate33inter0));
  nand2 gate2816(.a(gate33inter0), .b(s_324), .O(gate33inter1));
  and2  gate2817(.a(G21), .b(G17), .O(gate33inter2));
  inv1  gate2818(.a(s_324), .O(gate33inter3));
  inv1  gate2819(.a(s_325), .O(gate33inter4));
  nand2 gate2820(.a(gate33inter4), .b(gate33inter3), .O(gate33inter5));
  nor2  gate2821(.a(gate33inter5), .b(gate33inter2), .O(gate33inter6));
  inv1  gate2822(.a(G17), .O(gate33inter7));
  inv1  gate2823(.a(G21), .O(gate33inter8));
  nand2 gate2824(.a(gate33inter8), .b(gate33inter7), .O(gate33inter9));
  nand2 gate2825(.a(s_325), .b(gate33inter3), .O(gate33inter10));
  nor2  gate2826(.a(gate33inter10), .b(gate33inter9), .O(gate33inter11));
  nor2  gate2827(.a(gate33inter11), .b(gate33inter6), .O(gate33inter12));
  nand2 gate2828(.a(gate33inter12), .b(gate33inter1), .O(G338));
nand2 gate34( .a(G25), .b(G29), .O(G341) );
nand2 gate35( .a(G18), .b(G22), .O(G344) );

  xor2  gate1121(.a(G30), .b(G26), .O(gate36inter0));
  nand2 gate1122(.a(gate36inter0), .b(s_82), .O(gate36inter1));
  and2  gate1123(.a(G30), .b(G26), .O(gate36inter2));
  inv1  gate1124(.a(s_82), .O(gate36inter3));
  inv1  gate1125(.a(s_83), .O(gate36inter4));
  nand2 gate1126(.a(gate36inter4), .b(gate36inter3), .O(gate36inter5));
  nor2  gate1127(.a(gate36inter5), .b(gate36inter2), .O(gate36inter6));
  inv1  gate1128(.a(G26), .O(gate36inter7));
  inv1  gate1129(.a(G30), .O(gate36inter8));
  nand2 gate1130(.a(gate36inter8), .b(gate36inter7), .O(gate36inter9));
  nand2 gate1131(.a(s_83), .b(gate36inter3), .O(gate36inter10));
  nor2  gate1132(.a(gate36inter10), .b(gate36inter9), .O(gate36inter11));
  nor2  gate1133(.a(gate36inter11), .b(gate36inter6), .O(gate36inter12));
  nand2 gate1134(.a(gate36inter12), .b(gate36inter1), .O(G347));

  xor2  gate925(.a(G23), .b(G19), .O(gate37inter0));
  nand2 gate926(.a(gate37inter0), .b(s_54), .O(gate37inter1));
  and2  gate927(.a(G23), .b(G19), .O(gate37inter2));
  inv1  gate928(.a(s_54), .O(gate37inter3));
  inv1  gate929(.a(s_55), .O(gate37inter4));
  nand2 gate930(.a(gate37inter4), .b(gate37inter3), .O(gate37inter5));
  nor2  gate931(.a(gate37inter5), .b(gate37inter2), .O(gate37inter6));
  inv1  gate932(.a(G19), .O(gate37inter7));
  inv1  gate933(.a(G23), .O(gate37inter8));
  nand2 gate934(.a(gate37inter8), .b(gate37inter7), .O(gate37inter9));
  nand2 gate935(.a(s_55), .b(gate37inter3), .O(gate37inter10));
  nor2  gate936(.a(gate37inter10), .b(gate37inter9), .O(gate37inter11));
  nor2  gate937(.a(gate37inter11), .b(gate37inter6), .O(gate37inter12));
  nand2 gate938(.a(gate37inter12), .b(gate37inter1), .O(G350));

  xor2  gate1023(.a(G31), .b(G27), .O(gate38inter0));
  nand2 gate1024(.a(gate38inter0), .b(s_68), .O(gate38inter1));
  and2  gate1025(.a(G31), .b(G27), .O(gate38inter2));
  inv1  gate1026(.a(s_68), .O(gate38inter3));
  inv1  gate1027(.a(s_69), .O(gate38inter4));
  nand2 gate1028(.a(gate38inter4), .b(gate38inter3), .O(gate38inter5));
  nor2  gate1029(.a(gate38inter5), .b(gate38inter2), .O(gate38inter6));
  inv1  gate1030(.a(G27), .O(gate38inter7));
  inv1  gate1031(.a(G31), .O(gate38inter8));
  nand2 gate1032(.a(gate38inter8), .b(gate38inter7), .O(gate38inter9));
  nand2 gate1033(.a(s_69), .b(gate38inter3), .O(gate38inter10));
  nor2  gate1034(.a(gate38inter10), .b(gate38inter9), .O(gate38inter11));
  nor2  gate1035(.a(gate38inter11), .b(gate38inter6), .O(gate38inter12));
  nand2 gate1036(.a(gate38inter12), .b(gate38inter1), .O(G353));

  xor2  gate2353(.a(G24), .b(G20), .O(gate39inter0));
  nand2 gate2354(.a(gate39inter0), .b(s_258), .O(gate39inter1));
  and2  gate2355(.a(G24), .b(G20), .O(gate39inter2));
  inv1  gate2356(.a(s_258), .O(gate39inter3));
  inv1  gate2357(.a(s_259), .O(gate39inter4));
  nand2 gate2358(.a(gate39inter4), .b(gate39inter3), .O(gate39inter5));
  nor2  gate2359(.a(gate39inter5), .b(gate39inter2), .O(gate39inter6));
  inv1  gate2360(.a(G20), .O(gate39inter7));
  inv1  gate2361(.a(G24), .O(gate39inter8));
  nand2 gate2362(.a(gate39inter8), .b(gate39inter7), .O(gate39inter9));
  nand2 gate2363(.a(s_259), .b(gate39inter3), .O(gate39inter10));
  nor2  gate2364(.a(gate39inter10), .b(gate39inter9), .O(gate39inter11));
  nor2  gate2365(.a(gate39inter11), .b(gate39inter6), .O(gate39inter12));
  nand2 gate2366(.a(gate39inter12), .b(gate39inter1), .O(G356));
nand2 gate40( .a(G28), .b(G32), .O(G359) );
nand2 gate41( .a(G1), .b(G266), .O(G362) );
nand2 gate42( .a(G2), .b(G266), .O(G363) );

  xor2  gate911(.a(G269), .b(G3), .O(gate43inter0));
  nand2 gate912(.a(gate43inter0), .b(s_52), .O(gate43inter1));
  and2  gate913(.a(G269), .b(G3), .O(gate43inter2));
  inv1  gate914(.a(s_52), .O(gate43inter3));
  inv1  gate915(.a(s_53), .O(gate43inter4));
  nand2 gate916(.a(gate43inter4), .b(gate43inter3), .O(gate43inter5));
  nor2  gate917(.a(gate43inter5), .b(gate43inter2), .O(gate43inter6));
  inv1  gate918(.a(G3), .O(gate43inter7));
  inv1  gate919(.a(G269), .O(gate43inter8));
  nand2 gate920(.a(gate43inter8), .b(gate43inter7), .O(gate43inter9));
  nand2 gate921(.a(s_53), .b(gate43inter3), .O(gate43inter10));
  nor2  gate922(.a(gate43inter10), .b(gate43inter9), .O(gate43inter11));
  nor2  gate923(.a(gate43inter11), .b(gate43inter6), .O(gate43inter12));
  nand2 gate924(.a(gate43inter12), .b(gate43inter1), .O(G364));
nand2 gate44( .a(G4), .b(G269), .O(G365) );

  xor2  gate2297(.a(G272), .b(G5), .O(gate45inter0));
  nand2 gate2298(.a(gate45inter0), .b(s_250), .O(gate45inter1));
  and2  gate2299(.a(G272), .b(G5), .O(gate45inter2));
  inv1  gate2300(.a(s_250), .O(gate45inter3));
  inv1  gate2301(.a(s_251), .O(gate45inter4));
  nand2 gate2302(.a(gate45inter4), .b(gate45inter3), .O(gate45inter5));
  nor2  gate2303(.a(gate45inter5), .b(gate45inter2), .O(gate45inter6));
  inv1  gate2304(.a(G5), .O(gate45inter7));
  inv1  gate2305(.a(G272), .O(gate45inter8));
  nand2 gate2306(.a(gate45inter8), .b(gate45inter7), .O(gate45inter9));
  nand2 gate2307(.a(s_251), .b(gate45inter3), .O(gate45inter10));
  nor2  gate2308(.a(gate45inter10), .b(gate45inter9), .O(gate45inter11));
  nor2  gate2309(.a(gate45inter11), .b(gate45inter6), .O(gate45inter12));
  nand2 gate2310(.a(gate45inter12), .b(gate45inter1), .O(G366));
nand2 gate46( .a(G6), .b(G272), .O(G367) );
nand2 gate47( .a(G7), .b(G275), .O(G368) );

  xor2  gate2213(.a(G275), .b(G8), .O(gate48inter0));
  nand2 gate2214(.a(gate48inter0), .b(s_238), .O(gate48inter1));
  and2  gate2215(.a(G275), .b(G8), .O(gate48inter2));
  inv1  gate2216(.a(s_238), .O(gate48inter3));
  inv1  gate2217(.a(s_239), .O(gate48inter4));
  nand2 gate2218(.a(gate48inter4), .b(gate48inter3), .O(gate48inter5));
  nor2  gate2219(.a(gate48inter5), .b(gate48inter2), .O(gate48inter6));
  inv1  gate2220(.a(G8), .O(gate48inter7));
  inv1  gate2221(.a(G275), .O(gate48inter8));
  nand2 gate2222(.a(gate48inter8), .b(gate48inter7), .O(gate48inter9));
  nand2 gate2223(.a(s_239), .b(gate48inter3), .O(gate48inter10));
  nor2  gate2224(.a(gate48inter10), .b(gate48inter9), .O(gate48inter11));
  nor2  gate2225(.a(gate48inter11), .b(gate48inter6), .O(gate48inter12));
  nand2 gate2226(.a(gate48inter12), .b(gate48inter1), .O(G369));

  xor2  gate1765(.a(G278), .b(G9), .O(gate49inter0));
  nand2 gate1766(.a(gate49inter0), .b(s_174), .O(gate49inter1));
  and2  gate1767(.a(G278), .b(G9), .O(gate49inter2));
  inv1  gate1768(.a(s_174), .O(gate49inter3));
  inv1  gate1769(.a(s_175), .O(gate49inter4));
  nand2 gate1770(.a(gate49inter4), .b(gate49inter3), .O(gate49inter5));
  nor2  gate1771(.a(gate49inter5), .b(gate49inter2), .O(gate49inter6));
  inv1  gate1772(.a(G9), .O(gate49inter7));
  inv1  gate1773(.a(G278), .O(gate49inter8));
  nand2 gate1774(.a(gate49inter8), .b(gate49inter7), .O(gate49inter9));
  nand2 gate1775(.a(s_175), .b(gate49inter3), .O(gate49inter10));
  nor2  gate1776(.a(gate49inter10), .b(gate49inter9), .O(gate49inter11));
  nor2  gate1777(.a(gate49inter11), .b(gate49inter6), .O(gate49inter12));
  nand2 gate1778(.a(gate49inter12), .b(gate49inter1), .O(G370));
nand2 gate50( .a(G10), .b(G278), .O(G371) );
nand2 gate51( .a(G11), .b(G281), .O(G372) );
nand2 gate52( .a(G12), .b(G281), .O(G373) );

  xor2  gate1191(.a(G284), .b(G13), .O(gate53inter0));
  nand2 gate1192(.a(gate53inter0), .b(s_92), .O(gate53inter1));
  and2  gate1193(.a(G284), .b(G13), .O(gate53inter2));
  inv1  gate1194(.a(s_92), .O(gate53inter3));
  inv1  gate1195(.a(s_93), .O(gate53inter4));
  nand2 gate1196(.a(gate53inter4), .b(gate53inter3), .O(gate53inter5));
  nor2  gate1197(.a(gate53inter5), .b(gate53inter2), .O(gate53inter6));
  inv1  gate1198(.a(G13), .O(gate53inter7));
  inv1  gate1199(.a(G284), .O(gate53inter8));
  nand2 gate1200(.a(gate53inter8), .b(gate53inter7), .O(gate53inter9));
  nand2 gate1201(.a(s_93), .b(gate53inter3), .O(gate53inter10));
  nor2  gate1202(.a(gate53inter10), .b(gate53inter9), .O(gate53inter11));
  nor2  gate1203(.a(gate53inter11), .b(gate53inter6), .O(gate53inter12));
  nand2 gate1204(.a(gate53inter12), .b(gate53inter1), .O(G374));

  xor2  gate967(.a(G284), .b(G14), .O(gate54inter0));
  nand2 gate968(.a(gate54inter0), .b(s_60), .O(gate54inter1));
  and2  gate969(.a(G284), .b(G14), .O(gate54inter2));
  inv1  gate970(.a(s_60), .O(gate54inter3));
  inv1  gate971(.a(s_61), .O(gate54inter4));
  nand2 gate972(.a(gate54inter4), .b(gate54inter3), .O(gate54inter5));
  nor2  gate973(.a(gate54inter5), .b(gate54inter2), .O(gate54inter6));
  inv1  gate974(.a(G14), .O(gate54inter7));
  inv1  gate975(.a(G284), .O(gate54inter8));
  nand2 gate976(.a(gate54inter8), .b(gate54inter7), .O(gate54inter9));
  nand2 gate977(.a(s_61), .b(gate54inter3), .O(gate54inter10));
  nor2  gate978(.a(gate54inter10), .b(gate54inter9), .O(gate54inter11));
  nor2  gate979(.a(gate54inter11), .b(gate54inter6), .O(gate54inter12));
  nand2 gate980(.a(gate54inter12), .b(gate54inter1), .O(G375));

  xor2  gate2983(.a(G287), .b(G15), .O(gate55inter0));
  nand2 gate2984(.a(gate55inter0), .b(s_348), .O(gate55inter1));
  and2  gate2985(.a(G287), .b(G15), .O(gate55inter2));
  inv1  gate2986(.a(s_348), .O(gate55inter3));
  inv1  gate2987(.a(s_349), .O(gate55inter4));
  nand2 gate2988(.a(gate55inter4), .b(gate55inter3), .O(gate55inter5));
  nor2  gate2989(.a(gate55inter5), .b(gate55inter2), .O(gate55inter6));
  inv1  gate2990(.a(G15), .O(gate55inter7));
  inv1  gate2991(.a(G287), .O(gate55inter8));
  nand2 gate2992(.a(gate55inter8), .b(gate55inter7), .O(gate55inter9));
  nand2 gate2993(.a(s_349), .b(gate55inter3), .O(gate55inter10));
  nor2  gate2994(.a(gate55inter10), .b(gate55inter9), .O(gate55inter11));
  nor2  gate2995(.a(gate55inter11), .b(gate55inter6), .O(gate55inter12));
  nand2 gate2996(.a(gate55inter12), .b(gate55inter1), .O(G376));
nand2 gate56( .a(G16), .b(G287), .O(G377) );

  xor2  gate1107(.a(G290), .b(G17), .O(gate57inter0));
  nand2 gate1108(.a(gate57inter0), .b(s_80), .O(gate57inter1));
  and2  gate1109(.a(G290), .b(G17), .O(gate57inter2));
  inv1  gate1110(.a(s_80), .O(gate57inter3));
  inv1  gate1111(.a(s_81), .O(gate57inter4));
  nand2 gate1112(.a(gate57inter4), .b(gate57inter3), .O(gate57inter5));
  nor2  gate1113(.a(gate57inter5), .b(gate57inter2), .O(gate57inter6));
  inv1  gate1114(.a(G17), .O(gate57inter7));
  inv1  gate1115(.a(G290), .O(gate57inter8));
  nand2 gate1116(.a(gate57inter8), .b(gate57inter7), .O(gate57inter9));
  nand2 gate1117(.a(s_81), .b(gate57inter3), .O(gate57inter10));
  nor2  gate1118(.a(gate57inter10), .b(gate57inter9), .O(gate57inter11));
  nor2  gate1119(.a(gate57inter11), .b(gate57inter6), .O(gate57inter12));
  nand2 gate1120(.a(gate57inter12), .b(gate57inter1), .O(G378));

  xor2  gate1317(.a(G290), .b(G18), .O(gate58inter0));
  nand2 gate1318(.a(gate58inter0), .b(s_110), .O(gate58inter1));
  and2  gate1319(.a(G290), .b(G18), .O(gate58inter2));
  inv1  gate1320(.a(s_110), .O(gate58inter3));
  inv1  gate1321(.a(s_111), .O(gate58inter4));
  nand2 gate1322(.a(gate58inter4), .b(gate58inter3), .O(gate58inter5));
  nor2  gate1323(.a(gate58inter5), .b(gate58inter2), .O(gate58inter6));
  inv1  gate1324(.a(G18), .O(gate58inter7));
  inv1  gate1325(.a(G290), .O(gate58inter8));
  nand2 gate1326(.a(gate58inter8), .b(gate58inter7), .O(gate58inter9));
  nand2 gate1327(.a(s_111), .b(gate58inter3), .O(gate58inter10));
  nor2  gate1328(.a(gate58inter10), .b(gate58inter9), .O(gate58inter11));
  nor2  gate1329(.a(gate58inter11), .b(gate58inter6), .O(gate58inter12));
  nand2 gate1330(.a(gate58inter12), .b(gate58inter1), .O(G379));

  xor2  gate827(.a(G293), .b(G19), .O(gate59inter0));
  nand2 gate828(.a(gate59inter0), .b(s_40), .O(gate59inter1));
  and2  gate829(.a(G293), .b(G19), .O(gate59inter2));
  inv1  gate830(.a(s_40), .O(gate59inter3));
  inv1  gate831(.a(s_41), .O(gate59inter4));
  nand2 gate832(.a(gate59inter4), .b(gate59inter3), .O(gate59inter5));
  nor2  gate833(.a(gate59inter5), .b(gate59inter2), .O(gate59inter6));
  inv1  gate834(.a(G19), .O(gate59inter7));
  inv1  gate835(.a(G293), .O(gate59inter8));
  nand2 gate836(.a(gate59inter8), .b(gate59inter7), .O(gate59inter9));
  nand2 gate837(.a(s_41), .b(gate59inter3), .O(gate59inter10));
  nor2  gate838(.a(gate59inter10), .b(gate59inter9), .O(gate59inter11));
  nor2  gate839(.a(gate59inter11), .b(gate59inter6), .O(gate59inter12));
  nand2 gate840(.a(gate59inter12), .b(gate59inter1), .O(G380));

  xor2  gate1877(.a(G293), .b(G20), .O(gate60inter0));
  nand2 gate1878(.a(gate60inter0), .b(s_190), .O(gate60inter1));
  and2  gate1879(.a(G293), .b(G20), .O(gate60inter2));
  inv1  gate1880(.a(s_190), .O(gate60inter3));
  inv1  gate1881(.a(s_191), .O(gate60inter4));
  nand2 gate1882(.a(gate60inter4), .b(gate60inter3), .O(gate60inter5));
  nor2  gate1883(.a(gate60inter5), .b(gate60inter2), .O(gate60inter6));
  inv1  gate1884(.a(G20), .O(gate60inter7));
  inv1  gate1885(.a(G293), .O(gate60inter8));
  nand2 gate1886(.a(gate60inter8), .b(gate60inter7), .O(gate60inter9));
  nand2 gate1887(.a(s_191), .b(gate60inter3), .O(gate60inter10));
  nor2  gate1888(.a(gate60inter10), .b(gate60inter9), .O(gate60inter11));
  nor2  gate1889(.a(gate60inter11), .b(gate60inter6), .O(gate60inter12));
  nand2 gate1890(.a(gate60inter12), .b(gate60inter1), .O(G381));
nand2 gate61( .a(G21), .b(G296), .O(G382) );

  xor2  gate673(.a(G296), .b(G22), .O(gate62inter0));
  nand2 gate674(.a(gate62inter0), .b(s_18), .O(gate62inter1));
  and2  gate675(.a(G296), .b(G22), .O(gate62inter2));
  inv1  gate676(.a(s_18), .O(gate62inter3));
  inv1  gate677(.a(s_19), .O(gate62inter4));
  nand2 gate678(.a(gate62inter4), .b(gate62inter3), .O(gate62inter5));
  nor2  gate679(.a(gate62inter5), .b(gate62inter2), .O(gate62inter6));
  inv1  gate680(.a(G22), .O(gate62inter7));
  inv1  gate681(.a(G296), .O(gate62inter8));
  nand2 gate682(.a(gate62inter8), .b(gate62inter7), .O(gate62inter9));
  nand2 gate683(.a(s_19), .b(gate62inter3), .O(gate62inter10));
  nor2  gate684(.a(gate62inter10), .b(gate62inter9), .O(gate62inter11));
  nor2  gate685(.a(gate62inter11), .b(gate62inter6), .O(gate62inter12));
  nand2 gate686(.a(gate62inter12), .b(gate62inter1), .O(G383));

  xor2  gate1387(.a(G299), .b(G23), .O(gate63inter0));
  nand2 gate1388(.a(gate63inter0), .b(s_120), .O(gate63inter1));
  and2  gate1389(.a(G299), .b(G23), .O(gate63inter2));
  inv1  gate1390(.a(s_120), .O(gate63inter3));
  inv1  gate1391(.a(s_121), .O(gate63inter4));
  nand2 gate1392(.a(gate63inter4), .b(gate63inter3), .O(gate63inter5));
  nor2  gate1393(.a(gate63inter5), .b(gate63inter2), .O(gate63inter6));
  inv1  gate1394(.a(G23), .O(gate63inter7));
  inv1  gate1395(.a(G299), .O(gate63inter8));
  nand2 gate1396(.a(gate63inter8), .b(gate63inter7), .O(gate63inter9));
  nand2 gate1397(.a(s_121), .b(gate63inter3), .O(gate63inter10));
  nor2  gate1398(.a(gate63inter10), .b(gate63inter9), .O(gate63inter11));
  nor2  gate1399(.a(gate63inter11), .b(gate63inter6), .O(gate63inter12));
  nand2 gate1400(.a(gate63inter12), .b(gate63inter1), .O(G384));
nand2 gate64( .a(G24), .b(G299), .O(G385) );

  xor2  gate757(.a(G302), .b(G25), .O(gate65inter0));
  nand2 gate758(.a(gate65inter0), .b(s_30), .O(gate65inter1));
  and2  gate759(.a(G302), .b(G25), .O(gate65inter2));
  inv1  gate760(.a(s_30), .O(gate65inter3));
  inv1  gate761(.a(s_31), .O(gate65inter4));
  nand2 gate762(.a(gate65inter4), .b(gate65inter3), .O(gate65inter5));
  nor2  gate763(.a(gate65inter5), .b(gate65inter2), .O(gate65inter6));
  inv1  gate764(.a(G25), .O(gate65inter7));
  inv1  gate765(.a(G302), .O(gate65inter8));
  nand2 gate766(.a(gate65inter8), .b(gate65inter7), .O(gate65inter9));
  nand2 gate767(.a(s_31), .b(gate65inter3), .O(gate65inter10));
  nor2  gate768(.a(gate65inter10), .b(gate65inter9), .O(gate65inter11));
  nor2  gate769(.a(gate65inter11), .b(gate65inter6), .O(gate65inter12));
  nand2 gate770(.a(gate65inter12), .b(gate65inter1), .O(G386));

  xor2  gate1695(.a(G302), .b(G26), .O(gate66inter0));
  nand2 gate1696(.a(gate66inter0), .b(s_164), .O(gate66inter1));
  and2  gate1697(.a(G302), .b(G26), .O(gate66inter2));
  inv1  gate1698(.a(s_164), .O(gate66inter3));
  inv1  gate1699(.a(s_165), .O(gate66inter4));
  nand2 gate1700(.a(gate66inter4), .b(gate66inter3), .O(gate66inter5));
  nor2  gate1701(.a(gate66inter5), .b(gate66inter2), .O(gate66inter6));
  inv1  gate1702(.a(G26), .O(gate66inter7));
  inv1  gate1703(.a(G302), .O(gate66inter8));
  nand2 gate1704(.a(gate66inter8), .b(gate66inter7), .O(gate66inter9));
  nand2 gate1705(.a(s_165), .b(gate66inter3), .O(gate66inter10));
  nor2  gate1706(.a(gate66inter10), .b(gate66inter9), .O(gate66inter11));
  nor2  gate1707(.a(gate66inter11), .b(gate66inter6), .O(gate66inter12));
  nand2 gate1708(.a(gate66inter12), .b(gate66inter1), .O(G387));
nand2 gate67( .a(G27), .b(G305), .O(G388) );
nand2 gate68( .a(G28), .b(G305), .O(G389) );

  xor2  gate2283(.a(G308), .b(G29), .O(gate69inter0));
  nand2 gate2284(.a(gate69inter0), .b(s_248), .O(gate69inter1));
  and2  gate2285(.a(G308), .b(G29), .O(gate69inter2));
  inv1  gate2286(.a(s_248), .O(gate69inter3));
  inv1  gate2287(.a(s_249), .O(gate69inter4));
  nand2 gate2288(.a(gate69inter4), .b(gate69inter3), .O(gate69inter5));
  nor2  gate2289(.a(gate69inter5), .b(gate69inter2), .O(gate69inter6));
  inv1  gate2290(.a(G29), .O(gate69inter7));
  inv1  gate2291(.a(G308), .O(gate69inter8));
  nand2 gate2292(.a(gate69inter8), .b(gate69inter7), .O(gate69inter9));
  nand2 gate2293(.a(s_249), .b(gate69inter3), .O(gate69inter10));
  nor2  gate2294(.a(gate69inter10), .b(gate69inter9), .O(gate69inter11));
  nor2  gate2295(.a(gate69inter11), .b(gate69inter6), .O(gate69inter12));
  nand2 gate2296(.a(gate69inter12), .b(gate69inter1), .O(G390));
nand2 gate70( .a(G30), .b(G308), .O(G391) );

  xor2  gate2311(.a(G311), .b(G31), .O(gate71inter0));
  nand2 gate2312(.a(gate71inter0), .b(s_252), .O(gate71inter1));
  and2  gate2313(.a(G311), .b(G31), .O(gate71inter2));
  inv1  gate2314(.a(s_252), .O(gate71inter3));
  inv1  gate2315(.a(s_253), .O(gate71inter4));
  nand2 gate2316(.a(gate71inter4), .b(gate71inter3), .O(gate71inter5));
  nor2  gate2317(.a(gate71inter5), .b(gate71inter2), .O(gate71inter6));
  inv1  gate2318(.a(G31), .O(gate71inter7));
  inv1  gate2319(.a(G311), .O(gate71inter8));
  nand2 gate2320(.a(gate71inter8), .b(gate71inter7), .O(gate71inter9));
  nand2 gate2321(.a(s_253), .b(gate71inter3), .O(gate71inter10));
  nor2  gate2322(.a(gate71inter10), .b(gate71inter9), .O(gate71inter11));
  nor2  gate2323(.a(gate71inter11), .b(gate71inter6), .O(gate71inter12));
  nand2 gate2324(.a(gate71inter12), .b(gate71inter1), .O(G392));
nand2 gate72( .a(G32), .b(G311), .O(G393) );
nand2 gate73( .a(G1), .b(G314), .O(G394) );

  xor2  gate2087(.a(G314), .b(G5), .O(gate74inter0));
  nand2 gate2088(.a(gate74inter0), .b(s_220), .O(gate74inter1));
  and2  gate2089(.a(G314), .b(G5), .O(gate74inter2));
  inv1  gate2090(.a(s_220), .O(gate74inter3));
  inv1  gate2091(.a(s_221), .O(gate74inter4));
  nand2 gate2092(.a(gate74inter4), .b(gate74inter3), .O(gate74inter5));
  nor2  gate2093(.a(gate74inter5), .b(gate74inter2), .O(gate74inter6));
  inv1  gate2094(.a(G5), .O(gate74inter7));
  inv1  gate2095(.a(G314), .O(gate74inter8));
  nand2 gate2096(.a(gate74inter8), .b(gate74inter7), .O(gate74inter9));
  nand2 gate2097(.a(s_221), .b(gate74inter3), .O(gate74inter10));
  nor2  gate2098(.a(gate74inter10), .b(gate74inter9), .O(gate74inter11));
  nor2  gate2099(.a(gate74inter11), .b(gate74inter6), .O(gate74inter12));
  nand2 gate2100(.a(gate74inter12), .b(gate74inter1), .O(G395));

  xor2  gate1149(.a(G317), .b(G9), .O(gate75inter0));
  nand2 gate1150(.a(gate75inter0), .b(s_86), .O(gate75inter1));
  and2  gate1151(.a(G317), .b(G9), .O(gate75inter2));
  inv1  gate1152(.a(s_86), .O(gate75inter3));
  inv1  gate1153(.a(s_87), .O(gate75inter4));
  nand2 gate1154(.a(gate75inter4), .b(gate75inter3), .O(gate75inter5));
  nor2  gate1155(.a(gate75inter5), .b(gate75inter2), .O(gate75inter6));
  inv1  gate1156(.a(G9), .O(gate75inter7));
  inv1  gate1157(.a(G317), .O(gate75inter8));
  nand2 gate1158(.a(gate75inter8), .b(gate75inter7), .O(gate75inter9));
  nand2 gate1159(.a(s_87), .b(gate75inter3), .O(gate75inter10));
  nor2  gate1160(.a(gate75inter10), .b(gate75inter9), .O(gate75inter11));
  nor2  gate1161(.a(gate75inter11), .b(gate75inter6), .O(gate75inter12));
  nand2 gate1162(.a(gate75inter12), .b(gate75inter1), .O(G396));
nand2 gate76( .a(G13), .b(G317), .O(G397) );
nand2 gate77( .a(G2), .b(G320), .O(G398) );

  xor2  gate2997(.a(G320), .b(G6), .O(gate78inter0));
  nand2 gate2998(.a(gate78inter0), .b(s_350), .O(gate78inter1));
  and2  gate2999(.a(G320), .b(G6), .O(gate78inter2));
  inv1  gate3000(.a(s_350), .O(gate78inter3));
  inv1  gate3001(.a(s_351), .O(gate78inter4));
  nand2 gate3002(.a(gate78inter4), .b(gate78inter3), .O(gate78inter5));
  nor2  gate3003(.a(gate78inter5), .b(gate78inter2), .O(gate78inter6));
  inv1  gate3004(.a(G6), .O(gate78inter7));
  inv1  gate3005(.a(G320), .O(gate78inter8));
  nand2 gate3006(.a(gate78inter8), .b(gate78inter7), .O(gate78inter9));
  nand2 gate3007(.a(s_351), .b(gate78inter3), .O(gate78inter10));
  nor2  gate3008(.a(gate78inter10), .b(gate78inter9), .O(gate78inter11));
  nor2  gate3009(.a(gate78inter11), .b(gate78inter6), .O(gate78inter12));
  nand2 gate3010(.a(gate78inter12), .b(gate78inter1), .O(G399));
nand2 gate79( .a(G10), .b(G323), .O(G400) );
nand2 gate80( .a(G14), .b(G323), .O(G401) );
nand2 gate81( .a(G3), .b(G326), .O(G402) );
nand2 gate82( .a(G7), .b(G326), .O(G403) );

  xor2  gate1499(.a(G329), .b(G11), .O(gate83inter0));
  nand2 gate1500(.a(gate83inter0), .b(s_136), .O(gate83inter1));
  and2  gate1501(.a(G329), .b(G11), .O(gate83inter2));
  inv1  gate1502(.a(s_136), .O(gate83inter3));
  inv1  gate1503(.a(s_137), .O(gate83inter4));
  nand2 gate1504(.a(gate83inter4), .b(gate83inter3), .O(gate83inter5));
  nor2  gate1505(.a(gate83inter5), .b(gate83inter2), .O(gate83inter6));
  inv1  gate1506(.a(G11), .O(gate83inter7));
  inv1  gate1507(.a(G329), .O(gate83inter8));
  nand2 gate1508(.a(gate83inter8), .b(gate83inter7), .O(gate83inter9));
  nand2 gate1509(.a(s_137), .b(gate83inter3), .O(gate83inter10));
  nor2  gate1510(.a(gate83inter10), .b(gate83inter9), .O(gate83inter11));
  nor2  gate1511(.a(gate83inter11), .b(gate83inter6), .O(gate83inter12));
  nand2 gate1512(.a(gate83inter12), .b(gate83inter1), .O(G404));

  xor2  gate1205(.a(G329), .b(G15), .O(gate84inter0));
  nand2 gate1206(.a(gate84inter0), .b(s_94), .O(gate84inter1));
  and2  gate1207(.a(G329), .b(G15), .O(gate84inter2));
  inv1  gate1208(.a(s_94), .O(gate84inter3));
  inv1  gate1209(.a(s_95), .O(gate84inter4));
  nand2 gate1210(.a(gate84inter4), .b(gate84inter3), .O(gate84inter5));
  nor2  gate1211(.a(gate84inter5), .b(gate84inter2), .O(gate84inter6));
  inv1  gate1212(.a(G15), .O(gate84inter7));
  inv1  gate1213(.a(G329), .O(gate84inter8));
  nand2 gate1214(.a(gate84inter8), .b(gate84inter7), .O(gate84inter9));
  nand2 gate1215(.a(s_95), .b(gate84inter3), .O(gate84inter10));
  nor2  gate1216(.a(gate84inter10), .b(gate84inter9), .O(gate84inter11));
  nor2  gate1217(.a(gate84inter11), .b(gate84inter6), .O(gate84inter12));
  nand2 gate1218(.a(gate84inter12), .b(gate84inter1), .O(G405));

  xor2  gate785(.a(G332), .b(G4), .O(gate85inter0));
  nand2 gate786(.a(gate85inter0), .b(s_34), .O(gate85inter1));
  and2  gate787(.a(G332), .b(G4), .O(gate85inter2));
  inv1  gate788(.a(s_34), .O(gate85inter3));
  inv1  gate789(.a(s_35), .O(gate85inter4));
  nand2 gate790(.a(gate85inter4), .b(gate85inter3), .O(gate85inter5));
  nor2  gate791(.a(gate85inter5), .b(gate85inter2), .O(gate85inter6));
  inv1  gate792(.a(G4), .O(gate85inter7));
  inv1  gate793(.a(G332), .O(gate85inter8));
  nand2 gate794(.a(gate85inter8), .b(gate85inter7), .O(gate85inter9));
  nand2 gate795(.a(s_35), .b(gate85inter3), .O(gate85inter10));
  nor2  gate796(.a(gate85inter10), .b(gate85inter9), .O(gate85inter11));
  nor2  gate797(.a(gate85inter11), .b(gate85inter6), .O(gate85inter12));
  nand2 gate798(.a(gate85inter12), .b(gate85inter1), .O(G406));
nand2 gate86( .a(G8), .b(G332), .O(G407) );
nand2 gate87( .a(G12), .b(G335), .O(G408) );

  xor2  gate2563(.a(G335), .b(G16), .O(gate88inter0));
  nand2 gate2564(.a(gate88inter0), .b(s_288), .O(gate88inter1));
  and2  gate2565(.a(G335), .b(G16), .O(gate88inter2));
  inv1  gate2566(.a(s_288), .O(gate88inter3));
  inv1  gate2567(.a(s_289), .O(gate88inter4));
  nand2 gate2568(.a(gate88inter4), .b(gate88inter3), .O(gate88inter5));
  nor2  gate2569(.a(gate88inter5), .b(gate88inter2), .O(gate88inter6));
  inv1  gate2570(.a(G16), .O(gate88inter7));
  inv1  gate2571(.a(G335), .O(gate88inter8));
  nand2 gate2572(.a(gate88inter8), .b(gate88inter7), .O(gate88inter9));
  nand2 gate2573(.a(s_289), .b(gate88inter3), .O(gate88inter10));
  nor2  gate2574(.a(gate88inter10), .b(gate88inter9), .O(gate88inter11));
  nor2  gate2575(.a(gate88inter11), .b(gate88inter6), .O(gate88inter12));
  nand2 gate2576(.a(gate88inter12), .b(gate88inter1), .O(G409));
nand2 gate89( .a(G17), .b(G338), .O(G410) );
nand2 gate90( .a(G21), .b(G338), .O(G411) );
nand2 gate91( .a(G25), .b(G341), .O(G412) );
nand2 gate92( .a(G29), .b(G341), .O(G413) );

  xor2  gate2521(.a(G344), .b(G18), .O(gate93inter0));
  nand2 gate2522(.a(gate93inter0), .b(s_282), .O(gate93inter1));
  and2  gate2523(.a(G344), .b(G18), .O(gate93inter2));
  inv1  gate2524(.a(s_282), .O(gate93inter3));
  inv1  gate2525(.a(s_283), .O(gate93inter4));
  nand2 gate2526(.a(gate93inter4), .b(gate93inter3), .O(gate93inter5));
  nor2  gate2527(.a(gate93inter5), .b(gate93inter2), .O(gate93inter6));
  inv1  gate2528(.a(G18), .O(gate93inter7));
  inv1  gate2529(.a(G344), .O(gate93inter8));
  nand2 gate2530(.a(gate93inter8), .b(gate93inter7), .O(gate93inter9));
  nand2 gate2531(.a(s_283), .b(gate93inter3), .O(gate93inter10));
  nor2  gate2532(.a(gate93inter10), .b(gate93inter9), .O(gate93inter11));
  nor2  gate2533(.a(gate93inter11), .b(gate93inter6), .O(gate93inter12));
  nand2 gate2534(.a(gate93inter12), .b(gate93inter1), .O(G414));
nand2 gate94( .a(G22), .b(G344), .O(G415) );
nand2 gate95( .a(G26), .b(G347), .O(G416) );

  xor2  gate1177(.a(G347), .b(G30), .O(gate96inter0));
  nand2 gate1178(.a(gate96inter0), .b(s_90), .O(gate96inter1));
  and2  gate1179(.a(G347), .b(G30), .O(gate96inter2));
  inv1  gate1180(.a(s_90), .O(gate96inter3));
  inv1  gate1181(.a(s_91), .O(gate96inter4));
  nand2 gate1182(.a(gate96inter4), .b(gate96inter3), .O(gate96inter5));
  nor2  gate1183(.a(gate96inter5), .b(gate96inter2), .O(gate96inter6));
  inv1  gate1184(.a(G30), .O(gate96inter7));
  inv1  gate1185(.a(G347), .O(gate96inter8));
  nand2 gate1186(.a(gate96inter8), .b(gate96inter7), .O(gate96inter9));
  nand2 gate1187(.a(s_91), .b(gate96inter3), .O(gate96inter10));
  nor2  gate1188(.a(gate96inter10), .b(gate96inter9), .O(gate96inter11));
  nor2  gate1189(.a(gate96inter11), .b(gate96inter6), .O(gate96inter12));
  nand2 gate1190(.a(gate96inter12), .b(gate96inter1), .O(G417));
nand2 gate97( .a(G19), .b(G350), .O(G418) );

  xor2  gate2633(.a(G350), .b(G23), .O(gate98inter0));
  nand2 gate2634(.a(gate98inter0), .b(s_298), .O(gate98inter1));
  and2  gate2635(.a(G350), .b(G23), .O(gate98inter2));
  inv1  gate2636(.a(s_298), .O(gate98inter3));
  inv1  gate2637(.a(s_299), .O(gate98inter4));
  nand2 gate2638(.a(gate98inter4), .b(gate98inter3), .O(gate98inter5));
  nor2  gate2639(.a(gate98inter5), .b(gate98inter2), .O(gate98inter6));
  inv1  gate2640(.a(G23), .O(gate98inter7));
  inv1  gate2641(.a(G350), .O(gate98inter8));
  nand2 gate2642(.a(gate98inter8), .b(gate98inter7), .O(gate98inter9));
  nand2 gate2643(.a(s_299), .b(gate98inter3), .O(gate98inter10));
  nor2  gate2644(.a(gate98inter10), .b(gate98inter9), .O(gate98inter11));
  nor2  gate2645(.a(gate98inter11), .b(gate98inter6), .O(gate98inter12));
  nand2 gate2646(.a(gate98inter12), .b(gate98inter1), .O(G419));

  xor2  gate1079(.a(G353), .b(G27), .O(gate99inter0));
  nand2 gate1080(.a(gate99inter0), .b(s_76), .O(gate99inter1));
  and2  gate1081(.a(G353), .b(G27), .O(gate99inter2));
  inv1  gate1082(.a(s_76), .O(gate99inter3));
  inv1  gate1083(.a(s_77), .O(gate99inter4));
  nand2 gate1084(.a(gate99inter4), .b(gate99inter3), .O(gate99inter5));
  nor2  gate1085(.a(gate99inter5), .b(gate99inter2), .O(gate99inter6));
  inv1  gate1086(.a(G27), .O(gate99inter7));
  inv1  gate1087(.a(G353), .O(gate99inter8));
  nand2 gate1088(.a(gate99inter8), .b(gate99inter7), .O(gate99inter9));
  nand2 gate1089(.a(s_77), .b(gate99inter3), .O(gate99inter10));
  nor2  gate1090(.a(gate99inter10), .b(gate99inter9), .O(gate99inter11));
  nor2  gate1091(.a(gate99inter11), .b(gate99inter6), .O(gate99inter12));
  nand2 gate1092(.a(gate99inter12), .b(gate99inter1), .O(G420));
nand2 gate100( .a(G31), .b(G353), .O(G421) );

  xor2  gate1933(.a(G356), .b(G20), .O(gate101inter0));
  nand2 gate1934(.a(gate101inter0), .b(s_198), .O(gate101inter1));
  and2  gate1935(.a(G356), .b(G20), .O(gate101inter2));
  inv1  gate1936(.a(s_198), .O(gate101inter3));
  inv1  gate1937(.a(s_199), .O(gate101inter4));
  nand2 gate1938(.a(gate101inter4), .b(gate101inter3), .O(gate101inter5));
  nor2  gate1939(.a(gate101inter5), .b(gate101inter2), .O(gate101inter6));
  inv1  gate1940(.a(G20), .O(gate101inter7));
  inv1  gate1941(.a(G356), .O(gate101inter8));
  nand2 gate1942(.a(gate101inter8), .b(gate101inter7), .O(gate101inter9));
  nand2 gate1943(.a(s_199), .b(gate101inter3), .O(gate101inter10));
  nor2  gate1944(.a(gate101inter10), .b(gate101inter9), .O(gate101inter11));
  nor2  gate1945(.a(gate101inter11), .b(gate101inter6), .O(gate101inter12));
  nand2 gate1946(.a(gate101inter12), .b(gate101inter1), .O(G422));

  xor2  gate2269(.a(G356), .b(G24), .O(gate102inter0));
  nand2 gate2270(.a(gate102inter0), .b(s_246), .O(gate102inter1));
  and2  gate2271(.a(G356), .b(G24), .O(gate102inter2));
  inv1  gate2272(.a(s_246), .O(gate102inter3));
  inv1  gate2273(.a(s_247), .O(gate102inter4));
  nand2 gate2274(.a(gate102inter4), .b(gate102inter3), .O(gate102inter5));
  nor2  gate2275(.a(gate102inter5), .b(gate102inter2), .O(gate102inter6));
  inv1  gate2276(.a(G24), .O(gate102inter7));
  inv1  gate2277(.a(G356), .O(gate102inter8));
  nand2 gate2278(.a(gate102inter8), .b(gate102inter7), .O(gate102inter9));
  nand2 gate2279(.a(s_247), .b(gate102inter3), .O(gate102inter10));
  nor2  gate2280(.a(gate102inter10), .b(gate102inter9), .O(gate102inter11));
  nor2  gate2281(.a(gate102inter11), .b(gate102inter6), .O(gate102inter12));
  nand2 gate2282(.a(gate102inter12), .b(gate102inter1), .O(G423));

  xor2  gate1275(.a(G359), .b(G28), .O(gate103inter0));
  nand2 gate1276(.a(gate103inter0), .b(s_104), .O(gate103inter1));
  and2  gate1277(.a(G359), .b(G28), .O(gate103inter2));
  inv1  gate1278(.a(s_104), .O(gate103inter3));
  inv1  gate1279(.a(s_105), .O(gate103inter4));
  nand2 gate1280(.a(gate103inter4), .b(gate103inter3), .O(gate103inter5));
  nor2  gate1281(.a(gate103inter5), .b(gate103inter2), .O(gate103inter6));
  inv1  gate1282(.a(G28), .O(gate103inter7));
  inv1  gate1283(.a(G359), .O(gate103inter8));
  nand2 gate1284(.a(gate103inter8), .b(gate103inter7), .O(gate103inter9));
  nand2 gate1285(.a(s_105), .b(gate103inter3), .O(gate103inter10));
  nor2  gate1286(.a(gate103inter10), .b(gate103inter9), .O(gate103inter11));
  nor2  gate1287(.a(gate103inter11), .b(gate103inter6), .O(gate103inter12));
  nand2 gate1288(.a(gate103inter12), .b(gate103inter1), .O(G424));
nand2 gate104( .a(G32), .b(G359), .O(G425) );

  xor2  gate1037(.a(G363), .b(G362), .O(gate105inter0));
  nand2 gate1038(.a(gate105inter0), .b(s_70), .O(gate105inter1));
  and2  gate1039(.a(G363), .b(G362), .O(gate105inter2));
  inv1  gate1040(.a(s_70), .O(gate105inter3));
  inv1  gate1041(.a(s_71), .O(gate105inter4));
  nand2 gate1042(.a(gate105inter4), .b(gate105inter3), .O(gate105inter5));
  nor2  gate1043(.a(gate105inter5), .b(gate105inter2), .O(gate105inter6));
  inv1  gate1044(.a(G362), .O(gate105inter7));
  inv1  gate1045(.a(G363), .O(gate105inter8));
  nand2 gate1046(.a(gate105inter8), .b(gate105inter7), .O(gate105inter9));
  nand2 gate1047(.a(s_71), .b(gate105inter3), .O(gate105inter10));
  nor2  gate1048(.a(gate105inter10), .b(gate105inter9), .O(gate105inter11));
  nor2  gate1049(.a(gate105inter11), .b(gate105inter6), .O(gate105inter12));
  nand2 gate1050(.a(gate105inter12), .b(gate105inter1), .O(G426));
nand2 gate106( .a(G364), .b(G365), .O(G429) );
nand2 gate107( .a(G366), .b(G367), .O(G432) );
nand2 gate108( .a(G368), .b(G369), .O(G435) );

  xor2  gate659(.a(G371), .b(G370), .O(gate109inter0));
  nand2 gate660(.a(gate109inter0), .b(s_16), .O(gate109inter1));
  and2  gate661(.a(G371), .b(G370), .O(gate109inter2));
  inv1  gate662(.a(s_16), .O(gate109inter3));
  inv1  gate663(.a(s_17), .O(gate109inter4));
  nand2 gate664(.a(gate109inter4), .b(gate109inter3), .O(gate109inter5));
  nor2  gate665(.a(gate109inter5), .b(gate109inter2), .O(gate109inter6));
  inv1  gate666(.a(G370), .O(gate109inter7));
  inv1  gate667(.a(G371), .O(gate109inter8));
  nand2 gate668(.a(gate109inter8), .b(gate109inter7), .O(gate109inter9));
  nand2 gate669(.a(s_17), .b(gate109inter3), .O(gate109inter10));
  nor2  gate670(.a(gate109inter10), .b(gate109inter9), .O(gate109inter11));
  nor2  gate671(.a(gate109inter11), .b(gate109inter6), .O(gate109inter12));
  nand2 gate672(.a(gate109inter12), .b(gate109inter1), .O(G438));

  xor2  gate1135(.a(G373), .b(G372), .O(gate110inter0));
  nand2 gate1136(.a(gate110inter0), .b(s_84), .O(gate110inter1));
  and2  gate1137(.a(G373), .b(G372), .O(gate110inter2));
  inv1  gate1138(.a(s_84), .O(gate110inter3));
  inv1  gate1139(.a(s_85), .O(gate110inter4));
  nand2 gate1140(.a(gate110inter4), .b(gate110inter3), .O(gate110inter5));
  nor2  gate1141(.a(gate110inter5), .b(gate110inter2), .O(gate110inter6));
  inv1  gate1142(.a(G372), .O(gate110inter7));
  inv1  gate1143(.a(G373), .O(gate110inter8));
  nand2 gate1144(.a(gate110inter8), .b(gate110inter7), .O(gate110inter9));
  nand2 gate1145(.a(s_85), .b(gate110inter3), .O(gate110inter10));
  nor2  gate1146(.a(gate110inter10), .b(gate110inter9), .O(gate110inter11));
  nor2  gate1147(.a(gate110inter11), .b(gate110inter6), .O(gate110inter12));
  nand2 gate1148(.a(gate110inter12), .b(gate110inter1), .O(G441));
nand2 gate111( .a(G374), .b(G375), .O(G444) );

  xor2  gate2955(.a(G377), .b(G376), .O(gate112inter0));
  nand2 gate2956(.a(gate112inter0), .b(s_344), .O(gate112inter1));
  and2  gate2957(.a(G377), .b(G376), .O(gate112inter2));
  inv1  gate2958(.a(s_344), .O(gate112inter3));
  inv1  gate2959(.a(s_345), .O(gate112inter4));
  nand2 gate2960(.a(gate112inter4), .b(gate112inter3), .O(gate112inter5));
  nor2  gate2961(.a(gate112inter5), .b(gate112inter2), .O(gate112inter6));
  inv1  gate2962(.a(G376), .O(gate112inter7));
  inv1  gate2963(.a(G377), .O(gate112inter8));
  nand2 gate2964(.a(gate112inter8), .b(gate112inter7), .O(gate112inter9));
  nand2 gate2965(.a(s_345), .b(gate112inter3), .O(gate112inter10));
  nor2  gate2966(.a(gate112inter10), .b(gate112inter9), .O(gate112inter11));
  nor2  gate2967(.a(gate112inter11), .b(gate112inter6), .O(gate112inter12));
  nand2 gate2968(.a(gate112inter12), .b(gate112inter1), .O(G447));
nand2 gate113( .a(G378), .b(G379), .O(G450) );
nand2 gate114( .a(G380), .b(G381), .O(G453) );
nand2 gate115( .a(G382), .b(G383), .O(G456) );
nand2 gate116( .a(G384), .b(G385), .O(G459) );

  xor2  gate2759(.a(G387), .b(G386), .O(gate117inter0));
  nand2 gate2760(.a(gate117inter0), .b(s_316), .O(gate117inter1));
  and2  gate2761(.a(G387), .b(G386), .O(gate117inter2));
  inv1  gate2762(.a(s_316), .O(gate117inter3));
  inv1  gate2763(.a(s_317), .O(gate117inter4));
  nand2 gate2764(.a(gate117inter4), .b(gate117inter3), .O(gate117inter5));
  nor2  gate2765(.a(gate117inter5), .b(gate117inter2), .O(gate117inter6));
  inv1  gate2766(.a(G386), .O(gate117inter7));
  inv1  gate2767(.a(G387), .O(gate117inter8));
  nand2 gate2768(.a(gate117inter8), .b(gate117inter7), .O(gate117inter9));
  nand2 gate2769(.a(s_317), .b(gate117inter3), .O(gate117inter10));
  nor2  gate2770(.a(gate117inter10), .b(gate117inter9), .O(gate117inter11));
  nor2  gate2771(.a(gate117inter11), .b(gate117inter6), .O(gate117inter12));
  nand2 gate2772(.a(gate117inter12), .b(gate117inter1), .O(G462));

  xor2  gate1681(.a(G389), .b(G388), .O(gate118inter0));
  nand2 gate1682(.a(gate118inter0), .b(s_162), .O(gate118inter1));
  and2  gate1683(.a(G389), .b(G388), .O(gate118inter2));
  inv1  gate1684(.a(s_162), .O(gate118inter3));
  inv1  gate1685(.a(s_163), .O(gate118inter4));
  nand2 gate1686(.a(gate118inter4), .b(gate118inter3), .O(gate118inter5));
  nor2  gate1687(.a(gate118inter5), .b(gate118inter2), .O(gate118inter6));
  inv1  gate1688(.a(G388), .O(gate118inter7));
  inv1  gate1689(.a(G389), .O(gate118inter8));
  nand2 gate1690(.a(gate118inter8), .b(gate118inter7), .O(gate118inter9));
  nand2 gate1691(.a(s_163), .b(gate118inter3), .O(gate118inter10));
  nor2  gate1692(.a(gate118inter10), .b(gate118inter9), .O(gate118inter11));
  nor2  gate1693(.a(gate118inter11), .b(gate118inter6), .O(gate118inter12));
  nand2 gate1694(.a(gate118inter12), .b(gate118inter1), .O(G465));
nand2 gate119( .a(G390), .b(G391), .O(G468) );
nand2 gate120( .a(G392), .b(G393), .O(G471) );
nand2 gate121( .a(G394), .b(G395), .O(G474) );

  xor2  gate1485(.a(G397), .b(G396), .O(gate122inter0));
  nand2 gate1486(.a(gate122inter0), .b(s_134), .O(gate122inter1));
  and2  gate1487(.a(G397), .b(G396), .O(gate122inter2));
  inv1  gate1488(.a(s_134), .O(gate122inter3));
  inv1  gate1489(.a(s_135), .O(gate122inter4));
  nand2 gate1490(.a(gate122inter4), .b(gate122inter3), .O(gate122inter5));
  nor2  gate1491(.a(gate122inter5), .b(gate122inter2), .O(gate122inter6));
  inv1  gate1492(.a(G396), .O(gate122inter7));
  inv1  gate1493(.a(G397), .O(gate122inter8));
  nand2 gate1494(.a(gate122inter8), .b(gate122inter7), .O(gate122inter9));
  nand2 gate1495(.a(s_135), .b(gate122inter3), .O(gate122inter10));
  nor2  gate1496(.a(gate122inter10), .b(gate122inter9), .O(gate122inter11));
  nor2  gate1497(.a(gate122inter11), .b(gate122inter6), .O(gate122inter12));
  nand2 gate1498(.a(gate122inter12), .b(gate122inter1), .O(G477));
nand2 gate123( .a(G398), .b(G399), .O(G480) );
nand2 gate124( .a(G400), .b(G401), .O(G483) );
nand2 gate125( .a(G402), .b(G403), .O(G486) );

  xor2  gate2171(.a(G405), .b(G404), .O(gate126inter0));
  nand2 gate2172(.a(gate126inter0), .b(s_232), .O(gate126inter1));
  and2  gate2173(.a(G405), .b(G404), .O(gate126inter2));
  inv1  gate2174(.a(s_232), .O(gate126inter3));
  inv1  gate2175(.a(s_233), .O(gate126inter4));
  nand2 gate2176(.a(gate126inter4), .b(gate126inter3), .O(gate126inter5));
  nor2  gate2177(.a(gate126inter5), .b(gate126inter2), .O(gate126inter6));
  inv1  gate2178(.a(G404), .O(gate126inter7));
  inv1  gate2179(.a(G405), .O(gate126inter8));
  nand2 gate2180(.a(gate126inter8), .b(gate126inter7), .O(gate126inter9));
  nand2 gate2181(.a(s_233), .b(gate126inter3), .O(gate126inter10));
  nor2  gate2182(.a(gate126inter10), .b(gate126inter9), .O(gate126inter11));
  nor2  gate2183(.a(gate126inter11), .b(gate126inter6), .O(gate126inter12));
  nand2 gate2184(.a(gate126inter12), .b(gate126inter1), .O(G489));
nand2 gate127( .a(G406), .b(G407), .O(G492) );

  xor2  gate1009(.a(G409), .b(G408), .O(gate128inter0));
  nand2 gate1010(.a(gate128inter0), .b(s_66), .O(gate128inter1));
  and2  gate1011(.a(G409), .b(G408), .O(gate128inter2));
  inv1  gate1012(.a(s_66), .O(gate128inter3));
  inv1  gate1013(.a(s_67), .O(gate128inter4));
  nand2 gate1014(.a(gate128inter4), .b(gate128inter3), .O(gate128inter5));
  nor2  gate1015(.a(gate128inter5), .b(gate128inter2), .O(gate128inter6));
  inv1  gate1016(.a(G408), .O(gate128inter7));
  inv1  gate1017(.a(G409), .O(gate128inter8));
  nand2 gate1018(.a(gate128inter8), .b(gate128inter7), .O(gate128inter9));
  nand2 gate1019(.a(s_67), .b(gate128inter3), .O(gate128inter10));
  nor2  gate1020(.a(gate128inter10), .b(gate128inter9), .O(gate128inter11));
  nor2  gate1021(.a(gate128inter11), .b(gate128inter6), .O(gate128inter12));
  nand2 gate1022(.a(gate128inter12), .b(gate128inter1), .O(G495));

  xor2  gate2045(.a(G411), .b(G410), .O(gate129inter0));
  nand2 gate2046(.a(gate129inter0), .b(s_214), .O(gate129inter1));
  and2  gate2047(.a(G411), .b(G410), .O(gate129inter2));
  inv1  gate2048(.a(s_214), .O(gate129inter3));
  inv1  gate2049(.a(s_215), .O(gate129inter4));
  nand2 gate2050(.a(gate129inter4), .b(gate129inter3), .O(gate129inter5));
  nor2  gate2051(.a(gate129inter5), .b(gate129inter2), .O(gate129inter6));
  inv1  gate2052(.a(G410), .O(gate129inter7));
  inv1  gate2053(.a(G411), .O(gate129inter8));
  nand2 gate2054(.a(gate129inter8), .b(gate129inter7), .O(gate129inter9));
  nand2 gate2055(.a(s_215), .b(gate129inter3), .O(gate129inter10));
  nor2  gate2056(.a(gate129inter10), .b(gate129inter9), .O(gate129inter11));
  nor2  gate2057(.a(gate129inter11), .b(gate129inter6), .O(gate129inter12));
  nand2 gate2058(.a(gate129inter12), .b(gate129inter1), .O(G498));
nand2 gate130( .a(G412), .b(G413), .O(G501) );

  xor2  gate2899(.a(G415), .b(G414), .O(gate131inter0));
  nand2 gate2900(.a(gate131inter0), .b(s_336), .O(gate131inter1));
  and2  gate2901(.a(G415), .b(G414), .O(gate131inter2));
  inv1  gate2902(.a(s_336), .O(gate131inter3));
  inv1  gate2903(.a(s_337), .O(gate131inter4));
  nand2 gate2904(.a(gate131inter4), .b(gate131inter3), .O(gate131inter5));
  nor2  gate2905(.a(gate131inter5), .b(gate131inter2), .O(gate131inter6));
  inv1  gate2906(.a(G414), .O(gate131inter7));
  inv1  gate2907(.a(G415), .O(gate131inter8));
  nand2 gate2908(.a(gate131inter8), .b(gate131inter7), .O(gate131inter9));
  nand2 gate2909(.a(s_337), .b(gate131inter3), .O(gate131inter10));
  nor2  gate2910(.a(gate131inter10), .b(gate131inter9), .O(gate131inter11));
  nor2  gate2911(.a(gate131inter11), .b(gate131inter6), .O(gate131inter12));
  nand2 gate2912(.a(gate131inter12), .b(gate131inter1), .O(G504));

  xor2  gate1597(.a(G417), .b(G416), .O(gate132inter0));
  nand2 gate1598(.a(gate132inter0), .b(s_150), .O(gate132inter1));
  and2  gate1599(.a(G417), .b(G416), .O(gate132inter2));
  inv1  gate1600(.a(s_150), .O(gate132inter3));
  inv1  gate1601(.a(s_151), .O(gate132inter4));
  nand2 gate1602(.a(gate132inter4), .b(gate132inter3), .O(gate132inter5));
  nor2  gate1603(.a(gate132inter5), .b(gate132inter2), .O(gate132inter6));
  inv1  gate1604(.a(G416), .O(gate132inter7));
  inv1  gate1605(.a(G417), .O(gate132inter8));
  nand2 gate1606(.a(gate132inter8), .b(gate132inter7), .O(gate132inter9));
  nand2 gate1607(.a(s_151), .b(gate132inter3), .O(gate132inter10));
  nor2  gate1608(.a(gate132inter10), .b(gate132inter9), .O(gate132inter11));
  nor2  gate1609(.a(gate132inter11), .b(gate132inter6), .O(gate132inter12));
  nand2 gate1610(.a(gate132inter12), .b(gate132inter1), .O(G507));
nand2 gate133( .a(G418), .b(G419), .O(G510) );
nand2 gate134( .a(G420), .b(G421), .O(G513) );

  xor2  gate1527(.a(G423), .b(G422), .O(gate135inter0));
  nand2 gate1528(.a(gate135inter0), .b(s_140), .O(gate135inter1));
  and2  gate1529(.a(G423), .b(G422), .O(gate135inter2));
  inv1  gate1530(.a(s_140), .O(gate135inter3));
  inv1  gate1531(.a(s_141), .O(gate135inter4));
  nand2 gate1532(.a(gate135inter4), .b(gate135inter3), .O(gate135inter5));
  nor2  gate1533(.a(gate135inter5), .b(gate135inter2), .O(gate135inter6));
  inv1  gate1534(.a(G422), .O(gate135inter7));
  inv1  gate1535(.a(G423), .O(gate135inter8));
  nand2 gate1536(.a(gate135inter8), .b(gate135inter7), .O(gate135inter9));
  nand2 gate1537(.a(s_141), .b(gate135inter3), .O(gate135inter10));
  nor2  gate1538(.a(gate135inter10), .b(gate135inter9), .O(gate135inter11));
  nor2  gate1539(.a(gate135inter11), .b(gate135inter6), .O(gate135inter12));
  nand2 gate1540(.a(gate135inter12), .b(gate135inter1), .O(G516));

  xor2  gate1289(.a(G425), .b(G424), .O(gate136inter0));
  nand2 gate1290(.a(gate136inter0), .b(s_106), .O(gate136inter1));
  and2  gate1291(.a(G425), .b(G424), .O(gate136inter2));
  inv1  gate1292(.a(s_106), .O(gate136inter3));
  inv1  gate1293(.a(s_107), .O(gate136inter4));
  nand2 gate1294(.a(gate136inter4), .b(gate136inter3), .O(gate136inter5));
  nor2  gate1295(.a(gate136inter5), .b(gate136inter2), .O(gate136inter6));
  inv1  gate1296(.a(G424), .O(gate136inter7));
  inv1  gate1297(.a(G425), .O(gate136inter8));
  nand2 gate1298(.a(gate136inter8), .b(gate136inter7), .O(gate136inter9));
  nand2 gate1299(.a(s_107), .b(gate136inter3), .O(gate136inter10));
  nor2  gate1300(.a(gate136inter10), .b(gate136inter9), .O(gate136inter11));
  nor2  gate1301(.a(gate136inter11), .b(gate136inter6), .O(gate136inter12));
  nand2 gate1302(.a(gate136inter12), .b(gate136inter1), .O(G519));
nand2 gate137( .a(G426), .b(G429), .O(G522) );

  xor2  gate2773(.a(G435), .b(G432), .O(gate138inter0));
  nand2 gate2774(.a(gate138inter0), .b(s_318), .O(gate138inter1));
  and2  gate2775(.a(G435), .b(G432), .O(gate138inter2));
  inv1  gate2776(.a(s_318), .O(gate138inter3));
  inv1  gate2777(.a(s_319), .O(gate138inter4));
  nand2 gate2778(.a(gate138inter4), .b(gate138inter3), .O(gate138inter5));
  nor2  gate2779(.a(gate138inter5), .b(gate138inter2), .O(gate138inter6));
  inv1  gate2780(.a(G432), .O(gate138inter7));
  inv1  gate2781(.a(G435), .O(gate138inter8));
  nand2 gate2782(.a(gate138inter8), .b(gate138inter7), .O(gate138inter9));
  nand2 gate2783(.a(s_319), .b(gate138inter3), .O(gate138inter10));
  nor2  gate2784(.a(gate138inter10), .b(gate138inter9), .O(gate138inter11));
  nor2  gate2785(.a(gate138inter11), .b(gate138inter6), .O(gate138inter12));
  nand2 gate2786(.a(gate138inter12), .b(gate138inter1), .O(G525));

  xor2  gate1373(.a(G441), .b(G438), .O(gate139inter0));
  nand2 gate1374(.a(gate139inter0), .b(s_118), .O(gate139inter1));
  and2  gate1375(.a(G441), .b(G438), .O(gate139inter2));
  inv1  gate1376(.a(s_118), .O(gate139inter3));
  inv1  gate1377(.a(s_119), .O(gate139inter4));
  nand2 gate1378(.a(gate139inter4), .b(gate139inter3), .O(gate139inter5));
  nor2  gate1379(.a(gate139inter5), .b(gate139inter2), .O(gate139inter6));
  inv1  gate1380(.a(G438), .O(gate139inter7));
  inv1  gate1381(.a(G441), .O(gate139inter8));
  nand2 gate1382(.a(gate139inter8), .b(gate139inter7), .O(gate139inter9));
  nand2 gate1383(.a(s_119), .b(gate139inter3), .O(gate139inter10));
  nor2  gate1384(.a(gate139inter10), .b(gate139inter9), .O(gate139inter11));
  nor2  gate1385(.a(gate139inter11), .b(gate139inter6), .O(gate139inter12));
  nand2 gate1386(.a(gate139inter12), .b(gate139inter1), .O(G528));
nand2 gate140( .a(G444), .b(G447), .O(G531) );

  xor2  gate2227(.a(G453), .b(G450), .O(gate141inter0));
  nand2 gate2228(.a(gate141inter0), .b(s_240), .O(gate141inter1));
  and2  gate2229(.a(G453), .b(G450), .O(gate141inter2));
  inv1  gate2230(.a(s_240), .O(gate141inter3));
  inv1  gate2231(.a(s_241), .O(gate141inter4));
  nand2 gate2232(.a(gate141inter4), .b(gate141inter3), .O(gate141inter5));
  nor2  gate2233(.a(gate141inter5), .b(gate141inter2), .O(gate141inter6));
  inv1  gate2234(.a(G450), .O(gate141inter7));
  inv1  gate2235(.a(G453), .O(gate141inter8));
  nand2 gate2236(.a(gate141inter8), .b(gate141inter7), .O(gate141inter9));
  nand2 gate2237(.a(s_241), .b(gate141inter3), .O(gate141inter10));
  nor2  gate2238(.a(gate141inter10), .b(gate141inter9), .O(gate141inter11));
  nor2  gate2239(.a(gate141inter11), .b(gate141inter6), .O(gate141inter12));
  nand2 gate2240(.a(gate141inter12), .b(gate141inter1), .O(G534));
nand2 gate142( .a(G456), .b(G459), .O(G537) );
nand2 gate143( .a(G462), .b(G465), .O(G540) );

  xor2  gate2129(.a(G471), .b(G468), .O(gate144inter0));
  nand2 gate2130(.a(gate144inter0), .b(s_226), .O(gate144inter1));
  and2  gate2131(.a(G471), .b(G468), .O(gate144inter2));
  inv1  gate2132(.a(s_226), .O(gate144inter3));
  inv1  gate2133(.a(s_227), .O(gate144inter4));
  nand2 gate2134(.a(gate144inter4), .b(gate144inter3), .O(gate144inter5));
  nor2  gate2135(.a(gate144inter5), .b(gate144inter2), .O(gate144inter6));
  inv1  gate2136(.a(G468), .O(gate144inter7));
  inv1  gate2137(.a(G471), .O(gate144inter8));
  nand2 gate2138(.a(gate144inter8), .b(gate144inter7), .O(gate144inter9));
  nand2 gate2139(.a(s_227), .b(gate144inter3), .O(gate144inter10));
  nor2  gate2140(.a(gate144inter10), .b(gate144inter9), .O(gate144inter11));
  nor2  gate2141(.a(gate144inter11), .b(gate144inter6), .O(gate144inter12));
  nand2 gate2142(.a(gate144inter12), .b(gate144inter1), .O(G543));

  xor2  gate1065(.a(G477), .b(G474), .O(gate145inter0));
  nand2 gate1066(.a(gate145inter0), .b(s_74), .O(gate145inter1));
  and2  gate1067(.a(G477), .b(G474), .O(gate145inter2));
  inv1  gate1068(.a(s_74), .O(gate145inter3));
  inv1  gate1069(.a(s_75), .O(gate145inter4));
  nand2 gate1070(.a(gate145inter4), .b(gate145inter3), .O(gate145inter5));
  nor2  gate1071(.a(gate145inter5), .b(gate145inter2), .O(gate145inter6));
  inv1  gate1072(.a(G474), .O(gate145inter7));
  inv1  gate1073(.a(G477), .O(gate145inter8));
  nand2 gate1074(.a(gate145inter8), .b(gate145inter7), .O(gate145inter9));
  nand2 gate1075(.a(s_75), .b(gate145inter3), .O(gate145inter10));
  nor2  gate1076(.a(gate145inter10), .b(gate145inter9), .O(gate145inter11));
  nor2  gate1077(.a(gate145inter11), .b(gate145inter6), .O(gate145inter12));
  nand2 gate1078(.a(gate145inter12), .b(gate145inter1), .O(G546));

  xor2  gate1163(.a(G483), .b(G480), .O(gate146inter0));
  nand2 gate1164(.a(gate146inter0), .b(s_88), .O(gate146inter1));
  and2  gate1165(.a(G483), .b(G480), .O(gate146inter2));
  inv1  gate1166(.a(s_88), .O(gate146inter3));
  inv1  gate1167(.a(s_89), .O(gate146inter4));
  nand2 gate1168(.a(gate146inter4), .b(gate146inter3), .O(gate146inter5));
  nor2  gate1169(.a(gate146inter5), .b(gate146inter2), .O(gate146inter6));
  inv1  gate1170(.a(G480), .O(gate146inter7));
  inv1  gate1171(.a(G483), .O(gate146inter8));
  nand2 gate1172(.a(gate146inter8), .b(gate146inter7), .O(gate146inter9));
  nand2 gate1173(.a(s_89), .b(gate146inter3), .O(gate146inter10));
  nor2  gate1174(.a(gate146inter10), .b(gate146inter9), .O(gate146inter11));
  nor2  gate1175(.a(gate146inter11), .b(gate146inter6), .O(gate146inter12));
  nand2 gate1176(.a(gate146inter12), .b(gate146inter1), .O(G549));

  xor2  gate2031(.a(G489), .b(G486), .O(gate147inter0));
  nand2 gate2032(.a(gate147inter0), .b(s_212), .O(gate147inter1));
  and2  gate2033(.a(G489), .b(G486), .O(gate147inter2));
  inv1  gate2034(.a(s_212), .O(gate147inter3));
  inv1  gate2035(.a(s_213), .O(gate147inter4));
  nand2 gate2036(.a(gate147inter4), .b(gate147inter3), .O(gate147inter5));
  nor2  gate2037(.a(gate147inter5), .b(gate147inter2), .O(gate147inter6));
  inv1  gate2038(.a(G486), .O(gate147inter7));
  inv1  gate2039(.a(G489), .O(gate147inter8));
  nand2 gate2040(.a(gate147inter8), .b(gate147inter7), .O(gate147inter9));
  nand2 gate2041(.a(s_213), .b(gate147inter3), .O(gate147inter10));
  nor2  gate2042(.a(gate147inter10), .b(gate147inter9), .O(gate147inter11));
  nor2  gate2043(.a(gate147inter11), .b(gate147inter6), .O(gate147inter12));
  nand2 gate2044(.a(gate147inter12), .b(gate147inter1), .O(G552));
nand2 gate148( .a(G492), .b(G495), .O(G555) );
nand2 gate149( .a(G498), .b(G501), .O(G558) );
nand2 gate150( .a(G504), .b(G507), .O(G561) );
nand2 gate151( .a(G510), .b(G513), .O(G564) );

  xor2  gate2717(.a(G519), .b(G516), .O(gate152inter0));
  nand2 gate2718(.a(gate152inter0), .b(s_310), .O(gate152inter1));
  and2  gate2719(.a(G519), .b(G516), .O(gate152inter2));
  inv1  gate2720(.a(s_310), .O(gate152inter3));
  inv1  gate2721(.a(s_311), .O(gate152inter4));
  nand2 gate2722(.a(gate152inter4), .b(gate152inter3), .O(gate152inter5));
  nor2  gate2723(.a(gate152inter5), .b(gate152inter2), .O(gate152inter6));
  inv1  gate2724(.a(G516), .O(gate152inter7));
  inv1  gate2725(.a(G519), .O(gate152inter8));
  nand2 gate2726(.a(gate152inter8), .b(gate152inter7), .O(gate152inter9));
  nand2 gate2727(.a(s_311), .b(gate152inter3), .O(gate152inter10));
  nor2  gate2728(.a(gate152inter10), .b(gate152inter9), .O(gate152inter11));
  nor2  gate2729(.a(gate152inter11), .b(gate152inter6), .O(gate152inter12));
  nand2 gate2730(.a(gate152inter12), .b(gate152inter1), .O(G567));

  xor2  gate855(.a(G522), .b(G426), .O(gate153inter0));
  nand2 gate856(.a(gate153inter0), .b(s_44), .O(gate153inter1));
  and2  gate857(.a(G522), .b(G426), .O(gate153inter2));
  inv1  gate858(.a(s_44), .O(gate153inter3));
  inv1  gate859(.a(s_45), .O(gate153inter4));
  nand2 gate860(.a(gate153inter4), .b(gate153inter3), .O(gate153inter5));
  nor2  gate861(.a(gate153inter5), .b(gate153inter2), .O(gate153inter6));
  inv1  gate862(.a(G426), .O(gate153inter7));
  inv1  gate863(.a(G522), .O(gate153inter8));
  nand2 gate864(.a(gate153inter8), .b(gate153inter7), .O(gate153inter9));
  nand2 gate865(.a(s_45), .b(gate153inter3), .O(gate153inter10));
  nor2  gate866(.a(gate153inter10), .b(gate153inter9), .O(gate153inter11));
  nor2  gate867(.a(gate153inter11), .b(gate153inter6), .O(gate153inter12));
  nand2 gate868(.a(gate153inter12), .b(gate153inter1), .O(G570));

  xor2  gate2703(.a(G522), .b(G429), .O(gate154inter0));
  nand2 gate2704(.a(gate154inter0), .b(s_308), .O(gate154inter1));
  and2  gate2705(.a(G522), .b(G429), .O(gate154inter2));
  inv1  gate2706(.a(s_308), .O(gate154inter3));
  inv1  gate2707(.a(s_309), .O(gate154inter4));
  nand2 gate2708(.a(gate154inter4), .b(gate154inter3), .O(gate154inter5));
  nor2  gate2709(.a(gate154inter5), .b(gate154inter2), .O(gate154inter6));
  inv1  gate2710(.a(G429), .O(gate154inter7));
  inv1  gate2711(.a(G522), .O(gate154inter8));
  nand2 gate2712(.a(gate154inter8), .b(gate154inter7), .O(gate154inter9));
  nand2 gate2713(.a(s_309), .b(gate154inter3), .O(gate154inter10));
  nor2  gate2714(.a(gate154inter10), .b(gate154inter9), .O(gate154inter11));
  nor2  gate2715(.a(gate154inter11), .b(gate154inter6), .O(gate154inter12));
  nand2 gate2716(.a(gate154inter12), .b(gate154inter1), .O(G571));

  xor2  gate603(.a(G525), .b(G432), .O(gate155inter0));
  nand2 gate604(.a(gate155inter0), .b(s_8), .O(gate155inter1));
  and2  gate605(.a(G525), .b(G432), .O(gate155inter2));
  inv1  gate606(.a(s_8), .O(gate155inter3));
  inv1  gate607(.a(s_9), .O(gate155inter4));
  nand2 gate608(.a(gate155inter4), .b(gate155inter3), .O(gate155inter5));
  nor2  gate609(.a(gate155inter5), .b(gate155inter2), .O(gate155inter6));
  inv1  gate610(.a(G432), .O(gate155inter7));
  inv1  gate611(.a(G525), .O(gate155inter8));
  nand2 gate612(.a(gate155inter8), .b(gate155inter7), .O(gate155inter9));
  nand2 gate613(.a(s_9), .b(gate155inter3), .O(gate155inter10));
  nor2  gate614(.a(gate155inter10), .b(gate155inter9), .O(gate155inter11));
  nor2  gate615(.a(gate155inter11), .b(gate155inter6), .O(gate155inter12));
  nand2 gate616(.a(gate155inter12), .b(gate155inter1), .O(G572));
nand2 gate156( .a(G435), .b(G525), .O(G573) );
nand2 gate157( .a(G438), .b(G528), .O(G574) );
nand2 gate158( .a(G441), .b(G528), .O(G575) );

  xor2  gate1947(.a(G531), .b(G444), .O(gate159inter0));
  nand2 gate1948(.a(gate159inter0), .b(s_200), .O(gate159inter1));
  and2  gate1949(.a(G531), .b(G444), .O(gate159inter2));
  inv1  gate1950(.a(s_200), .O(gate159inter3));
  inv1  gate1951(.a(s_201), .O(gate159inter4));
  nand2 gate1952(.a(gate159inter4), .b(gate159inter3), .O(gate159inter5));
  nor2  gate1953(.a(gate159inter5), .b(gate159inter2), .O(gate159inter6));
  inv1  gate1954(.a(G444), .O(gate159inter7));
  inv1  gate1955(.a(G531), .O(gate159inter8));
  nand2 gate1956(.a(gate159inter8), .b(gate159inter7), .O(gate159inter9));
  nand2 gate1957(.a(s_201), .b(gate159inter3), .O(gate159inter10));
  nor2  gate1958(.a(gate159inter10), .b(gate159inter9), .O(gate159inter11));
  nor2  gate1959(.a(gate159inter11), .b(gate159inter6), .O(gate159inter12));
  nand2 gate1960(.a(gate159inter12), .b(gate159inter1), .O(G576));
nand2 gate160( .a(G447), .b(G531), .O(G577) );

  xor2  gate813(.a(G534), .b(G450), .O(gate161inter0));
  nand2 gate814(.a(gate161inter0), .b(s_38), .O(gate161inter1));
  and2  gate815(.a(G534), .b(G450), .O(gate161inter2));
  inv1  gate816(.a(s_38), .O(gate161inter3));
  inv1  gate817(.a(s_39), .O(gate161inter4));
  nand2 gate818(.a(gate161inter4), .b(gate161inter3), .O(gate161inter5));
  nor2  gate819(.a(gate161inter5), .b(gate161inter2), .O(gate161inter6));
  inv1  gate820(.a(G450), .O(gate161inter7));
  inv1  gate821(.a(G534), .O(gate161inter8));
  nand2 gate822(.a(gate161inter8), .b(gate161inter7), .O(gate161inter9));
  nand2 gate823(.a(s_39), .b(gate161inter3), .O(gate161inter10));
  nor2  gate824(.a(gate161inter10), .b(gate161inter9), .O(gate161inter11));
  nor2  gate825(.a(gate161inter11), .b(gate161inter6), .O(gate161inter12));
  nand2 gate826(.a(gate161inter12), .b(gate161inter1), .O(G578));

  xor2  gate1779(.a(G534), .b(G453), .O(gate162inter0));
  nand2 gate1780(.a(gate162inter0), .b(s_176), .O(gate162inter1));
  and2  gate1781(.a(G534), .b(G453), .O(gate162inter2));
  inv1  gate1782(.a(s_176), .O(gate162inter3));
  inv1  gate1783(.a(s_177), .O(gate162inter4));
  nand2 gate1784(.a(gate162inter4), .b(gate162inter3), .O(gate162inter5));
  nor2  gate1785(.a(gate162inter5), .b(gate162inter2), .O(gate162inter6));
  inv1  gate1786(.a(G453), .O(gate162inter7));
  inv1  gate1787(.a(G534), .O(gate162inter8));
  nand2 gate1788(.a(gate162inter8), .b(gate162inter7), .O(gate162inter9));
  nand2 gate1789(.a(s_177), .b(gate162inter3), .O(gate162inter10));
  nor2  gate1790(.a(gate162inter10), .b(gate162inter9), .O(gate162inter11));
  nor2  gate1791(.a(gate162inter11), .b(gate162inter6), .O(gate162inter12));
  nand2 gate1792(.a(gate162inter12), .b(gate162inter1), .O(G579));
nand2 gate163( .a(G456), .b(G537), .O(G580) );

  xor2  gate2661(.a(G537), .b(G459), .O(gate164inter0));
  nand2 gate2662(.a(gate164inter0), .b(s_302), .O(gate164inter1));
  and2  gate2663(.a(G537), .b(G459), .O(gate164inter2));
  inv1  gate2664(.a(s_302), .O(gate164inter3));
  inv1  gate2665(.a(s_303), .O(gate164inter4));
  nand2 gate2666(.a(gate164inter4), .b(gate164inter3), .O(gate164inter5));
  nor2  gate2667(.a(gate164inter5), .b(gate164inter2), .O(gate164inter6));
  inv1  gate2668(.a(G459), .O(gate164inter7));
  inv1  gate2669(.a(G537), .O(gate164inter8));
  nand2 gate2670(.a(gate164inter8), .b(gate164inter7), .O(gate164inter9));
  nand2 gate2671(.a(s_303), .b(gate164inter3), .O(gate164inter10));
  nor2  gate2672(.a(gate164inter10), .b(gate164inter9), .O(gate164inter11));
  nor2  gate2673(.a(gate164inter11), .b(gate164inter6), .O(gate164inter12));
  nand2 gate2674(.a(gate164inter12), .b(gate164inter1), .O(G581));
nand2 gate165( .a(G462), .b(G540), .O(G582) );

  xor2  gate2689(.a(G540), .b(G465), .O(gate166inter0));
  nand2 gate2690(.a(gate166inter0), .b(s_306), .O(gate166inter1));
  and2  gate2691(.a(G540), .b(G465), .O(gate166inter2));
  inv1  gate2692(.a(s_306), .O(gate166inter3));
  inv1  gate2693(.a(s_307), .O(gate166inter4));
  nand2 gate2694(.a(gate166inter4), .b(gate166inter3), .O(gate166inter5));
  nor2  gate2695(.a(gate166inter5), .b(gate166inter2), .O(gate166inter6));
  inv1  gate2696(.a(G465), .O(gate166inter7));
  inv1  gate2697(.a(G540), .O(gate166inter8));
  nand2 gate2698(.a(gate166inter8), .b(gate166inter7), .O(gate166inter9));
  nand2 gate2699(.a(s_307), .b(gate166inter3), .O(gate166inter10));
  nor2  gate2700(.a(gate166inter10), .b(gate166inter9), .O(gate166inter11));
  nor2  gate2701(.a(gate166inter11), .b(gate166inter6), .O(gate166inter12));
  nand2 gate2702(.a(gate166inter12), .b(gate166inter1), .O(G583));

  xor2  gate1513(.a(G543), .b(G468), .O(gate167inter0));
  nand2 gate1514(.a(gate167inter0), .b(s_138), .O(gate167inter1));
  and2  gate1515(.a(G543), .b(G468), .O(gate167inter2));
  inv1  gate1516(.a(s_138), .O(gate167inter3));
  inv1  gate1517(.a(s_139), .O(gate167inter4));
  nand2 gate1518(.a(gate167inter4), .b(gate167inter3), .O(gate167inter5));
  nor2  gate1519(.a(gate167inter5), .b(gate167inter2), .O(gate167inter6));
  inv1  gate1520(.a(G468), .O(gate167inter7));
  inv1  gate1521(.a(G543), .O(gate167inter8));
  nand2 gate1522(.a(gate167inter8), .b(gate167inter7), .O(gate167inter9));
  nand2 gate1523(.a(s_139), .b(gate167inter3), .O(gate167inter10));
  nor2  gate1524(.a(gate167inter10), .b(gate167inter9), .O(gate167inter11));
  nor2  gate1525(.a(gate167inter11), .b(gate167inter6), .O(gate167inter12));
  nand2 gate1526(.a(gate167inter12), .b(gate167inter1), .O(G584));

  xor2  gate2969(.a(G543), .b(G471), .O(gate168inter0));
  nand2 gate2970(.a(gate168inter0), .b(s_346), .O(gate168inter1));
  and2  gate2971(.a(G543), .b(G471), .O(gate168inter2));
  inv1  gate2972(.a(s_346), .O(gate168inter3));
  inv1  gate2973(.a(s_347), .O(gate168inter4));
  nand2 gate2974(.a(gate168inter4), .b(gate168inter3), .O(gate168inter5));
  nor2  gate2975(.a(gate168inter5), .b(gate168inter2), .O(gate168inter6));
  inv1  gate2976(.a(G471), .O(gate168inter7));
  inv1  gate2977(.a(G543), .O(gate168inter8));
  nand2 gate2978(.a(gate168inter8), .b(gate168inter7), .O(gate168inter9));
  nand2 gate2979(.a(s_347), .b(gate168inter3), .O(gate168inter10));
  nor2  gate2980(.a(gate168inter10), .b(gate168inter9), .O(gate168inter11));
  nor2  gate2981(.a(gate168inter11), .b(gate168inter6), .O(gate168inter12));
  nand2 gate2982(.a(gate168inter12), .b(gate168inter1), .O(G585));
nand2 gate169( .a(G474), .b(G546), .O(G586) );
nand2 gate170( .a(G477), .b(G546), .O(G587) );
nand2 gate171( .a(G480), .b(G549), .O(G588) );
nand2 gate172( .a(G483), .b(G549), .O(G589) );
nand2 gate173( .a(G486), .b(G552), .O(G590) );
nand2 gate174( .a(G489), .b(G552), .O(G591) );
nand2 gate175( .a(G492), .b(G555), .O(G592) );
nand2 gate176( .a(G495), .b(G555), .O(G593) );
nand2 gate177( .a(G498), .b(G558), .O(G594) );
nand2 gate178( .a(G501), .b(G558), .O(G595) );
nand2 gate179( .a(G504), .b(G561), .O(G596) );
nand2 gate180( .a(G507), .b(G561), .O(G597) );
nand2 gate181( .a(G510), .b(G564), .O(G598) );
nand2 gate182( .a(G513), .b(G564), .O(G599) );
nand2 gate183( .a(G516), .b(G567), .O(G600) );
nand2 gate184( .a(G519), .b(G567), .O(G601) );
nand2 gate185( .a(G570), .b(G571), .O(G602) );
nand2 gate186( .a(G572), .b(G573), .O(G607) );

  xor2  gate1989(.a(G575), .b(G574), .O(gate187inter0));
  nand2 gate1990(.a(gate187inter0), .b(s_206), .O(gate187inter1));
  and2  gate1991(.a(G575), .b(G574), .O(gate187inter2));
  inv1  gate1992(.a(s_206), .O(gate187inter3));
  inv1  gate1993(.a(s_207), .O(gate187inter4));
  nand2 gate1994(.a(gate187inter4), .b(gate187inter3), .O(gate187inter5));
  nor2  gate1995(.a(gate187inter5), .b(gate187inter2), .O(gate187inter6));
  inv1  gate1996(.a(G574), .O(gate187inter7));
  inv1  gate1997(.a(G575), .O(gate187inter8));
  nand2 gate1998(.a(gate187inter8), .b(gate187inter7), .O(gate187inter9));
  nand2 gate1999(.a(s_207), .b(gate187inter3), .O(gate187inter10));
  nor2  gate2000(.a(gate187inter10), .b(gate187inter9), .O(gate187inter11));
  nor2  gate2001(.a(gate187inter11), .b(gate187inter6), .O(gate187inter12));
  nand2 gate2002(.a(gate187inter12), .b(gate187inter1), .O(G612));
nand2 gate188( .a(G576), .b(G577), .O(G617) );
nand2 gate189( .a(G578), .b(G579), .O(G622) );
nand2 gate190( .a(G580), .b(G581), .O(G627) );
nand2 gate191( .a(G582), .b(G583), .O(G632) );

  xor2  gate2745(.a(G585), .b(G584), .O(gate192inter0));
  nand2 gate2746(.a(gate192inter0), .b(s_314), .O(gate192inter1));
  and2  gate2747(.a(G585), .b(G584), .O(gate192inter2));
  inv1  gate2748(.a(s_314), .O(gate192inter3));
  inv1  gate2749(.a(s_315), .O(gate192inter4));
  nand2 gate2750(.a(gate192inter4), .b(gate192inter3), .O(gate192inter5));
  nor2  gate2751(.a(gate192inter5), .b(gate192inter2), .O(gate192inter6));
  inv1  gate2752(.a(G584), .O(gate192inter7));
  inv1  gate2753(.a(G585), .O(gate192inter8));
  nand2 gate2754(.a(gate192inter8), .b(gate192inter7), .O(gate192inter9));
  nand2 gate2755(.a(s_315), .b(gate192inter3), .O(gate192inter10));
  nor2  gate2756(.a(gate192inter10), .b(gate192inter9), .O(gate192inter11));
  nor2  gate2757(.a(gate192inter11), .b(gate192inter6), .O(gate192inter12));
  nand2 gate2758(.a(gate192inter12), .b(gate192inter1), .O(G637));
nand2 gate193( .a(G586), .b(G587), .O(G642) );

  xor2  gate2003(.a(G589), .b(G588), .O(gate194inter0));
  nand2 gate2004(.a(gate194inter0), .b(s_208), .O(gate194inter1));
  and2  gate2005(.a(G589), .b(G588), .O(gate194inter2));
  inv1  gate2006(.a(s_208), .O(gate194inter3));
  inv1  gate2007(.a(s_209), .O(gate194inter4));
  nand2 gate2008(.a(gate194inter4), .b(gate194inter3), .O(gate194inter5));
  nor2  gate2009(.a(gate194inter5), .b(gate194inter2), .O(gate194inter6));
  inv1  gate2010(.a(G588), .O(gate194inter7));
  inv1  gate2011(.a(G589), .O(gate194inter8));
  nand2 gate2012(.a(gate194inter8), .b(gate194inter7), .O(gate194inter9));
  nand2 gate2013(.a(s_209), .b(gate194inter3), .O(gate194inter10));
  nor2  gate2014(.a(gate194inter10), .b(gate194inter9), .O(gate194inter11));
  nor2  gate2015(.a(gate194inter11), .b(gate194inter6), .O(gate194inter12));
  nand2 gate2016(.a(gate194inter12), .b(gate194inter1), .O(G645));
nand2 gate195( .a(G590), .b(G591), .O(G648) );
nand2 gate196( .a(G592), .b(G593), .O(G651) );
nand2 gate197( .a(G594), .b(G595), .O(G654) );
nand2 gate198( .a(G596), .b(G597), .O(G657) );
nand2 gate199( .a(G598), .b(G599), .O(G660) );
nand2 gate200( .a(G600), .b(G601), .O(G663) );

  xor2  gate1653(.a(G607), .b(G602), .O(gate201inter0));
  nand2 gate1654(.a(gate201inter0), .b(s_158), .O(gate201inter1));
  and2  gate1655(.a(G607), .b(G602), .O(gate201inter2));
  inv1  gate1656(.a(s_158), .O(gate201inter3));
  inv1  gate1657(.a(s_159), .O(gate201inter4));
  nand2 gate1658(.a(gate201inter4), .b(gate201inter3), .O(gate201inter5));
  nor2  gate1659(.a(gate201inter5), .b(gate201inter2), .O(gate201inter6));
  inv1  gate1660(.a(G602), .O(gate201inter7));
  inv1  gate1661(.a(G607), .O(gate201inter8));
  nand2 gate1662(.a(gate201inter8), .b(gate201inter7), .O(gate201inter9));
  nand2 gate1663(.a(s_159), .b(gate201inter3), .O(gate201inter10));
  nor2  gate1664(.a(gate201inter10), .b(gate201inter9), .O(gate201inter11));
  nor2  gate1665(.a(gate201inter11), .b(gate201inter6), .O(gate201inter12));
  nand2 gate1666(.a(gate201inter12), .b(gate201inter1), .O(G666));
nand2 gate202( .a(G612), .b(G617), .O(G669) );
nand2 gate203( .a(G602), .b(G612), .O(G672) );
nand2 gate204( .a(G607), .b(G617), .O(G675) );

  xor2  gate883(.a(G627), .b(G622), .O(gate205inter0));
  nand2 gate884(.a(gate205inter0), .b(s_48), .O(gate205inter1));
  and2  gate885(.a(G627), .b(G622), .O(gate205inter2));
  inv1  gate886(.a(s_48), .O(gate205inter3));
  inv1  gate887(.a(s_49), .O(gate205inter4));
  nand2 gate888(.a(gate205inter4), .b(gate205inter3), .O(gate205inter5));
  nor2  gate889(.a(gate205inter5), .b(gate205inter2), .O(gate205inter6));
  inv1  gate890(.a(G622), .O(gate205inter7));
  inv1  gate891(.a(G627), .O(gate205inter8));
  nand2 gate892(.a(gate205inter8), .b(gate205inter7), .O(gate205inter9));
  nand2 gate893(.a(s_49), .b(gate205inter3), .O(gate205inter10));
  nor2  gate894(.a(gate205inter10), .b(gate205inter9), .O(gate205inter11));
  nor2  gate895(.a(gate205inter11), .b(gate205inter6), .O(gate205inter12));
  nand2 gate896(.a(gate205inter12), .b(gate205inter1), .O(G678));

  xor2  gate1667(.a(G637), .b(G632), .O(gate206inter0));
  nand2 gate1668(.a(gate206inter0), .b(s_160), .O(gate206inter1));
  and2  gate1669(.a(G637), .b(G632), .O(gate206inter2));
  inv1  gate1670(.a(s_160), .O(gate206inter3));
  inv1  gate1671(.a(s_161), .O(gate206inter4));
  nand2 gate1672(.a(gate206inter4), .b(gate206inter3), .O(gate206inter5));
  nor2  gate1673(.a(gate206inter5), .b(gate206inter2), .O(gate206inter6));
  inv1  gate1674(.a(G632), .O(gate206inter7));
  inv1  gate1675(.a(G637), .O(gate206inter8));
  nand2 gate1676(.a(gate206inter8), .b(gate206inter7), .O(gate206inter9));
  nand2 gate1677(.a(s_161), .b(gate206inter3), .O(gate206inter10));
  nor2  gate1678(.a(gate206inter10), .b(gate206inter9), .O(gate206inter11));
  nor2  gate1679(.a(gate206inter11), .b(gate206inter6), .O(gate206inter12));
  nand2 gate1680(.a(gate206inter12), .b(gate206inter1), .O(G681));

  xor2  gate1821(.a(G632), .b(G622), .O(gate207inter0));
  nand2 gate1822(.a(gate207inter0), .b(s_182), .O(gate207inter1));
  and2  gate1823(.a(G632), .b(G622), .O(gate207inter2));
  inv1  gate1824(.a(s_182), .O(gate207inter3));
  inv1  gate1825(.a(s_183), .O(gate207inter4));
  nand2 gate1826(.a(gate207inter4), .b(gate207inter3), .O(gate207inter5));
  nor2  gate1827(.a(gate207inter5), .b(gate207inter2), .O(gate207inter6));
  inv1  gate1828(.a(G622), .O(gate207inter7));
  inv1  gate1829(.a(G632), .O(gate207inter8));
  nand2 gate1830(.a(gate207inter8), .b(gate207inter7), .O(gate207inter9));
  nand2 gate1831(.a(s_183), .b(gate207inter3), .O(gate207inter10));
  nor2  gate1832(.a(gate207inter10), .b(gate207inter9), .O(gate207inter11));
  nor2  gate1833(.a(gate207inter11), .b(gate207inter6), .O(gate207inter12));
  nand2 gate1834(.a(gate207inter12), .b(gate207inter1), .O(G684));

  xor2  gate743(.a(G637), .b(G627), .O(gate208inter0));
  nand2 gate744(.a(gate208inter0), .b(s_28), .O(gate208inter1));
  and2  gate745(.a(G637), .b(G627), .O(gate208inter2));
  inv1  gate746(.a(s_28), .O(gate208inter3));
  inv1  gate747(.a(s_29), .O(gate208inter4));
  nand2 gate748(.a(gate208inter4), .b(gate208inter3), .O(gate208inter5));
  nor2  gate749(.a(gate208inter5), .b(gate208inter2), .O(gate208inter6));
  inv1  gate750(.a(G627), .O(gate208inter7));
  inv1  gate751(.a(G637), .O(gate208inter8));
  nand2 gate752(.a(gate208inter8), .b(gate208inter7), .O(gate208inter9));
  nand2 gate753(.a(s_29), .b(gate208inter3), .O(gate208inter10));
  nor2  gate754(.a(gate208inter10), .b(gate208inter9), .O(gate208inter11));
  nor2  gate755(.a(gate208inter11), .b(gate208inter6), .O(gate208inter12));
  nand2 gate756(.a(gate208inter12), .b(gate208inter1), .O(G687));
nand2 gate209( .a(G602), .b(G666), .O(G690) );
nand2 gate210( .a(G607), .b(G666), .O(G691) );

  xor2  gate2871(.a(G669), .b(G612), .O(gate211inter0));
  nand2 gate2872(.a(gate211inter0), .b(s_332), .O(gate211inter1));
  and2  gate2873(.a(G669), .b(G612), .O(gate211inter2));
  inv1  gate2874(.a(s_332), .O(gate211inter3));
  inv1  gate2875(.a(s_333), .O(gate211inter4));
  nand2 gate2876(.a(gate211inter4), .b(gate211inter3), .O(gate211inter5));
  nor2  gate2877(.a(gate211inter5), .b(gate211inter2), .O(gate211inter6));
  inv1  gate2878(.a(G612), .O(gate211inter7));
  inv1  gate2879(.a(G669), .O(gate211inter8));
  nand2 gate2880(.a(gate211inter8), .b(gate211inter7), .O(gate211inter9));
  nand2 gate2881(.a(s_333), .b(gate211inter3), .O(gate211inter10));
  nor2  gate2882(.a(gate211inter10), .b(gate211inter9), .O(gate211inter11));
  nor2  gate2883(.a(gate211inter11), .b(gate211inter6), .O(gate211inter12));
  nand2 gate2884(.a(gate211inter12), .b(gate211inter1), .O(G692));
nand2 gate212( .a(G617), .b(G669), .O(G693) );
nand2 gate213( .a(G602), .b(G672), .O(G694) );
nand2 gate214( .a(G612), .b(G672), .O(G695) );
nand2 gate215( .a(G607), .b(G675), .O(G696) );

  xor2  gate953(.a(G675), .b(G617), .O(gate216inter0));
  nand2 gate954(.a(gate216inter0), .b(s_58), .O(gate216inter1));
  and2  gate955(.a(G675), .b(G617), .O(gate216inter2));
  inv1  gate956(.a(s_58), .O(gate216inter3));
  inv1  gate957(.a(s_59), .O(gate216inter4));
  nand2 gate958(.a(gate216inter4), .b(gate216inter3), .O(gate216inter5));
  nor2  gate959(.a(gate216inter5), .b(gate216inter2), .O(gate216inter6));
  inv1  gate960(.a(G617), .O(gate216inter7));
  inv1  gate961(.a(G675), .O(gate216inter8));
  nand2 gate962(.a(gate216inter8), .b(gate216inter7), .O(gate216inter9));
  nand2 gate963(.a(s_59), .b(gate216inter3), .O(gate216inter10));
  nor2  gate964(.a(gate216inter10), .b(gate216inter9), .O(gate216inter11));
  nor2  gate965(.a(gate216inter11), .b(gate216inter6), .O(gate216inter12));
  nand2 gate966(.a(gate216inter12), .b(gate216inter1), .O(G697));
nand2 gate217( .a(G622), .b(G678), .O(G698) );

  xor2  gate1807(.a(G678), .b(G627), .O(gate218inter0));
  nand2 gate1808(.a(gate218inter0), .b(s_180), .O(gate218inter1));
  and2  gate1809(.a(G678), .b(G627), .O(gate218inter2));
  inv1  gate1810(.a(s_180), .O(gate218inter3));
  inv1  gate1811(.a(s_181), .O(gate218inter4));
  nand2 gate1812(.a(gate218inter4), .b(gate218inter3), .O(gate218inter5));
  nor2  gate1813(.a(gate218inter5), .b(gate218inter2), .O(gate218inter6));
  inv1  gate1814(.a(G627), .O(gate218inter7));
  inv1  gate1815(.a(G678), .O(gate218inter8));
  nand2 gate1816(.a(gate218inter8), .b(gate218inter7), .O(gate218inter9));
  nand2 gate1817(.a(s_181), .b(gate218inter3), .O(gate218inter10));
  nor2  gate1818(.a(gate218inter10), .b(gate218inter9), .O(gate218inter11));
  nor2  gate1819(.a(gate218inter11), .b(gate218inter6), .O(gate218inter12));
  nand2 gate1820(.a(gate218inter12), .b(gate218inter1), .O(G699));
nand2 gate219( .a(G632), .b(G681), .O(G700) );
nand2 gate220( .a(G637), .b(G681), .O(G701) );

  xor2  gate2339(.a(G684), .b(G622), .O(gate221inter0));
  nand2 gate2340(.a(gate221inter0), .b(s_256), .O(gate221inter1));
  and2  gate2341(.a(G684), .b(G622), .O(gate221inter2));
  inv1  gate2342(.a(s_256), .O(gate221inter3));
  inv1  gate2343(.a(s_257), .O(gate221inter4));
  nand2 gate2344(.a(gate221inter4), .b(gate221inter3), .O(gate221inter5));
  nor2  gate2345(.a(gate221inter5), .b(gate221inter2), .O(gate221inter6));
  inv1  gate2346(.a(G622), .O(gate221inter7));
  inv1  gate2347(.a(G684), .O(gate221inter8));
  nand2 gate2348(.a(gate221inter8), .b(gate221inter7), .O(gate221inter9));
  nand2 gate2349(.a(s_257), .b(gate221inter3), .O(gate221inter10));
  nor2  gate2350(.a(gate221inter10), .b(gate221inter9), .O(gate221inter11));
  nor2  gate2351(.a(gate221inter11), .b(gate221inter6), .O(gate221inter12));
  nand2 gate2352(.a(gate221inter12), .b(gate221inter1), .O(G702));
nand2 gate222( .a(G632), .b(G684), .O(G703) );
nand2 gate223( .a(G627), .b(G687), .O(G704) );

  xor2  gate799(.a(G687), .b(G637), .O(gate224inter0));
  nand2 gate800(.a(gate224inter0), .b(s_36), .O(gate224inter1));
  and2  gate801(.a(G687), .b(G637), .O(gate224inter2));
  inv1  gate802(.a(s_36), .O(gate224inter3));
  inv1  gate803(.a(s_37), .O(gate224inter4));
  nand2 gate804(.a(gate224inter4), .b(gate224inter3), .O(gate224inter5));
  nor2  gate805(.a(gate224inter5), .b(gate224inter2), .O(gate224inter6));
  inv1  gate806(.a(G637), .O(gate224inter7));
  inv1  gate807(.a(G687), .O(gate224inter8));
  nand2 gate808(.a(gate224inter8), .b(gate224inter7), .O(gate224inter9));
  nand2 gate809(.a(s_37), .b(gate224inter3), .O(gate224inter10));
  nor2  gate810(.a(gate224inter10), .b(gate224inter9), .O(gate224inter11));
  nor2  gate811(.a(gate224inter11), .b(gate224inter6), .O(gate224inter12));
  nand2 gate812(.a(gate224inter12), .b(gate224inter1), .O(G705));
nand2 gate225( .a(G690), .b(G691), .O(G706) );
nand2 gate226( .a(G692), .b(G693), .O(G709) );
nand2 gate227( .a(G694), .b(G695), .O(G712) );
nand2 gate228( .a(G696), .b(G697), .O(G715) );
nand2 gate229( .a(G698), .b(G699), .O(G718) );

  xor2  gate2857(.a(G701), .b(G700), .O(gate230inter0));
  nand2 gate2858(.a(gate230inter0), .b(s_330), .O(gate230inter1));
  and2  gate2859(.a(G701), .b(G700), .O(gate230inter2));
  inv1  gate2860(.a(s_330), .O(gate230inter3));
  inv1  gate2861(.a(s_331), .O(gate230inter4));
  nand2 gate2862(.a(gate230inter4), .b(gate230inter3), .O(gate230inter5));
  nor2  gate2863(.a(gate230inter5), .b(gate230inter2), .O(gate230inter6));
  inv1  gate2864(.a(G700), .O(gate230inter7));
  inv1  gate2865(.a(G701), .O(gate230inter8));
  nand2 gate2866(.a(gate230inter8), .b(gate230inter7), .O(gate230inter9));
  nand2 gate2867(.a(s_331), .b(gate230inter3), .O(gate230inter10));
  nor2  gate2868(.a(gate230inter10), .b(gate230inter9), .O(gate230inter11));
  nor2  gate2869(.a(gate230inter11), .b(gate230inter6), .O(gate230inter12));
  nand2 gate2870(.a(gate230inter12), .b(gate230inter1), .O(G721));

  xor2  gate2787(.a(G703), .b(G702), .O(gate231inter0));
  nand2 gate2788(.a(gate231inter0), .b(s_320), .O(gate231inter1));
  and2  gate2789(.a(G703), .b(G702), .O(gate231inter2));
  inv1  gate2790(.a(s_320), .O(gate231inter3));
  inv1  gate2791(.a(s_321), .O(gate231inter4));
  nand2 gate2792(.a(gate231inter4), .b(gate231inter3), .O(gate231inter5));
  nor2  gate2793(.a(gate231inter5), .b(gate231inter2), .O(gate231inter6));
  inv1  gate2794(.a(G702), .O(gate231inter7));
  inv1  gate2795(.a(G703), .O(gate231inter8));
  nand2 gate2796(.a(gate231inter8), .b(gate231inter7), .O(gate231inter9));
  nand2 gate2797(.a(s_321), .b(gate231inter3), .O(gate231inter10));
  nor2  gate2798(.a(gate231inter10), .b(gate231inter9), .O(gate231inter11));
  nor2  gate2799(.a(gate231inter11), .b(gate231inter6), .O(gate231inter12));
  nand2 gate2800(.a(gate231inter12), .b(gate231inter1), .O(G724));
nand2 gate232( .a(G704), .b(G705), .O(G727) );
nand2 gate233( .a(G242), .b(G718), .O(G730) );
nand2 gate234( .a(G245), .b(G721), .O(G733) );
nand2 gate235( .a(G248), .b(G724), .O(G736) );

  xor2  gate1723(.a(G727), .b(G251), .O(gate236inter0));
  nand2 gate1724(.a(gate236inter0), .b(s_168), .O(gate236inter1));
  and2  gate1725(.a(G727), .b(G251), .O(gate236inter2));
  inv1  gate1726(.a(s_168), .O(gate236inter3));
  inv1  gate1727(.a(s_169), .O(gate236inter4));
  nand2 gate1728(.a(gate236inter4), .b(gate236inter3), .O(gate236inter5));
  nor2  gate1729(.a(gate236inter5), .b(gate236inter2), .O(gate236inter6));
  inv1  gate1730(.a(G251), .O(gate236inter7));
  inv1  gate1731(.a(G727), .O(gate236inter8));
  nand2 gate1732(.a(gate236inter8), .b(gate236inter7), .O(gate236inter9));
  nand2 gate1733(.a(s_169), .b(gate236inter3), .O(gate236inter10));
  nor2  gate1734(.a(gate236inter10), .b(gate236inter9), .O(gate236inter11));
  nor2  gate1735(.a(gate236inter11), .b(gate236inter6), .O(gate236inter12));
  nand2 gate1736(.a(gate236inter12), .b(gate236inter1), .O(G739));
nand2 gate237( .a(G254), .b(G706), .O(G742) );

  xor2  gate1303(.a(G709), .b(G257), .O(gate238inter0));
  nand2 gate1304(.a(gate238inter0), .b(s_108), .O(gate238inter1));
  and2  gate1305(.a(G709), .b(G257), .O(gate238inter2));
  inv1  gate1306(.a(s_108), .O(gate238inter3));
  inv1  gate1307(.a(s_109), .O(gate238inter4));
  nand2 gate1308(.a(gate238inter4), .b(gate238inter3), .O(gate238inter5));
  nor2  gate1309(.a(gate238inter5), .b(gate238inter2), .O(gate238inter6));
  inv1  gate1310(.a(G257), .O(gate238inter7));
  inv1  gate1311(.a(G709), .O(gate238inter8));
  nand2 gate1312(.a(gate238inter8), .b(gate238inter7), .O(gate238inter9));
  nand2 gate1313(.a(s_109), .b(gate238inter3), .O(gate238inter10));
  nor2  gate1314(.a(gate238inter10), .b(gate238inter9), .O(gate238inter11));
  nor2  gate1315(.a(gate238inter11), .b(gate238inter6), .O(gate238inter12));
  nand2 gate1316(.a(gate238inter12), .b(gate238inter1), .O(G745));

  xor2  gate1793(.a(G712), .b(G260), .O(gate239inter0));
  nand2 gate1794(.a(gate239inter0), .b(s_178), .O(gate239inter1));
  and2  gate1795(.a(G712), .b(G260), .O(gate239inter2));
  inv1  gate1796(.a(s_178), .O(gate239inter3));
  inv1  gate1797(.a(s_179), .O(gate239inter4));
  nand2 gate1798(.a(gate239inter4), .b(gate239inter3), .O(gate239inter5));
  nor2  gate1799(.a(gate239inter5), .b(gate239inter2), .O(gate239inter6));
  inv1  gate1800(.a(G260), .O(gate239inter7));
  inv1  gate1801(.a(G712), .O(gate239inter8));
  nand2 gate1802(.a(gate239inter8), .b(gate239inter7), .O(gate239inter9));
  nand2 gate1803(.a(s_179), .b(gate239inter3), .O(gate239inter10));
  nor2  gate1804(.a(gate239inter10), .b(gate239inter9), .O(gate239inter11));
  nor2  gate1805(.a(gate239inter11), .b(gate239inter6), .O(gate239inter12));
  nand2 gate1806(.a(gate239inter12), .b(gate239inter1), .O(G748));

  xor2  gate939(.a(G715), .b(G263), .O(gate240inter0));
  nand2 gate940(.a(gate240inter0), .b(s_56), .O(gate240inter1));
  and2  gate941(.a(G715), .b(G263), .O(gate240inter2));
  inv1  gate942(.a(s_56), .O(gate240inter3));
  inv1  gate943(.a(s_57), .O(gate240inter4));
  nand2 gate944(.a(gate240inter4), .b(gate240inter3), .O(gate240inter5));
  nor2  gate945(.a(gate240inter5), .b(gate240inter2), .O(gate240inter6));
  inv1  gate946(.a(G263), .O(gate240inter7));
  inv1  gate947(.a(G715), .O(gate240inter8));
  nand2 gate948(.a(gate240inter8), .b(gate240inter7), .O(gate240inter9));
  nand2 gate949(.a(s_57), .b(gate240inter3), .O(gate240inter10));
  nor2  gate950(.a(gate240inter10), .b(gate240inter9), .O(gate240inter11));
  nor2  gate951(.a(gate240inter11), .b(gate240inter6), .O(gate240inter12));
  nand2 gate952(.a(gate240inter12), .b(gate240inter1), .O(G751));
nand2 gate241( .a(G242), .b(G730), .O(G754) );
nand2 gate242( .a(G718), .b(G730), .O(G755) );
nand2 gate243( .a(G245), .b(G733), .O(G756) );
nand2 gate244( .a(G721), .b(G733), .O(G757) );
nand2 gate245( .a(G248), .b(G736), .O(G758) );

  xor2  gate1359(.a(G736), .b(G724), .O(gate246inter0));
  nand2 gate1360(.a(gate246inter0), .b(s_116), .O(gate246inter1));
  and2  gate1361(.a(G736), .b(G724), .O(gate246inter2));
  inv1  gate1362(.a(s_116), .O(gate246inter3));
  inv1  gate1363(.a(s_117), .O(gate246inter4));
  nand2 gate1364(.a(gate246inter4), .b(gate246inter3), .O(gate246inter5));
  nor2  gate1365(.a(gate246inter5), .b(gate246inter2), .O(gate246inter6));
  inv1  gate1366(.a(G724), .O(gate246inter7));
  inv1  gate1367(.a(G736), .O(gate246inter8));
  nand2 gate1368(.a(gate246inter8), .b(gate246inter7), .O(gate246inter9));
  nand2 gate1369(.a(s_117), .b(gate246inter3), .O(gate246inter10));
  nor2  gate1370(.a(gate246inter10), .b(gate246inter9), .O(gate246inter11));
  nor2  gate1371(.a(gate246inter11), .b(gate246inter6), .O(gate246inter12));
  nand2 gate1372(.a(gate246inter12), .b(gate246inter1), .O(G759));

  xor2  gate687(.a(G739), .b(G251), .O(gate247inter0));
  nand2 gate688(.a(gate247inter0), .b(s_20), .O(gate247inter1));
  and2  gate689(.a(G739), .b(G251), .O(gate247inter2));
  inv1  gate690(.a(s_20), .O(gate247inter3));
  inv1  gate691(.a(s_21), .O(gate247inter4));
  nand2 gate692(.a(gate247inter4), .b(gate247inter3), .O(gate247inter5));
  nor2  gate693(.a(gate247inter5), .b(gate247inter2), .O(gate247inter6));
  inv1  gate694(.a(G251), .O(gate247inter7));
  inv1  gate695(.a(G739), .O(gate247inter8));
  nand2 gate696(.a(gate247inter8), .b(gate247inter7), .O(gate247inter9));
  nand2 gate697(.a(s_21), .b(gate247inter3), .O(gate247inter10));
  nor2  gate698(.a(gate247inter10), .b(gate247inter9), .O(gate247inter11));
  nor2  gate699(.a(gate247inter11), .b(gate247inter6), .O(gate247inter12));
  nand2 gate700(.a(gate247inter12), .b(gate247inter1), .O(G760));
nand2 gate248( .a(G727), .b(G739), .O(G761) );
nand2 gate249( .a(G254), .b(G742), .O(G762) );
nand2 gate250( .a(G706), .b(G742), .O(G763) );

  xor2  gate2577(.a(G745), .b(G257), .O(gate251inter0));
  nand2 gate2578(.a(gate251inter0), .b(s_290), .O(gate251inter1));
  and2  gate2579(.a(G745), .b(G257), .O(gate251inter2));
  inv1  gate2580(.a(s_290), .O(gate251inter3));
  inv1  gate2581(.a(s_291), .O(gate251inter4));
  nand2 gate2582(.a(gate251inter4), .b(gate251inter3), .O(gate251inter5));
  nor2  gate2583(.a(gate251inter5), .b(gate251inter2), .O(gate251inter6));
  inv1  gate2584(.a(G257), .O(gate251inter7));
  inv1  gate2585(.a(G745), .O(gate251inter8));
  nand2 gate2586(.a(gate251inter8), .b(gate251inter7), .O(gate251inter9));
  nand2 gate2587(.a(s_291), .b(gate251inter3), .O(gate251inter10));
  nor2  gate2588(.a(gate251inter10), .b(gate251inter9), .O(gate251inter11));
  nor2  gate2589(.a(gate251inter11), .b(gate251inter6), .O(gate251inter12));
  nand2 gate2590(.a(gate251inter12), .b(gate251inter1), .O(G764));

  xor2  gate2493(.a(G745), .b(G709), .O(gate252inter0));
  nand2 gate2494(.a(gate252inter0), .b(s_278), .O(gate252inter1));
  and2  gate2495(.a(G745), .b(G709), .O(gate252inter2));
  inv1  gate2496(.a(s_278), .O(gate252inter3));
  inv1  gate2497(.a(s_279), .O(gate252inter4));
  nand2 gate2498(.a(gate252inter4), .b(gate252inter3), .O(gate252inter5));
  nor2  gate2499(.a(gate252inter5), .b(gate252inter2), .O(gate252inter6));
  inv1  gate2500(.a(G709), .O(gate252inter7));
  inv1  gate2501(.a(G745), .O(gate252inter8));
  nand2 gate2502(.a(gate252inter8), .b(gate252inter7), .O(gate252inter9));
  nand2 gate2503(.a(s_279), .b(gate252inter3), .O(gate252inter10));
  nor2  gate2504(.a(gate252inter10), .b(gate252inter9), .O(gate252inter11));
  nor2  gate2505(.a(gate252inter11), .b(gate252inter6), .O(gate252inter12));
  nand2 gate2506(.a(gate252inter12), .b(gate252inter1), .O(G765));
nand2 gate253( .a(G260), .b(G748), .O(G766) );

  xor2  gate897(.a(G748), .b(G712), .O(gate254inter0));
  nand2 gate898(.a(gate254inter0), .b(s_50), .O(gate254inter1));
  and2  gate899(.a(G748), .b(G712), .O(gate254inter2));
  inv1  gate900(.a(s_50), .O(gate254inter3));
  inv1  gate901(.a(s_51), .O(gate254inter4));
  nand2 gate902(.a(gate254inter4), .b(gate254inter3), .O(gate254inter5));
  nor2  gate903(.a(gate254inter5), .b(gate254inter2), .O(gate254inter6));
  inv1  gate904(.a(G712), .O(gate254inter7));
  inv1  gate905(.a(G748), .O(gate254inter8));
  nand2 gate906(.a(gate254inter8), .b(gate254inter7), .O(gate254inter9));
  nand2 gate907(.a(s_51), .b(gate254inter3), .O(gate254inter10));
  nor2  gate908(.a(gate254inter10), .b(gate254inter9), .O(gate254inter11));
  nor2  gate909(.a(gate254inter11), .b(gate254inter6), .O(gate254inter12));
  nand2 gate910(.a(gate254inter12), .b(gate254inter1), .O(G767));
nand2 gate255( .a(G263), .b(G751), .O(G768) );

  xor2  gate589(.a(G751), .b(G715), .O(gate256inter0));
  nand2 gate590(.a(gate256inter0), .b(s_6), .O(gate256inter1));
  and2  gate591(.a(G751), .b(G715), .O(gate256inter2));
  inv1  gate592(.a(s_6), .O(gate256inter3));
  inv1  gate593(.a(s_7), .O(gate256inter4));
  nand2 gate594(.a(gate256inter4), .b(gate256inter3), .O(gate256inter5));
  nor2  gate595(.a(gate256inter5), .b(gate256inter2), .O(gate256inter6));
  inv1  gate596(.a(G715), .O(gate256inter7));
  inv1  gate597(.a(G751), .O(gate256inter8));
  nand2 gate598(.a(gate256inter8), .b(gate256inter7), .O(gate256inter9));
  nand2 gate599(.a(s_7), .b(gate256inter3), .O(gate256inter10));
  nor2  gate600(.a(gate256inter10), .b(gate256inter9), .O(gate256inter11));
  nor2  gate601(.a(gate256inter11), .b(gate256inter6), .O(gate256inter12));
  nand2 gate602(.a(gate256inter12), .b(gate256inter1), .O(G769));
nand2 gate257( .a(G754), .b(G755), .O(G770) );
nand2 gate258( .a(G756), .b(G757), .O(G773) );
nand2 gate259( .a(G758), .b(G759), .O(G776) );

  xor2  gate1443(.a(G761), .b(G760), .O(gate260inter0));
  nand2 gate1444(.a(gate260inter0), .b(s_128), .O(gate260inter1));
  and2  gate1445(.a(G761), .b(G760), .O(gate260inter2));
  inv1  gate1446(.a(s_128), .O(gate260inter3));
  inv1  gate1447(.a(s_129), .O(gate260inter4));
  nand2 gate1448(.a(gate260inter4), .b(gate260inter3), .O(gate260inter5));
  nor2  gate1449(.a(gate260inter5), .b(gate260inter2), .O(gate260inter6));
  inv1  gate1450(.a(G760), .O(gate260inter7));
  inv1  gate1451(.a(G761), .O(gate260inter8));
  nand2 gate1452(.a(gate260inter8), .b(gate260inter7), .O(gate260inter9));
  nand2 gate1453(.a(s_129), .b(gate260inter3), .O(gate260inter10));
  nor2  gate1454(.a(gate260inter10), .b(gate260inter9), .O(gate260inter11));
  nor2  gate1455(.a(gate260inter11), .b(gate260inter6), .O(gate260inter12));
  nand2 gate1456(.a(gate260inter12), .b(gate260inter1), .O(G779));
nand2 gate261( .a(G762), .b(G763), .O(G782) );

  xor2  gate2479(.a(G765), .b(G764), .O(gate262inter0));
  nand2 gate2480(.a(gate262inter0), .b(s_276), .O(gate262inter1));
  and2  gate2481(.a(G765), .b(G764), .O(gate262inter2));
  inv1  gate2482(.a(s_276), .O(gate262inter3));
  inv1  gate2483(.a(s_277), .O(gate262inter4));
  nand2 gate2484(.a(gate262inter4), .b(gate262inter3), .O(gate262inter5));
  nor2  gate2485(.a(gate262inter5), .b(gate262inter2), .O(gate262inter6));
  inv1  gate2486(.a(G764), .O(gate262inter7));
  inv1  gate2487(.a(G765), .O(gate262inter8));
  nand2 gate2488(.a(gate262inter8), .b(gate262inter7), .O(gate262inter9));
  nand2 gate2489(.a(s_277), .b(gate262inter3), .O(gate262inter10));
  nor2  gate2490(.a(gate262inter10), .b(gate262inter9), .O(gate262inter11));
  nor2  gate2491(.a(gate262inter11), .b(gate262inter6), .O(gate262inter12));
  nand2 gate2492(.a(gate262inter12), .b(gate262inter1), .O(G785));

  xor2  gate771(.a(G767), .b(G766), .O(gate263inter0));
  nand2 gate772(.a(gate263inter0), .b(s_32), .O(gate263inter1));
  and2  gate773(.a(G767), .b(G766), .O(gate263inter2));
  inv1  gate774(.a(s_32), .O(gate263inter3));
  inv1  gate775(.a(s_33), .O(gate263inter4));
  nand2 gate776(.a(gate263inter4), .b(gate263inter3), .O(gate263inter5));
  nor2  gate777(.a(gate263inter5), .b(gate263inter2), .O(gate263inter6));
  inv1  gate778(.a(G766), .O(gate263inter7));
  inv1  gate779(.a(G767), .O(gate263inter8));
  nand2 gate780(.a(gate263inter8), .b(gate263inter7), .O(gate263inter9));
  nand2 gate781(.a(s_33), .b(gate263inter3), .O(gate263inter10));
  nor2  gate782(.a(gate263inter10), .b(gate263inter9), .O(gate263inter11));
  nor2  gate783(.a(gate263inter11), .b(gate263inter6), .O(gate263inter12));
  nand2 gate784(.a(gate263inter12), .b(gate263inter1), .O(G788));

  xor2  gate1401(.a(G769), .b(G768), .O(gate264inter0));
  nand2 gate1402(.a(gate264inter0), .b(s_122), .O(gate264inter1));
  and2  gate1403(.a(G769), .b(G768), .O(gate264inter2));
  inv1  gate1404(.a(s_122), .O(gate264inter3));
  inv1  gate1405(.a(s_123), .O(gate264inter4));
  nand2 gate1406(.a(gate264inter4), .b(gate264inter3), .O(gate264inter5));
  nor2  gate1407(.a(gate264inter5), .b(gate264inter2), .O(gate264inter6));
  inv1  gate1408(.a(G768), .O(gate264inter7));
  inv1  gate1409(.a(G769), .O(gate264inter8));
  nand2 gate1410(.a(gate264inter8), .b(gate264inter7), .O(gate264inter9));
  nand2 gate1411(.a(s_123), .b(gate264inter3), .O(gate264inter10));
  nor2  gate1412(.a(gate264inter10), .b(gate264inter9), .O(gate264inter11));
  nor2  gate1413(.a(gate264inter11), .b(gate264inter6), .O(gate264inter12));
  nand2 gate1414(.a(gate264inter12), .b(gate264inter1), .O(G791));
nand2 gate265( .a(G642), .b(G770), .O(G794) );
nand2 gate266( .a(G645), .b(G773), .O(G797) );
nand2 gate267( .a(G648), .b(G776), .O(G800) );

  xor2  gate2941(.a(G779), .b(G651), .O(gate268inter0));
  nand2 gate2942(.a(gate268inter0), .b(s_342), .O(gate268inter1));
  and2  gate2943(.a(G779), .b(G651), .O(gate268inter2));
  inv1  gate2944(.a(s_342), .O(gate268inter3));
  inv1  gate2945(.a(s_343), .O(gate268inter4));
  nand2 gate2946(.a(gate268inter4), .b(gate268inter3), .O(gate268inter5));
  nor2  gate2947(.a(gate268inter5), .b(gate268inter2), .O(gate268inter6));
  inv1  gate2948(.a(G651), .O(gate268inter7));
  inv1  gate2949(.a(G779), .O(gate268inter8));
  nand2 gate2950(.a(gate268inter8), .b(gate268inter7), .O(gate268inter9));
  nand2 gate2951(.a(s_343), .b(gate268inter3), .O(gate268inter10));
  nor2  gate2952(.a(gate268inter10), .b(gate268inter9), .O(gate268inter11));
  nor2  gate2953(.a(gate268inter11), .b(gate268inter6), .O(gate268inter12));
  nand2 gate2954(.a(gate268inter12), .b(gate268inter1), .O(G803));
nand2 gate269( .a(G654), .b(G782), .O(G806) );

  xor2  gate2591(.a(G785), .b(G657), .O(gate270inter0));
  nand2 gate2592(.a(gate270inter0), .b(s_292), .O(gate270inter1));
  and2  gate2593(.a(G785), .b(G657), .O(gate270inter2));
  inv1  gate2594(.a(s_292), .O(gate270inter3));
  inv1  gate2595(.a(s_293), .O(gate270inter4));
  nand2 gate2596(.a(gate270inter4), .b(gate270inter3), .O(gate270inter5));
  nor2  gate2597(.a(gate270inter5), .b(gate270inter2), .O(gate270inter6));
  inv1  gate2598(.a(G657), .O(gate270inter7));
  inv1  gate2599(.a(G785), .O(gate270inter8));
  nand2 gate2600(.a(gate270inter8), .b(gate270inter7), .O(gate270inter9));
  nand2 gate2601(.a(s_293), .b(gate270inter3), .O(gate270inter10));
  nor2  gate2602(.a(gate270inter10), .b(gate270inter9), .O(gate270inter11));
  nor2  gate2603(.a(gate270inter11), .b(gate270inter6), .O(gate270inter12));
  nand2 gate2604(.a(gate270inter12), .b(gate270inter1), .O(G809));
nand2 gate271( .a(G660), .b(G788), .O(G812) );
nand2 gate272( .a(G663), .b(G791), .O(G815) );

  xor2  gate575(.a(G794), .b(G642), .O(gate273inter0));
  nand2 gate576(.a(gate273inter0), .b(s_4), .O(gate273inter1));
  and2  gate577(.a(G794), .b(G642), .O(gate273inter2));
  inv1  gate578(.a(s_4), .O(gate273inter3));
  inv1  gate579(.a(s_5), .O(gate273inter4));
  nand2 gate580(.a(gate273inter4), .b(gate273inter3), .O(gate273inter5));
  nor2  gate581(.a(gate273inter5), .b(gate273inter2), .O(gate273inter6));
  inv1  gate582(.a(G642), .O(gate273inter7));
  inv1  gate583(.a(G794), .O(gate273inter8));
  nand2 gate584(.a(gate273inter8), .b(gate273inter7), .O(gate273inter9));
  nand2 gate585(.a(s_5), .b(gate273inter3), .O(gate273inter10));
  nor2  gate586(.a(gate273inter10), .b(gate273inter9), .O(gate273inter11));
  nor2  gate587(.a(gate273inter11), .b(gate273inter6), .O(gate273inter12));
  nand2 gate588(.a(gate273inter12), .b(gate273inter1), .O(G818));
nand2 gate274( .a(G770), .b(G794), .O(G819) );
nand2 gate275( .a(G645), .b(G797), .O(G820) );
nand2 gate276( .a(G773), .b(G797), .O(G821) );

  xor2  gate2059(.a(G800), .b(G648), .O(gate277inter0));
  nand2 gate2060(.a(gate277inter0), .b(s_216), .O(gate277inter1));
  and2  gate2061(.a(G800), .b(G648), .O(gate277inter2));
  inv1  gate2062(.a(s_216), .O(gate277inter3));
  inv1  gate2063(.a(s_217), .O(gate277inter4));
  nand2 gate2064(.a(gate277inter4), .b(gate277inter3), .O(gate277inter5));
  nor2  gate2065(.a(gate277inter5), .b(gate277inter2), .O(gate277inter6));
  inv1  gate2066(.a(G648), .O(gate277inter7));
  inv1  gate2067(.a(G800), .O(gate277inter8));
  nand2 gate2068(.a(gate277inter8), .b(gate277inter7), .O(gate277inter9));
  nand2 gate2069(.a(s_217), .b(gate277inter3), .O(gate277inter10));
  nor2  gate2070(.a(gate277inter10), .b(gate277inter9), .O(gate277inter11));
  nor2  gate2071(.a(gate277inter11), .b(gate277inter6), .O(gate277inter12));
  nand2 gate2072(.a(gate277inter12), .b(gate277inter1), .O(G822));

  xor2  gate2535(.a(G800), .b(G776), .O(gate278inter0));
  nand2 gate2536(.a(gate278inter0), .b(s_284), .O(gate278inter1));
  and2  gate2537(.a(G800), .b(G776), .O(gate278inter2));
  inv1  gate2538(.a(s_284), .O(gate278inter3));
  inv1  gate2539(.a(s_285), .O(gate278inter4));
  nand2 gate2540(.a(gate278inter4), .b(gate278inter3), .O(gate278inter5));
  nor2  gate2541(.a(gate278inter5), .b(gate278inter2), .O(gate278inter6));
  inv1  gate2542(.a(G776), .O(gate278inter7));
  inv1  gate2543(.a(G800), .O(gate278inter8));
  nand2 gate2544(.a(gate278inter8), .b(gate278inter7), .O(gate278inter9));
  nand2 gate2545(.a(s_285), .b(gate278inter3), .O(gate278inter10));
  nor2  gate2546(.a(gate278inter10), .b(gate278inter9), .O(gate278inter11));
  nor2  gate2547(.a(gate278inter11), .b(gate278inter6), .O(gate278inter12));
  nand2 gate2548(.a(gate278inter12), .b(gate278inter1), .O(G823));
nand2 gate279( .a(G651), .b(G803), .O(G824) );

  xor2  gate1919(.a(G803), .b(G779), .O(gate280inter0));
  nand2 gate1920(.a(gate280inter0), .b(s_196), .O(gate280inter1));
  and2  gate1921(.a(G803), .b(G779), .O(gate280inter2));
  inv1  gate1922(.a(s_196), .O(gate280inter3));
  inv1  gate1923(.a(s_197), .O(gate280inter4));
  nand2 gate1924(.a(gate280inter4), .b(gate280inter3), .O(gate280inter5));
  nor2  gate1925(.a(gate280inter5), .b(gate280inter2), .O(gate280inter6));
  inv1  gate1926(.a(G779), .O(gate280inter7));
  inv1  gate1927(.a(G803), .O(gate280inter8));
  nand2 gate1928(.a(gate280inter8), .b(gate280inter7), .O(gate280inter9));
  nand2 gate1929(.a(s_197), .b(gate280inter3), .O(gate280inter10));
  nor2  gate1930(.a(gate280inter10), .b(gate280inter9), .O(gate280inter11));
  nor2  gate1931(.a(gate280inter11), .b(gate280inter6), .O(gate280inter12));
  nand2 gate1932(.a(gate280inter12), .b(gate280inter1), .O(G825));

  xor2  gate729(.a(G806), .b(G654), .O(gate281inter0));
  nand2 gate730(.a(gate281inter0), .b(s_26), .O(gate281inter1));
  and2  gate731(.a(G806), .b(G654), .O(gate281inter2));
  inv1  gate732(.a(s_26), .O(gate281inter3));
  inv1  gate733(.a(s_27), .O(gate281inter4));
  nand2 gate734(.a(gate281inter4), .b(gate281inter3), .O(gate281inter5));
  nor2  gate735(.a(gate281inter5), .b(gate281inter2), .O(gate281inter6));
  inv1  gate736(.a(G654), .O(gate281inter7));
  inv1  gate737(.a(G806), .O(gate281inter8));
  nand2 gate738(.a(gate281inter8), .b(gate281inter7), .O(gate281inter9));
  nand2 gate739(.a(s_27), .b(gate281inter3), .O(gate281inter10));
  nor2  gate740(.a(gate281inter10), .b(gate281inter9), .O(gate281inter11));
  nor2  gate741(.a(gate281inter11), .b(gate281inter6), .O(gate281inter12));
  nand2 gate742(.a(gate281inter12), .b(gate281inter1), .O(G826));
nand2 gate282( .a(G782), .b(G806), .O(G827) );
nand2 gate283( .a(G657), .b(G809), .O(G828) );
nand2 gate284( .a(G785), .b(G809), .O(G829) );
nand2 gate285( .a(G660), .b(G812), .O(G830) );

  xor2  gate2409(.a(G812), .b(G788), .O(gate286inter0));
  nand2 gate2410(.a(gate286inter0), .b(s_266), .O(gate286inter1));
  and2  gate2411(.a(G812), .b(G788), .O(gate286inter2));
  inv1  gate2412(.a(s_266), .O(gate286inter3));
  inv1  gate2413(.a(s_267), .O(gate286inter4));
  nand2 gate2414(.a(gate286inter4), .b(gate286inter3), .O(gate286inter5));
  nor2  gate2415(.a(gate286inter5), .b(gate286inter2), .O(gate286inter6));
  inv1  gate2416(.a(G788), .O(gate286inter7));
  inv1  gate2417(.a(G812), .O(gate286inter8));
  nand2 gate2418(.a(gate286inter8), .b(gate286inter7), .O(gate286inter9));
  nand2 gate2419(.a(s_267), .b(gate286inter3), .O(gate286inter10));
  nor2  gate2420(.a(gate286inter10), .b(gate286inter9), .O(gate286inter11));
  nor2  gate2421(.a(gate286inter11), .b(gate286inter6), .O(gate286inter12));
  nand2 gate2422(.a(gate286inter12), .b(gate286inter1), .O(G831));
nand2 gate287( .a(G663), .b(G815), .O(G832) );

  xor2  gate1331(.a(G815), .b(G791), .O(gate288inter0));
  nand2 gate1332(.a(gate288inter0), .b(s_112), .O(gate288inter1));
  and2  gate1333(.a(G815), .b(G791), .O(gate288inter2));
  inv1  gate1334(.a(s_112), .O(gate288inter3));
  inv1  gate1335(.a(s_113), .O(gate288inter4));
  nand2 gate1336(.a(gate288inter4), .b(gate288inter3), .O(gate288inter5));
  nor2  gate1337(.a(gate288inter5), .b(gate288inter2), .O(gate288inter6));
  inv1  gate1338(.a(G791), .O(gate288inter7));
  inv1  gate1339(.a(G815), .O(gate288inter8));
  nand2 gate1340(.a(gate288inter8), .b(gate288inter7), .O(gate288inter9));
  nand2 gate1341(.a(s_113), .b(gate288inter3), .O(gate288inter10));
  nor2  gate1342(.a(gate288inter10), .b(gate288inter9), .O(gate288inter11));
  nor2  gate1343(.a(gate288inter11), .b(gate288inter6), .O(gate288inter12));
  nand2 gate1344(.a(gate288inter12), .b(gate288inter1), .O(G833));
nand2 gate289( .a(G818), .b(G819), .O(G834) );

  xor2  gate2843(.a(G821), .b(G820), .O(gate290inter0));
  nand2 gate2844(.a(gate290inter0), .b(s_328), .O(gate290inter1));
  and2  gate2845(.a(G821), .b(G820), .O(gate290inter2));
  inv1  gate2846(.a(s_328), .O(gate290inter3));
  inv1  gate2847(.a(s_329), .O(gate290inter4));
  nand2 gate2848(.a(gate290inter4), .b(gate290inter3), .O(gate290inter5));
  nor2  gate2849(.a(gate290inter5), .b(gate290inter2), .O(gate290inter6));
  inv1  gate2850(.a(G820), .O(gate290inter7));
  inv1  gate2851(.a(G821), .O(gate290inter8));
  nand2 gate2852(.a(gate290inter8), .b(gate290inter7), .O(gate290inter9));
  nand2 gate2853(.a(s_329), .b(gate290inter3), .O(gate290inter10));
  nor2  gate2854(.a(gate290inter10), .b(gate290inter9), .O(gate290inter11));
  nor2  gate2855(.a(gate290inter11), .b(gate290inter6), .O(gate290inter12));
  nand2 gate2856(.a(gate290inter12), .b(gate290inter1), .O(G847));
nand2 gate291( .a(G822), .b(G823), .O(G860) );

  xor2  gate1233(.a(G825), .b(G824), .O(gate292inter0));
  nand2 gate1234(.a(gate292inter0), .b(s_98), .O(gate292inter1));
  and2  gate1235(.a(G825), .b(G824), .O(gate292inter2));
  inv1  gate1236(.a(s_98), .O(gate292inter3));
  inv1  gate1237(.a(s_99), .O(gate292inter4));
  nand2 gate1238(.a(gate292inter4), .b(gate292inter3), .O(gate292inter5));
  nor2  gate1239(.a(gate292inter5), .b(gate292inter2), .O(gate292inter6));
  inv1  gate1240(.a(G824), .O(gate292inter7));
  inv1  gate1241(.a(G825), .O(gate292inter8));
  nand2 gate1242(.a(gate292inter8), .b(gate292inter7), .O(gate292inter9));
  nand2 gate1243(.a(s_99), .b(gate292inter3), .O(gate292inter10));
  nor2  gate1244(.a(gate292inter10), .b(gate292inter9), .O(gate292inter11));
  nor2  gate1245(.a(gate292inter11), .b(gate292inter6), .O(gate292inter12));
  nand2 gate1246(.a(gate292inter12), .b(gate292inter1), .O(G873));

  xor2  gate1541(.a(G829), .b(G828), .O(gate293inter0));
  nand2 gate1542(.a(gate293inter0), .b(s_142), .O(gate293inter1));
  and2  gate1543(.a(G829), .b(G828), .O(gate293inter2));
  inv1  gate1544(.a(s_142), .O(gate293inter3));
  inv1  gate1545(.a(s_143), .O(gate293inter4));
  nand2 gate1546(.a(gate293inter4), .b(gate293inter3), .O(gate293inter5));
  nor2  gate1547(.a(gate293inter5), .b(gate293inter2), .O(gate293inter6));
  inv1  gate1548(.a(G828), .O(gate293inter7));
  inv1  gate1549(.a(G829), .O(gate293inter8));
  nand2 gate1550(.a(gate293inter8), .b(gate293inter7), .O(gate293inter9));
  nand2 gate1551(.a(s_143), .b(gate293inter3), .O(gate293inter10));
  nor2  gate1552(.a(gate293inter10), .b(gate293inter9), .O(gate293inter11));
  nor2  gate1553(.a(gate293inter11), .b(gate293inter6), .O(gate293inter12));
  nand2 gate1554(.a(gate293inter12), .b(gate293inter1), .O(G886));
nand2 gate294( .a(G832), .b(G833), .O(G899) );

  xor2  gate1219(.a(G831), .b(G830), .O(gate295inter0));
  nand2 gate1220(.a(gate295inter0), .b(s_96), .O(gate295inter1));
  and2  gate1221(.a(G831), .b(G830), .O(gate295inter2));
  inv1  gate1222(.a(s_96), .O(gate295inter3));
  inv1  gate1223(.a(s_97), .O(gate295inter4));
  nand2 gate1224(.a(gate295inter4), .b(gate295inter3), .O(gate295inter5));
  nor2  gate1225(.a(gate295inter5), .b(gate295inter2), .O(gate295inter6));
  inv1  gate1226(.a(G830), .O(gate295inter7));
  inv1  gate1227(.a(G831), .O(gate295inter8));
  nand2 gate1228(.a(gate295inter8), .b(gate295inter7), .O(gate295inter9));
  nand2 gate1229(.a(s_97), .b(gate295inter3), .O(gate295inter10));
  nor2  gate1230(.a(gate295inter10), .b(gate295inter9), .O(gate295inter11));
  nor2  gate1231(.a(gate295inter11), .b(gate295inter6), .O(gate295inter12));
  nand2 gate1232(.a(gate295inter12), .b(gate295inter1), .O(G912));

  xor2  gate995(.a(G827), .b(G826), .O(gate296inter0));
  nand2 gate996(.a(gate296inter0), .b(s_64), .O(gate296inter1));
  and2  gate997(.a(G827), .b(G826), .O(gate296inter2));
  inv1  gate998(.a(s_64), .O(gate296inter3));
  inv1  gate999(.a(s_65), .O(gate296inter4));
  nand2 gate1000(.a(gate296inter4), .b(gate296inter3), .O(gate296inter5));
  nor2  gate1001(.a(gate296inter5), .b(gate296inter2), .O(gate296inter6));
  inv1  gate1002(.a(G826), .O(gate296inter7));
  inv1  gate1003(.a(G827), .O(gate296inter8));
  nand2 gate1004(.a(gate296inter8), .b(gate296inter7), .O(gate296inter9));
  nand2 gate1005(.a(s_65), .b(gate296inter3), .O(gate296inter10));
  nor2  gate1006(.a(gate296inter10), .b(gate296inter9), .O(gate296inter11));
  nor2  gate1007(.a(gate296inter11), .b(gate296inter6), .O(gate296inter12));
  nand2 gate1008(.a(gate296inter12), .b(gate296inter1), .O(G925));
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );
nand2 gate387( .a(G1), .b(G1036), .O(G1132) );
nand2 gate388( .a(G2), .b(G1039), .O(G1135) );

  xor2  gate1751(.a(G1042), .b(G3), .O(gate389inter0));
  nand2 gate1752(.a(gate389inter0), .b(s_172), .O(gate389inter1));
  and2  gate1753(.a(G1042), .b(G3), .O(gate389inter2));
  inv1  gate1754(.a(s_172), .O(gate389inter3));
  inv1  gate1755(.a(s_173), .O(gate389inter4));
  nand2 gate1756(.a(gate389inter4), .b(gate389inter3), .O(gate389inter5));
  nor2  gate1757(.a(gate389inter5), .b(gate389inter2), .O(gate389inter6));
  inv1  gate1758(.a(G3), .O(gate389inter7));
  inv1  gate1759(.a(G1042), .O(gate389inter8));
  nand2 gate1760(.a(gate389inter8), .b(gate389inter7), .O(gate389inter9));
  nand2 gate1761(.a(s_173), .b(gate389inter3), .O(gate389inter10));
  nor2  gate1762(.a(gate389inter10), .b(gate389inter9), .O(gate389inter11));
  nor2  gate1763(.a(gate389inter11), .b(gate389inter6), .O(gate389inter12));
  nand2 gate1764(.a(gate389inter12), .b(gate389inter1), .O(G1138));
nand2 gate390( .a(G4), .b(G1045), .O(G1141) );
nand2 gate391( .a(G5), .b(G1048), .O(G1144) );

  xor2  gate1555(.a(G1051), .b(G6), .O(gate392inter0));
  nand2 gate1556(.a(gate392inter0), .b(s_144), .O(gate392inter1));
  and2  gate1557(.a(G1051), .b(G6), .O(gate392inter2));
  inv1  gate1558(.a(s_144), .O(gate392inter3));
  inv1  gate1559(.a(s_145), .O(gate392inter4));
  nand2 gate1560(.a(gate392inter4), .b(gate392inter3), .O(gate392inter5));
  nor2  gate1561(.a(gate392inter5), .b(gate392inter2), .O(gate392inter6));
  inv1  gate1562(.a(G6), .O(gate392inter7));
  inv1  gate1563(.a(G1051), .O(gate392inter8));
  nand2 gate1564(.a(gate392inter8), .b(gate392inter7), .O(gate392inter9));
  nand2 gate1565(.a(s_145), .b(gate392inter3), .O(gate392inter10));
  nor2  gate1566(.a(gate392inter10), .b(gate392inter9), .O(gate392inter11));
  nor2  gate1567(.a(gate392inter11), .b(gate392inter6), .O(gate392inter12));
  nand2 gate1568(.a(gate392inter12), .b(gate392inter1), .O(G1147));

  xor2  gate2801(.a(G1054), .b(G7), .O(gate393inter0));
  nand2 gate2802(.a(gate393inter0), .b(s_322), .O(gate393inter1));
  and2  gate2803(.a(G1054), .b(G7), .O(gate393inter2));
  inv1  gate2804(.a(s_322), .O(gate393inter3));
  inv1  gate2805(.a(s_323), .O(gate393inter4));
  nand2 gate2806(.a(gate393inter4), .b(gate393inter3), .O(gate393inter5));
  nor2  gate2807(.a(gate393inter5), .b(gate393inter2), .O(gate393inter6));
  inv1  gate2808(.a(G7), .O(gate393inter7));
  inv1  gate2809(.a(G1054), .O(gate393inter8));
  nand2 gate2810(.a(gate393inter8), .b(gate393inter7), .O(gate393inter9));
  nand2 gate2811(.a(s_323), .b(gate393inter3), .O(gate393inter10));
  nor2  gate2812(.a(gate393inter10), .b(gate393inter9), .O(gate393inter11));
  nor2  gate2813(.a(gate393inter11), .b(gate393inter6), .O(gate393inter12));
  nand2 gate2814(.a(gate393inter12), .b(gate393inter1), .O(G1150));

  xor2  gate1709(.a(G1057), .b(G8), .O(gate394inter0));
  nand2 gate1710(.a(gate394inter0), .b(s_166), .O(gate394inter1));
  and2  gate1711(.a(G1057), .b(G8), .O(gate394inter2));
  inv1  gate1712(.a(s_166), .O(gate394inter3));
  inv1  gate1713(.a(s_167), .O(gate394inter4));
  nand2 gate1714(.a(gate394inter4), .b(gate394inter3), .O(gate394inter5));
  nor2  gate1715(.a(gate394inter5), .b(gate394inter2), .O(gate394inter6));
  inv1  gate1716(.a(G8), .O(gate394inter7));
  inv1  gate1717(.a(G1057), .O(gate394inter8));
  nand2 gate1718(.a(gate394inter8), .b(gate394inter7), .O(gate394inter9));
  nand2 gate1719(.a(s_167), .b(gate394inter3), .O(gate394inter10));
  nor2  gate1720(.a(gate394inter10), .b(gate394inter9), .O(gate394inter11));
  nor2  gate1721(.a(gate394inter11), .b(gate394inter6), .O(gate394inter12));
  nand2 gate1722(.a(gate394inter12), .b(gate394inter1), .O(G1153));
nand2 gate395( .a(G9), .b(G1060), .O(G1156) );

  xor2  gate2115(.a(G1063), .b(G10), .O(gate396inter0));
  nand2 gate2116(.a(gate396inter0), .b(s_224), .O(gate396inter1));
  and2  gate2117(.a(G1063), .b(G10), .O(gate396inter2));
  inv1  gate2118(.a(s_224), .O(gate396inter3));
  inv1  gate2119(.a(s_225), .O(gate396inter4));
  nand2 gate2120(.a(gate396inter4), .b(gate396inter3), .O(gate396inter5));
  nor2  gate2121(.a(gate396inter5), .b(gate396inter2), .O(gate396inter6));
  inv1  gate2122(.a(G10), .O(gate396inter7));
  inv1  gate2123(.a(G1063), .O(gate396inter8));
  nand2 gate2124(.a(gate396inter8), .b(gate396inter7), .O(gate396inter9));
  nand2 gate2125(.a(s_225), .b(gate396inter3), .O(gate396inter10));
  nor2  gate2126(.a(gate396inter10), .b(gate396inter9), .O(gate396inter11));
  nor2  gate2127(.a(gate396inter11), .b(gate396inter6), .O(gate396inter12));
  nand2 gate2128(.a(gate396inter12), .b(gate396inter1), .O(G1159));
nand2 gate397( .a(G11), .b(G1066), .O(G1162) );
nand2 gate398( .a(G12), .b(G1069), .O(G1165) );
nand2 gate399( .a(G13), .b(G1072), .O(G1168) );
nand2 gate400( .a(G14), .b(G1075), .O(G1171) );
nand2 gate401( .a(G15), .b(G1078), .O(G1174) );
nand2 gate402( .a(G16), .b(G1081), .O(G1177) );
nand2 gate403( .a(G17), .b(G1084), .O(G1180) );
nand2 gate404( .a(G18), .b(G1087), .O(G1183) );

  xor2  gate1611(.a(G1090), .b(G19), .O(gate405inter0));
  nand2 gate1612(.a(gate405inter0), .b(s_152), .O(gate405inter1));
  and2  gate1613(.a(G1090), .b(G19), .O(gate405inter2));
  inv1  gate1614(.a(s_152), .O(gate405inter3));
  inv1  gate1615(.a(s_153), .O(gate405inter4));
  nand2 gate1616(.a(gate405inter4), .b(gate405inter3), .O(gate405inter5));
  nor2  gate1617(.a(gate405inter5), .b(gate405inter2), .O(gate405inter6));
  inv1  gate1618(.a(G19), .O(gate405inter7));
  inv1  gate1619(.a(G1090), .O(gate405inter8));
  nand2 gate1620(.a(gate405inter8), .b(gate405inter7), .O(gate405inter9));
  nand2 gate1621(.a(s_153), .b(gate405inter3), .O(gate405inter10));
  nor2  gate1622(.a(gate405inter10), .b(gate405inter9), .O(gate405inter11));
  nor2  gate1623(.a(gate405inter11), .b(gate405inter6), .O(gate405inter12));
  nand2 gate1624(.a(gate405inter12), .b(gate405inter1), .O(G1186));
nand2 gate406( .a(G20), .b(G1093), .O(G1189) );
nand2 gate407( .a(G21), .b(G1096), .O(G1192) );
nand2 gate408( .a(G22), .b(G1099), .O(G1195) );

  xor2  gate1961(.a(G1102), .b(G23), .O(gate409inter0));
  nand2 gate1962(.a(gate409inter0), .b(s_202), .O(gate409inter1));
  and2  gate1963(.a(G1102), .b(G23), .O(gate409inter2));
  inv1  gate1964(.a(s_202), .O(gate409inter3));
  inv1  gate1965(.a(s_203), .O(gate409inter4));
  nand2 gate1966(.a(gate409inter4), .b(gate409inter3), .O(gate409inter5));
  nor2  gate1967(.a(gate409inter5), .b(gate409inter2), .O(gate409inter6));
  inv1  gate1968(.a(G23), .O(gate409inter7));
  inv1  gate1969(.a(G1102), .O(gate409inter8));
  nand2 gate1970(.a(gate409inter8), .b(gate409inter7), .O(gate409inter9));
  nand2 gate1971(.a(s_203), .b(gate409inter3), .O(gate409inter10));
  nor2  gate1972(.a(gate409inter10), .b(gate409inter9), .O(gate409inter11));
  nor2  gate1973(.a(gate409inter11), .b(gate409inter6), .O(gate409inter12));
  nand2 gate1974(.a(gate409inter12), .b(gate409inter1), .O(G1198));

  xor2  gate2017(.a(G1105), .b(G24), .O(gate410inter0));
  nand2 gate2018(.a(gate410inter0), .b(s_210), .O(gate410inter1));
  and2  gate2019(.a(G1105), .b(G24), .O(gate410inter2));
  inv1  gate2020(.a(s_210), .O(gate410inter3));
  inv1  gate2021(.a(s_211), .O(gate410inter4));
  nand2 gate2022(.a(gate410inter4), .b(gate410inter3), .O(gate410inter5));
  nor2  gate2023(.a(gate410inter5), .b(gate410inter2), .O(gate410inter6));
  inv1  gate2024(.a(G24), .O(gate410inter7));
  inv1  gate2025(.a(G1105), .O(gate410inter8));
  nand2 gate2026(.a(gate410inter8), .b(gate410inter7), .O(gate410inter9));
  nand2 gate2027(.a(s_211), .b(gate410inter3), .O(gate410inter10));
  nor2  gate2028(.a(gate410inter10), .b(gate410inter9), .O(gate410inter11));
  nor2  gate2029(.a(gate410inter11), .b(gate410inter6), .O(gate410inter12));
  nand2 gate2030(.a(gate410inter12), .b(gate410inter1), .O(G1201));
nand2 gate411( .a(G25), .b(G1108), .O(G1204) );

  xor2  gate2143(.a(G1111), .b(G26), .O(gate412inter0));
  nand2 gate2144(.a(gate412inter0), .b(s_228), .O(gate412inter1));
  and2  gate2145(.a(G1111), .b(G26), .O(gate412inter2));
  inv1  gate2146(.a(s_228), .O(gate412inter3));
  inv1  gate2147(.a(s_229), .O(gate412inter4));
  nand2 gate2148(.a(gate412inter4), .b(gate412inter3), .O(gate412inter5));
  nor2  gate2149(.a(gate412inter5), .b(gate412inter2), .O(gate412inter6));
  inv1  gate2150(.a(G26), .O(gate412inter7));
  inv1  gate2151(.a(G1111), .O(gate412inter8));
  nand2 gate2152(.a(gate412inter8), .b(gate412inter7), .O(gate412inter9));
  nand2 gate2153(.a(s_229), .b(gate412inter3), .O(gate412inter10));
  nor2  gate2154(.a(gate412inter10), .b(gate412inter9), .O(gate412inter11));
  nor2  gate2155(.a(gate412inter11), .b(gate412inter6), .O(gate412inter12));
  nand2 gate2156(.a(gate412inter12), .b(gate412inter1), .O(G1207));

  xor2  gate1247(.a(G1114), .b(G27), .O(gate413inter0));
  nand2 gate1248(.a(gate413inter0), .b(s_100), .O(gate413inter1));
  and2  gate1249(.a(G1114), .b(G27), .O(gate413inter2));
  inv1  gate1250(.a(s_100), .O(gate413inter3));
  inv1  gate1251(.a(s_101), .O(gate413inter4));
  nand2 gate1252(.a(gate413inter4), .b(gate413inter3), .O(gate413inter5));
  nor2  gate1253(.a(gate413inter5), .b(gate413inter2), .O(gate413inter6));
  inv1  gate1254(.a(G27), .O(gate413inter7));
  inv1  gate1255(.a(G1114), .O(gate413inter8));
  nand2 gate1256(.a(gate413inter8), .b(gate413inter7), .O(gate413inter9));
  nand2 gate1257(.a(s_101), .b(gate413inter3), .O(gate413inter10));
  nor2  gate1258(.a(gate413inter10), .b(gate413inter9), .O(gate413inter11));
  nor2  gate1259(.a(gate413inter11), .b(gate413inter6), .O(gate413inter12));
  nand2 gate1260(.a(gate413inter12), .b(gate413inter1), .O(G1210));
nand2 gate414( .a(G28), .b(G1117), .O(G1213) );

  xor2  gate2549(.a(G1120), .b(G29), .O(gate415inter0));
  nand2 gate2550(.a(gate415inter0), .b(s_286), .O(gate415inter1));
  and2  gate2551(.a(G1120), .b(G29), .O(gate415inter2));
  inv1  gate2552(.a(s_286), .O(gate415inter3));
  inv1  gate2553(.a(s_287), .O(gate415inter4));
  nand2 gate2554(.a(gate415inter4), .b(gate415inter3), .O(gate415inter5));
  nor2  gate2555(.a(gate415inter5), .b(gate415inter2), .O(gate415inter6));
  inv1  gate2556(.a(G29), .O(gate415inter7));
  inv1  gate2557(.a(G1120), .O(gate415inter8));
  nand2 gate2558(.a(gate415inter8), .b(gate415inter7), .O(gate415inter9));
  nand2 gate2559(.a(s_287), .b(gate415inter3), .O(gate415inter10));
  nor2  gate2560(.a(gate415inter10), .b(gate415inter9), .O(gate415inter11));
  nor2  gate2561(.a(gate415inter11), .b(gate415inter6), .O(gate415inter12));
  nand2 gate2562(.a(gate415inter12), .b(gate415inter1), .O(G1216));

  xor2  gate2465(.a(G1123), .b(G30), .O(gate416inter0));
  nand2 gate2466(.a(gate416inter0), .b(s_274), .O(gate416inter1));
  and2  gate2467(.a(G1123), .b(G30), .O(gate416inter2));
  inv1  gate2468(.a(s_274), .O(gate416inter3));
  inv1  gate2469(.a(s_275), .O(gate416inter4));
  nand2 gate2470(.a(gate416inter4), .b(gate416inter3), .O(gate416inter5));
  nor2  gate2471(.a(gate416inter5), .b(gate416inter2), .O(gate416inter6));
  inv1  gate2472(.a(G30), .O(gate416inter7));
  inv1  gate2473(.a(G1123), .O(gate416inter8));
  nand2 gate2474(.a(gate416inter8), .b(gate416inter7), .O(gate416inter9));
  nand2 gate2475(.a(s_275), .b(gate416inter3), .O(gate416inter10));
  nor2  gate2476(.a(gate416inter10), .b(gate416inter9), .O(gate416inter11));
  nor2  gate2477(.a(gate416inter11), .b(gate416inter6), .O(gate416inter12));
  nand2 gate2478(.a(gate416inter12), .b(gate416inter1), .O(G1219));
nand2 gate417( .a(G31), .b(G1126), .O(G1222) );
nand2 gate418( .a(G32), .b(G1129), .O(G1225) );
nand2 gate419( .a(G1), .b(G1132), .O(G1228) );
nand2 gate420( .a(G1036), .b(G1132), .O(G1229) );

  xor2  gate1583(.a(G1135), .b(G2), .O(gate421inter0));
  nand2 gate1584(.a(gate421inter0), .b(s_148), .O(gate421inter1));
  and2  gate1585(.a(G1135), .b(G2), .O(gate421inter2));
  inv1  gate1586(.a(s_148), .O(gate421inter3));
  inv1  gate1587(.a(s_149), .O(gate421inter4));
  nand2 gate1588(.a(gate421inter4), .b(gate421inter3), .O(gate421inter5));
  nor2  gate1589(.a(gate421inter5), .b(gate421inter2), .O(gate421inter6));
  inv1  gate1590(.a(G2), .O(gate421inter7));
  inv1  gate1591(.a(G1135), .O(gate421inter8));
  nand2 gate1592(.a(gate421inter8), .b(gate421inter7), .O(gate421inter9));
  nand2 gate1593(.a(s_149), .b(gate421inter3), .O(gate421inter10));
  nor2  gate1594(.a(gate421inter10), .b(gate421inter9), .O(gate421inter11));
  nor2  gate1595(.a(gate421inter11), .b(gate421inter6), .O(gate421inter12));
  nand2 gate1596(.a(gate421inter12), .b(gate421inter1), .O(G1230));
nand2 gate422( .a(G1039), .b(G1135), .O(G1231) );
nand2 gate423( .a(G3), .b(G1138), .O(G1232) );
nand2 gate424( .a(G1042), .b(G1138), .O(G1233) );

  xor2  gate2451(.a(G1141), .b(G4), .O(gate425inter0));
  nand2 gate2452(.a(gate425inter0), .b(s_272), .O(gate425inter1));
  and2  gate2453(.a(G1141), .b(G4), .O(gate425inter2));
  inv1  gate2454(.a(s_272), .O(gate425inter3));
  inv1  gate2455(.a(s_273), .O(gate425inter4));
  nand2 gate2456(.a(gate425inter4), .b(gate425inter3), .O(gate425inter5));
  nor2  gate2457(.a(gate425inter5), .b(gate425inter2), .O(gate425inter6));
  inv1  gate2458(.a(G4), .O(gate425inter7));
  inv1  gate2459(.a(G1141), .O(gate425inter8));
  nand2 gate2460(.a(gate425inter8), .b(gate425inter7), .O(gate425inter9));
  nand2 gate2461(.a(s_273), .b(gate425inter3), .O(gate425inter10));
  nor2  gate2462(.a(gate425inter10), .b(gate425inter9), .O(gate425inter11));
  nor2  gate2463(.a(gate425inter11), .b(gate425inter6), .O(gate425inter12));
  nand2 gate2464(.a(gate425inter12), .b(gate425inter1), .O(G1234));

  xor2  gate2423(.a(G1141), .b(G1045), .O(gate426inter0));
  nand2 gate2424(.a(gate426inter0), .b(s_268), .O(gate426inter1));
  and2  gate2425(.a(G1141), .b(G1045), .O(gate426inter2));
  inv1  gate2426(.a(s_268), .O(gate426inter3));
  inv1  gate2427(.a(s_269), .O(gate426inter4));
  nand2 gate2428(.a(gate426inter4), .b(gate426inter3), .O(gate426inter5));
  nor2  gate2429(.a(gate426inter5), .b(gate426inter2), .O(gate426inter6));
  inv1  gate2430(.a(G1045), .O(gate426inter7));
  inv1  gate2431(.a(G1141), .O(gate426inter8));
  nand2 gate2432(.a(gate426inter8), .b(gate426inter7), .O(gate426inter9));
  nand2 gate2433(.a(s_269), .b(gate426inter3), .O(gate426inter10));
  nor2  gate2434(.a(gate426inter10), .b(gate426inter9), .O(gate426inter11));
  nor2  gate2435(.a(gate426inter11), .b(gate426inter6), .O(gate426inter12));
  nand2 gate2436(.a(gate426inter12), .b(gate426inter1), .O(G1235));

  xor2  gate2157(.a(G1144), .b(G5), .O(gate427inter0));
  nand2 gate2158(.a(gate427inter0), .b(s_230), .O(gate427inter1));
  and2  gate2159(.a(G1144), .b(G5), .O(gate427inter2));
  inv1  gate2160(.a(s_230), .O(gate427inter3));
  inv1  gate2161(.a(s_231), .O(gate427inter4));
  nand2 gate2162(.a(gate427inter4), .b(gate427inter3), .O(gate427inter5));
  nor2  gate2163(.a(gate427inter5), .b(gate427inter2), .O(gate427inter6));
  inv1  gate2164(.a(G5), .O(gate427inter7));
  inv1  gate2165(.a(G1144), .O(gate427inter8));
  nand2 gate2166(.a(gate427inter8), .b(gate427inter7), .O(gate427inter9));
  nand2 gate2167(.a(s_231), .b(gate427inter3), .O(gate427inter10));
  nor2  gate2168(.a(gate427inter10), .b(gate427inter9), .O(gate427inter11));
  nor2  gate2169(.a(gate427inter11), .b(gate427inter6), .O(gate427inter12));
  nand2 gate2170(.a(gate427inter12), .b(gate427inter1), .O(G1236));

  xor2  gate1261(.a(G1144), .b(G1048), .O(gate428inter0));
  nand2 gate1262(.a(gate428inter0), .b(s_102), .O(gate428inter1));
  and2  gate1263(.a(G1144), .b(G1048), .O(gate428inter2));
  inv1  gate1264(.a(s_102), .O(gate428inter3));
  inv1  gate1265(.a(s_103), .O(gate428inter4));
  nand2 gate1266(.a(gate428inter4), .b(gate428inter3), .O(gate428inter5));
  nor2  gate1267(.a(gate428inter5), .b(gate428inter2), .O(gate428inter6));
  inv1  gate1268(.a(G1048), .O(gate428inter7));
  inv1  gate1269(.a(G1144), .O(gate428inter8));
  nand2 gate1270(.a(gate428inter8), .b(gate428inter7), .O(gate428inter9));
  nand2 gate1271(.a(s_103), .b(gate428inter3), .O(gate428inter10));
  nor2  gate1272(.a(gate428inter10), .b(gate428inter9), .O(gate428inter11));
  nor2  gate1273(.a(gate428inter11), .b(gate428inter6), .O(gate428inter12));
  nand2 gate1274(.a(gate428inter12), .b(gate428inter1), .O(G1237));
nand2 gate429( .a(G6), .b(G1147), .O(G1238) );
nand2 gate430( .a(G1051), .b(G1147), .O(G1239) );
nand2 gate431( .a(G7), .b(G1150), .O(G1240) );
nand2 gate432( .a(G1054), .b(G1150), .O(G1241) );

  xor2  gate645(.a(G1153), .b(G8), .O(gate433inter0));
  nand2 gate646(.a(gate433inter0), .b(s_14), .O(gate433inter1));
  and2  gate647(.a(G1153), .b(G8), .O(gate433inter2));
  inv1  gate648(.a(s_14), .O(gate433inter3));
  inv1  gate649(.a(s_15), .O(gate433inter4));
  nand2 gate650(.a(gate433inter4), .b(gate433inter3), .O(gate433inter5));
  nor2  gate651(.a(gate433inter5), .b(gate433inter2), .O(gate433inter6));
  inv1  gate652(.a(G8), .O(gate433inter7));
  inv1  gate653(.a(G1153), .O(gate433inter8));
  nand2 gate654(.a(gate433inter8), .b(gate433inter7), .O(gate433inter9));
  nand2 gate655(.a(s_15), .b(gate433inter3), .O(gate433inter10));
  nor2  gate656(.a(gate433inter10), .b(gate433inter9), .O(gate433inter11));
  nor2  gate657(.a(gate433inter11), .b(gate433inter6), .O(gate433inter12));
  nand2 gate658(.a(gate433inter12), .b(gate433inter1), .O(G1242));
nand2 gate434( .a(G1057), .b(G1153), .O(G1243) );
nand2 gate435( .a(G9), .b(G1156), .O(G1244) );
nand2 gate436( .a(G1060), .b(G1156), .O(G1245) );
nand2 gate437( .a(G10), .b(G1159), .O(G1246) );

  xor2  gate2619(.a(G1159), .b(G1063), .O(gate438inter0));
  nand2 gate2620(.a(gate438inter0), .b(s_296), .O(gate438inter1));
  and2  gate2621(.a(G1159), .b(G1063), .O(gate438inter2));
  inv1  gate2622(.a(s_296), .O(gate438inter3));
  inv1  gate2623(.a(s_297), .O(gate438inter4));
  nand2 gate2624(.a(gate438inter4), .b(gate438inter3), .O(gate438inter5));
  nor2  gate2625(.a(gate438inter5), .b(gate438inter2), .O(gate438inter6));
  inv1  gate2626(.a(G1063), .O(gate438inter7));
  inv1  gate2627(.a(G1159), .O(gate438inter8));
  nand2 gate2628(.a(gate438inter8), .b(gate438inter7), .O(gate438inter9));
  nand2 gate2629(.a(s_297), .b(gate438inter3), .O(gate438inter10));
  nor2  gate2630(.a(gate438inter10), .b(gate438inter9), .O(gate438inter11));
  nor2  gate2631(.a(gate438inter11), .b(gate438inter6), .O(gate438inter12));
  nand2 gate2632(.a(gate438inter12), .b(gate438inter1), .O(G1247));

  xor2  gate1905(.a(G1162), .b(G11), .O(gate439inter0));
  nand2 gate1906(.a(gate439inter0), .b(s_194), .O(gate439inter1));
  and2  gate1907(.a(G1162), .b(G11), .O(gate439inter2));
  inv1  gate1908(.a(s_194), .O(gate439inter3));
  inv1  gate1909(.a(s_195), .O(gate439inter4));
  nand2 gate1910(.a(gate439inter4), .b(gate439inter3), .O(gate439inter5));
  nor2  gate1911(.a(gate439inter5), .b(gate439inter2), .O(gate439inter6));
  inv1  gate1912(.a(G11), .O(gate439inter7));
  inv1  gate1913(.a(G1162), .O(gate439inter8));
  nand2 gate1914(.a(gate439inter8), .b(gate439inter7), .O(gate439inter9));
  nand2 gate1915(.a(s_195), .b(gate439inter3), .O(gate439inter10));
  nor2  gate1916(.a(gate439inter10), .b(gate439inter9), .O(gate439inter11));
  nor2  gate1917(.a(gate439inter11), .b(gate439inter6), .O(gate439inter12));
  nand2 gate1918(.a(gate439inter12), .b(gate439inter1), .O(G1248));
nand2 gate440( .a(G1066), .b(G1162), .O(G1249) );
nand2 gate441( .a(G12), .b(G1165), .O(G1250) );
nand2 gate442( .a(G1069), .b(G1165), .O(G1251) );

  xor2  gate2395(.a(G1168), .b(G13), .O(gate443inter0));
  nand2 gate2396(.a(gate443inter0), .b(s_264), .O(gate443inter1));
  and2  gate2397(.a(G1168), .b(G13), .O(gate443inter2));
  inv1  gate2398(.a(s_264), .O(gate443inter3));
  inv1  gate2399(.a(s_265), .O(gate443inter4));
  nand2 gate2400(.a(gate443inter4), .b(gate443inter3), .O(gate443inter5));
  nor2  gate2401(.a(gate443inter5), .b(gate443inter2), .O(gate443inter6));
  inv1  gate2402(.a(G13), .O(gate443inter7));
  inv1  gate2403(.a(G1168), .O(gate443inter8));
  nand2 gate2404(.a(gate443inter8), .b(gate443inter7), .O(gate443inter9));
  nand2 gate2405(.a(s_265), .b(gate443inter3), .O(gate443inter10));
  nor2  gate2406(.a(gate443inter10), .b(gate443inter9), .O(gate443inter11));
  nor2  gate2407(.a(gate443inter11), .b(gate443inter6), .O(gate443inter12));
  nand2 gate2408(.a(gate443inter12), .b(gate443inter1), .O(G1252));
nand2 gate444( .a(G1072), .b(G1168), .O(G1253) );

  xor2  gate547(.a(G1171), .b(G14), .O(gate445inter0));
  nand2 gate548(.a(gate445inter0), .b(s_0), .O(gate445inter1));
  and2  gate549(.a(G1171), .b(G14), .O(gate445inter2));
  inv1  gate550(.a(s_0), .O(gate445inter3));
  inv1  gate551(.a(s_1), .O(gate445inter4));
  nand2 gate552(.a(gate445inter4), .b(gate445inter3), .O(gate445inter5));
  nor2  gate553(.a(gate445inter5), .b(gate445inter2), .O(gate445inter6));
  inv1  gate554(.a(G14), .O(gate445inter7));
  inv1  gate555(.a(G1171), .O(gate445inter8));
  nand2 gate556(.a(gate445inter8), .b(gate445inter7), .O(gate445inter9));
  nand2 gate557(.a(s_1), .b(gate445inter3), .O(gate445inter10));
  nor2  gate558(.a(gate445inter10), .b(gate445inter9), .O(gate445inter11));
  nor2  gate559(.a(gate445inter11), .b(gate445inter6), .O(gate445inter12));
  nand2 gate560(.a(gate445inter12), .b(gate445inter1), .O(G1254));

  xor2  gate1625(.a(G1171), .b(G1075), .O(gate446inter0));
  nand2 gate1626(.a(gate446inter0), .b(s_154), .O(gate446inter1));
  and2  gate1627(.a(G1171), .b(G1075), .O(gate446inter2));
  inv1  gate1628(.a(s_154), .O(gate446inter3));
  inv1  gate1629(.a(s_155), .O(gate446inter4));
  nand2 gate1630(.a(gate446inter4), .b(gate446inter3), .O(gate446inter5));
  nor2  gate1631(.a(gate446inter5), .b(gate446inter2), .O(gate446inter6));
  inv1  gate1632(.a(G1075), .O(gate446inter7));
  inv1  gate1633(.a(G1171), .O(gate446inter8));
  nand2 gate1634(.a(gate446inter8), .b(gate446inter7), .O(gate446inter9));
  nand2 gate1635(.a(s_155), .b(gate446inter3), .O(gate446inter10));
  nor2  gate1636(.a(gate446inter10), .b(gate446inter9), .O(gate446inter11));
  nor2  gate1637(.a(gate446inter11), .b(gate446inter6), .O(gate446inter12));
  nand2 gate1638(.a(gate446inter12), .b(gate446inter1), .O(G1255));
nand2 gate447( .a(G15), .b(G1174), .O(G1256) );

  xor2  gate1975(.a(G1174), .b(G1078), .O(gate448inter0));
  nand2 gate1976(.a(gate448inter0), .b(s_204), .O(gate448inter1));
  and2  gate1977(.a(G1174), .b(G1078), .O(gate448inter2));
  inv1  gate1978(.a(s_204), .O(gate448inter3));
  inv1  gate1979(.a(s_205), .O(gate448inter4));
  nand2 gate1980(.a(gate448inter4), .b(gate448inter3), .O(gate448inter5));
  nor2  gate1981(.a(gate448inter5), .b(gate448inter2), .O(gate448inter6));
  inv1  gate1982(.a(G1078), .O(gate448inter7));
  inv1  gate1983(.a(G1174), .O(gate448inter8));
  nand2 gate1984(.a(gate448inter8), .b(gate448inter7), .O(gate448inter9));
  nand2 gate1985(.a(s_205), .b(gate448inter3), .O(gate448inter10));
  nor2  gate1986(.a(gate448inter10), .b(gate448inter9), .O(gate448inter11));
  nor2  gate1987(.a(gate448inter11), .b(gate448inter6), .O(gate448inter12));
  nand2 gate1988(.a(gate448inter12), .b(gate448inter1), .O(G1257));
nand2 gate449( .a(G16), .b(G1177), .O(G1258) );
nand2 gate450( .a(G1081), .b(G1177), .O(G1259) );
nand2 gate451( .a(G17), .b(G1180), .O(G1260) );
nand2 gate452( .a(G1084), .b(G1180), .O(G1261) );

  xor2  gate701(.a(G1183), .b(G18), .O(gate453inter0));
  nand2 gate702(.a(gate453inter0), .b(s_22), .O(gate453inter1));
  and2  gate703(.a(G1183), .b(G18), .O(gate453inter2));
  inv1  gate704(.a(s_22), .O(gate453inter3));
  inv1  gate705(.a(s_23), .O(gate453inter4));
  nand2 gate706(.a(gate453inter4), .b(gate453inter3), .O(gate453inter5));
  nor2  gate707(.a(gate453inter5), .b(gate453inter2), .O(gate453inter6));
  inv1  gate708(.a(G18), .O(gate453inter7));
  inv1  gate709(.a(G1183), .O(gate453inter8));
  nand2 gate710(.a(gate453inter8), .b(gate453inter7), .O(gate453inter9));
  nand2 gate711(.a(s_23), .b(gate453inter3), .O(gate453inter10));
  nor2  gate712(.a(gate453inter10), .b(gate453inter9), .O(gate453inter11));
  nor2  gate713(.a(gate453inter11), .b(gate453inter6), .O(gate453inter12));
  nand2 gate714(.a(gate453inter12), .b(gate453inter1), .O(G1262));
nand2 gate454( .a(G1087), .b(G1183), .O(G1263) );
nand2 gate455( .a(G19), .b(G1186), .O(G1264) );
nand2 gate456( .a(G1090), .b(G1186), .O(G1265) );
nand2 gate457( .a(G20), .b(G1189), .O(G1266) );
nand2 gate458( .a(G1093), .b(G1189), .O(G1267) );

  xor2  gate1471(.a(G1192), .b(G21), .O(gate459inter0));
  nand2 gate1472(.a(gate459inter0), .b(s_132), .O(gate459inter1));
  and2  gate1473(.a(G1192), .b(G21), .O(gate459inter2));
  inv1  gate1474(.a(s_132), .O(gate459inter3));
  inv1  gate1475(.a(s_133), .O(gate459inter4));
  nand2 gate1476(.a(gate459inter4), .b(gate459inter3), .O(gate459inter5));
  nor2  gate1477(.a(gate459inter5), .b(gate459inter2), .O(gate459inter6));
  inv1  gate1478(.a(G21), .O(gate459inter7));
  inv1  gate1479(.a(G1192), .O(gate459inter8));
  nand2 gate1480(.a(gate459inter8), .b(gate459inter7), .O(gate459inter9));
  nand2 gate1481(.a(s_133), .b(gate459inter3), .O(gate459inter10));
  nor2  gate1482(.a(gate459inter10), .b(gate459inter9), .O(gate459inter11));
  nor2  gate1483(.a(gate459inter11), .b(gate459inter6), .O(gate459inter12));
  nand2 gate1484(.a(gate459inter12), .b(gate459inter1), .O(G1268));

  xor2  gate617(.a(G1192), .b(G1096), .O(gate460inter0));
  nand2 gate618(.a(gate460inter0), .b(s_10), .O(gate460inter1));
  and2  gate619(.a(G1192), .b(G1096), .O(gate460inter2));
  inv1  gate620(.a(s_10), .O(gate460inter3));
  inv1  gate621(.a(s_11), .O(gate460inter4));
  nand2 gate622(.a(gate460inter4), .b(gate460inter3), .O(gate460inter5));
  nor2  gate623(.a(gate460inter5), .b(gate460inter2), .O(gate460inter6));
  inv1  gate624(.a(G1096), .O(gate460inter7));
  inv1  gate625(.a(G1192), .O(gate460inter8));
  nand2 gate626(.a(gate460inter8), .b(gate460inter7), .O(gate460inter9));
  nand2 gate627(.a(s_11), .b(gate460inter3), .O(gate460inter10));
  nor2  gate628(.a(gate460inter10), .b(gate460inter9), .O(gate460inter11));
  nor2  gate629(.a(gate460inter11), .b(gate460inter6), .O(gate460inter12));
  nand2 gate630(.a(gate460inter12), .b(gate460inter1), .O(G1269));
nand2 gate461( .a(G22), .b(G1195), .O(G1270) );

  xor2  gate1093(.a(G1195), .b(G1099), .O(gate462inter0));
  nand2 gate1094(.a(gate462inter0), .b(s_78), .O(gate462inter1));
  and2  gate1095(.a(G1195), .b(G1099), .O(gate462inter2));
  inv1  gate1096(.a(s_78), .O(gate462inter3));
  inv1  gate1097(.a(s_79), .O(gate462inter4));
  nand2 gate1098(.a(gate462inter4), .b(gate462inter3), .O(gate462inter5));
  nor2  gate1099(.a(gate462inter5), .b(gate462inter2), .O(gate462inter6));
  inv1  gate1100(.a(G1099), .O(gate462inter7));
  inv1  gate1101(.a(G1195), .O(gate462inter8));
  nand2 gate1102(.a(gate462inter8), .b(gate462inter7), .O(gate462inter9));
  nand2 gate1103(.a(s_79), .b(gate462inter3), .O(gate462inter10));
  nor2  gate1104(.a(gate462inter10), .b(gate462inter9), .O(gate462inter11));
  nor2  gate1105(.a(gate462inter11), .b(gate462inter6), .O(gate462inter12));
  nand2 gate1106(.a(gate462inter12), .b(gate462inter1), .O(G1271));
nand2 gate463( .a(G23), .b(G1198), .O(G1272) );
nand2 gate464( .a(G1102), .b(G1198), .O(G1273) );
nand2 gate465( .a(G24), .b(G1201), .O(G1274) );

  xor2  gate1835(.a(G1201), .b(G1105), .O(gate466inter0));
  nand2 gate1836(.a(gate466inter0), .b(s_184), .O(gate466inter1));
  and2  gate1837(.a(G1201), .b(G1105), .O(gate466inter2));
  inv1  gate1838(.a(s_184), .O(gate466inter3));
  inv1  gate1839(.a(s_185), .O(gate466inter4));
  nand2 gate1840(.a(gate466inter4), .b(gate466inter3), .O(gate466inter5));
  nor2  gate1841(.a(gate466inter5), .b(gate466inter2), .O(gate466inter6));
  inv1  gate1842(.a(G1105), .O(gate466inter7));
  inv1  gate1843(.a(G1201), .O(gate466inter8));
  nand2 gate1844(.a(gate466inter8), .b(gate466inter7), .O(gate466inter9));
  nand2 gate1845(.a(s_185), .b(gate466inter3), .O(gate466inter10));
  nor2  gate1846(.a(gate466inter10), .b(gate466inter9), .O(gate466inter11));
  nor2  gate1847(.a(gate466inter11), .b(gate466inter6), .O(gate466inter12));
  nand2 gate1848(.a(gate466inter12), .b(gate466inter1), .O(G1275));

  xor2  gate715(.a(G1204), .b(G25), .O(gate467inter0));
  nand2 gate716(.a(gate467inter0), .b(s_24), .O(gate467inter1));
  and2  gate717(.a(G1204), .b(G25), .O(gate467inter2));
  inv1  gate718(.a(s_24), .O(gate467inter3));
  inv1  gate719(.a(s_25), .O(gate467inter4));
  nand2 gate720(.a(gate467inter4), .b(gate467inter3), .O(gate467inter5));
  nor2  gate721(.a(gate467inter5), .b(gate467inter2), .O(gate467inter6));
  inv1  gate722(.a(G25), .O(gate467inter7));
  inv1  gate723(.a(G1204), .O(gate467inter8));
  nand2 gate724(.a(gate467inter8), .b(gate467inter7), .O(gate467inter9));
  nand2 gate725(.a(s_25), .b(gate467inter3), .O(gate467inter10));
  nor2  gate726(.a(gate467inter10), .b(gate467inter9), .O(gate467inter11));
  nor2  gate727(.a(gate467inter11), .b(gate467inter6), .O(gate467inter12));
  nand2 gate728(.a(gate467inter12), .b(gate467inter1), .O(G1276));
nand2 gate468( .a(G1108), .b(G1204), .O(G1277) );

  xor2  gate1863(.a(G1207), .b(G26), .O(gate469inter0));
  nand2 gate1864(.a(gate469inter0), .b(s_188), .O(gate469inter1));
  and2  gate1865(.a(G1207), .b(G26), .O(gate469inter2));
  inv1  gate1866(.a(s_188), .O(gate469inter3));
  inv1  gate1867(.a(s_189), .O(gate469inter4));
  nand2 gate1868(.a(gate469inter4), .b(gate469inter3), .O(gate469inter5));
  nor2  gate1869(.a(gate469inter5), .b(gate469inter2), .O(gate469inter6));
  inv1  gate1870(.a(G26), .O(gate469inter7));
  inv1  gate1871(.a(G1207), .O(gate469inter8));
  nand2 gate1872(.a(gate469inter8), .b(gate469inter7), .O(gate469inter9));
  nand2 gate1873(.a(s_189), .b(gate469inter3), .O(gate469inter10));
  nor2  gate1874(.a(gate469inter10), .b(gate469inter9), .O(gate469inter11));
  nor2  gate1875(.a(gate469inter11), .b(gate469inter6), .O(gate469inter12));
  nand2 gate1876(.a(gate469inter12), .b(gate469inter1), .O(G1278));

  xor2  gate2101(.a(G1207), .b(G1111), .O(gate470inter0));
  nand2 gate2102(.a(gate470inter0), .b(s_222), .O(gate470inter1));
  and2  gate2103(.a(G1207), .b(G1111), .O(gate470inter2));
  inv1  gate2104(.a(s_222), .O(gate470inter3));
  inv1  gate2105(.a(s_223), .O(gate470inter4));
  nand2 gate2106(.a(gate470inter4), .b(gate470inter3), .O(gate470inter5));
  nor2  gate2107(.a(gate470inter5), .b(gate470inter2), .O(gate470inter6));
  inv1  gate2108(.a(G1111), .O(gate470inter7));
  inv1  gate2109(.a(G1207), .O(gate470inter8));
  nand2 gate2110(.a(gate470inter8), .b(gate470inter7), .O(gate470inter9));
  nand2 gate2111(.a(s_223), .b(gate470inter3), .O(gate470inter10));
  nor2  gate2112(.a(gate470inter10), .b(gate470inter9), .O(gate470inter11));
  nor2  gate2113(.a(gate470inter11), .b(gate470inter6), .O(gate470inter12));
  nand2 gate2114(.a(gate470inter12), .b(gate470inter1), .O(G1279));
nand2 gate471( .a(G27), .b(G1210), .O(G1280) );
nand2 gate472( .a(G1114), .b(G1210), .O(G1281) );
nand2 gate473( .a(G28), .b(G1213), .O(G1282) );
nand2 gate474( .a(G1117), .b(G1213), .O(G1283) );
nand2 gate475( .a(G29), .b(G1216), .O(G1284) );
nand2 gate476( .a(G1120), .b(G1216), .O(G1285) );
nand2 gate477( .a(G30), .b(G1219), .O(G1286) );
nand2 gate478( .a(G1123), .b(G1219), .O(G1287) );
nand2 gate479( .a(G31), .b(G1222), .O(G1288) );

  xor2  gate1429(.a(G1222), .b(G1126), .O(gate480inter0));
  nand2 gate1430(.a(gate480inter0), .b(s_126), .O(gate480inter1));
  and2  gate1431(.a(G1222), .b(G1126), .O(gate480inter2));
  inv1  gate1432(.a(s_126), .O(gate480inter3));
  inv1  gate1433(.a(s_127), .O(gate480inter4));
  nand2 gate1434(.a(gate480inter4), .b(gate480inter3), .O(gate480inter5));
  nor2  gate1435(.a(gate480inter5), .b(gate480inter2), .O(gate480inter6));
  inv1  gate1436(.a(G1126), .O(gate480inter7));
  inv1  gate1437(.a(G1222), .O(gate480inter8));
  nand2 gate1438(.a(gate480inter8), .b(gate480inter7), .O(gate480inter9));
  nand2 gate1439(.a(s_127), .b(gate480inter3), .O(gate480inter10));
  nor2  gate1440(.a(gate480inter10), .b(gate480inter9), .O(gate480inter11));
  nor2  gate1441(.a(gate480inter11), .b(gate480inter6), .O(gate480inter12));
  nand2 gate1442(.a(gate480inter12), .b(gate480inter1), .O(G1289));

  xor2  gate1737(.a(G1225), .b(G32), .O(gate481inter0));
  nand2 gate1738(.a(gate481inter0), .b(s_170), .O(gate481inter1));
  and2  gate1739(.a(G1225), .b(G32), .O(gate481inter2));
  inv1  gate1740(.a(s_170), .O(gate481inter3));
  inv1  gate1741(.a(s_171), .O(gate481inter4));
  nand2 gate1742(.a(gate481inter4), .b(gate481inter3), .O(gate481inter5));
  nor2  gate1743(.a(gate481inter5), .b(gate481inter2), .O(gate481inter6));
  inv1  gate1744(.a(G32), .O(gate481inter7));
  inv1  gate1745(.a(G1225), .O(gate481inter8));
  nand2 gate1746(.a(gate481inter8), .b(gate481inter7), .O(gate481inter9));
  nand2 gate1747(.a(s_171), .b(gate481inter3), .O(gate481inter10));
  nor2  gate1748(.a(gate481inter10), .b(gate481inter9), .O(gate481inter11));
  nor2  gate1749(.a(gate481inter11), .b(gate481inter6), .O(gate481inter12));
  nand2 gate1750(.a(gate481inter12), .b(gate481inter1), .O(G1290));
nand2 gate482( .a(G1129), .b(G1225), .O(G1291) );

  xor2  gate2885(.a(G1229), .b(G1228), .O(gate483inter0));
  nand2 gate2886(.a(gate483inter0), .b(s_334), .O(gate483inter1));
  and2  gate2887(.a(G1229), .b(G1228), .O(gate483inter2));
  inv1  gate2888(.a(s_334), .O(gate483inter3));
  inv1  gate2889(.a(s_335), .O(gate483inter4));
  nand2 gate2890(.a(gate483inter4), .b(gate483inter3), .O(gate483inter5));
  nor2  gate2891(.a(gate483inter5), .b(gate483inter2), .O(gate483inter6));
  inv1  gate2892(.a(G1228), .O(gate483inter7));
  inv1  gate2893(.a(G1229), .O(gate483inter8));
  nand2 gate2894(.a(gate483inter8), .b(gate483inter7), .O(gate483inter9));
  nand2 gate2895(.a(s_335), .b(gate483inter3), .O(gate483inter10));
  nor2  gate2896(.a(gate483inter10), .b(gate483inter9), .O(gate483inter11));
  nor2  gate2897(.a(gate483inter11), .b(gate483inter6), .O(gate483inter12));
  nand2 gate2898(.a(gate483inter12), .b(gate483inter1), .O(G1292));
nand2 gate484( .a(G1230), .b(G1231), .O(G1293) );

  xor2  gate2829(.a(G1233), .b(G1232), .O(gate485inter0));
  nand2 gate2830(.a(gate485inter0), .b(s_326), .O(gate485inter1));
  and2  gate2831(.a(G1233), .b(G1232), .O(gate485inter2));
  inv1  gate2832(.a(s_326), .O(gate485inter3));
  inv1  gate2833(.a(s_327), .O(gate485inter4));
  nand2 gate2834(.a(gate485inter4), .b(gate485inter3), .O(gate485inter5));
  nor2  gate2835(.a(gate485inter5), .b(gate485inter2), .O(gate485inter6));
  inv1  gate2836(.a(G1232), .O(gate485inter7));
  inv1  gate2837(.a(G1233), .O(gate485inter8));
  nand2 gate2838(.a(gate485inter8), .b(gate485inter7), .O(gate485inter9));
  nand2 gate2839(.a(s_327), .b(gate485inter3), .O(gate485inter10));
  nor2  gate2840(.a(gate485inter10), .b(gate485inter9), .O(gate485inter11));
  nor2  gate2841(.a(gate485inter11), .b(gate485inter6), .O(gate485inter12));
  nand2 gate2842(.a(gate485inter12), .b(gate485inter1), .O(G1294));

  xor2  gate2073(.a(G1235), .b(G1234), .O(gate486inter0));
  nand2 gate2074(.a(gate486inter0), .b(s_218), .O(gate486inter1));
  and2  gate2075(.a(G1235), .b(G1234), .O(gate486inter2));
  inv1  gate2076(.a(s_218), .O(gate486inter3));
  inv1  gate2077(.a(s_219), .O(gate486inter4));
  nand2 gate2078(.a(gate486inter4), .b(gate486inter3), .O(gate486inter5));
  nor2  gate2079(.a(gate486inter5), .b(gate486inter2), .O(gate486inter6));
  inv1  gate2080(.a(G1234), .O(gate486inter7));
  inv1  gate2081(.a(G1235), .O(gate486inter8));
  nand2 gate2082(.a(gate486inter8), .b(gate486inter7), .O(gate486inter9));
  nand2 gate2083(.a(s_219), .b(gate486inter3), .O(gate486inter10));
  nor2  gate2084(.a(gate486inter10), .b(gate486inter9), .O(gate486inter11));
  nor2  gate2085(.a(gate486inter11), .b(gate486inter6), .O(gate486inter12));
  nand2 gate2086(.a(gate486inter12), .b(gate486inter1), .O(G1295));
nand2 gate487( .a(G1236), .b(G1237), .O(G1296) );

  xor2  gate2913(.a(G1239), .b(G1238), .O(gate488inter0));
  nand2 gate2914(.a(gate488inter0), .b(s_338), .O(gate488inter1));
  and2  gate2915(.a(G1239), .b(G1238), .O(gate488inter2));
  inv1  gate2916(.a(s_338), .O(gate488inter3));
  inv1  gate2917(.a(s_339), .O(gate488inter4));
  nand2 gate2918(.a(gate488inter4), .b(gate488inter3), .O(gate488inter5));
  nor2  gate2919(.a(gate488inter5), .b(gate488inter2), .O(gate488inter6));
  inv1  gate2920(.a(G1238), .O(gate488inter7));
  inv1  gate2921(.a(G1239), .O(gate488inter8));
  nand2 gate2922(.a(gate488inter8), .b(gate488inter7), .O(gate488inter9));
  nand2 gate2923(.a(s_339), .b(gate488inter3), .O(gate488inter10));
  nor2  gate2924(.a(gate488inter10), .b(gate488inter9), .O(gate488inter11));
  nor2  gate2925(.a(gate488inter11), .b(gate488inter6), .O(gate488inter12));
  nand2 gate2926(.a(gate488inter12), .b(gate488inter1), .O(G1297));

  xor2  gate1849(.a(G1241), .b(G1240), .O(gate489inter0));
  nand2 gate1850(.a(gate489inter0), .b(s_186), .O(gate489inter1));
  and2  gate1851(.a(G1241), .b(G1240), .O(gate489inter2));
  inv1  gate1852(.a(s_186), .O(gate489inter3));
  inv1  gate1853(.a(s_187), .O(gate489inter4));
  nand2 gate1854(.a(gate489inter4), .b(gate489inter3), .O(gate489inter5));
  nor2  gate1855(.a(gate489inter5), .b(gate489inter2), .O(gate489inter6));
  inv1  gate1856(.a(G1240), .O(gate489inter7));
  inv1  gate1857(.a(G1241), .O(gate489inter8));
  nand2 gate1858(.a(gate489inter8), .b(gate489inter7), .O(gate489inter9));
  nand2 gate1859(.a(s_187), .b(gate489inter3), .O(gate489inter10));
  nor2  gate1860(.a(gate489inter10), .b(gate489inter9), .O(gate489inter11));
  nor2  gate1861(.a(gate489inter11), .b(gate489inter6), .O(gate489inter12));
  nand2 gate1862(.a(gate489inter12), .b(gate489inter1), .O(G1298));
nand2 gate490( .a(G1242), .b(G1243), .O(G1299) );
nand2 gate491( .a(G1244), .b(G1245), .O(G1300) );

  xor2  gate2731(.a(G1247), .b(G1246), .O(gate492inter0));
  nand2 gate2732(.a(gate492inter0), .b(s_312), .O(gate492inter1));
  and2  gate2733(.a(G1247), .b(G1246), .O(gate492inter2));
  inv1  gate2734(.a(s_312), .O(gate492inter3));
  inv1  gate2735(.a(s_313), .O(gate492inter4));
  nand2 gate2736(.a(gate492inter4), .b(gate492inter3), .O(gate492inter5));
  nor2  gate2737(.a(gate492inter5), .b(gate492inter2), .O(gate492inter6));
  inv1  gate2738(.a(G1246), .O(gate492inter7));
  inv1  gate2739(.a(G1247), .O(gate492inter8));
  nand2 gate2740(.a(gate492inter8), .b(gate492inter7), .O(gate492inter9));
  nand2 gate2741(.a(s_313), .b(gate492inter3), .O(gate492inter10));
  nor2  gate2742(.a(gate492inter10), .b(gate492inter9), .O(gate492inter11));
  nor2  gate2743(.a(gate492inter11), .b(gate492inter6), .O(gate492inter12));
  nand2 gate2744(.a(gate492inter12), .b(gate492inter1), .O(G1301));

  xor2  gate2675(.a(G1249), .b(G1248), .O(gate493inter0));
  nand2 gate2676(.a(gate493inter0), .b(s_304), .O(gate493inter1));
  and2  gate2677(.a(G1249), .b(G1248), .O(gate493inter2));
  inv1  gate2678(.a(s_304), .O(gate493inter3));
  inv1  gate2679(.a(s_305), .O(gate493inter4));
  nand2 gate2680(.a(gate493inter4), .b(gate493inter3), .O(gate493inter5));
  nor2  gate2681(.a(gate493inter5), .b(gate493inter2), .O(gate493inter6));
  inv1  gate2682(.a(G1248), .O(gate493inter7));
  inv1  gate2683(.a(G1249), .O(gate493inter8));
  nand2 gate2684(.a(gate493inter8), .b(gate493inter7), .O(gate493inter9));
  nand2 gate2685(.a(s_305), .b(gate493inter3), .O(gate493inter10));
  nor2  gate2686(.a(gate493inter10), .b(gate493inter9), .O(gate493inter11));
  nor2  gate2687(.a(gate493inter11), .b(gate493inter6), .O(gate493inter12));
  nand2 gate2688(.a(gate493inter12), .b(gate493inter1), .O(G1302));

  xor2  gate2367(.a(G1251), .b(G1250), .O(gate494inter0));
  nand2 gate2368(.a(gate494inter0), .b(s_260), .O(gate494inter1));
  and2  gate2369(.a(G1251), .b(G1250), .O(gate494inter2));
  inv1  gate2370(.a(s_260), .O(gate494inter3));
  inv1  gate2371(.a(s_261), .O(gate494inter4));
  nand2 gate2372(.a(gate494inter4), .b(gate494inter3), .O(gate494inter5));
  nor2  gate2373(.a(gate494inter5), .b(gate494inter2), .O(gate494inter6));
  inv1  gate2374(.a(G1250), .O(gate494inter7));
  inv1  gate2375(.a(G1251), .O(gate494inter8));
  nand2 gate2376(.a(gate494inter8), .b(gate494inter7), .O(gate494inter9));
  nand2 gate2377(.a(s_261), .b(gate494inter3), .O(gate494inter10));
  nor2  gate2378(.a(gate494inter10), .b(gate494inter9), .O(gate494inter11));
  nor2  gate2379(.a(gate494inter11), .b(gate494inter6), .O(gate494inter12));
  nand2 gate2380(.a(gate494inter12), .b(gate494inter1), .O(G1303));

  xor2  gate2241(.a(G1253), .b(G1252), .O(gate495inter0));
  nand2 gate2242(.a(gate495inter0), .b(s_242), .O(gate495inter1));
  and2  gate2243(.a(G1253), .b(G1252), .O(gate495inter2));
  inv1  gate2244(.a(s_242), .O(gate495inter3));
  inv1  gate2245(.a(s_243), .O(gate495inter4));
  nand2 gate2246(.a(gate495inter4), .b(gate495inter3), .O(gate495inter5));
  nor2  gate2247(.a(gate495inter5), .b(gate495inter2), .O(gate495inter6));
  inv1  gate2248(.a(G1252), .O(gate495inter7));
  inv1  gate2249(.a(G1253), .O(gate495inter8));
  nand2 gate2250(.a(gate495inter8), .b(gate495inter7), .O(gate495inter9));
  nand2 gate2251(.a(s_243), .b(gate495inter3), .O(gate495inter10));
  nor2  gate2252(.a(gate495inter10), .b(gate495inter9), .O(gate495inter11));
  nor2  gate2253(.a(gate495inter11), .b(gate495inter6), .O(gate495inter12));
  nand2 gate2254(.a(gate495inter12), .b(gate495inter1), .O(G1304));
nand2 gate496( .a(G1254), .b(G1255), .O(G1305) );

  xor2  gate2437(.a(G1257), .b(G1256), .O(gate497inter0));
  nand2 gate2438(.a(gate497inter0), .b(s_270), .O(gate497inter1));
  and2  gate2439(.a(G1257), .b(G1256), .O(gate497inter2));
  inv1  gate2440(.a(s_270), .O(gate497inter3));
  inv1  gate2441(.a(s_271), .O(gate497inter4));
  nand2 gate2442(.a(gate497inter4), .b(gate497inter3), .O(gate497inter5));
  nor2  gate2443(.a(gate497inter5), .b(gate497inter2), .O(gate497inter6));
  inv1  gate2444(.a(G1256), .O(gate497inter7));
  inv1  gate2445(.a(G1257), .O(gate497inter8));
  nand2 gate2446(.a(gate497inter8), .b(gate497inter7), .O(gate497inter9));
  nand2 gate2447(.a(s_271), .b(gate497inter3), .O(gate497inter10));
  nor2  gate2448(.a(gate497inter10), .b(gate497inter9), .O(gate497inter11));
  nor2  gate2449(.a(gate497inter11), .b(gate497inter6), .O(gate497inter12));
  nand2 gate2450(.a(gate497inter12), .b(gate497inter1), .O(G1306));

  xor2  gate2507(.a(G1259), .b(G1258), .O(gate498inter0));
  nand2 gate2508(.a(gate498inter0), .b(s_280), .O(gate498inter1));
  and2  gate2509(.a(G1259), .b(G1258), .O(gate498inter2));
  inv1  gate2510(.a(s_280), .O(gate498inter3));
  inv1  gate2511(.a(s_281), .O(gate498inter4));
  nand2 gate2512(.a(gate498inter4), .b(gate498inter3), .O(gate498inter5));
  nor2  gate2513(.a(gate498inter5), .b(gate498inter2), .O(gate498inter6));
  inv1  gate2514(.a(G1258), .O(gate498inter7));
  inv1  gate2515(.a(G1259), .O(gate498inter8));
  nand2 gate2516(.a(gate498inter8), .b(gate498inter7), .O(gate498inter9));
  nand2 gate2517(.a(s_281), .b(gate498inter3), .O(gate498inter10));
  nor2  gate2518(.a(gate498inter10), .b(gate498inter9), .O(gate498inter11));
  nor2  gate2519(.a(gate498inter11), .b(gate498inter6), .O(gate498inter12));
  nand2 gate2520(.a(gate498inter12), .b(gate498inter1), .O(G1307));
nand2 gate499( .a(G1260), .b(G1261), .O(G1308) );
nand2 gate500( .a(G1262), .b(G1263), .O(G1309) );
nand2 gate501( .a(G1264), .b(G1265), .O(G1310) );
nand2 gate502( .a(G1266), .b(G1267), .O(G1311) );
nand2 gate503( .a(G1268), .b(G1269), .O(G1312) );
nand2 gate504( .a(G1270), .b(G1271), .O(G1313) );

  xor2  gate2647(.a(G1273), .b(G1272), .O(gate505inter0));
  nand2 gate2648(.a(gate505inter0), .b(s_300), .O(gate505inter1));
  and2  gate2649(.a(G1273), .b(G1272), .O(gate505inter2));
  inv1  gate2650(.a(s_300), .O(gate505inter3));
  inv1  gate2651(.a(s_301), .O(gate505inter4));
  nand2 gate2652(.a(gate505inter4), .b(gate505inter3), .O(gate505inter5));
  nor2  gate2653(.a(gate505inter5), .b(gate505inter2), .O(gate505inter6));
  inv1  gate2654(.a(G1272), .O(gate505inter7));
  inv1  gate2655(.a(G1273), .O(gate505inter8));
  nand2 gate2656(.a(gate505inter8), .b(gate505inter7), .O(gate505inter9));
  nand2 gate2657(.a(s_301), .b(gate505inter3), .O(gate505inter10));
  nor2  gate2658(.a(gate505inter10), .b(gate505inter9), .O(gate505inter11));
  nor2  gate2659(.a(gate505inter11), .b(gate505inter6), .O(gate505inter12));
  nand2 gate2660(.a(gate505inter12), .b(gate505inter1), .O(G1314));

  xor2  gate981(.a(G1275), .b(G1274), .O(gate506inter0));
  nand2 gate982(.a(gate506inter0), .b(s_62), .O(gate506inter1));
  and2  gate983(.a(G1275), .b(G1274), .O(gate506inter2));
  inv1  gate984(.a(s_62), .O(gate506inter3));
  inv1  gate985(.a(s_63), .O(gate506inter4));
  nand2 gate986(.a(gate506inter4), .b(gate506inter3), .O(gate506inter5));
  nor2  gate987(.a(gate506inter5), .b(gate506inter2), .O(gate506inter6));
  inv1  gate988(.a(G1274), .O(gate506inter7));
  inv1  gate989(.a(G1275), .O(gate506inter8));
  nand2 gate990(.a(gate506inter8), .b(gate506inter7), .O(gate506inter9));
  nand2 gate991(.a(s_63), .b(gate506inter3), .O(gate506inter10));
  nor2  gate992(.a(gate506inter10), .b(gate506inter9), .O(gate506inter11));
  nor2  gate993(.a(gate506inter11), .b(gate506inter6), .O(gate506inter12));
  nand2 gate994(.a(gate506inter12), .b(gate506inter1), .O(G1315));

  xor2  gate1457(.a(G1277), .b(G1276), .O(gate507inter0));
  nand2 gate1458(.a(gate507inter0), .b(s_130), .O(gate507inter1));
  and2  gate1459(.a(G1277), .b(G1276), .O(gate507inter2));
  inv1  gate1460(.a(s_130), .O(gate507inter3));
  inv1  gate1461(.a(s_131), .O(gate507inter4));
  nand2 gate1462(.a(gate507inter4), .b(gate507inter3), .O(gate507inter5));
  nor2  gate1463(.a(gate507inter5), .b(gate507inter2), .O(gate507inter6));
  inv1  gate1464(.a(G1276), .O(gate507inter7));
  inv1  gate1465(.a(G1277), .O(gate507inter8));
  nand2 gate1466(.a(gate507inter8), .b(gate507inter7), .O(gate507inter9));
  nand2 gate1467(.a(s_131), .b(gate507inter3), .O(gate507inter10));
  nor2  gate1468(.a(gate507inter10), .b(gate507inter9), .O(gate507inter11));
  nor2  gate1469(.a(gate507inter11), .b(gate507inter6), .O(gate507inter12));
  nand2 gate1470(.a(gate507inter12), .b(gate507inter1), .O(G1316));
nand2 gate508( .a(G1278), .b(G1279), .O(G1317) );

  xor2  gate631(.a(G1281), .b(G1280), .O(gate509inter0));
  nand2 gate632(.a(gate509inter0), .b(s_12), .O(gate509inter1));
  and2  gate633(.a(G1281), .b(G1280), .O(gate509inter2));
  inv1  gate634(.a(s_12), .O(gate509inter3));
  inv1  gate635(.a(s_13), .O(gate509inter4));
  nand2 gate636(.a(gate509inter4), .b(gate509inter3), .O(gate509inter5));
  nor2  gate637(.a(gate509inter5), .b(gate509inter2), .O(gate509inter6));
  inv1  gate638(.a(G1280), .O(gate509inter7));
  inv1  gate639(.a(G1281), .O(gate509inter8));
  nand2 gate640(.a(gate509inter8), .b(gate509inter7), .O(gate509inter9));
  nand2 gate641(.a(s_13), .b(gate509inter3), .O(gate509inter10));
  nor2  gate642(.a(gate509inter10), .b(gate509inter9), .O(gate509inter11));
  nor2  gate643(.a(gate509inter11), .b(gate509inter6), .O(gate509inter12));
  nand2 gate644(.a(gate509inter12), .b(gate509inter1), .O(G1318));

  xor2  gate561(.a(G1283), .b(G1282), .O(gate510inter0));
  nand2 gate562(.a(gate510inter0), .b(s_2), .O(gate510inter1));
  and2  gate563(.a(G1283), .b(G1282), .O(gate510inter2));
  inv1  gate564(.a(s_2), .O(gate510inter3));
  inv1  gate565(.a(s_3), .O(gate510inter4));
  nand2 gate566(.a(gate510inter4), .b(gate510inter3), .O(gate510inter5));
  nor2  gate567(.a(gate510inter5), .b(gate510inter2), .O(gate510inter6));
  inv1  gate568(.a(G1282), .O(gate510inter7));
  inv1  gate569(.a(G1283), .O(gate510inter8));
  nand2 gate570(.a(gate510inter8), .b(gate510inter7), .O(gate510inter9));
  nand2 gate571(.a(s_3), .b(gate510inter3), .O(gate510inter10));
  nor2  gate572(.a(gate510inter10), .b(gate510inter9), .O(gate510inter11));
  nor2  gate573(.a(gate510inter11), .b(gate510inter6), .O(gate510inter12));
  nand2 gate574(.a(gate510inter12), .b(gate510inter1), .O(G1319));

  xor2  gate2381(.a(G1285), .b(G1284), .O(gate511inter0));
  nand2 gate2382(.a(gate511inter0), .b(s_262), .O(gate511inter1));
  and2  gate2383(.a(G1285), .b(G1284), .O(gate511inter2));
  inv1  gate2384(.a(s_262), .O(gate511inter3));
  inv1  gate2385(.a(s_263), .O(gate511inter4));
  nand2 gate2386(.a(gate511inter4), .b(gate511inter3), .O(gate511inter5));
  nor2  gate2387(.a(gate511inter5), .b(gate511inter2), .O(gate511inter6));
  inv1  gate2388(.a(G1284), .O(gate511inter7));
  inv1  gate2389(.a(G1285), .O(gate511inter8));
  nand2 gate2390(.a(gate511inter8), .b(gate511inter7), .O(gate511inter9));
  nand2 gate2391(.a(s_263), .b(gate511inter3), .O(gate511inter10));
  nor2  gate2392(.a(gate511inter10), .b(gate511inter9), .O(gate511inter11));
  nor2  gate2393(.a(gate511inter11), .b(gate511inter6), .O(gate511inter12));
  nand2 gate2394(.a(gate511inter12), .b(gate511inter1), .O(G1320));
nand2 gate512( .a(G1286), .b(G1287), .O(G1321) );
nand2 gate513( .a(G1288), .b(G1289), .O(G1322) );

  xor2  gate2185(.a(G1291), .b(G1290), .O(gate514inter0));
  nand2 gate2186(.a(gate514inter0), .b(s_234), .O(gate514inter1));
  and2  gate2187(.a(G1291), .b(G1290), .O(gate514inter2));
  inv1  gate2188(.a(s_234), .O(gate514inter3));
  inv1  gate2189(.a(s_235), .O(gate514inter4));
  nand2 gate2190(.a(gate514inter4), .b(gate514inter3), .O(gate514inter5));
  nor2  gate2191(.a(gate514inter5), .b(gate514inter2), .O(gate514inter6));
  inv1  gate2192(.a(G1290), .O(gate514inter7));
  inv1  gate2193(.a(G1291), .O(gate514inter8));
  nand2 gate2194(.a(gate514inter8), .b(gate514inter7), .O(gate514inter9));
  nand2 gate2195(.a(s_235), .b(gate514inter3), .O(gate514inter10));
  nor2  gate2196(.a(gate514inter10), .b(gate514inter9), .O(gate514inter11));
  nor2  gate2197(.a(gate514inter11), .b(gate514inter6), .O(gate514inter12));
  nand2 gate2198(.a(gate514inter12), .b(gate514inter1), .O(G1323));
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule