module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);

input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;//RE__PI;

input s_0,s_1;//RE__ALLOW(00,01,10,11);
input s_2,s_3;//RE__ALLOW(00,01,10,11);
input s_4,s_5;//RE__ALLOW(00,01,10,11);
input s_6,s_7;//RE__ALLOW(00,01,10,11);
input s_8,s_9;//RE__ALLOW(00,01,10,11);
input s_10,s_11;//RE__ALLOW(00,01,10,11);
input s_12,s_13;//RE__ALLOW(00,01,10,11);
input s_14,s_15;//RE__ALLOW(00,01,10,11);
input s_16,s_17;//RE__ALLOW(00,01,10,11);
input s_18,s_19;//RE__ALLOW(00,01,10,11);
input s_20,s_21;//RE__ALLOW(00,01,10,11);
input s_22,s_23;//RE__ALLOW(00,01,10,11);
input s_24,s_25;//RE__ALLOW(00,01,10,11);
input s_26,s_27;//RE__ALLOW(00,01,10,11);
input s_28,s_29;//RE__ALLOW(00,01,10,11);
input s_30,s_31;//RE__ALLOW(00,01,10,11);
input s_32,s_33;//RE__ALLOW(00,01,10,11);
input s_34,s_35;//RE__ALLOW(00,01,10,11);
input s_36,s_37;//RE__ALLOW(00,01,10,11);
input s_38,s_39;//RE__ALLOW(00,01,10,11);
input s_40,s_41;//RE__ALLOW(00,01,10,11);
input s_42,s_43;//RE__ALLOW(00,01,10,11);
input s_44,s_45;//RE__ALLOW(00,01,10,11);
input s_46,s_47;//RE__ALLOW(00,01,10,11);
input s_48,s_49;//RE__ALLOW(00,01,10,11);
input s_50,s_51;//RE__ALLOW(00,01,10,11);
input s_52,s_53;//RE__ALLOW(00,01,10,11);
input s_54,s_55;//RE__ALLOW(00,01,10,11);
input s_56,s_57;//RE__ALLOW(00,01,10,11);
input s_58,s_59;//RE__ALLOW(00,01,10,11);
input s_60,s_61;//RE__ALLOW(00,01,10,11);
input s_62,s_63;//RE__ALLOW(00,01,10,11);
input s_64,s_65;//RE__ALLOW(00,01,10,11);
input s_66,s_67;//RE__ALLOW(00,01,10,11);
input s_68,s_69;//RE__ALLOW(00,01,10,11);
input s_70,s_71;//RE__ALLOW(00,01,10,11);
input s_72,s_73;//RE__ALLOW(00,01,10,11);
input s_74,s_75;//RE__ALLOW(00,01,10,11);
input s_76,s_77;//RE__ALLOW(00,01,10,11);
input s_78,s_79;//RE__ALLOW(00,01,10,11);
input s_80,s_81;//RE__ALLOW(00,01,10,11);
input s_82,s_83;//RE__ALLOW(00,01,10,11);
input s_84,s_85;//RE__ALLOW(00,01,10,11);
input s_86,s_87;//RE__ALLOW(00,01,10,11);
input s_88,s_89;//RE__ALLOW(00,01,10,11);
input s_90,s_91;//RE__ALLOW(00,01,10,11);
input s_92,s_93;//RE__ALLOW(00,01,10,11);
input s_94,s_95;//RE__ALLOW(00,01,10,11);
input s_96,s_97;//RE__ALLOW(00,01,10,11);
input s_98,s_99;//RE__ALLOW(00,01,10,11);
input s_100,s_101;//RE__ALLOW(00,01,10,11);
input s_102,s_103;//RE__ALLOW(00,01,10,11);
input s_104,s_105;//RE__ALLOW(00,01,10,11);
input s_106,s_107;//RE__ALLOW(00,01,10,11);
input s_108,s_109;//RE__ALLOW(00,01,10,11);
input s_110,s_111;//RE__ALLOW(00,01,10,11);
input s_112,s_113;//RE__ALLOW(00,01,10,11);
input s_114,s_115;//RE__ALLOW(00,01,10,11);
input s_116,s_117;//RE__ALLOW(00,01,10,11);
input s_118,s_119;//RE__ALLOW(00,01,10,11);
input s_120,s_121;//RE__ALLOW(00,01,10,11);
input s_122,s_123;//RE__ALLOW(00,01,10,11);
input s_124,s_125;//RE__ALLOW(00,01,10,11);
input s_126,s_127;//RE__ALLOW(00,01,10,11);
input s_128,s_129;//RE__ALLOW(00,01,10,11);
input s_130,s_131;//RE__ALLOW(00,01,10,11);
input s_132,s_133;//RE__ALLOW(00,01,10,11);
input s_134,s_135;//RE__ALLOW(00,01,10,11);
input s_136,s_137;//RE__ALLOW(00,01,10,11);
input s_138,s_139;//RE__ALLOW(00,01,10,11);
input s_140,s_141;//RE__ALLOW(00,01,10,11);
input s_142,s_143;//RE__ALLOW(00,01,10,11);
input s_144,s_145;//RE__ALLOW(00,01,10,11);
input s_146,s_147;//RE__ALLOW(00,01,10,11);
input s_148,s_149;//RE__ALLOW(00,01,10,11);
input s_150,s_151;//RE__ALLOW(00,01,10,11);
input s_152,s_153;//RE__ALLOW(00,01,10,11);
input s_154,s_155;//RE__ALLOW(00,01,10,11);
input s_156,s_157;//RE__ALLOW(00,01,10,11);
input s_158,s_159;//RE__ALLOW(00,01,10,11);
input s_160,s_161;//RE__ALLOW(00,01,10,11);
input s_162,s_163;//RE__ALLOW(00,01,10,11);
input s_164,s_165;//RE__ALLOW(00,01,10,11);
input s_166,s_167;//RE__ALLOW(00,01,10,11);
input s_168,s_169;//RE__ALLOW(00,01,10,11);
input s_170,s_171;//RE__ALLOW(00,01,10,11);
input s_172,s_173;//RE__ALLOW(00,01,10,11);
input s_174,s_175;//RE__ALLOW(00,01,10,11);
input s_176,s_177;//RE__ALLOW(00,01,10,11);
input s_178,s_179;//RE__ALLOW(00,01,10,11);
input s_180,s_181;//RE__ALLOW(00,01,10,11);
input s_182,s_183;//RE__ALLOW(00,01,10,11);
input s_184,s_185;//RE__ALLOW(00,01,10,11);
input s_186,s_187;//RE__ALLOW(00,01,10,11);
input s_188,s_189;//RE__ALLOW(00,01,10,11);
input s_190,s_191;//RE__ALLOW(00,01,10,11);
input s_192,s_193;//RE__ALLOW(00,01,10,11);
input s_194,s_195;//RE__ALLOW(00,01,10,11);
input s_196,s_197;//RE__ALLOW(00,01,10,11);
input s_198,s_199;//RE__ALLOW(00,01,10,11);
input s_200,s_201;//RE__ALLOW(00,01,10,11);
input s_202,s_203;//RE__ALLOW(00,01,10,11);
input s_204,s_205;//RE__ALLOW(00,01,10,11);
input s_206,s_207;//RE__ALLOW(00,01,10,11);
input s_208,s_209;//RE__ALLOW(00,01,10,11);
input s_210,s_211;//RE__ALLOW(00,01,10,11);
input s_212,s_213;//RE__ALLOW(00,01,10,11);
input s_214,s_215;//RE__ALLOW(00,01,10,11);
input s_216,s_217;//RE__ALLOW(00,01,10,11);
input s_218,s_219;//RE__ALLOW(00,01,10,11);
input s_220,s_221;//RE__ALLOW(00,01,10,11);
input s_222,s_223;//RE__ALLOW(00,01,10,11);
input s_224,s_225;//RE__ALLOW(00,01,10,11);
input s_226,s_227;//RE__ALLOW(00,01,10,11);
input s_228,s_229;//RE__ALLOW(00,01,10,11);
input s_230,s_231;//RE__ALLOW(00,01,10,11);
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;

  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate242inter0, gate242inter1, gate242inter2, gate242inter3, gate242inter4, gate242inter5, gate242inter6, gate242inter7, gate242inter8, gate242inter9, gate242inter10, gate242inter11, gate242inter12, gate394inter0, gate394inter1, gate394inter2, gate394inter3, gate394inter4, gate394inter5, gate394inter6, gate394inter7, gate394inter8, gate394inter9, gate394inter10, gate394inter11, gate394inter12, gate107inter0, gate107inter1, gate107inter2, gate107inter3, gate107inter4, gate107inter5, gate107inter6, gate107inter7, gate107inter8, gate107inter9, gate107inter10, gate107inter11, gate107inter12, gate157inter0, gate157inter1, gate157inter2, gate157inter3, gate157inter4, gate157inter5, gate157inter6, gate157inter7, gate157inter8, gate157inter9, gate157inter10, gate157inter11, gate157inter12, gate228inter0, gate228inter1, gate228inter2, gate228inter3, gate228inter4, gate228inter5, gate228inter6, gate228inter7, gate228inter8, gate228inter9, gate228inter10, gate228inter11, gate228inter12, gate29inter0, gate29inter1, gate29inter2, gate29inter3, gate29inter4, gate29inter5, gate29inter6, gate29inter7, gate29inter8, gate29inter9, gate29inter10, gate29inter11, gate29inter12, gate111inter0, gate111inter1, gate111inter2, gate111inter3, gate111inter4, gate111inter5, gate111inter6, gate111inter7, gate111inter8, gate111inter9, gate111inter10, gate111inter11, gate111inter12, gate500inter0, gate500inter1, gate500inter2, gate500inter3, gate500inter4, gate500inter5, gate500inter6, gate500inter7, gate500inter8, gate500inter9, gate500inter10, gate500inter11, gate500inter12, gate477inter0, gate477inter1, gate477inter2, gate477inter3, gate477inter4, gate477inter5, gate477inter6, gate477inter7, gate477inter8, gate477inter9, gate477inter10, gate477inter11, gate477inter12, gate264inter0, gate264inter1, gate264inter2, gate264inter3, gate264inter4, gate264inter5, gate264inter6, gate264inter7, gate264inter8, gate264inter9, gate264inter10, gate264inter11, gate264inter12, gate124inter0, gate124inter1, gate124inter2, gate124inter3, gate124inter4, gate124inter5, gate124inter6, gate124inter7, gate124inter8, gate124inter9, gate124inter10, gate124inter11, gate124inter12, gate101inter0, gate101inter1, gate101inter2, gate101inter3, gate101inter4, gate101inter5, gate101inter6, gate101inter7, gate101inter8, gate101inter9, gate101inter10, gate101inter11, gate101inter12, gate194inter0, gate194inter1, gate194inter2, gate194inter3, gate194inter4, gate194inter5, gate194inter6, gate194inter7, gate194inter8, gate194inter9, gate194inter10, gate194inter11, gate194inter12, gate267inter0, gate267inter1, gate267inter2, gate267inter3, gate267inter4, gate267inter5, gate267inter6, gate267inter7, gate267inter8, gate267inter9, gate267inter10, gate267inter11, gate267inter12, gate99inter0, gate99inter1, gate99inter2, gate99inter3, gate99inter4, gate99inter5, gate99inter6, gate99inter7, gate99inter8, gate99inter9, gate99inter10, gate99inter11, gate99inter12, gate260inter0, gate260inter1, gate260inter2, gate260inter3, gate260inter4, gate260inter5, gate260inter6, gate260inter7, gate260inter8, gate260inter9, gate260inter10, gate260inter11, gate260inter12, gate32inter0, gate32inter1, gate32inter2, gate32inter3, gate32inter4, gate32inter5, gate32inter6, gate32inter7, gate32inter8, gate32inter9, gate32inter10, gate32inter11, gate32inter12, gate213inter0, gate213inter1, gate213inter2, gate213inter3, gate213inter4, gate213inter5, gate213inter6, gate213inter7, gate213inter8, gate213inter9, gate213inter10, gate213inter11, gate213inter12, gate62inter0, gate62inter1, gate62inter2, gate62inter3, gate62inter4, gate62inter5, gate62inter6, gate62inter7, gate62inter8, gate62inter9, gate62inter10, gate62inter11, gate62inter12, gate21inter0, gate21inter1, gate21inter2, gate21inter3, gate21inter4, gate21inter5, gate21inter6, gate21inter7, gate21inter8, gate21inter9, gate21inter10, gate21inter11, gate21inter12, gate23inter0, gate23inter1, gate23inter2, gate23inter3, gate23inter4, gate23inter5, gate23inter6, gate23inter7, gate23inter8, gate23inter9, gate23inter10, gate23inter11, gate23inter12, gate273inter0, gate273inter1, gate273inter2, gate273inter3, gate273inter4, gate273inter5, gate273inter6, gate273inter7, gate273inter8, gate273inter9, gate273inter10, gate273inter11, gate273inter12, gate499inter0, gate499inter1, gate499inter2, gate499inter3, gate499inter4, gate499inter5, gate499inter6, gate499inter7, gate499inter8, gate499inter9, gate499inter10, gate499inter11, gate499inter12, gate56inter0, gate56inter1, gate56inter2, gate56inter3, gate56inter4, gate56inter5, gate56inter6, gate56inter7, gate56inter8, gate56inter9, gate56inter10, gate56inter11, gate56inter12, gate130inter0, gate130inter1, gate130inter2, gate130inter3, gate130inter4, gate130inter5, gate130inter6, gate130inter7, gate130inter8, gate130inter9, gate130inter10, gate130inter11, gate130inter12, gate417inter0, gate417inter1, gate417inter2, gate417inter3, gate417inter4, gate417inter5, gate417inter6, gate417inter7, gate417inter8, gate417inter9, gate417inter10, gate417inter11, gate417inter12, gate152inter0, gate152inter1, gate152inter2, gate152inter3, gate152inter4, gate152inter5, gate152inter6, gate152inter7, gate152inter8, gate152inter9, gate152inter10, gate152inter11, gate152inter12, gate463inter0, gate463inter1, gate463inter2, gate463inter3, gate463inter4, gate463inter5, gate463inter6, gate463inter7, gate463inter8, gate463inter9, gate463inter10, gate463inter11, gate463inter12, gate509inter0, gate509inter1, gate509inter2, gate509inter3, gate509inter4, gate509inter5, gate509inter6, gate509inter7, gate509inter8, gate509inter9, gate509inter10, gate509inter11, gate509inter12, gate292inter0, gate292inter1, gate292inter2, gate292inter3, gate292inter4, gate292inter5, gate292inter6, gate292inter7, gate292inter8, gate292inter9, gate292inter10, gate292inter11, gate292inter12, gate158inter0, gate158inter1, gate158inter2, gate158inter3, gate158inter4, gate158inter5, gate158inter6, gate158inter7, gate158inter8, gate158inter9, gate158inter10, gate158inter11, gate158inter12, gate59inter0, gate59inter1, gate59inter2, gate59inter3, gate59inter4, gate59inter5, gate59inter6, gate59inter7, gate59inter8, gate59inter9, gate59inter10, gate59inter11, gate59inter12, gate89inter0, gate89inter1, gate89inter2, gate89inter3, gate89inter4, gate89inter5, gate89inter6, gate89inter7, gate89inter8, gate89inter9, gate89inter10, gate89inter11, gate89inter12, gate39inter0, gate39inter1, gate39inter2, gate39inter3, gate39inter4, gate39inter5, gate39inter6, gate39inter7, gate39inter8, gate39inter9, gate39inter10, gate39inter11, gate39inter12, gate36inter0, gate36inter1, gate36inter2, gate36inter3, gate36inter4, gate36inter5, gate36inter6, gate36inter7, gate36inter8, gate36inter9, gate36inter10, gate36inter11, gate36inter12, gate427inter0, gate427inter1, gate427inter2, gate427inter3, gate427inter4, gate427inter5, gate427inter6, gate427inter7, gate427inter8, gate427inter9, gate427inter10, gate427inter11, gate427inter12, gate37inter0, gate37inter1, gate37inter2, gate37inter3, gate37inter4, gate37inter5, gate37inter6, gate37inter7, gate37inter8, gate37inter9, gate37inter10, gate37inter11, gate37inter12, gate388inter0, gate388inter1, gate388inter2, gate388inter3, gate388inter4, gate388inter5, gate388inter6, gate388inter7, gate388inter8, gate388inter9, gate388inter10, gate388inter11, gate388inter12, gate395inter0, gate395inter1, gate395inter2, gate395inter3, gate395inter4, gate395inter5, gate395inter6, gate395inter7, gate395inter8, gate395inter9, gate395inter10, gate395inter11, gate395inter12, gate195inter0, gate195inter1, gate195inter2, gate195inter3, gate195inter4, gate195inter5, gate195inter6, gate195inter7, gate195inter8, gate195inter9, gate195inter10, gate195inter11, gate195inter12, gate451inter0, gate451inter1, gate451inter2, gate451inter3, gate451inter4, gate451inter5, gate451inter6, gate451inter7, gate451inter8, gate451inter9, gate451inter10, gate451inter11, gate451inter12, gate467inter0, gate467inter1, gate467inter2, gate467inter3, gate467inter4, gate467inter5, gate467inter6, gate467inter7, gate467inter8, gate467inter9, gate467inter10, gate467inter11, gate467inter12, gate202inter0, gate202inter1, gate202inter2, gate202inter3, gate202inter4, gate202inter5, gate202inter6, gate202inter7, gate202inter8, gate202inter9, gate202inter10, gate202inter11, gate202inter12, gate409inter0, gate409inter1, gate409inter2, gate409inter3, gate409inter4, gate409inter5, gate409inter6, gate409inter7, gate409inter8, gate409inter9, gate409inter10, gate409inter11, gate409inter12, gate412inter0, gate412inter1, gate412inter2, gate412inter3, gate412inter4, gate412inter5, gate412inter6, gate412inter7, gate412inter8, gate412inter9, gate412inter10, gate412inter11, gate412inter12, gate411inter0, gate411inter1, gate411inter2, gate411inter3, gate411inter4, gate411inter5, gate411inter6, gate411inter7, gate411inter8, gate411inter9, gate411inter10, gate411inter11, gate411inter12, gate405inter0, gate405inter1, gate405inter2, gate405inter3, gate405inter4, gate405inter5, gate405inter6, gate405inter7, gate405inter8, gate405inter9, gate405inter10, gate405inter11, gate405inter12, gate286inter0, gate286inter1, gate286inter2, gate286inter3, gate286inter4, gate286inter5, gate286inter6, gate286inter7, gate286inter8, gate286inter9, gate286inter10, gate286inter11, gate286inter12, gate261inter0, gate261inter1, gate261inter2, gate261inter3, gate261inter4, gate261inter5, gate261inter6, gate261inter7, gate261inter8, gate261inter9, gate261inter10, gate261inter11, gate261inter12, gate174inter0, gate174inter1, gate174inter2, gate174inter3, gate174inter4, gate174inter5, gate174inter6, gate174inter7, gate174inter8, gate174inter9, gate174inter10, gate174inter11, gate174inter12, gate489inter0, gate489inter1, gate489inter2, gate489inter3, gate489inter4, gate489inter5, gate489inter6, gate489inter7, gate489inter8, gate489inter9, gate489inter10, gate489inter11, gate489inter12, gate33inter0, gate33inter1, gate33inter2, gate33inter3, gate33inter4, gate33inter5, gate33inter6, gate33inter7, gate33inter8, gate33inter9, gate33inter10, gate33inter11, gate33inter12, gate187inter0, gate187inter1, gate187inter2, gate187inter3, gate187inter4, gate187inter5, gate187inter6, gate187inter7, gate187inter8, gate187inter9, gate187inter10, gate187inter11, gate187inter12, gate484inter0, gate484inter1, gate484inter2, gate484inter3, gate484inter4, gate484inter5, gate484inter6, gate484inter7, gate484inter8, gate484inter9, gate484inter10, gate484inter11, gate484inter12, gate248inter0, gate248inter1, gate248inter2, gate248inter3, gate248inter4, gate248inter5, gate248inter6, gate248inter7, gate248inter8, gate248inter9, gate248inter10, gate248inter11, gate248inter12, gate291inter0, gate291inter1, gate291inter2, gate291inter3, gate291inter4, gate291inter5, gate291inter6, gate291inter7, gate291inter8, gate291inter9, gate291inter10, gate291inter11, gate291inter12, gate86inter0, gate86inter1, gate86inter2, gate86inter3, gate86inter4, gate86inter5, gate86inter6, gate86inter7, gate86inter8, gate86inter9, gate86inter10, gate86inter11, gate86inter12, gate240inter0, gate240inter1, gate240inter2, gate240inter3, gate240inter4, gate240inter5, gate240inter6, gate240inter7, gate240inter8, gate240inter9, gate240inter10, gate240inter11, gate240inter12, gate470inter0, gate470inter1, gate470inter2, gate470inter3, gate470inter4, gate470inter5, gate470inter6, gate470inter7, gate470inter8, gate470inter9, gate470inter10, gate470inter11, gate470inter12, gate407inter0, gate407inter1, gate407inter2, gate407inter3, gate407inter4, gate407inter5, gate407inter6, gate407inter7, gate407inter8, gate407inter9, gate407inter10, gate407inter11, gate407inter12, gate437inter0, gate437inter1, gate437inter2, gate437inter3, gate437inter4, gate437inter5, gate437inter6, gate437inter7, gate437inter8, gate437inter9, gate437inter10, gate437inter11, gate437inter12, gate247inter0, gate247inter1, gate247inter2, gate247inter3, gate247inter4, gate247inter5, gate247inter6, gate247inter7, gate247inter8, gate247inter9, gate247inter10, gate247inter11, gate247inter12, gate182inter0, gate182inter1, gate182inter2, gate182inter3, gate182inter4, gate182inter5, gate182inter6, gate182inter7, gate182inter8, gate182inter9, gate182inter10, gate182inter11, gate182inter12, gate51inter0, gate51inter1, gate51inter2, gate51inter3, gate51inter4, gate51inter5, gate51inter6, gate51inter7, gate51inter8, gate51inter9, gate51inter10, gate51inter11, gate51inter12, gate178inter0, gate178inter1, gate178inter2, gate178inter3, gate178inter4, gate178inter5, gate178inter6, gate178inter7, gate178inter8, gate178inter9, gate178inter10, gate178inter11, gate178inter12, gate415inter0, gate415inter1, gate415inter2, gate415inter3, gate415inter4, gate415inter5, gate415inter6, gate415inter7, gate415inter8, gate415inter9, gate415inter10, gate415inter11, gate415inter12, gate508inter0, gate508inter1, gate508inter2, gate508inter3, gate508inter4, gate508inter5, gate508inter6, gate508inter7, gate508inter8, gate508inter9, gate508inter10, gate508inter11, gate508inter12, gate14inter0, gate14inter1, gate14inter2, gate14inter3, gate14inter4, gate14inter5, gate14inter6, gate14inter7, gate14inter8, gate14inter9, gate14inter10, gate14inter11, gate14inter12, gate250inter0, gate250inter1, gate250inter2, gate250inter3, gate250inter4, gate250inter5, gate250inter6, gate250inter7, gate250inter8, gate250inter9, gate250inter10, gate250inter11, gate250inter12, gate488inter0, gate488inter1, gate488inter2, gate488inter3, gate488inter4, gate488inter5, gate488inter6, gate488inter7, gate488inter8, gate488inter9, gate488inter10, gate488inter11, gate488inter12, gate436inter0, gate436inter1, gate436inter2, gate436inter3, gate436inter4, gate436inter5, gate436inter6, gate436inter7, gate436inter8, gate436inter9, gate436inter10, gate436inter11, gate436inter12, gate44inter0, gate44inter1, gate44inter2, gate44inter3, gate44inter4, gate44inter5, gate44inter6, gate44inter7, gate44inter8, gate44inter9, gate44inter10, gate44inter11, gate44inter12, gate438inter0, gate438inter1, gate438inter2, gate438inter3, gate438inter4, gate438inter5, gate438inter6, gate438inter7, gate438inter8, gate438inter9, gate438inter10, gate438inter11, gate438inter12, gate227inter0, gate227inter1, gate227inter2, gate227inter3, gate227inter4, gate227inter5, gate227inter6, gate227inter7, gate227inter8, gate227inter9, gate227inter10, gate227inter11, gate227inter12, gate251inter0, gate251inter1, gate251inter2, gate251inter3, gate251inter4, gate251inter5, gate251inter6, gate251inter7, gate251inter8, gate251inter9, gate251inter10, gate251inter11, gate251inter12, gate19inter0, gate19inter1, gate19inter2, gate19inter3, gate19inter4, gate19inter5, gate19inter6, gate19inter7, gate19inter8, gate19inter9, gate19inter10, gate19inter11, gate19inter12, gate77inter0, gate77inter1, gate77inter2, gate77inter3, gate77inter4, gate77inter5, gate77inter6, gate77inter7, gate77inter8, gate77inter9, gate77inter10, gate77inter11, gate77inter12, gate465inter0, gate465inter1, gate465inter2, gate465inter3, gate465inter4, gate465inter5, gate465inter6, gate465inter7, gate465inter8, gate465inter9, gate465inter10, gate465inter11, gate465inter12, gate80inter0, gate80inter1, gate80inter2, gate80inter3, gate80inter4, gate80inter5, gate80inter6, gate80inter7, gate80inter8, gate80inter9, gate80inter10, gate80inter11, gate80inter12, gate208inter0, gate208inter1, gate208inter2, gate208inter3, gate208inter4, gate208inter5, gate208inter6, gate208inter7, gate208inter8, gate208inter9, gate208inter10, gate208inter11, gate208inter12, gate66inter0, gate66inter1, gate66inter2, gate66inter3, gate66inter4, gate66inter5, gate66inter6, gate66inter7, gate66inter8, gate66inter9, gate66inter10, gate66inter11, gate66inter12, gate220inter0, gate220inter1, gate220inter2, gate220inter3, gate220inter4, gate220inter5, gate220inter6, gate220inter7, gate220inter8, gate220inter9, gate220inter10, gate220inter11, gate220inter12, gate256inter0, gate256inter1, gate256inter2, gate256inter3, gate256inter4, gate256inter5, gate256inter6, gate256inter7, gate256inter8, gate256inter9, gate256inter10, gate256inter11, gate256inter12, gate54inter0, gate54inter1, gate54inter2, gate54inter3, gate54inter4, gate54inter5, gate54inter6, gate54inter7, gate54inter8, gate54inter9, gate54inter10, gate54inter11, gate54inter12, gate201inter0, gate201inter1, gate201inter2, gate201inter3, gate201inter4, gate201inter5, gate201inter6, gate201inter7, gate201inter8, gate201inter9, gate201inter10, gate201inter11, gate201inter12, gate433inter0, gate433inter1, gate433inter2, gate433inter3, gate433inter4, gate433inter5, gate433inter6, gate433inter7, gate433inter8, gate433inter9, gate433inter10, gate433inter11, gate433inter12, gate279inter0, gate279inter1, gate279inter2, gate279inter3, gate279inter4, gate279inter5, gate279inter6, gate279inter7, gate279inter8, gate279inter9, gate279inter10, gate279inter11, gate279inter12, gate191inter0, gate191inter1, gate191inter2, gate191inter3, gate191inter4, gate191inter5, gate191inter6, gate191inter7, gate191inter8, gate191inter9, gate191inter10, gate191inter11, gate191inter12, gate239inter0, gate239inter1, gate239inter2, gate239inter3, gate239inter4, gate239inter5, gate239inter6, gate239inter7, gate239inter8, gate239inter9, gate239inter10, gate239inter11, gate239inter12, gate70inter0, gate70inter1, gate70inter2, gate70inter3, gate70inter4, gate70inter5, gate70inter6, gate70inter7, gate70inter8, gate70inter9, gate70inter10, gate70inter11, gate70inter12, gate453inter0, gate453inter1, gate453inter2, gate453inter3, gate453inter4, gate453inter5, gate453inter6, gate453inter7, gate453inter8, gate453inter9, gate453inter10, gate453inter11, gate453inter12, gate140inter0, gate140inter1, gate140inter2, gate140inter3, gate140inter4, gate140inter5, gate140inter6, gate140inter7, gate140inter8, gate140inter9, gate140inter10, gate140inter11, gate140inter12, gate408inter0, gate408inter1, gate408inter2, gate408inter3, gate408inter4, gate408inter5, gate408inter6, gate408inter7, gate408inter8, gate408inter9, gate408inter10, gate408inter11, gate408inter12, gate146inter0, gate146inter1, gate146inter2, gate146inter3, gate146inter4, gate146inter5, gate146inter6, gate146inter7, gate146inter8, gate146inter9, gate146inter10, gate146inter11, gate146inter12, gate295inter0, gate295inter1, gate295inter2, gate295inter3, gate295inter4, gate295inter5, gate295inter6, gate295inter7, gate295inter8, gate295inter9, gate295inter10, gate295inter11, gate295inter12, gate416inter0, gate416inter1, gate416inter2, gate416inter3, gate416inter4, gate416inter5, gate416inter6, gate416inter7, gate416inter8, gate416inter9, gate416inter10, gate416inter11, gate416inter12, gate122inter0, gate122inter1, gate122inter2, gate122inter3, gate122inter4, gate122inter5, gate122inter6, gate122inter7, gate122inter8, gate122inter9, gate122inter10, gate122inter11, gate122inter12, gate169inter0, gate169inter1, gate169inter2, gate169inter3, gate169inter4, gate169inter5, gate169inter6, gate169inter7, gate169inter8, gate169inter9, gate169inter10, gate169inter11, gate169inter12, gate148inter0, gate148inter1, gate148inter2, gate148inter3, gate148inter4, gate148inter5, gate148inter6, gate148inter7, gate148inter8, gate148inter9, gate148inter10, gate148inter11, gate148inter12, gate434inter0, gate434inter1, gate434inter2, gate434inter3, gate434inter4, gate434inter5, gate434inter6, gate434inter7, gate434inter8, gate434inter9, gate434inter10, gate434inter11, gate434inter12, gate18inter0, gate18inter1, gate18inter2, gate18inter3, gate18inter4, gate18inter5, gate18inter6, gate18inter7, gate18inter8, gate18inter9, gate18inter10, gate18inter11, gate18inter12, gate390inter0, gate390inter1, gate390inter2, gate390inter3, gate390inter4, gate390inter5, gate390inter6, gate390inter7, gate390inter8, gate390inter9, gate390inter10, gate390inter11, gate390inter12, gate472inter0, gate472inter1, gate472inter2, gate472inter3, gate472inter4, gate472inter5, gate472inter6, gate472inter7, gate472inter8, gate472inter9, gate472inter10, gate472inter11, gate472inter12, gate263inter0, gate263inter1, gate263inter2, gate263inter3, gate263inter4, gate263inter5, gate263inter6, gate263inter7, gate263inter8, gate263inter9, gate263inter10, gate263inter11, gate263inter12, gate426inter0, gate426inter1, gate426inter2, gate426inter3, gate426inter4, gate426inter5, gate426inter6, gate426inter7, gate426inter8, gate426inter9, gate426inter10, gate426inter11, gate426inter12, gate218inter0, gate218inter1, gate218inter2, gate218inter3, gate218inter4, gate218inter5, gate218inter6, gate218inter7, gate218inter8, gate218inter9, gate218inter10, gate218inter11, gate218inter12, gate34inter0, gate34inter1, gate34inter2, gate34inter3, gate34inter4, gate34inter5, gate34inter6, gate34inter7, gate34inter8, gate34inter9, gate34inter10, gate34inter11, gate34inter12, gate121inter0, gate121inter1, gate121inter2, gate121inter3, gate121inter4, gate121inter5, gate121inter6, gate121inter7, gate121inter8, gate121inter9, gate121inter10, gate121inter11, gate121inter12, gate186inter0, gate186inter1, gate186inter2, gate186inter3, gate186inter4, gate186inter5, gate186inter6, gate186inter7, gate186inter8, gate186inter9, gate186inter10, gate186inter11, gate186inter12, gate514inter0, gate514inter1, gate514inter2, gate514inter3, gate514inter4, gate514inter5, gate514inter6, gate514inter7, gate514inter8, gate514inter9, gate514inter10, gate514inter11, gate514inter12, gate278inter0, gate278inter1, gate278inter2, gate278inter3, gate278inter4, gate278inter5, gate278inter6, gate278inter7, gate278inter8, gate278inter9, gate278inter10, gate278inter11, gate278inter12, gate406inter0, gate406inter1, gate406inter2, gate406inter3, gate406inter4, gate406inter5, gate406inter6, gate406inter7, gate406inter8, gate406inter9, gate406inter10, gate406inter11, gate406inter12, gate252inter0, gate252inter1, gate252inter2, gate252inter3, gate252inter4, gate252inter5, gate252inter6, gate252inter7, gate252inter8, gate252inter9, gate252inter10, gate252inter11, gate252inter12, gate271inter0, gate271inter1, gate271inter2, gate271inter3, gate271inter4, gate271inter5, gate271inter6, gate271inter7, gate271inter8, gate271inter9, gate271inter10, gate271inter11, gate271inter12, gate175inter0, gate175inter1, gate175inter2, gate175inter3, gate175inter4, gate175inter5, gate175inter6, gate175inter7, gate175inter8, gate175inter9, gate175inter10, gate175inter11, gate175inter12, gate274inter0, gate274inter1, gate274inter2, gate274inter3, gate274inter4, gate274inter5, gate274inter6, gate274inter7, gate274inter8, gate274inter9, gate274inter10, gate274inter11, gate274inter12;



and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );
nand2 gate9( .a(G1), .b(G2), .O(G266) );
nand2 gate10( .a(G3), .b(G4), .O(G269) );
nand2 gate11( .a(G5), .b(G6), .O(G272) );
nand2 gate12( .a(G7), .b(G8), .O(G275) );
nand2 gate13( .a(G9), .b(G10), .O(G278) );

  xor2  gate1485(.a(G12), .b(G11), .O(gate14inter0));
  nand2 gate1486(.a(gate14inter0), .b(s_134), .O(gate14inter1));
  and2  gate1487(.a(G12), .b(G11), .O(gate14inter2));
  inv1  gate1488(.a(s_134), .O(gate14inter3));
  inv1  gate1489(.a(s_135), .O(gate14inter4));
  nand2 gate1490(.a(gate14inter4), .b(gate14inter3), .O(gate14inter5));
  nor2  gate1491(.a(gate14inter5), .b(gate14inter2), .O(gate14inter6));
  inv1  gate1492(.a(G11), .O(gate14inter7));
  inv1  gate1493(.a(G12), .O(gate14inter8));
  nand2 gate1494(.a(gate14inter8), .b(gate14inter7), .O(gate14inter9));
  nand2 gate1495(.a(s_135), .b(gate14inter3), .O(gate14inter10));
  nor2  gate1496(.a(gate14inter10), .b(gate14inter9), .O(gate14inter11));
  nor2  gate1497(.a(gate14inter11), .b(gate14inter6), .O(gate14inter12));
  nand2 gate1498(.a(gate14inter12), .b(gate14inter1), .O(G281));
nand2 gate15( .a(G13), .b(G14), .O(G284) );
nand2 gate16( .a(G15), .b(G16), .O(G287) );
nand2 gate17( .a(G17), .b(G18), .O(G290) );

  xor2  gate1947(.a(G20), .b(G19), .O(gate18inter0));
  nand2 gate1948(.a(gate18inter0), .b(s_200), .O(gate18inter1));
  and2  gate1949(.a(G20), .b(G19), .O(gate18inter2));
  inv1  gate1950(.a(s_200), .O(gate18inter3));
  inv1  gate1951(.a(s_201), .O(gate18inter4));
  nand2 gate1952(.a(gate18inter4), .b(gate18inter3), .O(gate18inter5));
  nor2  gate1953(.a(gate18inter5), .b(gate18inter2), .O(gate18inter6));
  inv1  gate1954(.a(G19), .O(gate18inter7));
  inv1  gate1955(.a(G20), .O(gate18inter8));
  nand2 gate1956(.a(gate18inter8), .b(gate18inter7), .O(gate18inter9));
  nand2 gate1957(.a(s_201), .b(gate18inter3), .O(gate18inter10));
  nor2  gate1958(.a(gate18inter10), .b(gate18inter9), .O(gate18inter11));
  nor2  gate1959(.a(gate18inter11), .b(gate18inter6), .O(gate18inter12));
  nand2 gate1960(.a(gate18inter12), .b(gate18inter1), .O(G293));

  xor2  gate1597(.a(G22), .b(G21), .O(gate19inter0));
  nand2 gate1598(.a(gate19inter0), .b(s_150), .O(gate19inter1));
  and2  gate1599(.a(G22), .b(G21), .O(gate19inter2));
  inv1  gate1600(.a(s_150), .O(gate19inter3));
  inv1  gate1601(.a(s_151), .O(gate19inter4));
  nand2 gate1602(.a(gate19inter4), .b(gate19inter3), .O(gate19inter5));
  nor2  gate1603(.a(gate19inter5), .b(gate19inter2), .O(gate19inter6));
  inv1  gate1604(.a(G21), .O(gate19inter7));
  inv1  gate1605(.a(G22), .O(gate19inter8));
  nand2 gate1606(.a(gate19inter8), .b(gate19inter7), .O(gate19inter9));
  nand2 gate1607(.a(s_151), .b(gate19inter3), .O(gate19inter10));
  nor2  gate1608(.a(gate19inter10), .b(gate19inter9), .O(gate19inter11));
  nor2  gate1609(.a(gate19inter11), .b(gate19inter6), .O(gate19inter12));
  nand2 gate1610(.a(gate19inter12), .b(gate19inter1), .O(G296));
nand2 gate20( .a(G23), .b(G24), .O(G299) );

  xor2  gate813(.a(G26), .b(G25), .O(gate21inter0));
  nand2 gate814(.a(gate21inter0), .b(s_38), .O(gate21inter1));
  and2  gate815(.a(G26), .b(G25), .O(gate21inter2));
  inv1  gate816(.a(s_38), .O(gate21inter3));
  inv1  gate817(.a(s_39), .O(gate21inter4));
  nand2 gate818(.a(gate21inter4), .b(gate21inter3), .O(gate21inter5));
  nor2  gate819(.a(gate21inter5), .b(gate21inter2), .O(gate21inter6));
  inv1  gate820(.a(G25), .O(gate21inter7));
  inv1  gate821(.a(G26), .O(gate21inter8));
  nand2 gate822(.a(gate21inter8), .b(gate21inter7), .O(gate21inter9));
  nand2 gate823(.a(s_39), .b(gate21inter3), .O(gate21inter10));
  nor2  gate824(.a(gate21inter10), .b(gate21inter9), .O(gate21inter11));
  nor2  gate825(.a(gate21inter11), .b(gate21inter6), .O(gate21inter12));
  nand2 gate826(.a(gate21inter12), .b(gate21inter1), .O(G302));
nand2 gate22( .a(G27), .b(G28), .O(G305) );

  xor2  gate827(.a(G30), .b(G29), .O(gate23inter0));
  nand2 gate828(.a(gate23inter0), .b(s_40), .O(gate23inter1));
  and2  gate829(.a(G30), .b(G29), .O(gate23inter2));
  inv1  gate830(.a(s_40), .O(gate23inter3));
  inv1  gate831(.a(s_41), .O(gate23inter4));
  nand2 gate832(.a(gate23inter4), .b(gate23inter3), .O(gate23inter5));
  nor2  gate833(.a(gate23inter5), .b(gate23inter2), .O(gate23inter6));
  inv1  gate834(.a(G29), .O(gate23inter7));
  inv1  gate835(.a(G30), .O(gate23inter8));
  nand2 gate836(.a(gate23inter8), .b(gate23inter7), .O(gate23inter9));
  nand2 gate837(.a(s_41), .b(gate23inter3), .O(gate23inter10));
  nor2  gate838(.a(gate23inter10), .b(gate23inter9), .O(gate23inter11));
  nor2  gate839(.a(gate23inter11), .b(gate23inter6), .O(gate23inter12));
  nand2 gate840(.a(gate23inter12), .b(gate23inter1), .O(G308));
nand2 gate24( .a(G31), .b(G32), .O(G311) );
nand2 gate25( .a(G1), .b(G5), .O(G314) );
nand2 gate26( .a(G9), .b(G13), .O(G317) );
nand2 gate27( .a(G2), .b(G6), .O(G320) );
nand2 gate28( .a(G10), .b(G14), .O(G323) );

  xor2  gate617(.a(G7), .b(G3), .O(gate29inter0));
  nand2 gate618(.a(gate29inter0), .b(s_10), .O(gate29inter1));
  and2  gate619(.a(G7), .b(G3), .O(gate29inter2));
  inv1  gate620(.a(s_10), .O(gate29inter3));
  inv1  gate621(.a(s_11), .O(gate29inter4));
  nand2 gate622(.a(gate29inter4), .b(gate29inter3), .O(gate29inter5));
  nor2  gate623(.a(gate29inter5), .b(gate29inter2), .O(gate29inter6));
  inv1  gate624(.a(G3), .O(gate29inter7));
  inv1  gate625(.a(G7), .O(gate29inter8));
  nand2 gate626(.a(gate29inter8), .b(gate29inter7), .O(gate29inter9));
  nand2 gate627(.a(s_11), .b(gate29inter3), .O(gate29inter10));
  nor2  gate628(.a(gate29inter10), .b(gate29inter9), .O(gate29inter11));
  nor2  gate629(.a(gate29inter11), .b(gate29inter6), .O(gate29inter12));
  nand2 gate630(.a(gate29inter12), .b(gate29inter1), .O(G326));
nand2 gate30( .a(G11), .b(G15), .O(G329) );
nand2 gate31( .a(G4), .b(G8), .O(G332) );

  xor2  gate771(.a(G16), .b(G12), .O(gate32inter0));
  nand2 gate772(.a(gate32inter0), .b(s_32), .O(gate32inter1));
  and2  gate773(.a(G16), .b(G12), .O(gate32inter2));
  inv1  gate774(.a(s_32), .O(gate32inter3));
  inv1  gate775(.a(s_33), .O(gate32inter4));
  nand2 gate776(.a(gate32inter4), .b(gate32inter3), .O(gate32inter5));
  nor2  gate777(.a(gate32inter5), .b(gate32inter2), .O(gate32inter6));
  inv1  gate778(.a(G12), .O(gate32inter7));
  inv1  gate779(.a(G16), .O(gate32inter8));
  nand2 gate780(.a(gate32inter8), .b(gate32inter7), .O(gate32inter9));
  nand2 gate781(.a(s_33), .b(gate32inter3), .O(gate32inter10));
  nor2  gate782(.a(gate32inter10), .b(gate32inter9), .O(gate32inter11));
  nor2  gate783(.a(gate32inter11), .b(gate32inter6), .O(gate32inter12));
  nand2 gate784(.a(gate32inter12), .b(gate32inter1), .O(G335));

  xor2  gate1261(.a(G21), .b(G17), .O(gate33inter0));
  nand2 gate1262(.a(gate33inter0), .b(s_102), .O(gate33inter1));
  and2  gate1263(.a(G21), .b(G17), .O(gate33inter2));
  inv1  gate1264(.a(s_102), .O(gate33inter3));
  inv1  gate1265(.a(s_103), .O(gate33inter4));
  nand2 gate1266(.a(gate33inter4), .b(gate33inter3), .O(gate33inter5));
  nor2  gate1267(.a(gate33inter5), .b(gate33inter2), .O(gate33inter6));
  inv1  gate1268(.a(G17), .O(gate33inter7));
  inv1  gate1269(.a(G21), .O(gate33inter8));
  nand2 gate1270(.a(gate33inter8), .b(gate33inter7), .O(gate33inter9));
  nand2 gate1271(.a(s_103), .b(gate33inter3), .O(gate33inter10));
  nor2  gate1272(.a(gate33inter10), .b(gate33inter9), .O(gate33inter11));
  nor2  gate1273(.a(gate33inter11), .b(gate33inter6), .O(gate33inter12));
  nand2 gate1274(.a(gate33inter12), .b(gate33inter1), .O(G338));

  xor2  gate2031(.a(G29), .b(G25), .O(gate34inter0));
  nand2 gate2032(.a(gate34inter0), .b(s_212), .O(gate34inter1));
  and2  gate2033(.a(G29), .b(G25), .O(gate34inter2));
  inv1  gate2034(.a(s_212), .O(gate34inter3));
  inv1  gate2035(.a(s_213), .O(gate34inter4));
  nand2 gate2036(.a(gate34inter4), .b(gate34inter3), .O(gate34inter5));
  nor2  gate2037(.a(gate34inter5), .b(gate34inter2), .O(gate34inter6));
  inv1  gate2038(.a(G25), .O(gate34inter7));
  inv1  gate2039(.a(G29), .O(gate34inter8));
  nand2 gate2040(.a(gate34inter8), .b(gate34inter7), .O(gate34inter9));
  nand2 gate2041(.a(s_213), .b(gate34inter3), .O(gate34inter10));
  nor2  gate2042(.a(gate34inter10), .b(gate34inter9), .O(gate34inter11));
  nor2  gate2043(.a(gate34inter11), .b(gate34inter6), .O(gate34inter12));
  nand2 gate2044(.a(gate34inter12), .b(gate34inter1), .O(G341));
nand2 gate35( .a(G18), .b(G22), .O(G344) );

  xor2  gate1023(.a(G30), .b(G26), .O(gate36inter0));
  nand2 gate1024(.a(gate36inter0), .b(s_68), .O(gate36inter1));
  and2  gate1025(.a(G30), .b(G26), .O(gate36inter2));
  inv1  gate1026(.a(s_68), .O(gate36inter3));
  inv1  gate1027(.a(s_69), .O(gate36inter4));
  nand2 gate1028(.a(gate36inter4), .b(gate36inter3), .O(gate36inter5));
  nor2  gate1029(.a(gate36inter5), .b(gate36inter2), .O(gate36inter6));
  inv1  gate1030(.a(G26), .O(gate36inter7));
  inv1  gate1031(.a(G30), .O(gate36inter8));
  nand2 gate1032(.a(gate36inter8), .b(gate36inter7), .O(gate36inter9));
  nand2 gate1033(.a(s_69), .b(gate36inter3), .O(gate36inter10));
  nor2  gate1034(.a(gate36inter10), .b(gate36inter9), .O(gate36inter11));
  nor2  gate1035(.a(gate36inter11), .b(gate36inter6), .O(gate36inter12));
  nand2 gate1036(.a(gate36inter12), .b(gate36inter1), .O(G347));

  xor2  gate1051(.a(G23), .b(G19), .O(gate37inter0));
  nand2 gate1052(.a(gate37inter0), .b(s_72), .O(gate37inter1));
  and2  gate1053(.a(G23), .b(G19), .O(gate37inter2));
  inv1  gate1054(.a(s_72), .O(gate37inter3));
  inv1  gate1055(.a(s_73), .O(gate37inter4));
  nand2 gate1056(.a(gate37inter4), .b(gate37inter3), .O(gate37inter5));
  nor2  gate1057(.a(gate37inter5), .b(gate37inter2), .O(gate37inter6));
  inv1  gate1058(.a(G19), .O(gate37inter7));
  inv1  gate1059(.a(G23), .O(gate37inter8));
  nand2 gate1060(.a(gate37inter8), .b(gate37inter7), .O(gate37inter9));
  nand2 gate1061(.a(s_73), .b(gate37inter3), .O(gate37inter10));
  nor2  gate1062(.a(gate37inter10), .b(gate37inter9), .O(gate37inter11));
  nor2  gate1063(.a(gate37inter11), .b(gate37inter6), .O(gate37inter12));
  nand2 gate1064(.a(gate37inter12), .b(gate37inter1), .O(G350));
nand2 gate38( .a(G27), .b(G31), .O(G353) );

  xor2  gate1009(.a(G24), .b(G20), .O(gate39inter0));
  nand2 gate1010(.a(gate39inter0), .b(s_66), .O(gate39inter1));
  and2  gate1011(.a(G24), .b(G20), .O(gate39inter2));
  inv1  gate1012(.a(s_66), .O(gate39inter3));
  inv1  gate1013(.a(s_67), .O(gate39inter4));
  nand2 gate1014(.a(gate39inter4), .b(gate39inter3), .O(gate39inter5));
  nor2  gate1015(.a(gate39inter5), .b(gate39inter2), .O(gate39inter6));
  inv1  gate1016(.a(G20), .O(gate39inter7));
  inv1  gate1017(.a(G24), .O(gate39inter8));
  nand2 gate1018(.a(gate39inter8), .b(gate39inter7), .O(gate39inter9));
  nand2 gate1019(.a(s_67), .b(gate39inter3), .O(gate39inter10));
  nor2  gate1020(.a(gate39inter10), .b(gate39inter9), .O(gate39inter11));
  nor2  gate1021(.a(gate39inter11), .b(gate39inter6), .O(gate39inter12));
  nand2 gate1022(.a(gate39inter12), .b(gate39inter1), .O(G356));
nand2 gate40( .a(G28), .b(G32), .O(G359) );
nand2 gate41( .a(G1), .b(G266), .O(G362) );
nand2 gate42( .a(G2), .b(G266), .O(G363) );
nand2 gate43( .a(G3), .b(G269), .O(G364) );

  xor2  gate1541(.a(G269), .b(G4), .O(gate44inter0));
  nand2 gate1542(.a(gate44inter0), .b(s_142), .O(gate44inter1));
  and2  gate1543(.a(G269), .b(G4), .O(gate44inter2));
  inv1  gate1544(.a(s_142), .O(gate44inter3));
  inv1  gate1545(.a(s_143), .O(gate44inter4));
  nand2 gate1546(.a(gate44inter4), .b(gate44inter3), .O(gate44inter5));
  nor2  gate1547(.a(gate44inter5), .b(gate44inter2), .O(gate44inter6));
  inv1  gate1548(.a(G4), .O(gate44inter7));
  inv1  gate1549(.a(G269), .O(gate44inter8));
  nand2 gate1550(.a(gate44inter8), .b(gate44inter7), .O(gate44inter9));
  nand2 gate1551(.a(s_143), .b(gate44inter3), .O(gate44inter10));
  nor2  gate1552(.a(gate44inter10), .b(gate44inter9), .O(gate44inter11));
  nor2  gate1553(.a(gate44inter11), .b(gate44inter6), .O(gate44inter12));
  nand2 gate1554(.a(gate44inter12), .b(gate44inter1), .O(G365));
nand2 gate45( .a(G5), .b(G272), .O(G366) );
nand2 gate46( .a(G6), .b(G272), .O(G367) );
nand2 gate47( .a(G7), .b(G275), .O(G368) );
nand2 gate48( .a(G8), .b(G275), .O(G369) );
nand2 gate49( .a(G9), .b(G278), .O(G370) );
nand2 gate50( .a(G10), .b(G278), .O(G371) );

  xor2  gate1429(.a(G281), .b(G11), .O(gate51inter0));
  nand2 gate1430(.a(gate51inter0), .b(s_126), .O(gate51inter1));
  and2  gate1431(.a(G281), .b(G11), .O(gate51inter2));
  inv1  gate1432(.a(s_126), .O(gate51inter3));
  inv1  gate1433(.a(s_127), .O(gate51inter4));
  nand2 gate1434(.a(gate51inter4), .b(gate51inter3), .O(gate51inter5));
  nor2  gate1435(.a(gate51inter5), .b(gate51inter2), .O(gate51inter6));
  inv1  gate1436(.a(G11), .O(gate51inter7));
  inv1  gate1437(.a(G281), .O(gate51inter8));
  nand2 gate1438(.a(gate51inter8), .b(gate51inter7), .O(gate51inter9));
  nand2 gate1439(.a(s_127), .b(gate51inter3), .O(gate51inter10));
  nor2  gate1440(.a(gate51inter10), .b(gate51inter9), .O(gate51inter11));
  nor2  gate1441(.a(gate51inter11), .b(gate51inter6), .O(gate51inter12));
  nand2 gate1442(.a(gate51inter12), .b(gate51inter1), .O(G372));
nand2 gate52( .a(G12), .b(G281), .O(G373) );
nand2 gate53( .a(G13), .b(G284), .O(G374) );

  xor2  gate1709(.a(G284), .b(G14), .O(gate54inter0));
  nand2 gate1710(.a(gate54inter0), .b(s_166), .O(gate54inter1));
  and2  gate1711(.a(G284), .b(G14), .O(gate54inter2));
  inv1  gate1712(.a(s_166), .O(gate54inter3));
  inv1  gate1713(.a(s_167), .O(gate54inter4));
  nand2 gate1714(.a(gate54inter4), .b(gate54inter3), .O(gate54inter5));
  nor2  gate1715(.a(gate54inter5), .b(gate54inter2), .O(gate54inter6));
  inv1  gate1716(.a(G14), .O(gate54inter7));
  inv1  gate1717(.a(G284), .O(gate54inter8));
  nand2 gate1718(.a(gate54inter8), .b(gate54inter7), .O(gate54inter9));
  nand2 gate1719(.a(s_167), .b(gate54inter3), .O(gate54inter10));
  nor2  gate1720(.a(gate54inter10), .b(gate54inter9), .O(gate54inter11));
  nor2  gate1721(.a(gate54inter11), .b(gate54inter6), .O(gate54inter12));
  nand2 gate1722(.a(gate54inter12), .b(gate54inter1), .O(G375));
nand2 gate55( .a(G15), .b(G287), .O(G376) );

  xor2  gate869(.a(G287), .b(G16), .O(gate56inter0));
  nand2 gate870(.a(gate56inter0), .b(s_46), .O(gate56inter1));
  and2  gate871(.a(G287), .b(G16), .O(gate56inter2));
  inv1  gate872(.a(s_46), .O(gate56inter3));
  inv1  gate873(.a(s_47), .O(gate56inter4));
  nand2 gate874(.a(gate56inter4), .b(gate56inter3), .O(gate56inter5));
  nor2  gate875(.a(gate56inter5), .b(gate56inter2), .O(gate56inter6));
  inv1  gate876(.a(G16), .O(gate56inter7));
  inv1  gate877(.a(G287), .O(gate56inter8));
  nand2 gate878(.a(gate56inter8), .b(gate56inter7), .O(gate56inter9));
  nand2 gate879(.a(s_47), .b(gate56inter3), .O(gate56inter10));
  nor2  gate880(.a(gate56inter10), .b(gate56inter9), .O(gate56inter11));
  nor2  gate881(.a(gate56inter11), .b(gate56inter6), .O(gate56inter12));
  nand2 gate882(.a(gate56inter12), .b(gate56inter1), .O(G377));
nand2 gate57( .a(G17), .b(G290), .O(G378) );
nand2 gate58( .a(G18), .b(G290), .O(G379) );

  xor2  gate981(.a(G293), .b(G19), .O(gate59inter0));
  nand2 gate982(.a(gate59inter0), .b(s_62), .O(gate59inter1));
  and2  gate983(.a(G293), .b(G19), .O(gate59inter2));
  inv1  gate984(.a(s_62), .O(gate59inter3));
  inv1  gate985(.a(s_63), .O(gate59inter4));
  nand2 gate986(.a(gate59inter4), .b(gate59inter3), .O(gate59inter5));
  nor2  gate987(.a(gate59inter5), .b(gate59inter2), .O(gate59inter6));
  inv1  gate988(.a(G19), .O(gate59inter7));
  inv1  gate989(.a(G293), .O(gate59inter8));
  nand2 gate990(.a(gate59inter8), .b(gate59inter7), .O(gate59inter9));
  nand2 gate991(.a(s_63), .b(gate59inter3), .O(gate59inter10));
  nor2  gate992(.a(gate59inter10), .b(gate59inter9), .O(gate59inter11));
  nor2  gate993(.a(gate59inter11), .b(gate59inter6), .O(gate59inter12));
  nand2 gate994(.a(gate59inter12), .b(gate59inter1), .O(G380));
nand2 gate60( .a(G20), .b(G293), .O(G381) );
nand2 gate61( .a(G21), .b(G296), .O(G382) );

  xor2  gate799(.a(G296), .b(G22), .O(gate62inter0));
  nand2 gate800(.a(gate62inter0), .b(s_36), .O(gate62inter1));
  and2  gate801(.a(G296), .b(G22), .O(gate62inter2));
  inv1  gate802(.a(s_36), .O(gate62inter3));
  inv1  gate803(.a(s_37), .O(gate62inter4));
  nand2 gate804(.a(gate62inter4), .b(gate62inter3), .O(gate62inter5));
  nor2  gate805(.a(gate62inter5), .b(gate62inter2), .O(gate62inter6));
  inv1  gate806(.a(G22), .O(gate62inter7));
  inv1  gate807(.a(G296), .O(gate62inter8));
  nand2 gate808(.a(gate62inter8), .b(gate62inter7), .O(gate62inter9));
  nand2 gate809(.a(s_37), .b(gate62inter3), .O(gate62inter10));
  nor2  gate810(.a(gate62inter10), .b(gate62inter9), .O(gate62inter11));
  nor2  gate811(.a(gate62inter11), .b(gate62inter6), .O(gate62inter12));
  nand2 gate812(.a(gate62inter12), .b(gate62inter1), .O(G383));
nand2 gate63( .a(G23), .b(G299), .O(G384) );
nand2 gate64( .a(G24), .b(G299), .O(G385) );
nand2 gate65( .a(G25), .b(G302), .O(G386) );

  xor2  gate1667(.a(G302), .b(G26), .O(gate66inter0));
  nand2 gate1668(.a(gate66inter0), .b(s_160), .O(gate66inter1));
  and2  gate1669(.a(G302), .b(G26), .O(gate66inter2));
  inv1  gate1670(.a(s_160), .O(gate66inter3));
  inv1  gate1671(.a(s_161), .O(gate66inter4));
  nand2 gate1672(.a(gate66inter4), .b(gate66inter3), .O(gate66inter5));
  nor2  gate1673(.a(gate66inter5), .b(gate66inter2), .O(gate66inter6));
  inv1  gate1674(.a(G26), .O(gate66inter7));
  inv1  gate1675(.a(G302), .O(gate66inter8));
  nand2 gate1676(.a(gate66inter8), .b(gate66inter7), .O(gate66inter9));
  nand2 gate1677(.a(s_161), .b(gate66inter3), .O(gate66inter10));
  nor2  gate1678(.a(gate66inter10), .b(gate66inter9), .O(gate66inter11));
  nor2  gate1679(.a(gate66inter11), .b(gate66inter6), .O(gate66inter12));
  nand2 gate1680(.a(gate66inter12), .b(gate66inter1), .O(G387));
nand2 gate67( .a(G27), .b(G305), .O(G388) );
nand2 gate68( .a(G28), .b(G305), .O(G389) );
nand2 gate69( .a(G29), .b(G308), .O(G390) );

  xor2  gate1793(.a(G308), .b(G30), .O(gate70inter0));
  nand2 gate1794(.a(gate70inter0), .b(s_178), .O(gate70inter1));
  and2  gate1795(.a(G308), .b(G30), .O(gate70inter2));
  inv1  gate1796(.a(s_178), .O(gate70inter3));
  inv1  gate1797(.a(s_179), .O(gate70inter4));
  nand2 gate1798(.a(gate70inter4), .b(gate70inter3), .O(gate70inter5));
  nor2  gate1799(.a(gate70inter5), .b(gate70inter2), .O(gate70inter6));
  inv1  gate1800(.a(G30), .O(gate70inter7));
  inv1  gate1801(.a(G308), .O(gate70inter8));
  nand2 gate1802(.a(gate70inter8), .b(gate70inter7), .O(gate70inter9));
  nand2 gate1803(.a(s_179), .b(gate70inter3), .O(gate70inter10));
  nor2  gate1804(.a(gate70inter10), .b(gate70inter9), .O(gate70inter11));
  nor2  gate1805(.a(gate70inter11), .b(gate70inter6), .O(gate70inter12));
  nand2 gate1806(.a(gate70inter12), .b(gate70inter1), .O(G391));
nand2 gate71( .a(G31), .b(G311), .O(G392) );
nand2 gate72( .a(G32), .b(G311), .O(G393) );
nand2 gate73( .a(G1), .b(G314), .O(G394) );
nand2 gate74( .a(G5), .b(G314), .O(G395) );
nand2 gate75( .a(G9), .b(G317), .O(G396) );
nand2 gate76( .a(G13), .b(G317), .O(G397) );

  xor2  gate1611(.a(G320), .b(G2), .O(gate77inter0));
  nand2 gate1612(.a(gate77inter0), .b(s_152), .O(gate77inter1));
  and2  gate1613(.a(G320), .b(G2), .O(gate77inter2));
  inv1  gate1614(.a(s_152), .O(gate77inter3));
  inv1  gate1615(.a(s_153), .O(gate77inter4));
  nand2 gate1616(.a(gate77inter4), .b(gate77inter3), .O(gate77inter5));
  nor2  gate1617(.a(gate77inter5), .b(gate77inter2), .O(gate77inter6));
  inv1  gate1618(.a(G2), .O(gate77inter7));
  inv1  gate1619(.a(G320), .O(gate77inter8));
  nand2 gate1620(.a(gate77inter8), .b(gate77inter7), .O(gate77inter9));
  nand2 gate1621(.a(s_153), .b(gate77inter3), .O(gate77inter10));
  nor2  gate1622(.a(gate77inter10), .b(gate77inter9), .O(gate77inter11));
  nor2  gate1623(.a(gate77inter11), .b(gate77inter6), .O(gate77inter12));
  nand2 gate1624(.a(gate77inter12), .b(gate77inter1), .O(G398));
nand2 gate78( .a(G6), .b(G320), .O(G399) );
nand2 gate79( .a(G10), .b(G323), .O(G400) );

  xor2  gate1639(.a(G323), .b(G14), .O(gate80inter0));
  nand2 gate1640(.a(gate80inter0), .b(s_156), .O(gate80inter1));
  and2  gate1641(.a(G323), .b(G14), .O(gate80inter2));
  inv1  gate1642(.a(s_156), .O(gate80inter3));
  inv1  gate1643(.a(s_157), .O(gate80inter4));
  nand2 gate1644(.a(gate80inter4), .b(gate80inter3), .O(gate80inter5));
  nor2  gate1645(.a(gate80inter5), .b(gate80inter2), .O(gate80inter6));
  inv1  gate1646(.a(G14), .O(gate80inter7));
  inv1  gate1647(.a(G323), .O(gate80inter8));
  nand2 gate1648(.a(gate80inter8), .b(gate80inter7), .O(gate80inter9));
  nand2 gate1649(.a(s_157), .b(gate80inter3), .O(gate80inter10));
  nor2  gate1650(.a(gate80inter10), .b(gate80inter9), .O(gate80inter11));
  nor2  gate1651(.a(gate80inter11), .b(gate80inter6), .O(gate80inter12));
  nand2 gate1652(.a(gate80inter12), .b(gate80inter1), .O(G401));
nand2 gate81( .a(G3), .b(G326), .O(G402) );
nand2 gate82( .a(G7), .b(G326), .O(G403) );
nand2 gate83( .a(G11), .b(G329), .O(G404) );
nand2 gate84( .a(G15), .b(G329), .O(G405) );
nand2 gate85( .a(G4), .b(G332), .O(G406) );

  xor2  gate1331(.a(G332), .b(G8), .O(gate86inter0));
  nand2 gate1332(.a(gate86inter0), .b(s_112), .O(gate86inter1));
  and2  gate1333(.a(G332), .b(G8), .O(gate86inter2));
  inv1  gate1334(.a(s_112), .O(gate86inter3));
  inv1  gate1335(.a(s_113), .O(gate86inter4));
  nand2 gate1336(.a(gate86inter4), .b(gate86inter3), .O(gate86inter5));
  nor2  gate1337(.a(gate86inter5), .b(gate86inter2), .O(gate86inter6));
  inv1  gate1338(.a(G8), .O(gate86inter7));
  inv1  gate1339(.a(G332), .O(gate86inter8));
  nand2 gate1340(.a(gate86inter8), .b(gate86inter7), .O(gate86inter9));
  nand2 gate1341(.a(s_113), .b(gate86inter3), .O(gate86inter10));
  nor2  gate1342(.a(gate86inter10), .b(gate86inter9), .O(gate86inter11));
  nor2  gate1343(.a(gate86inter11), .b(gate86inter6), .O(gate86inter12));
  nand2 gate1344(.a(gate86inter12), .b(gate86inter1), .O(G407));
nand2 gate87( .a(G12), .b(G335), .O(G408) );
nand2 gate88( .a(G16), .b(G335), .O(G409) );

  xor2  gate995(.a(G338), .b(G17), .O(gate89inter0));
  nand2 gate996(.a(gate89inter0), .b(s_64), .O(gate89inter1));
  and2  gate997(.a(G338), .b(G17), .O(gate89inter2));
  inv1  gate998(.a(s_64), .O(gate89inter3));
  inv1  gate999(.a(s_65), .O(gate89inter4));
  nand2 gate1000(.a(gate89inter4), .b(gate89inter3), .O(gate89inter5));
  nor2  gate1001(.a(gate89inter5), .b(gate89inter2), .O(gate89inter6));
  inv1  gate1002(.a(G17), .O(gate89inter7));
  inv1  gate1003(.a(G338), .O(gate89inter8));
  nand2 gate1004(.a(gate89inter8), .b(gate89inter7), .O(gate89inter9));
  nand2 gate1005(.a(s_65), .b(gate89inter3), .O(gate89inter10));
  nor2  gate1006(.a(gate89inter10), .b(gate89inter9), .O(gate89inter11));
  nor2  gate1007(.a(gate89inter11), .b(gate89inter6), .O(gate89inter12));
  nand2 gate1008(.a(gate89inter12), .b(gate89inter1), .O(G410));
nand2 gate90( .a(G21), .b(G338), .O(G411) );
nand2 gate91( .a(G25), .b(G341), .O(G412) );
nand2 gate92( .a(G29), .b(G341), .O(G413) );
nand2 gate93( .a(G18), .b(G344), .O(G414) );
nand2 gate94( .a(G22), .b(G344), .O(G415) );
nand2 gate95( .a(G26), .b(G347), .O(G416) );
nand2 gate96( .a(G30), .b(G347), .O(G417) );
nand2 gate97( .a(G19), .b(G350), .O(G418) );
nand2 gate98( .a(G23), .b(G350), .O(G419) );

  xor2  gate743(.a(G353), .b(G27), .O(gate99inter0));
  nand2 gate744(.a(gate99inter0), .b(s_28), .O(gate99inter1));
  and2  gate745(.a(G353), .b(G27), .O(gate99inter2));
  inv1  gate746(.a(s_28), .O(gate99inter3));
  inv1  gate747(.a(s_29), .O(gate99inter4));
  nand2 gate748(.a(gate99inter4), .b(gate99inter3), .O(gate99inter5));
  nor2  gate749(.a(gate99inter5), .b(gate99inter2), .O(gate99inter6));
  inv1  gate750(.a(G27), .O(gate99inter7));
  inv1  gate751(.a(G353), .O(gate99inter8));
  nand2 gate752(.a(gate99inter8), .b(gate99inter7), .O(gate99inter9));
  nand2 gate753(.a(s_29), .b(gate99inter3), .O(gate99inter10));
  nor2  gate754(.a(gate99inter10), .b(gate99inter9), .O(gate99inter11));
  nor2  gate755(.a(gate99inter11), .b(gate99inter6), .O(gate99inter12));
  nand2 gate756(.a(gate99inter12), .b(gate99inter1), .O(G420));
nand2 gate100( .a(G31), .b(G353), .O(G421) );

  xor2  gate701(.a(G356), .b(G20), .O(gate101inter0));
  nand2 gate702(.a(gate101inter0), .b(s_22), .O(gate101inter1));
  and2  gate703(.a(G356), .b(G20), .O(gate101inter2));
  inv1  gate704(.a(s_22), .O(gate101inter3));
  inv1  gate705(.a(s_23), .O(gate101inter4));
  nand2 gate706(.a(gate101inter4), .b(gate101inter3), .O(gate101inter5));
  nor2  gate707(.a(gate101inter5), .b(gate101inter2), .O(gate101inter6));
  inv1  gate708(.a(G20), .O(gate101inter7));
  inv1  gate709(.a(G356), .O(gate101inter8));
  nand2 gate710(.a(gate101inter8), .b(gate101inter7), .O(gate101inter9));
  nand2 gate711(.a(s_23), .b(gate101inter3), .O(gate101inter10));
  nor2  gate712(.a(gate101inter10), .b(gate101inter9), .O(gate101inter11));
  nor2  gate713(.a(gate101inter11), .b(gate101inter6), .O(gate101inter12));
  nand2 gate714(.a(gate101inter12), .b(gate101inter1), .O(G422));
nand2 gate102( .a(G24), .b(G356), .O(G423) );
nand2 gate103( .a(G28), .b(G359), .O(G424) );
nand2 gate104( .a(G32), .b(G359), .O(G425) );
nand2 gate105( .a(G362), .b(G363), .O(G426) );
nand2 gate106( .a(G364), .b(G365), .O(G429) );

  xor2  gate575(.a(G367), .b(G366), .O(gate107inter0));
  nand2 gate576(.a(gate107inter0), .b(s_4), .O(gate107inter1));
  and2  gate577(.a(G367), .b(G366), .O(gate107inter2));
  inv1  gate578(.a(s_4), .O(gate107inter3));
  inv1  gate579(.a(s_5), .O(gate107inter4));
  nand2 gate580(.a(gate107inter4), .b(gate107inter3), .O(gate107inter5));
  nor2  gate581(.a(gate107inter5), .b(gate107inter2), .O(gate107inter6));
  inv1  gate582(.a(G366), .O(gate107inter7));
  inv1  gate583(.a(G367), .O(gate107inter8));
  nand2 gate584(.a(gate107inter8), .b(gate107inter7), .O(gate107inter9));
  nand2 gate585(.a(s_5), .b(gate107inter3), .O(gate107inter10));
  nor2  gate586(.a(gate107inter10), .b(gate107inter9), .O(gate107inter11));
  nor2  gate587(.a(gate107inter11), .b(gate107inter6), .O(gate107inter12));
  nand2 gate588(.a(gate107inter12), .b(gate107inter1), .O(G432));
nand2 gate108( .a(G368), .b(G369), .O(G435) );
nand2 gate109( .a(G370), .b(G371), .O(G438) );
nand2 gate110( .a(G372), .b(G373), .O(G441) );

  xor2  gate631(.a(G375), .b(G374), .O(gate111inter0));
  nand2 gate632(.a(gate111inter0), .b(s_12), .O(gate111inter1));
  and2  gate633(.a(G375), .b(G374), .O(gate111inter2));
  inv1  gate634(.a(s_12), .O(gate111inter3));
  inv1  gate635(.a(s_13), .O(gate111inter4));
  nand2 gate636(.a(gate111inter4), .b(gate111inter3), .O(gate111inter5));
  nor2  gate637(.a(gate111inter5), .b(gate111inter2), .O(gate111inter6));
  inv1  gate638(.a(G374), .O(gate111inter7));
  inv1  gate639(.a(G375), .O(gate111inter8));
  nand2 gate640(.a(gate111inter8), .b(gate111inter7), .O(gate111inter9));
  nand2 gate641(.a(s_13), .b(gate111inter3), .O(gate111inter10));
  nor2  gate642(.a(gate111inter10), .b(gate111inter9), .O(gate111inter11));
  nor2  gate643(.a(gate111inter11), .b(gate111inter6), .O(gate111inter12));
  nand2 gate644(.a(gate111inter12), .b(gate111inter1), .O(G444));
nand2 gate112( .a(G376), .b(G377), .O(G447) );
nand2 gate113( .a(G378), .b(G379), .O(G450) );
nand2 gate114( .a(G380), .b(G381), .O(G453) );
nand2 gate115( .a(G382), .b(G383), .O(G456) );
nand2 gate116( .a(G384), .b(G385), .O(G459) );
nand2 gate117( .a(G386), .b(G387), .O(G462) );
nand2 gate118( .a(G388), .b(G389), .O(G465) );
nand2 gate119( .a(G390), .b(G391), .O(G468) );
nand2 gate120( .a(G392), .b(G393), .O(G471) );

  xor2  gate2045(.a(G395), .b(G394), .O(gate121inter0));
  nand2 gate2046(.a(gate121inter0), .b(s_214), .O(gate121inter1));
  and2  gate2047(.a(G395), .b(G394), .O(gate121inter2));
  inv1  gate2048(.a(s_214), .O(gate121inter3));
  inv1  gate2049(.a(s_215), .O(gate121inter4));
  nand2 gate2050(.a(gate121inter4), .b(gate121inter3), .O(gate121inter5));
  nor2  gate2051(.a(gate121inter5), .b(gate121inter2), .O(gate121inter6));
  inv1  gate2052(.a(G394), .O(gate121inter7));
  inv1  gate2053(.a(G395), .O(gate121inter8));
  nand2 gate2054(.a(gate121inter8), .b(gate121inter7), .O(gate121inter9));
  nand2 gate2055(.a(s_215), .b(gate121inter3), .O(gate121inter10));
  nor2  gate2056(.a(gate121inter10), .b(gate121inter9), .O(gate121inter11));
  nor2  gate2057(.a(gate121inter11), .b(gate121inter6), .O(gate121inter12));
  nand2 gate2058(.a(gate121inter12), .b(gate121inter1), .O(G474));

  xor2  gate1891(.a(G397), .b(G396), .O(gate122inter0));
  nand2 gate1892(.a(gate122inter0), .b(s_192), .O(gate122inter1));
  and2  gate1893(.a(G397), .b(G396), .O(gate122inter2));
  inv1  gate1894(.a(s_192), .O(gate122inter3));
  inv1  gate1895(.a(s_193), .O(gate122inter4));
  nand2 gate1896(.a(gate122inter4), .b(gate122inter3), .O(gate122inter5));
  nor2  gate1897(.a(gate122inter5), .b(gate122inter2), .O(gate122inter6));
  inv1  gate1898(.a(G396), .O(gate122inter7));
  inv1  gate1899(.a(G397), .O(gate122inter8));
  nand2 gate1900(.a(gate122inter8), .b(gate122inter7), .O(gate122inter9));
  nand2 gate1901(.a(s_193), .b(gate122inter3), .O(gate122inter10));
  nor2  gate1902(.a(gate122inter10), .b(gate122inter9), .O(gate122inter11));
  nor2  gate1903(.a(gate122inter11), .b(gate122inter6), .O(gate122inter12));
  nand2 gate1904(.a(gate122inter12), .b(gate122inter1), .O(G477));
nand2 gate123( .a(G398), .b(G399), .O(G480) );

  xor2  gate687(.a(G401), .b(G400), .O(gate124inter0));
  nand2 gate688(.a(gate124inter0), .b(s_20), .O(gate124inter1));
  and2  gate689(.a(G401), .b(G400), .O(gate124inter2));
  inv1  gate690(.a(s_20), .O(gate124inter3));
  inv1  gate691(.a(s_21), .O(gate124inter4));
  nand2 gate692(.a(gate124inter4), .b(gate124inter3), .O(gate124inter5));
  nor2  gate693(.a(gate124inter5), .b(gate124inter2), .O(gate124inter6));
  inv1  gate694(.a(G400), .O(gate124inter7));
  inv1  gate695(.a(G401), .O(gate124inter8));
  nand2 gate696(.a(gate124inter8), .b(gate124inter7), .O(gate124inter9));
  nand2 gate697(.a(s_21), .b(gate124inter3), .O(gate124inter10));
  nor2  gate698(.a(gate124inter10), .b(gate124inter9), .O(gate124inter11));
  nor2  gate699(.a(gate124inter11), .b(gate124inter6), .O(gate124inter12));
  nand2 gate700(.a(gate124inter12), .b(gate124inter1), .O(G483));
nand2 gate125( .a(G402), .b(G403), .O(G486) );
nand2 gate126( .a(G404), .b(G405), .O(G489) );
nand2 gate127( .a(G406), .b(G407), .O(G492) );
nand2 gate128( .a(G408), .b(G409), .O(G495) );
nand2 gate129( .a(G410), .b(G411), .O(G498) );

  xor2  gate883(.a(G413), .b(G412), .O(gate130inter0));
  nand2 gate884(.a(gate130inter0), .b(s_48), .O(gate130inter1));
  and2  gate885(.a(G413), .b(G412), .O(gate130inter2));
  inv1  gate886(.a(s_48), .O(gate130inter3));
  inv1  gate887(.a(s_49), .O(gate130inter4));
  nand2 gate888(.a(gate130inter4), .b(gate130inter3), .O(gate130inter5));
  nor2  gate889(.a(gate130inter5), .b(gate130inter2), .O(gate130inter6));
  inv1  gate890(.a(G412), .O(gate130inter7));
  inv1  gate891(.a(G413), .O(gate130inter8));
  nand2 gate892(.a(gate130inter8), .b(gate130inter7), .O(gate130inter9));
  nand2 gate893(.a(s_49), .b(gate130inter3), .O(gate130inter10));
  nor2  gate894(.a(gate130inter10), .b(gate130inter9), .O(gate130inter11));
  nor2  gate895(.a(gate130inter11), .b(gate130inter6), .O(gate130inter12));
  nand2 gate896(.a(gate130inter12), .b(gate130inter1), .O(G501));
nand2 gate131( .a(G414), .b(G415), .O(G504) );
nand2 gate132( .a(G416), .b(G417), .O(G507) );
nand2 gate133( .a(G418), .b(G419), .O(G510) );
nand2 gate134( .a(G420), .b(G421), .O(G513) );
nand2 gate135( .a(G422), .b(G423), .O(G516) );
nand2 gate136( .a(G424), .b(G425), .O(G519) );
nand2 gate137( .a(G426), .b(G429), .O(G522) );
nand2 gate138( .a(G432), .b(G435), .O(G525) );
nand2 gate139( .a(G438), .b(G441), .O(G528) );

  xor2  gate1821(.a(G447), .b(G444), .O(gate140inter0));
  nand2 gate1822(.a(gate140inter0), .b(s_182), .O(gate140inter1));
  and2  gate1823(.a(G447), .b(G444), .O(gate140inter2));
  inv1  gate1824(.a(s_182), .O(gate140inter3));
  inv1  gate1825(.a(s_183), .O(gate140inter4));
  nand2 gate1826(.a(gate140inter4), .b(gate140inter3), .O(gate140inter5));
  nor2  gate1827(.a(gate140inter5), .b(gate140inter2), .O(gate140inter6));
  inv1  gate1828(.a(G444), .O(gate140inter7));
  inv1  gate1829(.a(G447), .O(gate140inter8));
  nand2 gate1830(.a(gate140inter8), .b(gate140inter7), .O(gate140inter9));
  nand2 gate1831(.a(s_183), .b(gate140inter3), .O(gate140inter10));
  nor2  gate1832(.a(gate140inter10), .b(gate140inter9), .O(gate140inter11));
  nor2  gate1833(.a(gate140inter11), .b(gate140inter6), .O(gate140inter12));
  nand2 gate1834(.a(gate140inter12), .b(gate140inter1), .O(G531));
nand2 gate141( .a(G450), .b(G453), .O(G534) );
nand2 gate142( .a(G456), .b(G459), .O(G537) );
nand2 gate143( .a(G462), .b(G465), .O(G540) );
nand2 gate144( .a(G468), .b(G471), .O(G543) );
nand2 gate145( .a(G474), .b(G477), .O(G546) );

  xor2  gate1849(.a(G483), .b(G480), .O(gate146inter0));
  nand2 gate1850(.a(gate146inter0), .b(s_186), .O(gate146inter1));
  and2  gate1851(.a(G483), .b(G480), .O(gate146inter2));
  inv1  gate1852(.a(s_186), .O(gate146inter3));
  inv1  gate1853(.a(s_187), .O(gate146inter4));
  nand2 gate1854(.a(gate146inter4), .b(gate146inter3), .O(gate146inter5));
  nor2  gate1855(.a(gate146inter5), .b(gate146inter2), .O(gate146inter6));
  inv1  gate1856(.a(G480), .O(gate146inter7));
  inv1  gate1857(.a(G483), .O(gate146inter8));
  nand2 gate1858(.a(gate146inter8), .b(gate146inter7), .O(gate146inter9));
  nand2 gate1859(.a(s_187), .b(gate146inter3), .O(gate146inter10));
  nor2  gate1860(.a(gate146inter10), .b(gate146inter9), .O(gate146inter11));
  nor2  gate1861(.a(gate146inter11), .b(gate146inter6), .O(gate146inter12));
  nand2 gate1862(.a(gate146inter12), .b(gate146inter1), .O(G549));
nand2 gate147( .a(G486), .b(G489), .O(G552) );

  xor2  gate1919(.a(G495), .b(G492), .O(gate148inter0));
  nand2 gate1920(.a(gate148inter0), .b(s_196), .O(gate148inter1));
  and2  gate1921(.a(G495), .b(G492), .O(gate148inter2));
  inv1  gate1922(.a(s_196), .O(gate148inter3));
  inv1  gate1923(.a(s_197), .O(gate148inter4));
  nand2 gate1924(.a(gate148inter4), .b(gate148inter3), .O(gate148inter5));
  nor2  gate1925(.a(gate148inter5), .b(gate148inter2), .O(gate148inter6));
  inv1  gate1926(.a(G492), .O(gate148inter7));
  inv1  gate1927(.a(G495), .O(gate148inter8));
  nand2 gate1928(.a(gate148inter8), .b(gate148inter7), .O(gate148inter9));
  nand2 gate1929(.a(s_197), .b(gate148inter3), .O(gate148inter10));
  nor2  gate1930(.a(gate148inter10), .b(gate148inter9), .O(gate148inter11));
  nor2  gate1931(.a(gate148inter11), .b(gate148inter6), .O(gate148inter12));
  nand2 gate1932(.a(gate148inter12), .b(gate148inter1), .O(G555));
nand2 gate149( .a(G498), .b(G501), .O(G558) );
nand2 gate150( .a(G504), .b(G507), .O(G561) );
nand2 gate151( .a(G510), .b(G513), .O(G564) );

  xor2  gate911(.a(G519), .b(G516), .O(gate152inter0));
  nand2 gate912(.a(gate152inter0), .b(s_52), .O(gate152inter1));
  and2  gate913(.a(G519), .b(G516), .O(gate152inter2));
  inv1  gate914(.a(s_52), .O(gate152inter3));
  inv1  gate915(.a(s_53), .O(gate152inter4));
  nand2 gate916(.a(gate152inter4), .b(gate152inter3), .O(gate152inter5));
  nor2  gate917(.a(gate152inter5), .b(gate152inter2), .O(gate152inter6));
  inv1  gate918(.a(G516), .O(gate152inter7));
  inv1  gate919(.a(G519), .O(gate152inter8));
  nand2 gate920(.a(gate152inter8), .b(gate152inter7), .O(gate152inter9));
  nand2 gate921(.a(s_53), .b(gate152inter3), .O(gate152inter10));
  nor2  gate922(.a(gate152inter10), .b(gate152inter9), .O(gate152inter11));
  nor2  gate923(.a(gate152inter11), .b(gate152inter6), .O(gate152inter12));
  nand2 gate924(.a(gate152inter12), .b(gate152inter1), .O(G567));
nand2 gate153( .a(G426), .b(G522), .O(G570) );
nand2 gate154( .a(G429), .b(G522), .O(G571) );
nand2 gate155( .a(G432), .b(G525), .O(G572) );
nand2 gate156( .a(G435), .b(G525), .O(G573) );

  xor2  gate589(.a(G528), .b(G438), .O(gate157inter0));
  nand2 gate590(.a(gate157inter0), .b(s_6), .O(gate157inter1));
  and2  gate591(.a(G528), .b(G438), .O(gate157inter2));
  inv1  gate592(.a(s_6), .O(gate157inter3));
  inv1  gate593(.a(s_7), .O(gate157inter4));
  nand2 gate594(.a(gate157inter4), .b(gate157inter3), .O(gate157inter5));
  nor2  gate595(.a(gate157inter5), .b(gate157inter2), .O(gate157inter6));
  inv1  gate596(.a(G438), .O(gate157inter7));
  inv1  gate597(.a(G528), .O(gate157inter8));
  nand2 gate598(.a(gate157inter8), .b(gate157inter7), .O(gate157inter9));
  nand2 gate599(.a(s_7), .b(gate157inter3), .O(gate157inter10));
  nor2  gate600(.a(gate157inter10), .b(gate157inter9), .O(gate157inter11));
  nor2  gate601(.a(gate157inter11), .b(gate157inter6), .O(gate157inter12));
  nand2 gate602(.a(gate157inter12), .b(gate157inter1), .O(G574));

  xor2  gate967(.a(G528), .b(G441), .O(gate158inter0));
  nand2 gate968(.a(gate158inter0), .b(s_60), .O(gate158inter1));
  and2  gate969(.a(G528), .b(G441), .O(gate158inter2));
  inv1  gate970(.a(s_60), .O(gate158inter3));
  inv1  gate971(.a(s_61), .O(gate158inter4));
  nand2 gate972(.a(gate158inter4), .b(gate158inter3), .O(gate158inter5));
  nor2  gate973(.a(gate158inter5), .b(gate158inter2), .O(gate158inter6));
  inv1  gate974(.a(G441), .O(gate158inter7));
  inv1  gate975(.a(G528), .O(gate158inter8));
  nand2 gate976(.a(gate158inter8), .b(gate158inter7), .O(gate158inter9));
  nand2 gate977(.a(s_61), .b(gate158inter3), .O(gate158inter10));
  nor2  gate978(.a(gate158inter10), .b(gate158inter9), .O(gate158inter11));
  nor2  gate979(.a(gate158inter11), .b(gate158inter6), .O(gate158inter12));
  nand2 gate980(.a(gate158inter12), .b(gate158inter1), .O(G575));
nand2 gate159( .a(G444), .b(G531), .O(G576) );
nand2 gate160( .a(G447), .b(G531), .O(G577) );
nand2 gate161( .a(G450), .b(G534), .O(G578) );
nand2 gate162( .a(G453), .b(G534), .O(G579) );
nand2 gate163( .a(G456), .b(G537), .O(G580) );
nand2 gate164( .a(G459), .b(G537), .O(G581) );
nand2 gate165( .a(G462), .b(G540), .O(G582) );
nand2 gate166( .a(G465), .b(G540), .O(G583) );
nand2 gate167( .a(G468), .b(G543), .O(G584) );
nand2 gate168( .a(G471), .b(G543), .O(G585) );

  xor2  gate1905(.a(G546), .b(G474), .O(gate169inter0));
  nand2 gate1906(.a(gate169inter0), .b(s_194), .O(gate169inter1));
  and2  gate1907(.a(G546), .b(G474), .O(gate169inter2));
  inv1  gate1908(.a(s_194), .O(gate169inter3));
  inv1  gate1909(.a(s_195), .O(gate169inter4));
  nand2 gate1910(.a(gate169inter4), .b(gate169inter3), .O(gate169inter5));
  nor2  gate1911(.a(gate169inter5), .b(gate169inter2), .O(gate169inter6));
  inv1  gate1912(.a(G474), .O(gate169inter7));
  inv1  gate1913(.a(G546), .O(gate169inter8));
  nand2 gate1914(.a(gate169inter8), .b(gate169inter7), .O(gate169inter9));
  nand2 gate1915(.a(s_195), .b(gate169inter3), .O(gate169inter10));
  nor2  gate1916(.a(gate169inter10), .b(gate169inter9), .O(gate169inter11));
  nor2  gate1917(.a(gate169inter11), .b(gate169inter6), .O(gate169inter12));
  nand2 gate1918(.a(gate169inter12), .b(gate169inter1), .O(G586));
nand2 gate170( .a(G477), .b(G546), .O(G587) );
nand2 gate171( .a(G480), .b(G549), .O(G588) );
nand2 gate172( .a(G483), .b(G549), .O(G589) );
nand2 gate173( .a(G486), .b(G552), .O(G590) );

  xor2  gate1233(.a(G552), .b(G489), .O(gate174inter0));
  nand2 gate1234(.a(gate174inter0), .b(s_98), .O(gate174inter1));
  and2  gate1235(.a(G552), .b(G489), .O(gate174inter2));
  inv1  gate1236(.a(s_98), .O(gate174inter3));
  inv1  gate1237(.a(s_99), .O(gate174inter4));
  nand2 gate1238(.a(gate174inter4), .b(gate174inter3), .O(gate174inter5));
  nor2  gate1239(.a(gate174inter5), .b(gate174inter2), .O(gate174inter6));
  inv1  gate1240(.a(G489), .O(gate174inter7));
  inv1  gate1241(.a(G552), .O(gate174inter8));
  nand2 gate1242(.a(gate174inter8), .b(gate174inter7), .O(gate174inter9));
  nand2 gate1243(.a(s_99), .b(gate174inter3), .O(gate174inter10));
  nor2  gate1244(.a(gate174inter10), .b(gate174inter9), .O(gate174inter11));
  nor2  gate1245(.a(gate174inter11), .b(gate174inter6), .O(gate174inter12));
  nand2 gate1246(.a(gate174inter12), .b(gate174inter1), .O(G591));

  xor2  gate2143(.a(G555), .b(G492), .O(gate175inter0));
  nand2 gate2144(.a(gate175inter0), .b(s_228), .O(gate175inter1));
  and2  gate2145(.a(G555), .b(G492), .O(gate175inter2));
  inv1  gate2146(.a(s_228), .O(gate175inter3));
  inv1  gate2147(.a(s_229), .O(gate175inter4));
  nand2 gate2148(.a(gate175inter4), .b(gate175inter3), .O(gate175inter5));
  nor2  gate2149(.a(gate175inter5), .b(gate175inter2), .O(gate175inter6));
  inv1  gate2150(.a(G492), .O(gate175inter7));
  inv1  gate2151(.a(G555), .O(gate175inter8));
  nand2 gate2152(.a(gate175inter8), .b(gate175inter7), .O(gate175inter9));
  nand2 gate2153(.a(s_229), .b(gate175inter3), .O(gate175inter10));
  nor2  gate2154(.a(gate175inter10), .b(gate175inter9), .O(gate175inter11));
  nor2  gate2155(.a(gate175inter11), .b(gate175inter6), .O(gate175inter12));
  nand2 gate2156(.a(gate175inter12), .b(gate175inter1), .O(G592));
nand2 gate176( .a(G495), .b(G555), .O(G593) );
nand2 gate177( .a(G498), .b(G558), .O(G594) );

  xor2  gate1443(.a(G558), .b(G501), .O(gate178inter0));
  nand2 gate1444(.a(gate178inter0), .b(s_128), .O(gate178inter1));
  and2  gate1445(.a(G558), .b(G501), .O(gate178inter2));
  inv1  gate1446(.a(s_128), .O(gate178inter3));
  inv1  gate1447(.a(s_129), .O(gate178inter4));
  nand2 gate1448(.a(gate178inter4), .b(gate178inter3), .O(gate178inter5));
  nor2  gate1449(.a(gate178inter5), .b(gate178inter2), .O(gate178inter6));
  inv1  gate1450(.a(G501), .O(gate178inter7));
  inv1  gate1451(.a(G558), .O(gate178inter8));
  nand2 gate1452(.a(gate178inter8), .b(gate178inter7), .O(gate178inter9));
  nand2 gate1453(.a(s_129), .b(gate178inter3), .O(gate178inter10));
  nor2  gate1454(.a(gate178inter10), .b(gate178inter9), .O(gate178inter11));
  nor2  gate1455(.a(gate178inter11), .b(gate178inter6), .O(gate178inter12));
  nand2 gate1456(.a(gate178inter12), .b(gate178inter1), .O(G595));
nand2 gate179( .a(G504), .b(G561), .O(G596) );
nand2 gate180( .a(G507), .b(G561), .O(G597) );
nand2 gate181( .a(G510), .b(G564), .O(G598) );

  xor2  gate1415(.a(G564), .b(G513), .O(gate182inter0));
  nand2 gate1416(.a(gate182inter0), .b(s_124), .O(gate182inter1));
  and2  gate1417(.a(G564), .b(G513), .O(gate182inter2));
  inv1  gate1418(.a(s_124), .O(gate182inter3));
  inv1  gate1419(.a(s_125), .O(gate182inter4));
  nand2 gate1420(.a(gate182inter4), .b(gate182inter3), .O(gate182inter5));
  nor2  gate1421(.a(gate182inter5), .b(gate182inter2), .O(gate182inter6));
  inv1  gate1422(.a(G513), .O(gate182inter7));
  inv1  gate1423(.a(G564), .O(gate182inter8));
  nand2 gate1424(.a(gate182inter8), .b(gate182inter7), .O(gate182inter9));
  nand2 gate1425(.a(s_125), .b(gate182inter3), .O(gate182inter10));
  nor2  gate1426(.a(gate182inter10), .b(gate182inter9), .O(gate182inter11));
  nor2  gate1427(.a(gate182inter11), .b(gate182inter6), .O(gate182inter12));
  nand2 gate1428(.a(gate182inter12), .b(gate182inter1), .O(G599));
nand2 gate183( .a(G516), .b(G567), .O(G600) );
nand2 gate184( .a(G519), .b(G567), .O(G601) );
nand2 gate185( .a(G570), .b(G571), .O(G602) );

  xor2  gate2059(.a(G573), .b(G572), .O(gate186inter0));
  nand2 gate2060(.a(gate186inter0), .b(s_216), .O(gate186inter1));
  and2  gate2061(.a(G573), .b(G572), .O(gate186inter2));
  inv1  gate2062(.a(s_216), .O(gate186inter3));
  inv1  gate2063(.a(s_217), .O(gate186inter4));
  nand2 gate2064(.a(gate186inter4), .b(gate186inter3), .O(gate186inter5));
  nor2  gate2065(.a(gate186inter5), .b(gate186inter2), .O(gate186inter6));
  inv1  gate2066(.a(G572), .O(gate186inter7));
  inv1  gate2067(.a(G573), .O(gate186inter8));
  nand2 gate2068(.a(gate186inter8), .b(gate186inter7), .O(gate186inter9));
  nand2 gate2069(.a(s_217), .b(gate186inter3), .O(gate186inter10));
  nor2  gate2070(.a(gate186inter10), .b(gate186inter9), .O(gate186inter11));
  nor2  gate2071(.a(gate186inter11), .b(gate186inter6), .O(gate186inter12));
  nand2 gate2072(.a(gate186inter12), .b(gate186inter1), .O(G607));

  xor2  gate1275(.a(G575), .b(G574), .O(gate187inter0));
  nand2 gate1276(.a(gate187inter0), .b(s_104), .O(gate187inter1));
  and2  gate1277(.a(G575), .b(G574), .O(gate187inter2));
  inv1  gate1278(.a(s_104), .O(gate187inter3));
  inv1  gate1279(.a(s_105), .O(gate187inter4));
  nand2 gate1280(.a(gate187inter4), .b(gate187inter3), .O(gate187inter5));
  nor2  gate1281(.a(gate187inter5), .b(gate187inter2), .O(gate187inter6));
  inv1  gate1282(.a(G574), .O(gate187inter7));
  inv1  gate1283(.a(G575), .O(gate187inter8));
  nand2 gate1284(.a(gate187inter8), .b(gate187inter7), .O(gate187inter9));
  nand2 gate1285(.a(s_105), .b(gate187inter3), .O(gate187inter10));
  nor2  gate1286(.a(gate187inter10), .b(gate187inter9), .O(gate187inter11));
  nor2  gate1287(.a(gate187inter11), .b(gate187inter6), .O(gate187inter12));
  nand2 gate1288(.a(gate187inter12), .b(gate187inter1), .O(G612));
nand2 gate188( .a(G576), .b(G577), .O(G617) );
nand2 gate189( .a(G578), .b(G579), .O(G622) );
nand2 gate190( .a(G580), .b(G581), .O(G627) );

  xor2  gate1765(.a(G583), .b(G582), .O(gate191inter0));
  nand2 gate1766(.a(gate191inter0), .b(s_174), .O(gate191inter1));
  and2  gate1767(.a(G583), .b(G582), .O(gate191inter2));
  inv1  gate1768(.a(s_174), .O(gate191inter3));
  inv1  gate1769(.a(s_175), .O(gate191inter4));
  nand2 gate1770(.a(gate191inter4), .b(gate191inter3), .O(gate191inter5));
  nor2  gate1771(.a(gate191inter5), .b(gate191inter2), .O(gate191inter6));
  inv1  gate1772(.a(G582), .O(gate191inter7));
  inv1  gate1773(.a(G583), .O(gate191inter8));
  nand2 gate1774(.a(gate191inter8), .b(gate191inter7), .O(gate191inter9));
  nand2 gate1775(.a(s_175), .b(gate191inter3), .O(gate191inter10));
  nor2  gate1776(.a(gate191inter10), .b(gate191inter9), .O(gate191inter11));
  nor2  gate1777(.a(gate191inter11), .b(gate191inter6), .O(gate191inter12));
  nand2 gate1778(.a(gate191inter12), .b(gate191inter1), .O(G632));
nand2 gate192( .a(G584), .b(G585), .O(G637) );
nand2 gate193( .a(G586), .b(G587), .O(G642) );

  xor2  gate715(.a(G589), .b(G588), .O(gate194inter0));
  nand2 gate716(.a(gate194inter0), .b(s_24), .O(gate194inter1));
  and2  gate717(.a(G589), .b(G588), .O(gate194inter2));
  inv1  gate718(.a(s_24), .O(gate194inter3));
  inv1  gate719(.a(s_25), .O(gate194inter4));
  nand2 gate720(.a(gate194inter4), .b(gate194inter3), .O(gate194inter5));
  nor2  gate721(.a(gate194inter5), .b(gate194inter2), .O(gate194inter6));
  inv1  gate722(.a(G588), .O(gate194inter7));
  inv1  gate723(.a(G589), .O(gate194inter8));
  nand2 gate724(.a(gate194inter8), .b(gate194inter7), .O(gate194inter9));
  nand2 gate725(.a(s_25), .b(gate194inter3), .O(gate194inter10));
  nor2  gate726(.a(gate194inter10), .b(gate194inter9), .O(gate194inter11));
  nor2  gate727(.a(gate194inter11), .b(gate194inter6), .O(gate194inter12));
  nand2 gate728(.a(gate194inter12), .b(gate194inter1), .O(G645));

  xor2  gate1093(.a(G591), .b(G590), .O(gate195inter0));
  nand2 gate1094(.a(gate195inter0), .b(s_78), .O(gate195inter1));
  and2  gate1095(.a(G591), .b(G590), .O(gate195inter2));
  inv1  gate1096(.a(s_78), .O(gate195inter3));
  inv1  gate1097(.a(s_79), .O(gate195inter4));
  nand2 gate1098(.a(gate195inter4), .b(gate195inter3), .O(gate195inter5));
  nor2  gate1099(.a(gate195inter5), .b(gate195inter2), .O(gate195inter6));
  inv1  gate1100(.a(G590), .O(gate195inter7));
  inv1  gate1101(.a(G591), .O(gate195inter8));
  nand2 gate1102(.a(gate195inter8), .b(gate195inter7), .O(gate195inter9));
  nand2 gate1103(.a(s_79), .b(gate195inter3), .O(gate195inter10));
  nor2  gate1104(.a(gate195inter10), .b(gate195inter9), .O(gate195inter11));
  nor2  gate1105(.a(gate195inter11), .b(gate195inter6), .O(gate195inter12));
  nand2 gate1106(.a(gate195inter12), .b(gate195inter1), .O(G648));
nand2 gate196( .a(G592), .b(G593), .O(G651) );
nand2 gate197( .a(G594), .b(G595), .O(G654) );
nand2 gate198( .a(G596), .b(G597), .O(G657) );
nand2 gate199( .a(G598), .b(G599), .O(G660) );
nand2 gate200( .a(G600), .b(G601), .O(G663) );

  xor2  gate1723(.a(G607), .b(G602), .O(gate201inter0));
  nand2 gate1724(.a(gate201inter0), .b(s_168), .O(gate201inter1));
  and2  gate1725(.a(G607), .b(G602), .O(gate201inter2));
  inv1  gate1726(.a(s_168), .O(gate201inter3));
  inv1  gate1727(.a(s_169), .O(gate201inter4));
  nand2 gate1728(.a(gate201inter4), .b(gate201inter3), .O(gate201inter5));
  nor2  gate1729(.a(gate201inter5), .b(gate201inter2), .O(gate201inter6));
  inv1  gate1730(.a(G602), .O(gate201inter7));
  inv1  gate1731(.a(G607), .O(gate201inter8));
  nand2 gate1732(.a(gate201inter8), .b(gate201inter7), .O(gate201inter9));
  nand2 gate1733(.a(s_169), .b(gate201inter3), .O(gate201inter10));
  nor2  gate1734(.a(gate201inter10), .b(gate201inter9), .O(gate201inter11));
  nor2  gate1735(.a(gate201inter11), .b(gate201inter6), .O(gate201inter12));
  nand2 gate1736(.a(gate201inter12), .b(gate201inter1), .O(G666));

  xor2  gate1135(.a(G617), .b(G612), .O(gate202inter0));
  nand2 gate1136(.a(gate202inter0), .b(s_84), .O(gate202inter1));
  and2  gate1137(.a(G617), .b(G612), .O(gate202inter2));
  inv1  gate1138(.a(s_84), .O(gate202inter3));
  inv1  gate1139(.a(s_85), .O(gate202inter4));
  nand2 gate1140(.a(gate202inter4), .b(gate202inter3), .O(gate202inter5));
  nor2  gate1141(.a(gate202inter5), .b(gate202inter2), .O(gate202inter6));
  inv1  gate1142(.a(G612), .O(gate202inter7));
  inv1  gate1143(.a(G617), .O(gate202inter8));
  nand2 gate1144(.a(gate202inter8), .b(gate202inter7), .O(gate202inter9));
  nand2 gate1145(.a(s_85), .b(gate202inter3), .O(gate202inter10));
  nor2  gate1146(.a(gate202inter10), .b(gate202inter9), .O(gate202inter11));
  nor2  gate1147(.a(gate202inter11), .b(gate202inter6), .O(gate202inter12));
  nand2 gate1148(.a(gate202inter12), .b(gate202inter1), .O(G669));
nand2 gate203( .a(G602), .b(G612), .O(G672) );
nand2 gate204( .a(G607), .b(G617), .O(G675) );
nand2 gate205( .a(G622), .b(G627), .O(G678) );
nand2 gate206( .a(G632), .b(G637), .O(G681) );
nand2 gate207( .a(G622), .b(G632), .O(G684) );

  xor2  gate1653(.a(G637), .b(G627), .O(gate208inter0));
  nand2 gate1654(.a(gate208inter0), .b(s_158), .O(gate208inter1));
  and2  gate1655(.a(G637), .b(G627), .O(gate208inter2));
  inv1  gate1656(.a(s_158), .O(gate208inter3));
  inv1  gate1657(.a(s_159), .O(gate208inter4));
  nand2 gate1658(.a(gate208inter4), .b(gate208inter3), .O(gate208inter5));
  nor2  gate1659(.a(gate208inter5), .b(gate208inter2), .O(gate208inter6));
  inv1  gate1660(.a(G627), .O(gate208inter7));
  inv1  gate1661(.a(G637), .O(gate208inter8));
  nand2 gate1662(.a(gate208inter8), .b(gate208inter7), .O(gate208inter9));
  nand2 gate1663(.a(s_159), .b(gate208inter3), .O(gate208inter10));
  nor2  gate1664(.a(gate208inter10), .b(gate208inter9), .O(gate208inter11));
  nor2  gate1665(.a(gate208inter11), .b(gate208inter6), .O(gate208inter12));
  nand2 gate1666(.a(gate208inter12), .b(gate208inter1), .O(G687));
nand2 gate209( .a(G602), .b(G666), .O(G690) );
nand2 gate210( .a(G607), .b(G666), .O(G691) );
nand2 gate211( .a(G612), .b(G669), .O(G692) );
nand2 gate212( .a(G617), .b(G669), .O(G693) );

  xor2  gate785(.a(G672), .b(G602), .O(gate213inter0));
  nand2 gate786(.a(gate213inter0), .b(s_34), .O(gate213inter1));
  and2  gate787(.a(G672), .b(G602), .O(gate213inter2));
  inv1  gate788(.a(s_34), .O(gate213inter3));
  inv1  gate789(.a(s_35), .O(gate213inter4));
  nand2 gate790(.a(gate213inter4), .b(gate213inter3), .O(gate213inter5));
  nor2  gate791(.a(gate213inter5), .b(gate213inter2), .O(gate213inter6));
  inv1  gate792(.a(G602), .O(gate213inter7));
  inv1  gate793(.a(G672), .O(gate213inter8));
  nand2 gate794(.a(gate213inter8), .b(gate213inter7), .O(gate213inter9));
  nand2 gate795(.a(s_35), .b(gate213inter3), .O(gate213inter10));
  nor2  gate796(.a(gate213inter10), .b(gate213inter9), .O(gate213inter11));
  nor2  gate797(.a(gate213inter11), .b(gate213inter6), .O(gate213inter12));
  nand2 gate798(.a(gate213inter12), .b(gate213inter1), .O(G694));
nand2 gate214( .a(G612), .b(G672), .O(G695) );
nand2 gate215( .a(G607), .b(G675), .O(G696) );
nand2 gate216( .a(G617), .b(G675), .O(G697) );
nand2 gate217( .a(G622), .b(G678), .O(G698) );

  xor2  gate2017(.a(G678), .b(G627), .O(gate218inter0));
  nand2 gate2018(.a(gate218inter0), .b(s_210), .O(gate218inter1));
  and2  gate2019(.a(G678), .b(G627), .O(gate218inter2));
  inv1  gate2020(.a(s_210), .O(gate218inter3));
  inv1  gate2021(.a(s_211), .O(gate218inter4));
  nand2 gate2022(.a(gate218inter4), .b(gate218inter3), .O(gate218inter5));
  nor2  gate2023(.a(gate218inter5), .b(gate218inter2), .O(gate218inter6));
  inv1  gate2024(.a(G627), .O(gate218inter7));
  inv1  gate2025(.a(G678), .O(gate218inter8));
  nand2 gate2026(.a(gate218inter8), .b(gate218inter7), .O(gate218inter9));
  nand2 gate2027(.a(s_211), .b(gate218inter3), .O(gate218inter10));
  nor2  gate2028(.a(gate218inter10), .b(gate218inter9), .O(gate218inter11));
  nor2  gate2029(.a(gate218inter11), .b(gate218inter6), .O(gate218inter12));
  nand2 gate2030(.a(gate218inter12), .b(gate218inter1), .O(G699));
nand2 gate219( .a(G632), .b(G681), .O(G700) );

  xor2  gate1681(.a(G681), .b(G637), .O(gate220inter0));
  nand2 gate1682(.a(gate220inter0), .b(s_162), .O(gate220inter1));
  and2  gate1683(.a(G681), .b(G637), .O(gate220inter2));
  inv1  gate1684(.a(s_162), .O(gate220inter3));
  inv1  gate1685(.a(s_163), .O(gate220inter4));
  nand2 gate1686(.a(gate220inter4), .b(gate220inter3), .O(gate220inter5));
  nor2  gate1687(.a(gate220inter5), .b(gate220inter2), .O(gate220inter6));
  inv1  gate1688(.a(G637), .O(gate220inter7));
  inv1  gate1689(.a(G681), .O(gate220inter8));
  nand2 gate1690(.a(gate220inter8), .b(gate220inter7), .O(gate220inter9));
  nand2 gate1691(.a(s_163), .b(gate220inter3), .O(gate220inter10));
  nor2  gate1692(.a(gate220inter10), .b(gate220inter9), .O(gate220inter11));
  nor2  gate1693(.a(gate220inter11), .b(gate220inter6), .O(gate220inter12));
  nand2 gate1694(.a(gate220inter12), .b(gate220inter1), .O(G701));
nand2 gate221( .a(G622), .b(G684), .O(G702) );
nand2 gate222( .a(G632), .b(G684), .O(G703) );
nand2 gate223( .a(G627), .b(G687), .O(G704) );
nand2 gate224( .a(G637), .b(G687), .O(G705) );
nand2 gate225( .a(G690), .b(G691), .O(G706) );
nand2 gate226( .a(G692), .b(G693), .O(G709) );

  xor2  gate1569(.a(G695), .b(G694), .O(gate227inter0));
  nand2 gate1570(.a(gate227inter0), .b(s_146), .O(gate227inter1));
  and2  gate1571(.a(G695), .b(G694), .O(gate227inter2));
  inv1  gate1572(.a(s_146), .O(gate227inter3));
  inv1  gate1573(.a(s_147), .O(gate227inter4));
  nand2 gate1574(.a(gate227inter4), .b(gate227inter3), .O(gate227inter5));
  nor2  gate1575(.a(gate227inter5), .b(gate227inter2), .O(gate227inter6));
  inv1  gate1576(.a(G694), .O(gate227inter7));
  inv1  gate1577(.a(G695), .O(gate227inter8));
  nand2 gate1578(.a(gate227inter8), .b(gate227inter7), .O(gate227inter9));
  nand2 gate1579(.a(s_147), .b(gate227inter3), .O(gate227inter10));
  nor2  gate1580(.a(gate227inter10), .b(gate227inter9), .O(gate227inter11));
  nor2  gate1581(.a(gate227inter11), .b(gate227inter6), .O(gate227inter12));
  nand2 gate1582(.a(gate227inter12), .b(gate227inter1), .O(G712));

  xor2  gate603(.a(G697), .b(G696), .O(gate228inter0));
  nand2 gate604(.a(gate228inter0), .b(s_8), .O(gate228inter1));
  and2  gate605(.a(G697), .b(G696), .O(gate228inter2));
  inv1  gate606(.a(s_8), .O(gate228inter3));
  inv1  gate607(.a(s_9), .O(gate228inter4));
  nand2 gate608(.a(gate228inter4), .b(gate228inter3), .O(gate228inter5));
  nor2  gate609(.a(gate228inter5), .b(gate228inter2), .O(gate228inter6));
  inv1  gate610(.a(G696), .O(gate228inter7));
  inv1  gate611(.a(G697), .O(gate228inter8));
  nand2 gate612(.a(gate228inter8), .b(gate228inter7), .O(gate228inter9));
  nand2 gate613(.a(s_9), .b(gate228inter3), .O(gate228inter10));
  nor2  gate614(.a(gate228inter10), .b(gate228inter9), .O(gate228inter11));
  nor2  gate615(.a(gate228inter11), .b(gate228inter6), .O(gate228inter12));
  nand2 gate616(.a(gate228inter12), .b(gate228inter1), .O(G715));
nand2 gate229( .a(G698), .b(G699), .O(G718) );
nand2 gate230( .a(G700), .b(G701), .O(G721) );
nand2 gate231( .a(G702), .b(G703), .O(G724) );
nand2 gate232( .a(G704), .b(G705), .O(G727) );
nand2 gate233( .a(G242), .b(G718), .O(G730) );
nand2 gate234( .a(G245), .b(G721), .O(G733) );
nand2 gate235( .a(G248), .b(G724), .O(G736) );
nand2 gate236( .a(G251), .b(G727), .O(G739) );
nand2 gate237( .a(G254), .b(G706), .O(G742) );
nand2 gate238( .a(G257), .b(G709), .O(G745) );

  xor2  gate1779(.a(G712), .b(G260), .O(gate239inter0));
  nand2 gate1780(.a(gate239inter0), .b(s_176), .O(gate239inter1));
  and2  gate1781(.a(G712), .b(G260), .O(gate239inter2));
  inv1  gate1782(.a(s_176), .O(gate239inter3));
  inv1  gate1783(.a(s_177), .O(gate239inter4));
  nand2 gate1784(.a(gate239inter4), .b(gate239inter3), .O(gate239inter5));
  nor2  gate1785(.a(gate239inter5), .b(gate239inter2), .O(gate239inter6));
  inv1  gate1786(.a(G260), .O(gate239inter7));
  inv1  gate1787(.a(G712), .O(gate239inter8));
  nand2 gate1788(.a(gate239inter8), .b(gate239inter7), .O(gate239inter9));
  nand2 gate1789(.a(s_177), .b(gate239inter3), .O(gate239inter10));
  nor2  gate1790(.a(gate239inter10), .b(gate239inter9), .O(gate239inter11));
  nor2  gate1791(.a(gate239inter11), .b(gate239inter6), .O(gate239inter12));
  nand2 gate1792(.a(gate239inter12), .b(gate239inter1), .O(G748));

  xor2  gate1345(.a(G715), .b(G263), .O(gate240inter0));
  nand2 gate1346(.a(gate240inter0), .b(s_114), .O(gate240inter1));
  and2  gate1347(.a(G715), .b(G263), .O(gate240inter2));
  inv1  gate1348(.a(s_114), .O(gate240inter3));
  inv1  gate1349(.a(s_115), .O(gate240inter4));
  nand2 gate1350(.a(gate240inter4), .b(gate240inter3), .O(gate240inter5));
  nor2  gate1351(.a(gate240inter5), .b(gate240inter2), .O(gate240inter6));
  inv1  gate1352(.a(G263), .O(gate240inter7));
  inv1  gate1353(.a(G715), .O(gate240inter8));
  nand2 gate1354(.a(gate240inter8), .b(gate240inter7), .O(gate240inter9));
  nand2 gate1355(.a(s_115), .b(gate240inter3), .O(gate240inter10));
  nor2  gate1356(.a(gate240inter10), .b(gate240inter9), .O(gate240inter11));
  nor2  gate1357(.a(gate240inter11), .b(gate240inter6), .O(gate240inter12));
  nand2 gate1358(.a(gate240inter12), .b(gate240inter1), .O(G751));
nand2 gate241( .a(G242), .b(G730), .O(G754) );

  xor2  gate547(.a(G730), .b(G718), .O(gate242inter0));
  nand2 gate548(.a(gate242inter0), .b(s_0), .O(gate242inter1));
  and2  gate549(.a(G730), .b(G718), .O(gate242inter2));
  inv1  gate550(.a(s_0), .O(gate242inter3));
  inv1  gate551(.a(s_1), .O(gate242inter4));
  nand2 gate552(.a(gate242inter4), .b(gate242inter3), .O(gate242inter5));
  nor2  gate553(.a(gate242inter5), .b(gate242inter2), .O(gate242inter6));
  inv1  gate554(.a(G718), .O(gate242inter7));
  inv1  gate555(.a(G730), .O(gate242inter8));
  nand2 gate556(.a(gate242inter8), .b(gate242inter7), .O(gate242inter9));
  nand2 gate557(.a(s_1), .b(gate242inter3), .O(gate242inter10));
  nor2  gate558(.a(gate242inter10), .b(gate242inter9), .O(gate242inter11));
  nor2  gate559(.a(gate242inter11), .b(gate242inter6), .O(gate242inter12));
  nand2 gate560(.a(gate242inter12), .b(gate242inter1), .O(G755));
nand2 gate243( .a(G245), .b(G733), .O(G756) );
nand2 gate244( .a(G721), .b(G733), .O(G757) );
nand2 gate245( .a(G248), .b(G736), .O(G758) );
nand2 gate246( .a(G724), .b(G736), .O(G759) );

  xor2  gate1401(.a(G739), .b(G251), .O(gate247inter0));
  nand2 gate1402(.a(gate247inter0), .b(s_122), .O(gate247inter1));
  and2  gate1403(.a(G739), .b(G251), .O(gate247inter2));
  inv1  gate1404(.a(s_122), .O(gate247inter3));
  inv1  gate1405(.a(s_123), .O(gate247inter4));
  nand2 gate1406(.a(gate247inter4), .b(gate247inter3), .O(gate247inter5));
  nor2  gate1407(.a(gate247inter5), .b(gate247inter2), .O(gate247inter6));
  inv1  gate1408(.a(G251), .O(gate247inter7));
  inv1  gate1409(.a(G739), .O(gate247inter8));
  nand2 gate1410(.a(gate247inter8), .b(gate247inter7), .O(gate247inter9));
  nand2 gate1411(.a(s_123), .b(gate247inter3), .O(gate247inter10));
  nor2  gate1412(.a(gate247inter10), .b(gate247inter9), .O(gate247inter11));
  nor2  gate1413(.a(gate247inter11), .b(gate247inter6), .O(gate247inter12));
  nand2 gate1414(.a(gate247inter12), .b(gate247inter1), .O(G760));

  xor2  gate1303(.a(G739), .b(G727), .O(gate248inter0));
  nand2 gate1304(.a(gate248inter0), .b(s_108), .O(gate248inter1));
  and2  gate1305(.a(G739), .b(G727), .O(gate248inter2));
  inv1  gate1306(.a(s_108), .O(gate248inter3));
  inv1  gate1307(.a(s_109), .O(gate248inter4));
  nand2 gate1308(.a(gate248inter4), .b(gate248inter3), .O(gate248inter5));
  nor2  gate1309(.a(gate248inter5), .b(gate248inter2), .O(gate248inter6));
  inv1  gate1310(.a(G727), .O(gate248inter7));
  inv1  gate1311(.a(G739), .O(gate248inter8));
  nand2 gate1312(.a(gate248inter8), .b(gate248inter7), .O(gate248inter9));
  nand2 gate1313(.a(s_109), .b(gate248inter3), .O(gate248inter10));
  nor2  gate1314(.a(gate248inter10), .b(gate248inter9), .O(gate248inter11));
  nor2  gate1315(.a(gate248inter11), .b(gate248inter6), .O(gate248inter12));
  nand2 gate1316(.a(gate248inter12), .b(gate248inter1), .O(G761));
nand2 gate249( .a(G254), .b(G742), .O(G762) );

  xor2  gate1499(.a(G742), .b(G706), .O(gate250inter0));
  nand2 gate1500(.a(gate250inter0), .b(s_136), .O(gate250inter1));
  and2  gate1501(.a(G742), .b(G706), .O(gate250inter2));
  inv1  gate1502(.a(s_136), .O(gate250inter3));
  inv1  gate1503(.a(s_137), .O(gate250inter4));
  nand2 gate1504(.a(gate250inter4), .b(gate250inter3), .O(gate250inter5));
  nor2  gate1505(.a(gate250inter5), .b(gate250inter2), .O(gate250inter6));
  inv1  gate1506(.a(G706), .O(gate250inter7));
  inv1  gate1507(.a(G742), .O(gate250inter8));
  nand2 gate1508(.a(gate250inter8), .b(gate250inter7), .O(gate250inter9));
  nand2 gate1509(.a(s_137), .b(gate250inter3), .O(gate250inter10));
  nor2  gate1510(.a(gate250inter10), .b(gate250inter9), .O(gate250inter11));
  nor2  gate1511(.a(gate250inter11), .b(gate250inter6), .O(gate250inter12));
  nand2 gate1512(.a(gate250inter12), .b(gate250inter1), .O(G763));

  xor2  gate1583(.a(G745), .b(G257), .O(gate251inter0));
  nand2 gate1584(.a(gate251inter0), .b(s_148), .O(gate251inter1));
  and2  gate1585(.a(G745), .b(G257), .O(gate251inter2));
  inv1  gate1586(.a(s_148), .O(gate251inter3));
  inv1  gate1587(.a(s_149), .O(gate251inter4));
  nand2 gate1588(.a(gate251inter4), .b(gate251inter3), .O(gate251inter5));
  nor2  gate1589(.a(gate251inter5), .b(gate251inter2), .O(gate251inter6));
  inv1  gate1590(.a(G257), .O(gate251inter7));
  inv1  gate1591(.a(G745), .O(gate251inter8));
  nand2 gate1592(.a(gate251inter8), .b(gate251inter7), .O(gate251inter9));
  nand2 gate1593(.a(s_149), .b(gate251inter3), .O(gate251inter10));
  nor2  gate1594(.a(gate251inter10), .b(gate251inter9), .O(gate251inter11));
  nor2  gate1595(.a(gate251inter11), .b(gate251inter6), .O(gate251inter12));
  nand2 gate1596(.a(gate251inter12), .b(gate251inter1), .O(G764));

  xor2  gate2115(.a(G745), .b(G709), .O(gate252inter0));
  nand2 gate2116(.a(gate252inter0), .b(s_224), .O(gate252inter1));
  and2  gate2117(.a(G745), .b(G709), .O(gate252inter2));
  inv1  gate2118(.a(s_224), .O(gate252inter3));
  inv1  gate2119(.a(s_225), .O(gate252inter4));
  nand2 gate2120(.a(gate252inter4), .b(gate252inter3), .O(gate252inter5));
  nor2  gate2121(.a(gate252inter5), .b(gate252inter2), .O(gate252inter6));
  inv1  gate2122(.a(G709), .O(gate252inter7));
  inv1  gate2123(.a(G745), .O(gate252inter8));
  nand2 gate2124(.a(gate252inter8), .b(gate252inter7), .O(gate252inter9));
  nand2 gate2125(.a(s_225), .b(gate252inter3), .O(gate252inter10));
  nor2  gate2126(.a(gate252inter10), .b(gate252inter9), .O(gate252inter11));
  nor2  gate2127(.a(gate252inter11), .b(gate252inter6), .O(gate252inter12));
  nand2 gate2128(.a(gate252inter12), .b(gate252inter1), .O(G765));
nand2 gate253( .a(G260), .b(G748), .O(G766) );
nand2 gate254( .a(G712), .b(G748), .O(G767) );
nand2 gate255( .a(G263), .b(G751), .O(G768) );

  xor2  gate1695(.a(G751), .b(G715), .O(gate256inter0));
  nand2 gate1696(.a(gate256inter0), .b(s_164), .O(gate256inter1));
  and2  gate1697(.a(G751), .b(G715), .O(gate256inter2));
  inv1  gate1698(.a(s_164), .O(gate256inter3));
  inv1  gate1699(.a(s_165), .O(gate256inter4));
  nand2 gate1700(.a(gate256inter4), .b(gate256inter3), .O(gate256inter5));
  nor2  gate1701(.a(gate256inter5), .b(gate256inter2), .O(gate256inter6));
  inv1  gate1702(.a(G715), .O(gate256inter7));
  inv1  gate1703(.a(G751), .O(gate256inter8));
  nand2 gate1704(.a(gate256inter8), .b(gate256inter7), .O(gate256inter9));
  nand2 gate1705(.a(s_165), .b(gate256inter3), .O(gate256inter10));
  nor2  gate1706(.a(gate256inter10), .b(gate256inter9), .O(gate256inter11));
  nor2  gate1707(.a(gate256inter11), .b(gate256inter6), .O(gate256inter12));
  nand2 gate1708(.a(gate256inter12), .b(gate256inter1), .O(G769));
nand2 gate257( .a(G754), .b(G755), .O(G770) );
nand2 gate258( .a(G756), .b(G757), .O(G773) );
nand2 gate259( .a(G758), .b(G759), .O(G776) );

  xor2  gate757(.a(G761), .b(G760), .O(gate260inter0));
  nand2 gate758(.a(gate260inter0), .b(s_30), .O(gate260inter1));
  and2  gate759(.a(G761), .b(G760), .O(gate260inter2));
  inv1  gate760(.a(s_30), .O(gate260inter3));
  inv1  gate761(.a(s_31), .O(gate260inter4));
  nand2 gate762(.a(gate260inter4), .b(gate260inter3), .O(gate260inter5));
  nor2  gate763(.a(gate260inter5), .b(gate260inter2), .O(gate260inter6));
  inv1  gate764(.a(G760), .O(gate260inter7));
  inv1  gate765(.a(G761), .O(gate260inter8));
  nand2 gate766(.a(gate260inter8), .b(gate260inter7), .O(gate260inter9));
  nand2 gate767(.a(s_31), .b(gate260inter3), .O(gate260inter10));
  nor2  gate768(.a(gate260inter10), .b(gate260inter9), .O(gate260inter11));
  nor2  gate769(.a(gate260inter11), .b(gate260inter6), .O(gate260inter12));
  nand2 gate770(.a(gate260inter12), .b(gate260inter1), .O(G779));

  xor2  gate1219(.a(G763), .b(G762), .O(gate261inter0));
  nand2 gate1220(.a(gate261inter0), .b(s_96), .O(gate261inter1));
  and2  gate1221(.a(G763), .b(G762), .O(gate261inter2));
  inv1  gate1222(.a(s_96), .O(gate261inter3));
  inv1  gate1223(.a(s_97), .O(gate261inter4));
  nand2 gate1224(.a(gate261inter4), .b(gate261inter3), .O(gate261inter5));
  nor2  gate1225(.a(gate261inter5), .b(gate261inter2), .O(gate261inter6));
  inv1  gate1226(.a(G762), .O(gate261inter7));
  inv1  gate1227(.a(G763), .O(gate261inter8));
  nand2 gate1228(.a(gate261inter8), .b(gate261inter7), .O(gate261inter9));
  nand2 gate1229(.a(s_97), .b(gate261inter3), .O(gate261inter10));
  nor2  gate1230(.a(gate261inter10), .b(gate261inter9), .O(gate261inter11));
  nor2  gate1231(.a(gate261inter11), .b(gate261inter6), .O(gate261inter12));
  nand2 gate1232(.a(gate261inter12), .b(gate261inter1), .O(G782));
nand2 gate262( .a(G764), .b(G765), .O(G785) );

  xor2  gate1989(.a(G767), .b(G766), .O(gate263inter0));
  nand2 gate1990(.a(gate263inter0), .b(s_206), .O(gate263inter1));
  and2  gate1991(.a(G767), .b(G766), .O(gate263inter2));
  inv1  gate1992(.a(s_206), .O(gate263inter3));
  inv1  gate1993(.a(s_207), .O(gate263inter4));
  nand2 gate1994(.a(gate263inter4), .b(gate263inter3), .O(gate263inter5));
  nor2  gate1995(.a(gate263inter5), .b(gate263inter2), .O(gate263inter6));
  inv1  gate1996(.a(G766), .O(gate263inter7));
  inv1  gate1997(.a(G767), .O(gate263inter8));
  nand2 gate1998(.a(gate263inter8), .b(gate263inter7), .O(gate263inter9));
  nand2 gate1999(.a(s_207), .b(gate263inter3), .O(gate263inter10));
  nor2  gate2000(.a(gate263inter10), .b(gate263inter9), .O(gate263inter11));
  nor2  gate2001(.a(gate263inter11), .b(gate263inter6), .O(gate263inter12));
  nand2 gate2002(.a(gate263inter12), .b(gate263inter1), .O(G788));

  xor2  gate673(.a(G769), .b(G768), .O(gate264inter0));
  nand2 gate674(.a(gate264inter0), .b(s_18), .O(gate264inter1));
  and2  gate675(.a(G769), .b(G768), .O(gate264inter2));
  inv1  gate676(.a(s_18), .O(gate264inter3));
  inv1  gate677(.a(s_19), .O(gate264inter4));
  nand2 gate678(.a(gate264inter4), .b(gate264inter3), .O(gate264inter5));
  nor2  gate679(.a(gate264inter5), .b(gate264inter2), .O(gate264inter6));
  inv1  gate680(.a(G768), .O(gate264inter7));
  inv1  gate681(.a(G769), .O(gate264inter8));
  nand2 gate682(.a(gate264inter8), .b(gate264inter7), .O(gate264inter9));
  nand2 gate683(.a(s_19), .b(gate264inter3), .O(gate264inter10));
  nor2  gate684(.a(gate264inter10), .b(gate264inter9), .O(gate264inter11));
  nor2  gate685(.a(gate264inter11), .b(gate264inter6), .O(gate264inter12));
  nand2 gate686(.a(gate264inter12), .b(gate264inter1), .O(G791));
nand2 gate265( .a(G642), .b(G770), .O(G794) );
nand2 gate266( .a(G645), .b(G773), .O(G797) );

  xor2  gate729(.a(G776), .b(G648), .O(gate267inter0));
  nand2 gate730(.a(gate267inter0), .b(s_26), .O(gate267inter1));
  and2  gate731(.a(G776), .b(G648), .O(gate267inter2));
  inv1  gate732(.a(s_26), .O(gate267inter3));
  inv1  gate733(.a(s_27), .O(gate267inter4));
  nand2 gate734(.a(gate267inter4), .b(gate267inter3), .O(gate267inter5));
  nor2  gate735(.a(gate267inter5), .b(gate267inter2), .O(gate267inter6));
  inv1  gate736(.a(G648), .O(gate267inter7));
  inv1  gate737(.a(G776), .O(gate267inter8));
  nand2 gate738(.a(gate267inter8), .b(gate267inter7), .O(gate267inter9));
  nand2 gate739(.a(s_27), .b(gate267inter3), .O(gate267inter10));
  nor2  gate740(.a(gate267inter10), .b(gate267inter9), .O(gate267inter11));
  nor2  gate741(.a(gate267inter11), .b(gate267inter6), .O(gate267inter12));
  nand2 gate742(.a(gate267inter12), .b(gate267inter1), .O(G800));
nand2 gate268( .a(G651), .b(G779), .O(G803) );
nand2 gate269( .a(G654), .b(G782), .O(G806) );
nand2 gate270( .a(G657), .b(G785), .O(G809) );

  xor2  gate2129(.a(G788), .b(G660), .O(gate271inter0));
  nand2 gate2130(.a(gate271inter0), .b(s_226), .O(gate271inter1));
  and2  gate2131(.a(G788), .b(G660), .O(gate271inter2));
  inv1  gate2132(.a(s_226), .O(gate271inter3));
  inv1  gate2133(.a(s_227), .O(gate271inter4));
  nand2 gate2134(.a(gate271inter4), .b(gate271inter3), .O(gate271inter5));
  nor2  gate2135(.a(gate271inter5), .b(gate271inter2), .O(gate271inter6));
  inv1  gate2136(.a(G660), .O(gate271inter7));
  inv1  gate2137(.a(G788), .O(gate271inter8));
  nand2 gate2138(.a(gate271inter8), .b(gate271inter7), .O(gate271inter9));
  nand2 gate2139(.a(s_227), .b(gate271inter3), .O(gate271inter10));
  nor2  gate2140(.a(gate271inter10), .b(gate271inter9), .O(gate271inter11));
  nor2  gate2141(.a(gate271inter11), .b(gate271inter6), .O(gate271inter12));
  nand2 gate2142(.a(gate271inter12), .b(gate271inter1), .O(G812));
nand2 gate272( .a(G663), .b(G791), .O(G815) );

  xor2  gate841(.a(G794), .b(G642), .O(gate273inter0));
  nand2 gate842(.a(gate273inter0), .b(s_42), .O(gate273inter1));
  and2  gate843(.a(G794), .b(G642), .O(gate273inter2));
  inv1  gate844(.a(s_42), .O(gate273inter3));
  inv1  gate845(.a(s_43), .O(gate273inter4));
  nand2 gate846(.a(gate273inter4), .b(gate273inter3), .O(gate273inter5));
  nor2  gate847(.a(gate273inter5), .b(gate273inter2), .O(gate273inter6));
  inv1  gate848(.a(G642), .O(gate273inter7));
  inv1  gate849(.a(G794), .O(gate273inter8));
  nand2 gate850(.a(gate273inter8), .b(gate273inter7), .O(gate273inter9));
  nand2 gate851(.a(s_43), .b(gate273inter3), .O(gate273inter10));
  nor2  gate852(.a(gate273inter10), .b(gate273inter9), .O(gate273inter11));
  nor2  gate853(.a(gate273inter11), .b(gate273inter6), .O(gate273inter12));
  nand2 gate854(.a(gate273inter12), .b(gate273inter1), .O(G818));

  xor2  gate2157(.a(G794), .b(G770), .O(gate274inter0));
  nand2 gate2158(.a(gate274inter0), .b(s_230), .O(gate274inter1));
  and2  gate2159(.a(G794), .b(G770), .O(gate274inter2));
  inv1  gate2160(.a(s_230), .O(gate274inter3));
  inv1  gate2161(.a(s_231), .O(gate274inter4));
  nand2 gate2162(.a(gate274inter4), .b(gate274inter3), .O(gate274inter5));
  nor2  gate2163(.a(gate274inter5), .b(gate274inter2), .O(gate274inter6));
  inv1  gate2164(.a(G770), .O(gate274inter7));
  inv1  gate2165(.a(G794), .O(gate274inter8));
  nand2 gate2166(.a(gate274inter8), .b(gate274inter7), .O(gate274inter9));
  nand2 gate2167(.a(s_231), .b(gate274inter3), .O(gate274inter10));
  nor2  gate2168(.a(gate274inter10), .b(gate274inter9), .O(gate274inter11));
  nor2  gate2169(.a(gate274inter11), .b(gate274inter6), .O(gate274inter12));
  nand2 gate2170(.a(gate274inter12), .b(gate274inter1), .O(G819));
nand2 gate275( .a(G645), .b(G797), .O(G820) );
nand2 gate276( .a(G773), .b(G797), .O(G821) );
nand2 gate277( .a(G648), .b(G800), .O(G822) );

  xor2  gate2087(.a(G800), .b(G776), .O(gate278inter0));
  nand2 gate2088(.a(gate278inter0), .b(s_220), .O(gate278inter1));
  and2  gate2089(.a(G800), .b(G776), .O(gate278inter2));
  inv1  gate2090(.a(s_220), .O(gate278inter3));
  inv1  gate2091(.a(s_221), .O(gate278inter4));
  nand2 gate2092(.a(gate278inter4), .b(gate278inter3), .O(gate278inter5));
  nor2  gate2093(.a(gate278inter5), .b(gate278inter2), .O(gate278inter6));
  inv1  gate2094(.a(G776), .O(gate278inter7));
  inv1  gate2095(.a(G800), .O(gate278inter8));
  nand2 gate2096(.a(gate278inter8), .b(gate278inter7), .O(gate278inter9));
  nand2 gate2097(.a(s_221), .b(gate278inter3), .O(gate278inter10));
  nor2  gate2098(.a(gate278inter10), .b(gate278inter9), .O(gate278inter11));
  nor2  gate2099(.a(gate278inter11), .b(gate278inter6), .O(gate278inter12));
  nand2 gate2100(.a(gate278inter12), .b(gate278inter1), .O(G823));

  xor2  gate1751(.a(G803), .b(G651), .O(gate279inter0));
  nand2 gate1752(.a(gate279inter0), .b(s_172), .O(gate279inter1));
  and2  gate1753(.a(G803), .b(G651), .O(gate279inter2));
  inv1  gate1754(.a(s_172), .O(gate279inter3));
  inv1  gate1755(.a(s_173), .O(gate279inter4));
  nand2 gate1756(.a(gate279inter4), .b(gate279inter3), .O(gate279inter5));
  nor2  gate1757(.a(gate279inter5), .b(gate279inter2), .O(gate279inter6));
  inv1  gate1758(.a(G651), .O(gate279inter7));
  inv1  gate1759(.a(G803), .O(gate279inter8));
  nand2 gate1760(.a(gate279inter8), .b(gate279inter7), .O(gate279inter9));
  nand2 gate1761(.a(s_173), .b(gate279inter3), .O(gate279inter10));
  nor2  gate1762(.a(gate279inter10), .b(gate279inter9), .O(gate279inter11));
  nor2  gate1763(.a(gate279inter11), .b(gate279inter6), .O(gate279inter12));
  nand2 gate1764(.a(gate279inter12), .b(gate279inter1), .O(G824));
nand2 gate280( .a(G779), .b(G803), .O(G825) );
nand2 gate281( .a(G654), .b(G806), .O(G826) );
nand2 gate282( .a(G782), .b(G806), .O(G827) );
nand2 gate283( .a(G657), .b(G809), .O(G828) );
nand2 gate284( .a(G785), .b(G809), .O(G829) );
nand2 gate285( .a(G660), .b(G812), .O(G830) );

  xor2  gate1205(.a(G812), .b(G788), .O(gate286inter0));
  nand2 gate1206(.a(gate286inter0), .b(s_94), .O(gate286inter1));
  and2  gate1207(.a(G812), .b(G788), .O(gate286inter2));
  inv1  gate1208(.a(s_94), .O(gate286inter3));
  inv1  gate1209(.a(s_95), .O(gate286inter4));
  nand2 gate1210(.a(gate286inter4), .b(gate286inter3), .O(gate286inter5));
  nor2  gate1211(.a(gate286inter5), .b(gate286inter2), .O(gate286inter6));
  inv1  gate1212(.a(G788), .O(gate286inter7));
  inv1  gate1213(.a(G812), .O(gate286inter8));
  nand2 gate1214(.a(gate286inter8), .b(gate286inter7), .O(gate286inter9));
  nand2 gate1215(.a(s_95), .b(gate286inter3), .O(gate286inter10));
  nor2  gate1216(.a(gate286inter10), .b(gate286inter9), .O(gate286inter11));
  nor2  gate1217(.a(gate286inter11), .b(gate286inter6), .O(gate286inter12));
  nand2 gate1218(.a(gate286inter12), .b(gate286inter1), .O(G831));
nand2 gate287( .a(G663), .b(G815), .O(G832) );
nand2 gate288( .a(G791), .b(G815), .O(G833) );
nand2 gate289( .a(G818), .b(G819), .O(G834) );
nand2 gate290( .a(G820), .b(G821), .O(G847) );

  xor2  gate1317(.a(G823), .b(G822), .O(gate291inter0));
  nand2 gate1318(.a(gate291inter0), .b(s_110), .O(gate291inter1));
  and2  gate1319(.a(G823), .b(G822), .O(gate291inter2));
  inv1  gate1320(.a(s_110), .O(gate291inter3));
  inv1  gate1321(.a(s_111), .O(gate291inter4));
  nand2 gate1322(.a(gate291inter4), .b(gate291inter3), .O(gate291inter5));
  nor2  gate1323(.a(gate291inter5), .b(gate291inter2), .O(gate291inter6));
  inv1  gate1324(.a(G822), .O(gate291inter7));
  inv1  gate1325(.a(G823), .O(gate291inter8));
  nand2 gate1326(.a(gate291inter8), .b(gate291inter7), .O(gate291inter9));
  nand2 gate1327(.a(s_111), .b(gate291inter3), .O(gate291inter10));
  nor2  gate1328(.a(gate291inter10), .b(gate291inter9), .O(gate291inter11));
  nor2  gate1329(.a(gate291inter11), .b(gate291inter6), .O(gate291inter12));
  nand2 gate1330(.a(gate291inter12), .b(gate291inter1), .O(G860));

  xor2  gate953(.a(G825), .b(G824), .O(gate292inter0));
  nand2 gate954(.a(gate292inter0), .b(s_58), .O(gate292inter1));
  and2  gate955(.a(G825), .b(G824), .O(gate292inter2));
  inv1  gate956(.a(s_58), .O(gate292inter3));
  inv1  gate957(.a(s_59), .O(gate292inter4));
  nand2 gate958(.a(gate292inter4), .b(gate292inter3), .O(gate292inter5));
  nor2  gate959(.a(gate292inter5), .b(gate292inter2), .O(gate292inter6));
  inv1  gate960(.a(G824), .O(gate292inter7));
  inv1  gate961(.a(G825), .O(gate292inter8));
  nand2 gate962(.a(gate292inter8), .b(gate292inter7), .O(gate292inter9));
  nand2 gate963(.a(s_59), .b(gate292inter3), .O(gate292inter10));
  nor2  gate964(.a(gate292inter10), .b(gate292inter9), .O(gate292inter11));
  nor2  gate965(.a(gate292inter11), .b(gate292inter6), .O(gate292inter12));
  nand2 gate966(.a(gate292inter12), .b(gate292inter1), .O(G873));
nand2 gate293( .a(G828), .b(G829), .O(G886) );
nand2 gate294( .a(G832), .b(G833), .O(G899) );

  xor2  gate1863(.a(G831), .b(G830), .O(gate295inter0));
  nand2 gate1864(.a(gate295inter0), .b(s_188), .O(gate295inter1));
  and2  gate1865(.a(G831), .b(G830), .O(gate295inter2));
  inv1  gate1866(.a(s_188), .O(gate295inter3));
  inv1  gate1867(.a(s_189), .O(gate295inter4));
  nand2 gate1868(.a(gate295inter4), .b(gate295inter3), .O(gate295inter5));
  nor2  gate1869(.a(gate295inter5), .b(gate295inter2), .O(gate295inter6));
  inv1  gate1870(.a(G830), .O(gate295inter7));
  inv1  gate1871(.a(G831), .O(gate295inter8));
  nand2 gate1872(.a(gate295inter8), .b(gate295inter7), .O(gate295inter9));
  nand2 gate1873(.a(s_189), .b(gate295inter3), .O(gate295inter10));
  nor2  gate1874(.a(gate295inter10), .b(gate295inter9), .O(gate295inter11));
  nor2  gate1875(.a(gate295inter11), .b(gate295inter6), .O(gate295inter12));
  nand2 gate1876(.a(gate295inter12), .b(gate295inter1), .O(G912));
nand2 gate296( .a(G826), .b(G827), .O(G925) );
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );
nand2 gate387( .a(G1), .b(G1036), .O(G1132) );

  xor2  gate1065(.a(G1039), .b(G2), .O(gate388inter0));
  nand2 gate1066(.a(gate388inter0), .b(s_74), .O(gate388inter1));
  and2  gate1067(.a(G1039), .b(G2), .O(gate388inter2));
  inv1  gate1068(.a(s_74), .O(gate388inter3));
  inv1  gate1069(.a(s_75), .O(gate388inter4));
  nand2 gate1070(.a(gate388inter4), .b(gate388inter3), .O(gate388inter5));
  nor2  gate1071(.a(gate388inter5), .b(gate388inter2), .O(gate388inter6));
  inv1  gate1072(.a(G2), .O(gate388inter7));
  inv1  gate1073(.a(G1039), .O(gate388inter8));
  nand2 gate1074(.a(gate388inter8), .b(gate388inter7), .O(gate388inter9));
  nand2 gate1075(.a(s_75), .b(gate388inter3), .O(gate388inter10));
  nor2  gate1076(.a(gate388inter10), .b(gate388inter9), .O(gate388inter11));
  nor2  gate1077(.a(gate388inter11), .b(gate388inter6), .O(gate388inter12));
  nand2 gate1078(.a(gate388inter12), .b(gate388inter1), .O(G1135));
nand2 gate389( .a(G3), .b(G1042), .O(G1138) );

  xor2  gate1961(.a(G1045), .b(G4), .O(gate390inter0));
  nand2 gate1962(.a(gate390inter0), .b(s_202), .O(gate390inter1));
  and2  gate1963(.a(G1045), .b(G4), .O(gate390inter2));
  inv1  gate1964(.a(s_202), .O(gate390inter3));
  inv1  gate1965(.a(s_203), .O(gate390inter4));
  nand2 gate1966(.a(gate390inter4), .b(gate390inter3), .O(gate390inter5));
  nor2  gate1967(.a(gate390inter5), .b(gate390inter2), .O(gate390inter6));
  inv1  gate1968(.a(G4), .O(gate390inter7));
  inv1  gate1969(.a(G1045), .O(gate390inter8));
  nand2 gate1970(.a(gate390inter8), .b(gate390inter7), .O(gate390inter9));
  nand2 gate1971(.a(s_203), .b(gate390inter3), .O(gate390inter10));
  nor2  gate1972(.a(gate390inter10), .b(gate390inter9), .O(gate390inter11));
  nor2  gate1973(.a(gate390inter11), .b(gate390inter6), .O(gate390inter12));
  nand2 gate1974(.a(gate390inter12), .b(gate390inter1), .O(G1141));
nand2 gate391( .a(G5), .b(G1048), .O(G1144) );
nand2 gate392( .a(G6), .b(G1051), .O(G1147) );
nand2 gate393( .a(G7), .b(G1054), .O(G1150) );

  xor2  gate561(.a(G1057), .b(G8), .O(gate394inter0));
  nand2 gate562(.a(gate394inter0), .b(s_2), .O(gate394inter1));
  and2  gate563(.a(G1057), .b(G8), .O(gate394inter2));
  inv1  gate564(.a(s_2), .O(gate394inter3));
  inv1  gate565(.a(s_3), .O(gate394inter4));
  nand2 gate566(.a(gate394inter4), .b(gate394inter3), .O(gate394inter5));
  nor2  gate567(.a(gate394inter5), .b(gate394inter2), .O(gate394inter6));
  inv1  gate568(.a(G8), .O(gate394inter7));
  inv1  gate569(.a(G1057), .O(gate394inter8));
  nand2 gate570(.a(gate394inter8), .b(gate394inter7), .O(gate394inter9));
  nand2 gate571(.a(s_3), .b(gate394inter3), .O(gate394inter10));
  nor2  gate572(.a(gate394inter10), .b(gate394inter9), .O(gate394inter11));
  nor2  gate573(.a(gate394inter11), .b(gate394inter6), .O(gate394inter12));
  nand2 gate574(.a(gate394inter12), .b(gate394inter1), .O(G1153));

  xor2  gate1079(.a(G1060), .b(G9), .O(gate395inter0));
  nand2 gate1080(.a(gate395inter0), .b(s_76), .O(gate395inter1));
  and2  gate1081(.a(G1060), .b(G9), .O(gate395inter2));
  inv1  gate1082(.a(s_76), .O(gate395inter3));
  inv1  gate1083(.a(s_77), .O(gate395inter4));
  nand2 gate1084(.a(gate395inter4), .b(gate395inter3), .O(gate395inter5));
  nor2  gate1085(.a(gate395inter5), .b(gate395inter2), .O(gate395inter6));
  inv1  gate1086(.a(G9), .O(gate395inter7));
  inv1  gate1087(.a(G1060), .O(gate395inter8));
  nand2 gate1088(.a(gate395inter8), .b(gate395inter7), .O(gate395inter9));
  nand2 gate1089(.a(s_77), .b(gate395inter3), .O(gate395inter10));
  nor2  gate1090(.a(gate395inter10), .b(gate395inter9), .O(gate395inter11));
  nor2  gate1091(.a(gate395inter11), .b(gate395inter6), .O(gate395inter12));
  nand2 gate1092(.a(gate395inter12), .b(gate395inter1), .O(G1156));
nand2 gate396( .a(G10), .b(G1063), .O(G1159) );
nand2 gate397( .a(G11), .b(G1066), .O(G1162) );
nand2 gate398( .a(G12), .b(G1069), .O(G1165) );
nand2 gate399( .a(G13), .b(G1072), .O(G1168) );
nand2 gate400( .a(G14), .b(G1075), .O(G1171) );
nand2 gate401( .a(G15), .b(G1078), .O(G1174) );
nand2 gate402( .a(G16), .b(G1081), .O(G1177) );
nand2 gate403( .a(G17), .b(G1084), .O(G1180) );
nand2 gate404( .a(G18), .b(G1087), .O(G1183) );

  xor2  gate1191(.a(G1090), .b(G19), .O(gate405inter0));
  nand2 gate1192(.a(gate405inter0), .b(s_92), .O(gate405inter1));
  and2  gate1193(.a(G1090), .b(G19), .O(gate405inter2));
  inv1  gate1194(.a(s_92), .O(gate405inter3));
  inv1  gate1195(.a(s_93), .O(gate405inter4));
  nand2 gate1196(.a(gate405inter4), .b(gate405inter3), .O(gate405inter5));
  nor2  gate1197(.a(gate405inter5), .b(gate405inter2), .O(gate405inter6));
  inv1  gate1198(.a(G19), .O(gate405inter7));
  inv1  gate1199(.a(G1090), .O(gate405inter8));
  nand2 gate1200(.a(gate405inter8), .b(gate405inter7), .O(gate405inter9));
  nand2 gate1201(.a(s_93), .b(gate405inter3), .O(gate405inter10));
  nor2  gate1202(.a(gate405inter10), .b(gate405inter9), .O(gate405inter11));
  nor2  gate1203(.a(gate405inter11), .b(gate405inter6), .O(gate405inter12));
  nand2 gate1204(.a(gate405inter12), .b(gate405inter1), .O(G1186));

  xor2  gate2101(.a(G1093), .b(G20), .O(gate406inter0));
  nand2 gate2102(.a(gate406inter0), .b(s_222), .O(gate406inter1));
  and2  gate2103(.a(G1093), .b(G20), .O(gate406inter2));
  inv1  gate2104(.a(s_222), .O(gate406inter3));
  inv1  gate2105(.a(s_223), .O(gate406inter4));
  nand2 gate2106(.a(gate406inter4), .b(gate406inter3), .O(gate406inter5));
  nor2  gate2107(.a(gate406inter5), .b(gate406inter2), .O(gate406inter6));
  inv1  gate2108(.a(G20), .O(gate406inter7));
  inv1  gate2109(.a(G1093), .O(gate406inter8));
  nand2 gate2110(.a(gate406inter8), .b(gate406inter7), .O(gate406inter9));
  nand2 gate2111(.a(s_223), .b(gate406inter3), .O(gate406inter10));
  nor2  gate2112(.a(gate406inter10), .b(gate406inter9), .O(gate406inter11));
  nor2  gate2113(.a(gate406inter11), .b(gate406inter6), .O(gate406inter12));
  nand2 gate2114(.a(gate406inter12), .b(gate406inter1), .O(G1189));

  xor2  gate1373(.a(G1096), .b(G21), .O(gate407inter0));
  nand2 gate1374(.a(gate407inter0), .b(s_118), .O(gate407inter1));
  and2  gate1375(.a(G1096), .b(G21), .O(gate407inter2));
  inv1  gate1376(.a(s_118), .O(gate407inter3));
  inv1  gate1377(.a(s_119), .O(gate407inter4));
  nand2 gate1378(.a(gate407inter4), .b(gate407inter3), .O(gate407inter5));
  nor2  gate1379(.a(gate407inter5), .b(gate407inter2), .O(gate407inter6));
  inv1  gate1380(.a(G21), .O(gate407inter7));
  inv1  gate1381(.a(G1096), .O(gate407inter8));
  nand2 gate1382(.a(gate407inter8), .b(gate407inter7), .O(gate407inter9));
  nand2 gate1383(.a(s_119), .b(gate407inter3), .O(gate407inter10));
  nor2  gate1384(.a(gate407inter10), .b(gate407inter9), .O(gate407inter11));
  nor2  gate1385(.a(gate407inter11), .b(gate407inter6), .O(gate407inter12));
  nand2 gate1386(.a(gate407inter12), .b(gate407inter1), .O(G1192));

  xor2  gate1835(.a(G1099), .b(G22), .O(gate408inter0));
  nand2 gate1836(.a(gate408inter0), .b(s_184), .O(gate408inter1));
  and2  gate1837(.a(G1099), .b(G22), .O(gate408inter2));
  inv1  gate1838(.a(s_184), .O(gate408inter3));
  inv1  gate1839(.a(s_185), .O(gate408inter4));
  nand2 gate1840(.a(gate408inter4), .b(gate408inter3), .O(gate408inter5));
  nor2  gate1841(.a(gate408inter5), .b(gate408inter2), .O(gate408inter6));
  inv1  gate1842(.a(G22), .O(gate408inter7));
  inv1  gate1843(.a(G1099), .O(gate408inter8));
  nand2 gate1844(.a(gate408inter8), .b(gate408inter7), .O(gate408inter9));
  nand2 gate1845(.a(s_185), .b(gate408inter3), .O(gate408inter10));
  nor2  gate1846(.a(gate408inter10), .b(gate408inter9), .O(gate408inter11));
  nor2  gate1847(.a(gate408inter11), .b(gate408inter6), .O(gate408inter12));
  nand2 gate1848(.a(gate408inter12), .b(gate408inter1), .O(G1195));

  xor2  gate1149(.a(G1102), .b(G23), .O(gate409inter0));
  nand2 gate1150(.a(gate409inter0), .b(s_86), .O(gate409inter1));
  and2  gate1151(.a(G1102), .b(G23), .O(gate409inter2));
  inv1  gate1152(.a(s_86), .O(gate409inter3));
  inv1  gate1153(.a(s_87), .O(gate409inter4));
  nand2 gate1154(.a(gate409inter4), .b(gate409inter3), .O(gate409inter5));
  nor2  gate1155(.a(gate409inter5), .b(gate409inter2), .O(gate409inter6));
  inv1  gate1156(.a(G23), .O(gate409inter7));
  inv1  gate1157(.a(G1102), .O(gate409inter8));
  nand2 gate1158(.a(gate409inter8), .b(gate409inter7), .O(gate409inter9));
  nand2 gate1159(.a(s_87), .b(gate409inter3), .O(gate409inter10));
  nor2  gate1160(.a(gate409inter10), .b(gate409inter9), .O(gate409inter11));
  nor2  gate1161(.a(gate409inter11), .b(gate409inter6), .O(gate409inter12));
  nand2 gate1162(.a(gate409inter12), .b(gate409inter1), .O(G1198));
nand2 gate410( .a(G24), .b(G1105), .O(G1201) );

  xor2  gate1177(.a(G1108), .b(G25), .O(gate411inter0));
  nand2 gate1178(.a(gate411inter0), .b(s_90), .O(gate411inter1));
  and2  gate1179(.a(G1108), .b(G25), .O(gate411inter2));
  inv1  gate1180(.a(s_90), .O(gate411inter3));
  inv1  gate1181(.a(s_91), .O(gate411inter4));
  nand2 gate1182(.a(gate411inter4), .b(gate411inter3), .O(gate411inter5));
  nor2  gate1183(.a(gate411inter5), .b(gate411inter2), .O(gate411inter6));
  inv1  gate1184(.a(G25), .O(gate411inter7));
  inv1  gate1185(.a(G1108), .O(gate411inter8));
  nand2 gate1186(.a(gate411inter8), .b(gate411inter7), .O(gate411inter9));
  nand2 gate1187(.a(s_91), .b(gate411inter3), .O(gate411inter10));
  nor2  gate1188(.a(gate411inter10), .b(gate411inter9), .O(gate411inter11));
  nor2  gate1189(.a(gate411inter11), .b(gate411inter6), .O(gate411inter12));
  nand2 gate1190(.a(gate411inter12), .b(gate411inter1), .O(G1204));

  xor2  gate1163(.a(G1111), .b(G26), .O(gate412inter0));
  nand2 gate1164(.a(gate412inter0), .b(s_88), .O(gate412inter1));
  and2  gate1165(.a(G1111), .b(G26), .O(gate412inter2));
  inv1  gate1166(.a(s_88), .O(gate412inter3));
  inv1  gate1167(.a(s_89), .O(gate412inter4));
  nand2 gate1168(.a(gate412inter4), .b(gate412inter3), .O(gate412inter5));
  nor2  gate1169(.a(gate412inter5), .b(gate412inter2), .O(gate412inter6));
  inv1  gate1170(.a(G26), .O(gate412inter7));
  inv1  gate1171(.a(G1111), .O(gate412inter8));
  nand2 gate1172(.a(gate412inter8), .b(gate412inter7), .O(gate412inter9));
  nand2 gate1173(.a(s_89), .b(gate412inter3), .O(gate412inter10));
  nor2  gate1174(.a(gate412inter10), .b(gate412inter9), .O(gate412inter11));
  nor2  gate1175(.a(gate412inter11), .b(gate412inter6), .O(gate412inter12));
  nand2 gate1176(.a(gate412inter12), .b(gate412inter1), .O(G1207));
nand2 gate413( .a(G27), .b(G1114), .O(G1210) );
nand2 gate414( .a(G28), .b(G1117), .O(G1213) );

  xor2  gate1457(.a(G1120), .b(G29), .O(gate415inter0));
  nand2 gate1458(.a(gate415inter0), .b(s_130), .O(gate415inter1));
  and2  gate1459(.a(G1120), .b(G29), .O(gate415inter2));
  inv1  gate1460(.a(s_130), .O(gate415inter3));
  inv1  gate1461(.a(s_131), .O(gate415inter4));
  nand2 gate1462(.a(gate415inter4), .b(gate415inter3), .O(gate415inter5));
  nor2  gate1463(.a(gate415inter5), .b(gate415inter2), .O(gate415inter6));
  inv1  gate1464(.a(G29), .O(gate415inter7));
  inv1  gate1465(.a(G1120), .O(gate415inter8));
  nand2 gate1466(.a(gate415inter8), .b(gate415inter7), .O(gate415inter9));
  nand2 gate1467(.a(s_131), .b(gate415inter3), .O(gate415inter10));
  nor2  gate1468(.a(gate415inter10), .b(gate415inter9), .O(gate415inter11));
  nor2  gate1469(.a(gate415inter11), .b(gate415inter6), .O(gate415inter12));
  nand2 gate1470(.a(gate415inter12), .b(gate415inter1), .O(G1216));

  xor2  gate1877(.a(G1123), .b(G30), .O(gate416inter0));
  nand2 gate1878(.a(gate416inter0), .b(s_190), .O(gate416inter1));
  and2  gate1879(.a(G1123), .b(G30), .O(gate416inter2));
  inv1  gate1880(.a(s_190), .O(gate416inter3));
  inv1  gate1881(.a(s_191), .O(gate416inter4));
  nand2 gate1882(.a(gate416inter4), .b(gate416inter3), .O(gate416inter5));
  nor2  gate1883(.a(gate416inter5), .b(gate416inter2), .O(gate416inter6));
  inv1  gate1884(.a(G30), .O(gate416inter7));
  inv1  gate1885(.a(G1123), .O(gate416inter8));
  nand2 gate1886(.a(gate416inter8), .b(gate416inter7), .O(gate416inter9));
  nand2 gate1887(.a(s_191), .b(gate416inter3), .O(gate416inter10));
  nor2  gate1888(.a(gate416inter10), .b(gate416inter9), .O(gate416inter11));
  nor2  gate1889(.a(gate416inter11), .b(gate416inter6), .O(gate416inter12));
  nand2 gate1890(.a(gate416inter12), .b(gate416inter1), .O(G1219));

  xor2  gate897(.a(G1126), .b(G31), .O(gate417inter0));
  nand2 gate898(.a(gate417inter0), .b(s_50), .O(gate417inter1));
  and2  gate899(.a(G1126), .b(G31), .O(gate417inter2));
  inv1  gate900(.a(s_50), .O(gate417inter3));
  inv1  gate901(.a(s_51), .O(gate417inter4));
  nand2 gate902(.a(gate417inter4), .b(gate417inter3), .O(gate417inter5));
  nor2  gate903(.a(gate417inter5), .b(gate417inter2), .O(gate417inter6));
  inv1  gate904(.a(G31), .O(gate417inter7));
  inv1  gate905(.a(G1126), .O(gate417inter8));
  nand2 gate906(.a(gate417inter8), .b(gate417inter7), .O(gate417inter9));
  nand2 gate907(.a(s_51), .b(gate417inter3), .O(gate417inter10));
  nor2  gate908(.a(gate417inter10), .b(gate417inter9), .O(gate417inter11));
  nor2  gate909(.a(gate417inter11), .b(gate417inter6), .O(gate417inter12));
  nand2 gate910(.a(gate417inter12), .b(gate417inter1), .O(G1222));
nand2 gate418( .a(G32), .b(G1129), .O(G1225) );
nand2 gate419( .a(G1), .b(G1132), .O(G1228) );
nand2 gate420( .a(G1036), .b(G1132), .O(G1229) );
nand2 gate421( .a(G2), .b(G1135), .O(G1230) );
nand2 gate422( .a(G1039), .b(G1135), .O(G1231) );
nand2 gate423( .a(G3), .b(G1138), .O(G1232) );
nand2 gate424( .a(G1042), .b(G1138), .O(G1233) );
nand2 gate425( .a(G4), .b(G1141), .O(G1234) );

  xor2  gate2003(.a(G1141), .b(G1045), .O(gate426inter0));
  nand2 gate2004(.a(gate426inter0), .b(s_208), .O(gate426inter1));
  and2  gate2005(.a(G1141), .b(G1045), .O(gate426inter2));
  inv1  gate2006(.a(s_208), .O(gate426inter3));
  inv1  gate2007(.a(s_209), .O(gate426inter4));
  nand2 gate2008(.a(gate426inter4), .b(gate426inter3), .O(gate426inter5));
  nor2  gate2009(.a(gate426inter5), .b(gate426inter2), .O(gate426inter6));
  inv1  gate2010(.a(G1045), .O(gate426inter7));
  inv1  gate2011(.a(G1141), .O(gate426inter8));
  nand2 gate2012(.a(gate426inter8), .b(gate426inter7), .O(gate426inter9));
  nand2 gate2013(.a(s_209), .b(gate426inter3), .O(gate426inter10));
  nor2  gate2014(.a(gate426inter10), .b(gate426inter9), .O(gate426inter11));
  nor2  gate2015(.a(gate426inter11), .b(gate426inter6), .O(gate426inter12));
  nand2 gate2016(.a(gate426inter12), .b(gate426inter1), .O(G1235));

  xor2  gate1037(.a(G1144), .b(G5), .O(gate427inter0));
  nand2 gate1038(.a(gate427inter0), .b(s_70), .O(gate427inter1));
  and2  gate1039(.a(G1144), .b(G5), .O(gate427inter2));
  inv1  gate1040(.a(s_70), .O(gate427inter3));
  inv1  gate1041(.a(s_71), .O(gate427inter4));
  nand2 gate1042(.a(gate427inter4), .b(gate427inter3), .O(gate427inter5));
  nor2  gate1043(.a(gate427inter5), .b(gate427inter2), .O(gate427inter6));
  inv1  gate1044(.a(G5), .O(gate427inter7));
  inv1  gate1045(.a(G1144), .O(gate427inter8));
  nand2 gate1046(.a(gate427inter8), .b(gate427inter7), .O(gate427inter9));
  nand2 gate1047(.a(s_71), .b(gate427inter3), .O(gate427inter10));
  nor2  gate1048(.a(gate427inter10), .b(gate427inter9), .O(gate427inter11));
  nor2  gate1049(.a(gate427inter11), .b(gate427inter6), .O(gate427inter12));
  nand2 gate1050(.a(gate427inter12), .b(gate427inter1), .O(G1236));
nand2 gate428( .a(G1048), .b(G1144), .O(G1237) );
nand2 gate429( .a(G6), .b(G1147), .O(G1238) );
nand2 gate430( .a(G1051), .b(G1147), .O(G1239) );
nand2 gate431( .a(G7), .b(G1150), .O(G1240) );
nand2 gate432( .a(G1054), .b(G1150), .O(G1241) );

  xor2  gate1737(.a(G1153), .b(G8), .O(gate433inter0));
  nand2 gate1738(.a(gate433inter0), .b(s_170), .O(gate433inter1));
  and2  gate1739(.a(G1153), .b(G8), .O(gate433inter2));
  inv1  gate1740(.a(s_170), .O(gate433inter3));
  inv1  gate1741(.a(s_171), .O(gate433inter4));
  nand2 gate1742(.a(gate433inter4), .b(gate433inter3), .O(gate433inter5));
  nor2  gate1743(.a(gate433inter5), .b(gate433inter2), .O(gate433inter6));
  inv1  gate1744(.a(G8), .O(gate433inter7));
  inv1  gate1745(.a(G1153), .O(gate433inter8));
  nand2 gate1746(.a(gate433inter8), .b(gate433inter7), .O(gate433inter9));
  nand2 gate1747(.a(s_171), .b(gate433inter3), .O(gate433inter10));
  nor2  gate1748(.a(gate433inter10), .b(gate433inter9), .O(gate433inter11));
  nor2  gate1749(.a(gate433inter11), .b(gate433inter6), .O(gate433inter12));
  nand2 gate1750(.a(gate433inter12), .b(gate433inter1), .O(G1242));

  xor2  gate1933(.a(G1153), .b(G1057), .O(gate434inter0));
  nand2 gate1934(.a(gate434inter0), .b(s_198), .O(gate434inter1));
  and2  gate1935(.a(G1153), .b(G1057), .O(gate434inter2));
  inv1  gate1936(.a(s_198), .O(gate434inter3));
  inv1  gate1937(.a(s_199), .O(gate434inter4));
  nand2 gate1938(.a(gate434inter4), .b(gate434inter3), .O(gate434inter5));
  nor2  gate1939(.a(gate434inter5), .b(gate434inter2), .O(gate434inter6));
  inv1  gate1940(.a(G1057), .O(gate434inter7));
  inv1  gate1941(.a(G1153), .O(gate434inter8));
  nand2 gate1942(.a(gate434inter8), .b(gate434inter7), .O(gate434inter9));
  nand2 gate1943(.a(s_199), .b(gate434inter3), .O(gate434inter10));
  nor2  gate1944(.a(gate434inter10), .b(gate434inter9), .O(gate434inter11));
  nor2  gate1945(.a(gate434inter11), .b(gate434inter6), .O(gate434inter12));
  nand2 gate1946(.a(gate434inter12), .b(gate434inter1), .O(G1243));
nand2 gate435( .a(G9), .b(G1156), .O(G1244) );

  xor2  gate1527(.a(G1156), .b(G1060), .O(gate436inter0));
  nand2 gate1528(.a(gate436inter0), .b(s_140), .O(gate436inter1));
  and2  gate1529(.a(G1156), .b(G1060), .O(gate436inter2));
  inv1  gate1530(.a(s_140), .O(gate436inter3));
  inv1  gate1531(.a(s_141), .O(gate436inter4));
  nand2 gate1532(.a(gate436inter4), .b(gate436inter3), .O(gate436inter5));
  nor2  gate1533(.a(gate436inter5), .b(gate436inter2), .O(gate436inter6));
  inv1  gate1534(.a(G1060), .O(gate436inter7));
  inv1  gate1535(.a(G1156), .O(gate436inter8));
  nand2 gate1536(.a(gate436inter8), .b(gate436inter7), .O(gate436inter9));
  nand2 gate1537(.a(s_141), .b(gate436inter3), .O(gate436inter10));
  nor2  gate1538(.a(gate436inter10), .b(gate436inter9), .O(gate436inter11));
  nor2  gate1539(.a(gate436inter11), .b(gate436inter6), .O(gate436inter12));
  nand2 gate1540(.a(gate436inter12), .b(gate436inter1), .O(G1245));

  xor2  gate1387(.a(G1159), .b(G10), .O(gate437inter0));
  nand2 gate1388(.a(gate437inter0), .b(s_120), .O(gate437inter1));
  and2  gate1389(.a(G1159), .b(G10), .O(gate437inter2));
  inv1  gate1390(.a(s_120), .O(gate437inter3));
  inv1  gate1391(.a(s_121), .O(gate437inter4));
  nand2 gate1392(.a(gate437inter4), .b(gate437inter3), .O(gate437inter5));
  nor2  gate1393(.a(gate437inter5), .b(gate437inter2), .O(gate437inter6));
  inv1  gate1394(.a(G10), .O(gate437inter7));
  inv1  gate1395(.a(G1159), .O(gate437inter8));
  nand2 gate1396(.a(gate437inter8), .b(gate437inter7), .O(gate437inter9));
  nand2 gate1397(.a(s_121), .b(gate437inter3), .O(gate437inter10));
  nor2  gate1398(.a(gate437inter10), .b(gate437inter9), .O(gate437inter11));
  nor2  gate1399(.a(gate437inter11), .b(gate437inter6), .O(gate437inter12));
  nand2 gate1400(.a(gate437inter12), .b(gate437inter1), .O(G1246));

  xor2  gate1555(.a(G1159), .b(G1063), .O(gate438inter0));
  nand2 gate1556(.a(gate438inter0), .b(s_144), .O(gate438inter1));
  and2  gate1557(.a(G1159), .b(G1063), .O(gate438inter2));
  inv1  gate1558(.a(s_144), .O(gate438inter3));
  inv1  gate1559(.a(s_145), .O(gate438inter4));
  nand2 gate1560(.a(gate438inter4), .b(gate438inter3), .O(gate438inter5));
  nor2  gate1561(.a(gate438inter5), .b(gate438inter2), .O(gate438inter6));
  inv1  gate1562(.a(G1063), .O(gate438inter7));
  inv1  gate1563(.a(G1159), .O(gate438inter8));
  nand2 gate1564(.a(gate438inter8), .b(gate438inter7), .O(gate438inter9));
  nand2 gate1565(.a(s_145), .b(gate438inter3), .O(gate438inter10));
  nor2  gate1566(.a(gate438inter10), .b(gate438inter9), .O(gate438inter11));
  nor2  gate1567(.a(gate438inter11), .b(gate438inter6), .O(gate438inter12));
  nand2 gate1568(.a(gate438inter12), .b(gate438inter1), .O(G1247));
nand2 gate439( .a(G11), .b(G1162), .O(G1248) );
nand2 gate440( .a(G1066), .b(G1162), .O(G1249) );
nand2 gate441( .a(G12), .b(G1165), .O(G1250) );
nand2 gate442( .a(G1069), .b(G1165), .O(G1251) );
nand2 gate443( .a(G13), .b(G1168), .O(G1252) );
nand2 gate444( .a(G1072), .b(G1168), .O(G1253) );
nand2 gate445( .a(G14), .b(G1171), .O(G1254) );
nand2 gate446( .a(G1075), .b(G1171), .O(G1255) );
nand2 gate447( .a(G15), .b(G1174), .O(G1256) );
nand2 gate448( .a(G1078), .b(G1174), .O(G1257) );
nand2 gate449( .a(G16), .b(G1177), .O(G1258) );
nand2 gate450( .a(G1081), .b(G1177), .O(G1259) );

  xor2  gate1107(.a(G1180), .b(G17), .O(gate451inter0));
  nand2 gate1108(.a(gate451inter0), .b(s_80), .O(gate451inter1));
  and2  gate1109(.a(G1180), .b(G17), .O(gate451inter2));
  inv1  gate1110(.a(s_80), .O(gate451inter3));
  inv1  gate1111(.a(s_81), .O(gate451inter4));
  nand2 gate1112(.a(gate451inter4), .b(gate451inter3), .O(gate451inter5));
  nor2  gate1113(.a(gate451inter5), .b(gate451inter2), .O(gate451inter6));
  inv1  gate1114(.a(G17), .O(gate451inter7));
  inv1  gate1115(.a(G1180), .O(gate451inter8));
  nand2 gate1116(.a(gate451inter8), .b(gate451inter7), .O(gate451inter9));
  nand2 gate1117(.a(s_81), .b(gate451inter3), .O(gate451inter10));
  nor2  gate1118(.a(gate451inter10), .b(gate451inter9), .O(gate451inter11));
  nor2  gate1119(.a(gate451inter11), .b(gate451inter6), .O(gate451inter12));
  nand2 gate1120(.a(gate451inter12), .b(gate451inter1), .O(G1260));
nand2 gate452( .a(G1084), .b(G1180), .O(G1261) );

  xor2  gate1807(.a(G1183), .b(G18), .O(gate453inter0));
  nand2 gate1808(.a(gate453inter0), .b(s_180), .O(gate453inter1));
  and2  gate1809(.a(G1183), .b(G18), .O(gate453inter2));
  inv1  gate1810(.a(s_180), .O(gate453inter3));
  inv1  gate1811(.a(s_181), .O(gate453inter4));
  nand2 gate1812(.a(gate453inter4), .b(gate453inter3), .O(gate453inter5));
  nor2  gate1813(.a(gate453inter5), .b(gate453inter2), .O(gate453inter6));
  inv1  gate1814(.a(G18), .O(gate453inter7));
  inv1  gate1815(.a(G1183), .O(gate453inter8));
  nand2 gate1816(.a(gate453inter8), .b(gate453inter7), .O(gate453inter9));
  nand2 gate1817(.a(s_181), .b(gate453inter3), .O(gate453inter10));
  nor2  gate1818(.a(gate453inter10), .b(gate453inter9), .O(gate453inter11));
  nor2  gate1819(.a(gate453inter11), .b(gate453inter6), .O(gate453inter12));
  nand2 gate1820(.a(gate453inter12), .b(gate453inter1), .O(G1262));
nand2 gate454( .a(G1087), .b(G1183), .O(G1263) );
nand2 gate455( .a(G19), .b(G1186), .O(G1264) );
nand2 gate456( .a(G1090), .b(G1186), .O(G1265) );
nand2 gate457( .a(G20), .b(G1189), .O(G1266) );
nand2 gate458( .a(G1093), .b(G1189), .O(G1267) );
nand2 gate459( .a(G21), .b(G1192), .O(G1268) );
nand2 gate460( .a(G1096), .b(G1192), .O(G1269) );
nand2 gate461( .a(G22), .b(G1195), .O(G1270) );
nand2 gate462( .a(G1099), .b(G1195), .O(G1271) );

  xor2  gate925(.a(G1198), .b(G23), .O(gate463inter0));
  nand2 gate926(.a(gate463inter0), .b(s_54), .O(gate463inter1));
  and2  gate927(.a(G1198), .b(G23), .O(gate463inter2));
  inv1  gate928(.a(s_54), .O(gate463inter3));
  inv1  gate929(.a(s_55), .O(gate463inter4));
  nand2 gate930(.a(gate463inter4), .b(gate463inter3), .O(gate463inter5));
  nor2  gate931(.a(gate463inter5), .b(gate463inter2), .O(gate463inter6));
  inv1  gate932(.a(G23), .O(gate463inter7));
  inv1  gate933(.a(G1198), .O(gate463inter8));
  nand2 gate934(.a(gate463inter8), .b(gate463inter7), .O(gate463inter9));
  nand2 gate935(.a(s_55), .b(gate463inter3), .O(gate463inter10));
  nor2  gate936(.a(gate463inter10), .b(gate463inter9), .O(gate463inter11));
  nor2  gate937(.a(gate463inter11), .b(gate463inter6), .O(gate463inter12));
  nand2 gate938(.a(gate463inter12), .b(gate463inter1), .O(G1272));
nand2 gate464( .a(G1102), .b(G1198), .O(G1273) );

  xor2  gate1625(.a(G1201), .b(G24), .O(gate465inter0));
  nand2 gate1626(.a(gate465inter0), .b(s_154), .O(gate465inter1));
  and2  gate1627(.a(G1201), .b(G24), .O(gate465inter2));
  inv1  gate1628(.a(s_154), .O(gate465inter3));
  inv1  gate1629(.a(s_155), .O(gate465inter4));
  nand2 gate1630(.a(gate465inter4), .b(gate465inter3), .O(gate465inter5));
  nor2  gate1631(.a(gate465inter5), .b(gate465inter2), .O(gate465inter6));
  inv1  gate1632(.a(G24), .O(gate465inter7));
  inv1  gate1633(.a(G1201), .O(gate465inter8));
  nand2 gate1634(.a(gate465inter8), .b(gate465inter7), .O(gate465inter9));
  nand2 gate1635(.a(s_155), .b(gate465inter3), .O(gate465inter10));
  nor2  gate1636(.a(gate465inter10), .b(gate465inter9), .O(gate465inter11));
  nor2  gate1637(.a(gate465inter11), .b(gate465inter6), .O(gate465inter12));
  nand2 gate1638(.a(gate465inter12), .b(gate465inter1), .O(G1274));
nand2 gate466( .a(G1105), .b(G1201), .O(G1275) );

  xor2  gate1121(.a(G1204), .b(G25), .O(gate467inter0));
  nand2 gate1122(.a(gate467inter0), .b(s_82), .O(gate467inter1));
  and2  gate1123(.a(G1204), .b(G25), .O(gate467inter2));
  inv1  gate1124(.a(s_82), .O(gate467inter3));
  inv1  gate1125(.a(s_83), .O(gate467inter4));
  nand2 gate1126(.a(gate467inter4), .b(gate467inter3), .O(gate467inter5));
  nor2  gate1127(.a(gate467inter5), .b(gate467inter2), .O(gate467inter6));
  inv1  gate1128(.a(G25), .O(gate467inter7));
  inv1  gate1129(.a(G1204), .O(gate467inter8));
  nand2 gate1130(.a(gate467inter8), .b(gate467inter7), .O(gate467inter9));
  nand2 gate1131(.a(s_83), .b(gate467inter3), .O(gate467inter10));
  nor2  gate1132(.a(gate467inter10), .b(gate467inter9), .O(gate467inter11));
  nor2  gate1133(.a(gate467inter11), .b(gate467inter6), .O(gate467inter12));
  nand2 gate1134(.a(gate467inter12), .b(gate467inter1), .O(G1276));
nand2 gate468( .a(G1108), .b(G1204), .O(G1277) );
nand2 gate469( .a(G26), .b(G1207), .O(G1278) );

  xor2  gate1359(.a(G1207), .b(G1111), .O(gate470inter0));
  nand2 gate1360(.a(gate470inter0), .b(s_116), .O(gate470inter1));
  and2  gate1361(.a(G1207), .b(G1111), .O(gate470inter2));
  inv1  gate1362(.a(s_116), .O(gate470inter3));
  inv1  gate1363(.a(s_117), .O(gate470inter4));
  nand2 gate1364(.a(gate470inter4), .b(gate470inter3), .O(gate470inter5));
  nor2  gate1365(.a(gate470inter5), .b(gate470inter2), .O(gate470inter6));
  inv1  gate1366(.a(G1111), .O(gate470inter7));
  inv1  gate1367(.a(G1207), .O(gate470inter8));
  nand2 gate1368(.a(gate470inter8), .b(gate470inter7), .O(gate470inter9));
  nand2 gate1369(.a(s_117), .b(gate470inter3), .O(gate470inter10));
  nor2  gate1370(.a(gate470inter10), .b(gate470inter9), .O(gate470inter11));
  nor2  gate1371(.a(gate470inter11), .b(gate470inter6), .O(gate470inter12));
  nand2 gate1372(.a(gate470inter12), .b(gate470inter1), .O(G1279));
nand2 gate471( .a(G27), .b(G1210), .O(G1280) );

  xor2  gate1975(.a(G1210), .b(G1114), .O(gate472inter0));
  nand2 gate1976(.a(gate472inter0), .b(s_204), .O(gate472inter1));
  and2  gate1977(.a(G1210), .b(G1114), .O(gate472inter2));
  inv1  gate1978(.a(s_204), .O(gate472inter3));
  inv1  gate1979(.a(s_205), .O(gate472inter4));
  nand2 gate1980(.a(gate472inter4), .b(gate472inter3), .O(gate472inter5));
  nor2  gate1981(.a(gate472inter5), .b(gate472inter2), .O(gate472inter6));
  inv1  gate1982(.a(G1114), .O(gate472inter7));
  inv1  gate1983(.a(G1210), .O(gate472inter8));
  nand2 gate1984(.a(gate472inter8), .b(gate472inter7), .O(gate472inter9));
  nand2 gate1985(.a(s_205), .b(gate472inter3), .O(gate472inter10));
  nor2  gate1986(.a(gate472inter10), .b(gate472inter9), .O(gate472inter11));
  nor2  gate1987(.a(gate472inter11), .b(gate472inter6), .O(gate472inter12));
  nand2 gate1988(.a(gate472inter12), .b(gate472inter1), .O(G1281));
nand2 gate473( .a(G28), .b(G1213), .O(G1282) );
nand2 gate474( .a(G1117), .b(G1213), .O(G1283) );
nand2 gate475( .a(G29), .b(G1216), .O(G1284) );
nand2 gate476( .a(G1120), .b(G1216), .O(G1285) );

  xor2  gate659(.a(G1219), .b(G30), .O(gate477inter0));
  nand2 gate660(.a(gate477inter0), .b(s_16), .O(gate477inter1));
  and2  gate661(.a(G1219), .b(G30), .O(gate477inter2));
  inv1  gate662(.a(s_16), .O(gate477inter3));
  inv1  gate663(.a(s_17), .O(gate477inter4));
  nand2 gate664(.a(gate477inter4), .b(gate477inter3), .O(gate477inter5));
  nor2  gate665(.a(gate477inter5), .b(gate477inter2), .O(gate477inter6));
  inv1  gate666(.a(G30), .O(gate477inter7));
  inv1  gate667(.a(G1219), .O(gate477inter8));
  nand2 gate668(.a(gate477inter8), .b(gate477inter7), .O(gate477inter9));
  nand2 gate669(.a(s_17), .b(gate477inter3), .O(gate477inter10));
  nor2  gate670(.a(gate477inter10), .b(gate477inter9), .O(gate477inter11));
  nor2  gate671(.a(gate477inter11), .b(gate477inter6), .O(gate477inter12));
  nand2 gate672(.a(gate477inter12), .b(gate477inter1), .O(G1286));
nand2 gate478( .a(G1123), .b(G1219), .O(G1287) );
nand2 gate479( .a(G31), .b(G1222), .O(G1288) );
nand2 gate480( .a(G1126), .b(G1222), .O(G1289) );
nand2 gate481( .a(G32), .b(G1225), .O(G1290) );
nand2 gate482( .a(G1129), .b(G1225), .O(G1291) );
nand2 gate483( .a(G1228), .b(G1229), .O(G1292) );

  xor2  gate1289(.a(G1231), .b(G1230), .O(gate484inter0));
  nand2 gate1290(.a(gate484inter0), .b(s_106), .O(gate484inter1));
  and2  gate1291(.a(G1231), .b(G1230), .O(gate484inter2));
  inv1  gate1292(.a(s_106), .O(gate484inter3));
  inv1  gate1293(.a(s_107), .O(gate484inter4));
  nand2 gate1294(.a(gate484inter4), .b(gate484inter3), .O(gate484inter5));
  nor2  gate1295(.a(gate484inter5), .b(gate484inter2), .O(gate484inter6));
  inv1  gate1296(.a(G1230), .O(gate484inter7));
  inv1  gate1297(.a(G1231), .O(gate484inter8));
  nand2 gate1298(.a(gate484inter8), .b(gate484inter7), .O(gate484inter9));
  nand2 gate1299(.a(s_107), .b(gate484inter3), .O(gate484inter10));
  nor2  gate1300(.a(gate484inter10), .b(gate484inter9), .O(gate484inter11));
  nor2  gate1301(.a(gate484inter11), .b(gate484inter6), .O(gate484inter12));
  nand2 gate1302(.a(gate484inter12), .b(gate484inter1), .O(G1293));
nand2 gate485( .a(G1232), .b(G1233), .O(G1294) );
nand2 gate486( .a(G1234), .b(G1235), .O(G1295) );
nand2 gate487( .a(G1236), .b(G1237), .O(G1296) );

  xor2  gate1513(.a(G1239), .b(G1238), .O(gate488inter0));
  nand2 gate1514(.a(gate488inter0), .b(s_138), .O(gate488inter1));
  and2  gate1515(.a(G1239), .b(G1238), .O(gate488inter2));
  inv1  gate1516(.a(s_138), .O(gate488inter3));
  inv1  gate1517(.a(s_139), .O(gate488inter4));
  nand2 gate1518(.a(gate488inter4), .b(gate488inter3), .O(gate488inter5));
  nor2  gate1519(.a(gate488inter5), .b(gate488inter2), .O(gate488inter6));
  inv1  gate1520(.a(G1238), .O(gate488inter7));
  inv1  gate1521(.a(G1239), .O(gate488inter8));
  nand2 gate1522(.a(gate488inter8), .b(gate488inter7), .O(gate488inter9));
  nand2 gate1523(.a(s_139), .b(gate488inter3), .O(gate488inter10));
  nor2  gate1524(.a(gate488inter10), .b(gate488inter9), .O(gate488inter11));
  nor2  gate1525(.a(gate488inter11), .b(gate488inter6), .O(gate488inter12));
  nand2 gate1526(.a(gate488inter12), .b(gate488inter1), .O(G1297));

  xor2  gate1247(.a(G1241), .b(G1240), .O(gate489inter0));
  nand2 gate1248(.a(gate489inter0), .b(s_100), .O(gate489inter1));
  and2  gate1249(.a(G1241), .b(G1240), .O(gate489inter2));
  inv1  gate1250(.a(s_100), .O(gate489inter3));
  inv1  gate1251(.a(s_101), .O(gate489inter4));
  nand2 gate1252(.a(gate489inter4), .b(gate489inter3), .O(gate489inter5));
  nor2  gate1253(.a(gate489inter5), .b(gate489inter2), .O(gate489inter6));
  inv1  gate1254(.a(G1240), .O(gate489inter7));
  inv1  gate1255(.a(G1241), .O(gate489inter8));
  nand2 gate1256(.a(gate489inter8), .b(gate489inter7), .O(gate489inter9));
  nand2 gate1257(.a(s_101), .b(gate489inter3), .O(gate489inter10));
  nor2  gate1258(.a(gate489inter10), .b(gate489inter9), .O(gate489inter11));
  nor2  gate1259(.a(gate489inter11), .b(gate489inter6), .O(gate489inter12));
  nand2 gate1260(.a(gate489inter12), .b(gate489inter1), .O(G1298));
nand2 gate490( .a(G1242), .b(G1243), .O(G1299) );
nand2 gate491( .a(G1244), .b(G1245), .O(G1300) );
nand2 gate492( .a(G1246), .b(G1247), .O(G1301) );
nand2 gate493( .a(G1248), .b(G1249), .O(G1302) );
nand2 gate494( .a(G1250), .b(G1251), .O(G1303) );
nand2 gate495( .a(G1252), .b(G1253), .O(G1304) );
nand2 gate496( .a(G1254), .b(G1255), .O(G1305) );
nand2 gate497( .a(G1256), .b(G1257), .O(G1306) );
nand2 gate498( .a(G1258), .b(G1259), .O(G1307) );

  xor2  gate855(.a(G1261), .b(G1260), .O(gate499inter0));
  nand2 gate856(.a(gate499inter0), .b(s_44), .O(gate499inter1));
  and2  gate857(.a(G1261), .b(G1260), .O(gate499inter2));
  inv1  gate858(.a(s_44), .O(gate499inter3));
  inv1  gate859(.a(s_45), .O(gate499inter4));
  nand2 gate860(.a(gate499inter4), .b(gate499inter3), .O(gate499inter5));
  nor2  gate861(.a(gate499inter5), .b(gate499inter2), .O(gate499inter6));
  inv1  gate862(.a(G1260), .O(gate499inter7));
  inv1  gate863(.a(G1261), .O(gate499inter8));
  nand2 gate864(.a(gate499inter8), .b(gate499inter7), .O(gate499inter9));
  nand2 gate865(.a(s_45), .b(gate499inter3), .O(gate499inter10));
  nor2  gate866(.a(gate499inter10), .b(gate499inter9), .O(gate499inter11));
  nor2  gate867(.a(gate499inter11), .b(gate499inter6), .O(gate499inter12));
  nand2 gate868(.a(gate499inter12), .b(gate499inter1), .O(G1308));

  xor2  gate645(.a(G1263), .b(G1262), .O(gate500inter0));
  nand2 gate646(.a(gate500inter0), .b(s_14), .O(gate500inter1));
  and2  gate647(.a(G1263), .b(G1262), .O(gate500inter2));
  inv1  gate648(.a(s_14), .O(gate500inter3));
  inv1  gate649(.a(s_15), .O(gate500inter4));
  nand2 gate650(.a(gate500inter4), .b(gate500inter3), .O(gate500inter5));
  nor2  gate651(.a(gate500inter5), .b(gate500inter2), .O(gate500inter6));
  inv1  gate652(.a(G1262), .O(gate500inter7));
  inv1  gate653(.a(G1263), .O(gate500inter8));
  nand2 gate654(.a(gate500inter8), .b(gate500inter7), .O(gate500inter9));
  nand2 gate655(.a(s_15), .b(gate500inter3), .O(gate500inter10));
  nor2  gate656(.a(gate500inter10), .b(gate500inter9), .O(gate500inter11));
  nor2  gate657(.a(gate500inter11), .b(gate500inter6), .O(gate500inter12));
  nand2 gate658(.a(gate500inter12), .b(gate500inter1), .O(G1309));
nand2 gate501( .a(G1264), .b(G1265), .O(G1310) );
nand2 gate502( .a(G1266), .b(G1267), .O(G1311) );
nand2 gate503( .a(G1268), .b(G1269), .O(G1312) );
nand2 gate504( .a(G1270), .b(G1271), .O(G1313) );
nand2 gate505( .a(G1272), .b(G1273), .O(G1314) );
nand2 gate506( .a(G1274), .b(G1275), .O(G1315) );
nand2 gate507( .a(G1276), .b(G1277), .O(G1316) );

  xor2  gate1471(.a(G1279), .b(G1278), .O(gate508inter0));
  nand2 gate1472(.a(gate508inter0), .b(s_132), .O(gate508inter1));
  and2  gate1473(.a(G1279), .b(G1278), .O(gate508inter2));
  inv1  gate1474(.a(s_132), .O(gate508inter3));
  inv1  gate1475(.a(s_133), .O(gate508inter4));
  nand2 gate1476(.a(gate508inter4), .b(gate508inter3), .O(gate508inter5));
  nor2  gate1477(.a(gate508inter5), .b(gate508inter2), .O(gate508inter6));
  inv1  gate1478(.a(G1278), .O(gate508inter7));
  inv1  gate1479(.a(G1279), .O(gate508inter8));
  nand2 gate1480(.a(gate508inter8), .b(gate508inter7), .O(gate508inter9));
  nand2 gate1481(.a(s_133), .b(gate508inter3), .O(gate508inter10));
  nor2  gate1482(.a(gate508inter10), .b(gate508inter9), .O(gate508inter11));
  nor2  gate1483(.a(gate508inter11), .b(gate508inter6), .O(gate508inter12));
  nand2 gate1484(.a(gate508inter12), .b(gate508inter1), .O(G1317));

  xor2  gate939(.a(G1281), .b(G1280), .O(gate509inter0));
  nand2 gate940(.a(gate509inter0), .b(s_56), .O(gate509inter1));
  and2  gate941(.a(G1281), .b(G1280), .O(gate509inter2));
  inv1  gate942(.a(s_56), .O(gate509inter3));
  inv1  gate943(.a(s_57), .O(gate509inter4));
  nand2 gate944(.a(gate509inter4), .b(gate509inter3), .O(gate509inter5));
  nor2  gate945(.a(gate509inter5), .b(gate509inter2), .O(gate509inter6));
  inv1  gate946(.a(G1280), .O(gate509inter7));
  inv1  gate947(.a(G1281), .O(gate509inter8));
  nand2 gate948(.a(gate509inter8), .b(gate509inter7), .O(gate509inter9));
  nand2 gate949(.a(s_57), .b(gate509inter3), .O(gate509inter10));
  nor2  gate950(.a(gate509inter10), .b(gate509inter9), .O(gate509inter11));
  nor2  gate951(.a(gate509inter11), .b(gate509inter6), .O(gate509inter12));
  nand2 gate952(.a(gate509inter12), .b(gate509inter1), .O(G1318));
nand2 gate510( .a(G1282), .b(G1283), .O(G1319) );
nand2 gate511( .a(G1284), .b(G1285), .O(G1320) );
nand2 gate512( .a(G1286), .b(G1287), .O(G1321) );
nand2 gate513( .a(G1288), .b(G1289), .O(G1322) );

  xor2  gate2073(.a(G1291), .b(G1290), .O(gate514inter0));
  nand2 gate2074(.a(gate514inter0), .b(s_218), .O(gate514inter1));
  and2  gate2075(.a(G1291), .b(G1290), .O(gate514inter2));
  inv1  gate2076(.a(s_218), .O(gate514inter3));
  inv1  gate2077(.a(s_219), .O(gate514inter4));
  nand2 gate2078(.a(gate514inter4), .b(gate514inter3), .O(gate514inter5));
  nor2  gate2079(.a(gate514inter5), .b(gate514inter2), .O(gate514inter6));
  inv1  gate2080(.a(G1290), .O(gate514inter7));
  inv1  gate2081(.a(G1291), .O(gate514inter8));
  nand2 gate2082(.a(gate514inter8), .b(gate514inter7), .O(gate514inter9));
  nand2 gate2083(.a(s_219), .b(gate514inter3), .O(gate514inter10));
  nor2  gate2084(.a(gate514inter10), .b(gate514inter9), .O(gate514inter11));
  nor2  gate2085(.a(gate514inter11), .b(gate514inter6), .O(gate514inter12));
  nand2 gate2086(.a(gate514inter12), .b(gate514inter1), .O(G1323));
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule