module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);

input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;//RE__PI;

input s_0,s_1;//RE__ALLOW(00,01,10,11);
input s_2,s_3;//RE__ALLOW(00,01,10,11);
input s_4,s_5;//RE__ALLOW(00,01,10,11);
input s_6,s_7;//RE__ALLOW(00,01,10,11);
input s_8,s_9;//RE__ALLOW(00,01,10,11);
input s_10,s_11;//RE__ALLOW(00,01,10,11);
input s_12,s_13;//RE__ALLOW(00,01,10,11);
input s_14,s_15;//RE__ALLOW(00,01,10,11);
input s_16,s_17;//RE__ALLOW(00,01,10,11);
input s_18,s_19;//RE__ALLOW(00,01,10,11);
input s_20,s_21;//RE__ALLOW(00,01,10,11);
input s_22,s_23;//RE__ALLOW(00,01,10,11);
input s_24,s_25;//RE__ALLOW(00,01,10,11);
input s_26,s_27;//RE__ALLOW(00,01,10,11);
input s_28,s_29;//RE__ALLOW(00,01,10,11);
input s_30,s_31;//RE__ALLOW(00,01,10,11);
input s_32,s_33;//RE__ALLOW(00,01,10,11);
input s_34,s_35;//RE__ALLOW(00,01,10,11);
input s_36,s_37;//RE__ALLOW(00,01,10,11);
input s_38,s_39;//RE__ALLOW(00,01,10,11);
input s_40,s_41;//RE__ALLOW(00,01,10,11);
input s_42,s_43;//RE__ALLOW(00,01,10,11);
input s_44,s_45;//RE__ALLOW(00,01,10,11);
input s_46,s_47;//RE__ALLOW(00,01,10,11);
input s_48,s_49;//RE__ALLOW(00,01,10,11);
input s_50,s_51;//RE__ALLOW(00,01,10,11);
input s_52,s_53;//RE__ALLOW(00,01,10,11);
input s_54,s_55;//RE__ALLOW(00,01,10,11);
input s_56,s_57;//RE__ALLOW(00,01,10,11);
input s_58,s_59;//RE__ALLOW(00,01,10,11);
input s_60,s_61;//RE__ALLOW(00,01,10,11);
input s_62,s_63;//RE__ALLOW(00,01,10,11);
input s_64,s_65;//RE__ALLOW(00,01,10,11);
input s_66,s_67;//RE__ALLOW(00,01,10,11);
input s_68,s_69;//RE__ALLOW(00,01,10,11);
input s_70,s_71;//RE__ALLOW(00,01,10,11);
input s_72,s_73;//RE__ALLOW(00,01,10,11);
input s_74,s_75;//RE__ALLOW(00,01,10,11);
input s_76,s_77;//RE__ALLOW(00,01,10,11);
input s_78,s_79;//RE__ALLOW(00,01,10,11);
input s_80,s_81;//RE__ALLOW(00,01,10,11);
input s_82,s_83;//RE__ALLOW(00,01,10,11);
input s_84,s_85;//RE__ALLOW(00,01,10,11);
input s_86,s_87;//RE__ALLOW(00,01,10,11);
input s_88,s_89;//RE__ALLOW(00,01,10,11);
input s_90,s_91;//RE__ALLOW(00,01,10,11);
input s_92,s_93;//RE__ALLOW(00,01,10,11);
input s_94,s_95;//RE__ALLOW(00,01,10,11);
input s_96,s_97;//RE__ALLOW(00,01,10,11);
input s_98,s_99;//RE__ALLOW(00,01,10,11);
input s_100,s_101;//RE__ALLOW(00,01,10,11);
input s_102,s_103;//RE__ALLOW(00,01,10,11);
input s_104,s_105;//RE__ALLOW(00,01,10,11);
input s_106,s_107;//RE__ALLOW(00,01,10,11);
input s_108,s_109;//RE__ALLOW(00,01,10,11);
input s_110,s_111;//RE__ALLOW(00,01,10,11);
input s_112,s_113;//RE__ALLOW(00,01,10,11);
input s_114,s_115;//RE__ALLOW(00,01,10,11);
input s_116,s_117;//RE__ALLOW(00,01,10,11);
input s_118,s_119;//RE__ALLOW(00,01,10,11);
input s_120,s_121;//RE__ALLOW(00,01,10,11);
input s_122,s_123;//RE__ALLOW(00,01,10,11);
input s_124,s_125;//RE__ALLOW(00,01,10,11);
input s_126,s_127;//RE__ALLOW(00,01,10,11);
input s_128,s_129;//RE__ALLOW(00,01,10,11);
input s_130,s_131;//RE__ALLOW(00,01,10,11);
input s_132,s_133;//RE__ALLOW(00,01,10,11);
input s_134,s_135;//RE__ALLOW(00,01,10,11);
input s_136,s_137;//RE__ALLOW(00,01,10,11);
input s_138,s_139;//RE__ALLOW(00,01,10,11);
input s_140,s_141;//RE__ALLOW(00,01,10,11);
input s_142,s_143;//RE__ALLOW(00,01,10,11);
input s_144,s_145;//RE__ALLOW(00,01,10,11);
input s_146,s_147;//RE__ALLOW(00,01,10,11);
input s_148,s_149;//RE__ALLOW(00,01,10,11);
input s_150,s_151;//RE__ALLOW(00,01,10,11);
input s_152,s_153;//RE__ALLOW(00,01,10,11);
input s_154,s_155;//RE__ALLOW(00,01,10,11);
input s_156,s_157;//RE__ALLOW(00,01,10,11);
input s_158,s_159;//RE__ALLOW(00,01,10,11);
input s_160,s_161;//RE__ALLOW(00,01,10,11);
input s_162,s_163;//RE__ALLOW(00,01,10,11);
input s_164,s_165;//RE__ALLOW(00,01,10,11);
input s_166,s_167;//RE__ALLOW(00,01,10,11);
input s_168,s_169;//RE__ALLOW(00,01,10,11);
input s_170,s_171;//RE__ALLOW(00,01,10,11);
input s_172,s_173;//RE__ALLOW(00,01,10,11);
input s_174,s_175;//RE__ALLOW(00,01,10,11);
input s_176,s_177;//RE__ALLOW(00,01,10,11);
input s_178,s_179;//RE__ALLOW(00,01,10,11);
input s_180,s_181;//RE__ALLOW(00,01,10,11);
input s_182,s_183;//RE__ALLOW(00,01,10,11);
input s_184,s_185;//RE__ALLOW(00,01,10,11);
input s_186,s_187;//RE__ALLOW(00,01,10,11);
input s_188,s_189;//RE__ALLOW(00,01,10,11);
input s_190,s_191;//RE__ALLOW(00,01,10,11);
input s_192,s_193;//RE__ALLOW(00,01,10,11);
input s_194,s_195;//RE__ALLOW(00,01,10,11);
input s_196,s_197;//RE__ALLOW(00,01,10,11);
input s_198,s_199;//RE__ALLOW(00,01,10,11);
input s_200,s_201;//RE__ALLOW(00,01,10,11);
input s_202,s_203;//RE__ALLOW(00,01,10,11);
input s_204,s_205;//RE__ALLOW(00,01,10,11);
input s_206,s_207;//RE__ALLOW(00,01,10,11);
input s_208,s_209;//RE__ALLOW(00,01,10,11);
input s_210,s_211;//RE__ALLOW(00,01,10,11);
input s_212,s_213;//RE__ALLOW(00,01,10,11);
input s_214,s_215;//RE__ALLOW(00,01,10,11);
input s_216,s_217;//RE__ALLOW(00,01,10,11);
input s_218,s_219;//RE__ALLOW(00,01,10,11);
input s_220,s_221;//RE__ALLOW(00,01,10,11);
input s_222,s_223;//RE__ALLOW(00,01,10,11);
input s_224,s_225;//RE__ALLOW(00,01,10,11);
input s_226,s_227;//RE__ALLOW(00,01,10,11);
input s_228,s_229;//RE__ALLOW(00,01,10,11);
input s_230,s_231;//RE__ALLOW(00,01,10,11);
input s_232,s_233;//RE__ALLOW(00,01,10,11);
input s_234,s_235;//RE__ALLOW(00,01,10,11);
input s_236,s_237;//RE__ALLOW(00,01,10,11);
input s_238,s_239;//RE__ALLOW(00,01,10,11);
input s_240,s_241;//RE__ALLOW(00,01,10,11);
input s_242,s_243;//RE__ALLOW(00,01,10,11);
input s_244,s_245;//RE__ALLOW(00,01,10,11);
input s_246,s_247;//RE__ALLOW(00,01,10,11);
input s_248,s_249;//RE__ALLOW(00,01,10,11);
input s_250,s_251;//RE__ALLOW(00,01,10,11);
input s_252,s_253;//RE__ALLOW(00,01,10,11);
input s_254,s_255;//RE__ALLOW(00,01,10,11);
input s_256,s_257;//RE__ALLOW(00,01,10,11);
input s_258,s_259;//RE__ALLOW(00,01,10,11);
input s_260,s_261;//RE__ALLOW(00,01,10,11);
input s_262,s_263;//RE__ALLOW(00,01,10,11);
input s_264,s_265;//RE__ALLOW(00,01,10,11);
input s_266,s_267;//RE__ALLOW(00,01,10,11);
input s_268,s_269;//RE__ALLOW(00,01,10,11);
input s_270,s_271;//RE__ALLOW(00,01,10,11);
input s_272,s_273;//RE__ALLOW(00,01,10,11);
input s_274,s_275;//RE__ALLOW(00,01,10,11);
input s_276,s_277;//RE__ALLOW(00,01,10,11);
input s_278,s_279;//RE__ALLOW(00,01,10,11);
input s_280,s_281;//RE__ALLOW(00,01,10,11);
input s_282,s_283;//RE__ALLOW(00,01,10,11);
input s_284,s_285;//RE__ALLOW(00,01,10,11);
input s_286,s_287;//RE__ALLOW(00,01,10,11);
input s_288,s_289;//RE__ALLOW(00,01,10,11);
input s_290,s_291;//RE__ALLOW(00,01,10,11);
input s_292,s_293;//RE__ALLOW(00,01,10,11);
input s_294,s_295;//RE__ALLOW(00,01,10,11);
input s_296,s_297;//RE__ALLOW(00,01,10,11);
input s_298,s_299;//RE__ALLOW(00,01,10,11);
input s_300,s_301;//RE__ALLOW(00,01,10,11);
input s_302,s_303;//RE__ALLOW(00,01,10,11);
input s_304,s_305;//RE__ALLOW(00,01,10,11);
input s_306,s_307;//RE__ALLOW(00,01,10,11);
input s_308,s_309;//RE__ALLOW(00,01,10,11);
input s_310,s_311;//RE__ALLOW(00,01,10,11);
input s_312,s_313;//RE__ALLOW(00,01,10,11);
input s_314,s_315;//RE__ALLOW(00,01,10,11);
input s_316,s_317;//RE__ALLOW(00,01,10,11);
input s_318,s_319;//RE__ALLOW(00,01,10,11);
input s_320,s_321;//RE__ALLOW(00,01,10,11);
input s_322,s_323;//RE__ALLOW(00,01,10,11);
input s_324,s_325;//RE__ALLOW(00,01,10,11);
input s_326,s_327;//RE__ALLOW(00,01,10,11);
input s_328,s_329;//RE__ALLOW(00,01,10,11);
input s_330,s_331;//RE__ALLOW(00,01,10,11);
input s_332,s_333;//RE__ALLOW(00,01,10,11);
input s_334,s_335;//RE__ALLOW(00,01,10,11);
input s_336,s_337;//RE__ALLOW(00,01,10,11);
input s_338,s_339;//RE__ALLOW(00,01,10,11);
input s_340,s_341;//RE__ALLOW(00,01,10,11);
input s_342,s_343;//RE__ALLOW(00,01,10,11);
input s_344,s_345;//RE__ALLOW(00,01,10,11);
input s_346,s_347;//RE__ALLOW(00,01,10,11);
input s_348,s_349;//RE__ALLOW(00,01,10,11);
input s_350,s_351;//RE__ALLOW(00,01,10,11);
input s_352,s_353;//RE__ALLOW(00,01,10,11);
input s_354,s_355;//RE__ALLOW(00,01,10,11);
input s_356,s_357;//RE__ALLOW(00,01,10,11);
input s_358,s_359;//RE__ALLOW(00,01,10,11);
input s_360,s_361;//RE__ALLOW(00,01,10,11);
input s_362,s_363;//RE__ALLOW(00,01,10,11);
input s_364,s_365;//RE__ALLOW(00,01,10,11);
input s_366,s_367;//RE__ALLOW(00,01,10,11);
input s_368,s_369;//RE__ALLOW(00,01,10,11);
input s_370,s_371;//RE__ALLOW(00,01,10,11);
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;

  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate55inter0, gate55inter1, gate55inter2, gate55inter3, gate55inter4, gate55inter5, gate55inter6, gate55inter7, gate55inter8, gate55inter9, gate55inter10, gate55inter11, gate55inter12, gate159inter0, gate159inter1, gate159inter2, gate159inter3, gate159inter4, gate159inter5, gate159inter6, gate159inter7, gate159inter8, gate159inter9, gate159inter10, gate159inter11, gate159inter12, gate207inter0, gate207inter1, gate207inter2, gate207inter3, gate207inter4, gate207inter5, gate207inter6, gate207inter7, gate207inter8, gate207inter9, gate207inter10, gate207inter11, gate207inter12, gate60inter0, gate60inter1, gate60inter2, gate60inter3, gate60inter4, gate60inter5, gate60inter6, gate60inter7, gate60inter8, gate60inter9, gate60inter10, gate60inter11, gate60inter12, gate94inter0, gate94inter1, gate94inter2, gate94inter3, gate94inter4, gate94inter5, gate94inter6, gate94inter7, gate94inter8, gate94inter9, gate94inter10, gate94inter11, gate94inter12, gate158inter0, gate158inter1, gate158inter2, gate158inter3, gate158inter4, gate158inter5, gate158inter6, gate158inter7, gate158inter8, gate158inter9, gate158inter10, gate158inter11, gate158inter12, gate19inter0, gate19inter1, gate19inter2, gate19inter3, gate19inter4, gate19inter5, gate19inter6, gate19inter7, gate19inter8, gate19inter9, gate19inter10, gate19inter11, gate19inter12, gate395inter0, gate395inter1, gate395inter2, gate395inter3, gate395inter4, gate395inter5, gate395inter6, gate395inter7, gate395inter8, gate395inter9, gate395inter10, gate395inter11, gate395inter12, gate129inter0, gate129inter1, gate129inter2, gate129inter3, gate129inter4, gate129inter5, gate129inter6, gate129inter7, gate129inter8, gate129inter9, gate129inter10, gate129inter11, gate129inter12, gate203inter0, gate203inter1, gate203inter2, gate203inter3, gate203inter4, gate203inter5, gate203inter6, gate203inter7, gate203inter8, gate203inter9, gate203inter10, gate203inter11, gate203inter12, gate222inter0, gate222inter1, gate222inter2, gate222inter3, gate222inter4, gate222inter5, gate222inter6, gate222inter7, gate222inter8, gate222inter9, gate222inter10, gate222inter11, gate222inter12, gate93inter0, gate93inter1, gate93inter2, gate93inter3, gate93inter4, gate93inter5, gate93inter6, gate93inter7, gate93inter8, gate93inter9, gate93inter10, gate93inter11, gate93inter12, gate392inter0, gate392inter1, gate392inter2, gate392inter3, gate392inter4, gate392inter5, gate392inter6, gate392inter7, gate392inter8, gate392inter9, gate392inter10, gate392inter11, gate392inter12, gate282inter0, gate282inter1, gate282inter2, gate282inter3, gate282inter4, gate282inter5, gate282inter6, gate282inter7, gate282inter8, gate282inter9, gate282inter10, gate282inter11, gate282inter12, gate211inter0, gate211inter1, gate211inter2, gate211inter3, gate211inter4, gate211inter5, gate211inter6, gate211inter7, gate211inter8, gate211inter9, gate211inter10, gate211inter11, gate211inter12, gate21inter0, gate21inter1, gate21inter2, gate21inter3, gate21inter4, gate21inter5, gate21inter6, gate21inter7, gate21inter8, gate21inter9, gate21inter10, gate21inter11, gate21inter12, gate210inter0, gate210inter1, gate210inter2, gate210inter3, gate210inter4, gate210inter5, gate210inter6, gate210inter7, gate210inter8, gate210inter9, gate210inter10, gate210inter11, gate210inter12, gate456inter0, gate456inter1, gate456inter2, gate456inter3, gate456inter4, gate456inter5, gate456inter6, gate456inter7, gate456inter8, gate456inter9, gate456inter10, gate456inter11, gate456inter12, gate118inter0, gate118inter1, gate118inter2, gate118inter3, gate118inter4, gate118inter5, gate118inter6, gate118inter7, gate118inter8, gate118inter9, gate118inter10, gate118inter11, gate118inter12, gate206inter0, gate206inter1, gate206inter2, gate206inter3, gate206inter4, gate206inter5, gate206inter6, gate206inter7, gate206inter8, gate206inter9, gate206inter10, gate206inter11, gate206inter12, gate240inter0, gate240inter1, gate240inter2, gate240inter3, gate240inter4, gate240inter5, gate240inter6, gate240inter7, gate240inter8, gate240inter9, gate240inter10, gate240inter11, gate240inter12, gate294inter0, gate294inter1, gate294inter2, gate294inter3, gate294inter4, gate294inter5, gate294inter6, gate294inter7, gate294inter8, gate294inter9, gate294inter10, gate294inter11, gate294inter12, gate387inter0, gate387inter1, gate387inter2, gate387inter3, gate387inter4, gate387inter5, gate387inter6, gate387inter7, gate387inter8, gate387inter9, gate387inter10, gate387inter11, gate387inter12, gate431inter0, gate431inter1, gate431inter2, gate431inter3, gate431inter4, gate431inter5, gate431inter6, gate431inter7, gate431inter8, gate431inter9, gate431inter10, gate431inter11, gate431inter12, gate197inter0, gate197inter1, gate197inter2, gate197inter3, gate197inter4, gate197inter5, gate197inter6, gate197inter7, gate197inter8, gate197inter9, gate197inter10, gate197inter11, gate197inter12, gate404inter0, gate404inter1, gate404inter2, gate404inter3, gate404inter4, gate404inter5, gate404inter6, gate404inter7, gate404inter8, gate404inter9, gate404inter10, gate404inter11, gate404inter12, gate410inter0, gate410inter1, gate410inter2, gate410inter3, gate410inter4, gate410inter5, gate410inter6, gate410inter7, gate410inter8, gate410inter9, gate410inter10, gate410inter11, gate410inter12, gate278inter0, gate278inter1, gate278inter2, gate278inter3, gate278inter4, gate278inter5, gate278inter6, gate278inter7, gate278inter8, gate278inter9, gate278inter10, gate278inter11, gate278inter12, gate122inter0, gate122inter1, gate122inter2, gate122inter3, gate122inter4, gate122inter5, gate122inter6, gate122inter7, gate122inter8, gate122inter9, gate122inter10, gate122inter11, gate122inter12, gate256inter0, gate256inter1, gate256inter2, gate256inter3, gate256inter4, gate256inter5, gate256inter6, gate256inter7, gate256inter8, gate256inter9, gate256inter10, gate256inter11, gate256inter12, gate243inter0, gate243inter1, gate243inter2, gate243inter3, gate243inter4, gate243inter5, gate243inter6, gate243inter7, gate243inter8, gate243inter9, gate243inter10, gate243inter11, gate243inter12, gate200inter0, gate200inter1, gate200inter2, gate200inter3, gate200inter4, gate200inter5, gate200inter6, gate200inter7, gate200inter8, gate200inter9, gate200inter10, gate200inter11, gate200inter12, gate18inter0, gate18inter1, gate18inter2, gate18inter3, gate18inter4, gate18inter5, gate18inter6, gate18inter7, gate18inter8, gate18inter9, gate18inter10, gate18inter11, gate18inter12, gate270inter0, gate270inter1, gate270inter2, gate270inter3, gate270inter4, gate270inter5, gate270inter6, gate270inter7, gate270inter8, gate270inter9, gate270inter10, gate270inter11, gate270inter12, gate87inter0, gate87inter1, gate87inter2, gate87inter3, gate87inter4, gate87inter5, gate87inter6, gate87inter7, gate87inter8, gate87inter9, gate87inter10, gate87inter11, gate87inter12, gate389inter0, gate389inter1, gate389inter2, gate389inter3, gate389inter4, gate389inter5, gate389inter6, gate389inter7, gate389inter8, gate389inter9, gate389inter10, gate389inter11, gate389inter12, gate179inter0, gate179inter1, gate179inter2, gate179inter3, gate179inter4, gate179inter5, gate179inter6, gate179inter7, gate179inter8, gate179inter9, gate179inter10, gate179inter11, gate179inter12, gate447inter0, gate447inter1, gate447inter2, gate447inter3, gate447inter4, gate447inter5, gate447inter6, gate447inter7, gate447inter8, gate447inter9, gate447inter10, gate447inter11, gate447inter12, gate154inter0, gate154inter1, gate154inter2, gate154inter3, gate154inter4, gate154inter5, gate154inter6, gate154inter7, gate154inter8, gate154inter9, gate154inter10, gate154inter11, gate154inter12, gate470inter0, gate470inter1, gate470inter2, gate470inter3, gate470inter4, gate470inter5, gate470inter6, gate470inter7, gate470inter8, gate470inter9, gate470inter10, gate470inter11, gate470inter12, gate57inter0, gate57inter1, gate57inter2, gate57inter3, gate57inter4, gate57inter5, gate57inter6, gate57inter7, gate57inter8, gate57inter9, gate57inter10, gate57inter11, gate57inter12, gate98inter0, gate98inter1, gate98inter2, gate98inter3, gate98inter4, gate98inter5, gate98inter6, gate98inter7, gate98inter8, gate98inter9, gate98inter10, gate98inter11, gate98inter12, gate265inter0, gate265inter1, gate265inter2, gate265inter3, gate265inter4, gate265inter5, gate265inter6, gate265inter7, gate265inter8, gate265inter9, gate265inter10, gate265inter11, gate265inter12, gate423inter0, gate423inter1, gate423inter2, gate423inter3, gate423inter4, gate423inter5, gate423inter6, gate423inter7, gate423inter8, gate423inter9, gate423inter10, gate423inter11, gate423inter12, gate491inter0, gate491inter1, gate491inter2, gate491inter3, gate491inter4, gate491inter5, gate491inter6, gate491inter7, gate491inter8, gate491inter9, gate491inter10, gate491inter11, gate491inter12, gate499inter0, gate499inter1, gate499inter2, gate499inter3, gate499inter4, gate499inter5, gate499inter6, gate499inter7, gate499inter8, gate499inter9, gate499inter10, gate499inter11, gate499inter12, gate183inter0, gate183inter1, gate183inter2, gate183inter3, gate183inter4, gate183inter5, gate183inter6, gate183inter7, gate183inter8, gate183inter9, gate183inter10, gate183inter11, gate183inter12, gate290inter0, gate290inter1, gate290inter2, gate290inter3, gate290inter4, gate290inter5, gate290inter6, gate290inter7, gate290inter8, gate290inter9, gate290inter10, gate290inter11, gate290inter12, gate45inter0, gate45inter1, gate45inter2, gate45inter3, gate45inter4, gate45inter5, gate45inter6, gate45inter7, gate45inter8, gate45inter9, gate45inter10, gate45inter11, gate45inter12, gate217inter0, gate217inter1, gate217inter2, gate217inter3, gate217inter4, gate217inter5, gate217inter6, gate217inter7, gate217inter8, gate217inter9, gate217inter10, gate217inter11, gate217inter12, gate492inter0, gate492inter1, gate492inter2, gate492inter3, gate492inter4, gate492inter5, gate492inter6, gate492inter7, gate492inter8, gate492inter9, gate492inter10, gate492inter11, gate492inter12, gate63inter0, gate63inter1, gate63inter2, gate63inter3, gate63inter4, gate63inter5, gate63inter6, gate63inter7, gate63inter8, gate63inter9, gate63inter10, gate63inter11, gate63inter12, gate485inter0, gate485inter1, gate485inter2, gate485inter3, gate485inter4, gate485inter5, gate485inter6, gate485inter7, gate485inter8, gate485inter9, gate485inter10, gate485inter11, gate485inter12, gate125inter0, gate125inter1, gate125inter2, gate125inter3, gate125inter4, gate125inter5, gate125inter6, gate125inter7, gate125inter8, gate125inter9, gate125inter10, gate125inter11, gate125inter12, gate61inter0, gate61inter1, gate61inter2, gate61inter3, gate61inter4, gate61inter5, gate61inter6, gate61inter7, gate61inter8, gate61inter9, gate61inter10, gate61inter11, gate61inter12, gate46inter0, gate46inter1, gate46inter2, gate46inter3, gate46inter4, gate46inter5, gate46inter6, gate46inter7, gate46inter8, gate46inter9, gate46inter10, gate46inter11, gate46inter12, gate453inter0, gate453inter1, gate453inter2, gate453inter3, gate453inter4, gate453inter5, gate453inter6, gate453inter7, gate453inter8, gate453inter9, gate453inter10, gate453inter11, gate453inter12, gate425inter0, gate425inter1, gate425inter2, gate425inter3, gate425inter4, gate425inter5, gate425inter6, gate425inter7, gate425inter8, gate425inter9, gate425inter10, gate425inter11, gate425inter12, gate424inter0, gate424inter1, gate424inter2, gate424inter3, gate424inter4, gate424inter5, gate424inter6, gate424inter7, gate424inter8, gate424inter9, gate424inter10, gate424inter11, gate424inter12, gate148inter0, gate148inter1, gate148inter2, gate148inter3, gate148inter4, gate148inter5, gate148inter6, gate148inter7, gate148inter8, gate148inter9, gate148inter10, gate148inter11, gate148inter12, gate28inter0, gate28inter1, gate28inter2, gate28inter3, gate28inter4, gate28inter5, gate28inter6, gate28inter7, gate28inter8, gate28inter9, gate28inter10, gate28inter11, gate28inter12, gate58inter0, gate58inter1, gate58inter2, gate58inter3, gate58inter4, gate58inter5, gate58inter6, gate58inter7, gate58inter8, gate58inter9, gate58inter10, gate58inter11, gate58inter12, gate443inter0, gate443inter1, gate443inter2, gate443inter3, gate443inter4, gate443inter5, gate443inter6, gate443inter7, gate443inter8, gate443inter9, gate443inter10, gate443inter11, gate443inter12, gate428inter0, gate428inter1, gate428inter2, gate428inter3, gate428inter4, gate428inter5, gate428inter6, gate428inter7, gate428inter8, gate428inter9, gate428inter10, gate428inter11, gate428inter12, gate25inter0, gate25inter1, gate25inter2, gate25inter3, gate25inter4, gate25inter5, gate25inter6, gate25inter7, gate25inter8, gate25inter9, gate25inter10, gate25inter11, gate25inter12, gate142inter0, gate142inter1, gate142inter2, gate142inter3, gate142inter4, gate142inter5, gate142inter6, gate142inter7, gate142inter8, gate142inter9, gate142inter10, gate142inter11, gate142inter12, gate466inter0, gate466inter1, gate466inter2, gate466inter3, gate466inter4, gate466inter5, gate466inter6, gate466inter7, gate466inter8, gate466inter9, gate466inter10, gate466inter11, gate466inter12, gate14inter0, gate14inter1, gate14inter2, gate14inter3, gate14inter4, gate14inter5, gate14inter6, gate14inter7, gate14inter8, gate14inter9, gate14inter10, gate14inter11, gate14inter12, gate249inter0, gate249inter1, gate249inter2, gate249inter3, gate249inter4, gate249inter5, gate249inter6, gate249inter7, gate249inter8, gate249inter9, gate249inter10, gate249inter11, gate249inter12, gate107inter0, gate107inter1, gate107inter2, gate107inter3, gate107inter4, gate107inter5, gate107inter6, gate107inter7, gate107inter8, gate107inter9, gate107inter10, gate107inter11, gate107inter12, gate108inter0, gate108inter1, gate108inter2, gate108inter3, gate108inter4, gate108inter5, gate108inter6, gate108inter7, gate108inter8, gate108inter9, gate108inter10, gate108inter11, gate108inter12, gate152inter0, gate152inter1, gate152inter2, gate152inter3, gate152inter4, gate152inter5, gate152inter6, gate152inter7, gate152inter8, gate152inter9, gate152inter10, gate152inter11, gate152inter12, gate109inter0, gate109inter1, gate109inter2, gate109inter3, gate109inter4, gate109inter5, gate109inter6, gate109inter7, gate109inter8, gate109inter9, gate109inter10, gate109inter11, gate109inter12, gate459inter0, gate459inter1, gate459inter2, gate459inter3, gate459inter4, gate459inter5, gate459inter6, gate459inter7, gate459inter8, gate459inter9, gate459inter10, gate459inter11, gate459inter12, gate70inter0, gate70inter1, gate70inter2, gate70inter3, gate70inter4, gate70inter5, gate70inter6, gate70inter7, gate70inter8, gate70inter9, gate70inter10, gate70inter11, gate70inter12, gate69inter0, gate69inter1, gate69inter2, gate69inter3, gate69inter4, gate69inter5, gate69inter6, gate69inter7, gate69inter8, gate69inter9, gate69inter10, gate69inter11, gate69inter12, gate31inter0, gate31inter1, gate31inter2, gate31inter3, gate31inter4, gate31inter5, gate31inter6, gate31inter7, gate31inter8, gate31inter9, gate31inter10, gate31inter11, gate31inter12, gate286inter0, gate286inter1, gate286inter2, gate286inter3, gate286inter4, gate286inter5, gate286inter6, gate286inter7, gate286inter8, gate286inter9, gate286inter10, gate286inter11, gate286inter12, gate244inter0, gate244inter1, gate244inter2, gate244inter3, gate244inter4, gate244inter5, gate244inter6, gate244inter7, gate244inter8, gate244inter9, gate244inter10, gate244inter11, gate244inter12, gate40inter0, gate40inter1, gate40inter2, gate40inter3, gate40inter4, gate40inter5, gate40inter6, gate40inter7, gate40inter8, gate40inter9, gate40inter10, gate40inter11, gate40inter12, gate38inter0, gate38inter1, gate38inter2, gate38inter3, gate38inter4, gate38inter5, gate38inter6, gate38inter7, gate38inter8, gate38inter9, gate38inter10, gate38inter11, gate38inter12, gate245inter0, gate245inter1, gate245inter2, gate245inter3, gate245inter4, gate245inter5, gate245inter6, gate245inter7, gate245inter8, gate245inter9, gate245inter10, gate245inter11, gate245inter12, gate433inter0, gate433inter1, gate433inter2, gate433inter3, gate433inter4, gate433inter5, gate433inter6, gate433inter7, gate433inter8, gate433inter9, gate433inter10, gate433inter11, gate433inter12, gate201inter0, gate201inter1, gate201inter2, gate201inter3, gate201inter4, gate201inter5, gate201inter6, gate201inter7, gate201inter8, gate201inter9, gate201inter10, gate201inter11, gate201inter12, gate236inter0, gate236inter1, gate236inter2, gate236inter3, gate236inter4, gate236inter5, gate236inter6, gate236inter7, gate236inter8, gate236inter9, gate236inter10, gate236inter11, gate236inter12, gate232inter0, gate232inter1, gate232inter2, gate232inter3, gate232inter4, gate232inter5, gate232inter6, gate232inter7, gate232inter8, gate232inter9, gate232inter10, gate232inter11, gate232inter12, gate113inter0, gate113inter1, gate113inter2, gate113inter3, gate113inter4, gate113inter5, gate113inter6, gate113inter7, gate113inter8, gate113inter9, gate113inter10, gate113inter11, gate113inter12, gate274inter0, gate274inter1, gate274inter2, gate274inter3, gate274inter4, gate274inter5, gate274inter6, gate274inter7, gate274inter8, gate274inter9, gate274inter10, gate274inter11, gate274inter12, gate262inter0, gate262inter1, gate262inter2, gate262inter3, gate262inter4, gate262inter5, gate262inter6, gate262inter7, gate262inter8, gate262inter9, gate262inter10, gate262inter11, gate262inter12, gate85inter0, gate85inter1, gate85inter2, gate85inter3, gate85inter4, gate85inter5, gate85inter6, gate85inter7, gate85inter8, gate85inter9, gate85inter10, gate85inter11, gate85inter12, gate196inter0, gate196inter1, gate196inter2, gate196inter3, gate196inter4, gate196inter5, gate196inter6, gate196inter7, gate196inter8, gate196inter9, gate196inter10, gate196inter11, gate196inter12, gate494inter0, gate494inter1, gate494inter2, gate494inter3, gate494inter4, gate494inter5, gate494inter6, gate494inter7, gate494inter8, gate494inter9, gate494inter10, gate494inter11, gate494inter12, gate507inter0, gate507inter1, gate507inter2, gate507inter3, gate507inter4, gate507inter5, gate507inter6, gate507inter7, gate507inter8, gate507inter9, gate507inter10, gate507inter11, gate507inter12, gate44inter0, gate44inter1, gate44inter2, gate44inter3, gate44inter4, gate44inter5, gate44inter6, gate44inter7, gate44inter8, gate44inter9, gate44inter10, gate44inter11, gate44inter12, gate504inter0, gate504inter1, gate504inter2, gate504inter3, gate504inter4, gate504inter5, gate504inter6, gate504inter7, gate504inter8, gate504inter9, gate504inter10, gate504inter11, gate504inter12, gate426inter0, gate426inter1, gate426inter2, gate426inter3, gate426inter4, gate426inter5, gate426inter6, gate426inter7, gate426inter8, gate426inter9, gate426inter10, gate426inter11, gate426inter12, gate29inter0, gate29inter1, gate29inter2, gate29inter3, gate29inter4, gate29inter5, gate29inter6, gate29inter7, gate29inter8, gate29inter9, gate29inter10, gate29inter11, gate29inter12, gate170inter0, gate170inter1, gate170inter2, gate170inter3, gate170inter4, gate170inter5, gate170inter6, gate170inter7, gate170inter8, gate170inter9, gate170inter10, gate170inter11, gate170inter12, gate138inter0, gate138inter1, gate138inter2, gate138inter3, gate138inter4, gate138inter5, gate138inter6, gate138inter7, gate138inter8, gate138inter9, gate138inter10, gate138inter11, gate138inter12, gate511inter0, gate511inter1, gate511inter2, gate511inter3, gate511inter4, gate511inter5, gate511inter6, gate511inter7, gate511inter8, gate511inter9, gate511inter10, gate511inter11, gate511inter12, gate411inter0, gate411inter1, gate411inter2, gate411inter3, gate411inter4, gate411inter5, gate411inter6, gate411inter7, gate411inter8, gate411inter9, gate411inter10, gate411inter11, gate411inter12, gate413inter0, gate413inter1, gate413inter2, gate413inter3, gate413inter4, gate413inter5, gate413inter6, gate413inter7, gate413inter8, gate413inter9, gate413inter10, gate413inter11, gate413inter12, gate288inter0, gate288inter1, gate288inter2, gate288inter3, gate288inter4, gate288inter5, gate288inter6, gate288inter7, gate288inter8, gate288inter9, gate288inter10, gate288inter11, gate288inter12, gate41inter0, gate41inter1, gate41inter2, gate41inter3, gate41inter4, gate41inter5, gate41inter6, gate41inter7, gate41inter8, gate41inter9, gate41inter10, gate41inter11, gate41inter12, gate400inter0, gate400inter1, gate400inter2, gate400inter3, gate400inter4, gate400inter5, gate400inter6, gate400inter7, gate400inter8, gate400inter9, gate400inter10, gate400inter11, gate400inter12, gate130inter0, gate130inter1, gate130inter2, gate130inter3, gate130inter4, gate130inter5, gate130inter6, gate130inter7, gate130inter8, gate130inter9, gate130inter10, gate130inter11, gate130inter12, gate15inter0, gate15inter1, gate15inter2, gate15inter3, gate15inter4, gate15inter5, gate15inter6, gate15inter7, gate15inter8, gate15inter9, gate15inter10, gate15inter11, gate15inter12, gate226inter0, gate226inter1, gate226inter2, gate226inter3, gate226inter4, gate226inter5, gate226inter6, gate226inter7, gate226inter8, gate226inter9, gate226inter10, gate226inter11, gate226inter12, gate505inter0, gate505inter1, gate505inter2, gate505inter3, gate505inter4, gate505inter5, gate505inter6, gate505inter7, gate505inter8, gate505inter9, gate505inter10, gate505inter11, gate505inter12, gate47inter0, gate47inter1, gate47inter2, gate47inter3, gate47inter4, gate47inter5, gate47inter6, gate47inter7, gate47inter8, gate47inter9, gate47inter10, gate47inter11, gate47inter12, gate95inter0, gate95inter1, gate95inter2, gate95inter3, gate95inter4, gate95inter5, gate95inter6, gate95inter7, gate95inter8, gate95inter9, gate95inter10, gate95inter11, gate95inter12, gate156inter0, gate156inter1, gate156inter2, gate156inter3, gate156inter4, gate156inter5, gate156inter6, gate156inter7, gate156inter8, gate156inter9, gate156inter10, gate156inter11, gate156inter12, gate146inter0, gate146inter1, gate146inter2, gate146inter3, gate146inter4, gate146inter5, gate146inter6, gate146inter7, gate146inter8, gate146inter9, gate146inter10, gate146inter11, gate146inter12, gate43inter0, gate43inter1, gate43inter2, gate43inter3, gate43inter4, gate43inter5, gate43inter6, gate43inter7, gate43inter8, gate43inter9, gate43inter10, gate43inter11, gate43inter12, gate394inter0, gate394inter1, gate394inter2, gate394inter3, gate394inter4, gate394inter5, gate394inter6, gate394inter7, gate394inter8, gate394inter9, gate394inter10, gate394inter11, gate394inter12, gate225inter0, gate225inter1, gate225inter2, gate225inter3, gate225inter4, gate225inter5, gate225inter6, gate225inter7, gate225inter8, gate225inter9, gate225inter10, gate225inter11, gate225inter12, gate66inter0, gate66inter1, gate66inter2, gate66inter3, gate66inter4, gate66inter5, gate66inter6, gate66inter7, gate66inter8, gate66inter9, gate66inter10, gate66inter11, gate66inter12, gate502inter0, gate502inter1, gate502inter2, gate502inter3, gate502inter4, gate502inter5, gate502inter6, gate502inter7, gate502inter8, gate502inter9, gate502inter10, gate502inter11, gate502inter12, gate62inter0, gate62inter1, gate62inter2, gate62inter3, gate62inter4, gate62inter5, gate62inter6, gate62inter7, gate62inter8, gate62inter9, gate62inter10, gate62inter11, gate62inter12, gate214inter0, gate214inter1, gate214inter2, gate214inter3, gate214inter4, gate214inter5, gate214inter6, gate214inter7, gate214inter8, gate214inter9, gate214inter10, gate214inter11, gate214inter12, gate149inter0, gate149inter1, gate149inter2, gate149inter3, gate149inter4, gate149inter5, gate149inter6, gate149inter7, gate149inter8, gate149inter9, gate149inter10, gate149inter11, gate149inter12, gate72inter0, gate72inter1, gate72inter2, gate72inter3, gate72inter4, gate72inter5, gate72inter6, gate72inter7, gate72inter8, gate72inter9, gate72inter10, gate72inter11, gate72inter12, gate405inter0, gate405inter1, gate405inter2, gate405inter3, gate405inter4, gate405inter5, gate405inter6, gate405inter7, gate405inter8, gate405inter9, gate405inter10, gate405inter11, gate405inter12, gate477inter0, gate477inter1, gate477inter2, gate477inter3, gate477inter4, gate477inter5, gate477inter6, gate477inter7, gate477inter8, gate477inter9, gate477inter10, gate477inter11, gate477inter12, gate289inter0, gate289inter1, gate289inter2, gate289inter3, gate289inter4, gate289inter5, gate289inter6, gate289inter7, gate289inter8, gate289inter9, gate289inter10, gate289inter11, gate289inter12, gate187inter0, gate187inter1, gate187inter2, gate187inter3, gate187inter4, gate187inter5, gate187inter6, gate187inter7, gate187inter8, gate187inter9, gate187inter10, gate187inter11, gate187inter12, gate17inter0, gate17inter1, gate17inter2, gate17inter3, gate17inter4, gate17inter5, gate17inter6, gate17inter7, gate17inter8, gate17inter9, gate17inter10, gate17inter11, gate17inter12, gate90inter0, gate90inter1, gate90inter2, gate90inter3, gate90inter4, gate90inter5, gate90inter6, gate90inter7, gate90inter8, gate90inter9, gate90inter10, gate90inter11, gate90inter12, gate71inter0, gate71inter1, gate71inter2, gate71inter3, gate71inter4, gate71inter5, gate71inter6, gate71inter7, gate71inter8, gate71inter9, gate71inter10, gate71inter11, gate71inter12, gate415inter0, gate415inter1, gate415inter2, gate415inter3, gate415inter4, gate415inter5, gate415inter6, gate415inter7, gate415inter8, gate415inter9, gate415inter10, gate415inter11, gate415inter12, gate417inter0, gate417inter1, gate417inter2, gate417inter3, gate417inter4, gate417inter5, gate417inter6, gate417inter7, gate417inter8, gate417inter9, gate417inter10, gate417inter11, gate417inter12, gate119inter0, gate119inter1, gate119inter2, gate119inter3, gate119inter4, gate119inter5, gate119inter6, gate119inter7, gate119inter8, gate119inter9, gate119inter10, gate119inter11, gate119inter12, gate250inter0, gate250inter1, gate250inter2, gate250inter3, gate250inter4, gate250inter5, gate250inter6, gate250inter7, gate250inter8, gate250inter9, gate250inter10, gate250inter11, gate250inter12, gate10inter0, gate10inter1, gate10inter2, gate10inter3, gate10inter4, gate10inter5, gate10inter6, gate10inter7, gate10inter8, gate10inter9, gate10inter10, gate10inter11, gate10inter12, gate101inter0, gate101inter1, gate101inter2, gate101inter3, gate101inter4, gate101inter5, gate101inter6, gate101inter7, gate101inter8, gate101inter9, gate101inter10, gate101inter11, gate101inter12, gate407inter0, gate407inter1, gate407inter2, gate407inter3, gate407inter4, gate407inter5, gate407inter6, gate407inter7, gate407inter8, gate407inter9, gate407inter10, gate407inter11, gate407inter12, gate175inter0, gate175inter1, gate175inter2, gate175inter3, gate175inter4, gate175inter5, gate175inter6, gate175inter7, gate175inter8, gate175inter9, gate175inter10, gate175inter11, gate175inter12, gate280inter0, gate280inter1, gate280inter2, gate280inter3, gate280inter4, gate280inter5, gate280inter6, gate280inter7, gate280inter8, gate280inter9, gate280inter10, gate280inter11, gate280inter12, gate512inter0, gate512inter1, gate512inter2, gate512inter3, gate512inter4, gate512inter5, gate512inter6, gate512inter7, gate512inter8, gate512inter9, gate512inter10, gate512inter11, gate512inter12, gate213inter0, gate213inter1, gate213inter2, gate213inter3, gate213inter4, gate213inter5, gate213inter6, gate213inter7, gate213inter8, gate213inter9, gate213inter10, gate213inter11, gate213inter12, gate460inter0, gate460inter1, gate460inter2, gate460inter3, gate460inter4, gate460inter5, gate460inter6, gate460inter7, gate460inter8, gate460inter9, gate460inter10, gate460inter11, gate460inter12, gate195inter0, gate195inter1, gate195inter2, gate195inter3, gate195inter4, gate195inter5, gate195inter6, gate195inter7, gate195inter8, gate195inter9, gate195inter10, gate195inter11, gate195inter12, gate449inter0, gate449inter1, gate449inter2, gate449inter3, gate449inter4, gate449inter5, gate449inter6, gate449inter7, gate449inter8, gate449inter9, gate449inter10, gate449inter11, gate449inter12, gate478inter0, gate478inter1, gate478inter2, gate478inter3, gate478inter4, gate478inter5, gate478inter6, gate478inter7, gate478inter8, gate478inter9, gate478inter10, gate478inter11, gate478inter12, gate114inter0, gate114inter1, gate114inter2, gate114inter3, gate114inter4, gate114inter5, gate114inter6, gate114inter7, gate114inter8, gate114inter9, gate114inter10, gate114inter11, gate114inter12, gate78inter0, gate78inter1, gate78inter2, gate78inter3, gate78inter4, gate78inter5, gate78inter6, gate78inter7, gate78inter8, gate78inter9, gate78inter10, gate78inter11, gate78inter12, gate64inter0, gate64inter1, gate64inter2, gate64inter3, gate64inter4, gate64inter5, gate64inter6, gate64inter7, gate64inter8, gate64inter9, gate64inter10, gate64inter11, gate64inter12, gate79inter0, gate79inter1, gate79inter2, gate79inter3, gate79inter4, gate79inter5, gate79inter6, gate79inter7, gate79inter8, gate79inter9, gate79inter10, gate79inter11, gate79inter12, gate399inter0, gate399inter1, gate399inter2, gate399inter3, gate399inter4, gate399inter5, gate399inter6, gate399inter7, gate399inter8, gate399inter9, gate399inter10, gate399inter11, gate399inter12, gate180inter0, gate180inter1, gate180inter2, gate180inter3, gate180inter4, gate180inter5, gate180inter6, gate180inter7, gate180inter8, gate180inter9, gate180inter10, gate180inter11, gate180inter12, gate414inter0, gate414inter1, gate414inter2, gate414inter3, gate414inter4, gate414inter5, gate414inter6, gate414inter7, gate414inter8, gate414inter9, gate414inter10, gate414inter11, gate414inter12, gate242inter0, gate242inter1, gate242inter2, gate242inter3, gate242inter4, gate242inter5, gate242inter6, gate242inter7, gate242inter8, gate242inter9, gate242inter10, gate242inter11, gate242inter12, gate194inter0, gate194inter1, gate194inter2, gate194inter3, gate194inter4, gate194inter5, gate194inter6, gate194inter7, gate194inter8, gate194inter9, gate194inter10, gate194inter11, gate194inter12, gate448inter0, gate448inter1, gate448inter2, gate448inter3, gate448inter4, gate448inter5, gate448inter6, gate448inter7, gate448inter8, gate448inter9, gate448inter10, gate448inter11, gate448inter12, gate139inter0, gate139inter1, gate139inter2, gate139inter3, gate139inter4, gate139inter5, gate139inter6, gate139inter7, gate139inter8, gate139inter9, gate139inter10, gate139inter11, gate139inter12, gate497inter0, gate497inter1, gate497inter2, gate497inter3, gate497inter4, gate497inter5, gate497inter6, gate497inter7, gate497inter8, gate497inter9, gate497inter10, gate497inter11, gate497inter12, gate48inter0, gate48inter1, gate48inter2, gate48inter3, gate48inter4, gate48inter5, gate48inter6, gate48inter7, gate48inter8, gate48inter9, gate48inter10, gate48inter11, gate48inter12, gate84inter0, gate84inter1, gate84inter2, gate84inter3, gate84inter4, gate84inter5, gate84inter6, gate84inter7, gate84inter8, gate84inter9, gate84inter10, gate84inter11, gate84inter12, gate277inter0, gate277inter1, gate277inter2, gate277inter3, gate277inter4, gate277inter5, gate277inter6, gate277inter7, gate277inter8, gate277inter9, gate277inter10, gate277inter11, gate277inter12, gate178inter0, gate178inter1, gate178inter2, gate178inter3, gate178inter4, gate178inter5, gate178inter6, gate178inter7, gate178inter8, gate178inter9, gate178inter10, gate178inter11, gate178inter12, gate76inter0, gate76inter1, gate76inter2, gate76inter3, gate76inter4, gate76inter5, gate76inter6, gate76inter7, gate76inter8, gate76inter9, gate76inter10, gate76inter11, gate76inter12, gate49inter0, gate49inter1, gate49inter2, gate49inter3, gate49inter4, gate49inter5, gate49inter6, gate49inter7, gate49inter8, gate49inter9, gate49inter10, gate49inter11, gate49inter12, gate30inter0, gate30inter1, gate30inter2, gate30inter3, gate30inter4, gate30inter5, gate30inter6, gate30inter7, gate30inter8, gate30inter9, gate30inter10, gate30inter11, gate30inter12, gate412inter0, gate412inter1, gate412inter2, gate412inter3, gate412inter4, gate412inter5, gate412inter6, gate412inter7, gate412inter8, gate412inter9, gate412inter10, gate412inter11, gate412inter12, gate285inter0, gate285inter1, gate285inter2, gate285inter3, gate285inter4, gate285inter5, gate285inter6, gate285inter7, gate285inter8, gate285inter9, gate285inter10, gate285inter11, gate285inter12, gate205inter0, gate205inter1, gate205inter2, gate205inter3, gate205inter4, gate205inter5, gate205inter6, gate205inter7, gate205inter8, gate205inter9, gate205inter10, gate205inter11, gate205inter12, gate422inter0, gate422inter1, gate422inter2, gate422inter3, gate422inter4, gate422inter5, gate422inter6, gate422inter7, gate422inter8, gate422inter9, gate422inter10, gate422inter11, gate422inter12, gate402inter0, gate402inter1, gate402inter2, gate402inter3, gate402inter4, gate402inter5, gate402inter6, gate402inter7, gate402inter8, gate402inter9, gate402inter10, gate402inter11, gate402inter12, gate287inter0, gate287inter1, gate287inter2, gate287inter3, gate287inter4, gate287inter5, gate287inter6, gate287inter7, gate287inter8, gate287inter9, gate287inter10, gate287inter11, gate287inter12, gate388inter0, gate388inter1, gate388inter2, gate388inter3, gate388inter4, gate388inter5, gate388inter6, gate388inter7, gate388inter8, gate388inter9, gate388inter10, gate388inter11, gate388inter12, gate258inter0, gate258inter1, gate258inter2, gate258inter3, gate258inter4, gate258inter5, gate258inter6, gate258inter7, gate258inter8, gate258inter9, gate258inter10, gate258inter11, gate258inter12, gate230inter0, gate230inter1, gate230inter2, gate230inter3, gate230inter4, gate230inter5, gate230inter6, gate230inter7, gate230inter8, gate230inter9, gate230inter10, gate230inter11, gate230inter12, gate34inter0, gate34inter1, gate34inter2, gate34inter3, gate34inter4, gate34inter5, gate34inter6, gate34inter7, gate34inter8, gate34inter9, gate34inter10, gate34inter11, gate34inter12, gate192inter0, gate192inter1, gate192inter2, gate192inter3, gate192inter4, gate192inter5, gate192inter6, gate192inter7, gate192inter8, gate192inter9, gate192inter10, gate192inter11, gate192inter12, gate233inter0, gate233inter1, gate233inter2, gate233inter3, gate233inter4, gate233inter5, gate233inter6, gate233inter7, gate233inter8, gate233inter9, gate233inter10, gate233inter11, gate233inter12, gate181inter0, gate181inter1, gate181inter2, gate181inter3, gate181inter4, gate181inter5, gate181inter6, gate181inter7, gate181inter8, gate181inter9, gate181inter10, gate181inter11, gate181inter12, gate54inter0, gate54inter1, gate54inter2, gate54inter3, gate54inter4, gate54inter5, gate54inter6, gate54inter7, gate54inter8, gate54inter9, gate54inter10, gate54inter11, gate54inter12, gate52inter0, gate52inter1, gate52inter2, gate52inter3, gate52inter4, gate52inter5, gate52inter6, gate52inter7, gate52inter8, gate52inter9, gate52inter10, gate52inter11, gate52inter12, gate416inter0, gate416inter1, gate416inter2, gate416inter3, gate416inter4, gate416inter5, gate416inter6, gate416inter7, gate416inter8, gate416inter9, gate416inter10, gate416inter11, gate416inter12, gate462inter0, gate462inter1, gate462inter2, gate462inter3, gate462inter4, gate462inter5, gate462inter6, gate462inter7, gate462inter8, gate462inter9, gate462inter10, gate462inter11, gate462inter12, gate498inter0, gate498inter1, gate498inter2, gate498inter3, gate498inter4, gate498inter5, gate498inter6, gate498inter7, gate498inter8, gate498inter9, gate498inter10, gate498inter11, gate498inter12, gate190inter0, gate190inter1, gate190inter2, gate190inter3, gate190inter4, gate190inter5, gate190inter6, gate190inter7, gate190inter8, gate190inter9, gate190inter10, gate190inter11, gate190inter12, gate508inter0, gate508inter1, gate508inter2, gate508inter3, gate508inter4, gate508inter5, gate508inter6, gate508inter7, gate508inter8, gate508inter9, gate508inter10, gate508inter11, gate508inter12, gate169inter0, gate169inter1, gate169inter2, gate169inter3, gate169inter4, gate169inter5, gate169inter6, gate169inter7, gate169inter8, gate169inter9, gate169inter10, gate169inter11, gate169inter12, gate220inter0, gate220inter1, gate220inter2, gate220inter3, gate220inter4, gate220inter5, gate220inter6, gate220inter7, gate220inter8, gate220inter9, gate220inter10, gate220inter11, gate220inter12, gate161inter0, gate161inter1, gate161inter2, gate161inter3, gate161inter4, gate161inter5, gate161inter6, gate161inter7, gate161inter8, gate161inter9, gate161inter10, gate161inter11, gate161inter12;



and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );
nand2 gate9( .a(G1), .b(G2), .O(G266) );

  xor2  gate2409(.a(G4), .b(G3), .O(gate10inter0));
  nand2 gate2410(.a(gate10inter0), .b(s_266), .O(gate10inter1));
  and2  gate2411(.a(G4), .b(G3), .O(gate10inter2));
  inv1  gate2412(.a(s_266), .O(gate10inter3));
  inv1  gate2413(.a(s_267), .O(gate10inter4));
  nand2 gate2414(.a(gate10inter4), .b(gate10inter3), .O(gate10inter5));
  nor2  gate2415(.a(gate10inter5), .b(gate10inter2), .O(gate10inter6));
  inv1  gate2416(.a(G3), .O(gate10inter7));
  inv1  gate2417(.a(G4), .O(gate10inter8));
  nand2 gate2418(.a(gate10inter8), .b(gate10inter7), .O(gate10inter9));
  nand2 gate2419(.a(s_267), .b(gate10inter3), .O(gate10inter10));
  nor2  gate2420(.a(gate10inter10), .b(gate10inter9), .O(gate10inter11));
  nor2  gate2421(.a(gate10inter11), .b(gate10inter6), .O(gate10inter12));
  nand2 gate2422(.a(gate10inter12), .b(gate10inter1), .O(G269));
nand2 gate11( .a(G5), .b(G6), .O(G272) );
nand2 gate12( .a(G7), .b(G8), .O(G275) );
nand2 gate13( .a(G9), .b(G10), .O(G278) );

  xor2  gate1485(.a(G12), .b(G11), .O(gate14inter0));
  nand2 gate1486(.a(gate14inter0), .b(s_134), .O(gate14inter1));
  and2  gate1487(.a(G12), .b(G11), .O(gate14inter2));
  inv1  gate1488(.a(s_134), .O(gate14inter3));
  inv1  gate1489(.a(s_135), .O(gate14inter4));
  nand2 gate1490(.a(gate14inter4), .b(gate14inter3), .O(gate14inter5));
  nor2  gate1491(.a(gate14inter5), .b(gate14inter2), .O(gate14inter6));
  inv1  gate1492(.a(G11), .O(gate14inter7));
  inv1  gate1493(.a(G12), .O(gate14inter8));
  nand2 gate1494(.a(gate14inter8), .b(gate14inter7), .O(gate14inter9));
  nand2 gate1495(.a(s_135), .b(gate14inter3), .O(gate14inter10));
  nor2  gate1496(.a(gate14inter10), .b(gate14inter9), .O(gate14inter11));
  nor2  gate1497(.a(gate14inter11), .b(gate14inter6), .O(gate14inter12));
  nand2 gate1498(.a(gate14inter12), .b(gate14inter1), .O(G281));

  xor2  gate2031(.a(G14), .b(G13), .O(gate15inter0));
  nand2 gate2032(.a(gate15inter0), .b(s_212), .O(gate15inter1));
  and2  gate2033(.a(G14), .b(G13), .O(gate15inter2));
  inv1  gate2034(.a(s_212), .O(gate15inter3));
  inv1  gate2035(.a(s_213), .O(gate15inter4));
  nand2 gate2036(.a(gate15inter4), .b(gate15inter3), .O(gate15inter5));
  nor2  gate2037(.a(gate15inter5), .b(gate15inter2), .O(gate15inter6));
  inv1  gate2038(.a(G13), .O(gate15inter7));
  inv1  gate2039(.a(G14), .O(gate15inter8));
  nand2 gate2040(.a(gate15inter8), .b(gate15inter7), .O(gate15inter9));
  nand2 gate2041(.a(s_213), .b(gate15inter3), .O(gate15inter10));
  nor2  gate2042(.a(gate15inter10), .b(gate15inter9), .O(gate15inter11));
  nor2  gate2043(.a(gate15inter11), .b(gate15inter6), .O(gate15inter12));
  nand2 gate2044(.a(gate15inter12), .b(gate15inter1), .O(G284));
nand2 gate16( .a(G15), .b(G16), .O(G287) );

  xor2  gate2311(.a(G18), .b(G17), .O(gate17inter0));
  nand2 gate2312(.a(gate17inter0), .b(s_252), .O(gate17inter1));
  and2  gate2313(.a(G18), .b(G17), .O(gate17inter2));
  inv1  gate2314(.a(s_252), .O(gate17inter3));
  inv1  gate2315(.a(s_253), .O(gate17inter4));
  nand2 gate2316(.a(gate17inter4), .b(gate17inter3), .O(gate17inter5));
  nor2  gate2317(.a(gate17inter5), .b(gate17inter2), .O(gate17inter6));
  inv1  gate2318(.a(G17), .O(gate17inter7));
  inv1  gate2319(.a(G18), .O(gate17inter8));
  nand2 gate2320(.a(gate17inter8), .b(gate17inter7), .O(gate17inter9));
  nand2 gate2321(.a(s_253), .b(gate17inter3), .O(gate17inter10));
  nor2  gate2322(.a(gate17inter10), .b(gate17inter9), .O(gate17inter11));
  nor2  gate2323(.a(gate17inter11), .b(gate17inter6), .O(gate17inter12));
  nand2 gate2324(.a(gate17inter12), .b(gate17inter1), .O(G290));

  xor2  gate995(.a(G20), .b(G19), .O(gate18inter0));
  nand2 gate996(.a(gate18inter0), .b(s_64), .O(gate18inter1));
  and2  gate997(.a(G20), .b(G19), .O(gate18inter2));
  inv1  gate998(.a(s_64), .O(gate18inter3));
  inv1  gate999(.a(s_65), .O(gate18inter4));
  nand2 gate1000(.a(gate18inter4), .b(gate18inter3), .O(gate18inter5));
  nor2  gate1001(.a(gate18inter5), .b(gate18inter2), .O(gate18inter6));
  inv1  gate1002(.a(G19), .O(gate18inter7));
  inv1  gate1003(.a(G20), .O(gate18inter8));
  nand2 gate1004(.a(gate18inter8), .b(gate18inter7), .O(gate18inter9));
  nand2 gate1005(.a(s_65), .b(gate18inter3), .O(gate18inter10));
  nor2  gate1006(.a(gate18inter10), .b(gate18inter9), .O(gate18inter11));
  nor2  gate1007(.a(gate18inter11), .b(gate18inter6), .O(gate18inter12));
  nand2 gate1008(.a(gate18inter12), .b(gate18inter1), .O(G293));

  xor2  gate631(.a(G22), .b(G21), .O(gate19inter0));
  nand2 gate632(.a(gate19inter0), .b(s_12), .O(gate19inter1));
  and2  gate633(.a(G22), .b(G21), .O(gate19inter2));
  inv1  gate634(.a(s_12), .O(gate19inter3));
  inv1  gate635(.a(s_13), .O(gate19inter4));
  nand2 gate636(.a(gate19inter4), .b(gate19inter3), .O(gate19inter5));
  nor2  gate637(.a(gate19inter5), .b(gate19inter2), .O(gate19inter6));
  inv1  gate638(.a(G21), .O(gate19inter7));
  inv1  gate639(.a(G22), .O(gate19inter8));
  nand2 gate640(.a(gate19inter8), .b(gate19inter7), .O(gate19inter9));
  nand2 gate641(.a(s_13), .b(gate19inter3), .O(gate19inter10));
  nor2  gate642(.a(gate19inter10), .b(gate19inter9), .O(gate19inter11));
  nor2  gate643(.a(gate19inter11), .b(gate19inter6), .O(gate19inter12));
  nand2 gate644(.a(gate19inter12), .b(gate19inter1), .O(G296));
nand2 gate20( .a(G23), .b(G24), .O(G299) );

  xor2  gate757(.a(G26), .b(G25), .O(gate21inter0));
  nand2 gate758(.a(gate21inter0), .b(s_30), .O(gate21inter1));
  and2  gate759(.a(G26), .b(G25), .O(gate21inter2));
  inv1  gate760(.a(s_30), .O(gate21inter3));
  inv1  gate761(.a(s_31), .O(gate21inter4));
  nand2 gate762(.a(gate21inter4), .b(gate21inter3), .O(gate21inter5));
  nor2  gate763(.a(gate21inter5), .b(gate21inter2), .O(gate21inter6));
  inv1  gate764(.a(G25), .O(gate21inter7));
  inv1  gate765(.a(G26), .O(gate21inter8));
  nand2 gate766(.a(gate21inter8), .b(gate21inter7), .O(gate21inter9));
  nand2 gate767(.a(s_31), .b(gate21inter3), .O(gate21inter10));
  nor2  gate768(.a(gate21inter10), .b(gate21inter9), .O(gate21inter11));
  nor2  gate769(.a(gate21inter11), .b(gate21inter6), .O(gate21inter12));
  nand2 gate770(.a(gate21inter12), .b(gate21inter1), .O(G302));
nand2 gate22( .a(G27), .b(G28), .O(G305) );
nand2 gate23( .a(G29), .b(G30), .O(G308) );
nand2 gate24( .a(G31), .b(G32), .O(G311) );

  xor2  gate1443(.a(G5), .b(G1), .O(gate25inter0));
  nand2 gate1444(.a(gate25inter0), .b(s_128), .O(gate25inter1));
  and2  gate1445(.a(G5), .b(G1), .O(gate25inter2));
  inv1  gate1446(.a(s_128), .O(gate25inter3));
  inv1  gate1447(.a(s_129), .O(gate25inter4));
  nand2 gate1448(.a(gate25inter4), .b(gate25inter3), .O(gate25inter5));
  nor2  gate1449(.a(gate25inter5), .b(gate25inter2), .O(gate25inter6));
  inv1  gate1450(.a(G1), .O(gate25inter7));
  inv1  gate1451(.a(G5), .O(gate25inter8));
  nand2 gate1452(.a(gate25inter8), .b(gate25inter7), .O(gate25inter9));
  nand2 gate1453(.a(s_129), .b(gate25inter3), .O(gate25inter10));
  nor2  gate1454(.a(gate25inter10), .b(gate25inter9), .O(gate25inter11));
  nor2  gate1455(.a(gate25inter11), .b(gate25inter6), .O(gate25inter12));
  nand2 gate1456(.a(gate25inter12), .b(gate25inter1), .O(G314));
nand2 gate26( .a(G9), .b(G13), .O(G317) );
nand2 gate27( .a(G2), .b(G6), .O(G320) );

  xor2  gate1387(.a(G14), .b(G10), .O(gate28inter0));
  nand2 gate1388(.a(gate28inter0), .b(s_120), .O(gate28inter1));
  and2  gate1389(.a(G14), .b(G10), .O(gate28inter2));
  inv1  gate1390(.a(s_120), .O(gate28inter3));
  inv1  gate1391(.a(s_121), .O(gate28inter4));
  nand2 gate1392(.a(gate28inter4), .b(gate28inter3), .O(gate28inter5));
  nor2  gate1393(.a(gate28inter5), .b(gate28inter2), .O(gate28inter6));
  inv1  gate1394(.a(G10), .O(gate28inter7));
  inv1  gate1395(.a(G14), .O(gate28inter8));
  nand2 gate1396(.a(gate28inter8), .b(gate28inter7), .O(gate28inter9));
  nand2 gate1397(.a(s_121), .b(gate28inter3), .O(gate28inter10));
  nor2  gate1398(.a(gate28inter10), .b(gate28inter9), .O(gate28inter11));
  nor2  gate1399(.a(gate28inter11), .b(gate28inter6), .O(gate28inter12));
  nand2 gate1400(.a(gate28inter12), .b(gate28inter1), .O(G323));

  xor2  gate1891(.a(G7), .b(G3), .O(gate29inter0));
  nand2 gate1892(.a(gate29inter0), .b(s_192), .O(gate29inter1));
  and2  gate1893(.a(G7), .b(G3), .O(gate29inter2));
  inv1  gate1894(.a(s_192), .O(gate29inter3));
  inv1  gate1895(.a(s_193), .O(gate29inter4));
  nand2 gate1896(.a(gate29inter4), .b(gate29inter3), .O(gate29inter5));
  nor2  gate1897(.a(gate29inter5), .b(gate29inter2), .O(gate29inter6));
  inv1  gate1898(.a(G3), .O(gate29inter7));
  inv1  gate1899(.a(G7), .O(gate29inter8));
  nand2 gate1900(.a(gate29inter8), .b(gate29inter7), .O(gate29inter9));
  nand2 gate1901(.a(s_193), .b(gate29inter3), .O(gate29inter10));
  nor2  gate1902(.a(gate29inter10), .b(gate29inter9), .O(gate29inter11));
  nor2  gate1903(.a(gate29inter11), .b(gate29inter6), .O(gate29inter12));
  nand2 gate1904(.a(gate29inter12), .b(gate29inter1), .O(G326));

  xor2  gate2815(.a(G15), .b(G11), .O(gate30inter0));
  nand2 gate2816(.a(gate30inter0), .b(s_324), .O(gate30inter1));
  and2  gate2817(.a(G15), .b(G11), .O(gate30inter2));
  inv1  gate2818(.a(s_324), .O(gate30inter3));
  inv1  gate2819(.a(s_325), .O(gate30inter4));
  nand2 gate2820(.a(gate30inter4), .b(gate30inter3), .O(gate30inter5));
  nor2  gate2821(.a(gate30inter5), .b(gate30inter2), .O(gate30inter6));
  inv1  gate2822(.a(G11), .O(gate30inter7));
  inv1  gate2823(.a(G15), .O(gate30inter8));
  nand2 gate2824(.a(gate30inter8), .b(gate30inter7), .O(gate30inter9));
  nand2 gate2825(.a(s_325), .b(gate30inter3), .O(gate30inter10));
  nor2  gate2826(.a(gate30inter10), .b(gate30inter9), .O(gate30inter11));
  nor2  gate2827(.a(gate30inter11), .b(gate30inter6), .O(gate30inter12));
  nand2 gate2828(.a(gate30inter12), .b(gate30inter1), .O(G329));

  xor2  gate1611(.a(G8), .b(G4), .O(gate31inter0));
  nand2 gate1612(.a(gate31inter0), .b(s_152), .O(gate31inter1));
  and2  gate1613(.a(G8), .b(G4), .O(gate31inter2));
  inv1  gate1614(.a(s_152), .O(gate31inter3));
  inv1  gate1615(.a(s_153), .O(gate31inter4));
  nand2 gate1616(.a(gate31inter4), .b(gate31inter3), .O(gate31inter5));
  nor2  gate1617(.a(gate31inter5), .b(gate31inter2), .O(gate31inter6));
  inv1  gate1618(.a(G4), .O(gate31inter7));
  inv1  gate1619(.a(G8), .O(gate31inter8));
  nand2 gate1620(.a(gate31inter8), .b(gate31inter7), .O(gate31inter9));
  nand2 gate1621(.a(s_153), .b(gate31inter3), .O(gate31inter10));
  nor2  gate1622(.a(gate31inter10), .b(gate31inter9), .O(gate31inter11));
  nor2  gate1623(.a(gate31inter11), .b(gate31inter6), .O(gate31inter12));
  nand2 gate1624(.a(gate31inter12), .b(gate31inter1), .O(G332));
nand2 gate32( .a(G12), .b(G16), .O(G335) );
nand2 gate33( .a(G17), .b(G21), .O(G338) );

  xor2  gate2955(.a(G29), .b(G25), .O(gate34inter0));
  nand2 gate2956(.a(gate34inter0), .b(s_344), .O(gate34inter1));
  and2  gate2957(.a(G29), .b(G25), .O(gate34inter2));
  inv1  gate2958(.a(s_344), .O(gate34inter3));
  inv1  gate2959(.a(s_345), .O(gate34inter4));
  nand2 gate2960(.a(gate34inter4), .b(gate34inter3), .O(gate34inter5));
  nor2  gate2961(.a(gate34inter5), .b(gate34inter2), .O(gate34inter6));
  inv1  gate2962(.a(G25), .O(gate34inter7));
  inv1  gate2963(.a(G29), .O(gate34inter8));
  nand2 gate2964(.a(gate34inter8), .b(gate34inter7), .O(gate34inter9));
  nand2 gate2965(.a(s_345), .b(gate34inter3), .O(gate34inter10));
  nor2  gate2966(.a(gate34inter10), .b(gate34inter9), .O(gate34inter11));
  nor2  gate2967(.a(gate34inter11), .b(gate34inter6), .O(gate34inter12));
  nand2 gate2968(.a(gate34inter12), .b(gate34inter1), .O(G341));
nand2 gate35( .a(G18), .b(G22), .O(G344) );
nand2 gate36( .a(G26), .b(G30), .O(G347) );
nand2 gate37( .a(G19), .b(G23), .O(G350) );

  xor2  gate1667(.a(G31), .b(G27), .O(gate38inter0));
  nand2 gate1668(.a(gate38inter0), .b(s_160), .O(gate38inter1));
  and2  gate1669(.a(G31), .b(G27), .O(gate38inter2));
  inv1  gate1670(.a(s_160), .O(gate38inter3));
  inv1  gate1671(.a(s_161), .O(gate38inter4));
  nand2 gate1672(.a(gate38inter4), .b(gate38inter3), .O(gate38inter5));
  nor2  gate1673(.a(gate38inter5), .b(gate38inter2), .O(gate38inter6));
  inv1  gate1674(.a(G27), .O(gate38inter7));
  inv1  gate1675(.a(G31), .O(gate38inter8));
  nand2 gate1676(.a(gate38inter8), .b(gate38inter7), .O(gate38inter9));
  nand2 gate1677(.a(s_161), .b(gate38inter3), .O(gate38inter10));
  nor2  gate1678(.a(gate38inter10), .b(gate38inter9), .O(gate38inter11));
  nor2  gate1679(.a(gate38inter11), .b(gate38inter6), .O(gate38inter12));
  nand2 gate1680(.a(gate38inter12), .b(gate38inter1), .O(G353));
nand2 gate39( .a(G20), .b(G24), .O(G356) );

  xor2  gate1653(.a(G32), .b(G28), .O(gate40inter0));
  nand2 gate1654(.a(gate40inter0), .b(s_158), .O(gate40inter1));
  and2  gate1655(.a(G32), .b(G28), .O(gate40inter2));
  inv1  gate1656(.a(s_158), .O(gate40inter3));
  inv1  gate1657(.a(s_159), .O(gate40inter4));
  nand2 gate1658(.a(gate40inter4), .b(gate40inter3), .O(gate40inter5));
  nor2  gate1659(.a(gate40inter5), .b(gate40inter2), .O(gate40inter6));
  inv1  gate1660(.a(G28), .O(gate40inter7));
  inv1  gate1661(.a(G32), .O(gate40inter8));
  nand2 gate1662(.a(gate40inter8), .b(gate40inter7), .O(gate40inter9));
  nand2 gate1663(.a(s_159), .b(gate40inter3), .O(gate40inter10));
  nor2  gate1664(.a(gate40inter10), .b(gate40inter9), .O(gate40inter11));
  nor2  gate1665(.a(gate40inter11), .b(gate40inter6), .O(gate40inter12));
  nand2 gate1666(.a(gate40inter12), .b(gate40inter1), .O(G359));

  xor2  gate1989(.a(G266), .b(G1), .O(gate41inter0));
  nand2 gate1990(.a(gate41inter0), .b(s_206), .O(gate41inter1));
  and2  gate1991(.a(G266), .b(G1), .O(gate41inter2));
  inv1  gate1992(.a(s_206), .O(gate41inter3));
  inv1  gate1993(.a(s_207), .O(gate41inter4));
  nand2 gate1994(.a(gate41inter4), .b(gate41inter3), .O(gate41inter5));
  nor2  gate1995(.a(gate41inter5), .b(gate41inter2), .O(gate41inter6));
  inv1  gate1996(.a(G1), .O(gate41inter7));
  inv1  gate1997(.a(G266), .O(gate41inter8));
  nand2 gate1998(.a(gate41inter8), .b(gate41inter7), .O(gate41inter9));
  nand2 gate1999(.a(s_207), .b(gate41inter3), .O(gate41inter10));
  nor2  gate2000(.a(gate41inter10), .b(gate41inter9), .O(gate41inter11));
  nor2  gate2001(.a(gate41inter11), .b(gate41inter6), .O(gate41inter12));
  nand2 gate2002(.a(gate41inter12), .b(gate41inter1), .O(G362));
nand2 gate42( .a(G2), .b(G266), .O(G363) );

  xor2  gate2129(.a(G269), .b(G3), .O(gate43inter0));
  nand2 gate2130(.a(gate43inter0), .b(s_226), .O(gate43inter1));
  and2  gate2131(.a(G269), .b(G3), .O(gate43inter2));
  inv1  gate2132(.a(s_226), .O(gate43inter3));
  inv1  gate2133(.a(s_227), .O(gate43inter4));
  nand2 gate2134(.a(gate43inter4), .b(gate43inter3), .O(gate43inter5));
  nor2  gate2135(.a(gate43inter5), .b(gate43inter2), .O(gate43inter6));
  inv1  gate2136(.a(G3), .O(gate43inter7));
  inv1  gate2137(.a(G269), .O(gate43inter8));
  nand2 gate2138(.a(gate43inter8), .b(gate43inter7), .O(gate43inter9));
  nand2 gate2139(.a(s_227), .b(gate43inter3), .O(gate43inter10));
  nor2  gate2140(.a(gate43inter10), .b(gate43inter9), .O(gate43inter11));
  nor2  gate2141(.a(gate43inter11), .b(gate43inter6), .O(gate43inter12));
  nand2 gate2142(.a(gate43inter12), .b(gate43inter1), .O(G364));

  xor2  gate1849(.a(G269), .b(G4), .O(gate44inter0));
  nand2 gate1850(.a(gate44inter0), .b(s_186), .O(gate44inter1));
  and2  gate1851(.a(G269), .b(G4), .O(gate44inter2));
  inv1  gate1852(.a(s_186), .O(gate44inter3));
  inv1  gate1853(.a(s_187), .O(gate44inter4));
  nand2 gate1854(.a(gate44inter4), .b(gate44inter3), .O(gate44inter5));
  nor2  gate1855(.a(gate44inter5), .b(gate44inter2), .O(gate44inter6));
  inv1  gate1856(.a(G4), .O(gate44inter7));
  inv1  gate1857(.a(G269), .O(gate44inter8));
  nand2 gate1858(.a(gate44inter8), .b(gate44inter7), .O(gate44inter9));
  nand2 gate1859(.a(s_187), .b(gate44inter3), .O(gate44inter10));
  nor2  gate1860(.a(gate44inter10), .b(gate44inter9), .O(gate44inter11));
  nor2  gate1861(.a(gate44inter11), .b(gate44inter6), .O(gate44inter12));
  nand2 gate1862(.a(gate44inter12), .b(gate44inter1), .O(G365));

  xor2  gate1219(.a(G272), .b(G5), .O(gate45inter0));
  nand2 gate1220(.a(gate45inter0), .b(s_96), .O(gate45inter1));
  and2  gate1221(.a(G272), .b(G5), .O(gate45inter2));
  inv1  gate1222(.a(s_96), .O(gate45inter3));
  inv1  gate1223(.a(s_97), .O(gate45inter4));
  nand2 gate1224(.a(gate45inter4), .b(gate45inter3), .O(gate45inter5));
  nor2  gate1225(.a(gate45inter5), .b(gate45inter2), .O(gate45inter6));
  inv1  gate1226(.a(G5), .O(gate45inter7));
  inv1  gate1227(.a(G272), .O(gate45inter8));
  nand2 gate1228(.a(gate45inter8), .b(gate45inter7), .O(gate45inter9));
  nand2 gate1229(.a(s_97), .b(gate45inter3), .O(gate45inter10));
  nor2  gate1230(.a(gate45inter10), .b(gate45inter9), .O(gate45inter11));
  nor2  gate1231(.a(gate45inter11), .b(gate45inter6), .O(gate45inter12));
  nand2 gate1232(.a(gate45inter12), .b(gate45inter1), .O(G366));

  xor2  gate1317(.a(G272), .b(G6), .O(gate46inter0));
  nand2 gate1318(.a(gate46inter0), .b(s_110), .O(gate46inter1));
  and2  gate1319(.a(G272), .b(G6), .O(gate46inter2));
  inv1  gate1320(.a(s_110), .O(gate46inter3));
  inv1  gate1321(.a(s_111), .O(gate46inter4));
  nand2 gate1322(.a(gate46inter4), .b(gate46inter3), .O(gate46inter5));
  nor2  gate1323(.a(gate46inter5), .b(gate46inter2), .O(gate46inter6));
  inv1  gate1324(.a(G6), .O(gate46inter7));
  inv1  gate1325(.a(G272), .O(gate46inter8));
  nand2 gate1326(.a(gate46inter8), .b(gate46inter7), .O(gate46inter9));
  nand2 gate1327(.a(s_111), .b(gate46inter3), .O(gate46inter10));
  nor2  gate1328(.a(gate46inter10), .b(gate46inter9), .O(gate46inter11));
  nor2  gate1329(.a(gate46inter11), .b(gate46inter6), .O(gate46inter12));
  nand2 gate1330(.a(gate46inter12), .b(gate46inter1), .O(G367));

  xor2  gate2073(.a(G275), .b(G7), .O(gate47inter0));
  nand2 gate2074(.a(gate47inter0), .b(s_218), .O(gate47inter1));
  and2  gate2075(.a(G275), .b(G7), .O(gate47inter2));
  inv1  gate2076(.a(s_218), .O(gate47inter3));
  inv1  gate2077(.a(s_219), .O(gate47inter4));
  nand2 gate2078(.a(gate47inter4), .b(gate47inter3), .O(gate47inter5));
  nor2  gate2079(.a(gate47inter5), .b(gate47inter2), .O(gate47inter6));
  inv1  gate2080(.a(G7), .O(gate47inter7));
  inv1  gate2081(.a(G275), .O(gate47inter8));
  nand2 gate2082(.a(gate47inter8), .b(gate47inter7), .O(gate47inter9));
  nand2 gate2083(.a(s_219), .b(gate47inter3), .O(gate47inter10));
  nor2  gate2084(.a(gate47inter10), .b(gate47inter9), .O(gate47inter11));
  nor2  gate2085(.a(gate47inter11), .b(gate47inter6), .O(gate47inter12));
  nand2 gate2086(.a(gate47inter12), .b(gate47inter1), .O(G368));

  xor2  gate2731(.a(G275), .b(G8), .O(gate48inter0));
  nand2 gate2732(.a(gate48inter0), .b(s_312), .O(gate48inter1));
  and2  gate2733(.a(G275), .b(G8), .O(gate48inter2));
  inv1  gate2734(.a(s_312), .O(gate48inter3));
  inv1  gate2735(.a(s_313), .O(gate48inter4));
  nand2 gate2736(.a(gate48inter4), .b(gate48inter3), .O(gate48inter5));
  nor2  gate2737(.a(gate48inter5), .b(gate48inter2), .O(gate48inter6));
  inv1  gate2738(.a(G8), .O(gate48inter7));
  inv1  gate2739(.a(G275), .O(gate48inter8));
  nand2 gate2740(.a(gate48inter8), .b(gate48inter7), .O(gate48inter9));
  nand2 gate2741(.a(s_313), .b(gate48inter3), .O(gate48inter10));
  nor2  gate2742(.a(gate48inter10), .b(gate48inter9), .O(gate48inter11));
  nor2  gate2743(.a(gate48inter11), .b(gate48inter6), .O(gate48inter12));
  nand2 gate2744(.a(gate48inter12), .b(gate48inter1), .O(G369));

  xor2  gate2801(.a(G278), .b(G9), .O(gate49inter0));
  nand2 gate2802(.a(gate49inter0), .b(s_322), .O(gate49inter1));
  and2  gate2803(.a(G278), .b(G9), .O(gate49inter2));
  inv1  gate2804(.a(s_322), .O(gate49inter3));
  inv1  gate2805(.a(s_323), .O(gate49inter4));
  nand2 gate2806(.a(gate49inter4), .b(gate49inter3), .O(gate49inter5));
  nor2  gate2807(.a(gate49inter5), .b(gate49inter2), .O(gate49inter6));
  inv1  gate2808(.a(G9), .O(gate49inter7));
  inv1  gate2809(.a(G278), .O(gate49inter8));
  nand2 gate2810(.a(gate49inter8), .b(gate49inter7), .O(gate49inter9));
  nand2 gate2811(.a(s_323), .b(gate49inter3), .O(gate49inter10));
  nor2  gate2812(.a(gate49inter10), .b(gate49inter9), .O(gate49inter11));
  nor2  gate2813(.a(gate49inter11), .b(gate49inter6), .O(gate49inter12));
  nand2 gate2814(.a(gate49inter12), .b(gate49inter1), .O(G370));
nand2 gate50( .a(G10), .b(G278), .O(G371) );
nand2 gate51( .a(G11), .b(G281), .O(G372) );

  xor2  gate3025(.a(G281), .b(G12), .O(gate52inter0));
  nand2 gate3026(.a(gate52inter0), .b(s_354), .O(gate52inter1));
  and2  gate3027(.a(G281), .b(G12), .O(gate52inter2));
  inv1  gate3028(.a(s_354), .O(gate52inter3));
  inv1  gate3029(.a(s_355), .O(gate52inter4));
  nand2 gate3030(.a(gate52inter4), .b(gate52inter3), .O(gate52inter5));
  nor2  gate3031(.a(gate52inter5), .b(gate52inter2), .O(gate52inter6));
  inv1  gate3032(.a(G12), .O(gate52inter7));
  inv1  gate3033(.a(G281), .O(gate52inter8));
  nand2 gate3034(.a(gate52inter8), .b(gate52inter7), .O(gate52inter9));
  nand2 gate3035(.a(s_355), .b(gate52inter3), .O(gate52inter10));
  nor2  gate3036(.a(gate52inter10), .b(gate52inter9), .O(gate52inter11));
  nor2  gate3037(.a(gate52inter11), .b(gate52inter6), .O(gate52inter12));
  nand2 gate3038(.a(gate52inter12), .b(gate52inter1), .O(G373));
nand2 gate53( .a(G13), .b(G284), .O(G374) );

  xor2  gate3011(.a(G284), .b(G14), .O(gate54inter0));
  nand2 gate3012(.a(gate54inter0), .b(s_352), .O(gate54inter1));
  and2  gate3013(.a(G284), .b(G14), .O(gate54inter2));
  inv1  gate3014(.a(s_352), .O(gate54inter3));
  inv1  gate3015(.a(s_353), .O(gate54inter4));
  nand2 gate3016(.a(gate54inter4), .b(gate54inter3), .O(gate54inter5));
  nor2  gate3017(.a(gate54inter5), .b(gate54inter2), .O(gate54inter6));
  inv1  gate3018(.a(G14), .O(gate54inter7));
  inv1  gate3019(.a(G284), .O(gate54inter8));
  nand2 gate3020(.a(gate54inter8), .b(gate54inter7), .O(gate54inter9));
  nand2 gate3021(.a(s_353), .b(gate54inter3), .O(gate54inter10));
  nor2  gate3022(.a(gate54inter10), .b(gate54inter9), .O(gate54inter11));
  nor2  gate3023(.a(gate54inter11), .b(gate54inter6), .O(gate54inter12));
  nand2 gate3024(.a(gate54inter12), .b(gate54inter1), .O(G375));

  xor2  gate547(.a(G287), .b(G15), .O(gate55inter0));
  nand2 gate548(.a(gate55inter0), .b(s_0), .O(gate55inter1));
  and2  gate549(.a(G287), .b(G15), .O(gate55inter2));
  inv1  gate550(.a(s_0), .O(gate55inter3));
  inv1  gate551(.a(s_1), .O(gate55inter4));
  nand2 gate552(.a(gate55inter4), .b(gate55inter3), .O(gate55inter5));
  nor2  gate553(.a(gate55inter5), .b(gate55inter2), .O(gate55inter6));
  inv1  gate554(.a(G15), .O(gate55inter7));
  inv1  gate555(.a(G287), .O(gate55inter8));
  nand2 gate556(.a(gate55inter8), .b(gate55inter7), .O(gate55inter9));
  nand2 gate557(.a(s_1), .b(gate55inter3), .O(gate55inter10));
  nor2  gate558(.a(gate55inter10), .b(gate55inter9), .O(gate55inter11));
  nor2  gate559(.a(gate55inter11), .b(gate55inter6), .O(gate55inter12));
  nand2 gate560(.a(gate55inter12), .b(gate55inter1), .O(G376));
nand2 gate56( .a(G16), .b(G287), .O(G377) );

  xor2  gate1107(.a(G290), .b(G17), .O(gate57inter0));
  nand2 gate1108(.a(gate57inter0), .b(s_80), .O(gate57inter1));
  and2  gate1109(.a(G290), .b(G17), .O(gate57inter2));
  inv1  gate1110(.a(s_80), .O(gate57inter3));
  inv1  gate1111(.a(s_81), .O(gate57inter4));
  nand2 gate1112(.a(gate57inter4), .b(gate57inter3), .O(gate57inter5));
  nor2  gate1113(.a(gate57inter5), .b(gate57inter2), .O(gate57inter6));
  inv1  gate1114(.a(G17), .O(gate57inter7));
  inv1  gate1115(.a(G290), .O(gate57inter8));
  nand2 gate1116(.a(gate57inter8), .b(gate57inter7), .O(gate57inter9));
  nand2 gate1117(.a(s_81), .b(gate57inter3), .O(gate57inter10));
  nor2  gate1118(.a(gate57inter10), .b(gate57inter9), .O(gate57inter11));
  nor2  gate1119(.a(gate57inter11), .b(gate57inter6), .O(gate57inter12));
  nand2 gate1120(.a(gate57inter12), .b(gate57inter1), .O(G378));

  xor2  gate1401(.a(G290), .b(G18), .O(gate58inter0));
  nand2 gate1402(.a(gate58inter0), .b(s_122), .O(gate58inter1));
  and2  gate1403(.a(G290), .b(G18), .O(gate58inter2));
  inv1  gate1404(.a(s_122), .O(gate58inter3));
  inv1  gate1405(.a(s_123), .O(gate58inter4));
  nand2 gate1406(.a(gate58inter4), .b(gate58inter3), .O(gate58inter5));
  nor2  gate1407(.a(gate58inter5), .b(gate58inter2), .O(gate58inter6));
  inv1  gate1408(.a(G18), .O(gate58inter7));
  inv1  gate1409(.a(G290), .O(gate58inter8));
  nand2 gate1410(.a(gate58inter8), .b(gate58inter7), .O(gate58inter9));
  nand2 gate1411(.a(s_123), .b(gate58inter3), .O(gate58inter10));
  nor2  gate1412(.a(gate58inter10), .b(gate58inter9), .O(gate58inter11));
  nor2  gate1413(.a(gate58inter11), .b(gate58inter6), .O(gate58inter12));
  nand2 gate1414(.a(gate58inter12), .b(gate58inter1), .O(G379));
nand2 gate59( .a(G19), .b(G293), .O(G380) );

  xor2  gate589(.a(G293), .b(G20), .O(gate60inter0));
  nand2 gate590(.a(gate60inter0), .b(s_6), .O(gate60inter1));
  and2  gate591(.a(G293), .b(G20), .O(gate60inter2));
  inv1  gate592(.a(s_6), .O(gate60inter3));
  inv1  gate593(.a(s_7), .O(gate60inter4));
  nand2 gate594(.a(gate60inter4), .b(gate60inter3), .O(gate60inter5));
  nor2  gate595(.a(gate60inter5), .b(gate60inter2), .O(gate60inter6));
  inv1  gate596(.a(G20), .O(gate60inter7));
  inv1  gate597(.a(G293), .O(gate60inter8));
  nand2 gate598(.a(gate60inter8), .b(gate60inter7), .O(gate60inter9));
  nand2 gate599(.a(s_7), .b(gate60inter3), .O(gate60inter10));
  nor2  gate600(.a(gate60inter10), .b(gate60inter9), .O(gate60inter11));
  nor2  gate601(.a(gate60inter11), .b(gate60inter6), .O(gate60inter12));
  nand2 gate602(.a(gate60inter12), .b(gate60inter1), .O(G381));

  xor2  gate1303(.a(G296), .b(G21), .O(gate61inter0));
  nand2 gate1304(.a(gate61inter0), .b(s_108), .O(gate61inter1));
  and2  gate1305(.a(G296), .b(G21), .O(gate61inter2));
  inv1  gate1306(.a(s_108), .O(gate61inter3));
  inv1  gate1307(.a(s_109), .O(gate61inter4));
  nand2 gate1308(.a(gate61inter4), .b(gate61inter3), .O(gate61inter5));
  nor2  gate1309(.a(gate61inter5), .b(gate61inter2), .O(gate61inter6));
  inv1  gate1310(.a(G21), .O(gate61inter7));
  inv1  gate1311(.a(G296), .O(gate61inter8));
  nand2 gate1312(.a(gate61inter8), .b(gate61inter7), .O(gate61inter9));
  nand2 gate1313(.a(s_109), .b(gate61inter3), .O(gate61inter10));
  nor2  gate1314(.a(gate61inter10), .b(gate61inter9), .O(gate61inter11));
  nor2  gate1315(.a(gate61inter11), .b(gate61inter6), .O(gate61inter12));
  nand2 gate1316(.a(gate61inter12), .b(gate61inter1), .O(G382));

  xor2  gate2199(.a(G296), .b(G22), .O(gate62inter0));
  nand2 gate2200(.a(gate62inter0), .b(s_236), .O(gate62inter1));
  and2  gate2201(.a(G296), .b(G22), .O(gate62inter2));
  inv1  gate2202(.a(s_236), .O(gate62inter3));
  inv1  gate2203(.a(s_237), .O(gate62inter4));
  nand2 gate2204(.a(gate62inter4), .b(gate62inter3), .O(gate62inter5));
  nor2  gate2205(.a(gate62inter5), .b(gate62inter2), .O(gate62inter6));
  inv1  gate2206(.a(G22), .O(gate62inter7));
  inv1  gate2207(.a(G296), .O(gate62inter8));
  nand2 gate2208(.a(gate62inter8), .b(gate62inter7), .O(gate62inter9));
  nand2 gate2209(.a(s_237), .b(gate62inter3), .O(gate62inter10));
  nor2  gate2210(.a(gate62inter10), .b(gate62inter9), .O(gate62inter11));
  nor2  gate2211(.a(gate62inter11), .b(gate62inter6), .O(gate62inter12));
  nand2 gate2212(.a(gate62inter12), .b(gate62inter1), .O(G383));

  xor2  gate1261(.a(G299), .b(G23), .O(gate63inter0));
  nand2 gate1262(.a(gate63inter0), .b(s_102), .O(gate63inter1));
  and2  gate1263(.a(G299), .b(G23), .O(gate63inter2));
  inv1  gate1264(.a(s_102), .O(gate63inter3));
  inv1  gate1265(.a(s_103), .O(gate63inter4));
  nand2 gate1266(.a(gate63inter4), .b(gate63inter3), .O(gate63inter5));
  nor2  gate1267(.a(gate63inter5), .b(gate63inter2), .O(gate63inter6));
  inv1  gate1268(.a(G23), .O(gate63inter7));
  inv1  gate1269(.a(G299), .O(gate63inter8));
  nand2 gate1270(.a(gate63inter8), .b(gate63inter7), .O(gate63inter9));
  nand2 gate1271(.a(s_103), .b(gate63inter3), .O(gate63inter10));
  nor2  gate1272(.a(gate63inter10), .b(gate63inter9), .O(gate63inter11));
  nor2  gate1273(.a(gate63inter11), .b(gate63inter6), .O(gate63inter12));
  nand2 gate1274(.a(gate63inter12), .b(gate63inter1), .O(G384));

  xor2  gate2591(.a(G299), .b(G24), .O(gate64inter0));
  nand2 gate2592(.a(gate64inter0), .b(s_292), .O(gate64inter1));
  and2  gate2593(.a(G299), .b(G24), .O(gate64inter2));
  inv1  gate2594(.a(s_292), .O(gate64inter3));
  inv1  gate2595(.a(s_293), .O(gate64inter4));
  nand2 gate2596(.a(gate64inter4), .b(gate64inter3), .O(gate64inter5));
  nor2  gate2597(.a(gate64inter5), .b(gate64inter2), .O(gate64inter6));
  inv1  gate2598(.a(G24), .O(gate64inter7));
  inv1  gate2599(.a(G299), .O(gate64inter8));
  nand2 gate2600(.a(gate64inter8), .b(gate64inter7), .O(gate64inter9));
  nand2 gate2601(.a(s_293), .b(gate64inter3), .O(gate64inter10));
  nor2  gate2602(.a(gate64inter10), .b(gate64inter9), .O(gate64inter11));
  nor2  gate2603(.a(gate64inter11), .b(gate64inter6), .O(gate64inter12));
  nand2 gate2604(.a(gate64inter12), .b(gate64inter1), .O(G385));
nand2 gate65( .a(G25), .b(G302), .O(G386) );

  xor2  gate2171(.a(G302), .b(G26), .O(gate66inter0));
  nand2 gate2172(.a(gate66inter0), .b(s_232), .O(gate66inter1));
  and2  gate2173(.a(G302), .b(G26), .O(gate66inter2));
  inv1  gate2174(.a(s_232), .O(gate66inter3));
  inv1  gate2175(.a(s_233), .O(gate66inter4));
  nand2 gate2176(.a(gate66inter4), .b(gate66inter3), .O(gate66inter5));
  nor2  gate2177(.a(gate66inter5), .b(gate66inter2), .O(gate66inter6));
  inv1  gate2178(.a(G26), .O(gate66inter7));
  inv1  gate2179(.a(G302), .O(gate66inter8));
  nand2 gate2180(.a(gate66inter8), .b(gate66inter7), .O(gate66inter9));
  nand2 gate2181(.a(s_233), .b(gate66inter3), .O(gate66inter10));
  nor2  gate2182(.a(gate66inter10), .b(gate66inter9), .O(gate66inter11));
  nor2  gate2183(.a(gate66inter11), .b(gate66inter6), .O(gate66inter12));
  nand2 gate2184(.a(gate66inter12), .b(gate66inter1), .O(G387));
nand2 gate67( .a(G27), .b(G305), .O(G388) );
nand2 gate68( .a(G28), .b(G305), .O(G389) );

  xor2  gate1597(.a(G308), .b(G29), .O(gate69inter0));
  nand2 gate1598(.a(gate69inter0), .b(s_150), .O(gate69inter1));
  and2  gate1599(.a(G308), .b(G29), .O(gate69inter2));
  inv1  gate1600(.a(s_150), .O(gate69inter3));
  inv1  gate1601(.a(s_151), .O(gate69inter4));
  nand2 gate1602(.a(gate69inter4), .b(gate69inter3), .O(gate69inter5));
  nor2  gate1603(.a(gate69inter5), .b(gate69inter2), .O(gate69inter6));
  inv1  gate1604(.a(G29), .O(gate69inter7));
  inv1  gate1605(.a(G308), .O(gate69inter8));
  nand2 gate1606(.a(gate69inter8), .b(gate69inter7), .O(gate69inter9));
  nand2 gate1607(.a(s_151), .b(gate69inter3), .O(gate69inter10));
  nor2  gate1608(.a(gate69inter10), .b(gate69inter9), .O(gate69inter11));
  nor2  gate1609(.a(gate69inter11), .b(gate69inter6), .O(gate69inter12));
  nand2 gate1610(.a(gate69inter12), .b(gate69inter1), .O(G390));

  xor2  gate1583(.a(G308), .b(G30), .O(gate70inter0));
  nand2 gate1584(.a(gate70inter0), .b(s_148), .O(gate70inter1));
  and2  gate1585(.a(G308), .b(G30), .O(gate70inter2));
  inv1  gate1586(.a(s_148), .O(gate70inter3));
  inv1  gate1587(.a(s_149), .O(gate70inter4));
  nand2 gate1588(.a(gate70inter4), .b(gate70inter3), .O(gate70inter5));
  nor2  gate1589(.a(gate70inter5), .b(gate70inter2), .O(gate70inter6));
  inv1  gate1590(.a(G30), .O(gate70inter7));
  inv1  gate1591(.a(G308), .O(gate70inter8));
  nand2 gate1592(.a(gate70inter8), .b(gate70inter7), .O(gate70inter9));
  nand2 gate1593(.a(s_149), .b(gate70inter3), .O(gate70inter10));
  nor2  gate1594(.a(gate70inter10), .b(gate70inter9), .O(gate70inter11));
  nor2  gate1595(.a(gate70inter11), .b(gate70inter6), .O(gate70inter12));
  nand2 gate1596(.a(gate70inter12), .b(gate70inter1), .O(G391));

  xor2  gate2339(.a(G311), .b(G31), .O(gate71inter0));
  nand2 gate2340(.a(gate71inter0), .b(s_256), .O(gate71inter1));
  and2  gate2341(.a(G311), .b(G31), .O(gate71inter2));
  inv1  gate2342(.a(s_256), .O(gate71inter3));
  inv1  gate2343(.a(s_257), .O(gate71inter4));
  nand2 gate2344(.a(gate71inter4), .b(gate71inter3), .O(gate71inter5));
  nor2  gate2345(.a(gate71inter5), .b(gate71inter2), .O(gate71inter6));
  inv1  gate2346(.a(G31), .O(gate71inter7));
  inv1  gate2347(.a(G311), .O(gate71inter8));
  nand2 gate2348(.a(gate71inter8), .b(gate71inter7), .O(gate71inter9));
  nand2 gate2349(.a(s_257), .b(gate71inter3), .O(gate71inter10));
  nor2  gate2350(.a(gate71inter10), .b(gate71inter9), .O(gate71inter11));
  nor2  gate2351(.a(gate71inter11), .b(gate71inter6), .O(gate71inter12));
  nand2 gate2352(.a(gate71inter12), .b(gate71inter1), .O(G392));

  xor2  gate2241(.a(G311), .b(G32), .O(gate72inter0));
  nand2 gate2242(.a(gate72inter0), .b(s_242), .O(gate72inter1));
  and2  gate2243(.a(G311), .b(G32), .O(gate72inter2));
  inv1  gate2244(.a(s_242), .O(gate72inter3));
  inv1  gate2245(.a(s_243), .O(gate72inter4));
  nand2 gate2246(.a(gate72inter4), .b(gate72inter3), .O(gate72inter5));
  nor2  gate2247(.a(gate72inter5), .b(gate72inter2), .O(gate72inter6));
  inv1  gate2248(.a(G32), .O(gate72inter7));
  inv1  gate2249(.a(G311), .O(gate72inter8));
  nand2 gate2250(.a(gate72inter8), .b(gate72inter7), .O(gate72inter9));
  nand2 gate2251(.a(s_243), .b(gate72inter3), .O(gate72inter10));
  nor2  gate2252(.a(gate72inter10), .b(gate72inter9), .O(gate72inter11));
  nor2  gate2253(.a(gate72inter11), .b(gate72inter6), .O(gate72inter12));
  nand2 gate2254(.a(gate72inter12), .b(gate72inter1), .O(G393));
nand2 gate73( .a(G1), .b(G314), .O(G394) );
nand2 gate74( .a(G5), .b(G314), .O(G395) );
nand2 gate75( .a(G9), .b(G317), .O(G396) );

  xor2  gate2787(.a(G317), .b(G13), .O(gate76inter0));
  nand2 gate2788(.a(gate76inter0), .b(s_320), .O(gate76inter1));
  and2  gate2789(.a(G317), .b(G13), .O(gate76inter2));
  inv1  gate2790(.a(s_320), .O(gate76inter3));
  inv1  gate2791(.a(s_321), .O(gate76inter4));
  nand2 gate2792(.a(gate76inter4), .b(gate76inter3), .O(gate76inter5));
  nor2  gate2793(.a(gate76inter5), .b(gate76inter2), .O(gate76inter6));
  inv1  gate2794(.a(G13), .O(gate76inter7));
  inv1  gate2795(.a(G317), .O(gate76inter8));
  nand2 gate2796(.a(gate76inter8), .b(gate76inter7), .O(gate76inter9));
  nand2 gate2797(.a(s_321), .b(gate76inter3), .O(gate76inter10));
  nor2  gate2798(.a(gate76inter10), .b(gate76inter9), .O(gate76inter11));
  nor2  gate2799(.a(gate76inter11), .b(gate76inter6), .O(gate76inter12));
  nand2 gate2800(.a(gate76inter12), .b(gate76inter1), .O(G397));
nand2 gate77( .a(G2), .b(G320), .O(G398) );

  xor2  gate2577(.a(G320), .b(G6), .O(gate78inter0));
  nand2 gate2578(.a(gate78inter0), .b(s_290), .O(gate78inter1));
  and2  gate2579(.a(G320), .b(G6), .O(gate78inter2));
  inv1  gate2580(.a(s_290), .O(gate78inter3));
  inv1  gate2581(.a(s_291), .O(gate78inter4));
  nand2 gate2582(.a(gate78inter4), .b(gate78inter3), .O(gate78inter5));
  nor2  gate2583(.a(gate78inter5), .b(gate78inter2), .O(gate78inter6));
  inv1  gate2584(.a(G6), .O(gate78inter7));
  inv1  gate2585(.a(G320), .O(gate78inter8));
  nand2 gate2586(.a(gate78inter8), .b(gate78inter7), .O(gate78inter9));
  nand2 gate2587(.a(s_291), .b(gate78inter3), .O(gate78inter10));
  nor2  gate2588(.a(gate78inter10), .b(gate78inter9), .O(gate78inter11));
  nor2  gate2589(.a(gate78inter11), .b(gate78inter6), .O(gate78inter12));
  nand2 gate2590(.a(gate78inter12), .b(gate78inter1), .O(G399));

  xor2  gate2605(.a(G323), .b(G10), .O(gate79inter0));
  nand2 gate2606(.a(gate79inter0), .b(s_294), .O(gate79inter1));
  and2  gate2607(.a(G323), .b(G10), .O(gate79inter2));
  inv1  gate2608(.a(s_294), .O(gate79inter3));
  inv1  gate2609(.a(s_295), .O(gate79inter4));
  nand2 gate2610(.a(gate79inter4), .b(gate79inter3), .O(gate79inter5));
  nor2  gate2611(.a(gate79inter5), .b(gate79inter2), .O(gate79inter6));
  inv1  gate2612(.a(G10), .O(gate79inter7));
  inv1  gate2613(.a(G323), .O(gate79inter8));
  nand2 gate2614(.a(gate79inter8), .b(gate79inter7), .O(gate79inter9));
  nand2 gate2615(.a(s_295), .b(gate79inter3), .O(gate79inter10));
  nor2  gate2616(.a(gate79inter10), .b(gate79inter9), .O(gate79inter11));
  nor2  gate2617(.a(gate79inter11), .b(gate79inter6), .O(gate79inter12));
  nand2 gate2618(.a(gate79inter12), .b(gate79inter1), .O(G400));
nand2 gate80( .a(G14), .b(G323), .O(G401) );
nand2 gate81( .a(G3), .b(G326), .O(G402) );
nand2 gate82( .a(G7), .b(G326), .O(G403) );
nand2 gate83( .a(G11), .b(G329), .O(G404) );

  xor2  gate2745(.a(G329), .b(G15), .O(gate84inter0));
  nand2 gate2746(.a(gate84inter0), .b(s_314), .O(gate84inter1));
  and2  gate2747(.a(G329), .b(G15), .O(gate84inter2));
  inv1  gate2748(.a(s_314), .O(gate84inter3));
  inv1  gate2749(.a(s_315), .O(gate84inter4));
  nand2 gate2750(.a(gate84inter4), .b(gate84inter3), .O(gate84inter5));
  nor2  gate2751(.a(gate84inter5), .b(gate84inter2), .O(gate84inter6));
  inv1  gate2752(.a(G15), .O(gate84inter7));
  inv1  gate2753(.a(G329), .O(gate84inter8));
  nand2 gate2754(.a(gate84inter8), .b(gate84inter7), .O(gate84inter9));
  nand2 gate2755(.a(s_315), .b(gate84inter3), .O(gate84inter10));
  nor2  gate2756(.a(gate84inter10), .b(gate84inter9), .O(gate84inter11));
  nor2  gate2757(.a(gate84inter11), .b(gate84inter6), .O(gate84inter12));
  nand2 gate2758(.a(gate84inter12), .b(gate84inter1), .O(G405));

  xor2  gate1793(.a(G332), .b(G4), .O(gate85inter0));
  nand2 gate1794(.a(gate85inter0), .b(s_178), .O(gate85inter1));
  and2  gate1795(.a(G332), .b(G4), .O(gate85inter2));
  inv1  gate1796(.a(s_178), .O(gate85inter3));
  inv1  gate1797(.a(s_179), .O(gate85inter4));
  nand2 gate1798(.a(gate85inter4), .b(gate85inter3), .O(gate85inter5));
  nor2  gate1799(.a(gate85inter5), .b(gate85inter2), .O(gate85inter6));
  inv1  gate1800(.a(G4), .O(gate85inter7));
  inv1  gate1801(.a(G332), .O(gate85inter8));
  nand2 gate1802(.a(gate85inter8), .b(gate85inter7), .O(gate85inter9));
  nand2 gate1803(.a(s_179), .b(gate85inter3), .O(gate85inter10));
  nor2  gate1804(.a(gate85inter10), .b(gate85inter9), .O(gate85inter11));
  nor2  gate1805(.a(gate85inter11), .b(gate85inter6), .O(gate85inter12));
  nand2 gate1806(.a(gate85inter12), .b(gate85inter1), .O(G406));
nand2 gate86( .a(G8), .b(G332), .O(G407) );

  xor2  gate1023(.a(G335), .b(G12), .O(gate87inter0));
  nand2 gate1024(.a(gate87inter0), .b(s_68), .O(gate87inter1));
  and2  gate1025(.a(G335), .b(G12), .O(gate87inter2));
  inv1  gate1026(.a(s_68), .O(gate87inter3));
  inv1  gate1027(.a(s_69), .O(gate87inter4));
  nand2 gate1028(.a(gate87inter4), .b(gate87inter3), .O(gate87inter5));
  nor2  gate1029(.a(gate87inter5), .b(gate87inter2), .O(gate87inter6));
  inv1  gate1030(.a(G12), .O(gate87inter7));
  inv1  gate1031(.a(G335), .O(gate87inter8));
  nand2 gate1032(.a(gate87inter8), .b(gate87inter7), .O(gate87inter9));
  nand2 gate1033(.a(s_69), .b(gate87inter3), .O(gate87inter10));
  nor2  gate1034(.a(gate87inter10), .b(gate87inter9), .O(gate87inter11));
  nor2  gate1035(.a(gate87inter11), .b(gate87inter6), .O(gate87inter12));
  nand2 gate1036(.a(gate87inter12), .b(gate87inter1), .O(G408));
nand2 gate88( .a(G16), .b(G335), .O(G409) );
nand2 gate89( .a(G17), .b(G338), .O(G410) );

  xor2  gate2325(.a(G338), .b(G21), .O(gate90inter0));
  nand2 gate2326(.a(gate90inter0), .b(s_254), .O(gate90inter1));
  and2  gate2327(.a(G338), .b(G21), .O(gate90inter2));
  inv1  gate2328(.a(s_254), .O(gate90inter3));
  inv1  gate2329(.a(s_255), .O(gate90inter4));
  nand2 gate2330(.a(gate90inter4), .b(gate90inter3), .O(gate90inter5));
  nor2  gate2331(.a(gate90inter5), .b(gate90inter2), .O(gate90inter6));
  inv1  gate2332(.a(G21), .O(gate90inter7));
  inv1  gate2333(.a(G338), .O(gate90inter8));
  nand2 gate2334(.a(gate90inter8), .b(gate90inter7), .O(gate90inter9));
  nand2 gate2335(.a(s_255), .b(gate90inter3), .O(gate90inter10));
  nor2  gate2336(.a(gate90inter10), .b(gate90inter9), .O(gate90inter11));
  nor2  gate2337(.a(gate90inter11), .b(gate90inter6), .O(gate90inter12));
  nand2 gate2338(.a(gate90inter12), .b(gate90inter1), .O(G411));
nand2 gate91( .a(G25), .b(G341), .O(G412) );
nand2 gate92( .a(G29), .b(G341), .O(G413) );

  xor2  gate701(.a(G344), .b(G18), .O(gate93inter0));
  nand2 gate702(.a(gate93inter0), .b(s_22), .O(gate93inter1));
  and2  gate703(.a(G344), .b(G18), .O(gate93inter2));
  inv1  gate704(.a(s_22), .O(gate93inter3));
  inv1  gate705(.a(s_23), .O(gate93inter4));
  nand2 gate706(.a(gate93inter4), .b(gate93inter3), .O(gate93inter5));
  nor2  gate707(.a(gate93inter5), .b(gate93inter2), .O(gate93inter6));
  inv1  gate708(.a(G18), .O(gate93inter7));
  inv1  gate709(.a(G344), .O(gate93inter8));
  nand2 gate710(.a(gate93inter8), .b(gate93inter7), .O(gate93inter9));
  nand2 gate711(.a(s_23), .b(gate93inter3), .O(gate93inter10));
  nor2  gate712(.a(gate93inter10), .b(gate93inter9), .O(gate93inter11));
  nor2  gate713(.a(gate93inter11), .b(gate93inter6), .O(gate93inter12));
  nand2 gate714(.a(gate93inter12), .b(gate93inter1), .O(G414));

  xor2  gate603(.a(G344), .b(G22), .O(gate94inter0));
  nand2 gate604(.a(gate94inter0), .b(s_8), .O(gate94inter1));
  and2  gate605(.a(G344), .b(G22), .O(gate94inter2));
  inv1  gate606(.a(s_8), .O(gate94inter3));
  inv1  gate607(.a(s_9), .O(gate94inter4));
  nand2 gate608(.a(gate94inter4), .b(gate94inter3), .O(gate94inter5));
  nor2  gate609(.a(gate94inter5), .b(gate94inter2), .O(gate94inter6));
  inv1  gate610(.a(G22), .O(gate94inter7));
  inv1  gate611(.a(G344), .O(gate94inter8));
  nand2 gate612(.a(gate94inter8), .b(gate94inter7), .O(gate94inter9));
  nand2 gate613(.a(s_9), .b(gate94inter3), .O(gate94inter10));
  nor2  gate614(.a(gate94inter10), .b(gate94inter9), .O(gate94inter11));
  nor2  gate615(.a(gate94inter11), .b(gate94inter6), .O(gate94inter12));
  nand2 gate616(.a(gate94inter12), .b(gate94inter1), .O(G415));

  xor2  gate2087(.a(G347), .b(G26), .O(gate95inter0));
  nand2 gate2088(.a(gate95inter0), .b(s_220), .O(gate95inter1));
  and2  gate2089(.a(G347), .b(G26), .O(gate95inter2));
  inv1  gate2090(.a(s_220), .O(gate95inter3));
  inv1  gate2091(.a(s_221), .O(gate95inter4));
  nand2 gate2092(.a(gate95inter4), .b(gate95inter3), .O(gate95inter5));
  nor2  gate2093(.a(gate95inter5), .b(gate95inter2), .O(gate95inter6));
  inv1  gate2094(.a(G26), .O(gate95inter7));
  inv1  gate2095(.a(G347), .O(gate95inter8));
  nand2 gate2096(.a(gate95inter8), .b(gate95inter7), .O(gate95inter9));
  nand2 gate2097(.a(s_221), .b(gate95inter3), .O(gate95inter10));
  nor2  gate2098(.a(gate95inter10), .b(gate95inter9), .O(gate95inter11));
  nor2  gate2099(.a(gate95inter11), .b(gate95inter6), .O(gate95inter12));
  nand2 gate2100(.a(gate95inter12), .b(gate95inter1), .O(G416));
nand2 gate96( .a(G30), .b(G347), .O(G417) );
nand2 gate97( .a(G19), .b(G350), .O(G418) );

  xor2  gate1121(.a(G350), .b(G23), .O(gate98inter0));
  nand2 gate1122(.a(gate98inter0), .b(s_82), .O(gate98inter1));
  and2  gate1123(.a(G350), .b(G23), .O(gate98inter2));
  inv1  gate1124(.a(s_82), .O(gate98inter3));
  inv1  gate1125(.a(s_83), .O(gate98inter4));
  nand2 gate1126(.a(gate98inter4), .b(gate98inter3), .O(gate98inter5));
  nor2  gate1127(.a(gate98inter5), .b(gate98inter2), .O(gate98inter6));
  inv1  gate1128(.a(G23), .O(gate98inter7));
  inv1  gate1129(.a(G350), .O(gate98inter8));
  nand2 gate1130(.a(gate98inter8), .b(gate98inter7), .O(gate98inter9));
  nand2 gate1131(.a(s_83), .b(gate98inter3), .O(gate98inter10));
  nor2  gate1132(.a(gate98inter10), .b(gate98inter9), .O(gate98inter11));
  nor2  gate1133(.a(gate98inter11), .b(gate98inter6), .O(gate98inter12));
  nand2 gate1134(.a(gate98inter12), .b(gate98inter1), .O(G419));
nand2 gate99( .a(G27), .b(G353), .O(G420) );
nand2 gate100( .a(G31), .b(G353), .O(G421) );

  xor2  gate2423(.a(G356), .b(G20), .O(gate101inter0));
  nand2 gate2424(.a(gate101inter0), .b(s_268), .O(gate101inter1));
  and2  gate2425(.a(G356), .b(G20), .O(gate101inter2));
  inv1  gate2426(.a(s_268), .O(gate101inter3));
  inv1  gate2427(.a(s_269), .O(gate101inter4));
  nand2 gate2428(.a(gate101inter4), .b(gate101inter3), .O(gate101inter5));
  nor2  gate2429(.a(gate101inter5), .b(gate101inter2), .O(gate101inter6));
  inv1  gate2430(.a(G20), .O(gate101inter7));
  inv1  gate2431(.a(G356), .O(gate101inter8));
  nand2 gate2432(.a(gate101inter8), .b(gate101inter7), .O(gate101inter9));
  nand2 gate2433(.a(s_269), .b(gate101inter3), .O(gate101inter10));
  nor2  gate2434(.a(gate101inter10), .b(gate101inter9), .O(gate101inter11));
  nor2  gate2435(.a(gate101inter11), .b(gate101inter6), .O(gate101inter12));
  nand2 gate2436(.a(gate101inter12), .b(gate101inter1), .O(G422));
nand2 gate102( .a(G24), .b(G356), .O(G423) );
nand2 gate103( .a(G28), .b(G359), .O(G424) );
nand2 gate104( .a(G32), .b(G359), .O(G425) );
nand2 gate105( .a(G362), .b(G363), .O(G426) );
nand2 gate106( .a(G364), .b(G365), .O(G429) );

  xor2  gate1513(.a(G367), .b(G366), .O(gate107inter0));
  nand2 gate1514(.a(gate107inter0), .b(s_138), .O(gate107inter1));
  and2  gate1515(.a(G367), .b(G366), .O(gate107inter2));
  inv1  gate1516(.a(s_138), .O(gate107inter3));
  inv1  gate1517(.a(s_139), .O(gate107inter4));
  nand2 gate1518(.a(gate107inter4), .b(gate107inter3), .O(gate107inter5));
  nor2  gate1519(.a(gate107inter5), .b(gate107inter2), .O(gate107inter6));
  inv1  gate1520(.a(G366), .O(gate107inter7));
  inv1  gate1521(.a(G367), .O(gate107inter8));
  nand2 gate1522(.a(gate107inter8), .b(gate107inter7), .O(gate107inter9));
  nand2 gate1523(.a(s_139), .b(gate107inter3), .O(gate107inter10));
  nor2  gate1524(.a(gate107inter10), .b(gate107inter9), .O(gate107inter11));
  nor2  gate1525(.a(gate107inter11), .b(gate107inter6), .O(gate107inter12));
  nand2 gate1526(.a(gate107inter12), .b(gate107inter1), .O(G432));

  xor2  gate1527(.a(G369), .b(G368), .O(gate108inter0));
  nand2 gate1528(.a(gate108inter0), .b(s_140), .O(gate108inter1));
  and2  gate1529(.a(G369), .b(G368), .O(gate108inter2));
  inv1  gate1530(.a(s_140), .O(gate108inter3));
  inv1  gate1531(.a(s_141), .O(gate108inter4));
  nand2 gate1532(.a(gate108inter4), .b(gate108inter3), .O(gate108inter5));
  nor2  gate1533(.a(gate108inter5), .b(gate108inter2), .O(gate108inter6));
  inv1  gate1534(.a(G368), .O(gate108inter7));
  inv1  gate1535(.a(G369), .O(gate108inter8));
  nand2 gate1536(.a(gate108inter8), .b(gate108inter7), .O(gate108inter9));
  nand2 gate1537(.a(s_141), .b(gate108inter3), .O(gate108inter10));
  nor2  gate1538(.a(gate108inter10), .b(gate108inter9), .O(gate108inter11));
  nor2  gate1539(.a(gate108inter11), .b(gate108inter6), .O(gate108inter12));
  nand2 gate1540(.a(gate108inter12), .b(gate108inter1), .O(G435));

  xor2  gate1555(.a(G371), .b(G370), .O(gate109inter0));
  nand2 gate1556(.a(gate109inter0), .b(s_144), .O(gate109inter1));
  and2  gate1557(.a(G371), .b(G370), .O(gate109inter2));
  inv1  gate1558(.a(s_144), .O(gate109inter3));
  inv1  gate1559(.a(s_145), .O(gate109inter4));
  nand2 gate1560(.a(gate109inter4), .b(gate109inter3), .O(gate109inter5));
  nor2  gate1561(.a(gate109inter5), .b(gate109inter2), .O(gate109inter6));
  inv1  gate1562(.a(G370), .O(gate109inter7));
  inv1  gate1563(.a(G371), .O(gate109inter8));
  nand2 gate1564(.a(gate109inter8), .b(gate109inter7), .O(gate109inter9));
  nand2 gate1565(.a(s_145), .b(gate109inter3), .O(gate109inter10));
  nor2  gate1566(.a(gate109inter10), .b(gate109inter9), .O(gate109inter11));
  nor2  gate1567(.a(gate109inter11), .b(gate109inter6), .O(gate109inter12));
  nand2 gate1568(.a(gate109inter12), .b(gate109inter1), .O(G438));
nand2 gate110( .a(G372), .b(G373), .O(G441) );
nand2 gate111( .a(G374), .b(G375), .O(G444) );
nand2 gate112( .a(G376), .b(G377), .O(G447) );

  xor2  gate1751(.a(G379), .b(G378), .O(gate113inter0));
  nand2 gate1752(.a(gate113inter0), .b(s_172), .O(gate113inter1));
  and2  gate1753(.a(G379), .b(G378), .O(gate113inter2));
  inv1  gate1754(.a(s_172), .O(gate113inter3));
  inv1  gate1755(.a(s_173), .O(gate113inter4));
  nand2 gate1756(.a(gate113inter4), .b(gate113inter3), .O(gate113inter5));
  nor2  gate1757(.a(gate113inter5), .b(gate113inter2), .O(gate113inter6));
  inv1  gate1758(.a(G378), .O(gate113inter7));
  inv1  gate1759(.a(G379), .O(gate113inter8));
  nand2 gate1760(.a(gate113inter8), .b(gate113inter7), .O(gate113inter9));
  nand2 gate1761(.a(s_173), .b(gate113inter3), .O(gate113inter10));
  nor2  gate1762(.a(gate113inter10), .b(gate113inter9), .O(gate113inter11));
  nor2  gate1763(.a(gate113inter11), .b(gate113inter6), .O(gate113inter12));
  nand2 gate1764(.a(gate113inter12), .b(gate113inter1), .O(G450));

  xor2  gate2563(.a(G381), .b(G380), .O(gate114inter0));
  nand2 gate2564(.a(gate114inter0), .b(s_288), .O(gate114inter1));
  and2  gate2565(.a(G381), .b(G380), .O(gate114inter2));
  inv1  gate2566(.a(s_288), .O(gate114inter3));
  inv1  gate2567(.a(s_289), .O(gate114inter4));
  nand2 gate2568(.a(gate114inter4), .b(gate114inter3), .O(gate114inter5));
  nor2  gate2569(.a(gate114inter5), .b(gate114inter2), .O(gate114inter6));
  inv1  gate2570(.a(G380), .O(gate114inter7));
  inv1  gate2571(.a(G381), .O(gate114inter8));
  nand2 gate2572(.a(gate114inter8), .b(gate114inter7), .O(gate114inter9));
  nand2 gate2573(.a(s_289), .b(gate114inter3), .O(gate114inter10));
  nor2  gate2574(.a(gate114inter10), .b(gate114inter9), .O(gate114inter11));
  nor2  gate2575(.a(gate114inter11), .b(gate114inter6), .O(gate114inter12));
  nand2 gate2576(.a(gate114inter12), .b(gate114inter1), .O(G453));
nand2 gate115( .a(G382), .b(G383), .O(G456) );
nand2 gate116( .a(G384), .b(G385), .O(G459) );
nand2 gate117( .a(G386), .b(G387), .O(G462) );

  xor2  gate799(.a(G389), .b(G388), .O(gate118inter0));
  nand2 gate800(.a(gate118inter0), .b(s_36), .O(gate118inter1));
  and2  gate801(.a(G389), .b(G388), .O(gate118inter2));
  inv1  gate802(.a(s_36), .O(gate118inter3));
  inv1  gate803(.a(s_37), .O(gate118inter4));
  nand2 gate804(.a(gate118inter4), .b(gate118inter3), .O(gate118inter5));
  nor2  gate805(.a(gate118inter5), .b(gate118inter2), .O(gate118inter6));
  inv1  gate806(.a(G388), .O(gate118inter7));
  inv1  gate807(.a(G389), .O(gate118inter8));
  nand2 gate808(.a(gate118inter8), .b(gate118inter7), .O(gate118inter9));
  nand2 gate809(.a(s_37), .b(gate118inter3), .O(gate118inter10));
  nor2  gate810(.a(gate118inter10), .b(gate118inter9), .O(gate118inter11));
  nor2  gate811(.a(gate118inter11), .b(gate118inter6), .O(gate118inter12));
  nand2 gate812(.a(gate118inter12), .b(gate118inter1), .O(G465));

  xor2  gate2381(.a(G391), .b(G390), .O(gate119inter0));
  nand2 gate2382(.a(gate119inter0), .b(s_262), .O(gate119inter1));
  and2  gate2383(.a(G391), .b(G390), .O(gate119inter2));
  inv1  gate2384(.a(s_262), .O(gate119inter3));
  inv1  gate2385(.a(s_263), .O(gate119inter4));
  nand2 gate2386(.a(gate119inter4), .b(gate119inter3), .O(gate119inter5));
  nor2  gate2387(.a(gate119inter5), .b(gate119inter2), .O(gate119inter6));
  inv1  gate2388(.a(G390), .O(gate119inter7));
  inv1  gate2389(.a(G391), .O(gate119inter8));
  nand2 gate2390(.a(gate119inter8), .b(gate119inter7), .O(gate119inter9));
  nand2 gate2391(.a(s_263), .b(gate119inter3), .O(gate119inter10));
  nor2  gate2392(.a(gate119inter10), .b(gate119inter9), .O(gate119inter11));
  nor2  gate2393(.a(gate119inter11), .b(gate119inter6), .O(gate119inter12));
  nand2 gate2394(.a(gate119inter12), .b(gate119inter1), .O(G468));
nand2 gate120( .a(G392), .b(G393), .O(G471) );
nand2 gate121( .a(G394), .b(G395), .O(G474) );

  xor2  gate939(.a(G397), .b(G396), .O(gate122inter0));
  nand2 gate940(.a(gate122inter0), .b(s_56), .O(gate122inter1));
  and2  gate941(.a(G397), .b(G396), .O(gate122inter2));
  inv1  gate942(.a(s_56), .O(gate122inter3));
  inv1  gate943(.a(s_57), .O(gate122inter4));
  nand2 gate944(.a(gate122inter4), .b(gate122inter3), .O(gate122inter5));
  nor2  gate945(.a(gate122inter5), .b(gate122inter2), .O(gate122inter6));
  inv1  gate946(.a(G396), .O(gate122inter7));
  inv1  gate947(.a(G397), .O(gate122inter8));
  nand2 gate948(.a(gate122inter8), .b(gate122inter7), .O(gate122inter9));
  nand2 gate949(.a(s_57), .b(gate122inter3), .O(gate122inter10));
  nor2  gate950(.a(gate122inter10), .b(gate122inter9), .O(gate122inter11));
  nor2  gate951(.a(gate122inter11), .b(gate122inter6), .O(gate122inter12));
  nand2 gate952(.a(gate122inter12), .b(gate122inter1), .O(G477));
nand2 gate123( .a(G398), .b(G399), .O(G480) );
nand2 gate124( .a(G400), .b(G401), .O(G483) );

  xor2  gate1289(.a(G403), .b(G402), .O(gate125inter0));
  nand2 gate1290(.a(gate125inter0), .b(s_106), .O(gate125inter1));
  and2  gate1291(.a(G403), .b(G402), .O(gate125inter2));
  inv1  gate1292(.a(s_106), .O(gate125inter3));
  inv1  gate1293(.a(s_107), .O(gate125inter4));
  nand2 gate1294(.a(gate125inter4), .b(gate125inter3), .O(gate125inter5));
  nor2  gate1295(.a(gate125inter5), .b(gate125inter2), .O(gate125inter6));
  inv1  gate1296(.a(G402), .O(gate125inter7));
  inv1  gate1297(.a(G403), .O(gate125inter8));
  nand2 gate1298(.a(gate125inter8), .b(gate125inter7), .O(gate125inter9));
  nand2 gate1299(.a(s_107), .b(gate125inter3), .O(gate125inter10));
  nor2  gate1300(.a(gate125inter10), .b(gate125inter9), .O(gate125inter11));
  nor2  gate1301(.a(gate125inter11), .b(gate125inter6), .O(gate125inter12));
  nand2 gate1302(.a(gate125inter12), .b(gate125inter1), .O(G486));
nand2 gate126( .a(G404), .b(G405), .O(G489) );
nand2 gate127( .a(G406), .b(G407), .O(G492) );
nand2 gate128( .a(G408), .b(G409), .O(G495) );

  xor2  gate659(.a(G411), .b(G410), .O(gate129inter0));
  nand2 gate660(.a(gate129inter0), .b(s_16), .O(gate129inter1));
  and2  gate661(.a(G411), .b(G410), .O(gate129inter2));
  inv1  gate662(.a(s_16), .O(gate129inter3));
  inv1  gate663(.a(s_17), .O(gate129inter4));
  nand2 gate664(.a(gate129inter4), .b(gate129inter3), .O(gate129inter5));
  nor2  gate665(.a(gate129inter5), .b(gate129inter2), .O(gate129inter6));
  inv1  gate666(.a(G410), .O(gate129inter7));
  inv1  gate667(.a(G411), .O(gate129inter8));
  nand2 gate668(.a(gate129inter8), .b(gate129inter7), .O(gate129inter9));
  nand2 gate669(.a(s_17), .b(gate129inter3), .O(gate129inter10));
  nor2  gate670(.a(gate129inter10), .b(gate129inter9), .O(gate129inter11));
  nor2  gate671(.a(gate129inter11), .b(gate129inter6), .O(gate129inter12));
  nand2 gate672(.a(gate129inter12), .b(gate129inter1), .O(G498));

  xor2  gate2017(.a(G413), .b(G412), .O(gate130inter0));
  nand2 gate2018(.a(gate130inter0), .b(s_210), .O(gate130inter1));
  and2  gate2019(.a(G413), .b(G412), .O(gate130inter2));
  inv1  gate2020(.a(s_210), .O(gate130inter3));
  inv1  gate2021(.a(s_211), .O(gate130inter4));
  nand2 gate2022(.a(gate130inter4), .b(gate130inter3), .O(gate130inter5));
  nor2  gate2023(.a(gate130inter5), .b(gate130inter2), .O(gate130inter6));
  inv1  gate2024(.a(G412), .O(gate130inter7));
  inv1  gate2025(.a(G413), .O(gate130inter8));
  nand2 gate2026(.a(gate130inter8), .b(gate130inter7), .O(gate130inter9));
  nand2 gate2027(.a(s_211), .b(gate130inter3), .O(gate130inter10));
  nor2  gate2028(.a(gate130inter10), .b(gate130inter9), .O(gate130inter11));
  nor2  gate2029(.a(gate130inter11), .b(gate130inter6), .O(gate130inter12));
  nand2 gate2030(.a(gate130inter12), .b(gate130inter1), .O(G501));
nand2 gate131( .a(G414), .b(G415), .O(G504) );
nand2 gate132( .a(G416), .b(G417), .O(G507) );
nand2 gate133( .a(G418), .b(G419), .O(G510) );
nand2 gate134( .a(G420), .b(G421), .O(G513) );
nand2 gate135( .a(G422), .b(G423), .O(G516) );
nand2 gate136( .a(G424), .b(G425), .O(G519) );
nand2 gate137( .a(G426), .b(G429), .O(G522) );

  xor2  gate1919(.a(G435), .b(G432), .O(gate138inter0));
  nand2 gate1920(.a(gate138inter0), .b(s_196), .O(gate138inter1));
  and2  gate1921(.a(G435), .b(G432), .O(gate138inter2));
  inv1  gate1922(.a(s_196), .O(gate138inter3));
  inv1  gate1923(.a(s_197), .O(gate138inter4));
  nand2 gate1924(.a(gate138inter4), .b(gate138inter3), .O(gate138inter5));
  nor2  gate1925(.a(gate138inter5), .b(gate138inter2), .O(gate138inter6));
  inv1  gate1926(.a(G432), .O(gate138inter7));
  inv1  gate1927(.a(G435), .O(gate138inter8));
  nand2 gate1928(.a(gate138inter8), .b(gate138inter7), .O(gate138inter9));
  nand2 gate1929(.a(s_197), .b(gate138inter3), .O(gate138inter10));
  nor2  gate1930(.a(gate138inter10), .b(gate138inter9), .O(gate138inter11));
  nor2  gate1931(.a(gate138inter11), .b(gate138inter6), .O(gate138inter12));
  nand2 gate1932(.a(gate138inter12), .b(gate138inter1), .O(G525));

  xor2  gate2703(.a(G441), .b(G438), .O(gate139inter0));
  nand2 gate2704(.a(gate139inter0), .b(s_308), .O(gate139inter1));
  and2  gate2705(.a(G441), .b(G438), .O(gate139inter2));
  inv1  gate2706(.a(s_308), .O(gate139inter3));
  inv1  gate2707(.a(s_309), .O(gate139inter4));
  nand2 gate2708(.a(gate139inter4), .b(gate139inter3), .O(gate139inter5));
  nor2  gate2709(.a(gate139inter5), .b(gate139inter2), .O(gate139inter6));
  inv1  gate2710(.a(G438), .O(gate139inter7));
  inv1  gate2711(.a(G441), .O(gate139inter8));
  nand2 gate2712(.a(gate139inter8), .b(gate139inter7), .O(gate139inter9));
  nand2 gate2713(.a(s_309), .b(gate139inter3), .O(gate139inter10));
  nor2  gate2714(.a(gate139inter10), .b(gate139inter9), .O(gate139inter11));
  nor2  gate2715(.a(gate139inter11), .b(gate139inter6), .O(gate139inter12));
  nand2 gate2716(.a(gate139inter12), .b(gate139inter1), .O(G528));
nand2 gate140( .a(G444), .b(G447), .O(G531) );
nand2 gate141( .a(G450), .b(G453), .O(G534) );

  xor2  gate1457(.a(G459), .b(G456), .O(gate142inter0));
  nand2 gate1458(.a(gate142inter0), .b(s_130), .O(gate142inter1));
  and2  gate1459(.a(G459), .b(G456), .O(gate142inter2));
  inv1  gate1460(.a(s_130), .O(gate142inter3));
  inv1  gate1461(.a(s_131), .O(gate142inter4));
  nand2 gate1462(.a(gate142inter4), .b(gate142inter3), .O(gate142inter5));
  nor2  gate1463(.a(gate142inter5), .b(gate142inter2), .O(gate142inter6));
  inv1  gate1464(.a(G456), .O(gate142inter7));
  inv1  gate1465(.a(G459), .O(gate142inter8));
  nand2 gate1466(.a(gate142inter8), .b(gate142inter7), .O(gate142inter9));
  nand2 gate1467(.a(s_131), .b(gate142inter3), .O(gate142inter10));
  nor2  gate1468(.a(gate142inter10), .b(gate142inter9), .O(gate142inter11));
  nor2  gate1469(.a(gate142inter11), .b(gate142inter6), .O(gate142inter12));
  nand2 gate1470(.a(gate142inter12), .b(gate142inter1), .O(G537));
nand2 gate143( .a(G462), .b(G465), .O(G540) );
nand2 gate144( .a(G468), .b(G471), .O(G543) );
nand2 gate145( .a(G474), .b(G477), .O(G546) );

  xor2  gate2115(.a(G483), .b(G480), .O(gate146inter0));
  nand2 gate2116(.a(gate146inter0), .b(s_224), .O(gate146inter1));
  and2  gate2117(.a(G483), .b(G480), .O(gate146inter2));
  inv1  gate2118(.a(s_224), .O(gate146inter3));
  inv1  gate2119(.a(s_225), .O(gate146inter4));
  nand2 gate2120(.a(gate146inter4), .b(gate146inter3), .O(gate146inter5));
  nor2  gate2121(.a(gate146inter5), .b(gate146inter2), .O(gate146inter6));
  inv1  gate2122(.a(G480), .O(gate146inter7));
  inv1  gate2123(.a(G483), .O(gate146inter8));
  nand2 gate2124(.a(gate146inter8), .b(gate146inter7), .O(gate146inter9));
  nand2 gate2125(.a(s_225), .b(gate146inter3), .O(gate146inter10));
  nor2  gate2126(.a(gate146inter10), .b(gate146inter9), .O(gate146inter11));
  nor2  gate2127(.a(gate146inter11), .b(gate146inter6), .O(gate146inter12));
  nand2 gate2128(.a(gate146inter12), .b(gate146inter1), .O(G549));
nand2 gate147( .a(G486), .b(G489), .O(G552) );

  xor2  gate1373(.a(G495), .b(G492), .O(gate148inter0));
  nand2 gate1374(.a(gate148inter0), .b(s_118), .O(gate148inter1));
  and2  gate1375(.a(G495), .b(G492), .O(gate148inter2));
  inv1  gate1376(.a(s_118), .O(gate148inter3));
  inv1  gate1377(.a(s_119), .O(gate148inter4));
  nand2 gate1378(.a(gate148inter4), .b(gate148inter3), .O(gate148inter5));
  nor2  gate1379(.a(gate148inter5), .b(gate148inter2), .O(gate148inter6));
  inv1  gate1380(.a(G492), .O(gate148inter7));
  inv1  gate1381(.a(G495), .O(gate148inter8));
  nand2 gate1382(.a(gate148inter8), .b(gate148inter7), .O(gate148inter9));
  nand2 gate1383(.a(s_119), .b(gate148inter3), .O(gate148inter10));
  nor2  gate1384(.a(gate148inter10), .b(gate148inter9), .O(gate148inter11));
  nor2  gate1385(.a(gate148inter11), .b(gate148inter6), .O(gate148inter12));
  nand2 gate1386(.a(gate148inter12), .b(gate148inter1), .O(G555));

  xor2  gate2227(.a(G501), .b(G498), .O(gate149inter0));
  nand2 gate2228(.a(gate149inter0), .b(s_240), .O(gate149inter1));
  and2  gate2229(.a(G501), .b(G498), .O(gate149inter2));
  inv1  gate2230(.a(s_240), .O(gate149inter3));
  inv1  gate2231(.a(s_241), .O(gate149inter4));
  nand2 gate2232(.a(gate149inter4), .b(gate149inter3), .O(gate149inter5));
  nor2  gate2233(.a(gate149inter5), .b(gate149inter2), .O(gate149inter6));
  inv1  gate2234(.a(G498), .O(gate149inter7));
  inv1  gate2235(.a(G501), .O(gate149inter8));
  nand2 gate2236(.a(gate149inter8), .b(gate149inter7), .O(gate149inter9));
  nand2 gate2237(.a(s_241), .b(gate149inter3), .O(gate149inter10));
  nor2  gate2238(.a(gate149inter10), .b(gate149inter9), .O(gate149inter11));
  nor2  gate2239(.a(gate149inter11), .b(gate149inter6), .O(gate149inter12));
  nand2 gate2240(.a(gate149inter12), .b(gate149inter1), .O(G558));
nand2 gate150( .a(G504), .b(G507), .O(G561) );
nand2 gate151( .a(G510), .b(G513), .O(G564) );

  xor2  gate1541(.a(G519), .b(G516), .O(gate152inter0));
  nand2 gate1542(.a(gate152inter0), .b(s_142), .O(gate152inter1));
  and2  gate1543(.a(G519), .b(G516), .O(gate152inter2));
  inv1  gate1544(.a(s_142), .O(gate152inter3));
  inv1  gate1545(.a(s_143), .O(gate152inter4));
  nand2 gate1546(.a(gate152inter4), .b(gate152inter3), .O(gate152inter5));
  nor2  gate1547(.a(gate152inter5), .b(gate152inter2), .O(gate152inter6));
  inv1  gate1548(.a(G516), .O(gate152inter7));
  inv1  gate1549(.a(G519), .O(gate152inter8));
  nand2 gate1550(.a(gate152inter8), .b(gate152inter7), .O(gate152inter9));
  nand2 gate1551(.a(s_143), .b(gate152inter3), .O(gate152inter10));
  nor2  gate1552(.a(gate152inter10), .b(gate152inter9), .O(gate152inter11));
  nor2  gate1553(.a(gate152inter11), .b(gate152inter6), .O(gate152inter12));
  nand2 gate1554(.a(gate152inter12), .b(gate152inter1), .O(G567));
nand2 gate153( .a(G426), .b(G522), .O(G570) );

  xor2  gate1079(.a(G522), .b(G429), .O(gate154inter0));
  nand2 gate1080(.a(gate154inter0), .b(s_76), .O(gate154inter1));
  and2  gate1081(.a(G522), .b(G429), .O(gate154inter2));
  inv1  gate1082(.a(s_76), .O(gate154inter3));
  inv1  gate1083(.a(s_77), .O(gate154inter4));
  nand2 gate1084(.a(gate154inter4), .b(gate154inter3), .O(gate154inter5));
  nor2  gate1085(.a(gate154inter5), .b(gate154inter2), .O(gate154inter6));
  inv1  gate1086(.a(G429), .O(gate154inter7));
  inv1  gate1087(.a(G522), .O(gate154inter8));
  nand2 gate1088(.a(gate154inter8), .b(gate154inter7), .O(gate154inter9));
  nand2 gate1089(.a(s_77), .b(gate154inter3), .O(gate154inter10));
  nor2  gate1090(.a(gate154inter10), .b(gate154inter9), .O(gate154inter11));
  nor2  gate1091(.a(gate154inter11), .b(gate154inter6), .O(gate154inter12));
  nand2 gate1092(.a(gate154inter12), .b(gate154inter1), .O(G571));
nand2 gate155( .a(G432), .b(G525), .O(G572) );

  xor2  gate2101(.a(G525), .b(G435), .O(gate156inter0));
  nand2 gate2102(.a(gate156inter0), .b(s_222), .O(gate156inter1));
  and2  gate2103(.a(G525), .b(G435), .O(gate156inter2));
  inv1  gate2104(.a(s_222), .O(gate156inter3));
  inv1  gate2105(.a(s_223), .O(gate156inter4));
  nand2 gate2106(.a(gate156inter4), .b(gate156inter3), .O(gate156inter5));
  nor2  gate2107(.a(gate156inter5), .b(gate156inter2), .O(gate156inter6));
  inv1  gate2108(.a(G435), .O(gate156inter7));
  inv1  gate2109(.a(G525), .O(gate156inter8));
  nand2 gate2110(.a(gate156inter8), .b(gate156inter7), .O(gate156inter9));
  nand2 gate2111(.a(s_223), .b(gate156inter3), .O(gate156inter10));
  nor2  gate2112(.a(gate156inter10), .b(gate156inter9), .O(gate156inter11));
  nor2  gate2113(.a(gate156inter11), .b(gate156inter6), .O(gate156inter12));
  nand2 gate2114(.a(gate156inter12), .b(gate156inter1), .O(G573));
nand2 gate157( .a(G438), .b(G528), .O(G574) );

  xor2  gate617(.a(G528), .b(G441), .O(gate158inter0));
  nand2 gate618(.a(gate158inter0), .b(s_10), .O(gate158inter1));
  and2  gate619(.a(G528), .b(G441), .O(gate158inter2));
  inv1  gate620(.a(s_10), .O(gate158inter3));
  inv1  gate621(.a(s_11), .O(gate158inter4));
  nand2 gate622(.a(gate158inter4), .b(gate158inter3), .O(gate158inter5));
  nor2  gate623(.a(gate158inter5), .b(gate158inter2), .O(gate158inter6));
  inv1  gate624(.a(G441), .O(gate158inter7));
  inv1  gate625(.a(G528), .O(gate158inter8));
  nand2 gate626(.a(gate158inter8), .b(gate158inter7), .O(gate158inter9));
  nand2 gate627(.a(s_11), .b(gate158inter3), .O(gate158inter10));
  nor2  gate628(.a(gate158inter10), .b(gate158inter9), .O(gate158inter11));
  nor2  gate629(.a(gate158inter11), .b(gate158inter6), .O(gate158inter12));
  nand2 gate630(.a(gate158inter12), .b(gate158inter1), .O(G575));

  xor2  gate561(.a(G531), .b(G444), .O(gate159inter0));
  nand2 gate562(.a(gate159inter0), .b(s_2), .O(gate159inter1));
  and2  gate563(.a(G531), .b(G444), .O(gate159inter2));
  inv1  gate564(.a(s_2), .O(gate159inter3));
  inv1  gate565(.a(s_3), .O(gate159inter4));
  nand2 gate566(.a(gate159inter4), .b(gate159inter3), .O(gate159inter5));
  nor2  gate567(.a(gate159inter5), .b(gate159inter2), .O(gate159inter6));
  inv1  gate568(.a(G444), .O(gate159inter7));
  inv1  gate569(.a(G531), .O(gate159inter8));
  nand2 gate570(.a(gate159inter8), .b(gate159inter7), .O(gate159inter9));
  nand2 gate571(.a(s_3), .b(gate159inter3), .O(gate159inter10));
  nor2  gate572(.a(gate159inter10), .b(gate159inter9), .O(gate159inter11));
  nor2  gate573(.a(gate159inter11), .b(gate159inter6), .O(gate159inter12));
  nand2 gate574(.a(gate159inter12), .b(gate159inter1), .O(G576));
nand2 gate160( .a(G447), .b(G531), .O(G577) );

  xor2  gate3137(.a(G534), .b(G450), .O(gate161inter0));
  nand2 gate3138(.a(gate161inter0), .b(s_370), .O(gate161inter1));
  and2  gate3139(.a(G534), .b(G450), .O(gate161inter2));
  inv1  gate3140(.a(s_370), .O(gate161inter3));
  inv1  gate3141(.a(s_371), .O(gate161inter4));
  nand2 gate3142(.a(gate161inter4), .b(gate161inter3), .O(gate161inter5));
  nor2  gate3143(.a(gate161inter5), .b(gate161inter2), .O(gate161inter6));
  inv1  gate3144(.a(G450), .O(gate161inter7));
  inv1  gate3145(.a(G534), .O(gate161inter8));
  nand2 gate3146(.a(gate161inter8), .b(gate161inter7), .O(gate161inter9));
  nand2 gate3147(.a(s_371), .b(gate161inter3), .O(gate161inter10));
  nor2  gate3148(.a(gate161inter10), .b(gate161inter9), .O(gate161inter11));
  nor2  gate3149(.a(gate161inter11), .b(gate161inter6), .O(gate161inter12));
  nand2 gate3150(.a(gate161inter12), .b(gate161inter1), .O(G578));
nand2 gate162( .a(G453), .b(G534), .O(G579) );
nand2 gate163( .a(G456), .b(G537), .O(G580) );
nand2 gate164( .a(G459), .b(G537), .O(G581) );
nand2 gate165( .a(G462), .b(G540), .O(G582) );
nand2 gate166( .a(G465), .b(G540), .O(G583) );
nand2 gate167( .a(G468), .b(G543), .O(G584) );
nand2 gate168( .a(G471), .b(G543), .O(G585) );

  xor2  gate3109(.a(G546), .b(G474), .O(gate169inter0));
  nand2 gate3110(.a(gate169inter0), .b(s_366), .O(gate169inter1));
  and2  gate3111(.a(G546), .b(G474), .O(gate169inter2));
  inv1  gate3112(.a(s_366), .O(gate169inter3));
  inv1  gate3113(.a(s_367), .O(gate169inter4));
  nand2 gate3114(.a(gate169inter4), .b(gate169inter3), .O(gate169inter5));
  nor2  gate3115(.a(gate169inter5), .b(gate169inter2), .O(gate169inter6));
  inv1  gate3116(.a(G474), .O(gate169inter7));
  inv1  gate3117(.a(G546), .O(gate169inter8));
  nand2 gate3118(.a(gate169inter8), .b(gate169inter7), .O(gate169inter9));
  nand2 gate3119(.a(s_367), .b(gate169inter3), .O(gate169inter10));
  nor2  gate3120(.a(gate169inter10), .b(gate169inter9), .O(gate169inter11));
  nor2  gate3121(.a(gate169inter11), .b(gate169inter6), .O(gate169inter12));
  nand2 gate3122(.a(gate169inter12), .b(gate169inter1), .O(G586));

  xor2  gate1905(.a(G546), .b(G477), .O(gate170inter0));
  nand2 gate1906(.a(gate170inter0), .b(s_194), .O(gate170inter1));
  and2  gate1907(.a(G546), .b(G477), .O(gate170inter2));
  inv1  gate1908(.a(s_194), .O(gate170inter3));
  inv1  gate1909(.a(s_195), .O(gate170inter4));
  nand2 gate1910(.a(gate170inter4), .b(gate170inter3), .O(gate170inter5));
  nor2  gate1911(.a(gate170inter5), .b(gate170inter2), .O(gate170inter6));
  inv1  gate1912(.a(G477), .O(gate170inter7));
  inv1  gate1913(.a(G546), .O(gate170inter8));
  nand2 gate1914(.a(gate170inter8), .b(gate170inter7), .O(gate170inter9));
  nand2 gate1915(.a(s_195), .b(gate170inter3), .O(gate170inter10));
  nor2  gate1916(.a(gate170inter10), .b(gate170inter9), .O(gate170inter11));
  nor2  gate1917(.a(gate170inter11), .b(gate170inter6), .O(gate170inter12));
  nand2 gate1918(.a(gate170inter12), .b(gate170inter1), .O(G587));
nand2 gate171( .a(G480), .b(G549), .O(G588) );
nand2 gate172( .a(G483), .b(G549), .O(G589) );
nand2 gate173( .a(G486), .b(G552), .O(G590) );
nand2 gate174( .a(G489), .b(G552), .O(G591) );

  xor2  gate2451(.a(G555), .b(G492), .O(gate175inter0));
  nand2 gate2452(.a(gate175inter0), .b(s_272), .O(gate175inter1));
  and2  gate2453(.a(G555), .b(G492), .O(gate175inter2));
  inv1  gate2454(.a(s_272), .O(gate175inter3));
  inv1  gate2455(.a(s_273), .O(gate175inter4));
  nand2 gate2456(.a(gate175inter4), .b(gate175inter3), .O(gate175inter5));
  nor2  gate2457(.a(gate175inter5), .b(gate175inter2), .O(gate175inter6));
  inv1  gate2458(.a(G492), .O(gate175inter7));
  inv1  gate2459(.a(G555), .O(gate175inter8));
  nand2 gate2460(.a(gate175inter8), .b(gate175inter7), .O(gate175inter9));
  nand2 gate2461(.a(s_273), .b(gate175inter3), .O(gate175inter10));
  nor2  gate2462(.a(gate175inter10), .b(gate175inter9), .O(gate175inter11));
  nor2  gate2463(.a(gate175inter11), .b(gate175inter6), .O(gate175inter12));
  nand2 gate2464(.a(gate175inter12), .b(gate175inter1), .O(G592));
nand2 gate176( .a(G495), .b(G555), .O(G593) );
nand2 gate177( .a(G498), .b(G558), .O(G594) );

  xor2  gate2773(.a(G558), .b(G501), .O(gate178inter0));
  nand2 gate2774(.a(gate178inter0), .b(s_318), .O(gate178inter1));
  and2  gate2775(.a(G558), .b(G501), .O(gate178inter2));
  inv1  gate2776(.a(s_318), .O(gate178inter3));
  inv1  gate2777(.a(s_319), .O(gate178inter4));
  nand2 gate2778(.a(gate178inter4), .b(gate178inter3), .O(gate178inter5));
  nor2  gate2779(.a(gate178inter5), .b(gate178inter2), .O(gate178inter6));
  inv1  gate2780(.a(G501), .O(gate178inter7));
  inv1  gate2781(.a(G558), .O(gate178inter8));
  nand2 gate2782(.a(gate178inter8), .b(gate178inter7), .O(gate178inter9));
  nand2 gate2783(.a(s_319), .b(gate178inter3), .O(gate178inter10));
  nor2  gate2784(.a(gate178inter10), .b(gate178inter9), .O(gate178inter11));
  nor2  gate2785(.a(gate178inter11), .b(gate178inter6), .O(gate178inter12));
  nand2 gate2786(.a(gate178inter12), .b(gate178inter1), .O(G595));

  xor2  gate1051(.a(G561), .b(G504), .O(gate179inter0));
  nand2 gate1052(.a(gate179inter0), .b(s_72), .O(gate179inter1));
  and2  gate1053(.a(G561), .b(G504), .O(gate179inter2));
  inv1  gate1054(.a(s_72), .O(gate179inter3));
  inv1  gate1055(.a(s_73), .O(gate179inter4));
  nand2 gate1056(.a(gate179inter4), .b(gate179inter3), .O(gate179inter5));
  nor2  gate1057(.a(gate179inter5), .b(gate179inter2), .O(gate179inter6));
  inv1  gate1058(.a(G504), .O(gate179inter7));
  inv1  gate1059(.a(G561), .O(gate179inter8));
  nand2 gate1060(.a(gate179inter8), .b(gate179inter7), .O(gate179inter9));
  nand2 gate1061(.a(s_73), .b(gate179inter3), .O(gate179inter10));
  nor2  gate1062(.a(gate179inter10), .b(gate179inter9), .O(gate179inter11));
  nor2  gate1063(.a(gate179inter11), .b(gate179inter6), .O(gate179inter12));
  nand2 gate1064(.a(gate179inter12), .b(gate179inter1), .O(G596));

  xor2  gate2633(.a(G561), .b(G507), .O(gate180inter0));
  nand2 gate2634(.a(gate180inter0), .b(s_298), .O(gate180inter1));
  and2  gate2635(.a(G561), .b(G507), .O(gate180inter2));
  inv1  gate2636(.a(s_298), .O(gate180inter3));
  inv1  gate2637(.a(s_299), .O(gate180inter4));
  nand2 gate2638(.a(gate180inter4), .b(gate180inter3), .O(gate180inter5));
  nor2  gate2639(.a(gate180inter5), .b(gate180inter2), .O(gate180inter6));
  inv1  gate2640(.a(G507), .O(gate180inter7));
  inv1  gate2641(.a(G561), .O(gate180inter8));
  nand2 gate2642(.a(gate180inter8), .b(gate180inter7), .O(gate180inter9));
  nand2 gate2643(.a(s_299), .b(gate180inter3), .O(gate180inter10));
  nor2  gate2644(.a(gate180inter10), .b(gate180inter9), .O(gate180inter11));
  nor2  gate2645(.a(gate180inter11), .b(gate180inter6), .O(gate180inter12));
  nand2 gate2646(.a(gate180inter12), .b(gate180inter1), .O(G597));

  xor2  gate2997(.a(G564), .b(G510), .O(gate181inter0));
  nand2 gate2998(.a(gate181inter0), .b(s_350), .O(gate181inter1));
  and2  gate2999(.a(G564), .b(G510), .O(gate181inter2));
  inv1  gate3000(.a(s_350), .O(gate181inter3));
  inv1  gate3001(.a(s_351), .O(gate181inter4));
  nand2 gate3002(.a(gate181inter4), .b(gate181inter3), .O(gate181inter5));
  nor2  gate3003(.a(gate181inter5), .b(gate181inter2), .O(gate181inter6));
  inv1  gate3004(.a(G510), .O(gate181inter7));
  inv1  gate3005(.a(G564), .O(gate181inter8));
  nand2 gate3006(.a(gate181inter8), .b(gate181inter7), .O(gate181inter9));
  nand2 gate3007(.a(s_351), .b(gate181inter3), .O(gate181inter10));
  nor2  gate3008(.a(gate181inter10), .b(gate181inter9), .O(gate181inter11));
  nor2  gate3009(.a(gate181inter11), .b(gate181inter6), .O(gate181inter12));
  nand2 gate3010(.a(gate181inter12), .b(gate181inter1), .O(G598));
nand2 gate182( .a(G513), .b(G564), .O(G599) );

  xor2  gate1191(.a(G567), .b(G516), .O(gate183inter0));
  nand2 gate1192(.a(gate183inter0), .b(s_92), .O(gate183inter1));
  and2  gate1193(.a(G567), .b(G516), .O(gate183inter2));
  inv1  gate1194(.a(s_92), .O(gate183inter3));
  inv1  gate1195(.a(s_93), .O(gate183inter4));
  nand2 gate1196(.a(gate183inter4), .b(gate183inter3), .O(gate183inter5));
  nor2  gate1197(.a(gate183inter5), .b(gate183inter2), .O(gate183inter6));
  inv1  gate1198(.a(G516), .O(gate183inter7));
  inv1  gate1199(.a(G567), .O(gate183inter8));
  nand2 gate1200(.a(gate183inter8), .b(gate183inter7), .O(gate183inter9));
  nand2 gate1201(.a(s_93), .b(gate183inter3), .O(gate183inter10));
  nor2  gate1202(.a(gate183inter10), .b(gate183inter9), .O(gate183inter11));
  nor2  gate1203(.a(gate183inter11), .b(gate183inter6), .O(gate183inter12));
  nand2 gate1204(.a(gate183inter12), .b(gate183inter1), .O(G600));
nand2 gate184( .a(G519), .b(G567), .O(G601) );
nand2 gate185( .a(G570), .b(G571), .O(G602) );
nand2 gate186( .a(G572), .b(G573), .O(G607) );

  xor2  gate2297(.a(G575), .b(G574), .O(gate187inter0));
  nand2 gate2298(.a(gate187inter0), .b(s_250), .O(gate187inter1));
  and2  gate2299(.a(G575), .b(G574), .O(gate187inter2));
  inv1  gate2300(.a(s_250), .O(gate187inter3));
  inv1  gate2301(.a(s_251), .O(gate187inter4));
  nand2 gate2302(.a(gate187inter4), .b(gate187inter3), .O(gate187inter5));
  nor2  gate2303(.a(gate187inter5), .b(gate187inter2), .O(gate187inter6));
  inv1  gate2304(.a(G574), .O(gate187inter7));
  inv1  gate2305(.a(G575), .O(gate187inter8));
  nand2 gate2306(.a(gate187inter8), .b(gate187inter7), .O(gate187inter9));
  nand2 gate2307(.a(s_251), .b(gate187inter3), .O(gate187inter10));
  nor2  gate2308(.a(gate187inter10), .b(gate187inter9), .O(gate187inter11));
  nor2  gate2309(.a(gate187inter11), .b(gate187inter6), .O(gate187inter12));
  nand2 gate2310(.a(gate187inter12), .b(gate187inter1), .O(G612));
nand2 gate188( .a(G576), .b(G577), .O(G617) );
nand2 gate189( .a(G578), .b(G579), .O(G622) );

  xor2  gate3081(.a(G581), .b(G580), .O(gate190inter0));
  nand2 gate3082(.a(gate190inter0), .b(s_362), .O(gate190inter1));
  and2  gate3083(.a(G581), .b(G580), .O(gate190inter2));
  inv1  gate3084(.a(s_362), .O(gate190inter3));
  inv1  gate3085(.a(s_363), .O(gate190inter4));
  nand2 gate3086(.a(gate190inter4), .b(gate190inter3), .O(gate190inter5));
  nor2  gate3087(.a(gate190inter5), .b(gate190inter2), .O(gate190inter6));
  inv1  gate3088(.a(G580), .O(gate190inter7));
  inv1  gate3089(.a(G581), .O(gate190inter8));
  nand2 gate3090(.a(gate190inter8), .b(gate190inter7), .O(gate190inter9));
  nand2 gate3091(.a(s_363), .b(gate190inter3), .O(gate190inter10));
  nor2  gate3092(.a(gate190inter10), .b(gate190inter9), .O(gate190inter11));
  nor2  gate3093(.a(gate190inter11), .b(gate190inter6), .O(gate190inter12));
  nand2 gate3094(.a(gate190inter12), .b(gate190inter1), .O(G627));
nand2 gate191( .a(G582), .b(G583), .O(G632) );

  xor2  gate2969(.a(G585), .b(G584), .O(gate192inter0));
  nand2 gate2970(.a(gate192inter0), .b(s_346), .O(gate192inter1));
  and2  gate2971(.a(G585), .b(G584), .O(gate192inter2));
  inv1  gate2972(.a(s_346), .O(gate192inter3));
  inv1  gate2973(.a(s_347), .O(gate192inter4));
  nand2 gate2974(.a(gate192inter4), .b(gate192inter3), .O(gate192inter5));
  nor2  gate2975(.a(gate192inter5), .b(gate192inter2), .O(gate192inter6));
  inv1  gate2976(.a(G584), .O(gate192inter7));
  inv1  gate2977(.a(G585), .O(gate192inter8));
  nand2 gate2978(.a(gate192inter8), .b(gate192inter7), .O(gate192inter9));
  nand2 gate2979(.a(s_347), .b(gate192inter3), .O(gate192inter10));
  nor2  gate2980(.a(gate192inter10), .b(gate192inter9), .O(gate192inter11));
  nor2  gate2981(.a(gate192inter11), .b(gate192inter6), .O(gate192inter12));
  nand2 gate2982(.a(gate192inter12), .b(gate192inter1), .O(G637));
nand2 gate193( .a(G586), .b(G587), .O(G642) );

  xor2  gate2675(.a(G589), .b(G588), .O(gate194inter0));
  nand2 gate2676(.a(gate194inter0), .b(s_304), .O(gate194inter1));
  and2  gate2677(.a(G589), .b(G588), .O(gate194inter2));
  inv1  gate2678(.a(s_304), .O(gate194inter3));
  inv1  gate2679(.a(s_305), .O(gate194inter4));
  nand2 gate2680(.a(gate194inter4), .b(gate194inter3), .O(gate194inter5));
  nor2  gate2681(.a(gate194inter5), .b(gate194inter2), .O(gate194inter6));
  inv1  gate2682(.a(G588), .O(gate194inter7));
  inv1  gate2683(.a(G589), .O(gate194inter8));
  nand2 gate2684(.a(gate194inter8), .b(gate194inter7), .O(gate194inter9));
  nand2 gate2685(.a(s_305), .b(gate194inter3), .O(gate194inter10));
  nor2  gate2686(.a(gate194inter10), .b(gate194inter9), .O(gate194inter11));
  nor2  gate2687(.a(gate194inter11), .b(gate194inter6), .O(gate194inter12));
  nand2 gate2688(.a(gate194inter12), .b(gate194inter1), .O(G645));

  xor2  gate2521(.a(G591), .b(G590), .O(gate195inter0));
  nand2 gate2522(.a(gate195inter0), .b(s_282), .O(gate195inter1));
  and2  gate2523(.a(G591), .b(G590), .O(gate195inter2));
  inv1  gate2524(.a(s_282), .O(gate195inter3));
  inv1  gate2525(.a(s_283), .O(gate195inter4));
  nand2 gate2526(.a(gate195inter4), .b(gate195inter3), .O(gate195inter5));
  nor2  gate2527(.a(gate195inter5), .b(gate195inter2), .O(gate195inter6));
  inv1  gate2528(.a(G590), .O(gate195inter7));
  inv1  gate2529(.a(G591), .O(gate195inter8));
  nand2 gate2530(.a(gate195inter8), .b(gate195inter7), .O(gate195inter9));
  nand2 gate2531(.a(s_283), .b(gate195inter3), .O(gate195inter10));
  nor2  gate2532(.a(gate195inter10), .b(gate195inter9), .O(gate195inter11));
  nor2  gate2533(.a(gate195inter11), .b(gate195inter6), .O(gate195inter12));
  nand2 gate2534(.a(gate195inter12), .b(gate195inter1), .O(G648));

  xor2  gate1807(.a(G593), .b(G592), .O(gate196inter0));
  nand2 gate1808(.a(gate196inter0), .b(s_180), .O(gate196inter1));
  and2  gate1809(.a(G593), .b(G592), .O(gate196inter2));
  inv1  gate1810(.a(s_180), .O(gate196inter3));
  inv1  gate1811(.a(s_181), .O(gate196inter4));
  nand2 gate1812(.a(gate196inter4), .b(gate196inter3), .O(gate196inter5));
  nor2  gate1813(.a(gate196inter5), .b(gate196inter2), .O(gate196inter6));
  inv1  gate1814(.a(G592), .O(gate196inter7));
  inv1  gate1815(.a(G593), .O(gate196inter8));
  nand2 gate1816(.a(gate196inter8), .b(gate196inter7), .O(gate196inter9));
  nand2 gate1817(.a(s_181), .b(gate196inter3), .O(gate196inter10));
  nor2  gate1818(.a(gate196inter10), .b(gate196inter9), .O(gate196inter11));
  nor2  gate1819(.a(gate196inter11), .b(gate196inter6), .O(gate196inter12));
  nand2 gate1820(.a(gate196inter12), .b(gate196inter1), .O(G651));

  xor2  gate883(.a(G595), .b(G594), .O(gate197inter0));
  nand2 gate884(.a(gate197inter0), .b(s_48), .O(gate197inter1));
  and2  gate885(.a(G595), .b(G594), .O(gate197inter2));
  inv1  gate886(.a(s_48), .O(gate197inter3));
  inv1  gate887(.a(s_49), .O(gate197inter4));
  nand2 gate888(.a(gate197inter4), .b(gate197inter3), .O(gate197inter5));
  nor2  gate889(.a(gate197inter5), .b(gate197inter2), .O(gate197inter6));
  inv1  gate890(.a(G594), .O(gate197inter7));
  inv1  gate891(.a(G595), .O(gate197inter8));
  nand2 gate892(.a(gate197inter8), .b(gate197inter7), .O(gate197inter9));
  nand2 gate893(.a(s_49), .b(gate197inter3), .O(gate197inter10));
  nor2  gate894(.a(gate197inter10), .b(gate197inter9), .O(gate197inter11));
  nor2  gate895(.a(gate197inter11), .b(gate197inter6), .O(gate197inter12));
  nand2 gate896(.a(gate197inter12), .b(gate197inter1), .O(G654));
nand2 gate198( .a(G596), .b(G597), .O(G657) );
nand2 gate199( .a(G598), .b(G599), .O(G660) );

  xor2  gate981(.a(G601), .b(G600), .O(gate200inter0));
  nand2 gate982(.a(gate200inter0), .b(s_62), .O(gate200inter1));
  and2  gate983(.a(G601), .b(G600), .O(gate200inter2));
  inv1  gate984(.a(s_62), .O(gate200inter3));
  inv1  gate985(.a(s_63), .O(gate200inter4));
  nand2 gate986(.a(gate200inter4), .b(gate200inter3), .O(gate200inter5));
  nor2  gate987(.a(gate200inter5), .b(gate200inter2), .O(gate200inter6));
  inv1  gate988(.a(G600), .O(gate200inter7));
  inv1  gate989(.a(G601), .O(gate200inter8));
  nand2 gate990(.a(gate200inter8), .b(gate200inter7), .O(gate200inter9));
  nand2 gate991(.a(s_63), .b(gate200inter3), .O(gate200inter10));
  nor2  gate992(.a(gate200inter10), .b(gate200inter9), .O(gate200inter11));
  nor2  gate993(.a(gate200inter11), .b(gate200inter6), .O(gate200inter12));
  nand2 gate994(.a(gate200inter12), .b(gate200inter1), .O(G663));

  xor2  gate1709(.a(G607), .b(G602), .O(gate201inter0));
  nand2 gate1710(.a(gate201inter0), .b(s_166), .O(gate201inter1));
  and2  gate1711(.a(G607), .b(G602), .O(gate201inter2));
  inv1  gate1712(.a(s_166), .O(gate201inter3));
  inv1  gate1713(.a(s_167), .O(gate201inter4));
  nand2 gate1714(.a(gate201inter4), .b(gate201inter3), .O(gate201inter5));
  nor2  gate1715(.a(gate201inter5), .b(gate201inter2), .O(gate201inter6));
  inv1  gate1716(.a(G602), .O(gate201inter7));
  inv1  gate1717(.a(G607), .O(gate201inter8));
  nand2 gate1718(.a(gate201inter8), .b(gate201inter7), .O(gate201inter9));
  nand2 gate1719(.a(s_167), .b(gate201inter3), .O(gate201inter10));
  nor2  gate1720(.a(gate201inter10), .b(gate201inter9), .O(gate201inter11));
  nor2  gate1721(.a(gate201inter11), .b(gate201inter6), .O(gate201inter12));
  nand2 gate1722(.a(gate201inter12), .b(gate201inter1), .O(G666));
nand2 gate202( .a(G612), .b(G617), .O(G669) );

  xor2  gate673(.a(G612), .b(G602), .O(gate203inter0));
  nand2 gate674(.a(gate203inter0), .b(s_18), .O(gate203inter1));
  and2  gate675(.a(G612), .b(G602), .O(gate203inter2));
  inv1  gate676(.a(s_18), .O(gate203inter3));
  inv1  gate677(.a(s_19), .O(gate203inter4));
  nand2 gate678(.a(gate203inter4), .b(gate203inter3), .O(gate203inter5));
  nor2  gate679(.a(gate203inter5), .b(gate203inter2), .O(gate203inter6));
  inv1  gate680(.a(G602), .O(gate203inter7));
  inv1  gate681(.a(G612), .O(gate203inter8));
  nand2 gate682(.a(gate203inter8), .b(gate203inter7), .O(gate203inter9));
  nand2 gate683(.a(s_19), .b(gate203inter3), .O(gate203inter10));
  nor2  gate684(.a(gate203inter10), .b(gate203inter9), .O(gate203inter11));
  nor2  gate685(.a(gate203inter11), .b(gate203inter6), .O(gate203inter12));
  nand2 gate686(.a(gate203inter12), .b(gate203inter1), .O(G672));
nand2 gate204( .a(G607), .b(G617), .O(G675) );

  xor2  gate2857(.a(G627), .b(G622), .O(gate205inter0));
  nand2 gate2858(.a(gate205inter0), .b(s_330), .O(gate205inter1));
  and2  gate2859(.a(G627), .b(G622), .O(gate205inter2));
  inv1  gate2860(.a(s_330), .O(gate205inter3));
  inv1  gate2861(.a(s_331), .O(gate205inter4));
  nand2 gate2862(.a(gate205inter4), .b(gate205inter3), .O(gate205inter5));
  nor2  gate2863(.a(gate205inter5), .b(gate205inter2), .O(gate205inter6));
  inv1  gate2864(.a(G622), .O(gate205inter7));
  inv1  gate2865(.a(G627), .O(gate205inter8));
  nand2 gate2866(.a(gate205inter8), .b(gate205inter7), .O(gate205inter9));
  nand2 gate2867(.a(s_331), .b(gate205inter3), .O(gate205inter10));
  nor2  gate2868(.a(gate205inter10), .b(gate205inter9), .O(gate205inter11));
  nor2  gate2869(.a(gate205inter11), .b(gate205inter6), .O(gate205inter12));
  nand2 gate2870(.a(gate205inter12), .b(gate205inter1), .O(G678));

  xor2  gate813(.a(G637), .b(G632), .O(gate206inter0));
  nand2 gate814(.a(gate206inter0), .b(s_38), .O(gate206inter1));
  and2  gate815(.a(G637), .b(G632), .O(gate206inter2));
  inv1  gate816(.a(s_38), .O(gate206inter3));
  inv1  gate817(.a(s_39), .O(gate206inter4));
  nand2 gate818(.a(gate206inter4), .b(gate206inter3), .O(gate206inter5));
  nor2  gate819(.a(gate206inter5), .b(gate206inter2), .O(gate206inter6));
  inv1  gate820(.a(G632), .O(gate206inter7));
  inv1  gate821(.a(G637), .O(gate206inter8));
  nand2 gate822(.a(gate206inter8), .b(gate206inter7), .O(gate206inter9));
  nand2 gate823(.a(s_39), .b(gate206inter3), .O(gate206inter10));
  nor2  gate824(.a(gate206inter10), .b(gate206inter9), .O(gate206inter11));
  nor2  gate825(.a(gate206inter11), .b(gate206inter6), .O(gate206inter12));
  nand2 gate826(.a(gate206inter12), .b(gate206inter1), .O(G681));

  xor2  gate575(.a(G632), .b(G622), .O(gate207inter0));
  nand2 gate576(.a(gate207inter0), .b(s_4), .O(gate207inter1));
  and2  gate577(.a(G632), .b(G622), .O(gate207inter2));
  inv1  gate578(.a(s_4), .O(gate207inter3));
  inv1  gate579(.a(s_5), .O(gate207inter4));
  nand2 gate580(.a(gate207inter4), .b(gate207inter3), .O(gate207inter5));
  nor2  gate581(.a(gate207inter5), .b(gate207inter2), .O(gate207inter6));
  inv1  gate582(.a(G622), .O(gate207inter7));
  inv1  gate583(.a(G632), .O(gate207inter8));
  nand2 gate584(.a(gate207inter8), .b(gate207inter7), .O(gate207inter9));
  nand2 gate585(.a(s_5), .b(gate207inter3), .O(gate207inter10));
  nor2  gate586(.a(gate207inter10), .b(gate207inter9), .O(gate207inter11));
  nor2  gate587(.a(gate207inter11), .b(gate207inter6), .O(gate207inter12));
  nand2 gate588(.a(gate207inter12), .b(gate207inter1), .O(G684));
nand2 gate208( .a(G627), .b(G637), .O(G687) );
nand2 gate209( .a(G602), .b(G666), .O(G690) );

  xor2  gate771(.a(G666), .b(G607), .O(gate210inter0));
  nand2 gate772(.a(gate210inter0), .b(s_32), .O(gate210inter1));
  and2  gate773(.a(G666), .b(G607), .O(gate210inter2));
  inv1  gate774(.a(s_32), .O(gate210inter3));
  inv1  gate775(.a(s_33), .O(gate210inter4));
  nand2 gate776(.a(gate210inter4), .b(gate210inter3), .O(gate210inter5));
  nor2  gate777(.a(gate210inter5), .b(gate210inter2), .O(gate210inter6));
  inv1  gate778(.a(G607), .O(gate210inter7));
  inv1  gate779(.a(G666), .O(gate210inter8));
  nand2 gate780(.a(gate210inter8), .b(gate210inter7), .O(gate210inter9));
  nand2 gate781(.a(s_33), .b(gate210inter3), .O(gate210inter10));
  nor2  gate782(.a(gate210inter10), .b(gate210inter9), .O(gate210inter11));
  nor2  gate783(.a(gate210inter11), .b(gate210inter6), .O(gate210inter12));
  nand2 gate784(.a(gate210inter12), .b(gate210inter1), .O(G691));

  xor2  gate743(.a(G669), .b(G612), .O(gate211inter0));
  nand2 gate744(.a(gate211inter0), .b(s_28), .O(gate211inter1));
  and2  gate745(.a(G669), .b(G612), .O(gate211inter2));
  inv1  gate746(.a(s_28), .O(gate211inter3));
  inv1  gate747(.a(s_29), .O(gate211inter4));
  nand2 gate748(.a(gate211inter4), .b(gate211inter3), .O(gate211inter5));
  nor2  gate749(.a(gate211inter5), .b(gate211inter2), .O(gate211inter6));
  inv1  gate750(.a(G612), .O(gate211inter7));
  inv1  gate751(.a(G669), .O(gate211inter8));
  nand2 gate752(.a(gate211inter8), .b(gate211inter7), .O(gate211inter9));
  nand2 gate753(.a(s_29), .b(gate211inter3), .O(gate211inter10));
  nor2  gate754(.a(gate211inter10), .b(gate211inter9), .O(gate211inter11));
  nor2  gate755(.a(gate211inter11), .b(gate211inter6), .O(gate211inter12));
  nand2 gate756(.a(gate211inter12), .b(gate211inter1), .O(G692));
nand2 gate212( .a(G617), .b(G669), .O(G693) );

  xor2  gate2493(.a(G672), .b(G602), .O(gate213inter0));
  nand2 gate2494(.a(gate213inter0), .b(s_278), .O(gate213inter1));
  and2  gate2495(.a(G672), .b(G602), .O(gate213inter2));
  inv1  gate2496(.a(s_278), .O(gate213inter3));
  inv1  gate2497(.a(s_279), .O(gate213inter4));
  nand2 gate2498(.a(gate213inter4), .b(gate213inter3), .O(gate213inter5));
  nor2  gate2499(.a(gate213inter5), .b(gate213inter2), .O(gate213inter6));
  inv1  gate2500(.a(G602), .O(gate213inter7));
  inv1  gate2501(.a(G672), .O(gate213inter8));
  nand2 gate2502(.a(gate213inter8), .b(gate213inter7), .O(gate213inter9));
  nand2 gate2503(.a(s_279), .b(gate213inter3), .O(gate213inter10));
  nor2  gate2504(.a(gate213inter10), .b(gate213inter9), .O(gate213inter11));
  nor2  gate2505(.a(gate213inter11), .b(gate213inter6), .O(gate213inter12));
  nand2 gate2506(.a(gate213inter12), .b(gate213inter1), .O(G694));

  xor2  gate2213(.a(G672), .b(G612), .O(gate214inter0));
  nand2 gate2214(.a(gate214inter0), .b(s_238), .O(gate214inter1));
  and2  gate2215(.a(G672), .b(G612), .O(gate214inter2));
  inv1  gate2216(.a(s_238), .O(gate214inter3));
  inv1  gate2217(.a(s_239), .O(gate214inter4));
  nand2 gate2218(.a(gate214inter4), .b(gate214inter3), .O(gate214inter5));
  nor2  gate2219(.a(gate214inter5), .b(gate214inter2), .O(gate214inter6));
  inv1  gate2220(.a(G612), .O(gate214inter7));
  inv1  gate2221(.a(G672), .O(gate214inter8));
  nand2 gate2222(.a(gate214inter8), .b(gate214inter7), .O(gate214inter9));
  nand2 gate2223(.a(s_239), .b(gate214inter3), .O(gate214inter10));
  nor2  gate2224(.a(gate214inter10), .b(gate214inter9), .O(gate214inter11));
  nor2  gate2225(.a(gate214inter11), .b(gate214inter6), .O(gate214inter12));
  nand2 gate2226(.a(gate214inter12), .b(gate214inter1), .O(G695));
nand2 gate215( .a(G607), .b(G675), .O(G696) );
nand2 gate216( .a(G617), .b(G675), .O(G697) );

  xor2  gate1233(.a(G678), .b(G622), .O(gate217inter0));
  nand2 gate1234(.a(gate217inter0), .b(s_98), .O(gate217inter1));
  and2  gate1235(.a(G678), .b(G622), .O(gate217inter2));
  inv1  gate1236(.a(s_98), .O(gate217inter3));
  inv1  gate1237(.a(s_99), .O(gate217inter4));
  nand2 gate1238(.a(gate217inter4), .b(gate217inter3), .O(gate217inter5));
  nor2  gate1239(.a(gate217inter5), .b(gate217inter2), .O(gate217inter6));
  inv1  gate1240(.a(G622), .O(gate217inter7));
  inv1  gate1241(.a(G678), .O(gate217inter8));
  nand2 gate1242(.a(gate217inter8), .b(gate217inter7), .O(gate217inter9));
  nand2 gate1243(.a(s_99), .b(gate217inter3), .O(gate217inter10));
  nor2  gate1244(.a(gate217inter10), .b(gate217inter9), .O(gate217inter11));
  nor2  gate1245(.a(gate217inter11), .b(gate217inter6), .O(gate217inter12));
  nand2 gate1246(.a(gate217inter12), .b(gate217inter1), .O(G698));
nand2 gate218( .a(G627), .b(G678), .O(G699) );
nand2 gate219( .a(G632), .b(G681), .O(G700) );

  xor2  gate3123(.a(G681), .b(G637), .O(gate220inter0));
  nand2 gate3124(.a(gate220inter0), .b(s_368), .O(gate220inter1));
  and2  gate3125(.a(G681), .b(G637), .O(gate220inter2));
  inv1  gate3126(.a(s_368), .O(gate220inter3));
  inv1  gate3127(.a(s_369), .O(gate220inter4));
  nand2 gate3128(.a(gate220inter4), .b(gate220inter3), .O(gate220inter5));
  nor2  gate3129(.a(gate220inter5), .b(gate220inter2), .O(gate220inter6));
  inv1  gate3130(.a(G637), .O(gate220inter7));
  inv1  gate3131(.a(G681), .O(gate220inter8));
  nand2 gate3132(.a(gate220inter8), .b(gate220inter7), .O(gate220inter9));
  nand2 gate3133(.a(s_369), .b(gate220inter3), .O(gate220inter10));
  nor2  gate3134(.a(gate220inter10), .b(gate220inter9), .O(gate220inter11));
  nor2  gate3135(.a(gate220inter11), .b(gate220inter6), .O(gate220inter12));
  nand2 gate3136(.a(gate220inter12), .b(gate220inter1), .O(G701));
nand2 gate221( .a(G622), .b(G684), .O(G702) );

  xor2  gate687(.a(G684), .b(G632), .O(gate222inter0));
  nand2 gate688(.a(gate222inter0), .b(s_20), .O(gate222inter1));
  and2  gate689(.a(G684), .b(G632), .O(gate222inter2));
  inv1  gate690(.a(s_20), .O(gate222inter3));
  inv1  gate691(.a(s_21), .O(gate222inter4));
  nand2 gate692(.a(gate222inter4), .b(gate222inter3), .O(gate222inter5));
  nor2  gate693(.a(gate222inter5), .b(gate222inter2), .O(gate222inter6));
  inv1  gate694(.a(G632), .O(gate222inter7));
  inv1  gate695(.a(G684), .O(gate222inter8));
  nand2 gate696(.a(gate222inter8), .b(gate222inter7), .O(gate222inter9));
  nand2 gate697(.a(s_21), .b(gate222inter3), .O(gate222inter10));
  nor2  gate698(.a(gate222inter10), .b(gate222inter9), .O(gate222inter11));
  nor2  gate699(.a(gate222inter11), .b(gate222inter6), .O(gate222inter12));
  nand2 gate700(.a(gate222inter12), .b(gate222inter1), .O(G703));
nand2 gate223( .a(G627), .b(G687), .O(G704) );
nand2 gate224( .a(G637), .b(G687), .O(G705) );

  xor2  gate2157(.a(G691), .b(G690), .O(gate225inter0));
  nand2 gate2158(.a(gate225inter0), .b(s_230), .O(gate225inter1));
  and2  gate2159(.a(G691), .b(G690), .O(gate225inter2));
  inv1  gate2160(.a(s_230), .O(gate225inter3));
  inv1  gate2161(.a(s_231), .O(gate225inter4));
  nand2 gate2162(.a(gate225inter4), .b(gate225inter3), .O(gate225inter5));
  nor2  gate2163(.a(gate225inter5), .b(gate225inter2), .O(gate225inter6));
  inv1  gate2164(.a(G690), .O(gate225inter7));
  inv1  gate2165(.a(G691), .O(gate225inter8));
  nand2 gate2166(.a(gate225inter8), .b(gate225inter7), .O(gate225inter9));
  nand2 gate2167(.a(s_231), .b(gate225inter3), .O(gate225inter10));
  nor2  gate2168(.a(gate225inter10), .b(gate225inter9), .O(gate225inter11));
  nor2  gate2169(.a(gate225inter11), .b(gate225inter6), .O(gate225inter12));
  nand2 gate2170(.a(gate225inter12), .b(gate225inter1), .O(G706));

  xor2  gate2045(.a(G693), .b(G692), .O(gate226inter0));
  nand2 gate2046(.a(gate226inter0), .b(s_214), .O(gate226inter1));
  and2  gate2047(.a(G693), .b(G692), .O(gate226inter2));
  inv1  gate2048(.a(s_214), .O(gate226inter3));
  inv1  gate2049(.a(s_215), .O(gate226inter4));
  nand2 gate2050(.a(gate226inter4), .b(gate226inter3), .O(gate226inter5));
  nor2  gate2051(.a(gate226inter5), .b(gate226inter2), .O(gate226inter6));
  inv1  gate2052(.a(G692), .O(gate226inter7));
  inv1  gate2053(.a(G693), .O(gate226inter8));
  nand2 gate2054(.a(gate226inter8), .b(gate226inter7), .O(gate226inter9));
  nand2 gate2055(.a(s_215), .b(gate226inter3), .O(gate226inter10));
  nor2  gate2056(.a(gate226inter10), .b(gate226inter9), .O(gate226inter11));
  nor2  gate2057(.a(gate226inter11), .b(gate226inter6), .O(gate226inter12));
  nand2 gate2058(.a(gate226inter12), .b(gate226inter1), .O(G709));
nand2 gate227( .a(G694), .b(G695), .O(G712) );
nand2 gate228( .a(G696), .b(G697), .O(G715) );
nand2 gate229( .a(G698), .b(G699), .O(G718) );

  xor2  gate2941(.a(G701), .b(G700), .O(gate230inter0));
  nand2 gate2942(.a(gate230inter0), .b(s_342), .O(gate230inter1));
  and2  gate2943(.a(G701), .b(G700), .O(gate230inter2));
  inv1  gate2944(.a(s_342), .O(gate230inter3));
  inv1  gate2945(.a(s_343), .O(gate230inter4));
  nand2 gate2946(.a(gate230inter4), .b(gate230inter3), .O(gate230inter5));
  nor2  gate2947(.a(gate230inter5), .b(gate230inter2), .O(gate230inter6));
  inv1  gate2948(.a(G700), .O(gate230inter7));
  inv1  gate2949(.a(G701), .O(gate230inter8));
  nand2 gate2950(.a(gate230inter8), .b(gate230inter7), .O(gate230inter9));
  nand2 gate2951(.a(s_343), .b(gate230inter3), .O(gate230inter10));
  nor2  gate2952(.a(gate230inter10), .b(gate230inter9), .O(gate230inter11));
  nor2  gate2953(.a(gate230inter11), .b(gate230inter6), .O(gate230inter12));
  nand2 gate2954(.a(gate230inter12), .b(gate230inter1), .O(G721));
nand2 gate231( .a(G702), .b(G703), .O(G724) );

  xor2  gate1737(.a(G705), .b(G704), .O(gate232inter0));
  nand2 gate1738(.a(gate232inter0), .b(s_170), .O(gate232inter1));
  and2  gate1739(.a(G705), .b(G704), .O(gate232inter2));
  inv1  gate1740(.a(s_170), .O(gate232inter3));
  inv1  gate1741(.a(s_171), .O(gate232inter4));
  nand2 gate1742(.a(gate232inter4), .b(gate232inter3), .O(gate232inter5));
  nor2  gate1743(.a(gate232inter5), .b(gate232inter2), .O(gate232inter6));
  inv1  gate1744(.a(G704), .O(gate232inter7));
  inv1  gate1745(.a(G705), .O(gate232inter8));
  nand2 gate1746(.a(gate232inter8), .b(gate232inter7), .O(gate232inter9));
  nand2 gate1747(.a(s_171), .b(gate232inter3), .O(gate232inter10));
  nor2  gate1748(.a(gate232inter10), .b(gate232inter9), .O(gate232inter11));
  nor2  gate1749(.a(gate232inter11), .b(gate232inter6), .O(gate232inter12));
  nand2 gate1750(.a(gate232inter12), .b(gate232inter1), .O(G727));

  xor2  gate2983(.a(G718), .b(G242), .O(gate233inter0));
  nand2 gate2984(.a(gate233inter0), .b(s_348), .O(gate233inter1));
  and2  gate2985(.a(G718), .b(G242), .O(gate233inter2));
  inv1  gate2986(.a(s_348), .O(gate233inter3));
  inv1  gate2987(.a(s_349), .O(gate233inter4));
  nand2 gate2988(.a(gate233inter4), .b(gate233inter3), .O(gate233inter5));
  nor2  gate2989(.a(gate233inter5), .b(gate233inter2), .O(gate233inter6));
  inv1  gate2990(.a(G242), .O(gate233inter7));
  inv1  gate2991(.a(G718), .O(gate233inter8));
  nand2 gate2992(.a(gate233inter8), .b(gate233inter7), .O(gate233inter9));
  nand2 gate2993(.a(s_349), .b(gate233inter3), .O(gate233inter10));
  nor2  gate2994(.a(gate233inter10), .b(gate233inter9), .O(gate233inter11));
  nor2  gate2995(.a(gate233inter11), .b(gate233inter6), .O(gate233inter12));
  nand2 gate2996(.a(gate233inter12), .b(gate233inter1), .O(G730));
nand2 gate234( .a(G245), .b(G721), .O(G733) );
nand2 gate235( .a(G248), .b(G724), .O(G736) );

  xor2  gate1723(.a(G727), .b(G251), .O(gate236inter0));
  nand2 gate1724(.a(gate236inter0), .b(s_168), .O(gate236inter1));
  and2  gate1725(.a(G727), .b(G251), .O(gate236inter2));
  inv1  gate1726(.a(s_168), .O(gate236inter3));
  inv1  gate1727(.a(s_169), .O(gate236inter4));
  nand2 gate1728(.a(gate236inter4), .b(gate236inter3), .O(gate236inter5));
  nor2  gate1729(.a(gate236inter5), .b(gate236inter2), .O(gate236inter6));
  inv1  gate1730(.a(G251), .O(gate236inter7));
  inv1  gate1731(.a(G727), .O(gate236inter8));
  nand2 gate1732(.a(gate236inter8), .b(gate236inter7), .O(gate236inter9));
  nand2 gate1733(.a(s_169), .b(gate236inter3), .O(gate236inter10));
  nor2  gate1734(.a(gate236inter10), .b(gate236inter9), .O(gate236inter11));
  nor2  gate1735(.a(gate236inter11), .b(gate236inter6), .O(gate236inter12));
  nand2 gate1736(.a(gate236inter12), .b(gate236inter1), .O(G739));
nand2 gate237( .a(G254), .b(G706), .O(G742) );
nand2 gate238( .a(G257), .b(G709), .O(G745) );
nand2 gate239( .a(G260), .b(G712), .O(G748) );

  xor2  gate827(.a(G715), .b(G263), .O(gate240inter0));
  nand2 gate828(.a(gate240inter0), .b(s_40), .O(gate240inter1));
  and2  gate829(.a(G715), .b(G263), .O(gate240inter2));
  inv1  gate830(.a(s_40), .O(gate240inter3));
  inv1  gate831(.a(s_41), .O(gate240inter4));
  nand2 gate832(.a(gate240inter4), .b(gate240inter3), .O(gate240inter5));
  nor2  gate833(.a(gate240inter5), .b(gate240inter2), .O(gate240inter6));
  inv1  gate834(.a(G263), .O(gate240inter7));
  inv1  gate835(.a(G715), .O(gate240inter8));
  nand2 gate836(.a(gate240inter8), .b(gate240inter7), .O(gate240inter9));
  nand2 gate837(.a(s_41), .b(gate240inter3), .O(gate240inter10));
  nor2  gate838(.a(gate240inter10), .b(gate240inter9), .O(gate240inter11));
  nor2  gate839(.a(gate240inter11), .b(gate240inter6), .O(gate240inter12));
  nand2 gate840(.a(gate240inter12), .b(gate240inter1), .O(G751));
nand2 gate241( .a(G242), .b(G730), .O(G754) );

  xor2  gate2661(.a(G730), .b(G718), .O(gate242inter0));
  nand2 gate2662(.a(gate242inter0), .b(s_302), .O(gate242inter1));
  and2  gate2663(.a(G730), .b(G718), .O(gate242inter2));
  inv1  gate2664(.a(s_302), .O(gate242inter3));
  inv1  gate2665(.a(s_303), .O(gate242inter4));
  nand2 gate2666(.a(gate242inter4), .b(gate242inter3), .O(gate242inter5));
  nor2  gate2667(.a(gate242inter5), .b(gate242inter2), .O(gate242inter6));
  inv1  gate2668(.a(G718), .O(gate242inter7));
  inv1  gate2669(.a(G730), .O(gate242inter8));
  nand2 gate2670(.a(gate242inter8), .b(gate242inter7), .O(gate242inter9));
  nand2 gate2671(.a(s_303), .b(gate242inter3), .O(gate242inter10));
  nor2  gate2672(.a(gate242inter10), .b(gate242inter9), .O(gate242inter11));
  nor2  gate2673(.a(gate242inter11), .b(gate242inter6), .O(gate242inter12));
  nand2 gate2674(.a(gate242inter12), .b(gate242inter1), .O(G755));

  xor2  gate967(.a(G733), .b(G245), .O(gate243inter0));
  nand2 gate968(.a(gate243inter0), .b(s_60), .O(gate243inter1));
  and2  gate969(.a(G733), .b(G245), .O(gate243inter2));
  inv1  gate970(.a(s_60), .O(gate243inter3));
  inv1  gate971(.a(s_61), .O(gate243inter4));
  nand2 gate972(.a(gate243inter4), .b(gate243inter3), .O(gate243inter5));
  nor2  gate973(.a(gate243inter5), .b(gate243inter2), .O(gate243inter6));
  inv1  gate974(.a(G245), .O(gate243inter7));
  inv1  gate975(.a(G733), .O(gate243inter8));
  nand2 gate976(.a(gate243inter8), .b(gate243inter7), .O(gate243inter9));
  nand2 gate977(.a(s_61), .b(gate243inter3), .O(gate243inter10));
  nor2  gate978(.a(gate243inter10), .b(gate243inter9), .O(gate243inter11));
  nor2  gate979(.a(gate243inter11), .b(gate243inter6), .O(gate243inter12));
  nand2 gate980(.a(gate243inter12), .b(gate243inter1), .O(G756));

  xor2  gate1639(.a(G733), .b(G721), .O(gate244inter0));
  nand2 gate1640(.a(gate244inter0), .b(s_156), .O(gate244inter1));
  and2  gate1641(.a(G733), .b(G721), .O(gate244inter2));
  inv1  gate1642(.a(s_156), .O(gate244inter3));
  inv1  gate1643(.a(s_157), .O(gate244inter4));
  nand2 gate1644(.a(gate244inter4), .b(gate244inter3), .O(gate244inter5));
  nor2  gate1645(.a(gate244inter5), .b(gate244inter2), .O(gate244inter6));
  inv1  gate1646(.a(G721), .O(gate244inter7));
  inv1  gate1647(.a(G733), .O(gate244inter8));
  nand2 gate1648(.a(gate244inter8), .b(gate244inter7), .O(gate244inter9));
  nand2 gate1649(.a(s_157), .b(gate244inter3), .O(gate244inter10));
  nor2  gate1650(.a(gate244inter10), .b(gate244inter9), .O(gate244inter11));
  nor2  gate1651(.a(gate244inter11), .b(gate244inter6), .O(gate244inter12));
  nand2 gate1652(.a(gate244inter12), .b(gate244inter1), .O(G757));

  xor2  gate1681(.a(G736), .b(G248), .O(gate245inter0));
  nand2 gate1682(.a(gate245inter0), .b(s_162), .O(gate245inter1));
  and2  gate1683(.a(G736), .b(G248), .O(gate245inter2));
  inv1  gate1684(.a(s_162), .O(gate245inter3));
  inv1  gate1685(.a(s_163), .O(gate245inter4));
  nand2 gate1686(.a(gate245inter4), .b(gate245inter3), .O(gate245inter5));
  nor2  gate1687(.a(gate245inter5), .b(gate245inter2), .O(gate245inter6));
  inv1  gate1688(.a(G248), .O(gate245inter7));
  inv1  gate1689(.a(G736), .O(gate245inter8));
  nand2 gate1690(.a(gate245inter8), .b(gate245inter7), .O(gate245inter9));
  nand2 gate1691(.a(s_163), .b(gate245inter3), .O(gate245inter10));
  nor2  gate1692(.a(gate245inter10), .b(gate245inter9), .O(gate245inter11));
  nor2  gate1693(.a(gate245inter11), .b(gate245inter6), .O(gate245inter12));
  nand2 gate1694(.a(gate245inter12), .b(gate245inter1), .O(G758));
nand2 gate246( .a(G724), .b(G736), .O(G759) );
nand2 gate247( .a(G251), .b(G739), .O(G760) );
nand2 gate248( .a(G727), .b(G739), .O(G761) );

  xor2  gate1499(.a(G742), .b(G254), .O(gate249inter0));
  nand2 gate1500(.a(gate249inter0), .b(s_136), .O(gate249inter1));
  and2  gate1501(.a(G742), .b(G254), .O(gate249inter2));
  inv1  gate1502(.a(s_136), .O(gate249inter3));
  inv1  gate1503(.a(s_137), .O(gate249inter4));
  nand2 gate1504(.a(gate249inter4), .b(gate249inter3), .O(gate249inter5));
  nor2  gate1505(.a(gate249inter5), .b(gate249inter2), .O(gate249inter6));
  inv1  gate1506(.a(G254), .O(gate249inter7));
  inv1  gate1507(.a(G742), .O(gate249inter8));
  nand2 gate1508(.a(gate249inter8), .b(gate249inter7), .O(gate249inter9));
  nand2 gate1509(.a(s_137), .b(gate249inter3), .O(gate249inter10));
  nor2  gate1510(.a(gate249inter10), .b(gate249inter9), .O(gate249inter11));
  nor2  gate1511(.a(gate249inter11), .b(gate249inter6), .O(gate249inter12));
  nand2 gate1512(.a(gate249inter12), .b(gate249inter1), .O(G762));

  xor2  gate2395(.a(G742), .b(G706), .O(gate250inter0));
  nand2 gate2396(.a(gate250inter0), .b(s_264), .O(gate250inter1));
  and2  gate2397(.a(G742), .b(G706), .O(gate250inter2));
  inv1  gate2398(.a(s_264), .O(gate250inter3));
  inv1  gate2399(.a(s_265), .O(gate250inter4));
  nand2 gate2400(.a(gate250inter4), .b(gate250inter3), .O(gate250inter5));
  nor2  gate2401(.a(gate250inter5), .b(gate250inter2), .O(gate250inter6));
  inv1  gate2402(.a(G706), .O(gate250inter7));
  inv1  gate2403(.a(G742), .O(gate250inter8));
  nand2 gate2404(.a(gate250inter8), .b(gate250inter7), .O(gate250inter9));
  nand2 gate2405(.a(s_265), .b(gate250inter3), .O(gate250inter10));
  nor2  gate2406(.a(gate250inter10), .b(gate250inter9), .O(gate250inter11));
  nor2  gate2407(.a(gate250inter11), .b(gate250inter6), .O(gate250inter12));
  nand2 gate2408(.a(gate250inter12), .b(gate250inter1), .O(G763));
nand2 gate251( .a(G257), .b(G745), .O(G764) );
nand2 gate252( .a(G709), .b(G745), .O(G765) );
nand2 gate253( .a(G260), .b(G748), .O(G766) );
nand2 gate254( .a(G712), .b(G748), .O(G767) );
nand2 gate255( .a(G263), .b(G751), .O(G768) );

  xor2  gate953(.a(G751), .b(G715), .O(gate256inter0));
  nand2 gate954(.a(gate256inter0), .b(s_58), .O(gate256inter1));
  and2  gate955(.a(G751), .b(G715), .O(gate256inter2));
  inv1  gate956(.a(s_58), .O(gate256inter3));
  inv1  gate957(.a(s_59), .O(gate256inter4));
  nand2 gate958(.a(gate256inter4), .b(gate256inter3), .O(gate256inter5));
  nor2  gate959(.a(gate256inter5), .b(gate256inter2), .O(gate256inter6));
  inv1  gate960(.a(G715), .O(gate256inter7));
  inv1  gate961(.a(G751), .O(gate256inter8));
  nand2 gate962(.a(gate256inter8), .b(gate256inter7), .O(gate256inter9));
  nand2 gate963(.a(s_59), .b(gate256inter3), .O(gate256inter10));
  nor2  gate964(.a(gate256inter10), .b(gate256inter9), .O(gate256inter11));
  nor2  gate965(.a(gate256inter11), .b(gate256inter6), .O(gate256inter12));
  nand2 gate966(.a(gate256inter12), .b(gate256inter1), .O(G769));
nand2 gate257( .a(G754), .b(G755), .O(G770) );

  xor2  gate2927(.a(G757), .b(G756), .O(gate258inter0));
  nand2 gate2928(.a(gate258inter0), .b(s_340), .O(gate258inter1));
  and2  gate2929(.a(G757), .b(G756), .O(gate258inter2));
  inv1  gate2930(.a(s_340), .O(gate258inter3));
  inv1  gate2931(.a(s_341), .O(gate258inter4));
  nand2 gate2932(.a(gate258inter4), .b(gate258inter3), .O(gate258inter5));
  nor2  gate2933(.a(gate258inter5), .b(gate258inter2), .O(gate258inter6));
  inv1  gate2934(.a(G756), .O(gate258inter7));
  inv1  gate2935(.a(G757), .O(gate258inter8));
  nand2 gate2936(.a(gate258inter8), .b(gate258inter7), .O(gate258inter9));
  nand2 gate2937(.a(s_341), .b(gate258inter3), .O(gate258inter10));
  nor2  gate2938(.a(gate258inter10), .b(gate258inter9), .O(gate258inter11));
  nor2  gate2939(.a(gate258inter11), .b(gate258inter6), .O(gate258inter12));
  nand2 gate2940(.a(gate258inter12), .b(gate258inter1), .O(G773));
nand2 gate259( .a(G758), .b(G759), .O(G776) );
nand2 gate260( .a(G760), .b(G761), .O(G779) );
nand2 gate261( .a(G762), .b(G763), .O(G782) );

  xor2  gate1779(.a(G765), .b(G764), .O(gate262inter0));
  nand2 gate1780(.a(gate262inter0), .b(s_176), .O(gate262inter1));
  and2  gate1781(.a(G765), .b(G764), .O(gate262inter2));
  inv1  gate1782(.a(s_176), .O(gate262inter3));
  inv1  gate1783(.a(s_177), .O(gate262inter4));
  nand2 gate1784(.a(gate262inter4), .b(gate262inter3), .O(gate262inter5));
  nor2  gate1785(.a(gate262inter5), .b(gate262inter2), .O(gate262inter6));
  inv1  gate1786(.a(G764), .O(gate262inter7));
  inv1  gate1787(.a(G765), .O(gate262inter8));
  nand2 gate1788(.a(gate262inter8), .b(gate262inter7), .O(gate262inter9));
  nand2 gate1789(.a(s_177), .b(gate262inter3), .O(gate262inter10));
  nor2  gate1790(.a(gate262inter10), .b(gate262inter9), .O(gate262inter11));
  nor2  gate1791(.a(gate262inter11), .b(gate262inter6), .O(gate262inter12));
  nand2 gate1792(.a(gate262inter12), .b(gate262inter1), .O(G785));
nand2 gate263( .a(G766), .b(G767), .O(G788) );
nand2 gate264( .a(G768), .b(G769), .O(G791) );

  xor2  gate1135(.a(G770), .b(G642), .O(gate265inter0));
  nand2 gate1136(.a(gate265inter0), .b(s_84), .O(gate265inter1));
  and2  gate1137(.a(G770), .b(G642), .O(gate265inter2));
  inv1  gate1138(.a(s_84), .O(gate265inter3));
  inv1  gate1139(.a(s_85), .O(gate265inter4));
  nand2 gate1140(.a(gate265inter4), .b(gate265inter3), .O(gate265inter5));
  nor2  gate1141(.a(gate265inter5), .b(gate265inter2), .O(gate265inter6));
  inv1  gate1142(.a(G642), .O(gate265inter7));
  inv1  gate1143(.a(G770), .O(gate265inter8));
  nand2 gate1144(.a(gate265inter8), .b(gate265inter7), .O(gate265inter9));
  nand2 gate1145(.a(s_85), .b(gate265inter3), .O(gate265inter10));
  nor2  gate1146(.a(gate265inter10), .b(gate265inter9), .O(gate265inter11));
  nor2  gate1147(.a(gate265inter11), .b(gate265inter6), .O(gate265inter12));
  nand2 gate1148(.a(gate265inter12), .b(gate265inter1), .O(G794));
nand2 gate266( .a(G645), .b(G773), .O(G797) );
nand2 gate267( .a(G648), .b(G776), .O(G800) );
nand2 gate268( .a(G651), .b(G779), .O(G803) );
nand2 gate269( .a(G654), .b(G782), .O(G806) );

  xor2  gate1009(.a(G785), .b(G657), .O(gate270inter0));
  nand2 gate1010(.a(gate270inter0), .b(s_66), .O(gate270inter1));
  and2  gate1011(.a(G785), .b(G657), .O(gate270inter2));
  inv1  gate1012(.a(s_66), .O(gate270inter3));
  inv1  gate1013(.a(s_67), .O(gate270inter4));
  nand2 gate1014(.a(gate270inter4), .b(gate270inter3), .O(gate270inter5));
  nor2  gate1015(.a(gate270inter5), .b(gate270inter2), .O(gate270inter6));
  inv1  gate1016(.a(G657), .O(gate270inter7));
  inv1  gate1017(.a(G785), .O(gate270inter8));
  nand2 gate1018(.a(gate270inter8), .b(gate270inter7), .O(gate270inter9));
  nand2 gate1019(.a(s_67), .b(gate270inter3), .O(gate270inter10));
  nor2  gate1020(.a(gate270inter10), .b(gate270inter9), .O(gate270inter11));
  nor2  gate1021(.a(gate270inter11), .b(gate270inter6), .O(gate270inter12));
  nand2 gate1022(.a(gate270inter12), .b(gate270inter1), .O(G809));
nand2 gate271( .a(G660), .b(G788), .O(G812) );
nand2 gate272( .a(G663), .b(G791), .O(G815) );
nand2 gate273( .a(G642), .b(G794), .O(G818) );

  xor2  gate1765(.a(G794), .b(G770), .O(gate274inter0));
  nand2 gate1766(.a(gate274inter0), .b(s_174), .O(gate274inter1));
  and2  gate1767(.a(G794), .b(G770), .O(gate274inter2));
  inv1  gate1768(.a(s_174), .O(gate274inter3));
  inv1  gate1769(.a(s_175), .O(gate274inter4));
  nand2 gate1770(.a(gate274inter4), .b(gate274inter3), .O(gate274inter5));
  nor2  gate1771(.a(gate274inter5), .b(gate274inter2), .O(gate274inter6));
  inv1  gate1772(.a(G770), .O(gate274inter7));
  inv1  gate1773(.a(G794), .O(gate274inter8));
  nand2 gate1774(.a(gate274inter8), .b(gate274inter7), .O(gate274inter9));
  nand2 gate1775(.a(s_175), .b(gate274inter3), .O(gate274inter10));
  nor2  gate1776(.a(gate274inter10), .b(gate274inter9), .O(gate274inter11));
  nor2  gate1777(.a(gate274inter11), .b(gate274inter6), .O(gate274inter12));
  nand2 gate1778(.a(gate274inter12), .b(gate274inter1), .O(G819));
nand2 gate275( .a(G645), .b(G797), .O(G820) );
nand2 gate276( .a(G773), .b(G797), .O(G821) );

  xor2  gate2759(.a(G800), .b(G648), .O(gate277inter0));
  nand2 gate2760(.a(gate277inter0), .b(s_316), .O(gate277inter1));
  and2  gate2761(.a(G800), .b(G648), .O(gate277inter2));
  inv1  gate2762(.a(s_316), .O(gate277inter3));
  inv1  gate2763(.a(s_317), .O(gate277inter4));
  nand2 gate2764(.a(gate277inter4), .b(gate277inter3), .O(gate277inter5));
  nor2  gate2765(.a(gate277inter5), .b(gate277inter2), .O(gate277inter6));
  inv1  gate2766(.a(G648), .O(gate277inter7));
  inv1  gate2767(.a(G800), .O(gate277inter8));
  nand2 gate2768(.a(gate277inter8), .b(gate277inter7), .O(gate277inter9));
  nand2 gate2769(.a(s_317), .b(gate277inter3), .O(gate277inter10));
  nor2  gate2770(.a(gate277inter10), .b(gate277inter9), .O(gate277inter11));
  nor2  gate2771(.a(gate277inter11), .b(gate277inter6), .O(gate277inter12));
  nand2 gate2772(.a(gate277inter12), .b(gate277inter1), .O(G822));

  xor2  gate925(.a(G800), .b(G776), .O(gate278inter0));
  nand2 gate926(.a(gate278inter0), .b(s_54), .O(gate278inter1));
  and2  gate927(.a(G800), .b(G776), .O(gate278inter2));
  inv1  gate928(.a(s_54), .O(gate278inter3));
  inv1  gate929(.a(s_55), .O(gate278inter4));
  nand2 gate930(.a(gate278inter4), .b(gate278inter3), .O(gate278inter5));
  nor2  gate931(.a(gate278inter5), .b(gate278inter2), .O(gate278inter6));
  inv1  gate932(.a(G776), .O(gate278inter7));
  inv1  gate933(.a(G800), .O(gate278inter8));
  nand2 gate934(.a(gate278inter8), .b(gate278inter7), .O(gate278inter9));
  nand2 gate935(.a(s_55), .b(gate278inter3), .O(gate278inter10));
  nor2  gate936(.a(gate278inter10), .b(gate278inter9), .O(gate278inter11));
  nor2  gate937(.a(gate278inter11), .b(gate278inter6), .O(gate278inter12));
  nand2 gate938(.a(gate278inter12), .b(gate278inter1), .O(G823));
nand2 gate279( .a(G651), .b(G803), .O(G824) );

  xor2  gate2465(.a(G803), .b(G779), .O(gate280inter0));
  nand2 gate2466(.a(gate280inter0), .b(s_274), .O(gate280inter1));
  and2  gate2467(.a(G803), .b(G779), .O(gate280inter2));
  inv1  gate2468(.a(s_274), .O(gate280inter3));
  inv1  gate2469(.a(s_275), .O(gate280inter4));
  nand2 gate2470(.a(gate280inter4), .b(gate280inter3), .O(gate280inter5));
  nor2  gate2471(.a(gate280inter5), .b(gate280inter2), .O(gate280inter6));
  inv1  gate2472(.a(G779), .O(gate280inter7));
  inv1  gate2473(.a(G803), .O(gate280inter8));
  nand2 gate2474(.a(gate280inter8), .b(gate280inter7), .O(gate280inter9));
  nand2 gate2475(.a(s_275), .b(gate280inter3), .O(gate280inter10));
  nor2  gate2476(.a(gate280inter10), .b(gate280inter9), .O(gate280inter11));
  nor2  gate2477(.a(gate280inter11), .b(gate280inter6), .O(gate280inter12));
  nand2 gate2478(.a(gate280inter12), .b(gate280inter1), .O(G825));
nand2 gate281( .a(G654), .b(G806), .O(G826) );

  xor2  gate729(.a(G806), .b(G782), .O(gate282inter0));
  nand2 gate730(.a(gate282inter0), .b(s_26), .O(gate282inter1));
  and2  gate731(.a(G806), .b(G782), .O(gate282inter2));
  inv1  gate732(.a(s_26), .O(gate282inter3));
  inv1  gate733(.a(s_27), .O(gate282inter4));
  nand2 gate734(.a(gate282inter4), .b(gate282inter3), .O(gate282inter5));
  nor2  gate735(.a(gate282inter5), .b(gate282inter2), .O(gate282inter6));
  inv1  gate736(.a(G782), .O(gate282inter7));
  inv1  gate737(.a(G806), .O(gate282inter8));
  nand2 gate738(.a(gate282inter8), .b(gate282inter7), .O(gate282inter9));
  nand2 gate739(.a(s_27), .b(gate282inter3), .O(gate282inter10));
  nor2  gate740(.a(gate282inter10), .b(gate282inter9), .O(gate282inter11));
  nor2  gate741(.a(gate282inter11), .b(gate282inter6), .O(gate282inter12));
  nand2 gate742(.a(gate282inter12), .b(gate282inter1), .O(G827));
nand2 gate283( .a(G657), .b(G809), .O(G828) );
nand2 gate284( .a(G785), .b(G809), .O(G829) );

  xor2  gate2843(.a(G812), .b(G660), .O(gate285inter0));
  nand2 gate2844(.a(gate285inter0), .b(s_328), .O(gate285inter1));
  and2  gate2845(.a(G812), .b(G660), .O(gate285inter2));
  inv1  gate2846(.a(s_328), .O(gate285inter3));
  inv1  gate2847(.a(s_329), .O(gate285inter4));
  nand2 gate2848(.a(gate285inter4), .b(gate285inter3), .O(gate285inter5));
  nor2  gate2849(.a(gate285inter5), .b(gate285inter2), .O(gate285inter6));
  inv1  gate2850(.a(G660), .O(gate285inter7));
  inv1  gate2851(.a(G812), .O(gate285inter8));
  nand2 gate2852(.a(gate285inter8), .b(gate285inter7), .O(gate285inter9));
  nand2 gate2853(.a(s_329), .b(gate285inter3), .O(gate285inter10));
  nor2  gate2854(.a(gate285inter10), .b(gate285inter9), .O(gate285inter11));
  nor2  gate2855(.a(gate285inter11), .b(gate285inter6), .O(gate285inter12));
  nand2 gate2856(.a(gate285inter12), .b(gate285inter1), .O(G830));

  xor2  gate1625(.a(G812), .b(G788), .O(gate286inter0));
  nand2 gate1626(.a(gate286inter0), .b(s_154), .O(gate286inter1));
  and2  gate1627(.a(G812), .b(G788), .O(gate286inter2));
  inv1  gate1628(.a(s_154), .O(gate286inter3));
  inv1  gate1629(.a(s_155), .O(gate286inter4));
  nand2 gate1630(.a(gate286inter4), .b(gate286inter3), .O(gate286inter5));
  nor2  gate1631(.a(gate286inter5), .b(gate286inter2), .O(gate286inter6));
  inv1  gate1632(.a(G788), .O(gate286inter7));
  inv1  gate1633(.a(G812), .O(gate286inter8));
  nand2 gate1634(.a(gate286inter8), .b(gate286inter7), .O(gate286inter9));
  nand2 gate1635(.a(s_155), .b(gate286inter3), .O(gate286inter10));
  nor2  gate1636(.a(gate286inter10), .b(gate286inter9), .O(gate286inter11));
  nor2  gate1637(.a(gate286inter11), .b(gate286inter6), .O(gate286inter12));
  nand2 gate1638(.a(gate286inter12), .b(gate286inter1), .O(G831));

  xor2  gate2899(.a(G815), .b(G663), .O(gate287inter0));
  nand2 gate2900(.a(gate287inter0), .b(s_336), .O(gate287inter1));
  and2  gate2901(.a(G815), .b(G663), .O(gate287inter2));
  inv1  gate2902(.a(s_336), .O(gate287inter3));
  inv1  gate2903(.a(s_337), .O(gate287inter4));
  nand2 gate2904(.a(gate287inter4), .b(gate287inter3), .O(gate287inter5));
  nor2  gate2905(.a(gate287inter5), .b(gate287inter2), .O(gate287inter6));
  inv1  gate2906(.a(G663), .O(gate287inter7));
  inv1  gate2907(.a(G815), .O(gate287inter8));
  nand2 gate2908(.a(gate287inter8), .b(gate287inter7), .O(gate287inter9));
  nand2 gate2909(.a(s_337), .b(gate287inter3), .O(gate287inter10));
  nor2  gate2910(.a(gate287inter10), .b(gate287inter9), .O(gate287inter11));
  nor2  gate2911(.a(gate287inter11), .b(gate287inter6), .O(gate287inter12));
  nand2 gate2912(.a(gate287inter12), .b(gate287inter1), .O(G832));

  xor2  gate1975(.a(G815), .b(G791), .O(gate288inter0));
  nand2 gate1976(.a(gate288inter0), .b(s_204), .O(gate288inter1));
  and2  gate1977(.a(G815), .b(G791), .O(gate288inter2));
  inv1  gate1978(.a(s_204), .O(gate288inter3));
  inv1  gate1979(.a(s_205), .O(gate288inter4));
  nand2 gate1980(.a(gate288inter4), .b(gate288inter3), .O(gate288inter5));
  nor2  gate1981(.a(gate288inter5), .b(gate288inter2), .O(gate288inter6));
  inv1  gate1982(.a(G791), .O(gate288inter7));
  inv1  gate1983(.a(G815), .O(gate288inter8));
  nand2 gate1984(.a(gate288inter8), .b(gate288inter7), .O(gate288inter9));
  nand2 gate1985(.a(s_205), .b(gate288inter3), .O(gate288inter10));
  nor2  gate1986(.a(gate288inter10), .b(gate288inter9), .O(gate288inter11));
  nor2  gate1987(.a(gate288inter11), .b(gate288inter6), .O(gate288inter12));
  nand2 gate1988(.a(gate288inter12), .b(gate288inter1), .O(G833));

  xor2  gate2283(.a(G819), .b(G818), .O(gate289inter0));
  nand2 gate2284(.a(gate289inter0), .b(s_248), .O(gate289inter1));
  and2  gate2285(.a(G819), .b(G818), .O(gate289inter2));
  inv1  gate2286(.a(s_248), .O(gate289inter3));
  inv1  gate2287(.a(s_249), .O(gate289inter4));
  nand2 gate2288(.a(gate289inter4), .b(gate289inter3), .O(gate289inter5));
  nor2  gate2289(.a(gate289inter5), .b(gate289inter2), .O(gate289inter6));
  inv1  gate2290(.a(G818), .O(gate289inter7));
  inv1  gate2291(.a(G819), .O(gate289inter8));
  nand2 gate2292(.a(gate289inter8), .b(gate289inter7), .O(gate289inter9));
  nand2 gate2293(.a(s_249), .b(gate289inter3), .O(gate289inter10));
  nor2  gate2294(.a(gate289inter10), .b(gate289inter9), .O(gate289inter11));
  nor2  gate2295(.a(gate289inter11), .b(gate289inter6), .O(gate289inter12));
  nand2 gate2296(.a(gate289inter12), .b(gate289inter1), .O(G834));

  xor2  gate1205(.a(G821), .b(G820), .O(gate290inter0));
  nand2 gate1206(.a(gate290inter0), .b(s_94), .O(gate290inter1));
  and2  gate1207(.a(G821), .b(G820), .O(gate290inter2));
  inv1  gate1208(.a(s_94), .O(gate290inter3));
  inv1  gate1209(.a(s_95), .O(gate290inter4));
  nand2 gate1210(.a(gate290inter4), .b(gate290inter3), .O(gate290inter5));
  nor2  gate1211(.a(gate290inter5), .b(gate290inter2), .O(gate290inter6));
  inv1  gate1212(.a(G820), .O(gate290inter7));
  inv1  gate1213(.a(G821), .O(gate290inter8));
  nand2 gate1214(.a(gate290inter8), .b(gate290inter7), .O(gate290inter9));
  nand2 gate1215(.a(s_95), .b(gate290inter3), .O(gate290inter10));
  nor2  gate1216(.a(gate290inter10), .b(gate290inter9), .O(gate290inter11));
  nor2  gate1217(.a(gate290inter11), .b(gate290inter6), .O(gate290inter12));
  nand2 gate1218(.a(gate290inter12), .b(gate290inter1), .O(G847));
nand2 gate291( .a(G822), .b(G823), .O(G860) );
nand2 gate292( .a(G824), .b(G825), .O(G873) );
nand2 gate293( .a(G828), .b(G829), .O(G886) );

  xor2  gate841(.a(G833), .b(G832), .O(gate294inter0));
  nand2 gate842(.a(gate294inter0), .b(s_42), .O(gate294inter1));
  and2  gate843(.a(G833), .b(G832), .O(gate294inter2));
  inv1  gate844(.a(s_42), .O(gate294inter3));
  inv1  gate845(.a(s_43), .O(gate294inter4));
  nand2 gate846(.a(gate294inter4), .b(gate294inter3), .O(gate294inter5));
  nor2  gate847(.a(gate294inter5), .b(gate294inter2), .O(gate294inter6));
  inv1  gate848(.a(G832), .O(gate294inter7));
  inv1  gate849(.a(G833), .O(gate294inter8));
  nand2 gate850(.a(gate294inter8), .b(gate294inter7), .O(gate294inter9));
  nand2 gate851(.a(s_43), .b(gate294inter3), .O(gate294inter10));
  nor2  gate852(.a(gate294inter10), .b(gate294inter9), .O(gate294inter11));
  nor2  gate853(.a(gate294inter11), .b(gate294inter6), .O(gate294inter12));
  nand2 gate854(.a(gate294inter12), .b(gate294inter1), .O(G899));
nand2 gate295( .a(G830), .b(G831), .O(G912) );
nand2 gate296( .a(G826), .b(G827), .O(G925) );
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );

  xor2  gate855(.a(G1036), .b(G1), .O(gate387inter0));
  nand2 gate856(.a(gate387inter0), .b(s_44), .O(gate387inter1));
  and2  gate857(.a(G1036), .b(G1), .O(gate387inter2));
  inv1  gate858(.a(s_44), .O(gate387inter3));
  inv1  gate859(.a(s_45), .O(gate387inter4));
  nand2 gate860(.a(gate387inter4), .b(gate387inter3), .O(gate387inter5));
  nor2  gate861(.a(gate387inter5), .b(gate387inter2), .O(gate387inter6));
  inv1  gate862(.a(G1), .O(gate387inter7));
  inv1  gate863(.a(G1036), .O(gate387inter8));
  nand2 gate864(.a(gate387inter8), .b(gate387inter7), .O(gate387inter9));
  nand2 gate865(.a(s_45), .b(gate387inter3), .O(gate387inter10));
  nor2  gate866(.a(gate387inter10), .b(gate387inter9), .O(gate387inter11));
  nor2  gate867(.a(gate387inter11), .b(gate387inter6), .O(gate387inter12));
  nand2 gate868(.a(gate387inter12), .b(gate387inter1), .O(G1132));

  xor2  gate2913(.a(G1039), .b(G2), .O(gate388inter0));
  nand2 gate2914(.a(gate388inter0), .b(s_338), .O(gate388inter1));
  and2  gate2915(.a(G1039), .b(G2), .O(gate388inter2));
  inv1  gate2916(.a(s_338), .O(gate388inter3));
  inv1  gate2917(.a(s_339), .O(gate388inter4));
  nand2 gate2918(.a(gate388inter4), .b(gate388inter3), .O(gate388inter5));
  nor2  gate2919(.a(gate388inter5), .b(gate388inter2), .O(gate388inter6));
  inv1  gate2920(.a(G2), .O(gate388inter7));
  inv1  gate2921(.a(G1039), .O(gate388inter8));
  nand2 gate2922(.a(gate388inter8), .b(gate388inter7), .O(gate388inter9));
  nand2 gate2923(.a(s_339), .b(gate388inter3), .O(gate388inter10));
  nor2  gate2924(.a(gate388inter10), .b(gate388inter9), .O(gate388inter11));
  nor2  gate2925(.a(gate388inter11), .b(gate388inter6), .O(gate388inter12));
  nand2 gate2926(.a(gate388inter12), .b(gate388inter1), .O(G1135));

  xor2  gate1037(.a(G1042), .b(G3), .O(gate389inter0));
  nand2 gate1038(.a(gate389inter0), .b(s_70), .O(gate389inter1));
  and2  gate1039(.a(G1042), .b(G3), .O(gate389inter2));
  inv1  gate1040(.a(s_70), .O(gate389inter3));
  inv1  gate1041(.a(s_71), .O(gate389inter4));
  nand2 gate1042(.a(gate389inter4), .b(gate389inter3), .O(gate389inter5));
  nor2  gate1043(.a(gate389inter5), .b(gate389inter2), .O(gate389inter6));
  inv1  gate1044(.a(G3), .O(gate389inter7));
  inv1  gate1045(.a(G1042), .O(gate389inter8));
  nand2 gate1046(.a(gate389inter8), .b(gate389inter7), .O(gate389inter9));
  nand2 gate1047(.a(s_71), .b(gate389inter3), .O(gate389inter10));
  nor2  gate1048(.a(gate389inter10), .b(gate389inter9), .O(gate389inter11));
  nor2  gate1049(.a(gate389inter11), .b(gate389inter6), .O(gate389inter12));
  nand2 gate1050(.a(gate389inter12), .b(gate389inter1), .O(G1138));
nand2 gate390( .a(G4), .b(G1045), .O(G1141) );
nand2 gate391( .a(G5), .b(G1048), .O(G1144) );

  xor2  gate715(.a(G1051), .b(G6), .O(gate392inter0));
  nand2 gate716(.a(gate392inter0), .b(s_24), .O(gate392inter1));
  and2  gate717(.a(G1051), .b(G6), .O(gate392inter2));
  inv1  gate718(.a(s_24), .O(gate392inter3));
  inv1  gate719(.a(s_25), .O(gate392inter4));
  nand2 gate720(.a(gate392inter4), .b(gate392inter3), .O(gate392inter5));
  nor2  gate721(.a(gate392inter5), .b(gate392inter2), .O(gate392inter6));
  inv1  gate722(.a(G6), .O(gate392inter7));
  inv1  gate723(.a(G1051), .O(gate392inter8));
  nand2 gate724(.a(gate392inter8), .b(gate392inter7), .O(gate392inter9));
  nand2 gate725(.a(s_25), .b(gate392inter3), .O(gate392inter10));
  nor2  gate726(.a(gate392inter10), .b(gate392inter9), .O(gate392inter11));
  nor2  gate727(.a(gate392inter11), .b(gate392inter6), .O(gate392inter12));
  nand2 gate728(.a(gate392inter12), .b(gate392inter1), .O(G1147));
nand2 gate393( .a(G7), .b(G1054), .O(G1150) );

  xor2  gate2143(.a(G1057), .b(G8), .O(gate394inter0));
  nand2 gate2144(.a(gate394inter0), .b(s_228), .O(gate394inter1));
  and2  gate2145(.a(G1057), .b(G8), .O(gate394inter2));
  inv1  gate2146(.a(s_228), .O(gate394inter3));
  inv1  gate2147(.a(s_229), .O(gate394inter4));
  nand2 gate2148(.a(gate394inter4), .b(gate394inter3), .O(gate394inter5));
  nor2  gate2149(.a(gate394inter5), .b(gate394inter2), .O(gate394inter6));
  inv1  gate2150(.a(G8), .O(gate394inter7));
  inv1  gate2151(.a(G1057), .O(gate394inter8));
  nand2 gate2152(.a(gate394inter8), .b(gate394inter7), .O(gate394inter9));
  nand2 gate2153(.a(s_229), .b(gate394inter3), .O(gate394inter10));
  nor2  gate2154(.a(gate394inter10), .b(gate394inter9), .O(gate394inter11));
  nor2  gate2155(.a(gate394inter11), .b(gate394inter6), .O(gate394inter12));
  nand2 gate2156(.a(gate394inter12), .b(gate394inter1), .O(G1153));

  xor2  gate645(.a(G1060), .b(G9), .O(gate395inter0));
  nand2 gate646(.a(gate395inter0), .b(s_14), .O(gate395inter1));
  and2  gate647(.a(G1060), .b(G9), .O(gate395inter2));
  inv1  gate648(.a(s_14), .O(gate395inter3));
  inv1  gate649(.a(s_15), .O(gate395inter4));
  nand2 gate650(.a(gate395inter4), .b(gate395inter3), .O(gate395inter5));
  nor2  gate651(.a(gate395inter5), .b(gate395inter2), .O(gate395inter6));
  inv1  gate652(.a(G9), .O(gate395inter7));
  inv1  gate653(.a(G1060), .O(gate395inter8));
  nand2 gate654(.a(gate395inter8), .b(gate395inter7), .O(gate395inter9));
  nand2 gate655(.a(s_15), .b(gate395inter3), .O(gate395inter10));
  nor2  gate656(.a(gate395inter10), .b(gate395inter9), .O(gate395inter11));
  nor2  gate657(.a(gate395inter11), .b(gate395inter6), .O(gate395inter12));
  nand2 gate658(.a(gate395inter12), .b(gate395inter1), .O(G1156));
nand2 gate396( .a(G10), .b(G1063), .O(G1159) );
nand2 gate397( .a(G11), .b(G1066), .O(G1162) );
nand2 gate398( .a(G12), .b(G1069), .O(G1165) );

  xor2  gate2619(.a(G1072), .b(G13), .O(gate399inter0));
  nand2 gate2620(.a(gate399inter0), .b(s_296), .O(gate399inter1));
  and2  gate2621(.a(G1072), .b(G13), .O(gate399inter2));
  inv1  gate2622(.a(s_296), .O(gate399inter3));
  inv1  gate2623(.a(s_297), .O(gate399inter4));
  nand2 gate2624(.a(gate399inter4), .b(gate399inter3), .O(gate399inter5));
  nor2  gate2625(.a(gate399inter5), .b(gate399inter2), .O(gate399inter6));
  inv1  gate2626(.a(G13), .O(gate399inter7));
  inv1  gate2627(.a(G1072), .O(gate399inter8));
  nand2 gate2628(.a(gate399inter8), .b(gate399inter7), .O(gate399inter9));
  nand2 gate2629(.a(s_297), .b(gate399inter3), .O(gate399inter10));
  nor2  gate2630(.a(gate399inter10), .b(gate399inter9), .O(gate399inter11));
  nor2  gate2631(.a(gate399inter11), .b(gate399inter6), .O(gate399inter12));
  nand2 gate2632(.a(gate399inter12), .b(gate399inter1), .O(G1168));

  xor2  gate2003(.a(G1075), .b(G14), .O(gate400inter0));
  nand2 gate2004(.a(gate400inter0), .b(s_208), .O(gate400inter1));
  and2  gate2005(.a(G1075), .b(G14), .O(gate400inter2));
  inv1  gate2006(.a(s_208), .O(gate400inter3));
  inv1  gate2007(.a(s_209), .O(gate400inter4));
  nand2 gate2008(.a(gate400inter4), .b(gate400inter3), .O(gate400inter5));
  nor2  gate2009(.a(gate400inter5), .b(gate400inter2), .O(gate400inter6));
  inv1  gate2010(.a(G14), .O(gate400inter7));
  inv1  gate2011(.a(G1075), .O(gate400inter8));
  nand2 gate2012(.a(gate400inter8), .b(gate400inter7), .O(gate400inter9));
  nand2 gate2013(.a(s_209), .b(gate400inter3), .O(gate400inter10));
  nor2  gate2014(.a(gate400inter10), .b(gate400inter9), .O(gate400inter11));
  nor2  gate2015(.a(gate400inter11), .b(gate400inter6), .O(gate400inter12));
  nand2 gate2016(.a(gate400inter12), .b(gate400inter1), .O(G1171));
nand2 gate401( .a(G15), .b(G1078), .O(G1174) );

  xor2  gate2885(.a(G1081), .b(G16), .O(gate402inter0));
  nand2 gate2886(.a(gate402inter0), .b(s_334), .O(gate402inter1));
  and2  gate2887(.a(G1081), .b(G16), .O(gate402inter2));
  inv1  gate2888(.a(s_334), .O(gate402inter3));
  inv1  gate2889(.a(s_335), .O(gate402inter4));
  nand2 gate2890(.a(gate402inter4), .b(gate402inter3), .O(gate402inter5));
  nor2  gate2891(.a(gate402inter5), .b(gate402inter2), .O(gate402inter6));
  inv1  gate2892(.a(G16), .O(gate402inter7));
  inv1  gate2893(.a(G1081), .O(gate402inter8));
  nand2 gate2894(.a(gate402inter8), .b(gate402inter7), .O(gate402inter9));
  nand2 gate2895(.a(s_335), .b(gate402inter3), .O(gate402inter10));
  nor2  gate2896(.a(gate402inter10), .b(gate402inter9), .O(gate402inter11));
  nor2  gate2897(.a(gate402inter11), .b(gate402inter6), .O(gate402inter12));
  nand2 gate2898(.a(gate402inter12), .b(gate402inter1), .O(G1177));
nand2 gate403( .a(G17), .b(G1084), .O(G1180) );

  xor2  gate897(.a(G1087), .b(G18), .O(gate404inter0));
  nand2 gate898(.a(gate404inter0), .b(s_50), .O(gate404inter1));
  and2  gate899(.a(G1087), .b(G18), .O(gate404inter2));
  inv1  gate900(.a(s_50), .O(gate404inter3));
  inv1  gate901(.a(s_51), .O(gate404inter4));
  nand2 gate902(.a(gate404inter4), .b(gate404inter3), .O(gate404inter5));
  nor2  gate903(.a(gate404inter5), .b(gate404inter2), .O(gate404inter6));
  inv1  gate904(.a(G18), .O(gate404inter7));
  inv1  gate905(.a(G1087), .O(gate404inter8));
  nand2 gate906(.a(gate404inter8), .b(gate404inter7), .O(gate404inter9));
  nand2 gate907(.a(s_51), .b(gate404inter3), .O(gate404inter10));
  nor2  gate908(.a(gate404inter10), .b(gate404inter9), .O(gate404inter11));
  nor2  gate909(.a(gate404inter11), .b(gate404inter6), .O(gate404inter12));
  nand2 gate910(.a(gate404inter12), .b(gate404inter1), .O(G1183));

  xor2  gate2255(.a(G1090), .b(G19), .O(gate405inter0));
  nand2 gate2256(.a(gate405inter0), .b(s_244), .O(gate405inter1));
  and2  gate2257(.a(G1090), .b(G19), .O(gate405inter2));
  inv1  gate2258(.a(s_244), .O(gate405inter3));
  inv1  gate2259(.a(s_245), .O(gate405inter4));
  nand2 gate2260(.a(gate405inter4), .b(gate405inter3), .O(gate405inter5));
  nor2  gate2261(.a(gate405inter5), .b(gate405inter2), .O(gate405inter6));
  inv1  gate2262(.a(G19), .O(gate405inter7));
  inv1  gate2263(.a(G1090), .O(gate405inter8));
  nand2 gate2264(.a(gate405inter8), .b(gate405inter7), .O(gate405inter9));
  nand2 gate2265(.a(s_245), .b(gate405inter3), .O(gate405inter10));
  nor2  gate2266(.a(gate405inter10), .b(gate405inter9), .O(gate405inter11));
  nor2  gate2267(.a(gate405inter11), .b(gate405inter6), .O(gate405inter12));
  nand2 gate2268(.a(gate405inter12), .b(gate405inter1), .O(G1186));
nand2 gate406( .a(G20), .b(G1093), .O(G1189) );

  xor2  gate2437(.a(G1096), .b(G21), .O(gate407inter0));
  nand2 gate2438(.a(gate407inter0), .b(s_270), .O(gate407inter1));
  and2  gate2439(.a(G1096), .b(G21), .O(gate407inter2));
  inv1  gate2440(.a(s_270), .O(gate407inter3));
  inv1  gate2441(.a(s_271), .O(gate407inter4));
  nand2 gate2442(.a(gate407inter4), .b(gate407inter3), .O(gate407inter5));
  nor2  gate2443(.a(gate407inter5), .b(gate407inter2), .O(gate407inter6));
  inv1  gate2444(.a(G21), .O(gate407inter7));
  inv1  gate2445(.a(G1096), .O(gate407inter8));
  nand2 gate2446(.a(gate407inter8), .b(gate407inter7), .O(gate407inter9));
  nand2 gate2447(.a(s_271), .b(gate407inter3), .O(gate407inter10));
  nor2  gate2448(.a(gate407inter10), .b(gate407inter9), .O(gate407inter11));
  nor2  gate2449(.a(gate407inter11), .b(gate407inter6), .O(gate407inter12));
  nand2 gate2450(.a(gate407inter12), .b(gate407inter1), .O(G1192));
nand2 gate408( .a(G22), .b(G1099), .O(G1195) );
nand2 gate409( .a(G23), .b(G1102), .O(G1198) );

  xor2  gate911(.a(G1105), .b(G24), .O(gate410inter0));
  nand2 gate912(.a(gate410inter0), .b(s_52), .O(gate410inter1));
  and2  gate913(.a(G1105), .b(G24), .O(gate410inter2));
  inv1  gate914(.a(s_52), .O(gate410inter3));
  inv1  gate915(.a(s_53), .O(gate410inter4));
  nand2 gate916(.a(gate410inter4), .b(gate410inter3), .O(gate410inter5));
  nor2  gate917(.a(gate410inter5), .b(gate410inter2), .O(gate410inter6));
  inv1  gate918(.a(G24), .O(gate410inter7));
  inv1  gate919(.a(G1105), .O(gate410inter8));
  nand2 gate920(.a(gate410inter8), .b(gate410inter7), .O(gate410inter9));
  nand2 gate921(.a(s_53), .b(gate410inter3), .O(gate410inter10));
  nor2  gate922(.a(gate410inter10), .b(gate410inter9), .O(gate410inter11));
  nor2  gate923(.a(gate410inter11), .b(gate410inter6), .O(gate410inter12));
  nand2 gate924(.a(gate410inter12), .b(gate410inter1), .O(G1201));

  xor2  gate1947(.a(G1108), .b(G25), .O(gate411inter0));
  nand2 gate1948(.a(gate411inter0), .b(s_200), .O(gate411inter1));
  and2  gate1949(.a(G1108), .b(G25), .O(gate411inter2));
  inv1  gate1950(.a(s_200), .O(gate411inter3));
  inv1  gate1951(.a(s_201), .O(gate411inter4));
  nand2 gate1952(.a(gate411inter4), .b(gate411inter3), .O(gate411inter5));
  nor2  gate1953(.a(gate411inter5), .b(gate411inter2), .O(gate411inter6));
  inv1  gate1954(.a(G25), .O(gate411inter7));
  inv1  gate1955(.a(G1108), .O(gate411inter8));
  nand2 gate1956(.a(gate411inter8), .b(gate411inter7), .O(gate411inter9));
  nand2 gate1957(.a(s_201), .b(gate411inter3), .O(gate411inter10));
  nor2  gate1958(.a(gate411inter10), .b(gate411inter9), .O(gate411inter11));
  nor2  gate1959(.a(gate411inter11), .b(gate411inter6), .O(gate411inter12));
  nand2 gate1960(.a(gate411inter12), .b(gate411inter1), .O(G1204));

  xor2  gate2829(.a(G1111), .b(G26), .O(gate412inter0));
  nand2 gate2830(.a(gate412inter0), .b(s_326), .O(gate412inter1));
  and2  gate2831(.a(G1111), .b(G26), .O(gate412inter2));
  inv1  gate2832(.a(s_326), .O(gate412inter3));
  inv1  gate2833(.a(s_327), .O(gate412inter4));
  nand2 gate2834(.a(gate412inter4), .b(gate412inter3), .O(gate412inter5));
  nor2  gate2835(.a(gate412inter5), .b(gate412inter2), .O(gate412inter6));
  inv1  gate2836(.a(G26), .O(gate412inter7));
  inv1  gate2837(.a(G1111), .O(gate412inter8));
  nand2 gate2838(.a(gate412inter8), .b(gate412inter7), .O(gate412inter9));
  nand2 gate2839(.a(s_327), .b(gate412inter3), .O(gate412inter10));
  nor2  gate2840(.a(gate412inter10), .b(gate412inter9), .O(gate412inter11));
  nor2  gate2841(.a(gate412inter11), .b(gate412inter6), .O(gate412inter12));
  nand2 gate2842(.a(gate412inter12), .b(gate412inter1), .O(G1207));

  xor2  gate1961(.a(G1114), .b(G27), .O(gate413inter0));
  nand2 gate1962(.a(gate413inter0), .b(s_202), .O(gate413inter1));
  and2  gate1963(.a(G1114), .b(G27), .O(gate413inter2));
  inv1  gate1964(.a(s_202), .O(gate413inter3));
  inv1  gate1965(.a(s_203), .O(gate413inter4));
  nand2 gate1966(.a(gate413inter4), .b(gate413inter3), .O(gate413inter5));
  nor2  gate1967(.a(gate413inter5), .b(gate413inter2), .O(gate413inter6));
  inv1  gate1968(.a(G27), .O(gate413inter7));
  inv1  gate1969(.a(G1114), .O(gate413inter8));
  nand2 gate1970(.a(gate413inter8), .b(gate413inter7), .O(gate413inter9));
  nand2 gate1971(.a(s_203), .b(gate413inter3), .O(gate413inter10));
  nor2  gate1972(.a(gate413inter10), .b(gate413inter9), .O(gate413inter11));
  nor2  gate1973(.a(gate413inter11), .b(gate413inter6), .O(gate413inter12));
  nand2 gate1974(.a(gate413inter12), .b(gate413inter1), .O(G1210));

  xor2  gate2647(.a(G1117), .b(G28), .O(gate414inter0));
  nand2 gate2648(.a(gate414inter0), .b(s_300), .O(gate414inter1));
  and2  gate2649(.a(G1117), .b(G28), .O(gate414inter2));
  inv1  gate2650(.a(s_300), .O(gate414inter3));
  inv1  gate2651(.a(s_301), .O(gate414inter4));
  nand2 gate2652(.a(gate414inter4), .b(gate414inter3), .O(gate414inter5));
  nor2  gate2653(.a(gate414inter5), .b(gate414inter2), .O(gate414inter6));
  inv1  gate2654(.a(G28), .O(gate414inter7));
  inv1  gate2655(.a(G1117), .O(gate414inter8));
  nand2 gate2656(.a(gate414inter8), .b(gate414inter7), .O(gate414inter9));
  nand2 gate2657(.a(s_301), .b(gate414inter3), .O(gate414inter10));
  nor2  gate2658(.a(gate414inter10), .b(gate414inter9), .O(gate414inter11));
  nor2  gate2659(.a(gate414inter11), .b(gate414inter6), .O(gate414inter12));
  nand2 gate2660(.a(gate414inter12), .b(gate414inter1), .O(G1213));

  xor2  gate2353(.a(G1120), .b(G29), .O(gate415inter0));
  nand2 gate2354(.a(gate415inter0), .b(s_258), .O(gate415inter1));
  and2  gate2355(.a(G1120), .b(G29), .O(gate415inter2));
  inv1  gate2356(.a(s_258), .O(gate415inter3));
  inv1  gate2357(.a(s_259), .O(gate415inter4));
  nand2 gate2358(.a(gate415inter4), .b(gate415inter3), .O(gate415inter5));
  nor2  gate2359(.a(gate415inter5), .b(gate415inter2), .O(gate415inter6));
  inv1  gate2360(.a(G29), .O(gate415inter7));
  inv1  gate2361(.a(G1120), .O(gate415inter8));
  nand2 gate2362(.a(gate415inter8), .b(gate415inter7), .O(gate415inter9));
  nand2 gate2363(.a(s_259), .b(gate415inter3), .O(gate415inter10));
  nor2  gate2364(.a(gate415inter10), .b(gate415inter9), .O(gate415inter11));
  nor2  gate2365(.a(gate415inter11), .b(gate415inter6), .O(gate415inter12));
  nand2 gate2366(.a(gate415inter12), .b(gate415inter1), .O(G1216));

  xor2  gate3039(.a(G1123), .b(G30), .O(gate416inter0));
  nand2 gate3040(.a(gate416inter0), .b(s_356), .O(gate416inter1));
  and2  gate3041(.a(G1123), .b(G30), .O(gate416inter2));
  inv1  gate3042(.a(s_356), .O(gate416inter3));
  inv1  gate3043(.a(s_357), .O(gate416inter4));
  nand2 gate3044(.a(gate416inter4), .b(gate416inter3), .O(gate416inter5));
  nor2  gate3045(.a(gate416inter5), .b(gate416inter2), .O(gate416inter6));
  inv1  gate3046(.a(G30), .O(gate416inter7));
  inv1  gate3047(.a(G1123), .O(gate416inter8));
  nand2 gate3048(.a(gate416inter8), .b(gate416inter7), .O(gate416inter9));
  nand2 gate3049(.a(s_357), .b(gate416inter3), .O(gate416inter10));
  nor2  gate3050(.a(gate416inter10), .b(gate416inter9), .O(gate416inter11));
  nor2  gate3051(.a(gate416inter11), .b(gate416inter6), .O(gate416inter12));
  nand2 gate3052(.a(gate416inter12), .b(gate416inter1), .O(G1219));

  xor2  gate2367(.a(G1126), .b(G31), .O(gate417inter0));
  nand2 gate2368(.a(gate417inter0), .b(s_260), .O(gate417inter1));
  and2  gate2369(.a(G1126), .b(G31), .O(gate417inter2));
  inv1  gate2370(.a(s_260), .O(gate417inter3));
  inv1  gate2371(.a(s_261), .O(gate417inter4));
  nand2 gate2372(.a(gate417inter4), .b(gate417inter3), .O(gate417inter5));
  nor2  gate2373(.a(gate417inter5), .b(gate417inter2), .O(gate417inter6));
  inv1  gate2374(.a(G31), .O(gate417inter7));
  inv1  gate2375(.a(G1126), .O(gate417inter8));
  nand2 gate2376(.a(gate417inter8), .b(gate417inter7), .O(gate417inter9));
  nand2 gate2377(.a(s_261), .b(gate417inter3), .O(gate417inter10));
  nor2  gate2378(.a(gate417inter10), .b(gate417inter9), .O(gate417inter11));
  nor2  gate2379(.a(gate417inter11), .b(gate417inter6), .O(gate417inter12));
  nand2 gate2380(.a(gate417inter12), .b(gate417inter1), .O(G1222));
nand2 gate418( .a(G32), .b(G1129), .O(G1225) );
nand2 gate419( .a(G1), .b(G1132), .O(G1228) );
nand2 gate420( .a(G1036), .b(G1132), .O(G1229) );
nand2 gate421( .a(G2), .b(G1135), .O(G1230) );

  xor2  gate2871(.a(G1135), .b(G1039), .O(gate422inter0));
  nand2 gate2872(.a(gate422inter0), .b(s_332), .O(gate422inter1));
  and2  gate2873(.a(G1135), .b(G1039), .O(gate422inter2));
  inv1  gate2874(.a(s_332), .O(gate422inter3));
  inv1  gate2875(.a(s_333), .O(gate422inter4));
  nand2 gate2876(.a(gate422inter4), .b(gate422inter3), .O(gate422inter5));
  nor2  gate2877(.a(gate422inter5), .b(gate422inter2), .O(gate422inter6));
  inv1  gate2878(.a(G1039), .O(gate422inter7));
  inv1  gate2879(.a(G1135), .O(gate422inter8));
  nand2 gate2880(.a(gate422inter8), .b(gate422inter7), .O(gate422inter9));
  nand2 gate2881(.a(s_333), .b(gate422inter3), .O(gate422inter10));
  nor2  gate2882(.a(gate422inter10), .b(gate422inter9), .O(gate422inter11));
  nor2  gate2883(.a(gate422inter11), .b(gate422inter6), .O(gate422inter12));
  nand2 gate2884(.a(gate422inter12), .b(gate422inter1), .O(G1231));

  xor2  gate1149(.a(G1138), .b(G3), .O(gate423inter0));
  nand2 gate1150(.a(gate423inter0), .b(s_86), .O(gate423inter1));
  and2  gate1151(.a(G1138), .b(G3), .O(gate423inter2));
  inv1  gate1152(.a(s_86), .O(gate423inter3));
  inv1  gate1153(.a(s_87), .O(gate423inter4));
  nand2 gate1154(.a(gate423inter4), .b(gate423inter3), .O(gate423inter5));
  nor2  gate1155(.a(gate423inter5), .b(gate423inter2), .O(gate423inter6));
  inv1  gate1156(.a(G3), .O(gate423inter7));
  inv1  gate1157(.a(G1138), .O(gate423inter8));
  nand2 gate1158(.a(gate423inter8), .b(gate423inter7), .O(gate423inter9));
  nand2 gate1159(.a(s_87), .b(gate423inter3), .O(gate423inter10));
  nor2  gate1160(.a(gate423inter10), .b(gate423inter9), .O(gate423inter11));
  nor2  gate1161(.a(gate423inter11), .b(gate423inter6), .O(gate423inter12));
  nand2 gate1162(.a(gate423inter12), .b(gate423inter1), .O(G1232));

  xor2  gate1359(.a(G1138), .b(G1042), .O(gate424inter0));
  nand2 gate1360(.a(gate424inter0), .b(s_116), .O(gate424inter1));
  and2  gate1361(.a(G1138), .b(G1042), .O(gate424inter2));
  inv1  gate1362(.a(s_116), .O(gate424inter3));
  inv1  gate1363(.a(s_117), .O(gate424inter4));
  nand2 gate1364(.a(gate424inter4), .b(gate424inter3), .O(gate424inter5));
  nor2  gate1365(.a(gate424inter5), .b(gate424inter2), .O(gate424inter6));
  inv1  gate1366(.a(G1042), .O(gate424inter7));
  inv1  gate1367(.a(G1138), .O(gate424inter8));
  nand2 gate1368(.a(gate424inter8), .b(gate424inter7), .O(gate424inter9));
  nand2 gate1369(.a(s_117), .b(gate424inter3), .O(gate424inter10));
  nor2  gate1370(.a(gate424inter10), .b(gate424inter9), .O(gate424inter11));
  nor2  gate1371(.a(gate424inter11), .b(gate424inter6), .O(gate424inter12));
  nand2 gate1372(.a(gate424inter12), .b(gate424inter1), .O(G1233));

  xor2  gate1345(.a(G1141), .b(G4), .O(gate425inter0));
  nand2 gate1346(.a(gate425inter0), .b(s_114), .O(gate425inter1));
  and2  gate1347(.a(G1141), .b(G4), .O(gate425inter2));
  inv1  gate1348(.a(s_114), .O(gate425inter3));
  inv1  gate1349(.a(s_115), .O(gate425inter4));
  nand2 gate1350(.a(gate425inter4), .b(gate425inter3), .O(gate425inter5));
  nor2  gate1351(.a(gate425inter5), .b(gate425inter2), .O(gate425inter6));
  inv1  gate1352(.a(G4), .O(gate425inter7));
  inv1  gate1353(.a(G1141), .O(gate425inter8));
  nand2 gate1354(.a(gate425inter8), .b(gate425inter7), .O(gate425inter9));
  nand2 gate1355(.a(s_115), .b(gate425inter3), .O(gate425inter10));
  nor2  gate1356(.a(gate425inter10), .b(gate425inter9), .O(gate425inter11));
  nor2  gate1357(.a(gate425inter11), .b(gate425inter6), .O(gate425inter12));
  nand2 gate1358(.a(gate425inter12), .b(gate425inter1), .O(G1234));

  xor2  gate1877(.a(G1141), .b(G1045), .O(gate426inter0));
  nand2 gate1878(.a(gate426inter0), .b(s_190), .O(gate426inter1));
  and2  gate1879(.a(G1141), .b(G1045), .O(gate426inter2));
  inv1  gate1880(.a(s_190), .O(gate426inter3));
  inv1  gate1881(.a(s_191), .O(gate426inter4));
  nand2 gate1882(.a(gate426inter4), .b(gate426inter3), .O(gate426inter5));
  nor2  gate1883(.a(gate426inter5), .b(gate426inter2), .O(gate426inter6));
  inv1  gate1884(.a(G1045), .O(gate426inter7));
  inv1  gate1885(.a(G1141), .O(gate426inter8));
  nand2 gate1886(.a(gate426inter8), .b(gate426inter7), .O(gate426inter9));
  nand2 gate1887(.a(s_191), .b(gate426inter3), .O(gate426inter10));
  nor2  gate1888(.a(gate426inter10), .b(gate426inter9), .O(gate426inter11));
  nor2  gate1889(.a(gate426inter11), .b(gate426inter6), .O(gate426inter12));
  nand2 gate1890(.a(gate426inter12), .b(gate426inter1), .O(G1235));
nand2 gate427( .a(G5), .b(G1144), .O(G1236) );

  xor2  gate1429(.a(G1144), .b(G1048), .O(gate428inter0));
  nand2 gate1430(.a(gate428inter0), .b(s_126), .O(gate428inter1));
  and2  gate1431(.a(G1144), .b(G1048), .O(gate428inter2));
  inv1  gate1432(.a(s_126), .O(gate428inter3));
  inv1  gate1433(.a(s_127), .O(gate428inter4));
  nand2 gate1434(.a(gate428inter4), .b(gate428inter3), .O(gate428inter5));
  nor2  gate1435(.a(gate428inter5), .b(gate428inter2), .O(gate428inter6));
  inv1  gate1436(.a(G1048), .O(gate428inter7));
  inv1  gate1437(.a(G1144), .O(gate428inter8));
  nand2 gate1438(.a(gate428inter8), .b(gate428inter7), .O(gate428inter9));
  nand2 gate1439(.a(s_127), .b(gate428inter3), .O(gate428inter10));
  nor2  gate1440(.a(gate428inter10), .b(gate428inter9), .O(gate428inter11));
  nor2  gate1441(.a(gate428inter11), .b(gate428inter6), .O(gate428inter12));
  nand2 gate1442(.a(gate428inter12), .b(gate428inter1), .O(G1237));
nand2 gate429( .a(G6), .b(G1147), .O(G1238) );
nand2 gate430( .a(G1051), .b(G1147), .O(G1239) );

  xor2  gate869(.a(G1150), .b(G7), .O(gate431inter0));
  nand2 gate870(.a(gate431inter0), .b(s_46), .O(gate431inter1));
  and2  gate871(.a(G1150), .b(G7), .O(gate431inter2));
  inv1  gate872(.a(s_46), .O(gate431inter3));
  inv1  gate873(.a(s_47), .O(gate431inter4));
  nand2 gate874(.a(gate431inter4), .b(gate431inter3), .O(gate431inter5));
  nor2  gate875(.a(gate431inter5), .b(gate431inter2), .O(gate431inter6));
  inv1  gate876(.a(G7), .O(gate431inter7));
  inv1  gate877(.a(G1150), .O(gate431inter8));
  nand2 gate878(.a(gate431inter8), .b(gate431inter7), .O(gate431inter9));
  nand2 gate879(.a(s_47), .b(gate431inter3), .O(gate431inter10));
  nor2  gate880(.a(gate431inter10), .b(gate431inter9), .O(gate431inter11));
  nor2  gate881(.a(gate431inter11), .b(gate431inter6), .O(gate431inter12));
  nand2 gate882(.a(gate431inter12), .b(gate431inter1), .O(G1240));
nand2 gate432( .a(G1054), .b(G1150), .O(G1241) );

  xor2  gate1695(.a(G1153), .b(G8), .O(gate433inter0));
  nand2 gate1696(.a(gate433inter0), .b(s_164), .O(gate433inter1));
  and2  gate1697(.a(G1153), .b(G8), .O(gate433inter2));
  inv1  gate1698(.a(s_164), .O(gate433inter3));
  inv1  gate1699(.a(s_165), .O(gate433inter4));
  nand2 gate1700(.a(gate433inter4), .b(gate433inter3), .O(gate433inter5));
  nor2  gate1701(.a(gate433inter5), .b(gate433inter2), .O(gate433inter6));
  inv1  gate1702(.a(G8), .O(gate433inter7));
  inv1  gate1703(.a(G1153), .O(gate433inter8));
  nand2 gate1704(.a(gate433inter8), .b(gate433inter7), .O(gate433inter9));
  nand2 gate1705(.a(s_165), .b(gate433inter3), .O(gate433inter10));
  nor2  gate1706(.a(gate433inter10), .b(gate433inter9), .O(gate433inter11));
  nor2  gate1707(.a(gate433inter11), .b(gate433inter6), .O(gate433inter12));
  nand2 gate1708(.a(gate433inter12), .b(gate433inter1), .O(G1242));
nand2 gate434( .a(G1057), .b(G1153), .O(G1243) );
nand2 gate435( .a(G9), .b(G1156), .O(G1244) );
nand2 gate436( .a(G1060), .b(G1156), .O(G1245) );
nand2 gate437( .a(G10), .b(G1159), .O(G1246) );
nand2 gate438( .a(G1063), .b(G1159), .O(G1247) );
nand2 gate439( .a(G11), .b(G1162), .O(G1248) );
nand2 gate440( .a(G1066), .b(G1162), .O(G1249) );
nand2 gate441( .a(G12), .b(G1165), .O(G1250) );
nand2 gate442( .a(G1069), .b(G1165), .O(G1251) );

  xor2  gate1415(.a(G1168), .b(G13), .O(gate443inter0));
  nand2 gate1416(.a(gate443inter0), .b(s_124), .O(gate443inter1));
  and2  gate1417(.a(G1168), .b(G13), .O(gate443inter2));
  inv1  gate1418(.a(s_124), .O(gate443inter3));
  inv1  gate1419(.a(s_125), .O(gate443inter4));
  nand2 gate1420(.a(gate443inter4), .b(gate443inter3), .O(gate443inter5));
  nor2  gate1421(.a(gate443inter5), .b(gate443inter2), .O(gate443inter6));
  inv1  gate1422(.a(G13), .O(gate443inter7));
  inv1  gate1423(.a(G1168), .O(gate443inter8));
  nand2 gate1424(.a(gate443inter8), .b(gate443inter7), .O(gate443inter9));
  nand2 gate1425(.a(s_125), .b(gate443inter3), .O(gate443inter10));
  nor2  gate1426(.a(gate443inter10), .b(gate443inter9), .O(gate443inter11));
  nor2  gate1427(.a(gate443inter11), .b(gate443inter6), .O(gate443inter12));
  nand2 gate1428(.a(gate443inter12), .b(gate443inter1), .O(G1252));
nand2 gate444( .a(G1072), .b(G1168), .O(G1253) );
nand2 gate445( .a(G14), .b(G1171), .O(G1254) );
nand2 gate446( .a(G1075), .b(G1171), .O(G1255) );

  xor2  gate1065(.a(G1174), .b(G15), .O(gate447inter0));
  nand2 gate1066(.a(gate447inter0), .b(s_74), .O(gate447inter1));
  and2  gate1067(.a(G1174), .b(G15), .O(gate447inter2));
  inv1  gate1068(.a(s_74), .O(gate447inter3));
  inv1  gate1069(.a(s_75), .O(gate447inter4));
  nand2 gate1070(.a(gate447inter4), .b(gate447inter3), .O(gate447inter5));
  nor2  gate1071(.a(gate447inter5), .b(gate447inter2), .O(gate447inter6));
  inv1  gate1072(.a(G15), .O(gate447inter7));
  inv1  gate1073(.a(G1174), .O(gate447inter8));
  nand2 gate1074(.a(gate447inter8), .b(gate447inter7), .O(gate447inter9));
  nand2 gate1075(.a(s_75), .b(gate447inter3), .O(gate447inter10));
  nor2  gate1076(.a(gate447inter10), .b(gate447inter9), .O(gate447inter11));
  nor2  gate1077(.a(gate447inter11), .b(gate447inter6), .O(gate447inter12));
  nand2 gate1078(.a(gate447inter12), .b(gate447inter1), .O(G1256));

  xor2  gate2689(.a(G1174), .b(G1078), .O(gate448inter0));
  nand2 gate2690(.a(gate448inter0), .b(s_306), .O(gate448inter1));
  and2  gate2691(.a(G1174), .b(G1078), .O(gate448inter2));
  inv1  gate2692(.a(s_306), .O(gate448inter3));
  inv1  gate2693(.a(s_307), .O(gate448inter4));
  nand2 gate2694(.a(gate448inter4), .b(gate448inter3), .O(gate448inter5));
  nor2  gate2695(.a(gate448inter5), .b(gate448inter2), .O(gate448inter6));
  inv1  gate2696(.a(G1078), .O(gate448inter7));
  inv1  gate2697(.a(G1174), .O(gate448inter8));
  nand2 gate2698(.a(gate448inter8), .b(gate448inter7), .O(gate448inter9));
  nand2 gate2699(.a(s_307), .b(gate448inter3), .O(gate448inter10));
  nor2  gate2700(.a(gate448inter10), .b(gate448inter9), .O(gate448inter11));
  nor2  gate2701(.a(gate448inter11), .b(gate448inter6), .O(gate448inter12));
  nand2 gate2702(.a(gate448inter12), .b(gate448inter1), .O(G1257));

  xor2  gate2535(.a(G1177), .b(G16), .O(gate449inter0));
  nand2 gate2536(.a(gate449inter0), .b(s_284), .O(gate449inter1));
  and2  gate2537(.a(G1177), .b(G16), .O(gate449inter2));
  inv1  gate2538(.a(s_284), .O(gate449inter3));
  inv1  gate2539(.a(s_285), .O(gate449inter4));
  nand2 gate2540(.a(gate449inter4), .b(gate449inter3), .O(gate449inter5));
  nor2  gate2541(.a(gate449inter5), .b(gate449inter2), .O(gate449inter6));
  inv1  gate2542(.a(G16), .O(gate449inter7));
  inv1  gate2543(.a(G1177), .O(gate449inter8));
  nand2 gate2544(.a(gate449inter8), .b(gate449inter7), .O(gate449inter9));
  nand2 gate2545(.a(s_285), .b(gate449inter3), .O(gate449inter10));
  nor2  gate2546(.a(gate449inter10), .b(gate449inter9), .O(gate449inter11));
  nor2  gate2547(.a(gate449inter11), .b(gate449inter6), .O(gate449inter12));
  nand2 gate2548(.a(gate449inter12), .b(gate449inter1), .O(G1258));
nand2 gate450( .a(G1081), .b(G1177), .O(G1259) );
nand2 gate451( .a(G17), .b(G1180), .O(G1260) );
nand2 gate452( .a(G1084), .b(G1180), .O(G1261) );

  xor2  gate1331(.a(G1183), .b(G18), .O(gate453inter0));
  nand2 gate1332(.a(gate453inter0), .b(s_112), .O(gate453inter1));
  and2  gate1333(.a(G1183), .b(G18), .O(gate453inter2));
  inv1  gate1334(.a(s_112), .O(gate453inter3));
  inv1  gate1335(.a(s_113), .O(gate453inter4));
  nand2 gate1336(.a(gate453inter4), .b(gate453inter3), .O(gate453inter5));
  nor2  gate1337(.a(gate453inter5), .b(gate453inter2), .O(gate453inter6));
  inv1  gate1338(.a(G18), .O(gate453inter7));
  inv1  gate1339(.a(G1183), .O(gate453inter8));
  nand2 gate1340(.a(gate453inter8), .b(gate453inter7), .O(gate453inter9));
  nand2 gate1341(.a(s_113), .b(gate453inter3), .O(gate453inter10));
  nor2  gate1342(.a(gate453inter10), .b(gate453inter9), .O(gate453inter11));
  nor2  gate1343(.a(gate453inter11), .b(gate453inter6), .O(gate453inter12));
  nand2 gate1344(.a(gate453inter12), .b(gate453inter1), .O(G1262));
nand2 gate454( .a(G1087), .b(G1183), .O(G1263) );
nand2 gate455( .a(G19), .b(G1186), .O(G1264) );

  xor2  gate785(.a(G1186), .b(G1090), .O(gate456inter0));
  nand2 gate786(.a(gate456inter0), .b(s_34), .O(gate456inter1));
  and2  gate787(.a(G1186), .b(G1090), .O(gate456inter2));
  inv1  gate788(.a(s_34), .O(gate456inter3));
  inv1  gate789(.a(s_35), .O(gate456inter4));
  nand2 gate790(.a(gate456inter4), .b(gate456inter3), .O(gate456inter5));
  nor2  gate791(.a(gate456inter5), .b(gate456inter2), .O(gate456inter6));
  inv1  gate792(.a(G1090), .O(gate456inter7));
  inv1  gate793(.a(G1186), .O(gate456inter8));
  nand2 gate794(.a(gate456inter8), .b(gate456inter7), .O(gate456inter9));
  nand2 gate795(.a(s_35), .b(gate456inter3), .O(gate456inter10));
  nor2  gate796(.a(gate456inter10), .b(gate456inter9), .O(gate456inter11));
  nor2  gate797(.a(gate456inter11), .b(gate456inter6), .O(gate456inter12));
  nand2 gate798(.a(gate456inter12), .b(gate456inter1), .O(G1265));
nand2 gate457( .a(G20), .b(G1189), .O(G1266) );
nand2 gate458( .a(G1093), .b(G1189), .O(G1267) );

  xor2  gate1569(.a(G1192), .b(G21), .O(gate459inter0));
  nand2 gate1570(.a(gate459inter0), .b(s_146), .O(gate459inter1));
  and2  gate1571(.a(G1192), .b(G21), .O(gate459inter2));
  inv1  gate1572(.a(s_146), .O(gate459inter3));
  inv1  gate1573(.a(s_147), .O(gate459inter4));
  nand2 gate1574(.a(gate459inter4), .b(gate459inter3), .O(gate459inter5));
  nor2  gate1575(.a(gate459inter5), .b(gate459inter2), .O(gate459inter6));
  inv1  gate1576(.a(G21), .O(gate459inter7));
  inv1  gate1577(.a(G1192), .O(gate459inter8));
  nand2 gate1578(.a(gate459inter8), .b(gate459inter7), .O(gate459inter9));
  nand2 gate1579(.a(s_147), .b(gate459inter3), .O(gate459inter10));
  nor2  gate1580(.a(gate459inter10), .b(gate459inter9), .O(gate459inter11));
  nor2  gate1581(.a(gate459inter11), .b(gate459inter6), .O(gate459inter12));
  nand2 gate1582(.a(gate459inter12), .b(gate459inter1), .O(G1268));

  xor2  gate2507(.a(G1192), .b(G1096), .O(gate460inter0));
  nand2 gate2508(.a(gate460inter0), .b(s_280), .O(gate460inter1));
  and2  gate2509(.a(G1192), .b(G1096), .O(gate460inter2));
  inv1  gate2510(.a(s_280), .O(gate460inter3));
  inv1  gate2511(.a(s_281), .O(gate460inter4));
  nand2 gate2512(.a(gate460inter4), .b(gate460inter3), .O(gate460inter5));
  nor2  gate2513(.a(gate460inter5), .b(gate460inter2), .O(gate460inter6));
  inv1  gate2514(.a(G1096), .O(gate460inter7));
  inv1  gate2515(.a(G1192), .O(gate460inter8));
  nand2 gate2516(.a(gate460inter8), .b(gate460inter7), .O(gate460inter9));
  nand2 gate2517(.a(s_281), .b(gate460inter3), .O(gate460inter10));
  nor2  gate2518(.a(gate460inter10), .b(gate460inter9), .O(gate460inter11));
  nor2  gate2519(.a(gate460inter11), .b(gate460inter6), .O(gate460inter12));
  nand2 gate2520(.a(gate460inter12), .b(gate460inter1), .O(G1269));
nand2 gate461( .a(G22), .b(G1195), .O(G1270) );

  xor2  gate3053(.a(G1195), .b(G1099), .O(gate462inter0));
  nand2 gate3054(.a(gate462inter0), .b(s_358), .O(gate462inter1));
  and2  gate3055(.a(G1195), .b(G1099), .O(gate462inter2));
  inv1  gate3056(.a(s_358), .O(gate462inter3));
  inv1  gate3057(.a(s_359), .O(gate462inter4));
  nand2 gate3058(.a(gate462inter4), .b(gate462inter3), .O(gate462inter5));
  nor2  gate3059(.a(gate462inter5), .b(gate462inter2), .O(gate462inter6));
  inv1  gate3060(.a(G1099), .O(gate462inter7));
  inv1  gate3061(.a(G1195), .O(gate462inter8));
  nand2 gate3062(.a(gate462inter8), .b(gate462inter7), .O(gate462inter9));
  nand2 gate3063(.a(s_359), .b(gate462inter3), .O(gate462inter10));
  nor2  gate3064(.a(gate462inter10), .b(gate462inter9), .O(gate462inter11));
  nor2  gate3065(.a(gate462inter11), .b(gate462inter6), .O(gate462inter12));
  nand2 gate3066(.a(gate462inter12), .b(gate462inter1), .O(G1271));
nand2 gate463( .a(G23), .b(G1198), .O(G1272) );
nand2 gate464( .a(G1102), .b(G1198), .O(G1273) );
nand2 gate465( .a(G24), .b(G1201), .O(G1274) );

  xor2  gate1471(.a(G1201), .b(G1105), .O(gate466inter0));
  nand2 gate1472(.a(gate466inter0), .b(s_132), .O(gate466inter1));
  and2  gate1473(.a(G1201), .b(G1105), .O(gate466inter2));
  inv1  gate1474(.a(s_132), .O(gate466inter3));
  inv1  gate1475(.a(s_133), .O(gate466inter4));
  nand2 gate1476(.a(gate466inter4), .b(gate466inter3), .O(gate466inter5));
  nor2  gate1477(.a(gate466inter5), .b(gate466inter2), .O(gate466inter6));
  inv1  gate1478(.a(G1105), .O(gate466inter7));
  inv1  gate1479(.a(G1201), .O(gate466inter8));
  nand2 gate1480(.a(gate466inter8), .b(gate466inter7), .O(gate466inter9));
  nand2 gate1481(.a(s_133), .b(gate466inter3), .O(gate466inter10));
  nor2  gate1482(.a(gate466inter10), .b(gate466inter9), .O(gate466inter11));
  nor2  gate1483(.a(gate466inter11), .b(gate466inter6), .O(gate466inter12));
  nand2 gate1484(.a(gate466inter12), .b(gate466inter1), .O(G1275));
nand2 gate467( .a(G25), .b(G1204), .O(G1276) );
nand2 gate468( .a(G1108), .b(G1204), .O(G1277) );
nand2 gate469( .a(G26), .b(G1207), .O(G1278) );

  xor2  gate1093(.a(G1207), .b(G1111), .O(gate470inter0));
  nand2 gate1094(.a(gate470inter0), .b(s_78), .O(gate470inter1));
  and2  gate1095(.a(G1207), .b(G1111), .O(gate470inter2));
  inv1  gate1096(.a(s_78), .O(gate470inter3));
  inv1  gate1097(.a(s_79), .O(gate470inter4));
  nand2 gate1098(.a(gate470inter4), .b(gate470inter3), .O(gate470inter5));
  nor2  gate1099(.a(gate470inter5), .b(gate470inter2), .O(gate470inter6));
  inv1  gate1100(.a(G1111), .O(gate470inter7));
  inv1  gate1101(.a(G1207), .O(gate470inter8));
  nand2 gate1102(.a(gate470inter8), .b(gate470inter7), .O(gate470inter9));
  nand2 gate1103(.a(s_79), .b(gate470inter3), .O(gate470inter10));
  nor2  gate1104(.a(gate470inter10), .b(gate470inter9), .O(gate470inter11));
  nor2  gate1105(.a(gate470inter11), .b(gate470inter6), .O(gate470inter12));
  nand2 gate1106(.a(gate470inter12), .b(gate470inter1), .O(G1279));
nand2 gate471( .a(G27), .b(G1210), .O(G1280) );
nand2 gate472( .a(G1114), .b(G1210), .O(G1281) );
nand2 gate473( .a(G28), .b(G1213), .O(G1282) );
nand2 gate474( .a(G1117), .b(G1213), .O(G1283) );
nand2 gate475( .a(G29), .b(G1216), .O(G1284) );
nand2 gate476( .a(G1120), .b(G1216), .O(G1285) );

  xor2  gate2269(.a(G1219), .b(G30), .O(gate477inter0));
  nand2 gate2270(.a(gate477inter0), .b(s_246), .O(gate477inter1));
  and2  gate2271(.a(G1219), .b(G30), .O(gate477inter2));
  inv1  gate2272(.a(s_246), .O(gate477inter3));
  inv1  gate2273(.a(s_247), .O(gate477inter4));
  nand2 gate2274(.a(gate477inter4), .b(gate477inter3), .O(gate477inter5));
  nor2  gate2275(.a(gate477inter5), .b(gate477inter2), .O(gate477inter6));
  inv1  gate2276(.a(G30), .O(gate477inter7));
  inv1  gate2277(.a(G1219), .O(gate477inter8));
  nand2 gate2278(.a(gate477inter8), .b(gate477inter7), .O(gate477inter9));
  nand2 gate2279(.a(s_247), .b(gate477inter3), .O(gate477inter10));
  nor2  gate2280(.a(gate477inter10), .b(gate477inter9), .O(gate477inter11));
  nor2  gate2281(.a(gate477inter11), .b(gate477inter6), .O(gate477inter12));
  nand2 gate2282(.a(gate477inter12), .b(gate477inter1), .O(G1286));

  xor2  gate2549(.a(G1219), .b(G1123), .O(gate478inter0));
  nand2 gate2550(.a(gate478inter0), .b(s_286), .O(gate478inter1));
  and2  gate2551(.a(G1219), .b(G1123), .O(gate478inter2));
  inv1  gate2552(.a(s_286), .O(gate478inter3));
  inv1  gate2553(.a(s_287), .O(gate478inter4));
  nand2 gate2554(.a(gate478inter4), .b(gate478inter3), .O(gate478inter5));
  nor2  gate2555(.a(gate478inter5), .b(gate478inter2), .O(gate478inter6));
  inv1  gate2556(.a(G1123), .O(gate478inter7));
  inv1  gate2557(.a(G1219), .O(gate478inter8));
  nand2 gate2558(.a(gate478inter8), .b(gate478inter7), .O(gate478inter9));
  nand2 gate2559(.a(s_287), .b(gate478inter3), .O(gate478inter10));
  nor2  gate2560(.a(gate478inter10), .b(gate478inter9), .O(gate478inter11));
  nor2  gate2561(.a(gate478inter11), .b(gate478inter6), .O(gate478inter12));
  nand2 gate2562(.a(gate478inter12), .b(gate478inter1), .O(G1287));
nand2 gate479( .a(G31), .b(G1222), .O(G1288) );
nand2 gate480( .a(G1126), .b(G1222), .O(G1289) );
nand2 gate481( .a(G32), .b(G1225), .O(G1290) );
nand2 gate482( .a(G1129), .b(G1225), .O(G1291) );
nand2 gate483( .a(G1228), .b(G1229), .O(G1292) );
nand2 gate484( .a(G1230), .b(G1231), .O(G1293) );

  xor2  gate1275(.a(G1233), .b(G1232), .O(gate485inter0));
  nand2 gate1276(.a(gate485inter0), .b(s_104), .O(gate485inter1));
  and2  gate1277(.a(G1233), .b(G1232), .O(gate485inter2));
  inv1  gate1278(.a(s_104), .O(gate485inter3));
  inv1  gate1279(.a(s_105), .O(gate485inter4));
  nand2 gate1280(.a(gate485inter4), .b(gate485inter3), .O(gate485inter5));
  nor2  gate1281(.a(gate485inter5), .b(gate485inter2), .O(gate485inter6));
  inv1  gate1282(.a(G1232), .O(gate485inter7));
  inv1  gate1283(.a(G1233), .O(gate485inter8));
  nand2 gate1284(.a(gate485inter8), .b(gate485inter7), .O(gate485inter9));
  nand2 gate1285(.a(s_105), .b(gate485inter3), .O(gate485inter10));
  nor2  gate1286(.a(gate485inter10), .b(gate485inter9), .O(gate485inter11));
  nor2  gate1287(.a(gate485inter11), .b(gate485inter6), .O(gate485inter12));
  nand2 gate1288(.a(gate485inter12), .b(gate485inter1), .O(G1294));
nand2 gate486( .a(G1234), .b(G1235), .O(G1295) );
nand2 gate487( .a(G1236), .b(G1237), .O(G1296) );
nand2 gate488( .a(G1238), .b(G1239), .O(G1297) );
nand2 gate489( .a(G1240), .b(G1241), .O(G1298) );
nand2 gate490( .a(G1242), .b(G1243), .O(G1299) );

  xor2  gate1163(.a(G1245), .b(G1244), .O(gate491inter0));
  nand2 gate1164(.a(gate491inter0), .b(s_88), .O(gate491inter1));
  and2  gate1165(.a(G1245), .b(G1244), .O(gate491inter2));
  inv1  gate1166(.a(s_88), .O(gate491inter3));
  inv1  gate1167(.a(s_89), .O(gate491inter4));
  nand2 gate1168(.a(gate491inter4), .b(gate491inter3), .O(gate491inter5));
  nor2  gate1169(.a(gate491inter5), .b(gate491inter2), .O(gate491inter6));
  inv1  gate1170(.a(G1244), .O(gate491inter7));
  inv1  gate1171(.a(G1245), .O(gate491inter8));
  nand2 gate1172(.a(gate491inter8), .b(gate491inter7), .O(gate491inter9));
  nand2 gate1173(.a(s_89), .b(gate491inter3), .O(gate491inter10));
  nor2  gate1174(.a(gate491inter10), .b(gate491inter9), .O(gate491inter11));
  nor2  gate1175(.a(gate491inter11), .b(gate491inter6), .O(gate491inter12));
  nand2 gate1176(.a(gate491inter12), .b(gate491inter1), .O(G1300));

  xor2  gate1247(.a(G1247), .b(G1246), .O(gate492inter0));
  nand2 gate1248(.a(gate492inter0), .b(s_100), .O(gate492inter1));
  and2  gate1249(.a(G1247), .b(G1246), .O(gate492inter2));
  inv1  gate1250(.a(s_100), .O(gate492inter3));
  inv1  gate1251(.a(s_101), .O(gate492inter4));
  nand2 gate1252(.a(gate492inter4), .b(gate492inter3), .O(gate492inter5));
  nor2  gate1253(.a(gate492inter5), .b(gate492inter2), .O(gate492inter6));
  inv1  gate1254(.a(G1246), .O(gate492inter7));
  inv1  gate1255(.a(G1247), .O(gate492inter8));
  nand2 gate1256(.a(gate492inter8), .b(gate492inter7), .O(gate492inter9));
  nand2 gate1257(.a(s_101), .b(gate492inter3), .O(gate492inter10));
  nor2  gate1258(.a(gate492inter10), .b(gate492inter9), .O(gate492inter11));
  nor2  gate1259(.a(gate492inter11), .b(gate492inter6), .O(gate492inter12));
  nand2 gate1260(.a(gate492inter12), .b(gate492inter1), .O(G1301));
nand2 gate493( .a(G1248), .b(G1249), .O(G1302) );

  xor2  gate1821(.a(G1251), .b(G1250), .O(gate494inter0));
  nand2 gate1822(.a(gate494inter0), .b(s_182), .O(gate494inter1));
  and2  gate1823(.a(G1251), .b(G1250), .O(gate494inter2));
  inv1  gate1824(.a(s_182), .O(gate494inter3));
  inv1  gate1825(.a(s_183), .O(gate494inter4));
  nand2 gate1826(.a(gate494inter4), .b(gate494inter3), .O(gate494inter5));
  nor2  gate1827(.a(gate494inter5), .b(gate494inter2), .O(gate494inter6));
  inv1  gate1828(.a(G1250), .O(gate494inter7));
  inv1  gate1829(.a(G1251), .O(gate494inter8));
  nand2 gate1830(.a(gate494inter8), .b(gate494inter7), .O(gate494inter9));
  nand2 gate1831(.a(s_183), .b(gate494inter3), .O(gate494inter10));
  nor2  gate1832(.a(gate494inter10), .b(gate494inter9), .O(gate494inter11));
  nor2  gate1833(.a(gate494inter11), .b(gate494inter6), .O(gate494inter12));
  nand2 gate1834(.a(gate494inter12), .b(gate494inter1), .O(G1303));
nand2 gate495( .a(G1252), .b(G1253), .O(G1304) );
nand2 gate496( .a(G1254), .b(G1255), .O(G1305) );

  xor2  gate2717(.a(G1257), .b(G1256), .O(gate497inter0));
  nand2 gate2718(.a(gate497inter0), .b(s_310), .O(gate497inter1));
  and2  gate2719(.a(G1257), .b(G1256), .O(gate497inter2));
  inv1  gate2720(.a(s_310), .O(gate497inter3));
  inv1  gate2721(.a(s_311), .O(gate497inter4));
  nand2 gate2722(.a(gate497inter4), .b(gate497inter3), .O(gate497inter5));
  nor2  gate2723(.a(gate497inter5), .b(gate497inter2), .O(gate497inter6));
  inv1  gate2724(.a(G1256), .O(gate497inter7));
  inv1  gate2725(.a(G1257), .O(gate497inter8));
  nand2 gate2726(.a(gate497inter8), .b(gate497inter7), .O(gate497inter9));
  nand2 gate2727(.a(s_311), .b(gate497inter3), .O(gate497inter10));
  nor2  gate2728(.a(gate497inter10), .b(gate497inter9), .O(gate497inter11));
  nor2  gate2729(.a(gate497inter11), .b(gate497inter6), .O(gate497inter12));
  nand2 gate2730(.a(gate497inter12), .b(gate497inter1), .O(G1306));

  xor2  gate3067(.a(G1259), .b(G1258), .O(gate498inter0));
  nand2 gate3068(.a(gate498inter0), .b(s_360), .O(gate498inter1));
  and2  gate3069(.a(G1259), .b(G1258), .O(gate498inter2));
  inv1  gate3070(.a(s_360), .O(gate498inter3));
  inv1  gate3071(.a(s_361), .O(gate498inter4));
  nand2 gate3072(.a(gate498inter4), .b(gate498inter3), .O(gate498inter5));
  nor2  gate3073(.a(gate498inter5), .b(gate498inter2), .O(gate498inter6));
  inv1  gate3074(.a(G1258), .O(gate498inter7));
  inv1  gate3075(.a(G1259), .O(gate498inter8));
  nand2 gate3076(.a(gate498inter8), .b(gate498inter7), .O(gate498inter9));
  nand2 gate3077(.a(s_361), .b(gate498inter3), .O(gate498inter10));
  nor2  gate3078(.a(gate498inter10), .b(gate498inter9), .O(gate498inter11));
  nor2  gate3079(.a(gate498inter11), .b(gate498inter6), .O(gate498inter12));
  nand2 gate3080(.a(gate498inter12), .b(gate498inter1), .O(G1307));

  xor2  gate1177(.a(G1261), .b(G1260), .O(gate499inter0));
  nand2 gate1178(.a(gate499inter0), .b(s_90), .O(gate499inter1));
  and2  gate1179(.a(G1261), .b(G1260), .O(gate499inter2));
  inv1  gate1180(.a(s_90), .O(gate499inter3));
  inv1  gate1181(.a(s_91), .O(gate499inter4));
  nand2 gate1182(.a(gate499inter4), .b(gate499inter3), .O(gate499inter5));
  nor2  gate1183(.a(gate499inter5), .b(gate499inter2), .O(gate499inter6));
  inv1  gate1184(.a(G1260), .O(gate499inter7));
  inv1  gate1185(.a(G1261), .O(gate499inter8));
  nand2 gate1186(.a(gate499inter8), .b(gate499inter7), .O(gate499inter9));
  nand2 gate1187(.a(s_91), .b(gate499inter3), .O(gate499inter10));
  nor2  gate1188(.a(gate499inter10), .b(gate499inter9), .O(gate499inter11));
  nor2  gate1189(.a(gate499inter11), .b(gate499inter6), .O(gate499inter12));
  nand2 gate1190(.a(gate499inter12), .b(gate499inter1), .O(G1308));
nand2 gate500( .a(G1262), .b(G1263), .O(G1309) );
nand2 gate501( .a(G1264), .b(G1265), .O(G1310) );

  xor2  gate2185(.a(G1267), .b(G1266), .O(gate502inter0));
  nand2 gate2186(.a(gate502inter0), .b(s_234), .O(gate502inter1));
  and2  gate2187(.a(G1267), .b(G1266), .O(gate502inter2));
  inv1  gate2188(.a(s_234), .O(gate502inter3));
  inv1  gate2189(.a(s_235), .O(gate502inter4));
  nand2 gate2190(.a(gate502inter4), .b(gate502inter3), .O(gate502inter5));
  nor2  gate2191(.a(gate502inter5), .b(gate502inter2), .O(gate502inter6));
  inv1  gate2192(.a(G1266), .O(gate502inter7));
  inv1  gate2193(.a(G1267), .O(gate502inter8));
  nand2 gate2194(.a(gate502inter8), .b(gate502inter7), .O(gate502inter9));
  nand2 gate2195(.a(s_235), .b(gate502inter3), .O(gate502inter10));
  nor2  gate2196(.a(gate502inter10), .b(gate502inter9), .O(gate502inter11));
  nor2  gate2197(.a(gate502inter11), .b(gate502inter6), .O(gate502inter12));
  nand2 gate2198(.a(gate502inter12), .b(gate502inter1), .O(G1311));
nand2 gate503( .a(G1268), .b(G1269), .O(G1312) );

  xor2  gate1863(.a(G1271), .b(G1270), .O(gate504inter0));
  nand2 gate1864(.a(gate504inter0), .b(s_188), .O(gate504inter1));
  and2  gate1865(.a(G1271), .b(G1270), .O(gate504inter2));
  inv1  gate1866(.a(s_188), .O(gate504inter3));
  inv1  gate1867(.a(s_189), .O(gate504inter4));
  nand2 gate1868(.a(gate504inter4), .b(gate504inter3), .O(gate504inter5));
  nor2  gate1869(.a(gate504inter5), .b(gate504inter2), .O(gate504inter6));
  inv1  gate1870(.a(G1270), .O(gate504inter7));
  inv1  gate1871(.a(G1271), .O(gate504inter8));
  nand2 gate1872(.a(gate504inter8), .b(gate504inter7), .O(gate504inter9));
  nand2 gate1873(.a(s_189), .b(gate504inter3), .O(gate504inter10));
  nor2  gate1874(.a(gate504inter10), .b(gate504inter9), .O(gate504inter11));
  nor2  gate1875(.a(gate504inter11), .b(gate504inter6), .O(gate504inter12));
  nand2 gate1876(.a(gate504inter12), .b(gate504inter1), .O(G1313));

  xor2  gate2059(.a(G1273), .b(G1272), .O(gate505inter0));
  nand2 gate2060(.a(gate505inter0), .b(s_216), .O(gate505inter1));
  and2  gate2061(.a(G1273), .b(G1272), .O(gate505inter2));
  inv1  gate2062(.a(s_216), .O(gate505inter3));
  inv1  gate2063(.a(s_217), .O(gate505inter4));
  nand2 gate2064(.a(gate505inter4), .b(gate505inter3), .O(gate505inter5));
  nor2  gate2065(.a(gate505inter5), .b(gate505inter2), .O(gate505inter6));
  inv1  gate2066(.a(G1272), .O(gate505inter7));
  inv1  gate2067(.a(G1273), .O(gate505inter8));
  nand2 gate2068(.a(gate505inter8), .b(gate505inter7), .O(gate505inter9));
  nand2 gate2069(.a(s_217), .b(gate505inter3), .O(gate505inter10));
  nor2  gate2070(.a(gate505inter10), .b(gate505inter9), .O(gate505inter11));
  nor2  gate2071(.a(gate505inter11), .b(gate505inter6), .O(gate505inter12));
  nand2 gate2072(.a(gate505inter12), .b(gate505inter1), .O(G1314));
nand2 gate506( .a(G1274), .b(G1275), .O(G1315) );

  xor2  gate1835(.a(G1277), .b(G1276), .O(gate507inter0));
  nand2 gate1836(.a(gate507inter0), .b(s_184), .O(gate507inter1));
  and2  gate1837(.a(G1277), .b(G1276), .O(gate507inter2));
  inv1  gate1838(.a(s_184), .O(gate507inter3));
  inv1  gate1839(.a(s_185), .O(gate507inter4));
  nand2 gate1840(.a(gate507inter4), .b(gate507inter3), .O(gate507inter5));
  nor2  gate1841(.a(gate507inter5), .b(gate507inter2), .O(gate507inter6));
  inv1  gate1842(.a(G1276), .O(gate507inter7));
  inv1  gate1843(.a(G1277), .O(gate507inter8));
  nand2 gate1844(.a(gate507inter8), .b(gate507inter7), .O(gate507inter9));
  nand2 gate1845(.a(s_185), .b(gate507inter3), .O(gate507inter10));
  nor2  gate1846(.a(gate507inter10), .b(gate507inter9), .O(gate507inter11));
  nor2  gate1847(.a(gate507inter11), .b(gate507inter6), .O(gate507inter12));
  nand2 gate1848(.a(gate507inter12), .b(gate507inter1), .O(G1316));

  xor2  gate3095(.a(G1279), .b(G1278), .O(gate508inter0));
  nand2 gate3096(.a(gate508inter0), .b(s_364), .O(gate508inter1));
  and2  gate3097(.a(G1279), .b(G1278), .O(gate508inter2));
  inv1  gate3098(.a(s_364), .O(gate508inter3));
  inv1  gate3099(.a(s_365), .O(gate508inter4));
  nand2 gate3100(.a(gate508inter4), .b(gate508inter3), .O(gate508inter5));
  nor2  gate3101(.a(gate508inter5), .b(gate508inter2), .O(gate508inter6));
  inv1  gate3102(.a(G1278), .O(gate508inter7));
  inv1  gate3103(.a(G1279), .O(gate508inter8));
  nand2 gate3104(.a(gate508inter8), .b(gate508inter7), .O(gate508inter9));
  nand2 gate3105(.a(s_365), .b(gate508inter3), .O(gate508inter10));
  nor2  gate3106(.a(gate508inter10), .b(gate508inter9), .O(gate508inter11));
  nor2  gate3107(.a(gate508inter11), .b(gate508inter6), .O(gate508inter12));
  nand2 gate3108(.a(gate508inter12), .b(gate508inter1), .O(G1317));
nand2 gate509( .a(G1280), .b(G1281), .O(G1318) );
nand2 gate510( .a(G1282), .b(G1283), .O(G1319) );

  xor2  gate1933(.a(G1285), .b(G1284), .O(gate511inter0));
  nand2 gate1934(.a(gate511inter0), .b(s_198), .O(gate511inter1));
  and2  gate1935(.a(G1285), .b(G1284), .O(gate511inter2));
  inv1  gate1936(.a(s_198), .O(gate511inter3));
  inv1  gate1937(.a(s_199), .O(gate511inter4));
  nand2 gate1938(.a(gate511inter4), .b(gate511inter3), .O(gate511inter5));
  nor2  gate1939(.a(gate511inter5), .b(gate511inter2), .O(gate511inter6));
  inv1  gate1940(.a(G1284), .O(gate511inter7));
  inv1  gate1941(.a(G1285), .O(gate511inter8));
  nand2 gate1942(.a(gate511inter8), .b(gate511inter7), .O(gate511inter9));
  nand2 gate1943(.a(s_199), .b(gate511inter3), .O(gate511inter10));
  nor2  gate1944(.a(gate511inter10), .b(gate511inter9), .O(gate511inter11));
  nor2  gate1945(.a(gate511inter11), .b(gate511inter6), .O(gate511inter12));
  nand2 gate1946(.a(gate511inter12), .b(gate511inter1), .O(G1320));

  xor2  gate2479(.a(G1287), .b(G1286), .O(gate512inter0));
  nand2 gate2480(.a(gate512inter0), .b(s_276), .O(gate512inter1));
  and2  gate2481(.a(G1287), .b(G1286), .O(gate512inter2));
  inv1  gate2482(.a(s_276), .O(gate512inter3));
  inv1  gate2483(.a(s_277), .O(gate512inter4));
  nand2 gate2484(.a(gate512inter4), .b(gate512inter3), .O(gate512inter5));
  nor2  gate2485(.a(gate512inter5), .b(gate512inter2), .O(gate512inter6));
  inv1  gate2486(.a(G1286), .O(gate512inter7));
  inv1  gate2487(.a(G1287), .O(gate512inter8));
  nand2 gate2488(.a(gate512inter8), .b(gate512inter7), .O(gate512inter9));
  nand2 gate2489(.a(s_277), .b(gate512inter3), .O(gate512inter10));
  nor2  gate2490(.a(gate512inter10), .b(gate512inter9), .O(gate512inter11));
  nor2  gate2491(.a(gate512inter11), .b(gate512inter6), .O(gate512inter12));
  nand2 gate2492(.a(gate512inter12), .b(gate512inter1), .O(G1321));
nand2 gate513( .a(G1288), .b(G1289), .O(G1322) );
nand2 gate514( .a(G1290), .b(G1291), .O(G1323) );
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule