module c499 (N1,N5,N9,N13,N17,N21,N25,N29,N33,N37,
             N41,N45,N49,N53,N57,N61,N65,N69,N73,N77,
             N81,N85,N89,N93,N97,N101,N105,N109,N113,N117,
             N121,N125,N129,N130,N131,N132,N133,N134,N135,N136,
             N137,N724,N725,N726,N727,N728,N729,N730,N731,N732,
             N733,N734,N735,N736,N737,N738,N739,N740,N741,N742,
             N743,N744,N745,N746,N747,N748,N749,N750,N751,N752,
             N753,N754,N755);

input N1,N5,N9,N13,N17,N21,N25,N29,N33,N37,
      N41,N45,N49,N53,N57,N61,N65,N69,N73,N77,
      N81,N85,N89,N93,N97,N101,N105,N109,N113,N117,
      N121,N125,N129,N130,N131,N132,N133,N134,N135,N136,
      N137;//RE__PI;

input s_0,s_1;//RE__ALLOW(00,01,10,11);
input s_2,s_3;//RE__ALLOW(00,01,10,11);
input s_4,s_5;//RE__ALLOW(00,01,10,11);
input s_6,s_7;//RE__ALLOW(00,01,10,11);
input s_8,s_9;//RE__ALLOW(00,01,10,11);
input s_10,s_11;//RE__ALLOW(00,01,10,11);
input s_12,s_13;//RE__ALLOW(00,01,10,11);
input s_14,s_15;//RE__ALLOW(00,01,10,11);
input s_16,s_17;//RE__ALLOW(00,01,10,11);
input s_18,s_19;//RE__ALLOW(00,01,10,11);
input s_20,s_21;//RE__ALLOW(00,01,10,11);
input s_22,s_23;//RE__ALLOW(00,01,10,11);
input s_24,s_25;//RE__ALLOW(00,01,10,11);
input s_26,s_27;//RE__ALLOW(00,01,10,11);
input s_28,s_29;//RE__ALLOW(00,01,10,11);
input s_30,s_31;//RE__ALLOW(00,01,10,11);
input s_32,s_33;//RE__ALLOW(00,01,10,11);
input s_34,s_35;//RE__ALLOW(00,01,10,11);
input s_36,s_37;//RE__ALLOW(00,01,10,11);
input s_38,s_39;//RE__ALLOW(00,01,10,11);
input s_40,s_41;//RE__ALLOW(00,01,10,11);
output N724,N725,N726,N727,N728,N729,N730,N731,N732,N733,
       N734,N735,N736,N737,N738,N739,N740,N741,N742,N743,
       N744,N745,N746,N747,N748,N749,N750,N751,N752,N753,
       N754,N755;

wire N250,N251,N252,N253,N254,N255,N256,N257,N258,N259,
     N260,N261,N262,N263,N264,N265,N266,N267,N268,N269,
     N270,N271,N272,N273,N274,N275,N276,N277,N278,N279,
     N280,N281,N282,N283,N284,N285,N286,N287,N288,N289,
     N290,N293,N296,N299,N302,N305,N308,N311,N314,N315,
     N316,N317,N318,N319,N320,N321,N338,N339,N340,N341,
     N342,N343,N344,N345,N346,N347,N348,N349,N350,N351,
     N352,N353,N354,N367,N380,N393,N406,N419,N432,N445,
     N554,N555,N556,N557,N558,N559,N560,N561,N562,N563,
     N564,N565,N566,N567,N568,N569,N570,N571,N572,N573,
     N574,N575,N576,N577,N578,N579,N580,N581,N582,N583,
     N584,N585,N586,N587,N588,N589,N590,N591,N592,N593,
     N594,N595,N596,N597,N598,N599,N600,N601,N602,N607,
     N620,N625,N630,N635,N640,N645,N650,N655,N692,N693,
     N694,N695,N696,N697,N698,N699,N700,N701,N702,N703,
     N704,N705,N706,N707,N708,N709,N710,N711,N712,N713,
     N714,N715,N716,N717,N718,N719,N720,N721,N722,N723, gate42inter0, gate42inter1, gate42inter2, gate42inter3, gate42inter4, gate42inter5, gate42inter6, gate42inter7, gate42inter8, gate42inter9, gate42inter10, gate42inter11, gate42inter12, gate79inter0, gate79inter1, gate79inter2, gate79inter3, gate79inter4, gate79inter5, gate79inter6, gate79inter7, gate79inter8, gate79inter9, gate79inter10, gate79inter11, gate79inter12, gate63inter0, gate63inter1, gate63inter2, gate63inter3, gate63inter4, gate63inter5, gate63inter6, gate63inter7, gate63inter8, gate63inter9, gate63inter10, gate63inter11, gate63inter12, gate176inter0, gate176inter1, gate176inter2, gate176inter3, gate176inter4, gate176inter5, gate176inter6, gate176inter7, gate176inter8, gate176inter9, gate176inter10, gate176inter11, gate176inter12, gate181inter0, gate181inter1, gate181inter2, gate181inter3, gate181inter4, gate181inter5, gate181inter6, gate181inter7, gate181inter8, gate181inter9, gate181inter10, gate181inter11, gate181inter12, gate188inter0, gate188inter1, gate188inter2, gate188inter3, gate188inter4, gate188inter5, gate188inter6, gate188inter7, gate188inter8, gate188inter9, gate188inter10, gate188inter11, gate188inter12, gate55inter0, gate55inter1, gate55inter2, gate55inter3, gate55inter4, gate55inter5, gate55inter6, gate55inter7, gate55inter8, gate55inter9, gate55inter10, gate55inter11, gate55inter12, gate31inter0, gate31inter1, gate31inter2, gate31inter3, gate31inter4, gate31inter5, gate31inter6, gate31inter7, gate31inter8, gate31inter9, gate31inter10, gate31inter11, gate31inter12, gate197inter0, gate197inter1, gate197inter2, gate197inter3, gate197inter4, gate197inter5, gate197inter6, gate197inter7, gate197inter8, gate197inter9, gate197inter10, gate197inter11, gate197inter12, gate2inter0, gate2inter1, gate2inter2, gate2inter3, gate2inter4, gate2inter5, gate2inter6, gate2inter7, gate2inter8, gate2inter9, gate2inter10, gate2inter11, gate2inter12, gate186inter0, gate186inter1, gate186inter2, gate186inter3, gate186inter4, gate186inter5, gate186inter6, gate186inter7, gate186inter8, gate186inter9, gate186inter10, gate186inter11, gate186inter12, gate52inter0, gate52inter1, gate52inter2, gate52inter3, gate52inter4, gate52inter5, gate52inter6, gate52inter7, gate52inter8, gate52inter9, gate52inter10, gate52inter11, gate52inter12, gate45inter0, gate45inter1, gate45inter2, gate45inter3, gate45inter4, gate45inter5, gate45inter6, gate45inter7, gate45inter8, gate45inter9, gate45inter10, gate45inter11, gate45inter12, gate200inter0, gate200inter1, gate200inter2, gate200inter3, gate200inter4, gate200inter5, gate200inter6, gate200inter7, gate200inter8, gate200inter9, gate200inter10, gate200inter11, gate200inter12, gate173inter0, gate173inter1, gate173inter2, gate173inter3, gate173inter4, gate173inter5, gate173inter6, gate173inter7, gate173inter8, gate173inter9, gate173inter10, gate173inter11, gate173inter12, gate27inter0, gate27inter1, gate27inter2, gate27inter3, gate27inter4, gate27inter5, gate27inter6, gate27inter7, gate27inter8, gate27inter9, gate27inter10, gate27inter11, gate27inter12, gate187inter0, gate187inter1, gate187inter2, gate187inter3, gate187inter4, gate187inter5, gate187inter6, gate187inter7, gate187inter8, gate187inter9, gate187inter10, gate187inter11, gate187inter12, gate49inter0, gate49inter1, gate49inter2, gate49inter3, gate49inter4, gate49inter5, gate49inter6, gate49inter7, gate49inter8, gate49inter9, gate49inter10, gate49inter11, gate49inter12, gate71inter0, gate71inter1, gate71inter2, gate71inter3, gate71inter4, gate71inter5, gate71inter6, gate71inter7, gate71inter8, gate71inter9, gate71inter10, gate71inter11, gate71inter12, gate178inter0, gate178inter1, gate178inter2, gate178inter3, gate178inter4, gate178inter5, gate178inter6, gate178inter7, gate178inter8, gate178inter9, gate178inter10, gate178inter11, gate178inter12, gate61inter0, gate61inter1, gate61inter2, gate61inter3, gate61inter4, gate61inter5, gate61inter6, gate61inter7, gate61inter8, gate61inter9, gate61inter10, gate61inter11, gate61inter12;



xor2 gate1( .a(N1), .b(N5), .O(N250) );

  xor2  gate329(.a(N13), .b(N9), .O(gate2inter0));
  nand2 gate330(.a(gate2inter0), .b(s_18), .O(gate2inter1));
  and2  gate331(.a(N13), .b(N9), .O(gate2inter2));
  inv1  gate332(.a(s_18), .O(gate2inter3));
  inv1  gate333(.a(s_19), .O(gate2inter4));
  nand2 gate334(.a(gate2inter4), .b(gate2inter3), .O(gate2inter5));
  nor2  gate335(.a(gate2inter5), .b(gate2inter2), .O(gate2inter6));
  inv1  gate336(.a(N9), .O(gate2inter7));
  inv1  gate337(.a(N13), .O(gate2inter8));
  nand2 gate338(.a(gate2inter8), .b(gate2inter7), .O(gate2inter9));
  nand2 gate339(.a(s_19), .b(gate2inter3), .O(gate2inter10));
  nor2  gate340(.a(gate2inter10), .b(gate2inter9), .O(gate2inter11));
  nor2  gate341(.a(gate2inter11), .b(gate2inter6), .O(gate2inter12));
  nand2 gate342(.a(gate2inter12), .b(gate2inter1), .O(N251));
xor2 gate3( .a(N17), .b(N21), .O(N252) );
xor2 gate4( .a(N25), .b(N29), .O(N253) );
xor2 gate5( .a(N33), .b(N37), .O(N254) );
xor2 gate6( .a(N41), .b(N45), .O(N255) );
xor2 gate7( .a(N49), .b(N53), .O(N256) );
xor2 gate8( .a(N57), .b(N61), .O(N257) );
xor2 gate9( .a(N65), .b(N69), .O(N258) );
xor2 gate10( .a(N73), .b(N77), .O(N259) );
xor2 gate11( .a(N81), .b(N85), .O(N260) );
xor2 gate12( .a(N89), .b(N93), .O(N261) );
xor2 gate13( .a(N97), .b(N101), .O(N262) );
xor2 gate14( .a(N105), .b(N109), .O(N263) );
xor2 gate15( .a(N113), .b(N117), .O(N264) );
xor2 gate16( .a(N121), .b(N125), .O(N265) );
and2 gate17( .a(N129), .b(N137), .O(N266) );
and2 gate18( .a(N130), .b(N137), .O(N267) );
and2 gate19( .a(N131), .b(N137), .O(N268) );
and2 gate20( .a(N132), .b(N137), .O(N269) );
and2 gate21( .a(N133), .b(N137), .O(N270) );
and2 gate22( .a(N134), .b(N137), .O(N271) );
and2 gate23( .a(N135), .b(N137), .O(N272) );
and2 gate24( .a(N136), .b(N137), .O(N273) );
xor2 gate25( .a(N1), .b(N17), .O(N274) );
xor2 gate26( .a(N33), .b(N49), .O(N275) );

  xor2  gate413(.a(N21), .b(N5), .O(gate27inter0));
  nand2 gate414(.a(gate27inter0), .b(s_30), .O(gate27inter1));
  and2  gate415(.a(N21), .b(N5), .O(gate27inter2));
  inv1  gate416(.a(s_30), .O(gate27inter3));
  inv1  gate417(.a(s_31), .O(gate27inter4));
  nand2 gate418(.a(gate27inter4), .b(gate27inter3), .O(gate27inter5));
  nor2  gate419(.a(gate27inter5), .b(gate27inter2), .O(gate27inter6));
  inv1  gate420(.a(N5), .O(gate27inter7));
  inv1  gate421(.a(N21), .O(gate27inter8));
  nand2 gate422(.a(gate27inter8), .b(gate27inter7), .O(gate27inter9));
  nand2 gate423(.a(s_31), .b(gate27inter3), .O(gate27inter10));
  nor2  gate424(.a(gate27inter10), .b(gate27inter9), .O(gate27inter11));
  nor2  gate425(.a(gate27inter11), .b(gate27inter6), .O(gate27inter12));
  nand2 gate426(.a(gate27inter12), .b(gate27inter1), .O(N276));
xor2 gate28( .a(N37), .b(N53), .O(N277) );
xor2 gate29( .a(N9), .b(N25), .O(N278) );
xor2 gate30( .a(N41), .b(N57), .O(N279) );

  xor2  gate301(.a(N29), .b(N13), .O(gate31inter0));
  nand2 gate302(.a(gate31inter0), .b(s_14), .O(gate31inter1));
  and2  gate303(.a(N29), .b(N13), .O(gate31inter2));
  inv1  gate304(.a(s_14), .O(gate31inter3));
  inv1  gate305(.a(s_15), .O(gate31inter4));
  nand2 gate306(.a(gate31inter4), .b(gate31inter3), .O(gate31inter5));
  nor2  gate307(.a(gate31inter5), .b(gate31inter2), .O(gate31inter6));
  inv1  gate308(.a(N13), .O(gate31inter7));
  inv1  gate309(.a(N29), .O(gate31inter8));
  nand2 gate310(.a(gate31inter8), .b(gate31inter7), .O(gate31inter9));
  nand2 gate311(.a(s_15), .b(gate31inter3), .O(gate31inter10));
  nor2  gate312(.a(gate31inter10), .b(gate31inter9), .O(gate31inter11));
  nor2  gate313(.a(gate31inter11), .b(gate31inter6), .O(gate31inter12));
  nand2 gate314(.a(gate31inter12), .b(gate31inter1), .O(N280));
xor2 gate32( .a(N45), .b(N61), .O(N281) );
xor2 gate33( .a(N65), .b(N81), .O(N282) );
xor2 gate34( .a(N97), .b(N113), .O(N283) );
xor2 gate35( .a(N69), .b(N85), .O(N284) );
xor2 gate36( .a(N101), .b(N117), .O(N285) );
xor2 gate37( .a(N73), .b(N89), .O(N286) );
xor2 gate38( .a(N105), .b(N121), .O(N287) );
xor2 gate39( .a(N77), .b(N93), .O(N288) );
xor2 gate40( .a(N109), .b(N125), .O(N289) );
xor2 gate41( .a(N250), .b(N251), .O(N290) );

  xor2  gate203(.a(N253), .b(N252), .O(gate42inter0));
  nand2 gate204(.a(gate42inter0), .b(s_0), .O(gate42inter1));
  and2  gate205(.a(N253), .b(N252), .O(gate42inter2));
  inv1  gate206(.a(s_0), .O(gate42inter3));
  inv1  gate207(.a(s_1), .O(gate42inter4));
  nand2 gate208(.a(gate42inter4), .b(gate42inter3), .O(gate42inter5));
  nor2  gate209(.a(gate42inter5), .b(gate42inter2), .O(gate42inter6));
  inv1  gate210(.a(N252), .O(gate42inter7));
  inv1  gate211(.a(N253), .O(gate42inter8));
  nand2 gate212(.a(gate42inter8), .b(gate42inter7), .O(gate42inter9));
  nand2 gate213(.a(s_1), .b(gate42inter3), .O(gate42inter10));
  nor2  gate214(.a(gate42inter10), .b(gate42inter9), .O(gate42inter11));
  nor2  gate215(.a(gate42inter11), .b(gate42inter6), .O(gate42inter12));
  nand2 gate216(.a(gate42inter12), .b(gate42inter1), .O(N293));
xor2 gate43( .a(N254), .b(N255), .O(N296) );
xor2 gate44( .a(N256), .b(N257), .O(N299) );

  xor2  gate371(.a(N259), .b(N258), .O(gate45inter0));
  nand2 gate372(.a(gate45inter0), .b(s_24), .O(gate45inter1));
  and2  gate373(.a(N259), .b(N258), .O(gate45inter2));
  inv1  gate374(.a(s_24), .O(gate45inter3));
  inv1  gate375(.a(s_25), .O(gate45inter4));
  nand2 gate376(.a(gate45inter4), .b(gate45inter3), .O(gate45inter5));
  nor2  gate377(.a(gate45inter5), .b(gate45inter2), .O(gate45inter6));
  inv1  gate378(.a(N258), .O(gate45inter7));
  inv1  gate379(.a(N259), .O(gate45inter8));
  nand2 gate380(.a(gate45inter8), .b(gate45inter7), .O(gate45inter9));
  nand2 gate381(.a(s_25), .b(gate45inter3), .O(gate45inter10));
  nor2  gate382(.a(gate45inter10), .b(gate45inter9), .O(gate45inter11));
  nor2  gate383(.a(gate45inter11), .b(gate45inter6), .O(gate45inter12));
  nand2 gate384(.a(gate45inter12), .b(gate45inter1), .O(N302));
xor2 gate46( .a(N260), .b(N261), .O(N305) );
xor2 gate47( .a(N262), .b(N263), .O(N308) );
xor2 gate48( .a(N264), .b(N265), .O(N311) );

  xor2  gate441(.a(N275), .b(N274), .O(gate49inter0));
  nand2 gate442(.a(gate49inter0), .b(s_34), .O(gate49inter1));
  and2  gate443(.a(N275), .b(N274), .O(gate49inter2));
  inv1  gate444(.a(s_34), .O(gate49inter3));
  inv1  gate445(.a(s_35), .O(gate49inter4));
  nand2 gate446(.a(gate49inter4), .b(gate49inter3), .O(gate49inter5));
  nor2  gate447(.a(gate49inter5), .b(gate49inter2), .O(gate49inter6));
  inv1  gate448(.a(N274), .O(gate49inter7));
  inv1  gate449(.a(N275), .O(gate49inter8));
  nand2 gate450(.a(gate49inter8), .b(gate49inter7), .O(gate49inter9));
  nand2 gate451(.a(s_35), .b(gate49inter3), .O(gate49inter10));
  nor2  gate452(.a(gate49inter10), .b(gate49inter9), .O(gate49inter11));
  nor2  gate453(.a(gate49inter11), .b(gate49inter6), .O(gate49inter12));
  nand2 gate454(.a(gate49inter12), .b(gate49inter1), .O(N314));
xor2 gate50( .a(N276), .b(N277), .O(N315) );
xor2 gate51( .a(N278), .b(N279), .O(N316) );

  xor2  gate357(.a(N281), .b(N280), .O(gate52inter0));
  nand2 gate358(.a(gate52inter0), .b(s_22), .O(gate52inter1));
  and2  gate359(.a(N281), .b(N280), .O(gate52inter2));
  inv1  gate360(.a(s_22), .O(gate52inter3));
  inv1  gate361(.a(s_23), .O(gate52inter4));
  nand2 gate362(.a(gate52inter4), .b(gate52inter3), .O(gate52inter5));
  nor2  gate363(.a(gate52inter5), .b(gate52inter2), .O(gate52inter6));
  inv1  gate364(.a(N280), .O(gate52inter7));
  inv1  gate365(.a(N281), .O(gate52inter8));
  nand2 gate366(.a(gate52inter8), .b(gate52inter7), .O(gate52inter9));
  nand2 gate367(.a(s_23), .b(gate52inter3), .O(gate52inter10));
  nor2  gate368(.a(gate52inter10), .b(gate52inter9), .O(gate52inter11));
  nor2  gate369(.a(gate52inter11), .b(gate52inter6), .O(gate52inter12));
  nand2 gate370(.a(gate52inter12), .b(gate52inter1), .O(N317));
xor2 gate53( .a(N282), .b(N283), .O(N318) );
xor2 gate54( .a(N284), .b(N285), .O(N319) );

  xor2  gate287(.a(N287), .b(N286), .O(gate55inter0));
  nand2 gate288(.a(gate55inter0), .b(s_12), .O(gate55inter1));
  and2  gate289(.a(N287), .b(N286), .O(gate55inter2));
  inv1  gate290(.a(s_12), .O(gate55inter3));
  inv1  gate291(.a(s_13), .O(gate55inter4));
  nand2 gate292(.a(gate55inter4), .b(gate55inter3), .O(gate55inter5));
  nor2  gate293(.a(gate55inter5), .b(gate55inter2), .O(gate55inter6));
  inv1  gate294(.a(N286), .O(gate55inter7));
  inv1  gate295(.a(N287), .O(gate55inter8));
  nand2 gate296(.a(gate55inter8), .b(gate55inter7), .O(gate55inter9));
  nand2 gate297(.a(s_13), .b(gate55inter3), .O(gate55inter10));
  nor2  gate298(.a(gate55inter10), .b(gate55inter9), .O(gate55inter11));
  nor2  gate299(.a(gate55inter11), .b(gate55inter6), .O(gate55inter12));
  nand2 gate300(.a(gate55inter12), .b(gate55inter1), .O(N320));
xor2 gate56( .a(N288), .b(N289), .O(N321) );
xor2 gate57( .a(N290), .b(N293), .O(N338) );
xor2 gate58( .a(N296), .b(N299), .O(N339) );
xor2 gate59( .a(N290), .b(N296), .O(N340) );
xor2 gate60( .a(N293), .b(N299), .O(N341) );

  xor2  gate483(.a(N305), .b(N302), .O(gate61inter0));
  nand2 gate484(.a(gate61inter0), .b(s_40), .O(gate61inter1));
  and2  gate485(.a(N305), .b(N302), .O(gate61inter2));
  inv1  gate486(.a(s_40), .O(gate61inter3));
  inv1  gate487(.a(s_41), .O(gate61inter4));
  nand2 gate488(.a(gate61inter4), .b(gate61inter3), .O(gate61inter5));
  nor2  gate489(.a(gate61inter5), .b(gate61inter2), .O(gate61inter6));
  inv1  gate490(.a(N302), .O(gate61inter7));
  inv1  gate491(.a(N305), .O(gate61inter8));
  nand2 gate492(.a(gate61inter8), .b(gate61inter7), .O(gate61inter9));
  nand2 gate493(.a(s_41), .b(gate61inter3), .O(gate61inter10));
  nor2  gate494(.a(gate61inter10), .b(gate61inter9), .O(gate61inter11));
  nor2  gate495(.a(gate61inter11), .b(gate61inter6), .O(gate61inter12));
  nand2 gate496(.a(gate61inter12), .b(gate61inter1), .O(N342));
xor2 gate62( .a(N308), .b(N311), .O(N343) );

  xor2  gate231(.a(N308), .b(N302), .O(gate63inter0));
  nand2 gate232(.a(gate63inter0), .b(s_4), .O(gate63inter1));
  and2  gate233(.a(N308), .b(N302), .O(gate63inter2));
  inv1  gate234(.a(s_4), .O(gate63inter3));
  inv1  gate235(.a(s_5), .O(gate63inter4));
  nand2 gate236(.a(gate63inter4), .b(gate63inter3), .O(gate63inter5));
  nor2  gate237(.a(gate63inter5), .b(gate63inter2), .O(gate63inter6));
  inv1  gate238(.a(N302), .O(gate63inter7));
  inv1  gate239(.a(N308), .O(gate63inter8));
  nand2 gate240(.a(gate63inter8), .b(gate63inter7), .O(gate63inter9));
  nand2 gate241(.a(s_5), .b(gate63inter3), .O(gate63inter10));
  nor2  gate242(.a(gate63inter10), .b(gate63inter9), .O(gate63inter11));
  nor2  gate243(.a(gate63inter11), .b(gate63inter6), .O(gate63inter12));
  nand2 gate244(.a(gate63inter12), .b(gate63inter1), .O(N344));
xor2 gate64( .a(N305), .b(N311), .O(N345) );
xor2 gate65( .a(N266), .b(N342), .O(N346) );
xor2 gate66( .a(N267), .b(N343), .O(N347) );
xor2 gate67( .a(N268), .b(N344), .O(N348) );
xor2 gate68( .a(N269), .b(N345), .O(N349) );
xor2 gate69( .a(N270), .b(N338), .O(N350) );
xor2 gate70( .a(N271), .b(N339), .O(N351) );

  xor2  gate455(.a(N340), .b(N272), .O(gate71inter0));
  nand2 gate456(.a(gate71inter0), .b(s_36), .O(gate71inter1));
  and2  gate457(.a(N340), .b(N272), .O(gate71inter2));
  inv1  gate458(.a(s_36), .O(gate71inter3));
  inv1  gate459(.a(s_37), .O(gate71inter4));
  nand2 gate460(.a(gate71inter4), .b(gate71inter3), .O(gate71inter5));
  nor2  gate461(.a(gate71inter5), .b(gate71inter2), .O(gate71inter6));
  inv1  gate462(.a(N272), .O(gate71inter7));
  inv1  gate463(.a(N340), .O(gate71inter8));
  nand2 gate464(.a(gate71inter8), .b(gate71inter7), .O(gate71inter9));
  nand2 gate465(.a(s_37), .b(gate71inter3), .O(gate71inter10));
  nor2  gate466(.a(gate71inter10), .b(gate71inter9), .O(gate71inter11));
  nor2  gate467(.a(gate71inter11), .b(gate71inter6), .O(gate71inter12));
  nand2 gate468(.a(gate71inter12), .b(gate71inter1), .O(N352));
xor2 gate72( .a(N273), .b(N341), .O(N353) );
xor2 gate73( .a(N314), .b(N346), .O(N354) );
xor2 gate74( .a(N315), .b(N347), .O(N367) );
xor2 gate75( .a(N316), .b(N348), .O(N380) );
xor2 gate76( .a(N317), .b(N349), .O(N393) );
xor2 gate77( .a(N318), .b(N350), .O(N406) );
xor2 gate78( .a(N319), .b(N351), .O(N419) );

  xor2  gate217(.a(N352), .b(N320), .O(gate79inter0));
  nand2 gate218(.a(gate79inter0), .b(s_2), .O(gate79inter1));
  and2  gate219(.a(N352), .b(N320), .O(gate79inter2));
  inv1  gate220(.a(s_2), .O(gate79inter3));
  inv1  gate221(.a(s_3), .O(gate79inter4));
  nand2 gate222(.a(gate79inter4), .b(gate79inter3), .O(gate79inter5));
  nor2  gate223(.a(gate79inter5), .b(gate79inter2), .O(gate79inter6));
  inv1  gate224(.a(N320), .O(gate79inter7));
  inv1  gate225(.a(N352), .O(gate79inter8));
  nand2 gate226(.a(gate79inter8), .b(gate79inter7), .O(gate79inter9));
  nand2 gate227(.a(s_3), .b(gate79inter3), .O(gate79inter10));
  nor2  gate228(.a(gate79inter10), .b(gate79inter9), .O(gate79inter11));
  nor2  gate229(.a(gate79inter11), .b(gate79inter6), .O(gate79inter12));
  nand2 gate230(.a(gate79inter12), .b(gate79inter1), .O(N432));
xor2 gate80( .a(N321), .b(N353), .O(N445) );
inv1 gate81( .a(N354), .O(N554) );
inv1 gate82( .a(N367), .O(N555) );
inv1 gate83( .a(N380), .O(N556) );
inv1 gate84( .a(N354), .O(N557) );
inv1 gate85( .a(N367), .O(N558) );
inv1 gate86( .a(N393), .O(N559) );
inv1 gate87( .a(N354), .O(N560) );
inv1 gate88( .a(N380), .O(N561) );
inv1 gate89( .a(N393), .O(N562) );
inv1 gate90( .a(N367), .O(N563) );
inv1 gate91( .a(N380), .O(N564) );
inv1 gate92( .a(N393), .O(N565) );
inv1 gate93( .a(N419), .O(N566) );
inv1 gate94( .a(N445), .O(N567) );
inv1 gate95( .a(N419), .O(N568) );
inv1 gate96( .a(N432), .O(N569) );
inv1 gate97( .a(N406), .O(N570) );
inv1 gate98( .a(N445), .O(N571) );
inv1 gate99( .a(N406), .O(N572) );
inv1 gate100( .a(N432), .O(N573) );
inv1 gate101( .a(N406), .O(N574) );
inv1 gate102( .a(N419), .O(N575) );
inv1 gate103( .a(N432), .O(N576) );
inv1 gate104( .a(N406), .O(N577) );
inv1 gate105( .a(N419), .O(N578) );
inv1 gate106( .a(N445), .O(N579) );
inv1 gate107( .a(N406), .O(N580) );
inv1 gate108( .a(N432), .O(N581) );
inv1 gate109( .a(N445), .O(N582) );
inv1 gate110( .a(N419), .O(N583) );
inv1 gate111( .a(N432), .O(N584) );
inv1 gate112( .a(N445), .O(N585) );
inv1 gate113( .a(N367), .O(N586) );
inv1 gate114( .a(N393), .O(N587) );
inv1 gate115( .a(N367), .O(N588) );
inv1 gate116( .a(N380), .O(N589) );
inv1 gate117( .a(N354), .O(N590) );
inv1 gate118( .a(N393), .O(N591) );
inv1 gate119( .a(N354), .O(N592) );
inv1 gate120( .a(N380), .O(N593) );
and4 gate121( .a(N554), .b(N555), .c(N556), .d(N393), .O(N594) );
and4 gate122( .a(N557), .b(N558), .c(N380), .d(N559), .O(N595) );
and4 gate123( .a(N560), .b(N367), .c(N561), .d(N562), .O(N596) );
and4 gate124( .a(N354), .b(N563), .c(N564), .d(N565), .O(N597) );
and4 gate125( .a(N574), .b(N575), .c(N576), .d(N445), .O(N598) );
and4 gate126( .a(N577), .b(N578), .c(N432), .d(N579), .O(N599) );
and4 gate127( .a(N580), .b(N419), .c(N581), .d(N582), .O(N600) );
and4 gate128( .a(N406), .b(N583), .c(N584), .d(N585), .O(N601) );
or4 gate129( .a(N594), .b(N595), .c(N596), .d(N597), .O(N602) );
or4 gate130( .a(N598), .b(N599), .c(N600), .d(N601), .O(N607) );
and5 gate131( .a(N406), .b(N566), .c(N432), .d(N567), .e(N602), .O(N620) );
and5 gate132( .a(N406), .b(N568), .c(N569), .d(N445), .e(N602), .O(N625) );
and5 gate133( .a(N570), .b(N419), .c(N432), .d(N571), .e(N602), .O(N630) );
and5 gate134( .a(N572), .b(N419), .c(N573), .d(N445), .e(N602), .O(N635) );
and5 gate135( .a(N354), .b(N586), .c(N380), .d(N587), .e(N607), .O(N640) );
and5 gate136( .a(N354), .b(N588), .c(N589), .d(N393), .e(N607), .O(N645) );
and5 gate137( .a(N590), .b(N367), .c(N380), .d(N591), .e(N607), .O(N650) );
and5 gate138( .a(N592), .b(N367), .c(N593), .d(N393), .e(N607), .O(N655) );
and2 gate139( .a(N354), .b(N620), .O(N692) );
and2 gate140( .a(N367), .b(N620), .O(N693) );
and2 gate141( .a(N380), .b(N620), .O(N694) );
and2 gate142( .a(N393), .b(N620), .O(N695) );
and2 gate143( .a(N354), .b(N625), .O(N696) );
and2 gate144( .a(N367), .b(N625), .O(N697) );
and2 gate145( .a(N380), .b(N625), .O(N698) );
and2 gate146( .a(N393), .b(N625), .O(N699) );
and2 gate147( .a(N354), .b(N630), .O(N700) );
and2 gate148( .a(N367), .b(N630), .O(N701) );
and2 gate149( .a(N380), .b(N630), .O(N702) );
and2 gate150( .a(N393), .b(N630), .O(N703) );
and2 gate151( .a(N354), .b(N635), .O(N704) );
and2 gate152( .a(N367), .b(N635), .O(N705) );
and2 gate153( .a(N380), .b(N635), .O(N706) );
and2 gate154( .a(N393), .b(N635), .O(N707) );
and2 gate155( .a(N406), .b(N640), .O(N708) );
and2 gate156( .a(N419), .b(N640), .O(N709) );
and2 gate157( .a(N432), .b(N640), .O(N710) );
and2 gate158( .a(N445), .b(N640), .O(N711) );
and2 gate159( .a(N406), .b(N645), .O(N712) );
and2 gate160( .a(N419), .b(N645), .O(N713) );
and2 gate161( .a(N432), .b(N645), .O(N714) );
and2 gate162( .a(N445), .b(N645), .O(N715) );
and2 gate163( .a(N406), .b(N650), .O(N716) );
and2 gate164( .a(N419), .b(N650), .O(N717) );
and2 gate165( .a(N432), .b(N650), .O(N718) );
and2 gate166( .a(N445), .b(N650), .O(N719) );
and2 gate167( .a(N406), .b(N655), .O(N720) );
and2 gate168( .a(N419), .b(N655), .O(N721) );
and2 gate169( .a(N432), .b(N655), .O(N722) );
and2 gate170( .a(N445), .b(N655), .O(N723) );
xor2 gate171( .a(N1), .b(N692), .O(N724) );
xor2 gate172( .a(N5), .b(N693), .O(N725) );

  xor2  gate399(.a(N694), .b(N9), .O(gate173inter0));
  nand2 gate400(.a(gate173inter0), .b(s_28), .O(gate173inter1));
  and2  gate401(.a(N694), .b(N9), .O(gate173inter2));
  inv1  gate402(.a(s_28), .O(gate173inter3));
  inv1  gate403(.a(s_29), .O(gate173inter4));
  nand2 gate404(.a(gate173inter4), .b(gate173inter3), .O(gate173inter5));
  nor2  gate405(.a(gate173inter5), .b(gate173inter2), .O(gate173inter6));
  inv1  gate406(.a(N9), .O(gate173inter7));
  inv1  gate407(.a(N694), .O(gate173inter8));
  nand2 gate408(.a(gate173inter8), .b(gate173inter7), .O(gate173inter9));
  nand2 gate409(.a(s_29), .b(gate173inter3), .O(gate173inter10));
  nor2  gate410(.a(gate173inter10), .b(gate173inter9), .O(gate173inter11));
  nor2  gate411(.a(gate173inter11), .b(gate173inter6), .O(gate173inter12));
  nand2 gate412(.a(gate173inter12), .b(gate173inter1), .O(N726));
xor2 gate174( .a(N13), .b(N695), .O(N727) );
xor2 gate175( .a(N17), .b(N696), .O(N728) );

  xor2  gate245(.a(N697), .b(N21), .O(gate176inter0));
  nand2 gate246(.a(gate176inter0), .b(s_6), .O(gate176inter1));
  and2  gate247(.a(N697), .b(N21), .O(gate176inter2));
  inv1  gate248(.a(s_6), .O(gate176inter3));
  inv1  gate249(.a(s_7), .O(gate176inter4));
  nand2 gate250(.a(gate176inter4), .b(gate176inter3), .O(gate176inter5));
  nor2  gate251(.a(gate176inter5), .b(gate176inter2), .O(gate176inter6));
  inv1  gate252(.a(N21), .O(gate176inter7));
  inv1  gate253(.a(N697), .O(gate176inter8));
  nand2 gate254(.a(gate176inter8), .b(gate176inter7), .O(gate176inter9));
  nand2 gate255(.a(s_7), .b(gate176inter3), .O(gate176inter10));
  nor2  gate256(.a(gate176inter10), .b(gate176inter9), .O(gate176inter11));
  nor2  gate257(.a(gate176inter11), .b(gate176inter6), .O(gate176inter12));
  nand2 gate258(.a(gate176inter12), .b(gate176inter1), .O(N729));
xor2 gate177( .a(N25), .b(N698), .O(N730) );

  xor2  gate469(.a(N699), .b(N29), .O(gate178inter0));
  nand2 gate470(.a(gate178inter0), .b(s_38), .O(gate178inter1));
  and2  gate471(.a(N699), .b(N29), .O(gate178inter2));
  inv1  gate472(.a(s_38), .O(gate178inter3));
  inv1  gate473(.a(s_39), .O(gate178inter4));
  nand2 gate474(.a(gate178inter4), .b(gate178inter3), .O(gate178inter5));
  nor2  gate475(.a(gate178inter5), .b(gate178inter2), .O(gate178inter6));
  inv1  gate476(.a(N29), .O(gate178inter7));
  inv1  gate477(.a(N699), .O(gate178inter8));
  nand2 gate478(.a(gate178inter8), .b(gate178inter7), .O(gate178inter9));
  nand2 gate479(.a(s_39), .b(gate178inter3), .O(gate178inter10));
  nor2  gate480(.a(gate178inter10), .b(gate178inter9), .O(gate178inter11));
  nor2  gate481(.a(gate178inter11), .b(gate178inter6), .O(gate178inter12));
  nand2 gate482(.a(gate178inter12), .b(gate178inter1), .O(N731));
xor2 gate179( .a(N33), .b(N700), .O(N732) );
xor2 gate180( .a(N37), .b(N701), .O(N733) );

  xor2  gate259(.a(N702), .b(N41), .O(gate181inter0));
  nand2 gate260(.a(gate181inter0), .b(s_8), .O(gate181inter1));
  and2  gate261(.a(N702), .b(N41), .O(gate181inter2));
  inv1  gate262(.a(s_8), .O(gate181inter3));
  inv1  gate263(.a(s_9), .O(gate181inter4));
  nand2 gate264(.a(gate181inter4), .b(gate181inter3), .O(gate181inter5));
  nor2  gate265(.a(gate181inter5), .b(gate181inter2), .O(gate181inter6));
  inv1  gate266(.a(N41), .O(gate181inter7));
  inv1  gate267(.a(N702), .O(gate181inter8));
  nand2 gate268(.a(gate181inter8), .b(gate181inter7), .O(gate181inter9));
  nand2 gate269(.a(s_9), .b(gate181inter3), .O(gate181inter10));
  nor2  gate270(.a(gate181inter10), .b(gate181inter9), .O(gate181inter11));
  nor2  gate271(.a(gate181inter11), .b(gate181inter6), .O(gate181inter12));
  nand2 gate272(.a(gate181inter12), .b(gate181inter1), .O(N734));
xor2 gate182( .a(N45), .b(N703), .O(N735) );
xor2 gate183( .a(N49), .b(N704), .O(N736) );
xor2 gate184( .a(N53), .b(N705), .O(N737) );
xor2 gate185( .a(N57), .b(N706), .O(N738) );

  xor2  gate343(.a(N707), .b(N61), .O(gate186inter0));
  nand2 gate344(.a(gate186inter0), .b(s_20), .O(gate186inter1));
  and2  gate345(.a(N707), .b(N61), .O(gate186inter2));
  inv1  gate346(.a(s_20), .O(gate186inter3));
  inv1  gate347(.a(s_21), .O(gate186inter4));
  nand2 gate348(.a(gate186inter4), .b(gate186inter3), .O(gate186inter5));
  nor2  gate349(.a(gate186inter5), .b(gate186inter2), .O(gate186inter6));
  inv1  gate350(.a(N61), .O(gate186inter7));
  inv1  gate351(.a(N707), .O(gate186inter8));
  nand2 gate352(.a(gate186inter8), .b(gate186inter7), .O(gate186inter9));
  nand2 gate353(.a(s_21), .b(gate186inter3), .O(gate186inter10));
  nor2  gate354(.a(gate186inter10), .b(gate186inter9), .O(gate186inter11));
  nor2  gate355(.a(gate186inter11), .b(gate186inter6), .O(gate186inter12));
  nand2 gate356(.a(gate186inter12), .b(gate186inter1), .O(N739));

  xor2  gate427(.a(N708), .b(N65), .O(gate187inter0));
  nand2 gate428(.a(gate187inter0), .b(s_32), .O(gate187inter1));
  and2  gate429(.a(N708), .b(N65), .O(gate187inter2));
  inv1  gate430(.a(s_32), .O(gate187inter3));
  inv1  gate431(.a(s_33), .O(gate187inter4));
  nand2 gate432(.a(gate187inter4), .b(gate187inter3), .O(gate187inter5));
  nor2  gate433(.a(gate187inter5), .b(gate187inter2), .O(gate187inter6));
  inv1  gate434(.a(N65), .O(gate187inter7));
  inv1  gate435(.a(N708), .O(gate187inter8));
  nand2 gate436(.a(gate187inter8), .b(gate187inter7), .O(gate187inter9));
  nand2 gate437(.a(s_33), .b(gate187inter3), .O(gate187inter10));
  nor2  gate438(.a(gate187inter10), .b(gate187inter9), .O(gate187inter11));
  nor2  gate439(.a(gate187inter11), .b(gate187inter6), .O(gate187inter12));
  nand2 gate440(.a(gate187inter12), .b(gate187inter1), .O(N740));

  xor2  gate273(.a(N709), .b(N69), .O(gate188inter0));
  nand2 gate274(.a(gate188inter0), .b(s_10), .O(gate188inter1));
  and2  gate275(.a(N709), .b(N69), .O(gate188inter2));
  inv1  gate276(.a(s_10), .O(gate188inter3));
  inv1  gate277(.a(s_11), .O(gate188inter4));
  nand2 gate278(.a(gate188inter4), .b(gate188inter3), .O(gate188inter5));
  nor2  gate279(.a(gate188inter5), .b(gate188inter2), .O(gate188inter6));
  inv1  gate280(.a(N69), .O(gate188inter7));
  inv1  gate281(.a(N709), .O(gate188inter8));
  nand2 gate282(.a(gate188inter8), .b(gate188inter7), .O(gate188inter9));
  nand2 gate283(.a(s_11), .b(gate188inter3), .O(gate188inter10));
  nor2  gate284(.a(gate188inter10), .b(gate188inter9), .O(gate188inter11));
  nor2  gate285(.a(gate188inter11), .b(gate188inter6), .O(gate188inter12));
  nand2 gate286(.a(gate188inter12), .b(gate188inter1), .O(N741));
xor2 gate189( .a(N73), .b(N710), .O(N742) );
xor2 gate190( .a(N77), .b(N711), .O(N743) );
xor2 gate191( .a(N81), .b(N712), .O(N744) );
xor2 gate192( .a(N85), .b(N713), .O(N745) );
xor2 gate193( .a(N89), .b(N714), .O(N746) );
xor2 gate194( .a(N93), .b(N715), .O(N747) );
xor2 gate195( .a(N97), .b(N716), .O(N748) );
xor2 gate196( .a(N101), .b(N717), .O(N749) );

  xor2  gate315(.a(N718), .b(N105), .O(gate197inter0));
  nand2 gate316(.a(gate197inter0), .b(s_16), .O(gate197inter1));
  and2  gate317(.a(N718), .b(N105), .O(gate197inter2));
  inv1  gate318(.a(s_16), .O(gate197inter3));
  inv1  gate319(.a(s_17), .O(gate197inter4));
  nand2 gate320(.a(gate197inter4), .b(gate197inter3), .O(gate197inter5));
  nor2  gate321(.a(gate197inter5), .b(gate197inter2), .O(gate197inter6));
  inv1  gate322(.a(N105), .O(gate197inter7));
  inv1  gate323(.a(N718), .O(gate197inter8));
  nand2 gate324(.a(gate197inter8), .b(gate197inter7), .O(gate197inter9));
  nand2 gate325(.a(s_17), .b(gate197inter3), .O(gate197inter10));
  nor2  gate326(.a(gate197inter10), .b(gate197inter9), .O(gate197inter11));
  nor2  gate327(.a(gate197inter11), .b(gate197inter6), .O(gate197inter12));
  nand2 gate328(.a(gate197inter12), .b(gate197inter1), .O(N750));
xor2 gate198( .a(N109), .b(N719), .O(N751) );
xor2 gate199( .a(N113), .b(N720), .O(N752) );

  xor2  gate385(.a(N721), .b(N117), .O(gate200inter0));
  nand2 gate386(.a(gate200inter0), .b(s_26), .O(gate200inter1));
  and2  gate387(.a(N721), .b(N117), .O(gate200inter2));
  inv1  gate388(.a(s_26), .O(gate200inter3));
  inv1  gate389(.a(s_27), .O(gate200inter4));
  nand2 gate390(.a(gate200inter4), .b(gate200inter3), .O(gate200inter5));
  nor2  gate391(.a(gate200inter5), .b(gate200inter2), .O(gate200inter6));
  inv1  gate392(.a(N117), .O(gate200inter7));
  inv1  gate393(.a(N721), .O(gate200inter8));
  nand2 gate394(.a(gate200inter8), .b(gate200inter7), .O(gate200inter9));
  nand2 gate395(.a(s_27), .b(gate200inter3), .O(gate200inter10));
  nor2  gate396(.a(gate200inter10), .b(gate200inter9), .O(gate200inter11));
  nor2  gate397(.a(gate200inter11), .b(gate200inter6), .O(gate200inter12));
  nand2 gate398(.a(gate200inter12), .b(gate200inter1), .O(N753));
xor2 gate201( .a(N121), .b(N722), .O(N754) );
xor2 gate202( .a(N125), .b(N723), .O(N755) );

endmodule