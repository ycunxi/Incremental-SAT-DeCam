module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);

input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;//RE__PI;

input s_0,s_1;//RE__ALLOW(00,01,10,11);
input s_2,s_3;//RE__ALLOW(00,01,10,11);
input s_4,s_5;//RE__ALLOW(00,01,10,11);
input s_6,s_7;//RE__ALLOW(00,01,10,11);
input s_8,s_9;//RE__ALLOW(00,01,10,11);
input s_10,s_11;//RE__ALLOW(00,01,10,11);
input s_12,s_13;//RE__ALLOW(00,01,10,11);
input s_14,s_15;//RE__ALLOW(00,01,10,11);
input s_16,s_17;//RE__ALLOW(00,01,10,11);
input s_18,s_19;//RE__ALLOW(00,01,10,11);
input s_20,s_21;//RE__ALLOW(00,01,10,11);
input s_22,s_23;//RE__ALLOW(00,01,10,11);
input s_24,s_25;//RE__ALLOW(00,01,10,11);
input s_26,s_27;//RE__ALLOW(00,01,10,11);
input s_28,s_29;//RE__ALLOW(00,01,10,11);
input s_30,s_31;//RE__ALLOW(00,01,10,11);
input s_32,s_33;//RE__ALLOW(00,01,10,11);
input s_34,s_35;//RE__ALLOW(00,01,10,11);
input s_36,s_37;//RE__ALLOW(00,01,10,11);
input s_38,s_39;//RE__ALLOW(00,01,10,11);
input s_40,s_41;//RE__ALLOW(00,01,10,11);
input s_42,s_43;//RE__ALLOW(00,01,10,11);
input s_44,s_45;//RE__ALLOW(00,01,10,11);
input s_46,s_47;//RE__ALLOW(00,01,10,11);
input s_48,s_49;//RE__ALLOW(00,01,10,11);
input s_50,s_51;//RE__ALLOW(00,01,10,11);
input s_52,s_53;//RE__ALLOW(00,01,10,11);
input s_54,s_55;//RE__ALLOW(00,01,10,11);
input s_56,s_57;//RE__ALLOW(00,01,10,11);
input s_58,s_59;//RE__ALLOW(00,01,10,11);
input s_60,s_61;//RE__ALLOW(00,01,10,11);
input s_62,s_63;//RE__ALLOW(00,01,10,11);
input s_64,s_65;//RE__ALLOW(00,01,10,11);
input s_66,s_67;//RE__ALLOW(00,01,10,11);
input s_68,s_69;//RE__ALLOW(00,01,10,11);
input s_70,s_71;//RE__ALLOW(00,01,10,11);
input s_72,s_73;//RE__ALLOW(00,01,10,11);
input s_74,s_75;//RE__ALLOW(00,01,10,11);
input s_76,s_77;//RE__ALLOW(00,01,10,11);
input s_78,s_79;//RE__ALLOW(00,01,10,11);
input s_80,s_81;//RE__ALLOW(00,01,10,11);
input s_82,s_83;//RE__ALLOW(00,01,10,11);
input s_84,s_85;//RE__ALLOW(00,01,10,11);
input s_86,s_87;//RE__ALLOW(00,01,10,11);
input s_88,s_89;//RE__ALLOW(00,01,10,11);
input s_90,s_91;//RE__ALLOW(00,01,10,11);
input s_92,s_93;//RE__ALLOW(00,01,10,11);
input s_94,s_95;//RE__ALLOW(00,01,10,11);
input s_96,s_97;//RE__ALLOW(00,01,10,11);
input s_98,s_99;//RE__ALLOW(00,01,10,11);
input s_100,s_101;//RE__ALLOW(00,01,10,11);
input s_102,s_103;//RE__ALLOW(00,01,10,11);
input s_104,s_105;//RE__ALLOW(00,01,10,11);
input s_106,s_107;//RE__ALLOW(00,01,10,11);
input s_108,s_109;//RE__ALLOW(00,01,10,11);
input s_110,s_111;//RE__ALLOW(00,01,10,11);
input s_112,s_113;//RE__ALLOW(00,01,10,11);
input s_114,s_115;//RE__ALLOW(00,01,10,11);
input s_116,s_117;//RE__ALLOW(00,01,10,11);
input s_118,s_119;//RE__ALLOW(00,01,10,11);
input s_120,s_121;//RE__ALLOW(00,01,10,11);
input s_122,s_123;//RE__ALLOW(00,01,10,11);
input s_124,s_125;//RE__ALLOW(00,01,10,11);
input s_126,s_127;//RE__ALLOW(00,01,10,11);
input s_128,s_129;//RE__ALLOW(00,01,10,11);
input s_130,s_131;//RE__ALLOW(00,01,10,11);
input s_132,s_133;//RE__ALLOW(00,01,10,11);
input s_134,s_135;//RE__ALLOW(00,01,10,11);
input s_136,s_137;//RE__ALLOW(00,01,10,11);
input s_138,s_139;//RE__ALLOW(00,01,10,11);
input s_140,s_141;//RE__ALLOW(00,01,10,11);
input s_142,s_143;//RE__ALLOW(00,01,10,11);
input s_144,s_145;//RE__ALLOW(00,01,10,11);
input s_146,s_147;//RE__ALLOW(00,01,10,11);
input s_148,s_149;//RE__ALLOW(00,01,10,11);
input s_150,s_151;//RE__ALLOW(00,01,10,11);
input s_152,s_153;//RE__ALLOW(00,01,10,11);
input s_154,s_155;//RE__ALLOW(00,01,10,11);
input s_156,s_157;//RE__ALLOW(00,01,10,11);
input s_158,s_159;//RE__ALLOW(00,01,10,11);
input s_160,s_161;//RE__ALLOW(00,01,10,11);
input s_162,s_163;//RE__ALLOW(00,01,10,11);
input s_164,s_165;//RE__ALLOW(00,01,10,11);
input s_166,s_167;//RE__ALLOW(00,01,10,11);
input s_168,s_169;//RE__ALLOW(00,01,10,11);
input s_170,s_171;//RE__ALLOW(00,01,10,11);
input s_172,s_173;//RE__ALLOW(00,01,10,11);
input s_174,s_175;//RE__ALLOW(00,01,10,11);
input s_176,s_177;//RE__ALLOW(00,01,10,11);
input s_178,s_179;//RE__ALLOW(00,01,10,11);
input s_180,s_181;//RE__ALLOW(00,01,10,11);
input s_182,s_183;//RE__ALLOW(00,01,10,11);
input s_184,s_185;//RE__ALLOW(00,01,10,11);
input s_186,s_187;//RE__ALLOW(00,01,10,11);
input s_188,s_189;//RE__ALLOW(00,01,10,11);
input s_190,s_191;//RE__ALLOW(00,01,10,11);
input s_192,s_193;//RE__ALLOW(00,01,10,11);
input s_194,s_195;//RE__ALLOW(00,01,10,11);
input s_196,s_197;//RE__ALLOW(00,01,10,11);
input s_198,s_199;//RE__ALLOW(00,01,10,11);
input s_200,s_201;//RE__ALLOW(00,01,10,11);
input s_202,s_203;//RE__ALLOW(00,01,10,11);
input s_204,s_205;//RE__ALLOW(00,01,10,11);
input s_206,s_207;//RE__ALLOW(00,01,10,11);
input s_208,s_209;//RE__ALLOW(00,01,10,11);
input s_210,s_211;//RE__ALLOW(00,01,10,11);
input s_212,s_213;//RE__ALLOW(00,01,10,11);
input s_214,s_215;//RE__ALLOW(00,01,10,11);
input s_216,s_217;//RE__ALLOW(00,01,10,11);
input s_218,s_219;//RE__ALLOW(00,01,10,11);
input s_220,s_221;//RE__ALLOW(00,01,10,11);
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;

  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate139inter0, gate139inter1, gate139inter2, gate139inter3, gate139inter4, gate139inter5, gate139inter6, gate139inter7, gate139inter8, gate139inter9, gate139inter10, gate139inter11, gate139inter12, gate73inter0, gate73inter1, gate73inter2, gate73inter3, gate73inter4, gate73inter5, gate73inter6, gate73inter7, gate73inter8, gate73inter9, gate73inter10, gate73inter11, gate73inter12, gate277inter0, gate277inter1, gate277inter2, gate277inter3, gate277inter4, gate277inter5, gate277inter6, gate277inter7, gate277inter8, gate277inter9, gate277inter10, gate277inter11, gate277inter12, gate150inter0, gate150inter1, gate150inter2, gate150inter3, gate150inter4, gate150inter5, gate150inter6, gate150inter7, gate150inter8, gate150inter9, gate150inter10, gate150inter11, gate150inter12, gate395inter0, gate395inter1, gate395inter2, gate395inter3, gate395inter4, gate395inter5, gate395inter6, gate395inter7, gate395inter8, gate395inter9, gate395inter10, gate395inter11, gate395inter12, gate224inter0, gate224inter1, gate224inter2, gate224inter3, gate224inter4, gate224inter5, gate224inter6, gate224inter7, gate224inter8, gate224inter9, gate224inter10, gate224inter11, gate224inter12, gate183inter0, gate183inter1, gate183inter2, gate183inter3, gate183inter4, gate183inter5, gate183inter6, gate183inter7, gate183inter8, gate183inter9, gate183inter10, gate183inter11, gate183inter12, gate226inter0, gate226inter1, gate226inter2, gate226inter3, gate226inter4, gate226inter5, gate226inter6, gate226inter7, gate226inter8, gate226inter9, gate226inter10, gate226inter11, gate226inter12, gate441inter0, gate441inter1, gate441inter2, gate441inter3, gate441inter4, gate441inter5, gate441inter6, gate441inter7, gate441inter8, gate441inter9, gate441inter10, gate441inter11, gate441inter12, gate145inter0, gate145inter1, gate145inter2, gate145inter3, gate145inter4, gate145inter5, gate145inter6, gate145inter7, gate145inter8, gate145inter9, gate145inter10, gate145inter11, gate145inter12, gate513inter0, gate513inter1, gate513inter2, gate513inter3, gate513inter4, gate513inter5, gate513inter6, gate513inter7, gate513inter8, gate513inter9, gate513inter10, gate513inter11, gate513inter12, gate56inter0, gate56inter1, gate56inter2, gate56inter3, gate56inter4, gate56inter5, gate56inter6, gate56inter7, gate56inter8, gate56inter9, gate56inter10, gate56inter11, gate56inter12, gate86inter0, gate86inter1, gate86inter2, gate86inter3, gate86inter4, gate86inter5, gate86inter6, gate86inter7, gate86inter8, gate86inter9, gate86inter10, gate86inter11, gate86inter12, gate41inter0, gate41inter1, gate41inter2, gate41inter3, gate41inter4, gate41inter5, gate41inter6, gate41inter7, gate41inter8, gate41inter9, gate41inter10, gate41inter11, gate41inter12, gate170inter0, gate170inter1, gate170inter2, gate170inter3, gate170inter4, gate170inter5, gate170inter6, gate170inter7, gate170inter8, gate170inter9, gate170inter10, gate170inter11, gate170inter12, gate109inter0, gate109inter1, gate109inter2, gate109inter3, gate109inter4, gate109inter5, gate109inter6, gate109inter7, gate109inter8, gate109inter9, gate109inter10, gate109inter11, gate109inter12, gate35inter0, gate35inter1, gate35inter2, gate35inter3, gate35inter4, gate35inter5, gate35inter6, gate35inter7, gate35inter8, gate35inter9, gate35inter10, gate35inter11, gate35inter12, gate32inter0, gate32inter1, gate32inter2, gate32inter3, gate32inter4, gate32inter5, gate32inter6, gate32inter7, gate32inter8, gate32inter9, gate32inter10, gate32inter11, gate32inter12, gate186inter0, gate186inter1, gate186inter2, gate186inter3, gate186inter4, gate186inter5, gate186inter6, gate186inter7, gate186inter8, gate186inter9, gate186inter10, gate186inter11, gate186inter12, gate71inter0, gate71inter1, gate71inter2, gate71inter3, gate71inter4, gate71inter5, gate71inter6, gate71inter7, gate71inter8, gate71inter9, gate71inter10, gate71inter11, gate71inter12, gate174inter0, gate174inter1, gate174inter2, gate174inter3, gate174inter4, gate174inter5, gate174inter6, gate174inter7, gate174inter8, gate174inter9, gate174inter10, gate174inter11, gate174inter12, gate405inter0, gate405inter1, gate405inter2, gate405inter3, gate405inter4, gate405inter5, gate405inter6, gate405inter7, gate405inter8, gate405inter9, gate405inter10, gate405inter11, gate405inter12, gate449inter0, gate449inter1, gate449inter2, gate449inter3, gate449inter4, gate449inter5, gate449inter6, gate449inter7, gate449inter8, gate449inter9, gate449inter10, gate449inter11, gate449inter12, gate387inter0, gate387inter1, gate387inter2, gate387inter3, gate387inter4, gate387inter5, gate387inter6, gate387inter7, gate387inter8, gate387inter9, gate387inter10, gate387inter11, gate387inter12, gate24inter0, gate24inter1, gate24inter2, gate24inter3, gate24inter4, gate24inter5, gate24inter6, gate24inter7, gate24inter8, gate24inter9, gate24inter10, gate24inter11, gate24inter12, gate77inter0, gate77inter1, gate77inter2, gate77inter3, gate77inter4, gate77inter5, gate77inter6, gate77inter7, gate77inter8, gate77inter9, gate77inter10, gate77inter11, gate77inter12, gate409inter0, gate409inter1, gate409inter2, gate409inter3, gate409inter4, gate409inter5, gate409inter6, gate409inter7, gate409inter8, gate409inter9, gate409inter10, gate409inter11, gate409inter12, gate215inter0, gate215inter1, gate215inter2, gate215inter3, gate215inter4, gate215inter5, gate215inter6, gate215inter7, gate215inter8, gate215inter9, gate215inter10, gate215inter11, gate215inter12, gate65inter0, gate65inter1, gate65inter2, gate65inter3, gate65inter4, gate65inter5, gate65inter6, gate65inter7, gate65inter8, gate65inter9, gate65inter10, gate65inter11, gate65inter12, gate245inter0, gate245inter1, gate245inter2, gate245inter3, gate245inter4, gate245inter5, gate245inter6, gate245inter7, gate245inter8, gate245inter9, gate245inter10, gate245inter11, gate245inter12, gate37inter0, gate37inter1, gate37inter2, gate37inter3, gate37inter4, gate37inter5, gate37inter6, gate37inter7, gate37inter8, gate37inter9, gate37inter10, gate37inter11, gate37inter12, gate178inter0, gate178inter1, gate178inter2, gate178inter3, gate178inter4, gate178inter5, gate178inter6, gate178inter7, gate178inter8, gate178inter9, gate178inter10, gate178inter11, gate178inter12, gate120inter0, gate120inter1, gate120inter2, gate120inter3, gate120inter4, gate120inter5, gate120inter6, gate120inter7, gate120inter8, gate120inter9, gate120inter10, gate120inter11, gate120inter12, gate481inter0, gate481inter1, gate481inter2, gate481inter3, gate481inter4, gate481inter5, gate481inter6, gate481inter7, gate481inter8, gate481inter9, gate481inter10, gate481inter11, gate481inter12, gate388inter0, gate388inter1, gate388inter2, gate388inter3, gate388inter4, gate388inter5, gate388inter6, gate388inter7, gate388inter8, gate388inter9, gate388inter10, gate388inter11, gate388inter12, gate111inter0, gate111inter1, gate111inter2, gate111inter3, gate111inter4, gate111inter5, gate111inter6, gate111inter7, gate111inter8, gate111inter9, gate111inter10, gate111inter11, gate111inter12, gate185inter0, gate185inter1, gate185inter2, gate185inter3, gate185inter4, gate185inter5, gate185inter6, gate185inter7, gate185inter8, gate185inter9, gate185inter10, gate185inter11, gate185inter12, gate275inter0, gate275inter1, gate275inter2, gate275inter3, gate275inter4, gate275inter5, gate275inter6, gate275inter7, gate275inter8, gate275inter9, gate275inter10, gate275inter11, gate275inter12, gate119inter0, gate119inter1, gate119inter2, gate119inter3, gate119inter4, gate119inter5, gate119inter6, gate119inter7, gate119inter8, gate119inter9, gate119inter10, gate119inter11, gate119inter12, gate129inter0, gate129inter1, gate129inter2, gate129inter3, gate129inter4, gate129inter5, gate129inter6, gate129inter7, gate129inter8, gate129inter9, gate129inter10, gate129inter11, gate129inter12, gate294inter0, gate294inter1, gate294inter2, gate294inter3, gate294inter4, gate294inter5, gate294inter6, gate294inter7, gate294inter8, gate294inter9, gate294inter10, gate294inter11, gate294inter12, gate406inter0, gate406inter1, gate406inter2, gate406inter3, gate406inter4, gate406inter5, gate406inter6, gate406inter7, gate406inter8, gate406inter9, gate406inter10, gate406inter11, gate406inter12, gate397inter0, gate397inter1, gate397inter2, gate397inter3, gate397inter4, gate397inter5, gate397inter6, gate397inter7, gate397inter8, gate397inter9, gate397inter10, gate397inter11, gate397inter12, gate124inter0, gate124inter1, gate124inter2, gate124inter3, gate124inter4, gate124inter5, gate124inter6, gate124inter7, gate124inter8, gate124inter9, gate124inter10, gate124inter11, gate124inter12, gate203inter0, gate203inter1, gate203inter2, gate203inter3, gate203inter4, gate203inter5, gate203inter6, gate203inter7, gate203inter8, gate203inter9, gate203inter10, gate203inter11, gate203inter12, gate118inter0, gate118inter1, gate118inter2, gate118inter3, gate118inter4, gate118inter5, gate118inter6, gate118inter7, gate118inter8, gate118inter9, gate118inter10, gate118inter11, gate118inter12, gate490inter0, gate490inter1, gate490inter2, gate490inter3, gate490inter4, gate490inter5, gate490inter6, gate490inter7, gate490inter8, gate490inter9, gate490inter10, gate490inter11, gate490inter12, gate84inter0, gate84inter1, gate84inter2, gate84inter3, gate84inter4, gate84inter5, gate84inter6, gate84inter7, gate84inter8, gate84inter9, gate84inter10, gate84inter11, gate84inter12, gate122inter0, gate122inter1, gate122inter2, gate122inter3, gate122inter4, gate122inter5, gate122inter6, gate122inter7, gate122inter8, gate122inter9, gate122inter10, gate122inter11, gate122inter12, gate133inter0, gate133inter1, gate133inter2, gate133inter3, gate133inter4, gate133inter5, gate133inter6, gate133inter7, gate133inter8, gate133inter9, gate133inter10, gate133inter11, gate133inter12, gate54inter0, gate54inter1, gate54inter2, gate54inter3, gate54inter4, gate54inter5, gate54inter6, gate54inter7, gate54inter8, gate54inter9, gate54inter10, gate54inter11, gate54inter12, gate293inter0, gate293inter1, gate293inter2, gate293inter3, gate293inter4, gate293inter5, gate293inter6, gate293inter7, gate293inter8, gate293inter9, gate293inter10, gate293inter11, gate293inter12, gate507inter0, gate507inter1, gate507inter2, gate507inter3, gate507inter4, gate507inter5, gate507inter6, gate507inter7, gate507inter8, gate507inter9, gate507inter10, gate507inter11, gate507inter12, gate442inter0, gate442inter1, gate442inter2, gate442inter3, gate442inter4, gate442inter5, gate442inter6, gate442inter7, gate442inter8, gate442inter9, gate442inter10, gate442inter11, gate442inter12, gate143inter0, gate143inter1, gate143inter2, gate143inter3, gate143inter4, gate143inter5, gate143inter6, gate143inter7, gate143inter8, gate143inter9, gate143inter10, gate143inter11, gate143inter12, gate91inter0, gate91inter1, gate91inter2, gate91inter3, gate91inter4, gate91inter5, gate91inter6, gate91inter7, gate91inter8, gate91inter9, gate91inter10, gate91inter11, gate91inter12, gate415inter0, gate415inter1, gate415inter2, gate415inter3, gate415inter4, gate415inter5, gate415inter6, gate415inter7, gate415inter8, gate415inter9, gate415inter10, gate415inter11, gate415inter12, gate439inter0, gate439inter1, gate439inter2, gate439inter3, gate439inter4, gate439inter5, gate439inter6, gate439inter7, gate439inter8, gate439inter9, gate439inter10, gate439inter11, gate439inter12, gate140inter0, gate140inter1, gate140inter2, gate140inter3, gate140inter4, gate140inter5, gate140inter6, gate140inter7, gate140inter8, gate140inter9, gate140inter10, gate140inter11, gate140inter12, gate14inter0, gate14inter1, gate14inter2, gate14inter3, gate14inter4, gate14inter5, gate14inter6, gate14inter7, gate14inter8, gate14inter9, gate14inter10, gate14inter11, gate14inter12, gate22inter0, gate22inter1, gate22inter2, gate22inter3, gate22inter4, gate22inter5, gate22inter6, gate22inter7, gate22inter8, gate22inter9, gate22inter10, gate22inter11, gate22inter12, gate424inter0, gate424inter1, gate424inter2, gate424inter3, gate424inter4, gate424inter5, gate424inter6, gate424inter7, gate424inter8, gate424inter9, gate424inter10, gate424inter11, gate424inter12, gate31inter0, gate31inter1, gate31inter2, gate31inter3, gate31inter4, gate31inter5, gate31inter6, gate31inter7, gate31inter8, gate31inter9, gate31inter10, gate31inter11, gate31inter12, gate440inter0, gate440inter1, gate440inter2, gate440inter3, gate440inter4, gate440inter5, gate440inter6, gate440inter7, gate440inter8, gate440inter9, gate440inter10, gate440inter11, gate440inter12, gate190inter0, gate190inter1, gate190inter2, gate190inter3, gate190inter4, gate190inter5, gate190inter6, gate190inter7, gate190inter8, gate190inter9, gate190inter10, gate190inter11, gate190inter12, gate100inter0, gate100inter1, gate100inter2, gate100inter3, gate100inter4, gate100inter5, gate100inter6, gate100inter7, gate100inter8, gate100inter9, gate100inter10, gate100inter11, gate100inter12, gate34inter0, gate34inter1, gate34inter2, gate34inter3, gate34inter4, gate34inter5, gate34inter6, gate34inter7, gate34inter8, gate34inter9, gate34inter10, gate34inter11, gate34inter12, gate278inter0, gate278inter1, gate278inter2, gate278inter3, gate278inter4, gate278inter5, gate278inter6, gate278inter7, gate278inter8, gate278inter9, gate278inter10, gate278inter11, gate278inter12, gate252inter0, gate252inter1, gate252inter2, gate252inter3, gate252inter4, gate252inter5, gate252inter6, gate252inter7, gate252inter8, gate252inter9, gate252inter10, gate252inter11, gate252inter12, gate504inter0, gate504inter1, gate504inter2, gate504inter3, gate504inter4, gate504inter5, gate504inter6, gate504inter7, gate504inter8, gate504inter9, gate504inter10, gate504inter11, gate504inter12, gate102inter0, gate102inter1, gate102inter2, gate102inter3, gate102inter4, gate102inter5, gate102inter6, gate102inter7, gate102inter8, gate102inter9, gate102inter10, gate102inter11, gate102inter12, gate287inter0, gate287inter1, gate287inter2, gate287inter3, gate287inter4, gate287inter5, gate287inter6, gate287inter7, gate287inter8, gate287inter9, gate287inter10, gate287inter11, gate287inter12, gate51inter0, gate51inter1, gate51inter2, gate51inter3, gate51inter4, gate51inter5, gate51inter6, gate51inter7, gate51inter8, gate51inter9, gate51inter10, gate51inter11, gate51inter12, gate85inter0, gate85inter1, gate85inter2, gate85inter3, gate85inter4, gate85inter5, gate85inter6, gate85inter7, gate85inter8, gate85inter9, gate85inter10, gate85inter11, gate85inter12, gate79inter0, gate79inter1, gate79inter2, gate79inter3, gate79inter4, gate79inter5, gate79inter6, gate79inter7, gate79inter8, gate79inter9, gate79inter10, gate79inter11, gate79inter12, gate33inter0, gate33inter1, gate33inter2, gate33inter3, gate33inter4, gate33inter5, gate33inter6, gate33inter7, gate33inter8, gate33inter9, gate33inter10, gate33inter11, gate33inter12, gate445inter0, gate445inter1, gate445inter2, gate445inter3, gate445inter4, gate445inter5, gate445inter6, gate445inter7, gate445inter8, gate445inter9, gate445inter10, gate445inter11, gate445inter12, gate125inter0, gate125inter1, gate125inter2, gate125inter3, gate125inter4, gate125inter5, gate125inter6, gate125inter7, gate125inter8, gate125inter9, gate125inter10, gate125inter11, gate125inter12, gate70inter0, gate70inter1, gate70inter2, gate70inter3, gate70inter4, gate70inter5, gate70inter6, gate70inter7, gate70inter8, gate70inter9, gate70inter10, gate70inter11, gate70inter12, gate172inter0, gate172inter1, gate172inter2, gate172inter3, gate172inter4, gate172inter5, gate172inter6, gate172inter7, gate172inter8, gate172inter9, gate172inter10, gate172inter11, gate172inter12, gate461inter0, gate461inter1, gate461inter2, gate461inter3, gate461inter4, gate461inter5, gate461inter6, gate461inter7, gate461inter8, gate461inter9, gate461inter10, gate461inter11, gate461inter12, gate402inter0, gate402inter1, gate402inter2, gate402inter3, gate402inter4, gate402inter5, gate402inter6, gate402inter7, gate402inter8, gate402inter9, gate402inter10, gate402inter11, gate402inter12, gate63inter0, gate63inter1, gate63inter2, gate63inter3, gate63inter4, gate63inter5, gate63inter6, gate63inter7, gate63inter8, gate63inter9, gate63inter10, gate63inter11, gate63inter12, gate220inter0, gate220inter1, gate220inter2, gate220inter3, gate220inter4, gate220inter5, gate220inter6, gate220inter7, gate220inter8, gate220inter9, gate220inter10, gate220inter11, gate220inter12, gate117inter0, gate117inter1, gate117inter2, gate117inter3, gate117inter4, gate117inter5, gate117inter6, gate117inter7, gate117inter8, gate117inter9, gate117inter10, gate117inter11, gate117inter12, gate72inter0, gate72inter1, gate72inter2, gate72inter3, gate72inter4, gate72inter5, gate72inter6, gate72inter7, gate72inter8, gate72inter9, gate72inter10, gate72inter11, gate72inter12, gate108inter0, gate108inter1, gate108inter2, gate108inter3, gate108inter4, gate108inter5, gate108inter6, gate108inter7, gate108inter8, gate108inter9, gate108inter10, gate108inter11, gate108inter12, gate420inter0, gate420inter1, gate420inter2, gate420inter3, gate420inter4, gate420inter5, gate420inter6, gate420inter7, gate420inter8, gate420inter9, gate420inter10, gate420inter11, gate420inter12, gate193inter0, gate193inter1, gate193inter2, gate193inter3, gate193inter4, gate193inter5, gate193inter6, gate193inter7, gate193inter8, gate193inter9, gate193inter10, gate193inter11, gate193inter12, gate236inter0, gate236inter1, gate236inter2, gate236inter3, gate236inter4, gate236inter5, gate236inter6, gate236inter7, gate236inter8, gate236inter9, gate236inter10, gate236inter11, gate236inter12, gate25inter0, gate25inter1, gate25inter2, gate25inter3, gate25inter4, gate25inter5, gate25inter6, gate25inter7, gate25inter8, gate25inter9, gate25inter10, gate25inter11, gate25inter12, gate17inter0, gate17inter1, gate17inter2, gate17inter3, gate17inter4, gate17inter5, gate17inter6, gate17inter7, gate17inter8, gate17inter9, gate17inter10, gate17inter11, gate17inter12, gate116inter0, gate116inter1, gate116inter2, gate116inter3, gate116inter4, gate116inter5, gate116inter6, gate116inter7, gate116inter8, gate116inter9, gate116inter10, gate116inter11, gate116inter12, gate239inter0, gate239inter1, gate239inter2, gate239inter3, gate239inter4, gate239inter5, gate239inter6, gate239inter7, gate239inter8, gate239inter9, gate239inter10, gate239inter11, gate239inter12, gate187inter0, gate187inter1, gate187inter2, gate187inter3, gate187inter4, gate187inter5, gate187inter6, gate187inter7, gate187inter8, gate187inter9, gate187inter10, gate187inter11, gate187inter12, gate74inter0, gate74inter1, gate74inter2, gate74inter3, gate74inter4, gate74inter5, gate74inter6, gate74inter7, gate74inter8, gate74inter9, gate74inter10, gate74inter11, gate74inter12, gate223inter0, gate223inter1, gate223inter2, gate223inter3, gate223inter4, gate223inter5, gate223inter6, gate223inter7, gate223inter8, gate223inter9, gate223inter10, gate223inter11, gate223inter12, gate479inter0, gate479inter1, gate479inter2, gate479inter3, gate479inter4, gate479inter5, gate479inter6, gate479inter7, gate479inter8, gate479inter9, gate479inter10, gate479inter11, gate479inter12, gate67inter0, gate67inter1, gate67inter2, gate67inter3, gate67inter4, gate67inter5, gate67inter6, gate67inter7, gate67inter8, gate67inter9, gate67inter10, gate67inter11, gate67inter12, gate494inter0, gate494inter1, gate494inter2, gate494inter3, gate494inter4, gate494inter5, gate494inter6, gate494inter7, gate494inter8, gate494inter9, gate494inter10, gate494inter11, gate494inter12, gate512inter0, gate512inter1, gate512inter2, gate512inter3, gate512inter4, gate512inter5, gate512inter6, gate512inter7, gate512inter8, gate512inter9, gate512inter10, gate512inter11, gate512inter12, gate198inter0, gate198inter1, gate198inter2, gate198inter3, gate198inter4, gate198inter5, gate198inter6, gate198inter7, gate198inter8, gate198inter9, gate198inter10, gate198inter11, gate198inter12, gate250inter0, gate250inter1, gate250inter2, gate250inter3, gate250inter4, gate250inter5, gate250inter6, gate250inter7, gate250inter8, gate250inter9, gate250inter10, gate250inter11, gate250inter12, gate437inter0, gate437inter1, gate437inter2, gate437inter3, gate437inter4, gate437inter5, gate437inter6, gate437inter7, gate437inter8, gate437inter9, gate437inter10, gate437inter11, gate437inter12, gate432inter0, gate432inter1, gate432inter2, gate432inter3, gate432inter4, gate432inter5, gate432inter6, gate432inter7, gate432inter8, gate432inter9, gate432inter10, gate432inter11, gate432inter12, gate497inter0, gate497inter1, gate497inter2, gate497inter3, gate497inter4, gate497inter5, gate497inter6, gate497inter7, gate497inter8, gate497inter9, gate497inter10, gate497inter11, gate497inter12, gate291inter0, gate291inter1, gate291inter2, gate291inter3, gate291inter4, gate291inter5, gate291inter6, gate291inter7, gate291inter8, gate291inter9, gate291inter10, gate291inter11, gate291inter12, gate261inter0, gate261inter1, gate261inter2, gate261inter3, gate261inter4, gate261inter5, gate261inter6, gate261inter7, gate261inter8, gate261inter9, gate261inter10, gate261inter11, gate261inter12, gate191inter0, gate191inter1, gate191inter2, gate191inter3, gate191inter4, gate191inter5, gate191inter6, gate191inter7, gate191inter8, gate191inter9, gate191inter10, gate191inter11, gate191inter12, gate81inter0, gate81inter1, gate81inter2, gate81inter3, gate81inter4, gate81inter5, gate81inter6, gate81inter7, gate81inter8, gate81inter9, gate81inter10, gate81inter11, gate81inter12, gate138inter0, gate138inter1, gate138inter2, gate138inter3, gate138inter4, gate138inter5, gate138inter6, gate138inter7, gate138inter8, gate138inter9, gate138inter10, gate138inter11, gate138inter12;



and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );
nand2 gate9( .a(G1), .b(G2), .O(G266) );
nand2 gate10( .a(G3), .b(G4), .O(G269) );
nand2 gate11( .a(G5), .b(G6), .O(G272) );
nand2 gate12( .a(G7), .b(G8), .O(G275) );
nand2 gate13( .a(G9), .b(G10), .O(G278) );

  xor2  gate1373(.a(G12), .b(G11), .O(gate14inter0));
  nand2 gate1374(.a(gate14inter0), .b(s_118), .O(gate14inter1));
  and2  gate1375(.a(G12), .b(G11), .O(gate14inter2));
  inv1  gate1376(.a(s_118), .O(gate14inter3));
  inv1  gate1377(.a(s_119), .O(gate14inter4));
  nand2 gate1378(.a(gate14inter4), .b(gate14inter3), .O(gate14inter5));
  nor2  gate1379(.a(gate14inter5), .b(gate14inter2), .O(gate14inter6));
  inv1  gate1380(.a(G11), .O(gate14inter7));
  inv1  gate1381(.a(G12), .O(gate14inter8));
  nand2 gate1382(.a(gate14inter8), .b(gate14inter7), .O(gate14inter9));
  nand2 gate1383(.a(s_119), .b(gate14inter3), .O(gate14inter10));
  nor2  gate1384(.a(gate14inter10), .b(gate14inter9), .O(gate14inter11));
  nor2  gate1385(.a(gate14inter11), .b(gate14inter6), .O(gate14inter12));
  nand2 gate1386(.a(gate14inter12), .b(gate14inter1), .O(G281));
nand2 gate15( .a(G13), .b(G14), .O(G284) );
nand2 gate16( .a(G15), .b(G16), .O(G287) );

  xor2  gate1821(.a(G18), .b(G17), .O(gate17inter0));
  nand2 gate1822(.a(gate17inter0), .b(s_182), .O(gate17inter1));
  and2  gate1823(.a(G18), .b(G17), .O(gate17inter2));
  inv1  gate1824(.a(s_182), .O(gate17inter3));
  inv1  gate1825(.a(s_183), .O(gate17inter4));
  nand2 gate1826(.a(gate17inter4), .b(gate17inter3), .O(gate17inter5));
  nor2  gate1827(.a(gate17inter5), .b(gate17inter2), .O(gate17inter6));
  inv1  gate1828(.a(G17), .O(gate17inter7));
  inv1  gate1829(.a(G18), .O(gate17inter8));
  nand2 gate1830(.a(gate17inter8), .b(gate17inter7), .O(gate17inter9));
  nand2 gate1831(.a(s_183), .b(gate17inter3), .O(gate17inter10));
  nor2  gate1832(.a(gate17inter10), .b(gate17inter9), .O(gate17inter11));
  nor2  gate1833(.a(gate17inter11), .b(gate17inter6), .O(gate17inter12));
  nand2 gate1834(.a(gate17inter12), .b(gate17inter1), .O(G290));
nand2 gate18( .a(G19), .b(G20), .O(G293) );
nand2 gate19( .a(G21), .b(G22), .O(G296) );
nand2 gate20( .a(G23), .b(G24), .O(G299) );
nand2 gate21( .a(G25), .b(G26), .O(G302) );

  xor2  gate1387(.a(G28), .b(G27), .O(gate22inter0));
  nand2 gate1388(.a(gate22inter0), .b(s_120), .O(gate22inter1));
  and2  gate1389(.a(G28), .b(G27), .O(gate22inter2));
  inv1  gate1390(.a(s_120), .O(gate22inter3));
  inv1  gate1391(.a(s_121), .O(gate22inter4));
  nand2 gate1392(.a(gate22inter4), .b(gate22inter3), .O(gate22inter5));
  nor2  gate1393(.a(gate22inter5), .b(gate22inter2), .O(gate22inter6));
  inv1  gate1394(.a(G27), .O(gate22inter7));
  inv1  gate1395(.a(G28), .O(gate22inter8));
  nand2 gate1396(.a(gate22inter8), .b(gate22inter7), .O(gate22inter9));
  nand2 gate1397(.a(s_121), .b(gate22inter3), .O(gate22inter10));
  nor2  gate1398(.a(gate22inter10), .b(gate22inter9), .O(gate22inter11));
  nor2  gate1399(.a(gate22inter11), .b(gate22inter6), .O(gate22inter12));
  nand2 gate1400(.a(gate22inter12), .b(gate22inter1), .O(G305));
nand2 gate23( .a(G29), .b(G30), .O(G308) );

  xor2  gate883(.a(G32), .b(G31), .O(gate24inter0));
  nand2 gate884(.a(gate24inter0), .b(s_48), .O(gate24inter1));
  and2  gate885(.a(G32), .b(G31), .O(gate24inter2));
  inv1  gate886(.a(s_48), .O(gate24inter3));
  inv1  gate887(.a(s_49), .O(gate24inter4));
  nand2 gate888(.a(gate24inter4), .b(gate24inter3), .O(gate24inter5));
  nor2  gate889(.a(gate24inter5), .b(gate24inter2), .O(gate24inter6));
  inv1  gate890(.a(G31), .O(gate24inter7));
  inv1  gate891(.a(G32), .O(gate24inter8));
  nand2 gate892(.a(gate24inter8), .b(gate24inter7), .O(gate24inter9));
  nand2 gate893(.a(s_49), .b(gate24inter3), .O(gate24inter10));
  nor2  gate894(.a(gate24inter10), .b(gate24inter9), .O(gate24inter11));
  nor2  gate895(.a(gate24inter11), .b(gate24inter6), .O(gate24inter12));
  nand2 gate896(.a(gate24inter12), .b(gate24inter1), .O(G311));

  xor2  gate1807(.a(G5), .b(G1), .O(gate25inter0));
  nand2 gate1808(.a(gate25inter0), .b(s_180), .O(gate25inter1));
  and2  gate1809(.a(G5), .b(G1), .O(gate25inter2));
  inv1  gate1810(.a(s_180), .O(gate25inter3));
  inv1  gate1811(.a(s_181), .O(gate25inter4));
  nand2 gate1812(.a(gate25inter4), .b(gate25inter3), .O(gate25inter5));
  nor2  gate1813(.a(gate25inter5), .b(gate25inter2), .O(gate25inter6));
  inv1  gate1814(.a(G1), .O(gate25inter7));
  inv1  gate1815(.a(G5), .O(gate25inter8));
  nand2 gate1816(.a(gate25inter8), .b(gate25inter7), .O(gate25inter9));
  nand2 gate1817(.a(s_181), .b(gate25inter3), .O(gate25inter10));
  nor2  gate1818(.a(gate25inter10), .b(gate25inter9), .O(gate25inter11));
  nor2  gate1819(.a(gate25inter11), .b(gate25inter6), .O(gate25inter12));
  nand2 gate1820(.a(gate25inter12), .b(gate25inter1), .O(G314));
nand2 gate26( .a(G9), .b(G13), .O(G317) );
nand2 gate27( .a(G2), .b(G6), .O(G320) );
nand2 gate28( .a(G10), .b(G14), .O(G323) );
nand2 gate29( .a(G3), .b(G7), .O(G326) );
nand2 gate30( .a(G11), .b(G15), .O(G329) );

  xor2  gate1415(.a(G8), .b(G4), .O(gate31inter0));
  nand2 gate1416(.a(gate31inter0), .b(s_124), .O(gate31inter1));
  and2  gate1417(.a(G8), .b(G4), .O(gate31inter2));
  inv1  gate1418(.a(s_124), .O(gate31inter3));
  inv1  gate1419(.a(s_125), .O(gate31inter4));
  nand2 gate1420(.a(gate31inter4), .b(gate31inter3), .O(gate31inter5));
  nor2  gate1421(.a(gate31inter5), .b(gate31inter2), .O(gate31inter6));
  inv1  gate1422(.a(G4), .O(gate31inter7));
  inv1  gate1423(.a(G8), .O(gate31inter8));
  nand2 gate1424(.a(gate31inter8), .b(gate31inter7), .O(gate31inter9));
  nand2 gate1425(.a(s_125), .b(gate31inter3), .O(gate31inter10));
  nor2  gate1426(.a(gate31inter10), .b(gate31inter9), .O(gate31inter11));
  nor2  gate1427(.a(gate31inter11), .b(gate31inter6), .O(gate31inter12));
  nand2 gate1428(.a(gate31inter12), .b(gate31inter1), .O(G332));

  xor2  gate785(.a(G16), .b(G12), .O(gate32inter0));
  nand2 gate786(.a(gate32inter0), .b(s_34), .O(gate32inter1));
  and2  gate787(.a(G16), .b(G12), .O(gate32inter2));
  inv1  gate788(.a(s_34), .O(gate32inter3));
  inv1  gate789(.a(s_35), .O(gate32inter4));
  nand2 gate790(.a(gate32inter4), .b(gate32inter3), .O(gate32inter5));
  nor2  gate791(.a(gate32inter5), .b(gate32inter2), .O(gate32inter6));
  inv1  gate792(.a(G12), .O(gate32inter7));
  inv1  gate793(.a(G16), .O(gate32inter8));
  nand2 gate794(.a(gate32inter8), .b(gate32inter7), .O(gate32inter9));
  nand2 gate795(.a(s_35), .b(gate32inter3), .O(gate32inter10));
  nor2  gate796(.a(gate32inter10), .b(gate32inter9), .O(gate32inter11));
  nor2  gate797(.a(gate32inter11), .b(gate32inter6), .O(gate32inter12));
  nand2 gate798(.a(gate32inter12), .b(gate32inter1), .O(G335));

  xor2  gate1597(.a(G21), .b(G17), .O(gate33inter0));
  nand2 gate1598(.a(gate33inter0), .b(s_150), .O(gate33inter1));
  and2  gate1599(.a(G21), .b(G17), .O(gate33inter2));
  inv1  gate1600(.a(s_150), .O(gate33inter3));
  inv1  gate1601(.a(s_151), .O(gate33inter4));
  nand2 gate1602(.a(gate33inter4), .b(gate33inter3), .O(gate33inter5));
  nor2  gate1603(.a(gate33inter5), .b(gate33inter2), .O(gate33inter6));
  inv1  gate1604(.a(G17), .O(gate33inter7));
  inv1  gate1605(.a(G21), .O(gate33inter8));
  nand2 gate1606(.a(gate33inter8), .b(gate33inter7), .O(gate33inter9));
  nand2 gate1607(.a(s_151), .b(gate33inter3), .O(gate33inter10));
  nor2  gate1608(.a(gate33inter10), .b(gate33inter9), .O(gate33inter11));
  nor2  gate1609(.a(gate33inter11), .b(gate33inter6), .O(gate33inter12));
  nand2 gate1610(.a(gate33inter12), .b(gate33inter1), .O(G338));

  xor2  gate1471(.a(G29), .b(G25), .O(gate34inter0));
  nand2 gate1472(.a(gate34inter0), .b(s_132), .O(gate34inter1));
  and2  gate1473(.a(G29), .b(G25), .O(gate34inter2));
  inv1  gate1474(.a(s_132), .O(gate34inter3));
  inv1  gate1475(.a(s_133), .O(gate34inter4));
  nand2 gate1476(.a(gate34inter4), .b(gate34inter3), .O(gate34inter5));
  nor2  gate1477(.a(gate34inter5), .b(gate34inter2), .O(gate34inter6));
  inv1  gate1478(.a(G25), .O(gate34inter7));
  inv1  gate1479(.a(G29), .O(gate34inter8));
  nand2 gate1480(.a(gate34inter8), .b(gate34inter7), .O(gate34inter9));
  nand2 gate1481(.a(s_133), .b(gate34inter3), .O(gate34inter10));
  nor2  gate1482(.a(gate34inter10), .b(gate34inter9), .O(gate34inter11));
  nor2  gate1483(.a(gate34inter11), .b(gate34inter6), .O(gate34inter12));
  nand2 gate1484(.a(gate34inter12), .b(gate34inter1), .O(G341));

  xor2  gate771(.a(G22), .b(G18), .O(gate35inter0));
  nand2 gate772(.a(gate35inter0), .b(s_32), .O(gate35inter1));
  and2  gate773(.a(G22), .b(G18), .O(gate35inter2));
  inv1  gate774(.a(s_32), .O(gate35inter3));
  inv1  gate775(.a(s_33), .O(gate35inter4));
  nand2 gate776(.a(gate35inter4), .b(gate35inter3), .O(gate35inter5));
  nor2  gate777(.a(gate35inter5), .b(gate35inter2), .O(gate35inter6));
  inv1  gate778(.a(G18), .O(gate35inter7));
  inv1  gate779(.a(G22), .O(gate35inter8));
  nand2 gate780(.a(gate35inter8), .b(gate35inter7), .O(gate35inter9));
  nand2 gate781(.a(s_33), .b(gate35inter3), .O(gate35inter10));
  nor2  gate782(.a(gate35inter10), .b(gate35inter9), .O(gate35inter11));
  nor2  gate783(.a(gate35inter11), .b(gate35inter6), .O(gate35inter12));
  nand2 gate784(.a(gate35inter12), .b(gate35inter1), .O(G344));
nand2 gate36( .a(G26), .b(G30), .O(G347) );

  xor2  gate967(.a(G23), .b(G19), .O(gate37inter0));
  nand2 gate968(.a(gate37inter0), .b(s_60), .O(gate37inter1));
  and2  gate969(.a(G23), .b(G19), .O(gate37inter2));
  inv1  gate970(.a(s_60), .O(gate37inter3));
  inv1  gate971(.a(s_61), .O(gate37inter4));
  nand2 gate972(.a(gate37inter4), .b(gate37inter3), .O(gate37inter5));
  nor2  gate973(.a(gate37inter5), .b(gate37inter2), .O(gate37inter6));
  inv1  gate974(.a(G19), .O(gate37inter7));
  inv1  gate975(.a(G23), .O(gate37inter8));
  nand2 gate976(.a(gate37inter8), .b(gate37inter7), .O(gate37inter9));
  nand2 gate977(.a(s_61), .b(gate37inter3), .O(gate37inter10));
  nor2  gate978(.a(gate37inter10), .b(gate37inter9), .O(gate37inter11));
  nor2  gate979(.a(gate37inter11), .b(gate37inter6), .O(gate37inter12));
  nand2 gate980(.a(gate37inter12), .b(gate37inter1), .O(G350));
nand2 gate38( .a(G27), .b(G31), .O(G353) );
nand2 gate39( .a(G20), .b(G24), .O(G356) );
nand2 gate40( .a(G28), .b(G32), .O(G359) );

  xor2  gate729(.a(G266), .b(G1), .O(gate41inter0));
  nand2 gate730(.a(gate41inter0), .b(s_26), .O(gate41inter1));
  and2  gate731(.a(G266), .b(G1), .O(gate41inter2));
  inv1  gate732(.a(s_26), .O(gate41inter3));
  inv1  gate733(.a(s_27), .O(gate41inter4));
  nand2 gate734(.a(gate41inter4), .b(gate41inter3), .O(gate41inter5));
  nor2  gate735(.a(gate41inter5), .b(gate41inter2), .O(gate41inter6));
  inv1  gate736(.a(G1), .O(gate41inter7));
  inv1  gate737(.a(G266), .O(gate41inter8));
  nand2 gate738(.a(gate41inter8), .b(gate41inter7), .O(gate41inter9));
  nand2 gate739(.a(s_27), .b(gate41inter3), .O(gate41inter10));
  nor2  gate740(.a(gate41inter10), .b(gate41inter9), .O(gate41inter11));
  nor2  gate741(.a(gate41inter11), .b(gate41inter6), .O(gate41inter12));
  nand2 gate742(.a(gate41inter12), .b(gate41inter1), .O(G362));
nand2 gate42( .a(G2), .b(G266), .O(G363) );
nand2 gate43( .a(G3), .b(G269), .O(G364) );
nand2 gate44( .a(G4), .b(G269), .O(G365) );
nand2 gate45( .a(G5), .b(G272), .O(G366) );
nand2 gate46( .a(G6), .b(G272), .O(G367) );
nand2 gate47( .a(G7), .b(G275), .O(G368) );
nand2 gate48( .a(G8), .b(G275), .O(G369) );
nand2 gate49( .a(G9), .b(G278), .O(G370) );
nand2 gate50( .a(G10), .b(G278), .O(G371) );

  xor2  gate1555(.a(G281), .b(G11), .O(gate51inter0));
  nand2 gate1556(.a(gate51inter0), .b(s_144), .O(gate51inter1));
  and2  gate1557(.a(G281), .b(G11), .O(gate51inter2));
  inv1  gate1558(.a(s_144), .O(gate51inter3));
  inv1  gate1559(.a(s_145), .O(gate51inter4));
  nand2 gate1560(.a(gate51inter4), .b(gate51inter3), .O(gate51inter5));
  nor2  gate1561(.a(gate51inter5), .b(gate51inter2), .O(gate51inter6));
  inv1  gate1562(.a(G11), .O(gate51inter7));
  inv1  gate1563(.a(G281), .O(gate51inter8));
  nand2 gate1564(.a(gate51inter8), .b(gate51inter7), .O(gate51inter9));
  nand2 gate1565(.a(s_145), .b(gate51inter3), .O(gate51inter10));
  nor2  gate1566(.a(gate51inter10), .b(gate51inter9), .O(gate51inter11));
  nor2  gate1567(.a(gate51inter11), .b(gate51inter6), .O(gate51inter12));
  nand2 gate1568(.a(gate51inter12), .b(gate51inter1), .O(G372));
nand2 gate52( .a(G12), .b(G281), .O(G373) );
nand2 gate53( .a(G13), .b(G284), .O(G374) );

  xor2  gate1247(.a(G284), .b(G14), .O(gate54inter0));
  nand2 gate1248(.a(gate54inter0), .b(s_100), .O(gate54inter1));
  and2  gate1249(.a(G284), .b(G14), .O(gate54inter2));
  inv1  gate1250(.a(s_100), .O(gate54inter3));
  inv1  gate1251(.a(s_101), .O(gate54inter4));
  nand2 gate1252(.a(gate54inter4), .b(gate54inter3), .O(gate54inter5));
  nor2  gate1253(.a(gate54inter5), .b(gate54inter2), .O(gate54inter6));
  inv1  gate1254(.a(G14), .O(gate54inter7));
  inv1  gate1255(.a(G284), .O(gate54inter8));
  nand2 gate1256(.a(gate54inter8), .b(gate54inter7), .O(gate54inter9));
  nand2 gate1257(.a(s_101), .b(gate54inter3), .O(gate54inter10));
  nor2  gate1258(.a(gate54inter10), .b(gate54inter9), .O(gate54inter11));
  nor2  gate1259(.a(gate54inter11), .b(gate54inter6), .O(gate54inter12));
  nand2 gate1260(.a(gate54inter12), .b(gate54inter1), .O(G375));
nand2 gate55( .a(G15), .b(G287), .O(G376) );

  xor2  gate701(.a(G287), .b(G16), .O(gate56inter0));
  nand2 gate702(.a(gate56inter0), .b(s_22), .O(gate56inter1));
  and2  gate703(.a(G287), .b(G16), .O(gate56inter2));
  inv1  gate704(.a(s_22), .O(gate56inter3));
  inv1  gate705(.a(s_23), .O(gate56inter4));
  nand2 gate706(.a(gate56inter4), .b(gate56inter3), .O(gate56inter5));
  nor2  gate707(.a(gate56inter5), .b(gate56inter2), .O(gate56inter6));
  inv1  gate708(.a(G16), .O(gate56inter7));
  inv1  gate709(.a(G287), .O(gate56inter8));
  nand2 gate710(.a(gate56inter8), .b(gate56inter7), .O(gate56inter9));
  nand2 gate711(.a(s_23), .b(gate56inter3), .O(gate56inter10));
  nor2  gate712(.a(gate56inter10), .b(gate56inter9), .O(gate56inter11));
  nor2  gate713(.a(gate56inter11), .b(gate56inter6), .O(gate56inter12));
  nand2 gate714(.a(gate56inter12), .b(gate56inter1), .O(G377));
nand2 gate57( .a(G17), .b(G290), .O(G378) );
nand2 gate58( .a(G18), .b(G290), .O(G379) );
nand2 gate59( .a(G19), .b(G293), .O(G380) );
nand2 gate60( .a(G20), .b(G293), .O(G381) );
nand2 gate61( .a(G21), .b(G296), .O(G382) );
nand2 gate62( .a(G22), .b(G296), .O(G383) );

  xor2  gate1695(.a(G299), .b(G23), .O(gate63inter0));
  nand2 gate1696(.a(gate63inter0), .b(s_164), .O(gate63inter1));
  and2  gate1697(.a(G299), .b(G23), .O(gate63inter2));
  inv1  gate1698(.a(s_164), .O(gate63inter3));
  inv1  gate1699(.a(s_165), .O(gate63inter4));
  nand2 gate1700(.a(gate63inter4), .b(gate63inter3), .O(gate63inter5));
  nor2  gate1701(.a(gate63inter5), .b(gate63inter2), .O(gate63inter6));
  inv1  gate1702(.a(G23), .O(gate63inter7));
  inv1  gate1703(.a(G299), .O(gate63inter8));
  nand2 gate1704(.a(gate63inter8), .b(gate63inter7), .O(gate63inter9));
  nand2 gate1705(.a(s_165), .b(gate63inter3), .O(gate63inter10));
  nor2  gate1706(.a(gate63inter10), .b(gate63inter9), .O(gate63inter11));
  nor2  gate1707(.a(gate63inter11), .b(gate63inter6), .O(gate63inter12));
  nand2 gate1708(.a(gate63inter12), .b(gate63inter1), .O(G384));
nand2 gate64( .a(G24), .b(G299), .O(G385) );

  xor2  gate939(.a(G302), .b(G25), .O(gate65inter0));
  nand2 gate940(.a(gate65inter0), .b(s_56), .O(gate65inter1));
  and2  gate941(.a(G302), .b(G25), .O(gate65inter2));
  inv1  gate942(.a(s_56), .O(gate65inter3));
  inv1  gate943(.a(s_57), .O(gate65inter4));
  nand2 gate944(.a(gate65inter4), .b(gate65inter3), .O(gate65inter5));
  nor2  gate945(.a(gate65inter5), .b(gate65inter2), .O(gate65inter6));
  inv1  gate946(.a(G25), .O(gate65inter7));
  inv1  gate947(.a(G302), .O(gate65inter8));
  nand2 gate948(.a(gate65inter8), .b(gate65inter7), .O(gate65inter9));
  nand2 gate949(.a(s_57), .b(gate65inter3), .O(gate65inter10));
  nor2  gate950(.a(gate65inter10), .b(gate65inter9), .O(gate65inter11));
  nor2  gate951(.a(gate65inter11), .b(gate65inter6), .O(gate65inter12));
  nand2 gate952(.a(gate65inter12), .b(gate65inter1), .O(G386));
nand2 gate66( .a(G26), .b(G302), .O(G387) );

  xor2  gate1919(.a(G305), .b(G27), .O(gate67inter0));
  nand2 gate1920(.a(gate67inter0), .b(s_196), .O(gate67inter1));
  and2  gate1921(.a(G305), .b(G27), .O(gate67inter2));
  inv1  gate1922(.a(s_196), .O(gate67inter3));
  inv1  gate1923(.a(s_197), .O(gate67inter4));
  nand2 gate1924(.a(gate67inter4), .b(gate67inter3), .O(gate67inter5));
  nor2  gate1925(.a(gate67inter5), .b(gate67inter2), .O(gate67inter6));
  inv1  gate1926(.a(G27), .O(gate67inter7));
  inv1  gate1927(.a(G305), .O(gate67inter8));
  nand2 gate1928(.a(gate67inter8), .b(gate67inter7), .O(gate67inter9));
  nand2 gate1929(.a(s_197), .b(gate67inter3), .O(gate67inter10));
  nor2  gate1930(.a(gate67inter10), .b(gate67inter9), .O(gate67inter11));
  nor2  gate1931(.a(gate67inter11), .b(gate67inter6), .O(gate67inter12));
  nand2 gate1932(.a(gate67inter12), .b(gate67inter1), .O(G388));
nand2 gate68( .a(G28), .b(G305), .O(G389) );
nand2 gate69( .a(G29), .b(G308), .O(G390) );

  xor2  gate1639(.a(G308), .b(G30), .O(gate70inter0));
  nand2 gate1640(.a(gate70inter0), .b(s_156), .O(gate70inter1));
  and2  gate1641(.a(G308), .b(G30), .O(gate70inter2));
  inv1  gate1642(.a(s_156), .O(gate70inter3));
  inv1  gate1643(.a(s_157), .O(gate70inter4));
  nand2 gate1644(.a(gate70inter4), .b(gate70inter3), .O(gate70inter5));
  nor2  gate1645(.a(gate70inter5), .b(gate70inter2), .O(gate70inter6));
  inv1  gate1646(.a(G30), .O(gate70inter7));
  inv1  gate1647(.a(G308), .O(gate70inter8));
  nand2 gate1648(.a(gate70inter8), .b(gate70inter7), .O(gate70inter9));
  nand2 gate1649(.a(s_157), .b(gate70inter3), .O(gate70inter10));
  nor2  gate1650(.a(gate70inter10), .b(gate70inter9), .O(gate70inter11));
  nor2  gate1651(.a(gate70inter11), .b(gate70inter6), .O(gate70inter12));
  nand2 gate1652(.a(gate70inter12), .b(gate70inter1), .O(G391));

  xor2  gate813(.a(G311), .b(G31), .O(gate71inter0));
  nand2 gate814(.a(gate71inter0), .b(s_38), .O(gate71inter1));
  and2  gate815(.a(G311), .b(G31), .O(gate71inter2));
  inv1  gate816(.a(s_38), .O(gate71inter3));
  inv1  gate817(.a(s_39), .O(gate71inter4));
  nand2 gate818(.a(gate71inter4), .b(gate71inter3), .O(gate71inter5));
  nor2  gate819(.a(gate71inter5), .b(gate71inter2), .O(gate71inter6));
  inv1  gate820(.a(G31), .O(gate71inter7));
  inv1  gate821(.a(G311), .O(gate71inter8));
  nand2 gate822(.a(gate71inter8), .b(gate71inter7), .O(gate71inter9));
  nand2 gate823(.a(s_39), .b(gate71inter3), .O(gate71inter10));
  nor2  gate824(.a(gate71inter10), .b(gate71inter9), .O(gate71inter11));
  nor2  gate825(.a(gate71inter11), .b(gate71inter6), .O(gate71inter12));
  nand2 gate826(.a(gate71inter12), .b(gate71inter1), .O(G392));

  xor2  gate1737(.a(G311), .b(G32), .O(gate72inter0));
  nand2 gate1738(.a(gate72inter0), .b(s_170), .O(gate72inter1));
  and2  gate1739(.a(G311), .b(G32), .O(gate72inter2));
  inv1  gate1740(.a(s_170), .O(gate72inter3));
  inv1  gate1741(.a(s_171), .O(gate72inter4));
  nand2 gate1742(.a(gate72inter4), .b(gate72inter3), .O(gate72inter5));
  nor2  gate1743(.a(gate72inter5), .b(gate72inter2), .O(gate72inter6));
  inv1  gate1744(.a(G32), .O(gate72inter7));
  inv1  gate1745(.a(G311), .O(gate72inter8));
  nand2 gate1746(.a(gate72inter8), .b(gate72inter7), .O(gate72inter9));
  nand2 gate1747(.a(s_171), .b(gate72inter3), .O(gate72inter10));
  nor2  gate1748(.a(gate72inter10), .b(gate72inter9), .O(gate72inter11));
  nor2  gate1749(.a(gate72inter11), .b(gate72inter6), .O(gate72inter12));
  nand2 gate1750(.a(gate72inter12), .b(gate72inter1), .O(G393));

  xor2  gate561(.a(G314), .b(G1), .O(gate73inter0));
  nand2 gate562(.a(gate73inter0), .b(s_2), .O(gate73inter1));
  and2  gate563(.a(G314), .b(G1), .O(gate73inter2));
  inv1  gate564(.a(s_2), .O(gate73inter3));
  inv1  gate565(.a(s_3), .O(gate73inter4));
  nand2 gate566(.a(gate73inter4), .b(gate73inter3), .O(gate73inter5));
  nor2  gate567(.a(gate73inter5), .b(gate73inter2), .O(gate73inter6));
  inv1  gate568(.a(G1), .O(gate73inter7));
  inv1  gate569(.a(G314), .O(gate73inter8));
  nand2 gate570(.a(gate73inter8), .b(gate73inter7), .O(gate73inter9));
  nand2 gate571(.a(s_3), .b(gate73inter3), .O(gate73inter10));
  nor2  gate572(.a(gate73inter10), .b(gate73inter9), .O(gate73inter11));
  nor2  gate573(.a(gate73inter11), .b(gate73inter6), .O(gate73inter12));
  nand2 gate574(.a(gate73inter12), .b(gate73inter1), .O(G394));

  xor2  gate1877(.a(G314), .b(G5), .O(gate74inter0));
  nand2 gate1878(.a(gate74inter0), .b(s_190), .O(gate74inter1));
  and2  gate1879(.a(G314), .b(G5), .O(gate74inter2));
  inv1  gate1880(.a(s_190), .O(gate74inter3));
  inv1  gate1881(.a(s_191), .O(gate74inter4));
  nand2 gate1882(.a(gate74inter4), .b(gate74inter3), .O(gate74inter5));
  nor2  gate1883(.a(gate74inter5), .b(gate74inter2), .O(gate74inter6));
  inv1  gate1884(.a(G5), .O(gate74inter7));
  inv1  gate1885(.a(G314), .O(gate74inter8));
  nand2 gate1886(.a(gate74inter8), .b(gate74inter7), .O(gate74inter9));
  nand2 gate1887(.a(s_191), .b(gate74inter3), .O(gate74inter10));
  nor2  gate1888(.a(gate74inter10), .b(gate74inter9), .O(gate74inter11));
  nor2  gate1889(.a(gate74inter11), .b(gate74inter6), .O(gate74inter12));
  nand2 gate1890(.a(gate74inter12), .b(gate74inter1), .O(G395));
nand2 gate75( .a(G9), .b(G317), .O(G396) );
nand2 gate76( .a(G13), .b(G317), .O(G397) );

  xor2  gate897(.a(G320), .b(G2), .O(gate77inter0));
  nand2 gate898(.a(gate77inter0), .b(s_50), .O(gate77inter1));
  and2  gate899(.a(G320), .b(G2), .O(gate77inter2));
  inv1  gate900(.a(s_50), .O(gate77inter3));
  inv1  gate901(.a(s_51), .O(gate77inter4));
  nand2 gate902(.a(gate77inter4), .b(gate77inter3), .O(gate77inter5));
  nor2  gate903(.a(gate77inter5), .b(gate77inter2), .O(gate77inter6));
  inv1  gate904(.a(G2), .O(gate77inter7));
  inv1  gate905(.a(G320), .O(gate77inter8));
  nand2 gate906(.a(gate77inter8), .b(gate77inter7), .O(gate77inter9));
  nand2 gate907(.a(s_51), .b(gate77inter3), .O(gate77inter10));
  nor2  gate908(.a(gate77inter10), .b(gate77inter9), .O(gate77inter11));
  nor2  gate909(.a(gate77inter11), .b(gate77inter6), .O(gate77inter12));
  nand2 gate910(.a(gate77inter12), .b(gate77inter1), .O(G398));
nand2 gate78( .a(G6), .b(G320), .O(G399) );

  xor2  gate1583(.a(G323), .b(G10), .O(gate79inter0));
  nand2 gate1584(.a(gate79inter0), .b(s_148), .O(gate79inter1));
  and2  gate1585(.a(G323), .b(G10), .O(gate79inter2));
  inv1  gate1586(.a(s_148), .O(gate79inter3));
  inv1  gate1587(.a(s_149), .O(gate79inter4));
  nand2 gate1588(.a(gate79inter4), .b(gate79inter3), .O(gate79inter5));
  nor2  gate1589(.a(gate79inter5), .b(gate79inter2), .O(gate79inter6));
  inv1  gate1590(.a(G10), .O(gate79inter7));
  inv1  gate1591(.a(G323), .O(gate79inter8));
  nand2 gate1592(.a(gate79inter8), .b(gate79inter7), .O(gate79inter9));
  nand2 gate1593(.a(s_149), .b(gate79inter3), .O(gate79inter10));
  nor2  gate1594(.a(gate79inter10), .b(gate79inter9), .O(gate79inter11));
  nor2  gate1595(.a(gate79inter11), .b(gate79inter6), .O(gate79inter12));
  nand2 gate1596(.a(gate79inter12), .b(gate79inter1), .O(G400));
nand2 gate80( .a(G14), .b(G323), .O(G401) );

  xor2  gate2073(.a(G326), .b(G3), .O(gate81inter0));
  nand2 gate2074(.a(gate81inter0), .b(s_218), .O(gate81inter1));
  and2  gate2075(.a(G326), .b(G3), .O(gate81inter2));
  inv1  gate2076(.a(s_218), .O(gate81inter3));
  inv1  gate2077(.a(s_219), .O(gate81inter4));
  nand2 gate2078(.a(gate81inter4), .b(gate81inter3), .O(gate81inter5));
  nor2  gate2079(.a(gate81inter5), .b(gate81inter2), .O(gate81inter6));
  inv1  gate2080(.a(G3), .O(gate81inter7));
  inv1  gate2081(.a(G326), .O(gate81inter8));
  nand2 gate2082(.a(gate81inter8), .b(gate81inter7), .O(gate81inter9));
  nand2 gate2083(.a(s_219), .b(gate81inter3), .O(gate81inter10));
  nor2  gate2084(.a(gate81inter10), .b(gate81inter9), .O(gate81inter11));
  nor2  gate2085(.a(gate81inter11), .b(gate81inter6), .O(gate81inter12));
  nand2 gate2086(.a(gate81inter12), .b(gate81inter1), .O(G402));
nand2 gate82( .a(G7), .b(G326), .O(G403) );
nand2 gate83( .a(G11), .b(G329), .O(G404) );

  xor2  gate1205(.a(G329), .b(G15), .O(gate84inter0));
  nand2 gate1206(.a(gate84inter0), .b(s_94), .O(gate84inter1));
  and2  gate1207(.a(G329), .b(G15), .O(gate84inter2));
  inv1  gate1208(.a(s_94), .O(gate84inter3));
  inv1  gate1209(.a(s_95), .O(gate84inter4));
  nand2 gate1210(.a(gate84inter4), .b(gate84inter3), .O(gate84inter5));
  nor2  gate1211(.a(gate84inter5), .b(gate84inter2), .O(gate84inter6));
  inv1  gate1212(.a(G15), .O(gate84inter7));
  inv1  gate1213(.a(G329), .O(gate84inter8));
  nand2 gate1214(.a(gate84inter8), .b(gate84inter7), .O(gate84inter9));
  nand2 gate1215(.a(s_95), .b(gate84inter3), .O(gate84inter10));
  nor2  gate1216(.a(gate84inter10), .b(gate84inter9), .O(gate84inter11));
  nor2  gate1217(.a(gate84inter11), .b(gate84inter6), .O(gate84inter12));
  nand2 gate1218(.a(gate84inter12), .b(gate84inter1), .O(G405));

  xor2  gate1569(.a(G332), .b(G4), .O(gate85inter0));
  nand2 gate1570(.a(gate85inter0), .b(s_146), .O(gate85inter1));
  and2  gate1571(.a(G332), .b(G4), .O(gate85inter2));
  inv1  gate1572(.a(s_146), .O(gate85inter3));
  inv1  gate1573(.a(s_147), .O(gate85inter4));
  nand2 gate1574(.a(gate85inter4), .b(gate85inter3), .O(gate85inter5));
  nor2  gate1575(.a(gate85inter5), .b(gate85inter2), .O(gate85inter6));
  inv1  gate1576(.a(G4), .O(gate85inter7));
  inv1  gate1577(.a(G332), .O(gate85inter8));
  nand2 gate1578(.a(gate85inter8), .b(gate85inter7), .O(gate85inter9));
  nand2 gate1579(.a(s_147), .b(gate85inter3), .O(gate85inter10));
  nor2  gate1580(.a(gate85inter10), .b(gate85inter9), .O(gate85inter11));
  nor2  gate1581(.a(gate85inter11), .b(gate85inter6), .O(gate85inter12));
  nand2 gate1582(.a(gate85inter12), .b(gate85inter1), .O(G406));

  xor2  gate715(.a(G332), .b(G8), .O(gate86inter0));
  nand2 gate716(.a(gate86inter0), .b(s_24), .O(gate86inter1));
  and2  gate717(.a(G332), .b(G8), .O(gate86inter2));
  inv1  gate718(.a(s_24), .O(gate86inter3));
  inv1  gate719(.a(s_25), .O(gate86inter4));
  nand2 gate720(.a(gate86inter4), .b(gate86inter3), .O(gate86inter5));
  nor2  gate721(.a(gate86inter5), .b(gate86inter2), .O(gate86inter6));
  inv1  gate722(.a(G8), .O(gate86inter7));
  inv1  gate723(.a(G332), .O(gate86inter8));
  nand2 gate724(.a(gate86inter8), .b(gate86inter7), .O(gate86inter9));
  nand2 gate725(.a(s_25), .b(gate86inter3), .O(gate86inter10));
  nor2  gate726(.a(gate86inter10), .b(gate86inter9), .O(gate86inter11));
  nor2  gate727(.a(gate86inter11), .b(gate86inter6), .O(gate86inter12));
  nand2 gate728(.a(gate86inter12), .b(gate86inter1), .O(G407));
nand2 gate87( .a(G12), .b(G335), .O(G408) );
nand2 gate88( .a(G16), .b(G335), .O(G409) );
nand2 gate89( .a(G17), .b(G338), .O(G410) );
nand2 gate90( .a(G21), .b(G338), .O(G411) );

  xor2  gate1317(.a(G341), .b(G25), .O(gate91inter0));
  nand2 gate1318(.a(gate91inter0), .b(s_110), .O(gate91inter1));
  and2  gate1319(.a(G341), .b(G25), .O(gate91inter2));
  inv1  gate1320(.a(s_110), .O(gate91inter3));
  inv1  gate1321(.a(s_111), .O(gate91inter4));
  nand2 gate1322(.a(gate91inter4), .b(gate91inter3), .O(gate91inter5));
  nor2  gate1323(.a(gate91inter5), .b(gate91inter2), .O(gate91inter6));
  inv1  gate1324(.a(G25), .O(gate91inter7));
  inv1  gate1325(.a(G341), .O(gate91inter8));
  nand2 gate1326(.a(gate91inter8), .b(gate91inter7), .O(gate91inter9));
  nand2 gate1327(.a(s_111), .b(gate91inter3), .O(gate91inter10));
  nor2  gate1328(.a(gate91inter10), .b(gate91inter9), .O(gate91inter11));
  nor2  gate1329(.a(gate91inter11), .b(gate91inter6), .O(gate91inter12));
  nand2 gate1330(.a(gate91inter12), .b(gate91inter1), .O(G412));
nand2 gate92( .a(G29), .b(G341), .O(G413) );
nand2 gate93( .a(G18), .b(G344), .O(G414) );
nand2 gate94( .a(G22), .b(G344), .O(G415) );
nand2 gate95( .a(G26), .b(G347), .O(G416) );
nand2 gate96( .a(G30), .b(G347), .O(G417) );
nand2 gate97( .a(G19), .b(G350), .O(G418) );
nand2 gate98( .a(G23), .b(G350), .O(G419) );
nand2 gate99( .a(G27), .b(G353), .O(G420) );

  xor2  gate1457(.a(G353), .b(G31), .O(gate100inter0));
  nand2 gate1458(.a(gate100inter0), .b(s_130), .O(gate100inter1));
  and2  gate1459(.a(G353), .b(G31), .O(gate100inter2));
  inv1  gate1460(.a(s_130), .O(gate100inter3));
  inv1  gate1461(.a(s_131), .O(gate100inter4));
  nand2 gate1462(.a(gate100inter4), .b(gate100inter3), .O(gate100inter5));
  nor2  gate1463(.a(gate100inter5), .b(gate100inter2), .O(gate100inter6));
  inv1  gate1464(.a(G31), .O(gate100inter7));
  inv1  gate1465(.a(G353), .O(gate100inter8));
  nand2 gate1466(.a(gate100inter8), .b(gate100inter7), .O(gate100inter9));
  nand2 gate1467(.a(s_131), .b(gate100inter3), .O(gate100inter10));
  nor2  gate1468(.a(gate100inter10), .b(gate100inter9), .O(gate100inter11));
  nor2  gate1469(.a(gate100inter11), .b(gate100inter6), .O(gate100inter12));
  nand2 gate1470(.a(gate100inter12), .b(gate100inter1), .O(G421));
nand2 gate101( .a(G20), .b(G356), .O(G422) );

  xor2  gate1527(.a(G356), .b(G24), .O(gate102inter0));
  nand2 gate1528(.a(gate102inter0), .b(s_140), .O(gate102inter1));
  and2  gate1529(.a(G356), .b(G24), .O(gate102inter2));
  inv1  gate1530(.a(s_140), .O(gate102inter3));
  inv1  gate1531(.a(s_141), .O(gate102inter4));
  nand2 gate1532(.a(gate102inter4), .b(gate102inter3), .O(gate102inter5));
  nor2  gate1533(.a(gate102inter5), .b(gate102inter2), .O(gate102inter6));
  inv1  gate1534(.a(G24), .O(gate102inter7));
  inv1  gate1535(.a(G356), .O(gate102inter8));
  nand2 gate1536(.a(gate102inter8), .b(gate102inter7), .O(gate102inter9));
  nand2 gate1537(.a(s_141), .b(gate102inter3), .O(gate102inter10));
  nor2  gate1538(.a(gate102inter10), .b(gate102inter9), .O(gate102inter11));
  nor2  gate1539(.a(gate102inter11), .b(gate102inter6), .O(gate102inter12));
  nand2 gate1540(.a(gate102inter12), .b(gate102inter1), .O(G423));
nand2 gate103( .a(G28), .b(G359), .O(G424) );
nand2 gate104( .a(G32), .b(G359), .O(G425) );
nand2 gate105( .a(G362), .b(G363), .O(G426) );
nand2 gate106( .a(G364), .b(G365), .O(G429) );
nand2 gate107( .a(G366), .b(G367), .O(G432) );

  xor2  gate1751(.a(G369), .b(G368), .O(gate108inter0));
  nand2 gate1752(.a(gate108inter0), .b(s_172), .O(gate108inter1));
  and2  gate1753(.a(G369), .b(G368), .O(gate108inter2));
  inv1  gate1754(.a(s_172), .O(gate108inter3));
  inv1  gate1755(.a(s_173), .O(gate108inter4));
  nand2 gate1756(.a(gate108inter4), .b(gate108inter3), .O(gate108inter5));
  nor2  gate1757(.a(gate108inter5), .b(gate108inter2), .O(gate108inter6));
  inv1  gate1758(.a(G368), .O(gate108inter7));
  inv1  gate1759(.a(G369), .O(gate108inter8));
  nand2 gate1760(.a(gate108inter8), .b(gate108inter7), .O(gate108inter9));
  nand2 gate1761(.a(s_173), .b(gate108inter3), .O(gate108inter10));
  nor2  gate1762(.a(gate108inter10), .b(gate108inter9), .O(gate108inter11));
  nor2  gate1763(.a(gate108inter11), .b(gate108inter6), .O(gate108inter12));
  nand2 gate1764(.a(gate108inter12), .b(gate108inter1), .O(G435));

  xor2  gate757(.a(G371), .b(G370), .O(gate109inter0));
  nand2 gate758(.a(gate109inter0), .b(s_30), .O(gate109inter1));
  and2  gate759(.a(G371), .b(G370), .O(gate109inter2));
  inv1  gate760(.a(s_30), .O(gate109inter3));
  inv1  gate761(.a(s_31), .O(gate109inter4));
  nand2 gate762(.a(gate109inter4), .b(gate109inter3), .O(gate109inter5));
  nor2  gate763(.a(gate109inter5), .b(gate109inter2), .O(gate109inter6));
  inv1  gate764(.a(G370), .O(gate109inter7));
  inv1  gate765(.a(G371), .O(gate109inter8));
  nand2 gate766(.a(gate109inter8), .b(gate109inter7), .O(gate109inter9));
  nand2 gate767(.a(s_31), .b(gate109inter3), .O(gate109inter10));
  nor2  gate768(.a(gate109inter10), .b(gate109inter9), .O(gate109inter11));
  nor2  gate769(.a(gate109inter11), .b(gate109inter6), .O(gate109inter12));
  nand2 gate770(.a(gate109inter12), .b(gate109inter1), .O(G438));
nand2 gate110( .a(G372), .b(G373), .O(G441) );

  xor2  gate1037(.a(G375), .b(G374), .O(gate111inter0));
  nand2 gate1038(.a(gate111inter0), .b(s_70), .O(gate111inter1));
  and2  gate1039(.a(G375), .b(G374), .O(gate111inter2));
  inv1  gate1040(.a(s_70), .O(gate111inter3));
  inv1  gate1041(.a(s_71), .O(gate111inter4));
  nand2 gate1042(.a(gate111inter4), .b(gate111inter3), .O(gate111inter5));
  nor2  gate1043(.a(gate111inter5), .b(gate111inter2), .O(gate111inter6));
  inv1  gate1044(.a(G374), .O(gate111inter7));
  inv1  gate1045(.a(G375), .O(gate111inter8));
  nand2 gate1046(.a(gate111inter8), .b(gate111inter7), .O(gate111inter9));
  nand2 gate1047(.a(s_71), .b(gate111inter3), .O(gate111inter10));
  nor2  gate1048(.a(gate111inter10), .b(gate111inter9), .O(gate111inter11));
  nor2  gate1049(.a(gate111inter11), .b(gate111inter6), .O(gate111inter12));
  nand2 gate1050(.a(gate111inter12), .b(gate111inter1), .O(G444));
nand2 gate112( .a(G376), .b(G377), .O(G447) );
nand2 gate113( .a(G378), .b(G379), .O(G450) );
nand2 gate114( .a(G380), .b(G381), .O(G453) );
nand2 gate115( .a(G382), .b(G383), .O(G456) );

  xor2  gate1835(.a(G385), .b(G384), .O(gate116inter0));
  nand2 gate1836(.a(gate116inter0), .b(s_184), .O(gate116inter1));
  and2  gate1837(.a(G385), .b(G384), .O(gate116inter2));
  inv1  gate1838(.a(s_184), .O(gate116inter3));
  inv1  gate1839(.a(s_185), .O(gate116inter4));
  nand2 gate1840(.a(gate116inter4), .b(gate116inter3), .O(gate116inter5));
  nor2  gate1841(.a(gate116inter5), .b(gate116inter2), .O(gate116inter6));
  inv1  gate1842(.a(G384), .O(gate116inter7));
  inv1  gate1843(.a(G385), .O(gate116inter8));
  nand2 gate1844(.a(gate116inter8), .b(gate116inter7), .O(gate116inter9));
  nand2 gate1845(.a(s_185), .b(gate116inter3), .O(gate116inter10));
  nor2  gate1846(.a(gate116inter10), .b(gate116inter9), .O(gate116inter11));
  nor2  gate1847(.a(gate116inter11), .b(gate116inter6), .O(gate116inter12));
  nand2 gate1848(.a(gate116inter12), .b(gate116inter1), .O(G459));

  xor2  gate1723(.a(G387), .b(G386), .O(gate117inter0));
  nand2 gate1724(.a(gate117inter0), .b(s_168), .O(gate117inter1));
  and2  gate1725(.a(G387), .b(G386), .O(gate117inter2));
  inv1  gate1726(.a(s_168), .O(gate117inter3));
  inv1  gate1727(.a(s_169), .O(gate117inter4));
  nand2 gate1728(.a(gate117inter4), .b(gate117inter3), .O(gate117inter5));
  nor2  gate1729(.a(gate117inter5), .b(gate117inter2), .O(gate117inter6));
  inv1  gate1730(.a(G386), .O(gate117inter7));
  inv1  gate1731(.a(G387), .O(gate117inter8));
  nand2 gate1732(.a(gate117inter8), .b(gate117inter7), .O(gate117inter9));
  nand2 gate1733(.a(s_169), .b(gate117inter3), .O(gate117inter10));
  nor2  gate1734(.a(gate117inter10), .b(gate117inter9), .O(gate117inter11));
  nor2  gate1735(.a(gate117inter11), .b(gate117inter6), .O(gate117inter12));
  nand2 gate1736(.a(gate117inter12), .b(gate117inter1), .O(G462));

  xor2  gate1177(.a(G389), .b(G388), .O(gate118inter0));
  nand2 gate1178(.a(gate118inter0), .b(s_90), .O(gate118inter1));
  and2  gate1179(.a(G389), .b(G388), .O(gate118inter2));
  inv1  gate1180(.a(s_90), .O(gate118inter3));
  inv1  gate1181(.a(s_91), .O(gate118inter4));
  nand2 gate1182(.a(gate118inter4), .b(gate118inter3), .O(gate118inter5));
  nor2  gate1183(.a(gate118inter5), .b(gate118inter2), .O(gate118inter6));
  inv1  gate1184(.a(G388), .O(gate118inter7));
  inv1  gate1185(.a(G389), .O(gate118inter8));
  nand2 gate1186(.a(gate118inter8), .b(gate118inter7), .O(gate118inter9));
  nand2 gate1187(.a(s_91), .b(gate118inter3), .O(gate118inter10));
  nor2  gate1188(.a(gate118inter10), .b(gate118inter9), .O(gate118inter11));
  nor2  gate1189(.a(gate118inter11), .b(gate118inter6), .O(gate118inter12));
  nand2 gate1190(.a(gate118inter12), .b(gate118inter1), .O(G465));

  xor2  gate1079(.a(G391), .b(G390), .O(gate119inter0));
  nand2 gate1080(.a(gate119inter0), .b(s_76), .O(gate119inter1));
  and2  gate1081(.a(G391), .b(G390), .O(gate119inter2));
  inv1  gate1082(.a(s_76), .O(gate119inter3));
  inv1  gate1083(.a(s_77), .O(gate119inter4));
  nand2 gate1084(.a(gate119inter4), .b(gate119inter3), .O(gate119inter5));
  nor2  gate1085(.a(gate119inter5), .b(gate119inter2), .O(gate119inter6));
  inv1  gate1086(.a(G390), .O(gate119inter7));
  inv1  gate1087(.a(G391), .O(gate119inter8));
  nand2 gate1088(.a(gate119inter8), .b(gate119inter7), .O(gate119inter9));
  nand2 gate1089(.a(s_77), .b(gate119inter3), .O(gate119inter10));
  nor2  gate1090(.a(gate119inter10), .b(gate119inter9), .O(gate119inter11));
  nor2  gate1091(.a(gate119inter11), .b(gate119inter6), .O(gate119inter12));
  nand2 gate1092(.a(gate119inter12), .b(gate119inter1), .O(G468));

  xor2  gate995(.a(G393), .b(G392), .O(gate120inter0));
  nand2 gate996(.a(gate120inter0), .b(s_64), .O(gate120inter1));
  and2  gate997(.a(G393), .b(G392), .O(gate120inter2));
  inv1  gate998(.a(s_64), .O(gate120inter3));
  inv1  gate999(.a(s_65), .O(gate120inter4));
  nand2 gate1000(.a(gate120inter4), .b(gate120inter3), .O(gate120inter5));
  nor2  gate1001(.a(gate120inter5), .b(gate120inter2), .O(gate120inter6));
  inv1  gate1002(.a(G392), .O(gate120inter7));
  inv1  gate1003(.a(G393), .O(gate120inter8));
  nand2 gate1004(.a(gate120inter8), .b(gate120inter7), .O(gate120inter9));
  nand2 gate1005(.a(s_65), .b(gate120inter3), .O(gate120inter10));
  nor2  gate1006(.a(gate120inter10), .b(gate120inter9), .O(gate120inter11));
  nor2  gate1007(.a(gate120inter11), .b(gate120inter6), .O(gate120inter12));
  nand2 gate1008(.a(gate120inter12), .b(gate120inter1), .O(G471));
nand2 gate121( .a(G394), .b(G395), .O(G474) );

  xor2  gate1219(.a(G397), .b(G396), .O(gate122inter0));
  nand2 gate1220(.a(gate122inter0), .b(s_96), .O(gate122inter1));
  and2  gate1221(.a(G397), .b(G396), .O(gate122inter2));
  inv1  gate1222(.a(s_96), .O(gate122inter3));
  inv1  gate1223(.a(s_97), .O(gate122inter4));
  nand2 gate1224(.a(gate122inter4), .b(gate122inter3), .O(gate122inter5));
  nor2  gate1225(.a(gate122inter5), .b(gate122inter2), .O(gate122inter6));
  inv1  gate1226(.a(G396), .O(gate122inter7));
  inv1  gate1227(.a(G397), .O(gate122inter8));
  nand2 gate1228(.a(gate122inter8), .b(gate122inter7), .O(gate122inter9));
  nand2 gate1229(.a(s_97), .b(gate122inter3), .O(gate122inter10));
  nor2  gate1230(.a(gate122inter10), .b(gate122inter9), .O(gate122inter11));
  nor2  gate1231(.a(gate122inter11), .b(gate122inter6), .O(gate122inter12));
  nand2 gate1232(.a(gate122inter12), .b(gate122inter1), .O(G477));
nand2 gate123( .a(G398), .b(G399), .O(G480) );

  xor2  gate1149(.a(G401), .b(G400), .O(gate124inter0));
  nand2 gate1150(.a(gate124inter0), .b(s_86), .O(gate124inter1));
  and2  gate1151(.a(G401), .b(G400), .O(gate124inter2));
  inv1  gate1152(.a(s_86), .O(gate124inter3));
  inv1  gate1153(.a(s_87), .O(gate124inter4));
  nand2 gate1154(.a(gate124inter4), .b(gate124inter3), .O(gate124inter5));
  nor2  gate1155(.a(gate124inter5), .b(gate124inter2), .O(gate124inter6));
  inv1  gate1156(.a(G400), .O(gate124inter7));
  inv1  gate1157(.a(G401), .O(gate124inter8));
  nand2 gate1158(.a(gate124inter8), .b(gate124inter7), .O(gate124inter9));
  nand2 gate1159(.a(s_87), .b(gate124inter3), .O(gate124inter10));
  nor2  gate1160(.a(gate124inter10), .b(gate124inter9), .O(gate124inter11));
  nor2  gate1161(.a(gate124inter11), .b(gate124inter6), .O(gate124inter12));
  nand2 gate1162(.a(gate124inter12), .b(gate124inter1), .O(G483));

  xor2  gate1625(.a(G403), .b(G402), .O(gate125inter0));
  nand2 gate1626(.a(gate125inter0), .b(s_154), .O(gate125inter1));
  and2  gate1627(.a(G403), .b(G402), .O(gate125inter2));
  inv1  gate1628(.a(s_154), .O(gate125inter3));
  inv1  gate1629(.a(s_155), .O(gate125inter4));
  nand2 gate1630(.a(gate125inter4), .b(gate125inter3), .O(gate125inter5));
  nor2  gate1631(.a(gate125inter5), .b(gate125inter2), .O(gate125inter6));
  inv1  gate1632(.a(G402), .O(gate125inter7));
  inv1  gate1633(.a(G403), .O(gate125inter8));
  nand2 gate1634(.a(gate125inter8), .b(gate125inter7), .O(gate125inter9));
  nand2 gate1635(.a(s_155), .b(gate125inter3), .O(gate125inter10));
  nor2  gate1636(.a(gate125inter10), .b(gate125inter9), .O(gate125inter11));
  nor2  gate1637(.a(gate125inter11), .b(gate125inter6), .O(gate125inter12));
  nand2 gate1638(.a(gate125inter12), .b(gate125inter1), .O(G486));
nand2 gate126( .a(G404), .b(G405), .O(G489) );
nand2 gate127( .a(G406), .b(G407), .O(G492) );
nand2 gate128( .a(G408), .b(G409), .O(G495) );

  xor2  gate1093(.a(G411), .b(G410), .O(gate129inter0));
  nand2 gate1094(.a(gate129inter0), .b(s_78), .O(gate129inter1));
  and2  gate1095(.a(G411), .b(G410), .O(gate129inter2));
  inv1  gate1096(.a(s_78), .O(gate129inter3));
  inv1  gate1097(.a(s_79), .O(gate129inter4));
  nand2 gate1098(.a(gate129inter4), .b(gate129inter3), .O(gate129inter5));
  nor2  gate1099(.a(gate129inter5), .b(gate129inter2), .O(gate129inter6));
  inv1  gate1100(.a(G410), .O(gate129inter7));
  inv1  gate1101(.a(G411), .O(gate129inter8));
  nand2 gate1102(.a(gate129inter8), .b(gate129inter7), .O(gate129inter9));
  nand2 gate1103(.a(s_79), .b(gate129inter3), .O(gate129inter10));
  nor2  gate1104(.a(gate129inter10), .b(gate129inter9), .O(gate129inter11));
  nor2  gate1105(.a(gate129inter11), .b(gate129inter6), .O(gate129inter12));
  nand2 gate1106(.a(gate129inter12), .b(gate129inter1), .O(G498));
nand2 gate130( .a(G412), .b(G413), .O(G501) );
nand2 gate131( .a(G414), .b(G415), .O(G504) );
nand2 gate132( .a(G416), .b(G417), .O(G507) );

  xor2  gate1233(.a(G419), .b(G418), .O(gate133inter0));
  nand2 gate1234(.a(gate133inter0), .b(s_98), .O(gate133inter1));
  and2  gate1235(.a(G419), .b(G418), .O(gate133inter2));
  inv1  gate1236(.a(s_98), .O(gate133inter3));
  inv1  gate1237(.a(s_99), .O(gate133inter4));
  nand2 gate1238(.a(gate133inter4), .b(gate133inter3), .O(gate133inter5));
  nor2  gate1239(.a(gate133inter5), .b(gate133inter2), .O(gate133inter6));
  inv1  gate1240(.a(G418), .O(gate133inter7));
  inv1  gate1241(.a(G419), .O(gate133inter8));
  nand2 gate1242(.a(gate133inter8), .b(gate133inter7), .O(gate133inter9));
  nand2 gate1243(.a(s_99), .b(gate133inter3), .O(gate133inter10));
  nor2  gate1244(.a(gate133inter10), .b(gate133inter9), .O(gate133inter11));
  nor2  gate1245(.a(gate133inter11), .b(gate133inter6), .O(gate133inter12));
  nand2 gate1246(.a(gate133inter12), .b(gate133inter1), .O(G510));
nand2 gate134( .a(G420), .b(G421), .O(G513) );
nand2 gate135( .a(G422), .b(G423), .O(G516) );
nand2 gate136( .a(G424), .b(G425), .O(G519) );
nand2 gate137( .a(G426), .b(G429), .O(G522) );

  xor2  gate2087(.a(G435), .b(G432), .O(gate138inter0));
  nand2 gate2088(.a(gate138inter0), .b(s_220), .O(gate138inter1));
  and2  gate2089(.a(G435), .b(G432), .O(gate138inter2));
  inv1  gate2090(.a(s_220), .O(gate138inter3));
  inv1  gate2091(.a(s_221), .O(gate138inter4));
  nand2 gate2092(.a(gate138inter4), .b(gate138inter3), .O(gate138inter5));
  nor2  gate2093(.a(gate138inter5), .b(gate138inter2), .O(gate138inter6));
  inv1  gate2094(.a(G432), .O(gate138inter7));
  inv1  gate2095(.a(G435), .O(gate138inter8));
  nand2 gate2096(.a(gate138inter8), .b(gate138inter7), .O(gate138inter9));
  nand2 gate2097(.a(s_221), .b(gate138inter3), .O(gate138inter10));
  nor2  gate2098(.a(gate138inter10), .b(gate138inter9), .O(gate138inter11));
  nor2  gate2099(.a(gate138inter11), .b(gate138inter6), .O(gate138inter12));
  nand2 gate2100(.a(gate138inter12), .b(gate138inter1), .O(G525));

  xor2  gate547(.a(G441), .b(G438), .O(gate139inter0));
  nand2 gate548(.a(gate139inter0), .b(s_0), .O(gate139inter1));
  and2  gate549(.a(G441), .b(G438), .O(gate139inter2));
  inv1  gate550(.a(s_0), .O(gate139inter3));
  inv1  gate551(.a(s_1), .O(gate139inter4));
  nand2 gate552(.a(gate139inter4), .b(gate139inter3), .O(gate139inter5));
  nor2  gate553(.a(gate139inter5), .b(gate139inter2), .O(gate139inter6));
  inv1  gate554(.a(G438), .O(gate139inter7));
  inv1  gate555(.a(G441), .O(gate139inter8));
  nand2 gate556(.a(gate139inter8), .b(gate139inter7), .O(gate139inter9));
  nand2 gate557(.a(s_1), .b(gate139inter3), .O(gate139inter10));
  nor2  gate558(.a(gate139inter10), .b(gate139inter9), .O(gate139inter11));
  nor2  gate559(.a(gate139inter11), .b(gate139inter6), .O(gate139inter12));
  nand2 gate560(.a(gate139inter12), .b(gate139inter1), .O(G528));

  xor2  gate1359(.a(G447), .b(G444), .O(gate140inter0));
  nand2 gate1360(.a(gate140inter0), .b(s_116), .O(gate140inter1));
  and2  gate1361(.a(G447), .b(G444), .O(gate140inter2));
  inv1  gate1362(.a(s_116), .O(gate140inter3));
  inv1  gate1363(.a(s_117), .O(gate140inter4));
  nand2 gate1364(.a(gate140inter4), .b(gate140inter3), .O(gate140inter5));
  nor2  gate1365(.a(gate140inter5), .b(gate140inter2), .O(gate140inter6));
  inv1  gate1366(.a(G444), .O(gate140inter7));
  inv1  gate1367(.a(G447), .O(gate140inter8));
  nand2 gate1368(.a(gate140inter8), .b(gate140inter7), .O(gate140inter9));
  nand2 gate1369(.a(s_117), .b(gate140inter3), .O(gate140inter10));
  nor2  gate1370(.a(gate140inter10), .b(gate140inter9), .O(gate140inter11));
  nor2  gate1371(.a(gate140inter11), .b(gate140inter6), .O(gate140inter12));
  nand2 gate1372(.a(gate140inter12), .b(gate140inter1), .O(G531));
nand2 gate141( .a(G450), .b(G453), .O(G534) );
nand2 gate142( .a(G456), .b(G459), .O(G537) );

  xor2  gate1303(.a(G465), .b(G462), .O(gate143inter0));
  nand2 gate1304(.a(gate143inter0), .b(s_108), .O(gate143inter1));
  and2  gate1305(.a(G465), .b(G462), .O(gate143inter2));
  inv1  gate1306(.a(s_108), .O(gate143inter3));
  inv1  gate1307(.a(s_109), .O(gate143inter4));
  nand2 gate1308(.a(gate143inter4), .b(gate143inter3), .O(gate143inter5));
  nor2  gate1309(.a(gate143inter5), .b(gate143inter2), .O(gate143inter6));
  inv1  gate1310(.a(G462), .O(gate143inter7));
  inv1  gate1311(.a(G465), .O(gate143inter8));
  nand2 gate1312(.a(gate143inter8), .b(gate143inter7), .O(gate143inter9));
  nand2 gate1313(.a(s_109), .b(gate143inter3), .O(gate143inter10));
  nor2  gate1314(.a(gate143inter10), .b(gate143inter9), .O(gate143inter11));
  nor2  gate1315(.a(gate143inter11), .b(gate143inter6), .O(gate143inter12));
  nand2 gate1316(.a(gate143inter12), .b(gate143inter1), .O(G540));
nand2 gate144( .a(G468), .b(G471), .O(G543) );

  xor2  gate673(.a(G477), .b(G474), .O(gate145inter0));
  nand2 gate674(.a(gate145inter0), .b(s_18), .O(gate145inter1));
  and2  gate675(.a(G477), .b(G474), .O(gate145inter2));
  inv1  gate676(.a(s_18), .O(gate145inter3));
  inv1  gate677(.a(s_19), .O(gate145inter4));
  nand2 gate678(.a(gate145inter4), .b(gate145inter3), .O(gate145inter5));
  nor2  gate679(.a(gate145inter5), .b(gate145inter2), .O(gate145inter6));
  inv1  gate680(.a(G474), .O(gate145inter7));
  inv1  gate681(.a(G477), .O(gate145inter8));
  nand2 gate682(.a(gate145inter8), .b(gate145inter7), .O(gate145inter9));
  nand2 gate683(.a(s_19), .b(gate145inter3), .O(gate145inter10));
  nor2  gate684(.a(gate145inter10), .b(gate145inter9), .O(gate145inter11));
  nor2  gate685(.a(gate145inter11), .b(gate145inter6), .O(gate145inter12));
  nand2 gate686(.a(gate145inter12), .b(gate145inter1), .O(G546));
nand2 gate146( .a(G480), .b(G483), .O(G549) );
nand2 gate147( .a(G486), .b(G489), .O(G552) );
nand2 gate148( .a(G492), .b(G495), .O(G555) );
nand2 gate149( .a(G498), .b(G501), .O(G558) );

  xor2  gate589(.a(G507), .b(G504), .O(gate150inter0));
  nand2 gate590(.a(gate150inter0), .b(s_6), .O(gate150inter1));
  and2  gate591(.a(G507), .b(G504), .O(gate150inter2));
  inv1  gate592(.a(s_6), .O(gate150inter3));
  inv1  gate593(.a(s_7), .O(gate150inter4));
  nand2 gate594(.a(gate150inter4), .b(gate150inter3), .O(gate150inter5));
  nor2  gate595(.a(gate150inter5), .b(gate150inter2), .O(gate150inter6));
  inv1  gate596(.a(G504), .O(gate150inter7));
  inv1  gate597(.a(G507), .O(gate150inter8));
  nand2 gate598(.a(gate150inter8), .b(gate150inter7), .O(gate150inter9));
  nand2 gate599(.a(s_7), .b(gate150inter3), .O(gate150inter10));
  nor2  gate600(.a(gate150inter10), .b(gate150inter9), .O(gate150inter11));
  nor2  gate601(.a(gate150inter11), .b(gate150inter6), .O(gate150inter12));
  nand2 gate602(.a(gate150inter12), .b(gate150inter1), .O(G561));
nand2 gate151( .a(G510), .b(G513), .O(G564) );
nand2 gate152( .a(G516), .b(G519), .O(G567) );
nand2 gate153( .a(G426), .b(G522), .O(G570) );
nand2 gate154( .a(G429), .b(G522), .O(G571) );
nand2 gate155( .a(G432), .b(G525), .O(G572) );
nand2 gate156( .a(G435), .b(G525), .O(G573) );
nand2 gate157( .a(G438), .b(G528), .O(G574) );
nand2 gate158( .a(G441), .b(G528), .O(G575) );
nand2 gate159( .a(G444), .b(G531), .O(G576) );
nand2 gate160( .a(G447), .b(G531), .O(G577) );
nand2 gate161( .a(G450), .b(G534), .O(G578) );
nand2 gate162( .a(G453), .b(G534), .O(G579) );
nand2 gate163( .a(G456), .b(G537), .O(G580) );
nand2 gate164( .a(G459), .b(G537), .O(G581) );
nand2 gate165( .a(G462), .b(G540), .O(G582) );
nand2 gate166( .a(G465), .b(G540), .O(G583) );
nand2 gate167( .a(G468), .b(G543), .O(G584) );
nand2 gate168( .a(G471), .b(G543), .O(G585) );
nand2 gate169( .a(G474), .b(G546), .O(G586) );

  xor2  gate743(.a(G546), .b(G477), .O(gate170inter0));
  nand2 gate744(.a(gate170inter0), .b(s_28), .O(gate170inter1));
  and2  gate745(.a(G546), .b(G477), .O(gate170inter2));
  inv1  gate746(.a(s_28), .O(gate170inter3));
  inv1  gate747(.a(s_29), .O(gate170inter4));
  nand2 gate748(.a(gate170inter4), .b(gate170inter3), .O(gate170inter5));
  nor2  gate749(.a(gate170inter5), .b(gate170inter2), .O(gate170inter6));
  inv1  gate750(.a(G477), .O(gate170inter7));
  inv1  gate751(.a(G546), .O(gate170inter8));
  nand2 gate752(.a(gate170inter8), .b(gate170inter7), .O(gate170inter9));
  nand2 gate753(.a(s_29), .b(gate170inter3), .O(gate170inter10));
  nor2  gate754(.a(gate170inter10), .b(gate170inter9), .O(gate170inter11));
  nor2  gate755(.a(gate170inter11), .b(gate170inter6), .O(gate170inter12));
  nand2 gate756(.a(gate170inter12), .b(gate170inter1), .O(G587));
nand2 gate171( .a(G480), .b(G549), .O(G588) );

  xor2  gate1653(.a(G549), .b(G483), .O(gate172inter0));
  nand2 gate1654(.a(gate172inter0), .b(s_158), .O(gate172inter1));
  and2  gate1655(.a(G549), .b(G483), .O(gate172inter2));
  inv1  gate1656(.a(s_158), .O(gate172inter3));
  inv1  gate1657(.a(s_159), .O(gate172inter4));
  nand2 gate1658(.a(gate172inter4), .b(gate172inter3), .O(gate172inter5));
  nor2  gate1659(.a(gate172inter5), .b(gate172inter2), .O(gate172inter6));
  inv1  gate1660(.a(G483), .O(gate172inter7));
  inv1  gate1661(.a(G549), .O(gate172inter8));
  nand2 gate1662(.a(gate172inter8), .b(gate172inter7), .O(gate172inter9));
  nand2 gate1663(.a(s_159), .b(gate172inter3), .O(gate172inter10));
  nor2  gate1664(.a(gate172inter10), .b(gate172inter9), .O(gate172inter11));
  nor2  gate1665(.a(gate172inter11), .b(gate172inter6), .O(gate172inter12));
  nand2 gate1666(.a(gate172inter12), .b(gate172inter1), .O(G589));
nand2 gate173( .a(G486), .b(G552), .O(G590) );

  xor2  gate827(.a(G552), .b(G489), .O(gate174inter0));
  nand2 gate828(.a(gate174inter0), .b(s_40), .O(gate174inter1));
  and2  gate829(.a(G552), .b(G489), .O(gate174inter2));
  inv1  gate830(.a(s_40), .O(gate174inter3));
  inv1  gate831(.a(s_41), .O(gate174inter4));
  nand2 gate832(.a(gate174inter4), .b(gate174inter3), .O(gate174inter5));
  nor2  gate833(.a(gate174inter5), .b(gate174inter2), .O(gate174inter6));
  inv1  gate834(.a(G489), .O(gate174inter7));
  inv1  gate835(.a(G552), .O(gate174inter8));
  nand2 gate836(.a(gate174inter8), .b(gate174inter7), .O(gate174inter9));
  nand2 gate837(.a(s_41), .b(gate174inter3), .O(gate174inter10));
  nor2  gate838(.a(gate174inter10), .b(gate174inter9), .O(gate174inter11));
  nor2  gate839(.a(gate174inter11), .b(gate174inter6), .O(gate174inter12));
  nand2 gate840(.a(gate174inter12), .b(gate174inter1), .O(G591));
nand2 gate175( .a(G492), .b(G555), .O(G592) );
nand2 gate176( .a(G495), .b(G555), .O(G593) );
nand2 gate177( .a(G498), .b(G558), .O(G594) );

  xor2  gate981(.a(G558), .b(G501), .O(gate178inter0));
  nand2 gate982(.a(gate178inter0), .b(s_62), .O(gate178inter1));
  and2  gate983(.a(G558), .b(G501), .O(gate178inter2));
  inv1  gate984(.a(s_62), .O(gate178inter3));
  inv1  gate985(.a(s_63), .O(gate178inter4));
  nand2 gate986(.a(gate178inter4), .b(gate178inter3), .O(gate178inter5));
  nor2  gate987(.a(gate178inter5), .b(gate178inter2), .O(gate178inter6));
  inv1  gate988(.a(G501), .O(gate178inter7));
  inv1  gate989(.a(G558), .O(gate178inter8));
  nand2 gate990(.a(gate178inter8), .b(gate178inter7), .O(gate178inter9));
  nand2 gate991(.a(s_63), .b(gate178inter3), .O(gate178inter10));
  nor2  gate992(.a(gate178inter10), .b(gate178inter9), .O(gate178inter11));
  nor2  gate993(.a(gate178inter11), .b(gate178inter6), .O(gate178inter12));
  nand2 gate994(.a(gate178inter12), .b(gate178inter1), .O(G595));
nand2 gate179( .a(G504), .b(G561), .O(G596) );
nand2 gate180( .a(G507), .b(G561), .O(G597) );
nand2 gate181( .a(G510), .b(G564), .O(G598) );
nand2 gate182( .a(G513), .b(G564), .O(G599) );

  xor2  gate631(.a(G567), .b(G516), .O(gate183inter0));
  nand2 gate632(.a(gate183inter0), .b(s_12), .O(gate183inter1));
  and2  gate633(.a(G567), .b(G516), .O(gate183inter2));
  inv1  gate634(.a(s_12), .O(gate183inter3));
  inv1  gate635(.a(s_13), .O(gate183inter4));
  nand2 gate636(.a(gate183inter4), .b(gate183inter3), .O(gate183inter5));
  nor2  gate637(.a(gate183inter5), .b(gate183inter2), .O(gate183inter6));
  inv1  gate638(.a(G516), .O(gate183inter7));
  inv1  gate639(.a(G567), .O(gate183inter8));
  nand2 gate640(.a(gate183inter8), .b(gate183inter7), .O(gate183inter9));
  nand2 gate641(.a(s_13), .b(gate183inter3), .O(gate183inter10));
  nor2  gate642(.a(gate183inter10), .b(gate183inter9), .O(gate183inter11));
  nor2  gate643(.a(gate183inter11), .b(gate183inter6), .O(gate183inter12));
  nand2 gate644(.a(gate183inter12), .b(gate183inter1), .O(G600));
nand2 gate184( .a(G519), .b(G567), .O(G601) );

  xor2  gate1051(.a(G571), .b(G570), .O(gate185inter0));
  nand2 gate1052(.a(gate185inter0), .b(s_72), .O(gate185inter1));
  and2  gate1053(.a(G571), .b(G570), .O(gate185inter2));
  inv1  gate1054(.a(s_72), .O(gate185inter3));
  inv1  gate1055(.a(s_73), .O(gate185inter4));
  nand2 gate1056(.a(gate185inter4), .b(gate185inter3), .O(gate185inter5));
  nor2  gate1057(.a(gate185inter5), .b(gate185inter2), .O(gate185inter6));
  inv1  gate1058(.a(G570), .O(gate185inter7));
  inv1  gate1059(.a(G571), .O(gate185inter8));
  nand2 gate1060(.a(gate185inter8), .b(gate185inter7), .O(gate185inter9));
  nand2 gate1061(.a(s_73), .b(gate185inter3), .O(gate185inter10));
  nor2  gate1062(.a(gate185inter10), .b(gate185inter9), .O(gate185inter11));
  nor2  gate1063(.a(gate185inter11), .b(gate185inter6), .O(gate185inter12));
  nand2 gate1064(.a(gate185inter12), .b(gate185inter1), .O(G602));

  xor2  gate799(.a(G573), .b(G572), .O(gate186inter0));
  nand2 gate800(.a(gate186inter0), .b(s_36), .O(gate186inter1));
  and2  gate801(.a(G573), .b(G572), .O(gate186inter2));
  inv1  gate802(.a(s_36), .O(gate186inter3));
  inv1  gate803(.a(s_37), .O(gate186inter4));
  nand2 gate804(.a(gate186inter4), .b(gate186inter3), .O(gate186inter5));
  nor2  gate805(.a(gate186inter5), .b(gate186inter2), .O(gate186inter6));
  inv1  gate806(.a(G572), .O(gate186inter7));
  inv1  gate807(.a(G573), .O(gate186inter8));
  nand2 gate808(.a(gate186inter8), .b(gate186inter7), .O(gate186inter9));
  nand2 gate809(.a(s_37), .b(gate186inter3), .O(gate186inter10));
  nor2  gate810(.a(gate186inter10), .b(gate186inter9), .O(gate186inter11));
  nor2  gate811(.a(gate186inter11), .b(gate186inter6), .O(gate186inter12));
  nand2 gate812(.a(gate186inter12), .b(gate186inter1), .O(G607));

  xor2  gate1863(.a(G575), .b(G574), .O(gate187inter0));
  nand2 gate1864(.a(gate187inter0), .b(s_188), .O(gate187inter1));
  and2  gate1865(.a(G575), .b(G574), .O(gate187inter2));
  inv1  gate1866(.a(s_188), .O(gate187inter3));
  inv1  gate1867(.a(s_189), .O(gate187inter4));
  nand2 gate1868(.a(gate187inter4), .b(gate187inter3), .O(gate187inter5));
  nor2  gate1869(.a(gate187inter5), .b(gate187inter2), .O(gate187inter6));
  inv1  gate1870(.a(G574), .O(gate187inter7));
  inv1  gate1871(.a(G575), .O(gate187inter8));
  nand2 gate1872(.a(gate187inter8), .b(gate187inter7), .O(gate187inter9));
  nand2 gate1873(.a(s_189), .b(gate187inter3), .O(gate187inter10));
  nor2  gate1874(.a(gate187inter10), .b(gate187inter9), .O(gate187inter11));
  nor2  gate1875(.a(gate187inter11), .b(gate187inter6), .O(gate187inter12));
  nand2 gate1876(.a(gate187inter12), .b(gate187inter1), .O(G612));
nand2 gate188( .a(G576), .b(G577), .O(G617) );
nand2 gate189( .a(G578), .b(G579), .O(G622) );

  xor2  gate1443(.a(G581), .b(G580), .O(gate190inter0));
  nand2 gate1444(.a(gate190inter0), .b(s_128), .O(gate190inter1));
  and2  gate1445(.a(G581), .b(G580), .O(gate190inter2));
  inv1  gate1446(.a(s_128), .O(gate190inter3));
  inv1  gate1447(.a(s_129), .O(gate190inter4));
  nand2 gate1448(.a(gate190inter4), .b(gate190inter3), .O(gate190inter5));
  nor2  gate1449(.a(gate190inter5), .b(gate190inter2), .O(gate190inter6));
  inv1  gate1450(.a(G580), .O(gate190inter7));
  inv1  gate1451(.a(G581), .O(gate190inter8));
  nand2 gate1452(.a(gate190inter8), .b(gate190inter7), .O(gate190inter9));
  nand2 gate1453(.a(s_129), .b(gate190inter3), .O(gate190inter10));
  nor2  gate1454(.a(gate190inter10), .b(gate190inter9), .O(gate190inter11));
  nor2  gate1455(.a(gate190inter11), .b(gate190inter6), .O(gate190inter12));
  nand2 gate1456(.a(gate190inter12), .b(gate190inter1), .O(G627));

  xor2  gate2059(.a(G583), .b(G582), .O(gate191inter0));
  nand2 gate2060(.a(gate191inter0), .b(s_216), .O(gate191inter1));
  and2  gate2061(.a(G583), .b(G582), .O(gate191inter2));
  inv1  gate2062(.a(s_216), .O(gate191inter3));
  inv1  gate2063(.a(s_217), .O(gate191inter4));
  nand2 gate2064(.a(gate191inter4), .b(gate191inter3), .O(gate191inter5));
  nor2  gate2065(.a(gate191inter5), .b(gate191inter2), .O(gate191inter6));
  inv1  gate2066(.a(G582), .O(gate191inter7));
  inv1  gate2067(.a(G583), .O(gate191inter8));
  nand2 gate2068(.a(gate191inter8), .b(gate191inter7), .O(gate191inter9));
  nand2 gate2069(.a(s_217), .b(gate191inter3), .O(gate191inter10));
  nor2  gate2070(.a(gate191inter10), .b(gate191inter9), .O(gate191inter11));
  nor2  gate2071(.a(gate191inter11), .b(gate191inter6), .O(gate191inter12));
  nand2 gate2072(.a(gate191inter12), .b(gate191inter1), .O(G632));
nand2 gate192( .a(G584), .b(G585), .O(G637) );

  xor2  gate1779(.a(G587), .b(G586), .O(gate193inter0));
  nand2 gate1780(.a(gate193inter0), .b(s_176), .O(gate193inter1));
  and2  gate1781(.a(G587), .b(G586), .O(gate193inter2));
  inv1  gate1782(.a(s_176), .O(gate193inter3));
  inv1  gate1783(.a(s_177), .O(gate193inter4));
  nand2 gate1784(.a(gate193inter4), .b(gate193inter3), .O(gate193inter5));
  nor2  gate1785(.a(gate193inter5), .b(gate193inter2), .O(gate193inter6));
  inv1  gate1786(.a(G586), .O(gate193inter7));
  inv1  gate1787(.a(G587), .O(gate193inter8));
  nand2 gate1788(.a(gate193inter8), .b(gate193inter7), .O(gate193inter9));
  nand2 gate1789(.a(s_177), .b(gate193inter3), .O(gate193inter10));
  nor2  gate1790(.a(gate193inter10), .b(gate193inter9), .O(gate193inter11));
  nor2  gate1791(.a(gate193inter11), .b(gate193inter6), .O(gate193inter12));
  nand2 gate1792(.a(gate193inter12), .b(gate193inter1), .O(G642));
nand2 gate194( .a(G588), .b(G589), .O(G645) );
nand2 gate195( .a(G590), .b(G591), .O(G648) );
nand2 gate196( .a(G592), .b(G593), .O(G651) );
nand2 gate197( .a(G594), .b(G595), .O(G654) );

  xor2  gate1961(.a(G597), .b(G596), .O(gate198inter0));
  nand2 gate1962(.a(gate198inter0), .b(s_202), .O(gate198inter1));
  and2  gate1963(.a(G597), .b(G596), .O(gate198inter2));
  inv1  gate1964(.a(s_202), .O(gate198inter3));
  inv1  gate1965(.a(s_203), .O(gate198inter4));
  nand2 gate1966(.a(gate198inter4), .b(gate198inter3), .O(gate198inter5));
  nor2  gate1967(.a(gate198inter5), .b(gate198inter2), .O(gate198inter6));
  inv1  gate1968(.a(G596), .O(gate198inter7));
  inv1  gate1969(.a(G597), .O(gate198inter8));
  nand2 gate1970(.a(gate198inter8), .b(gate198inter7), .O(gate198inter9));
  nand2 gate1971(.a(s_203), .b(gate198inter3), .O(gate198inter10));
  nor2  gate1972(.a(gate198inter10), .b(gate198inter9), .O(gate198inter11));
  nor2  gate1973(.a(gate198inter11), .b(gate198inter6), .O(gate198inter12));
  nand2 gate1974(.a(gate198inter12), .b(gate198inter1), .O(G657));
nand2 gate199( .a(G598), .b(G599), .O(G660) );
nand2 gate200( .a(G600), .b(G601), .O(G663) );
nand2 gate201( .a(G602), .b(G607), .O(G666) );
nand2 gate202( .a(G612), .b(G617), .O(G669) );

  xor2  gate1163(.a(G612), .b(G602), .O(gate203inter0));
  nand2 gate1164(.a(gate203inter0), .b(s_88), .O(gate203inter1));
  and2  gate1165(.a(G612), .b(G602), .O(gate203inter2));
  inv1  gate1166(.a(s_88), .O(gate203inter3));
  inv1  gate1167(.a(s_89), .O(gate203inter4));
  nand2 gate1168(.a(gate203inter4), .b(gate203inter3), .O(gate203inter5));
  nor2  gate1169(.a(gate203inter5), .b(gate203inter2), .O(gate203inter6));
  inv1  gate1170(.a(G602), .O(gate203inter7));
  inv1  gate1171(.a(G612), .O(gate203inter8));
  nand2 gate1172(.a(gate203inter8), .b(gate203inter7), .O(gate203inter9));
  nand2 gate1173(.a(s_89), .b(gate203inter3), .O(gate203inter10));
  nor2  gate1174(.a(gate203inter10), .b(gate203inter9), .O(gate203inter11));
  nor2  gate1175(.a(gate203inter11), .b(gate203inter6), .O(gate203inter12));
  nand2 gate1176(.a(gate203inter12), .b(gate203inter1), .O(G672));
nand2 gate204( .a(G607), .b(G617), .O(G675) );
nand2 gate205( .a(G622), .b(G627), .O(G678) );
nand2 gate206( .a(G632), .b(G637), .O(G681) );
nand2 gate207( .a(G622), .b(G632), .O(G684) );
nand2 gate208( .a(G627), .b(G637), .O(G687) );
nand2 gate209( .a(G602), .b(G666), .O(G690) );
nand2 gate210( .a(G607), .b(G666), .O(G691) );
nand2 gate211( .a(G612), .b(G669), .O(G692) );
nand2 gate212( .a(G617), .b(G669), .O(G693) );
nand2 gate213( .a(G602), .b(G672), .O(G694) );
nand2 gate214( .a(G612), .b(G672), .O(G695) );

  xor2  gate925(.a(G675), .b(G607), .O(gate215inter0));
  nand2 gate926(.a(gate215inter0), .b(s_54), .O(gate215inter1));
  and2  gate927(.a(G675), .b(G607), .O(gate215inter2));
  inv1  gate928(.a(s_54), .O(gate215inter3));
  inv1  gate929(.a(s_55), .O(gate215inter4));
  nand2 gate930(.a(gate215inter4), .b(gate215inter3), .O(gate215inter5));
  nor2  gate931(.a(gate215inter5), .b(gate215inter2), .O(gate215inter6));
  inv1  gate932(.a(G607), .O(gate215inter7));
  inv1  gate933(.a(G675), .O(gate215inter8));
  nand2 gate934(.a(gate215inter8), .b(gate215inter7), .O(gate215inter9));
  nand2 gate935(.a(s_55), .b(gate215inter3), .O(gate215inter10));
  nor2  gate936(.a(gate215inter10), .b(gate215inter9), .O(gate215inter11));
  nor2  gate937(.a(gate215inter11), .b(gate215inter6), .O(gate215inter12));
  nand2 gate938(.a(gate215inter12), .b(gate215inter1), .O(G696));
nand2 gate216( .a(G617), .b(G675), .O(G697) );
nand2 gate217( .a(G622), .b(G678), .O(G698) );
nand2 gate218( .a(G627), .b(G678), .O(G699) );
nand2 gate219( .a(G632), .b(G681), .O(G700) );

  xor2  gate1709(.a(G681), .b(G637), .O(gate220inter0));
  nand2 gate1710(.a(gate220inter0), .b(s_166), .O(gate220inter1));
  and2  gate1711(.a(G681), .b(G637), .O(gate220inter2));
  inv1  gate1712(.a(s_166), .O(gate220inter3));
  inv1  gate1713(.a(s_167), .O(gate220inter4));
  nand2 gate1714(.a(gate220inter4), .b(gate220inter3), .O(gate220inter5));
  nor2  gate1715(.a(gate220inter5), .b(gate220inter2), .O(gate220inter6));
  inv1  gate1716(.a(G637), .O(gate220inter7));
  inv1  gate1717(.a(G681), .O(gate220inter8));
  nand2 gate1718(.a(gate220inter8), .b(gate220inter7), .O(gate220inter9));
  nand2 gate1719(.a(s_167), .b(gate220inter3), .O(gate220inter10));
  nor2  gate1720(.a(gate220inter10), .b(gate220inter9), .O(gate220inter11));
  nor2  gate1721(.a(gate220inter11), .b(gate220inter6), .O(gate220inter12));
  nand2 gate1722(.a(gate220inter12), .b(gate220inter1), .O(G701));
nand2 gate221( .a(G622), .b(G684), .O(G702) );
nand2 gate222( .a(G632), .b(G684), .O(G703) );

  xor2  gate1891(.a(G687), .b(G627), .O(gate223inter0));
  nand2 gate1892(.a(gate223inter0), .b(s_192), .O(gate223inter1));
  and2  gate1893(.a(G687), .b(G627), .O(gate223inter2));
  inv1  gate1894(.a(s_192), .O(gate223inter3));
  inv1  gate1895(.a(s_193), .O(gate223inter4));
  nand2 gate1896(.a(gate223inter4), .b(gate223inter3), .O(gate223inter5));
  nor2  gate1897(.a(gate223inter5), .b(gate223inter2), .O(gate223inter6));
  inv1  gate1898(.a(G627), .O(gate223inter7));
  inv1  gate1899(.a(G687), .O(gate223inter8));
  nand2 gate1900(.a(gate223inter8), .b(gate223inter7), .O(gate223inter9));
  nand2 gate1901(.a(s_193), .b(gate223inter3), .O(gate223inter10));
  nor2  gate1902(.a(gate223inter10), .b(gate223inter9), .O(gate223inter11));
  nor2  gate1903(.a(gate223inter11), .b(gate223inter6), .O(gate223inter12));
  nand2 gate1904(.a(gate223inter12), .b(gate223inter1), .O(G704));

  xor2  gate617(.a(G687), .b(G637), .O(gate224inter0));
  nand2 gate618(.a(gate224inter0), .b(s_10), .O(gate224inter1));
  and2  gate619(.a(G687), .b(G637), .O(gate224inter2));
  inv1  gate620(.a(s_10), .O(gate224inter3));
  inv1  gate621(.a(s_11), .O(gate224inter4));
  nand2 gate622(.a(gate224inter4), .b(gate224inter3), .O(gate224inter5));
  nor2  gate623(.a(gate224inter5), .b(gate224inter2), .O(gate224inter6));
  inv1  gate624(.a(G637), .O(gate224inter7));
  inv1  gate625(.a(G687), .O(gate224inter8));
  nand2 gate626(.a(gate224inter8), .b(gate224inter7), .O(gate224inter9));
  nand2 gate627(.a(s_11), .b(gate224inter3), .O(gate224inter10));
  nor2  gate628(.a(gate224inter10), .b(gate224inter9), .O(gate224inter11));
  nor2  gate629(.a(gate224inter11), .b(gate224inter6), .O(gate224inter12));
  nand2 gate630(.a(gate224inter12), .b(gate224inter1), .O(G705));
nand2 gate225( .a(G690), .b(G691), .O(G706) );

  xor2  gate645(.a(G693), .b(G692), .O(gate226inter0));
  nand2 gate646(.a(gate226inter0), .b(s_14), .O(gate226inter1));
  and2  gate647(.a(G693), .b(G692), .O(gate226inter2));
  inv1  gate648(.a(s_14), .O(gate226inter3));
  inv1  gate649(.a(s_15), .O(gate226inter4));
  nand2 gate650(.a(gate226inter4), .b(gate226inter3), .O(gate226inter5));
  nor2  gate651(.a(gate226inter5), .b(gate226inter2), .O(gate226inter6));
  inv1  gate652(.a(G692), .O(gate226inter7));
  inv1  gate653(.a(G693), .O(gate226inter8));
  nand2 gate654(.a(gate226inter8), .b(gate226inter7), .O(gate226inter9));
  nand2 gate655(.a(s_15), .b(gate226inter3), .O(gate226inter10));
  nor2  gate656(.a(gate226inter10), .b(gate226inter9), .O(gate226inter11));
  nor2  gate657(.a(gate226inter11), .b(gate226inter6), .O(gate226inter12));
  nand2 gate658(.a(gate226inter12), .b(gate226inter1), .O(G709));
nand2 gate227( .a(G694), .b(G695), .O(G712) );
nand2 gate228( .a(G696), .b(G697), .O(G715) );
nand2 gate229( .a(G698), .b(G699), .O(G718) );
nand2 gate230( .a(G700), .b(G701), .O(G721) );
nand2 gate231( .a(G702), .b(G703), .O(G724) );
nand2 gate232( .a(G704), .b(G705), .O(G727) );
nand2 gate233( .a(G242), .b(G718), .O(G730) );
nand2 gate234( .a(G245), .b(G721), .O(G733) );
nand2 gate235( .a(G248), .b(G724), .O(G736) );

  xor2  gate1793(.a(G727), .b(G251), .O(gate236inter0));
  nand2 gate1794(.a(gate236inter0), .b(s_178), .O(gate236inter1));
  and2  gate1795(.a(G727), .b(G251), .O(gate236inter2));
  inv1  gate1796(.a(s_178), .O(gate236inter3));
  inv1  gate1797(.a(s_179), .O(gate236inter4));
  nand2 gate1798(.a(gate236inter4), .b(gate236inter3), .O(gate236inter5));
  nor2  gate1799(.a(gate236inter5), .b(gate236inter2), .O(gate236inter6));
  inv1  gate1800(.a(G251), .O(gate236inter7));
  inv1  gate1801(.a(G727), .O(gate236inter8));
  nand2 gate1802(.a(gate236inter8), .b(gate236inter7), .O(gate236inter9));
  nand2 gate1803(.a(s_179), .b(gate236inter3), .O(gate236inter10));
  nor2  gate1804(.a(gate236inter10), .b(gate236inter9), .O(gate236inter11));
  nor2  gate1805(.a(gate236inter11), .b(gate236inter6), .O(gate236inter12));
  nand2 gate1806(.a(gate236inter12), .b(gate236inter1), .O(G739));
nand2 gate237( .a(G254), .b(G706), .O(G742) );
nand2 gate238( .a(G257), .b(G709), .O(G745) );

  xor2  gate1849(.a(G712), .b(G260), .O(gate239inter0));
  nand2 gate1850(.a(gate239inter0), .b(s_186), .O(gate239inter1));
  and2  gate1851(.a(G712), .b(G260), .O(gate239inter2));
  inv1  gate1852(.a(s_186), .O(gate239inter3));
  inv1  gate1853(.a(s_187), .O(gate239inter4));
  nand2 gate1854(.a(gate239inter4), .b(gate239inter3), .O(gate239inter5));
  nor2  gate1855(.a(gate239inter5), .b(gate239inter2), .O(gate239inter6));
  inv1  gate1856(.a(G260), .O(gate239inter7));
  inv1  gate1857(.a(G712), .O(gate239inter8));
  nand2 gate1858(.a(gate239inter8), .b(gate239inter7), .O(gate239inter9));
  nand2 gate1859(.a(s_187), .b(gate239inter3), .O(gate239inter10));
  nor2  gate1860(.a(gate239inter10), .b(gate239inter9), .O(gate239inter11));
  nor2  gate1861(.a(gate239inter11), .b(gate239inter6), .O(gate239inter12));
  nand2 gate1862(.a(gate239inter12), .b(gate239inter1), .O(G748));
nand2 gate240( .a(G263), .b(G715), .O(G751) );
nand2 gate241( .a(G242), .b(G730), .O(G754) );
nand2 gate242( .a(G718), .b(G730), .O(G755) );
nand2 gate243( .a(G245), .b(G733), .O(G756) );
nand2 gate244( .a(G721), .b(G733), .O(G757) );

  xor2  gate953(.a(G736), .b(G248), .O(gate245inter0));
  nand2 gate954(.a(gate245inter0), .b(s_58), .O(gate245inter1));
  and2  gate955(.a(G736), .b(G248), .O(gate245inter2));
  inv1  gate956(.a(s_58), .O(gate245inter3));
  inv1  gate957(.a(s_59), .O(gate245inter4));
  nand2 gate958(.a(gate245inter4), .b(gate245inter3), .O(gate245inter5));
  nor2  gate959(.a(gate245inter5), .b(gate245inter2), .O(gate245inter6));
  inv1  gate960(.a(G248), .O(gate245inter7));
  inv1  gate961(.a(G736), .O(gate245inter8));
  nand2 gate962(.a(gate245inter8), .b(gate245inter7), .O(gate245inter9));
  nand2 gate963(.a(s_59), .b(gate245inter3), .O(gate245inter10));
  nor2  gate964(.a(gate245inter10), .b(gate245inter9), .O(gate245inter11));
  nor2  gate965(.a(gate245inter11), .b(gate245inter6), .O(gate245inter12));
  nand2 gate966(.a(gate245inter12), .b(gate245inter1), .O(G758));
nand2 gate246( .a(G724), .b(G736), .O(G759) );
nand2 gate247( .a(G251), .b(G739), .O(G760) );
nand2 gate248( .a(G727), .b(G739), .O(G761) );
nand2 gate249( .a(G254), .b(G742), .O(G762) );

  xor2  gate1975(.a(G742), .b(G706), .O(gate250inter0));
  nand2 gate1976(.a(gate250inter0), .b(s_204), .O(gate250inter1));
  and2  gate1977(.a(G742), .b(G706), .O(gate250inter2));
  inv1  gate1978(.a(s_204), .O(gate250inter3));
  inv1  gate1979(.a(s_205), .O(gate250inter4));
  nand2 gate1980(.a(gate250inter4), .b(gate250inter3), .O(gate250inter5));
  nor2  gate1981(.a(gate250inter5), .b(gate250inter2), .O(gate250inter6));
  inv1  gate1982(.a(G706), .O(gate250inter7));
  inv1  gate1983(.a(G742), .O(gate250inter8));
  nand2 gate1984(.a(gate250inter8), .b(gate250inter7), .O(gate250inter9));
  nand2 gate1985(.a(s_205), .b(gate250inter3), .O(gate250inter10));
  nor2  gate1986(.a(gate250inter10), .b(gate250inter9), .O(gate250inter11));
  nor2  gate1987(.a(gate250inter11), .b(gate250inter6), .O(gate250inter12));
  nand2 gate1988(.a(gate250inter12), .b(gate250inter1), .O(G763));
nand2 gate251( .a(G257), .b(G745), .O(G764) );

  xor2  gate1499(.a(G745), .b(G709), .O(gate252inter0));
  nand2 gate1500(.a(gate252inter0), .b(s_136), .O(gate252inter1));
  and2  gate1501(.a(G745), .b(G709), .O(gate252inter2));
  inv1  gate1502(.a(s_136), .O(gate252inter3));
  inv1  gate1503(.a(s_137), .O(gate252inter4));
  nand2 gate1504(.a(gate252inter4), .b(gate252inter3), .O(gate252inter5));
  nor2  gate1505(.a(gate252inter5), .b(gate252inter2), .O(gate252inter6));
  inv1  gate1506(.a(G709), .O(gate252inter7));
  inv1  gate1507(.a(G745), .O(gate252inter8));
  nand2 gate1508(.a(gate252inter8), .b(gate252inter7), .O(gate252inter9));
  nand2 gate1509(.a(s_137), .b(gate252inter3), .O(gate252inter10));
  nor2  gate1510(.a(gate252inter10), .b(gate252inter9), .O(gate252inter11));
  nor2  gate1511(.a(gate252inter11), .b(gate252inter6), .O(gate252inter12));
  nand2 gate1512(.a(gate252inter12), .b(gate252inter1), .O(G765));
nand2 gate253( .a(G260), .b(G748), .O(G766) );
nand2 gate254( .a(G712), .b(G748), .O(G767) );
nand2 gate255( .a(G263), .b(G751), .O(G768) );
nand2 gate256( .a(G715), .b(G751), .O(G769) );
nand2 gate257( .a(G754), .b(G755), .O(G770) );
nand2 gate258( .a(G756), .b(G757), .O(G773) );
nand2 gate259( .a(G758), .b(G759), .O(G776) );
nand2 gate260( .a(G760), .b(G761), .O(G779) );

  xor2  gate2045(.a(G763), .b(G762), .O(gate261inter0));
  nand2 gate2046(.a(gate261inter0), .b(s_214), .O(gate261inter1));
  and2  gate2047(.a(G763), .b(G762), .O(gate261inter2));
  inv1  gate2048(.a(s_214), .O(gate261inter3));
  inv1  gate2049(.a(s_215), .O(gate261inter4));
  nand2 gate2050(.a(gate261inter4), .b(gate261inter3), .O(gate261inter5));
  nor2  gate2051(.a(gate261inter5), .b(gate261inter2), .O(gate261inter6));
  inv1  gate2052(.a(G762), .O(gate261inter7));
  inv1  gate2053(.a(G763), .O(gate261inter8));
  nand2 gate2054(.a(gate261inter8), .b(gate261inter7), .O(gate261inter9));
  nand2 gate2055(.a(s_215), .b(gate261inter3), .O(gate261inter10));
  nor2  gate2056(.a(gate261inter10), .b(gate261inter9), .O(gate261inter11));
  nor2  gate2057(.a(gate261inter11), .b(gate261inter6), .O(gate261inter12));
  nand2 gate2058(.a(gate261inter12), .b(gate261inter1), .O(G782));
nand2 gate262( .a(G764), .b(G765), .O(G785) );
nand2 gate263( .a(G766), .b(G767), .O(G788) );
nand2 gate264( .a(G768), .b(G769), .O(G791) );
nand2 gate265( .a(G642), .b(G770), .O(G794) );
nand2 gate266( .a(G645), .b(G773), .O(G797) );
nand2 gate267( .a(G648), .b(G776), .O(G800) );
nand2 gate268( .a(G651), .b(G779), .O(G803) );
nand2 gate269( .a(G654), .b(G782), .O(G806) );
nand2 gate270( .a(G657), .b(G785), .O(G809) );
nand2 gate271( .a(G660), .b(G788), .O(G812) );
nand2 gate272( .a(G663), .b(G791), .O(G815) );
nand2 gate273( .a(G642), .b(G794), .O(G818) );
nand2 gate274( .a(G770), .b(G794), .O(G819) );

  xor2  gate1065(.a(G797), .b(G645), .O(gate275inter0));
  nand2 gate1066(.a(gate275inter0), .b(s_74), .O(gate275inter1));
  and2  gate1067(.a(G797), .b(G645), .O(gate275inter2));
  inv1  gate1068(.a(s_74), .O(gate275inter3));
  inv1  gate1069(.a(s_75), .O(gate275inter4));
  nand2 gate1070(.a(gate275inter4), .b(gate275inter3), .O(gate275inter5));
  nor2  gate1071(.a(gate275inter5), .b(gate275inter2), .O(gate275inter6));
  inv1  gate1072(.a(G645), .O(gate275inter7));
  inv1  gate1073(.a(G797), .O(gate275inter8));
  nand2 gate1074(.a(gate275inter8), .b(gate275inter7), .O(gate275inter9));
  nand2 gate1075(.a(s_75), .b(gate275inter3), .O(gate275inter10));
  nor2  gate1076(.a(gate275inter10), .b(gate275inter9), .O(gate275inter11));
  nor2  gate1077(.a(gate275inter11), .b(gate275inter6), .O(gate275inter12));
  nand2 gate1078(.a(gate275inter12), .b(gate275inter1), .O(G820));
nand2 gate276( .a(G773), .b(G797), .O(G821) );

  xor2  gate575(.a(G800), .b(G648), .O(gate277inter0));
  nand2 gate576(.a(gate277inter0), .b(s_4), .O(gate277inter1));
  and2  gate577(.a(G800), .b(G648), .O(gate277inter2));
  inv1  gate578(.a(s_4), .O(gate277inter3));
  inv1  gate579(.a(s_5), .O(gate277inter4));
  nand2 gate580(.a(gate277inter4), .b(gate277inter3), .O(gate277inter5));
  nor2  gate581(.a(gate277inter5), .b(gate277inter2), .O(gate277inter6));
  inv1  gate582(.a(G648), .O(gate277inter7));
  inv1  gate583(.a(G800), .O(gate277inter8));
  nand2 gate584(.a(gate277inter8), .b(gate277inter7), .O(gate277inter9));
  nand2 gate585(.a(s_5), .b(gate277inter3), .O(gate277inter10));
  nor2  gate586(.a(gate277inter10), .b(gate277inter9), .O(gate277inter11));
  nor2  gate587(.a(gate277inter11), .b(gate277inter6), .O(gate277inter12));
  nand2 gate588(.a(gate277inter12), .b(gate277inter1), .O(G822));

  xor2  gate1485(.a(G800), .b(G776), .O(gate278inter0));
  nand2 gate1486(.a(gate278inter0), .b(s_134), .O(gate278inter1));
  and2  gate1487(.a(G800), .b(G776), .O(gate278inter2));
  inv1  gate1488(.a(s_134), .O(gate278inter3));
  inv1  gate1489(.a(s_135), .O(gate278inter4));
  nand2 gate1490(.a(gate278inter4), .b(gate278inter3), .O(gate278inter5));
  nor2  gate1491(.a(gate278inter5), .b(gate278inter2), .O(gate278inter6));
  inv1  gate1492(.a(G776), .O(gate278inter7));
  inv1  gate1493(.a(G800), .O(gate278inter8));
  nand2 gate1494(.a(gate278inter8), .b(gate278inter7), .O(gate278inter9));
  nand2 gate1495(.a(s_135), .b(gate278inter3), .O(gate278inter10));
  nor2  gate1496(.a(gate278inter10), .b(gate278inter9), .O(gate278inter11));
  nor2  gate1497(.a(gate278inter11), .b(gate278inter6), .O(gate278inter12));
  nand2 gate1498(.a(gate278inter12), .b(gate278inter1), .O(G823));
nand2 gate279( .a(G651), .b(G803), .O(G824) );
nand2 gate280( .a(G779), .b(G803), .O(G825) );
nand2 gate281( .a(G654), .b(G806), .O(G826) );
nand2 gate282( .a(G782), .b(G806), .O(G827) );
nand2 gate283( .a(G657), .b(G809), .O(G828) );
nand2 gate284( .a(G785), .b(G809), .O(G829) );
nand2 gate285( .a(G660), .b(G812), .O(G830) );
nand2 gate286( .a(G788), .b(G812), .O(G831) );

  xor2  gate1541(.a(G815), .b(G663), .O(gate287inter0));
  nand2 gate1542(.a(gate287inter0), .b(s_142), .O(gate287inter1));
  and2  gate1543(.a(G815), .b(G663), .O(gate287inter2));
  inv1  gate1544(.a(s_142), .O(gate287inter3));
  inv1  gate1545(.a(s_143), .O(gate287inter4));
  nand2 gate1546(.a(gate287inter4), .b(gate287inter3), .O(gate287inter5));
  nor2  gate1547(.a(gate287inter5), .b(gate287inter2), .O(gate287inter6));
  inv1  gate1548(.a(G663), .O(gate287inter7));
  inv1  gate1549(.a(G815), .O(gate287inter8));
  nand2 gate1550(.a(gate287inter8), .b(gate287inter7), .O(gate287inter9));
  nand2 gate1551(.a(s_143), .b(gate287inter3), .O(gate287inter10));
  nor2  gate1552(.a(gate287inter10), .b(gate287inter9), .O(gate287inter11));
  nor2  gate1553(.a(gate287inter11), .b(gate287inter6), .O(gate287inter12));
  nand2 gate1554(.a(gate287inter12), .b(gate287inter1), .O(G832));
nand2 gate288( .a(G791), .b(G815), .O(G833) );
nand2 gate289( .a(G818), .b(G819), .O(G834) );
nand2 gate290( .a(G820), .b(G821), .O(G847) );

  xor2  gate2031(.a(G823), .b(G822), .O(gate291inter0));
  nand2 gate2032(.a(gate291inter0), .b(s_212), .O(gate291inter1));
  and2  gate2033(.a(G823), .b(G822), .O(gate291inter2));
  inv1  gate2034(.a(s_212), .O(gate291inter3));
  inv1  gate2035(.a(s_213), .O(gate291inter4));
  nand2 gate2036(.a(gate291inter4), .b(gate291inter3), .O(gate291inter5));
  nor2  gate2037(.a(gate291inter5), .b(gate291inter2), .O(gate291inter6));
  inv1  gate2038(.a(G822), .O(gate291inter7));
  inv1  gate2039(.a(G823), .O(gate291inter8));
  nand2 gate2040(.a(gate291inter8), .b(gate291inter7), .O(gate291inter9));
  nand2 gate2041(.a(s_213), .b(gate291inter3), .O(gate291inter10));
  nor2  gate2042(.a(gate291inter10), .b(gate291inter9), .O(gate291inter11));
  nor2  gate2043(.a(gate291inter11), .b(gate291inter6), .O(gate291inter12));
  nand2 gate2044(.a(gate291inter12), .b(gate291inter1), .O(G860));
nand2 gate292( .a(G824), .b(G825), .O(G873) );

  xor2  gate1261(.a(G829), .b(G828), .O(gate293inter0));
  nand2 gate1262(.a(gate293inter0), .b(s_102), .O(gate293inter1));
  and2  gate1263(.a(G829), .b(G828), .O(gate293inter2));
  inv1  gate1264(.a(s_102), .O(gate293inter3));
  inv1  gate1265(.a(s_103), .O(gate293inter4));
  nand2 gate1266(.a(gate293inter4), .b(gate293inter3), .O(gate293inter5));
  nor2  gate1267(.a(gate293inter5), .b(gate293inter2), .O(gate293inter6));
  inv1  gate1268(.a(G828), .O(gate293inter7));
  inv1  gate1269(.a(G829), .O(gate293inter8));
  nand2 gate1270(.a(gate293inter8), .b(gate293inter7), .O(gate293inter9));
  nand2 gate1271(.a(s_103), .b(gate293inter3), .O(gate293inter10));
  nor2  gate1272(.a(gate293inter10), .b(gate293inter9), .O(gate293inter11));
  nor2  gate1273(.a(gate293inter11), .b(gate293inter6), .O(gate293inter12));
  nand2 gate1274(.a(gate293inter12), .b(gate293inter1), .O(G886));

  xor2  gate1107(.a(G833), .b(G832), .O(gate294inter0));
  nand2 gate1108(.a(gate294inter0), .b(s_80), .O(gate294inter1));
  and2  gate1109(.a(G833), .b(G832), .O(gate294inter2));
  inv1  gate1110(.a(s_80), .O(gate294inter3));
  inv1  gate1111(.a(s_81), .O(gate294inter4));
  nand2 gate1112(.a(gate294inter4), .b(gate294inter3), .O(gate294inter5));
  nor2  gate1113(.a(gate294inter5), .b(gate294inter2), .O(gate294inter6));
  inv1  gate1114(.a(G832), .O(gate294inter7));
  inv1  gate1115(.a(G833), .O(gate294inter8));
  nand2 gate1116(.a(gate294inter8), .b(gate294inter7), .O(gate294inter9));
  nand2 gate1117(.a(s_81), .b(gate294inter3), .O(gate294inter10));
  nor2  gate1118(.a(gate294inter10), .b(gate294inter9), .O(gate294inter11));
  nor2  gate1119(.a(gate294inter11), .b(gate294inter6), .O(gate294inter12));
  nand2 gate1120(.a(gate294inter12), .b(gate294inter1), .O(G899));
nand2 gate295( .a(G830), .b(G831), .O(G912) );
nand2 gate296( .a(G826), .b(G827), .O(G925) );
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );

  xor2  gate869(.a(G1036), .b(G1), .O(gate387inter0));
  nand2 gate870(.a(gate387inter0), .b(s_46), .O(gate387inter1));
  and2  gate871(.a(G1036), .b(G1), .O(gate387inter2));
  inv1  gate872(.a(s_46), .O(gate387inter3));
  inv1  gate873(.a(s_47), .O(gate387inter4));
  nand2 gate874(.a(gate387inter4), .b(gate387inter3), .O(gate387inter5));
  nor2  gate875(.a(gate387inter5), .b(gate387inter2), .O(gate387inter6));
  inv1  gate876(.a(G1), .O(gate387inter7));
  inv1  gate877(.a(G1036), .O(gate387inter8));
  nand2 gate878(.a(gate387inter8), .b(gate387inter7), .O(gate387inter9));
  nand2 gate879(.a(s_47), .b(gate387inter3), .O(gate387inter10));
  nor2  gate880(.a(gate387inter10), .b(gate387inter9), .O(gate387inter11));
  nor2  gate881(.a(gate387inter11), .b(gate387inter6), .O(gate387inter12));
  nand2 gate882(.a(gate387inter12), .b(gate387inter1), .O(G1132));

  xor2  gate1023(.a(G1039), .b(G2), .O(gate388inter0));
  nand2 gate1024(.a(gate388inter0), .b(s_68), .O(gate388inter1));
  and2  gate1025(.a(G1039), .b(G2), .O(gate388inter2));
  inv1  gate1026(.a(s_68), .O(gate388inter3));
  inv1  gate1027(.a(s_69), .O(gate388inter4));
  nand2 gate1028(.a(gate388inter4), .b(gate388inter3), .O(gate388inter5));
  nor2  gate1029(.a(gate388inter5), .b(gate388inter2), .O(gate388inter6));
  inv1  gate1030(.a(G2), .O(gate388inter7));
  inv1  gate1031(.a(G1039), .O(gate388inter8));
  nand2 gate1032(.a(gate388inter8), .b(gate388inter7), .O(gate388inter9));
  nand2 gate1033(.a(s_69), .b(gate388inter3), .O(gate388inter10));
  nor2  gate1034(.a(gate388inter10), .b(gate388inter9), .O(gate388inter11));
  nor2  gate1035(.a(gate388inter11), .b(gate388inter6), .O(gate388inter12));
  nand2 gate1036(.a(gate388inter12), .b(gate388inter1), .O(G1135));
nand2 gate389( .a(G3), .b(G1042), .O(G1138) );
nand2 gate390( .a(G4), .b(G1045), .O(G1141) );
nand2 gate391( .a(G5), .b(G1048), .O(G1144) );
nand2 gate392( .a(G6), .b(G1051), .O(G1147) );
nand2 gate393( .a(G7), .b(G1054), .O(G1150) );
nand2 gate394( .a(G8), .b(G1057), .O(G1153) );

  xor2  gate603(.a(G1060), .b(G9), .O(gate395inter0));
  nand2 gate604(.a(gate395inter0), .b(s_8), .O(gate395inter1));
  and2  gate605(.a(G1060), .b(G9), .O(gate395inter2));
  inv1  gate606(.a(s_8), .O(gate395inter3));
  inv1  gate607(.a(s_9), .O(gate395inter4));
  nand2 gate608(.a(gate395inter4), .b(gate395inter3), .O(gate395inter5));
  nor2  gate609(.a(gate395inter5), .b(gate395inter2), .O(gate395inter6));
  inv1  gate610(.a(G9), .O(gate395inter7));
  inv1  gate611(.a(G1060), .O(gate395inter8));
  nand2 gate612(.a(gate395inter8), .b(gate395inter7), .O(gate395inter9));
  nand2 gate613(.a(s_9), .b(gate395inter3), .O(gate395inter10));
  nor2  gate614(.a(gate395inter10), .b(gate395inter9), .O(gate395inter11));
  nor2  gate615(.a(gate395inter11), .b(gate395inter6), .O(gate395inter12));
  nand2 gate616(.a(gate395inter12), .b(gate395inter1), .O(G1156));
nand2 gate396( .a(G10), .b(G1063), .O(G1159) );

  xor2  gate1135(.a(G1066), .b(G11), .O(gate397inter0));
  nand2 gate1136(.a(gate397inter0), .b(s_84), .O(gate397inter1));
  and2  gate1137(.a(G1066), .b(G11), .O(gate397inter2));
  inv1  gate1138(.a(s_84), .O(gate397inter3));
  inv1  gate1139(.a(s_85), .O(gate397inter4));
  nand2 gate1140(.a(gate397inter4), .b(gate397inter3), .O(gate397inter5));
  nor2  gate1141(.a(gate397inter5), .b(gate397inter2), .O(gate397inter6));
  inv1  gate1142(.a(G11), .O(gate397inter7));
  inv1  gate1143(.a(G1066), .O(gate397inter8));
  nand2 gate1144(.a(gate397inter8), .b(gate397inter7), .O(gate397inter9));
  nand2 gate1145(.a(s_85), .b(gate397inter3), .O(gate397inter10));
  nor2  gate1146(.a(gate397inter10), .b(gate397inter9), .O(gate397inter11));
  nor2  gate1147(.a(gate397inter11), .b(gate397inter6), .O(gate397inter12));
  nand2 gate1148(.a(gate397inter12), .b(gate397inter1), .O(G1162));
nand2 gate398( .a(G12), .b(G1069), .O(G1165) );
nand2 gate399( .a(G13), .b(G1072), .O(G1168) );
nand2 gate400( .a(G14), .b(G1075), .O(G1171) );
nand2 gate401( .a(G15), .b(G1078), .O(G1174) );

  xor2  gate1681(.a(G1081), .b(G16), .O(gate402inter0));
  nand2 gate1682(.a(gate402inter0), .b(s_162), .O(gate402inter1));
  and2  gate1683(.a(G1081), .b(G16), .O(gate402inter2));
  inv1  gate1684(.a(s_162), .O(gate402inter3));
  inv1  gate1685(.a(s_163), .O(gate402inter4));
  nand2 gate1686(.a(gate402inter4), .b(gate402inter3), .O(gate402inter5));
  nor2  gate1687(.a(gate402inter5), .b(gate402inter2), .O(gate402inter6));
  inv1  gate1688(.a(G16), .O(gate402inter7));
  inv1  gate1689(.a(G1081), .O(gate402inter8));
  nand2 gate1690(.a(gate402inter8), .b(gate402inter7), .O(gate402inter9));
  nand2 gate1691(.a(s_163), .b(gate402inter3), .O(gate402inter10));
  nor2  gate1692(.a(gate402inter10), .b(gate402inter9), .O(gate402inter11));
  nor2  gate1693(.a(gate402inter11), .b(gate402inter6), .O(gate402inter12));
  nand2 gate1694(.a(gate402inter12), .b(gate402inter1), .O(G1177));
nand2 gate403( .a(G17), .b(G1084), .O(G1180) );
nand2 gate404( .a(G18), .b(G1087), .O(G1183) );

  xor2  gate841(.a(G1090), .b(G19), .O(gate405inter0));
  nand2 gate842(.a(gate405inter0), .b(s_42), .O(gate405inter1));
  and2  gate843(.a(G1090), .b(G19), .O(gate405inter2));
  inv1  gate844(.a(s_42), .O(gate405inter3));
  inv1  gate845(.a(s_43), .O(gate405inter4));
  nand2 gate846(.a(gate405inter4), .b(gate405inter3), .O(gate405inter5));
  nor2  gate847(.a(gate405inter5), .b(gate405inter2), .O(gate405inter6));
  inv1  gate848(.a(G19), .O(gate405inter7));
  inv1  gate849(.a(G1090), .O(gate405inter8));
  nand2 gate850(.a(gate405inter8), .b(gate405inter7), .O(gate405inter9));
  nand2 gate851(.a(s_43), .b(gate405inter3), .O(gate405inter10));
  nor2  gate852(.a(gate405inter10), .b(gate405inter9), .O(gate405inter11));
  nor2  gate853(.a(gate405inter11), .b(gate405inter6), .O(gate405inter12));
  nand2 gate854(.a(gate405inter12), .b(gate405inter1), .O(G1186));

  xor2  gate1121(.a(G1093), .b(G20), .O(gate406inter0));
  nand2 gate1122(.a(gate406inter0), .b(s_82), .O(gate406inter1));
  and2  gate1123(.a(G1093), .b(G20), .O(gate406inter2));
  inv1  gate1124(.a(s_82), .O(gate406inter3));
  inv1  gate1125(.a(s_83), .O(gate406inter4));
  nand2 gate1126(.a(gate406inter4), .b(gate406inter3), .O(gate406inter5));
  nor2  gate1127(.a(gate406inter5), .b(gate406inter2), .O(gate406inter6));
  inv1  gate1128(.a(G20), .O(gate406inter7));
  inv1  gate1129(.a(G1093), .O(gate406inter8));
  nand2 gate1130(.a(gate406inter8), .b(gate406inter7), .O(gate406inter9));
  nand2 gate1131(.a(s_83), .b(gate406inter3), .O(gate406inter10));
  nor2  gate1132(.a(gate406inter10), .b(gate406inter9), .O(gate406inter11));
  nor2  gate1133(.a(gate406inter11), .b(gate406inter6), .O(gate406inter12));
  nand2 gate1134(.a(gate406inter12), .b(gate406inter1), .O(G1189));
nand2 gate407( .a(G21), .b(G1096), .O(G1192) );
nand2 gate408( .a(G22), .b(G1099), .O(G1195) );

  xor2  gate911(.a(G1102), .b(G23), .O(gate409inter0));
  nand2 gate912(.a(gate409inter0), .b(s_52), .O(gate409inter1));
  and2  gate913(.a(G1102), .b(G23), .O(gate409inter2));
  inv1  gate914(.a(s_52), .O(gate409inter3));
  inv1  gate915(.a(s_53), .O(gate409inter4));
  nand2 gate916(.a(gate409inter4), .b(gate409inter3), .O(gate409inter5));
  nor2  gate917(.a(gate409inter5), .b(gate409inter2), .O(gate409inter6));
  inv1  gate918(.a(G23), .O(gate409inter7));
  inv1  gate919(.a(G1102), .O(gate409inter8));
  nand2 gate920(.a(gate409inter8), .b(gate409inter7), .O(gate409inter9));
  nand2 gate921(.a(s_53), .b(gate409inter3), .O(gate409inter10));
  nor2  gate922(.a(gate409inter10), .b(gate409inter9), .O(gate409inter11));
  nor2  gate923(.a(gate409inter11), .b(gate409inter6), .O(gate409inter12));
  nand2 gate924(.a(gate409inter12), .b(gate409inter1), .O(G1198));
nand2 gate410( .a(G24), .b(G1105), .O(G1201) );
nand2 gate411( .a(G25), .b(G1108), .O(G1204) );
nand2 gate412( .a(G26), .b(G1111), .O(G1207) );
nand2 gate413( .a(G27), .b(G1114), .O(G1210) );
nand2 gate414( .a(G28), .b(G1117), .O(G1213) );

  xor2  gate1331(.a(G1120), .b(G29), .O(gate415inter0));
  nand2 gate1332(.a(gate415inter0), .b(s_112), .O(gate415inter1));
  and2  gate1333(.a(G1120), .b(G29), .O(gate415inter2));
  inv1  gate1334(.a(s_112), .O(gate415inter3));
  inv1  gate1335(.a(s_113), .O(gate415inter4));
  nand2 gate1336(.a(gate415inter4), .b(gate415inter3), .O(gate415inter5));
  nor2  gate1337(.a(gate415inter5), .b(gate415inter2), .O(gate415inter6));
  inv1  gate1338(.a(G29), .O(gate415inter7));
  inv1  gate1339(.a(G1120), .O(gate415inter8));
  nand2 gate1340(.a(gate415inter8), .b(gate415inter7), .O(gate415inter9));
  nand2 gate1341(.a(s_113), .b(gate415inter3), .O(gate415inter10));
  nor2  gate1342(.a(gate415inter10), .b(gate415inter9), .O(gate415inter11));
  nor2  gate1343(.a(gate415inter11), .b(gate415inter6), .O(gate415inter12));
  nand2 gate1344(.a(gate415inter12), .b(gate415inter1), .O(G1216));
nand2 gate416( .a(G30), .b(G1123), .O(G1219) );
nand2 gate417( .a(G31), .b(G1126), .O(G1222) );
nand2 gate418( .a(G32), .b(G1129), .O(G1225) );
nand2 gate419( .a(G1), .b(G1132), .O(G1228) );

  xor2  gate1765(.a(G1132), .b(G1036), .O(gate420inter0));
  nand2 gate1766(.a(gate420inter0), .b(s_174), .O(gate420inter1));
  and2  gate1767(.a(G1132), .b(G1036), .O(gate420inter2));
  inv1  gate1768(.a(s_174), .O(gate420inter3));
  inv1  gate1769(.a(s_175), .O(gate420inter4));
  nand2 gate1770(.a(gate420inter4), .b(gate420inter3), .O(gate420inter5));
  nor2  gate1771(.a(gate420inter5), .b(gate420inter2), .O(gate420inter6));
  inv1  gate1772(.a(G1036), .O(gate420inter7));
  inv1  gate1773(.a(G1132), .O(gate420inter8));
  nand2 gate1774(.a(gate420inter8), .b(gate420inter7), .O(gate420inter9));
  nand2 gate1775(.a(s_175), .b(gate420inter3), .O(gate420inter10));
  nor2  gate1776(.a(gate420inter10), .b(gate420inter9), .O(gate420inter11));
  nor2  gate1777(.a(gate420inter11), .b(gate420inter6), .O(gate420inter12));
  nand2 gate1778(.a(gate420inter12), .b(gate420inter1), .O(G1229));
nand2 gate421( .a(G2), .b(G1135), .O(G1230) );
nand2 gate422( .a(G1039), .b(G1135), .O(G1231) );
nand2 gate423( .a(G3), .b(G1138), .O(G1232) );

  xor2  gate1401(.a(G1138), .b(G1042), .O(gate424inter0));
  nand2 gate1402(.a(gate424inter0), .b(s_122), .O(gate424inter1));
  and2  gate1403(.a(G1138), .b(G1042), .O(gate424inter2));
  inv1  gate1404(.a(s_122), .O(gate424inter3));
  inv1  gate1405(.a(s_123), .O(gate424inter4));
  nand2 gate1406(.a(gate424inter4), .b(gate424inter3), .O(gate424inter5));
  nor2  gate1407(.a(gate424inter5), .b(gate424inter2), .O(gate424inter6));
  inv1  gate1408(.a(G1042), .O(gate424inter7));
  inv1  gate1409(.a(G1138), .O(gate424inter8));
  nand2 gate1410(.a(gate424inter8), .b(gate424inter7), .O(gate424inter9));
  nand2 gate1411(.a(s_123), .b(gate424inter3), .O(gate424inter10));
  nor2  gate1412(.a(gate424inter10), .b(gate424inter9), .O(gate424inter11));
  nor2  gate1413(.a(gate424inter11), .b(gate424inter6), .O(gate424inter12));
  nand2 gate1414(.a(gate424inter12), .b(gate424inter1), .O(G1233));
nand2 gate425( .a(G4), .b(G1141), .O(G1234) );
nand2 gate426( .a(G1045), .b(G1141), .O(G1235) );
nand2 gate427( .a(G5), .b(G1144), .O(G1236) );
nand2 gate428( .a(G1048), .b(G1144), .O(G1237) );
nand2 gate429( .a(G6), .b(G1147), .O(G1238) );
nand2 gate430( .a(G1051), .b(G1147), .O(G1239) );
nand2 gate431( .a(G7), .b(G1150), .O(G1240) );

  xor2  gate2003(.a(G1150), .b(G1054), .O(gate432inter0));
  nand2 gate2004(.a(gate432inter0), .b(s_208), .O(gate432inter1));
  and2  gate2005(.a(G1150), .b(G1054), .O(gate432inter2));
  inv1  gate2006(.a(s_208), .O(gate432inter3));
  inv1  gate2007(.a(s_209), .O(gate432inter4));
  nand2 gate2008(.a(gate432inter4), .b(gate432inter3), .O(gate432inter5));
  nor2  gate2009(.a(gate432inter5), .b(gate432inter2), .O(gate432inter6));
  inv1  gate2010(.a(G1054), .O(gate432inter7));
  inv1  gate2011(.a(G1150), .O(gate432inter8));
  nand2 gate2012(.a(gate432inter8), .b(gate432inter7), .O(gate432inter9));
  nand2 gate2013(.a(s_209), .b(gate432inter3), .O(gate432inter10));
  nor2  gate2014(.a(gate432inter10), .b(gate432inter9), .O(gate432inter11));
  nor2  gate2015(.a(gate432inter11), .b(gate432inter6), .O(gate432inter12));
  nand2 gate2016(.a(gate432inter12), .b(gate432inter1), .O(G1241));
nand2 gate433( .a(G8), .b(G1153), .O(G1242) );
nand2 gate434( .a(G1057), .b(G1153), .O(G1243) );
nand2 gate435( .a(G9), .b(G1156), .O(G1244) );
nand2 gate436( .a(G1060), .b(G1156), .O(G1245) );

  xor2  gate1989(.a(G1159), .b(G10), .O(gate437inter0));
  nand2 gate1990(.a(gate437inter0), .b(s_206), .O(gate437inter1));
  and2  gate1991(.a(G1159), .b(G10), .O(gate437inter2));
  inv1  gate1992(.a(s_206), .O(gate437inter3));
  inv1  gate1993(.a(s_207), .O(gate437inter4));
  nand2 gate1994(.a(gate437inter4), .b(gate437inter3), .O(gate437inter5));
  nor2  gate1995(.a(gate437inter5), .b(gate437inter2), .O(gate437inter6));
  inv1  gate1996(.a(G10), .O(gate437inter7));
  inv1  gate1997(.a(G1159), .O(gate437inter8));
  nand2 gate1998(.a(gate437inter8), .b(gate437inter7), .O(gate437inter9));
  nand2 gate1999(.a(s_207), .b(gate437inter3), .O(gate437inter10));
  nor2  gate2000(.a(gate437inter10), .b(gate437inter9), .O(gate437inter11));
  nor2  gate2001(.a(gate437inter11), .b(gate437inter6), .O(gate437inter12));
  nand2 gate2002(.a(gate437inter12), .b(gate437inter1), .O(G1246));
nand2 gate438( .a(G1063), .b(G1159), .O(G1247) );

  xor2  gate1345(.a(G1162), .b(G11), .O(gate439inter0));
  nand2 gate1346(.a(gate439inter0), .b(s_114), .O(gate439inter1));
  and2  gate1347(.a(G1162), .b(G11), .O(gate439inter2));
  inv1  gate1348(.a(s_114), .O(gate439inter3));
  inv1  gate1349(.a(s_115), .O(gate439inter4));
  nand2 gate1350(.a(gate439inter4), .b(gate439inter3), .O(gate439inter5));
  nor2  gate1351(.a(gate439inter5), .b(gate439inter2), .O(gate439inter6));
  inv1  gate1352(.a(G11), .O(gate439inter7));
  inv1  gate1353(.a(G1162), .O(gate439inter8));
  nand2 gate1354(.a(gate439inter8), .b(gate439inter7), .O(gate439inter9));
  nand2 gate1355(.a(s_115), .b(gate439inter3), .O(gate439inter10));
  nor2  gate1356(.a(gate439inter10), .b(gate439inter9), .O(gate439inter11));
  nor2  gate1357(.a(gate439inter11), .b(gate439inter6), .O(gate439inter12));
  nand2 gate1358(.a(gate439inter12), .b(gate439inter1), .O(G1248));

  xor2  gate1429(.a(G1162), .b(G1066), .O(gate440inter0));
  nand2 gate1430(.a(gate440inter0), .b(s_126), .O(gate440inter1));
  and2  gate1431(.a(G1162), .b(G1066), .O(gate440inter2));
  inv1  gate1432(.a(s_126), .O(gate440inter3));
  inv1  gate1433(.a(s_127), .O(gate440inter4));
  nand2 gate1434(.a(gate440inter4), .b(gate440inter3), .O(gate440inter5));
  nor2  gate1435(.a(gate440inter5), .b(gate440inter2), .O(gate440inter6));
  inv1  gate1436(.a(G1066), .O(gate440inter7));
  inv1  gate1437(.a(G1162), .O(gate440inter8));
  nand2 gate1438(.a(gate440inter8), .b(gate440inter7), .O(gate440inter9));
  nand2 gate1439(.a(s_127), .b(gate440inter3), .O(gate440inter10));
  nor2  gate1440(.a(gate440inter10), .b(gate440inter9), .O(gate440inter11));
  nor2  gate1441(.a(gate440inter11), .b(gate440inter6), .O(gate440inter12));
  nand2 gate1442(.a(gate440inter12), .b(gate440inter1), .O(G1249));

  xor2  gate659(.a(G1165), .b(G12), .O(gate441inter0));
  nand2 gate660(.a(gate441inter0), .b(s_16), .O(gate441inter1));
  and2  gate661(.a(G1165), .b(G12), .O(gate441inter2));
  inv1  gate662(.a(s_16), .O(gate441inter3));
  inv1  gate663(.a(s_17), .O(gate441inter4));
  nand2 gate664(.a(gate441inter4), .b(gate441inter3), .O(gate441inter5));
  nor2  gate665(.a(gate441inter5), .b(gate441inter2), .O(gate441inter6));
  inv1  gate666(.a(G12), .O(gate441inter7));
  inv1  gate667(.a(G1165), .O(gate441inter8));
  nand2 gate668(.a(gate441inter8), .b(gate441inter7), .O(gate441inter9));
  nand2 gate669(.a(s_17), .b(gate441inter3), .O(gate441inter10));
  nor2  gate670(.a(gate441inter10), .b(gate441inter9), .O(gate441inter11));
  nor2  gate671(.a(gate441inter11), .b(gate441inter6), .O(gate441inter12));
  nand2 gate672(.a(gate441inter12), .b(gate441inter1), .O(G1250));

  xor2  gate1289(.a(G1165), .b(G1069), .O(gate442inter0));
  nand2 gate1290(.a(gate442inter0), .b(s_106), .O(gate442inter1));
  and2  gate1291(.a(G1165), .b(G1069), .O(gate442inter2));
  inv1  gate1292(.a(s_106), .O(gate442inter3));
  inv1  gate1293(.a(s_107), .O(gate442inter4));
  nand2 gate1294(.a(gate442inter4), .b(gate442inter3), .O(gate442inter5));
  nor2  gate1295(.a(gate442inter5), .b(gate442inter2), .O(gate442inter6));
  inv1  gate1296(.a(G1069), .O(gate442inter7));
  inv1  gate1297(.a(G1165), .O(gate442inter8));
  nand2 gate1298(.a(gate442inter8), .b(gate442inter7), .O(gate442inter9));
  nand2 gate1299(.a(s_107), .b(gate442inter3), .O(gate442inter10));
  nor2  gate1300(.a(gate442inter10), .b(gate442inter9), .O(gate442inter11));
  nor2  gate1301(.a(gate442inter11), .b(gate442inter6), .O(gate442inter12));
  nand2 gate1302(.a(gate442inter12), .b(gate442inter1), .O(G1251));
nand2 gate443( .a(G13), .b(G1168), .O(G1252) );
nand2 gate444( .a(G1072), .b(G1168), .O(G1253) );

  xor2  gate1611(.a(G1171), .b(G14), .O(gate445inter0));
  nand2 gate1612(.a(gate445inter0), .b(s_152), .O(gate445inter1));
  and2  gate1613(.a(G1171), .b(G14), .O(gate445inter2));
  inv1  gate1614(.a(s_152), .O(gate445inter3));
  inv1  gate1615(.a(s_153), .O(gate445inter4));
  nand2 gate1616(.a(gate445inter4), .b(gate445inter3), .O(gate445inter5));
  nor2  gate1617(.a(gate445inter5), .b(gate445inter2), .O(gate445inter6));
  inv1  gate1618(.a(G14), .O(gate445inter7));
  inv1  gate1619(.a(G1171), .O(gate445inter8));
  nand2 gate1620(.a(gate445inter8), .b(gate445inter7), .O(gate445inter9));
  nand2 gate1621(.a(s_153), .b(gate445inter3), .O(gate445inter10));
  nor2  gate1622(.a(gate445inter10), .b(gate445inter9), .O(gate445inter11));
  nor2  gate1623(.a(gate445inter11), .b(gate445inter6), .O(gate445inter12));
  nand2 gate1624(.a(gate445inter12), .b(gate445inter1), .O(G1254));
nand2 gate446( .a(G1075), .b(G1171), .O(G1255) );
nand2 gate447( .a(G15), .b(G1174), .O(G1256) );
nand2 gate448( .a(G1078), .b(G1174), .O(G1257) );

  xor2  gate855(.a(G1177), .b(G16), .O(gate449inter0));
  nand2 gate856(.a(gate449inter0), .b(s_44), .O(gate449inter1));
  and2  gate857(.a(G1177), .b(G16), .O(gate449inter2));
  inv1  gate858(.a(s_44), .O(gate449inter3));
  inv1  gate859(.a(s_45), .O(gate449inter4));
  nand2 gate860(.a(gate449inter4), .b(gate449inter3), .O(gate449inter5));
  nor2  gate861(.a(gate449inter5), .b(gate449inter2), .O(gate449inter6));
  inv1  gate862(.a(G16), .O(gate449inter7));
  inv1  gate863(.a(G1177), .O(gate449inter8));
  nand2 gate864(.a(gate449inter8), .b(gate449inter7), .O(gate449inter9));
  nand2 gate865(.a(s_45), .b(gate449inter3), .O(gate449inter10));
  nor2  gate866(.a(gate449inter10), .b(gate449inter9), .O(gate449inter11));
  nor2  gate867(.a(gate449inter11), .b(gate449inter6), .O(gate449inter12));
  nand2 gate868(.a(gate449inter12), .b(gate449inter1), .O(G1258));
nand2 gate450( .a(G1081), .b(G1177), .O(G1259) );
nand2 gate451( .a(G17), .b(G1180), .O(G1260) );
nand2 gate452( .a(G1084), .b(G1180), .O(G1261) );
nand2 gate453( .a(G18), .b(G1183), .O(G1262) );
nand2 gate454( .a(G1087), .b(G1183), .O(G1263) );
nand2 gate455( .a(G19), .b(G1186), .O(G1264) );
nand2 gate456( .a(G1090), .b(G1186), .O(G1265) );
nand2 gate457( .a(G20), .b(G1189), .O(G1266) );
nand2 gate458( .a(G1093), .b(G1189), .O(G1267) );
nand2 gate459( .a(G21), .b(G1192), .O(G1268) );
nand2 gate460( .a(G1096), .b(G1192), .O(G1269) );

  xor2  gate1667(.a(G1195), .b(G22), .O(gate461inter0));
  nand2 gate1668(.a(gate461inter0), .b(s_160), .O(gate461inter1));
  and2  gate1669(.a(G1195), .b(G22), .O(gate461inter2));
  inv1  gate1670(.a(s_160), .O(gate461inter3));
  inv1  gate1671(.a(s_161), .O(gate461inter4));
  nand2 gate1672(.a(gate461inter4), .b(gate461inter3), .O(gate461inter5));
  nor2  gate1673(.a(gate461inter5), .b(gate461inter2), .O(gate461inter6));
  inv1  gate1674(.a(G22), .O(gate461inter7));
  inv1  gate1675(.a(G1195), .O(gate461inter8));
  nand2 gate1676(.a(gate461inter8), .b(gate461inter7), .O(gate461inter9));
  nand2 gate1677(.a(s_161), .b(gate461inter3), .O(gate461inter10));
  nor2  gate1678(.a(gate461inter10), .b(gate461inter9), .O(gate461inter11));
  nor2  gate1679(.a(gate461inter11), .b(gate461inter6), .O(gate461inter12));
  nand2 gate1680(.a(gate461inter12), .b(gate461inter1), .O(G1270));
nand2 gate462( .a(G1099), .b(G1195), .O(G1271) );
nand2 gate463( .a(G23), .b(G1198), .O(G1272) );
nand2 gate464( .a(G1102), .b(G1198), .O(G1273) );
nand2 gate465( .a(G24), .b(G1201), .O(G1274) );
nand2 gate466( .a(G1105), .b(G1201), .O(G1275) );
nand2 gate467( .a(G25), .b(G1204), .O(G1276) );
nand2 gate468( .a(G1108), .b(G1204), .O(G1277) );
nand2 gate469( .a(G26), .b(G1207), .O(G1278) );
nand2 gate470( .a(G1111), .b(G1207), .O(G1279) );
nand2 gate471( .a(G27), .b(G1210), .O(G1280) );
nand2 gate472( .a(G1114), .b(G1210), .O(G1281) );
nand2 gate473( .a(G28), .b(G1213), .O(G1282) );
nand2 gate474( .a(G1117), .b(G1213), .O(G1283) );
nand2 gate475( .a(G29), .b(G1216), .O(G1284) );
nand2 gate476( .a(G1120), .b(G1216), .O(G1285) );
nand2 gate477( .a(G30), .b(G1219), .O(G1286) );
nand2 gate478( .a(G1123), .b(G1219), .O(G1287) );

  xor2  gate1905(.a(G1222), .b(G31), .O(gate479inter0));
  nand2 gate1906(.a(gate479inter0), .b(s_194), .O(gate479inter1));
  and2  gate1907(.a(G1222), .b(G31), .O(gate479inter2));
  inv1  gate1908(.a(s_194), .O(gate479inter3));
  inv1  gate1909(.a(s_195), .O(gate479inter4));
  nand2 gate1910(.a(gate479inter4), .b(gate479inter3), .O(gate479inter5));
  nor2  gate1911(.a(gate479inter5), .b(gate479inter2), .O(gate479inter6));
  inv1  gate1912(.a(G31), .O(gate479inter7));
  inv1  gate1913(.a(G1222), .O(gate479inter8));
  nand2 gate1914(.a(gate479inter8), .b(gate479inter7), .O(gate479inter9));
  nand2 gate1915(.a(s_195), .b(gate479inter3), .O(gate479inter10));
  nor2  gate1916(.a(gate479inter10), .b(gate479inter9), .O(gate479inter11));
  nor2  gate1917(.a(gate479inter11), .b(gate479inter6), .O(gate479inter12));
  nand2 gate1918(.a(gate479inter12), .b(gate479inter1), .O(G1288));
nand2 gate480( .a(G1126), .b(G1222), .O(G1289) );

  xor2  gate1009(.a(G1225), .b(G32), .O(gate481inter0));
  nand2 gate1010(.a(gate481inter0), .b(s_66), .O(gate481inter1));
  and2  gate1011(.a(G1225), .b(G32), .O(gate481inter2));
  inv1  gate1012(.a(s_66), .O(gate481inter3));
  inv1  gate1013(.a(s_67), .O(gate481inter4));
  nand2 gate1014(.a(gate481inter4), .b(gate481inter3), .O(gate481inter5));
  nor2  gate1015(.a(gate481inter5), .b(gate481inter2), .O(gate481inter6));
  inv1  gate1016(.a(G32), .O(gate481inter7));
  inv1  gate1017(.a(G1225), .O(gate481inter8));
  nand2 gate1018(.a(gate481inter8), .b(gate481inter7), .O(gate481inter9));
  nand2 gate1019(.a(s_67), .b(gate481inter3), .O(gate481inter10));
  nor2  gate1020(.a(gate481inter10), .b(gate481inter9), .O(gate481inter11));
  nor2  gate1021(.a(gate481inter11), .b(gate481inter6), .O(gate481inter12));
  nand2 gate1022(.a(gate481inter12), .b(gate481inter1), .O(G1290));
nand2 gate482( .a(G1129), .b(G1225), .O(G1291) );
nand2 gate483( .a(G1228), .b(G1229), .O(G1292) );
nand2 gate484( .a(G1230), .b(G1231), .O(G1293) );
nand2 gate485( .a(G1232), .b(G1233), .O(G1294) );
nand2 gate486( .a(G1234), .b(G1235), .O(G1295) );
nand2 gate487( .a(G1236), .b(G1237), .O(G1296) );
nand2 gate488( .a(G1238), .b(G1239), .O(G1297) );
nand2 gate489( .a(G1240), .b(G1241), .O(G1298) );

  xor2  gate1191(.a(G1243), .b(G1242), .O(gate490inter0));
  nand2 gate1192(.a(gate490inter0), .b(s_92), .O(gate490inter1));
  and2  gate1193(.a(G1243), .b(G1242), .O(gate490inter2));
  inv1  gate1194(.a(s_92), .O(gate490inter3));
  inv1  gate1195(.a(s_93), .O(gate490inter4));
  nand2 gate1196(.a(gate490inter4), .b(gate490inter3), .O(gate490inter5));
  nor2  gate1197(.a(gate490inter5), .b(gate490inter2), .O(gate490inter6));
  inv1  gate1198(.a(G1242), .O(gate490inter7));
  inv1  gate1199(.a(G1243), .O(gate490inter8));
  nand2 gate1200(.a(gate490inter8), .b(gate490inter7), .O(gate490inter9));
  nand2 gate1201(.a(s_93), .b(gate490inter3), .O(gate490inter10));
  nor2  gate1202(.a(gate490inter10), .b(gate490inter9), .O(gate490inter11));
  nor2  gate1203(.a(gate490inter11), .b(gate490inter6), .O(gate490inter12));
  nand2 gate1204(.a(gate490inter12), .b(gate490inter1), .O(G1299));
nand2 gate491( .a(G1244), .b(G1245), .O(G1300) );
nand2 gate492( .a(G1246), .b(G1247), .O(G1301) );
nand2 gate493( .a(G1248), .b(G1249), .O(G1302) );

  xor2  gate1933(.a(G1251), .b(G1250), .O(gate494inter0));
  nand2 gate1934(.a(gate494inter0), .b(s_198), .O(gate494inter1));
  and2  gate1935(.a(G1251), .b(G1250), .O(gate494inter2));
  inv1  gate1936(.a(s_198), .O(gate494inter3));
  inv1  gate1937(.a(s_199), .O(gate494inter4));
  nand2 gate1938(.a(gate494inter4), .b(gate494inter3), .O(gate494inter5));
  nor2  gate1939(.a(gate494inter5), .b(gate494inter2), .O(gate494inter6));
  inv1  gate1940(.a(G1250), .O(gate494inter7));
  inv1  gate1941(.a(G1251), .O(gate494inter8));
  nand2 gate1942(.a(gate494inter8), .b(gate494inter7), .O(gate494inter9));
  nand2 gate1943(.a(s_199), .b(gate494inter3), .O(gate494inter10));
  nor2  gate1944(.a(gate494inter10), .b(gate494inter9), .O(gate494inter11));
  nor2  gate1945(.a(gate494inter11), .b(gate494inter6), .O(gate494inter12));
  nand2 gate1946(.a(gate494inter12), .b(gate494inter1), .O(G1303));
nand2 gate495( .a(G1252), .b(G1253), .O(G1304) );
nand2 gate496( .a(G1254), .b(G1255), .O(G1305) );

  xor2  gate2017(.a(G1257), .b(G1256), .O(gate497inter0));
  nand2 gate2018(.a(gate497inter0), .b(s_210), .O(gate497inter1));
  and2  gate2019(.a(G1257), .b(G1256), .O(gate497inter2));
  inv1  gate2020(.a(s_210), .O(gate497inter3));
  inv1  gate2021(.a(s_211), .O(gate497inter4));
  nand2 gate2022(.a(gate497inter4), .b(gate497inter3), .O(gate497inter5));
  nor2  gate2023(.a(gate497inter5), .b(gate497inter2), .O(gate497inter6));
  inv1  gate2024(.a(G1256), .O(gate497inter7));
  inv1  gate2025(.a(G1257), .O(gate497inter8));
  nand2 gate2026(.a(gate497inter8), .b(gate497inter7), .O(gate497inter9));
  nand2 gate2027(.a(s_211), .b(gate497inter3), .O(gate497inter10));
  nor2  gate2028(.a(gate497inter10), .b(gate497inter9), .O(gate497inter11));
  nor2  gate2029(.a(gate497inter11), .b(gate497inter6), .O(gate497inter12));
  nand2 gate2030(.a(gate497inter12), .b(gate497inter1), .O(G1306));
nand2 gate498( .a(G1258), .b(G1259), .O(G1307) );
nand2 gate499( .a(G1260), .b(G1261), .O(G1308) );
nand2 gate500( .a(G1262), .b(G1263), .O(G1309) );
nand2 gate501( .a(G1264), .b(G1265), .O(G1310) );
nand2 gate502( .a(G1266), .b(G1267), .O(G1311) );
nand2 gate503( .a(G1268), .b(G1269), .O(G1312) );

  xor2  gate1513(.a(G1271), .b(G1270), .O(gate504inter0));
  nand2 gate1514(.a(gate504inter0), .b(s_138), .O(gate504inter1));
  and2  gate1515(.a(G1271), .b(G1270), .O(gate504inter2));
  inv1  gate1516(.a(s_138), .O(gate504inter3));
  inv1  gate1517(.a(s_139), .O(gate504inter4));
  nand2 gate1518(.a(gate504inter4), .b(gate504inter3), .O(gate504inter5));
  nor2  gate1519(.a(gate504inter5), .b(gate504inter2), .O(gate504inter6));
  inv1  gate1520(.a(G1270), .O(gate504inter7));
  inv1  gate1521(.a(G1271), .O(gate504inter8));
  nand2 gate1522(.a(gate504inter8), .b(gate504inter7), .O(gate504inter9));
  nand2 gate1523(.a(s_139), .b(gate504inter3), .O(gate504inter10));
  nor2  gate1524(.a(gate504inter10), .b(gate504inter9), .O(gate504inter11));
  nor2  gate1525(.a(gate504inter11), .b(gate504inter6), .O(gate504inter12));
  nand2 gate1526(.a(gate504inter12), .b(gate504inter1), .O(G1313));
nand2 gate505( .a(G1272), .b(G1273), .O(G1314) );
nand2 gate506( .a(G1274), .b(G1275), .O(G1315) );

  xor2  gate1275(.a(G1277), .b(G1276), .O(gate507inter0));
  nand2 gate1276(.a(gate507inter0), .b(s_104), .O(gate507inter1));
  and2  gate1277(.a(G1277), .b(G1276), .O(gate507inter2));
  inv1  gate1278(.a(s_104), .O(gate507inter3));
  inv1  gate1279(.a(s_105), .O(gate507inter4));
  nand2 gate1280(.a(gate507inter4), .b(gate507inter3), .O(gate507inter5));
  nor2  gate1281(.a(gate507inter5), .b(gate507inter2), .O(gate507inter6));
  inv1  gate1282(.a(G1276), .O(gate507inter7));
  inv1  gate1283(.a(G1277), .O(gate507inter8));
  nand2 gate1284(.a(gate507inter8), .b(gate507inter7), .O(gate507inter9));
  nand2 gate1285(.a(s_105), .b(gate507inter3), .O(gate507inter10));
  nor2  gate1286(.a(gate507inter10), .b(gate507inter9), .O(gate507inter11));
  nor2  gate1287(.a(gate507inter11), .b(gate507inter6), .O(gate507inter12));
  nand2 gate1288(.a(gate507inter12), .b(gate507inter1), .O(G1316));
nand2 gate508( .a(G1278), .b(G1279), .O(G1317) );
nand2 gate509( .a(G1280), .b(G1281), .O(G1318) );
nand2 gate510( .a(G1282), .b(G1283), .O(G1319) );
nand2 gate511( .a(G1284), .b(G1285), .O(G1320) );

  xor2  gate1947(.a(G1287), .b(G1286), .O(gate512inter0));
  nand2 gate1948(.a(gate512inter0), .b(s_200), .O(gate512inter1));
  and2  gate1949(.a(G1287), .b(G1286), .O(gate512inter2));
  inv1  gate1950(.a(s_200), .O(gate512inter3));
  inv1  gate1951(.a(s_201), .O(gate512inter4));
  nand2 gate1952(.a(gate512inter4), .b(gate512inter3), .O(gate512inter5));
  nor2  gate1953(.a(gate512inter5), .b(gate512inter2), .O(gate512inter6));
  inv1  gate1954(.a(G1286), .O(gate512inter7));
  inv1  gate1955(.a(G1287), .O(gate512inter8));
  nand2 gate1956(.a(gate512inter8), .b(gate512inter7), .O(gate512inter9));
  nand2 gate1957(.a(s_201), .b(gate512inter3), .O(gate512inter10));
  nor2  gate1958(.a(gate512inter10), .b(gate512inter9), .O(gate512inter11));
  nor2  gate1959(.a(gate512inter11), .b(gate512inter6), .O(gate512inter12));
  nand2 gate1960(.a(gate512inter12), .b(gate512inter1), .O(G1321));

  xor2  gate687(.a(G1289), .b(G1288), .O(gate513inter0));
  nand2 gate688(.a(gate513inter0), .b(s_20), .O(gate513inter1));
  and2  gate689(.a(G1289), .b(G1288), .O(gate513inter2));
  inv1  gate690(.a(s_20), .O(gate513inter3));
  inv1  gate691(.a(s_21), .O(gate513inter4));
  nand2 gate692(.a(gate513inter4), .b(gate513inter3), .O(gate513inter5));
  nor2  gate693(.a(gate513inter5), .b(gate513inter2), .O(gate513inter6));
  inv1  gate694(.a(G1288), .O(gate513inter7));
  inv1  gate695(.a(G1289), .O(gate513inter8));
  nand2 gate696(.a(gate513inter8), .b(gate513inter7), .O(gate513inter9));
  nand2 gate697(.a(s_21), .b(gate513inter3), .O(gate513inter10));
  nor2  gate698(.a(gate513inter10), .b(gate513inter9), .O(gate513inter11));
  nor2  gate699(.a(gate513inter11), .b(gate513inter6), .O(gate513inter12));
  nand2 gate700(.a(gate513inter12), .b(gate513inter1), .O(G1322));
nand2 gate514( .a(G1290), .b(G1291), .O(G1323) );
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule