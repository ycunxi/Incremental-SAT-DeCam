module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);

input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;//RE__PI;

input s_0,s_1;//RE__ALLOW(00,01,10,11);
input s_2,s_3;//RE__ALLOW(00,01,10,11);
input s_4,s_5;//RE__ALLOW(00,01,10,11);
input s_6,s_7;//RE__ALLOW(00,01,10,11);
input s_8,s_9;//RE__ALLOW(00,01,10,11);
input s_10,s_11;//RE__ALLOW(00,01,10,11);
input s_12,s_13;//RE__ALLOW(00,01,10,11);
input s_14,s_15;//RE__ALLOW(00,01,10,11);
input s_16,s_17;//RE__ALLOW(00,01,10,11);
input s_18,s_19;//RE__ALLOW(00,01,10,11);
input s_20,s_21;//RE__ALLOW(00,01,10,11);
input s_22,s_23;//RE__ALLOW(00,01,10,11);
input s_24,s_25;//RE__ALLOW(00,01,10,11);
input s_26,s_27;//RE__ALLOW(00,01,10,11);
input s_28,s_29;//RE__ALLOW(00,01,10,11);
input s_30,s_31;//RE__ALLOW(00,01,10,11);
input s_32,s_33;//RE__ALLOW(00,01,10,11);
input s_34,s_35;//RE__ALLOW(00,01,10,11);
input s_36,s_37;//RE__ALLOW(00,01,10,11);
input s_38,s_39;//RE__ALLOW(00,01,10,11);
input s_40,s_41;//RE__ALLOW(00,01,10,11);
input s_42,s_43;//RE__ALLOW(00,01,10,11);
input s_44,s_45;//RE__ALLOW(00,01,10,11);
input s_46,s_47;//RE__ALLOW(00,01,10,11);
input s_48,s_49;//RE__ALLOW(00,01,10,11);
input s_50,s_51;//RE__ALLOW(00,01,10,11);
input s_52,s_53;//RE__ALLOW(00,01,10,11);
input s_54,s_55;//RE__ALLOW(00,01,10,11);
input s_56,s_57;//RE__ALLOW(00,01,10,11);
input s_58,s_59;//RE__ALLOW(00,01,10,11);
input s_60,s_61;//RE__ALLOW(00,01,10,11);
input s_62,s_63;//RE__ALLOW(00,01,10,11);
input s_64,s_65;//RE__ALLOW(00,01,10,11);
input s_66,s_67;//RE__ALLOW(00,01,10,11);
input s_68,s_69;//RE__ALLOW(00,01,10,11);
input s_70,s_71;//RE__ALLOW(00,01,10,11);
input s_72,s_73;//RE__ALLOW(00,01,10,11);
input s_74,s_75;//RE__ALLOW(00,01,10,11);
input s_76,s_77;//RE__ALLOW(00,01,10,11);
input s_78,s_79;//RE__ALLOW(00,01,10,11);
input s_80,s_81;//RE__ALLOW(00,01,10,11);
input s_82,s_83;//RE__ALLOW(00,01,10,11);
input s_84,s_85;//RE__ALLOW(00,01,10,11);
input s_86,s_87;//RE__ALLOW(00,01,10,11);
input s_88,s_89;//RE__ALLOW(00,01,10,11);
input s_90,s_91;//RE__ALLOW(00,01,10,11);
input s_92,s_93;//RE__ALLOW(00,01,10,11);
input s_94,s_95;//RE__ALLOW(00,01,10,11);
input s_96,s_97;//RE__ALLOW(00,01,10,11);
input s_98,s_99;//RE__ALLOW(00,01,10,11);
input s_100,s_101;//RE__ALLOW(00,01,10,11);
input s_102,s_103;//RE__ALLOW(00,01,10,11);
input s_104,s_105;//RE__ALLOW(00,01,10,11);
input s_106,s_107;//RE__ALLOW(00,01,10,11);
input s_108,s_109;//RE__ALLOW(00,01,10,11);
input s_110,s_111;//RE__ALLOW(00,01,10,11);
input s_112,s_113;//RE__ALLOW(00,01,10,11);
input s_114,s_115;//RE__ALLOW(00,01,10,11);
input s_116,s_117;//RE__ALLOW(00,01,10,11);
input s_118,s_119;//RE__ALLOW(00,01,10,11);
input s_120,s_121;//RE__ALLOW(00,01,10,11);
input s_122,s_123;//RE__ALLOW(00,01,10,11);
input s_124,s_125;//RE__ALLOW(00,01,10,11);
input s_126,s_127;//RE__ALLOW(00,01,10,11);
input s_128,s_129;//RE__ALLOW(00,01,10,11);
input s_130,s_131;//RE__ALLOW(00,01,10,11);
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;

  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate206inter0, gate206inter1, gate206inter2, gate206inter3, gate206inter4, gate206inter5, gate206inter6, gate206inter7, gate206inter8, gate206inter9, gate206inter10, gate206inter11, gate206inter12, gate296inter0, gate296inter1, gate296inter2, gate296inter3, gate296inter4, gate296inter5, gate296inter6, gate296inter7, gate296inter8, gate296inter9, gate296inter10, gate296inter11, gate296inter12, gate29inter0, gate29inter1, gate29inter2, gate29inter3, gate29inter4, gate29inter5, gate29inter6, gate29inter7, gate29inter8, gate29inter9, gate29inter10, gate29inter11, gate29inter12, gate412inter0, gate412inter1, gate412inter2, gate412inter3, gate412inter4, gate412inter5, gate412inter6, gate412inter7, gate412inter8, gate412inter9, gate412inter10, gate412inter11, gate412inter12, gate115inter0, gate115inter1, gate115inter2, gate115inter3, gate115inter4, gate115inter5, gate115inter6, gate115inter7, gate115inter8, gate115inter9, gate115inter10, gate115inter11, gate115inter12, gate264inter0, gate264inter1, gate264inter2, gate264inter3, gate264inter4, gate264inter5, gate264inter6, gate264inter7, gate264inter8, gate264inter9, gate264inter10, gate264inter11, gate264inter12, gate398inter0, gate398inter1, gate398inter2, gate398inter3, gate398inter4, gate398inter5, gate398inter6, gate398inter7, gate398inter8, gate398inter9, gate398inter10, gate398inter11, gate398inter12, gate24inter0, gate24inter1, gate24inter2, gate24inter3, gate24inter4, gate24inter5, gate24inter6, gate24inter7, gate24inter8, gate24inter9, gate24inter10, gate24inter11, gate24inter12, gate460inter0, gate460inter1, gate460inter2, gate460inter3, gate460inter4, gate460inter5, gate460inter6, gate460inter7, gate460inter8, gate460inter9, gate460inter10, gate460inter11, gate460inter12, gate197inter0, gate197inter1, gate197inter2, gate197inter3, gate197inter4, gate197inter5, gate197inter6, gate197inter7, gate197inter8, gate197inter9, gate197inter10, gate197inter11, gate197inter12, gate141inter0, gate141inter1, gate141inter2, gate141inter3, gate141inter4, gate141inter5, gate141inter6, gate141inter7, gate141inter8, gate141inter9, gate141inter10, gate141inter11, gate141inter12, gate491inter0, gate491inter1, gate491inter2, gate491inter3, gate491inter4, gate491inter5, gate491inter6, gate491inter7, gate491inter8, gate491inter9, gate491inter10, gate491inter11, gate491inter12, gate410inter0, gate410inter1, gate410inter2, gate410inter3, gate410inter4, gate410inter5, gate410inter6, gate410inter7, gate410inter8, gate410inter9, gate410inter10, gate410inter11, gate410inter12, gate278inter0, gate278inter1, gate278inter2, gate278inter3, gate278inter4, gate278inter5, gate278inter6, gate278inter7, gate278inter8, gate278inter9, gate278inter10, gate278inter11, gate278inter12, gate110inter0, gate110inter1, gate110inter2, gate110inter3, gate110inter4, gate110inter5, gate110inter6, gate110inter7, gate110inter8, gate110inter9, gate110inter10, gate110inter11, gate110inter12, gate464inter0, gate464inter1, gate464inter2, gate464inter3, gate464inter4, gate464inter5, gate464inter6, gate464inter7, gate464inter8, gate464inter9, gate464inter10, gate464inter11, gate464inter12, gate417inter0, gate417inter1, gate417inter2, gate417inter3, gate417inter4, gate417inter5, gate417inter6, gate417inter7, gate417inter8, gate417inter9, gate417inter10, gate417inter11, gate417inter12, gate471inter0, gate471inter1, gate471inter2, gate471inter3, gate471inter4, gate471inter5, gate471inter6, gate471inter7, gate471inter8, gate471inter9, gate471inter10, gate471inter11, gate471inter12, gate131inter0, gate131inter1, gate131inter2, gate131inter3, gate131inter4, gate131inter5, gate131inter6, gate131inter7, gate131inter8, gate131inter9, gate131inter10, gate131inter11, gate131inter12, gate403inter0, gate403inter1, gate403inter2, gate403inter3, gate403inter4, gate403inter5, gate403inter6, gate403inter7, gate403inter8, gate403inter9, gate403inter10, gate403inter11, gate403inter12, gate111inter0, gate111inter1, gate111inter2, gate111inter3, gate111inter4, gate111inter5, gate111inter6, gate111inter7, gate111inter8, gate111inter9, gate111inter10, gate111inter11, gate111inter12, gate84inter0, gate84inter1, gate84inter2, gate84inter3, gate84inter4, gate84inter5, gate84inter6, gate84inter7, gate84inter8, gate84inter9, gate84inter10, gate84inter11, gate84inter12, gate187inter0, gate187inter1, gate187inter2, gate187inter3, gate187inter4, gate187inter5, gate187inter6, gate187inter7, gate187inter8, gate187inter9, gate187inter10, gate187inter11, gate187inter12, gate154inter0, gate154inter1, gate154inter2, gate154inter3, gate154inter4, gate154inter5, gate154inter6, gate154inter7, gate154inter8, gate154inter9, gate154inter10, gate154inter11, gate154inter12, gate218inter0, gate218inter1, gate218inter2, gate218inter3, gate218inter4, gate218inter5, gate218inter6, gate218inter7, gate218inter8, gate218inter9, gate218inter10, gate218inter11, gate218inter12, gate38inter0, gate38inter1, gate38inter2, gate38inter3, gate38inter4, gate38inter5, gate38inter6, gate38inter7, gate38inter8, gate38inter9, gate38inter10, gate38inter11, gate38inter12, gate489inter0, gate489inter1, gate489inter2, gate489inter3, gate489inter4, gate489inter5, gate489inter6, gate489inter7, gate489inter8, gate489inter9, gate489inter10, gate489inter11, gate489inter12, gate432inter0, gate432inter1, gate432inter2, gate432inter3, gate432inter4, gate432inter5, gate432inter6, gate432inter7, gate432inter8, gate432inter9, gate432inter10, gate432inter11, gate432inter12, gate291inter0, gate291inter1, gate291inter2, gate291inter3, gate291inter4, gate291inter5, gate291inter6, gate291inter7, gate291inter8, gate291inter9, gate291inter10, gate291inter11, gate291inter12, gate484inter0, gate484inter1, gate484inter2, gate484inter3, gate484inter4, gate484inter5, gate484inter6, gate484inter7, gate484inter8, gate484inter9, gate484inter10, gate484inter11, gate484inter12, gate23inter0, gate23inter1, gate23inter2, gate23inter3, gate23inter4, gate23inter5, gate23inter6, gate23inter7, gate23inter8, gate23inter9, gate23inter10, gate23inter11, gate23inter12, gate27inter0, gate27inter1, gate27inter2, gate27inter3, gate27inter4, gate27inter5, gate27inter6, gate27inter7, gate27inter8, gate27inter9, gate27inter10, gate27inter11, gate27inter12, gate98inter0, gate98inter1, gate98inter2, gate98inter3, gate98inter4, gate98inter5, gate98inter6, gate98inter7, gate98inter8, gate98inter9, gate98inter10, gate98inter11, gate98inter12, gate231inter0, gate231inter1, gate231inter2, gate231inter3, gate231inter4, gate231inter5, gate231inter6, gate231inter7, gate231inter8, gate231inter9, gate231inter10, gate231inter11, gate231inter12, gate237inter0, gate237inter1, gate237inter2, gate237inter3, gate237inter4, gate237inter5, gate237inter6, gate237inter7, gate237inter8, gate237inter9, gate237inter10, gate237inter11, gate237inter12, gate95inter0, gate95inter1, gate95inter2, gate95inter3, gate95inter4, gate95inter5, gate95inter6, gate95inter7, gate95inter8, gate95inter9, gate95inter10, gate95inter11, gate95inter12, gate413inter0, gate413inter1, gate413inter2, gate413inter3, gate413inter4, gate413inter5, gate413inter6, gate413inter7, gate413inter8, gate413inter9, gate413inter10, gate413inter11, gate413inter12, gate132inter0, gate132inter1, gate132inter2, gate132inter3, gate132inter4, gate132inter5, gate132inter6, gate132inter7, gate132inter8, gate132inter9, gate132inter10, gate132inter11, gate132inter12, gate107inter0, gate107inter1, gate107inter2, gate107inter3, gate107inter4, gate107inter5, gate107inter6, gate107inter7, gate107inter8, gate107inter9, gate107inter10, gate107inter11, gate107inter12, gate53inter0, gate53inter1, gate53inter2, gate53inter3, gate53inter4, gate53inter5, gate53inter6, gate53inter7, gate53inter8, gate53inter9, gate53inter10, gate53inter11, gate53inter12, gate180inter0, gate180inter1, gate180inter2, gate180inter3, gate180inter4, gate180inter5, gate180inter6, gate180inter7, gate180inter8, gate180inter9, gate180inter10, gate180inter11, gate180inter12, gate189inter0, gate189inter1, gate189inter2, gate189inter3, gate189inter4, gate189inter5, gate189inter6, gate189inter7, gate189inter8, gate189inter9, gate189inter10, gate189inter11, gate189inter12, gate170inter0, gate170inter1, gate170inter2, gate170inter3, gate170inter4, gate170inter5, gate170inter6, gate170inter7, gate170inter8, gate170inter9, gate170inter10, gate170inter11, gate170inter12, gate66inter0, gate66inter1, gate66inter2, gate66inter3, gate66inter4, gate66inter5, gate66inter6, gate66inter7, gate66inter8, gate66inter9, gate66inter10, gate66inter11, gate66inter12, gate43inter0, gate43inter1, gate43inter2, gate43inter3, gate43inter4, gate43inter5, gate43inter6, gate43inter7, gate43inter8, gate43inter9, gate43inter10, gate43inter11, gate43inter12, gate11inter0, gate11inter1, gate11inter2, gate11inter3, gate11inter4, gate11inter5, gate11inter6, gate11inter7, gate11inter8, gate11inter9, gate11inter10, gate11inter11, gate11inter12, gate255inter0, gate255inter1, gate255inter2, gate255inter3, gate255inter4, gate255inter5, gate255inter6, gate255inter7, gate255inter8, gate255inter9, gate255inter10, gate255inter11, gate255inter12, gate34inter0, gate34inter1, gate34inter2, gate34inter3, gate34inter4, gate34inter5, gate34inter6, gate34inter7, gate34inter8, gate34inter9, gate34inter10, gate34inter11, gate34inter12, gate106inter0, gate106inter1, gate106inter2, gate106inter3, gate106inter4, gate106inter5, gate106inter6, gate106inter7, gate106inter8, gate106inter9, gate106inter10, gate106inter11, gate106inter12, gate435inter0, gate435inter1, gate435inter2, gate435inter3, gate435inter4, gate435inter5, gate435inter6, gate435inter7, gate435inter8, gate435inter9, gate435inter10, gate435inter11, gate435inter12, gate468inter0, gate468inter1, gate468inter2, gate468inter3, gate468inter4, gate468inter5, gate468inter6, gate468inter7, gate468inter8, gate468inter9, gate468inter10, gate468inter11, gate468inter12, gate81inter0, gate81inter1, gate81inter2, gate81inter3, gate81inter4, gate81inter5, gate81inter6, gate81inter7, gate81inter8, gate81inter9, gate81inter10, gate81inter11, gate81inter12, gate51inter0, gate51inter1, gate51inter2, gate51inter3, gate51inter4, gate51inter5, gate51inter6, gate51inter7, gate51inter8, gate51inter9, gate51inter10, gate51inter11, gate51inter12, gate177inter0, gate177inter1, gate177inter2, gate177inter3, gate177inter4, gate177inter5, gate177inter6, gate177inter7, gate177inter8, gate177inter9, gate177inter10, gate177inter11, gate177inter12, gate488inter0, gate488inter1, gate488inter2, gate488inter3, gate488inter4, gate488inter5, gate488inter6, gate488inter7, gate488inter8, gate488inter9, gate488inter10, gate488inter11, gate488inter12, gate232inter0, gate232inter1, gate232inter2, gate232inter3, gate232inter4, gate232inter5, gate232inter6, gate232inter7, gate232inter8, gate232inter9, gate232inter10, gate232inter11, gate232inter12, gate235inter0, gate235inter1, gate235inter2, gate235inter3, gate235inter4, gate235inter5, gate235inter6, gate235inter7, gate235inter8, gate235inter9, gate235inter10, gate235inter11, gate235inter12, gate234inter0, gate234inter1, gate234inter2, gate234inter3, gate234inter4, gate234inter5, gate234inter6, gate234inter7, gate234inter8, gate234inter9, gate234inter10, gate234inter11, gate234inter12, gate501inter0, gate501inter1, gate501inter2, gate501inter3, gate501inter4, gate501inter5, gate501inter6, gate501inter7, gate501inter8, gate501inter9, gate501inter10, gate501inter11, gate501inter12, gate139inter0, gate139inter1, gate139inter2, gate139inter3, gate139inter4, gate139inter5, gate139inter6, gate139inter7, gate139inter8, gate139inter9, gate139inter10, gate139inter11, gate139inter12, gate242inter0, gate242inter1, gate242inter2, gate242inter3, gate242inter4, gate242inter5, gate242inter6, gate242inter7, gate242inter8, gate242inter9, gate242inter10, gate242inter11, gate242inter12, gate268inter0, gate268inter1, gate268inter2, gate268inter3, gate268inter4, gate268inter5, gate268inter6, gate268inter7, gate268inter8, gate268inter9, gate268inter10, gate268inter11, gate268inter12, gate91inter0, gate91inter1, gate91inter2, gate91inter3, gate91inter4, gate91inter5, gate91inter6, gate91inter7, gate91inter8, gate91inter9, gate91inter10, gate91inter11, gate91inter12, gate175inter0, gate175inter1, gate175inter2, gate175inter3, gate175inter4, gate175inter5, gate175inter6, gate175inter7, gate175inter8, gate175inter9, gate175inter10, gate175inter11, gate175inter12, gate183inter0, gate183inter1, gate183inter2, gate183inter3, gate183inter4, gate183inter5, gate183inter6, gate183inter7, gate183inter8, gate183inter9, gate183inter10, gate183inter11, gate183inter12, gate133inter0, gate133inter1, gate133inter2, gate133inter3, gate133inter4, gate133inter5, gate133inter6, gate133inter7, gate133inter8, gate133inter9, gate133inter10, gate133inter11, gate133inter12;



and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );
nand2 gate9( .a(G1), .b(G2), .O(G266) );
nand2 gate10( .a(G3), .b(G4), .O(G269) );

  xor2  gate1177(.a(G6), .b(G5), .O(gate11inter0));
  nand2 gate1178(.a(gate11inter0), .b(s_90), .O(gate11inter1));
  and2  gate1179(.a(G6), .b(G5), .O(gate11inter2));
  inv1  gate1180(.a(s_90), .O(gate11inter3));
  inv1  gate1181(.a(s_91), .O(gate11inter4));
  nand2 gate1182(.a(gate11inter4), .b(gate11inter3), .O(gate11inter5));
  nor2  gate1183(.a(gate11inter5), .b(gate11inter2), .O(gate11inter6));
  inv1  gate1184(.a(G5), .O(gate11inter7));
  inv1  gate1185(.a(G6), .O(gate11inter8));
  nand2 gate1186(.a(gate11inter8), .b(gate11inter7), .O(gate11inter9));
  nand2 gate1187(.a(s_91), .b(gate11inter3), .O(gate11inter10));
  nor2  gate1188(.a(gate11inter10), .b(gate11inter9), .O(gate11inter11));
  nor2  gate1189(.a(gate11inter11), .b(gate11inter6), .O(gate11inter12));
  nand2 gate1190(.a(gate11inter12), .b(gate11inter1), .O(G272));
nand2 gate12( .a(G7), .b(G8), .O(G275) );
nand2 gate13( .a(G9), .b(G10), .O(G278) );
nand2 gate14( .a(G11), .b(G12), .O(G281) );
nand2 gate15( .a(G13), .b(G14), .O(G284) );
nand2 gate16( .a(G15), .b(G16), .O(G287) );
nand2 gate17( .a(G17), .b(G18), .O(G290) );
nand2 gate18( .a(G19), .b(G20), .O(G293) );
nand2 gate19( .a(G21), .b(G22), .O(G296) );
nand2 gate20( .a(G23), .b(G24), .O(G299) );
nand2 gate21( .a(G25), .b(G26), .O(G302) );
nand2 gate22( .a(G27), .b(G28), .O(G305) );

  xor2  gate967(.a(G30), .b(G29), .O(gate23inter0));
  nand2 gate968(.a(gate23inter0), .b(s_60), .O(gate23inter1));
  and2  gate969(.a(G30), .b(G29), .O(gate23inter2));
  inv1  gate970(.a(s_60), .O(gate23inter3));
  inv1  gate971(.a(s_61), .O(gate23inter4));
  nand2 gate972(.a(gate23inter4), .b(gate23inter3), .O(gate23inter5));
  nor2  gate973(.a(gate23inter5), .b(gate23inter2), .O(gate23inter6));
  inv1  gate974(.a(G29), .O(gate23inter7));
  inv1  gate975(.a(G30), .O(gate23inter8));
  nand2 gate976(.a(gate23inter8), .b(gate23inter7), .O(gate23inter9));
  nand2 gate977(.a(s_61), .b(gate23inter3), .O(gate23inter10));
  nor2  gate978(.a(gate23inter10), .b(gate23inter9), .O(gate23inter11));
  nor2  gate979(.a(gate23inter11), .b(gate23inter6), .O(gate23inter12));
  nand2 gate980(.a(gate23inter12), .b(gate23inter1), .O(G308));

  xor2  gate645(.a(G32), .b(G31), .O(gate24inter0));
  nand2 gate646(.a(gate24inter0), .b(s_14), .O(gate24inter1));
  and2  gate647(.a(G32), .b(G31), .O(gate24inter2));
  inv1  gate648(.a(s_14), .O(gate24inter3));
  inv1  gate649(.a(s_15), .O(gate24inter4));
  nand2 gate650(.a(gate24inter4), .b(gate24inter3), .O(gate24inter5));
  nor2  gate651(.a(gate24inter5), .b(gate24inter2), .O(gate24inter6));
  inv1  gate652(.a(G31), .O(gate24inter7));
  inv1  gate653(.a(G32), .O(gate24inter8));
  nand2 gate654(.a(gate24inter8), .b(gate24inter7), .O(gate24inter9));
  nand2 gate655(.a(s_15), .b(gate24inter3), .O(gate24inter10));
  nor2  gate656(.a(gate24inter10), .b(gate24inter9), .O(gate24inter11));
  nor2  gate657(.a(gate24inter11), .b(gate24inter6), .O(gate24inter12));
  nand2 gate658(.a(gate24inter12), .b(gate24inter1), .O(G311));
nand2 gate25( .a(G1), .b(G5), .O(G314) );
nand2 gate26( .a(G9), .b(G13), .O(G317) );

  xor2  gate981(.a(G6), .b(G2), .O(gate27inter0));
  nand2 gate982(.a(gate27inter0), .b(s_62), .O(gate27inter1));
  and2  gate983(.a(G6), .b(G2), .O(gate27inter2));
  inv1  gate984(.a(s_62), .O(gate27inter3));
  inv1  gate985(.a(s_63), .O(gate27inter4));
  nand2 gate986(.a(gate27inter4), .b(gate27inter3), .O(gate27inter5));
  nor2  gate987(.a(gate27inter5), .b(gate27inter2), .O(gate27inter6));
  inv1  gate988(.a(G2), .O(gate27inter7));
  inv1  gate989(.a(G6), .O(gate27inter8));
  nand2 gate990(.a(gate27inter8), .b(gate27inter7), .O(gate27inter9));
  nand2 gate991(.a(s_63), .b(gate27inter3), .O(gate27inter10));
  nor2  gate992(.a(gate27inter10), .b(gate27inter9), .O(gate27inter11));
  nor2  gate993(.a(gate27inter11), .b(gate27inter6), .O(gate27inter12));
  nand2 gate994(.a(gate27inter12), .b(gate27inter1), .O(G320));
nand2 gate28( .a(G10), .b(G14), .O(G323) );

  xor2  gate575(.a(G7), .b(G3), .O(gate29inter0));
  nand2 gate576(.a(gate29inter0), .b(s_4), .O(gate29inter1));
  and2  gate577(.a(G7), .b(G3), .O(gate29inter2));
  inv1  gate578(.a(s_4), .O(gate29inter3));
  inv1  gate579(.a(s_5), .O(gate29inter4));
  nand2 gate580(.a(gate29inter4), .b(gate29inter3), .O(gate29inter5));
  nor2  gate581(.a(gate29inter5), .b(gate29inter2), .O(gate29inter6));
  inv1  gate582(.a(G3), .O(gate29inter7));
  inv1  gate583(.a(G7), .O(gate29inter8));
  nand2 gate584(.a(gate29inter8), .b(gate29inter7), .O(gate29inter9));
  nand2 gate585(.a(s_5), .b(gate29inter3), .O(gate29inter10));
  nor2  gate586(.a(gate29inter10), .b(gate29inter9), .O(gate29inter11));
  nor2  gate587(.a(gate29inter11), .b(gate29inter6), .O(gate29inter12));
  nand2 gate588(.a(gate29inter12), .b(gate29inter1), .O(G326));
nand2 gate30( .a(G11), .b(G15), .O(G329) );
nand2 gate31( .a(G4), .b(G8), .O(G332) );
nand2 gate32( .a(G12), .b(G16), .O(G335) );
nand2 gate33( .a(G17), .b(G21), .O(G338) );

  xor2  gate1205(.a(G29), .b(G25), .O(gate34inter0));
  nand2 gate1206(.a(gate34inter0), .b(s_94), .O(gate34inter1));
  and2  gate1207(.a(G29), .b(G25), .O(gate34inter2));
  inv1  gate1208(.a(s_94), .O(gate34inter3));
  inv1  gate1209(.a(s_95), .O(gate34inter4));
  nand2 gate1210(.a(gate34inter4), .b(gate34inter3), .O(gate34inter5));
  nor2  gate1211(.a(gate34inter5), .b(gate34inter2), .O(gate34inter6));
  inv1  gate1212(.a(G25), .O(gate34inter7));
  inv1  gate1213(.a(G29), .O(gate34inter8));
  nand2 gate1214(.a(gate34inter8), .b(gate34inter7), .O(gate34inter9));
  nand2 gate1215(.a(s_95), .b(gate34inter3), .O(gate34inter10));
  nor2  gate1216(.a(gate34inter10), .b(gate34inter9), .O(gate34inter11));
  nor2  gate1217(.a(gate34inter11), .b(gate34inter6), .O(gate34inter12));
  nand2 gate1218(.a(gate34inter12), .b(gate34inter1), .O(G341));
nand2 gate35( .a(G18), .b(G22), .O(G344) );
nand2 gate36( .a(G26), .b(G30), .O(G347) );
nand2 gate37( .a(G19), .b(G23), .O(G350) );

  xor2  gate897(.a(G31), .b(G27), .O(gate38inter0));
  nand2 gate898(.a(gate38inter0), .b(s_50), .O(gate38inter1));
  and2  gate899(.a(G31), .b(G27), .O(gate38inter2));
  inv1  gate900(.a(s_50), .O(gate38inter3));
  inv1  gate901(.a(s_51), .O(gate38inter4));
  nand2 gate902(.a(gate38inter4), .b(gate38inter3), .O(gate38inter5));
  nor2  gate903(.a(gate38inter5), .b(gate38inter2), .O(gate38inter6));
  inv1  gate904(.a(G27), .O(gate38inter7));
  inv1  gate905(.a(G31), .O(gate38inter8));
  nand2 gate906(.a(gate38inter8), .b(gate38inter7), .O(gate38inter9));
  nand2 gate907(.a(s_51), .b(gate38inter3), .O(gate38inter10));
  nor2  gate908(.a(gate38inter10), .b(gate38inter9), .O(gate38inter11));
  nor2  gate909(.a(gate38inter11), .b(gate38inter6), .O(gate38inter12));
  nand2 gate910(.a(gate38inter12), .b(gate38inter1), .O(G353));
nand2 gate39( .a(G20), .b(G24), .O(G356) );
nand2 gate40( .a(G28), .b(G32), .O(G359) );
nand2 gate41( .a(G1), .b(G266), .O(G362) );
nand2 gate42( .a(G2), .b(G266), .O(G363) );

  xor2  gate1163(.a(G269), .b(G3), .O(gate43inter0));
  nand2 gate1164(.a(gate43inter0), .b(s_88), .O(gate43inter1));
  and2  gate1165(.a(G269), .b(G3), .O(gate43inter2));
  inv1  gate1166(.a(s_88), .O(gate43inter3));
  inv1  gate1167(.a(s_89), .O(gate43inter4));
  nand2 gate1168(.a(gate43inter4), .b(gate43inter3), .O(gate43inter5));
  nor2  gate1169(.a(gate43inter5), .b(gate43inter2), .O(gate43inter6));
  inv1  gate1170(.a(G3), .O(gate43inter7));
  inv1  gate1171(.a(G269), .O(gate43inter8));
  nand2 gate1172(.a(gate43inter8), .b(gate43inter7), .O(gate43inter9));
  nand2 gate1173(.a(s_89), .b(gate43inter3), .O(gate43inter10));
  nor2  gate1174(.a(gate43inter10), .b(gate43inter9), .O(gate43inter11));
  nor2  gate1175(.a(gate43inter11), .b(gate43inter6), .O(gate43inter12));
  nand2 gate1176(.a(gate43inter12), .b(gate43inter1), .O(G364));
nand2 gate44( .a(G4), .b(G269), .O(G365) );
nand2 gate45( .a(G5), .b(G272), .O(G366) );
nand2 gate46( .a(G6), .b(G272), .O(G367) );
nand2 gate47( .a(G7), .b(G275), .O(G368) );
nand2 gate48( .a(G8), .b(G275), .O(G369) );
nand2 gate49( .a(G9), .b(G278), .O(G370) );
nand2 gate50( .a(G10), .b(G278), .O(G371) );

  xor2  gate1275(.a(G281), .b(G11), .O(gate51inter0));
  nand2 gate1276(.a(gate51inter0), .b(s_104), .O(gate51inter1));
  and2  gate1277(.a(G281), .b(G11), .O(gate51inter2));
  inv1  gate1278(.a(s_104), .O(gate51inter3));
  inv1  gate1279(.a(s_105), .O(gate51inter4));
  nand2 gate1280(.a(gate51inter4), .b(gate51inter3), .O(gate51inter5));
  nor2  gate1281(.a(gate51inter5), .b(gate51inter2), .O(gate51inter6));
  inv1  gate1282(.a(G11), .O(gate51inter7));
  inv1  gate1283(.a(G281), .O(gate51inter8));
  nand2 gate1284(.a(gate51inter8), .b(gate51inter7), .O(gate51inter9));
  nand2 gate1285(.a(s_105), .b(gate51inter3), .O(gate51inter10));
  nor2  gate1286(.a(gate51inter10), .b(gate51inter9), .O(gate51inter11));
  nor2  gate1287(.a(gate51inter11), .b(gate51inter6), .O(gate51inter12));
  nand2 gate1288(.a(gate51inter12), .b(gate51inter1), .O(G372));
nand2 gate52( .a(G12), .b(G281), .O(G373) );

  xor2  gate1093(.a(G284), .b(G13), .O(gate53inter0));
  nand2 gate1094(.a(gate53inter0), .b(s_78), .O(gate53inter1));
  and2  gate1095(.a(G284), .b(G13), .O(gate53inter2));
  inv1  gate1096(.a(s_78), .O(gate53inter3));
  inv1  gate1097(.a(s_79), .O(gate53inter4));
  nand2 gate1098(.a(gate53inter4), .b(gate53inter3), .O(gate53inter5));
  nor2  gate1099(.a(gate53inter5), .b(gate53inter2), .O(gate53inter6));
  inv1  gate1100(.a(G13), .O(gate53inter7));
  inv1  gate1101(.a(G284), .O(gate53inter8));
  nand2 gate1102(.a(gate53inter8), .b(gate53inter7), .O(gate53inter9));
  nand2 gate1103(.a(s_79), .b(gate53inter3), .O(gate53inter10));
  nor2  gate1104(.a(gate53inter10), .b(gate53inter9), .O(gate53inter11));
  nor2  gate1105(.a(gate53inter11), .b(gate53inter6), .O(gate53inter12));
  nand2 gate1106(.a(gate53inter12), .b(gate53inter1), .O(G374));
nand2 gate54( .a(G14), .b(G284), .O(G375) );
nand2 gate55( .a(G15), .b(G287), .O(G376) );
nand2 gate56( .a(G16), .b(G287), .O(G377) );
nand2 gate57( .a(G17), .b(G290), .O(G378) );
nand2 gate58( .a(G18), .b(G290), .O(G379) );
nand2 gate59( .a(G19), .b(G293), .O(G380) );
nand2 gate60( .a(G20), .b(G293), .O(G381) );
nand2 gate61( .a(G21), .b(G296), .O(G382) );
nand2 gate62( .a(G22), .b(G296), .O(G383) );
nand2 gate63( .a(G23), .b(G299), .O(G384) );
nand2 gate64( .a(G24), .b(G299), .O(G385) );
nand2 gate65( .a(G25), .b(G302), .O(G386) );

  xor2  gate1149(.a(G302), .b(G26), .O(gate66inter0));
  nand2 gate1150(.a(gate66inter0), .b(s_86), .O(gate66inter1));
  and2  gate1151(.a(G302), .b(G26), .O(gate66inter2));
  inv1  gate1152(.a(s_86), .O(gate66inter3));
  inv1  gate1153(.a(s_87), .O(gate66inter4));
  nand2 gate1154(.a(gate66inter4), .b(gate66inter3), .O(gate66inter5));
  nor2  gate1155(.a(gate66inter5), .b(gate66inter2), .O(gate66inter6));
  inv1  gate1156(.a(G26), .O(gate66inter7));
  inv1  gate1157(.a(G302), .O(gate66inter8));
  nand2 gate1158(.a(gate66inter8), .b(gate66inter7), .O(gate66inter9));
  nand2 gate1159(.a(s_87), .b(gate66inter3), .O(gate66inter10));
  nor2  gate1160(.a(gate66inter10), .b(gate66inter9), .O(gate66inter11));
  nor2  gate1161(.a(gate66inter11), .b(gate66inter6), .O(gate66inter12));
  nand2 gate1162(.a(gate66inter12), .b(gate66inter1), .O(G387));
nand2 gate67( .a(G27), .b(G305), .O(G388) );
nand2 gate68( .a(G28), .b(G305), .O(G389) );
nand2 gate69( .a(G29), .b(G308), .O(G390) );
nand2 gate70( .a(G30), .b(G308), .O(G391) );
nand2 gate71( .a(G31), .b(G311), .O(G392) );
nand2 gate72( .a(G32), .b(G311), .O(G393) );
nand2 gate73( .a(G1), .b(G314), .O(G394) );
nand2 gate74( .a(G5), .b(G314), .O(G395) );
nand2 gate75( .a(G9), .b(G317), .O(G396) );
nand2 gate76( .a(G13), .b(G317), .O(G397) );
nand2 gate77( .a(G2), .b(G320), .O(G398) );
nand2 gate78( .a(G6), .b(G320), .O(G399) );
nand2 gate79( .a(G10), .b(G323), .O(G400) );
nand2 gate80( .a(G14), .b(G323), .O(G401) );

  xor2  gate1261(.a(G326), .b(G3), .O(gate81inter0));
  nand2 gate1262(.a(gate81inter0), .b(s_102), .O(gate81inter1));
  and2  gate1263(.a(G326), .b(G3), .O(gate81inter2));
  inv1  gate1264(.a(s_102), .O(gate81inter3));
  inv1  gate1265(.a(s_103), .O(gate81inter4));
  nand2 gate1266(.a(gate81inter4), .b(gate81inter3), .O(gate81inter5));
  nor2  gate1267(.a(gate81inter5), .b(gate81inter2), .O(gate81inter6));
  inv1  gate1268(.a(G3), .O(gate81inter7));
  inv1  gate1269(.a(G326), .O(gate81inter8));
  nand2 gate1270(.a(gate81inter8), .b(gate81inter7), .O(gate81inter9));
  nand2 gate1271(.a(s_103), .b(gate81inter3), .O(gate81inter10));
  nor2  gate1272(.a(gate81inter10), .b(gate81inter9), .O(gate81inter11));
  nor2  gate1273(.a(gate81inter11), .b(gate81inter6), .O(gate81inter12));
  nand2 gate1274(.a(gate81inter12), .b(gate81inter1), .O(G402));
nand2 gate82( .a(G7), .b(G326), .O(G403) );
nand2 gate83( .a(G11), .b(G329), .O(G404) );

  xor2  gate841(.a(G329), .b(G15), .O(gate84inter0));
  nand2 gate842(.a(gate84inter0), .b(s_42), .O(gate84inter1));
  and2  gate843(.a(G329), .b(G15), .O(gate84inter2));
  inv1  gate844(.a(s_42), .O(gate84inter3));
  inv1  gate845(.a(s_43), .O(gate84inter4));
  nand2 gate846(.a(gate84inter4), .b(gate84inter3), .O(gate84inter5));
  nor2  gate847(.a(gate84inter5), .b(gate84inter2), .O(gate84inter6));
  inv1  gate848(.a(G15), .O(gate84inter7));
  inv1  gate849(.a(G329), .O(gate84inter8));
  nand2 gate850(.a(gate84inter8), .b(gate84inter7), .O(gate84inter9));
  nand2 gate851(.a(s_43), .b(gate84inter3), .O(gate84inter10));
  nor2  gate852(.a(gate84inter10), .b(gate84inter9), .O(gate84inter11));
  nor2  gate853(.a(gate84inter11), .b(gate84inter6), .O(gate84inter12));
  nand2 gate854(.a(gate84inter12), .b(gate84inter1), .O(G405));
nand2 gate85( .a(G4), .b(G332), .O(G406) );
nand2 gate86( .a(G8), .b(G332), .O(G407) );
nand2 gate87( .a(G12), .b(G335), .O(G408) );
nand2 gate88( .a(G16), .b(G335), .O(G409) );
nand2 gate89( .a(G17), .b(G338), .O(G410) );
nand2 gate90( .a(G21), .b(G338), .O(G411) );

  xor2  gate1415(.a(G341), .b(G25), .O(gate91inter0));
  nand2 gate1416(.a(gate91inter0), .b(s_124), .O(gate91inter1));
  and2  gate1417(.a(G341), .b(G25), .O(gate91inter2));
  inv1  gate1418(.a(s_124), .O(gate91inter3));
  inv1  gate1419(.a(s_125), .O(gate91inter4));
  nand2 gate1420(.a(gate91inter4), .b(gate91inter3), .O(gate91inter5));
  nor2  gate1421(.a(gate91inter5), .b(gate91inter2), .O(gate91inter6));
  inv1  gate1422(.a(G25), .O(gate91inter7));
  inv1  gate1423(.a(G341), .O(gate91inter8));
  nand2 gate1424(.a(gate91inter8), .b(gate91inter7), .O(gate91inter9));
  nand2 gate1425(.a(s_125), .b(gate91inter3), .O(gate91inter10));
  nor2  gate1426(.a(gate91inter10), .b(gate91inter9), .O(gate91inter11));
  nor2  gate1427(.a(gate91inter11), .b(gate91inter6), .O(gate91inter12));
  nand2 gate1428(.a(gate91inter12), .b(gate91inter1), .O(G412));
nand2 gate92( .a(G29), .b(G341), .O(G413) );
nand2 gate93( .a(G18), .b(G344), .O(G414) );
nand2 gate94( .a(G22), .b(G344), .O(G415) );

  xor2  gate1037(.a(G347), .b(G26), .O(gate95inter0));
  nand2 gate1038(.a(gate95inter0), .b(s_70), .O(gate95inter1));
  and2  gate1039(.a(G347), .b(G26), .O(gate95inter2));
  inv1  gate1040(.a(s_70), .O(gate95inter3));
  inv1  gate1041(.a(s_71), .O(gate95inter4));
  nand2 gate1042(.a(gate95inter4), .b(gate95inter3), .O(gate95inter5));
  nor2  gate1043(.a(gate95inter5), .b(gate95inter2), .O(gate95inter6));
  inv1  gate1044(.a(G26), .O(gate95inter7));
  inv1  gate1045(.a(G347), .O(gate95inter8));
  nand2 gate1046(.a(gate95inter8), .b(gate95inter7), .O(gate95inter9));
  nand2 gate1047(.a(s_71), .b(gate95inter3), .O(gate95inter10));
  nor2  gate1048(.a(gate95inter10), .b(gate95inter9), .O(gate95inter11));
  nor2  gate1049(.a(gate95inter11), .b(gate95inter6), .O(gate95inter12));
  nand2 gate1050(.a(gate95inter12), .b(gate95inter1), .O(G416));
nand2 gate96( .a(G30), .b(G347), .O(G417) );
nand2 gate97( .a(G19), .b(G350), .O(G418) );

  xor2  gate995(.a(G350), .b(G23), .O(gate98inter0));
  nand2 gate996(.a(gate98inter0), .b(s_64), .O(gate98inter1));
  and2  gate997(.a(G350), .b(G23), .O(gate98inter2));
  inv1  gate998(.a(s_64), .O(gate98inter3));
  inv1  gate999(.a(s_65), .O(gate98inter4));
  nand2 gate1000(.a(gate98inter4), .b(gate98inter3), .O(gate98inter5));
  nor2  gate1001(.a(gate98inter5), .b(gate98inter2), .O(gate98inter6));
  inv1  gate1002(.a(G23), .O(gate98inter7));
  inv1  gate1003(.a(G350), .O(gate98inter8));
  nand2 gate1004(.a(gate98inter8), .b(gate98inter7), .O(gate98inter9));
  nand2 gate1005(.a(s_65), .b(gate98inter3), .O(gate98inter10));
  nor2  gate1006(.a(gate98inter10), .b(gate98inter9), .O(gate98inter11));
  nor2  gate1007(.a(gate98inter11), .b(gate98inter6), .O(gate98inter12));
  nand2 gate1008(.a(gate98inter12), .b(gate98inter1), .O(G419));
nand2 gate99( .a(G27), .b(G353), .O(G420) );
nand2 gate100( .a(G31), .b(G353), .O(G421) );
nand2 gate101( .a(G20), .b(G356), .O(G422) );
nand2 gate102( .a(G24), .b(G356), .O(G423) );
nand2 gate103( .a(G28), .b(G359), .O(G424) );
nand2 gate104( .a(G32), .b(G359), .O(G425) );
nand2 gate105( .a(G362), .b(G363), .O(G426) );

  xor2  gate1219(.a(G365), .b(G364), .O(gate106inter0));
  nand2 gate1220(.a(gate106inter0), .b(s_96), .O(gate106inter1));
  and2  gate1221(.a(G365), .b(G364), .O(gate106inter2));
  inv1  gate1222(.a(s_96), .O(gate106inter3));
  inv1  gate1223(.a(s_97), .O(gate106inter4));
  nand2 gate1224(.a(gate106inter4), .b(gate106inter3), .O(gate106inter5));
  nor2  gate1225(.a(gate106inter5), .b(gate106inter2), .O(gate106inter6));
  inv1  gate1226(.a(G364), .O(gate106inter7));
  inv1  gate1227(.a(G365), .O(gate106inter8));
  nand2 gate1228(.a(gate106inter8), .b(gate106inter7), .O(gate106inter9));
  nand2 gate1229(.a(s_97), .b(gate106inter3), .O(gate106inter10));
  nor2  gate1230(.a(gate106inter10), .b(gate106inter9), .O(gate106inter11));
  nor2  gate1231(.a(gate106inter11), .b(gate106inter6), .O(gate106inter12));
  nand2 gate1232(.a(gate106inter12), .b(gate106inter1), .O(G429));

  xor2  gate1079(.a(G367), .b(G366), .O(gate107inter0));
  nand2 gate1080(.a(gate107inter0), .b(s_76), .O(gate107inter1));
  and2  gate1081(.a(G367), .b(G366), .O(gate107inter2));
  inv1  gate1082(.a(s_76), .O(gate107inter3));
  inv1  gate1083(.a(s_77), .O(gate107inter4));
  nand2 gate1084(.a(gate107inter4), .b(gate107inter3), .O(gate107inter5));
  nor2  gate1085(.a(gate107inter5), .b(gate107inter2), .O(gate107inter6));
  inv1  gate1086(.a(G366), .O(gate107inter7));
  inv1  gate1087(.a(G367), .O(gate107inter8));
  nand2 gate1088(.a(gate107inter8), .b(gate107inter7), .O(gate107inter9));
  nand2 gate1089(.a(s_77), .b(gate107inter3), .O(gate107inter10));
  nor2  gate1090(.a(gate107inter10), .b(gate107inter9), .O(gate107inter11));
  nor2  gate1091(.a(gate107inter11), .b(gate107inter6), .O(gate107inter12));
  nand2 gate1092(.a(gate107inter12), .b(gate107inter1), .O(G432));
nand2 gate108( .a(G368), .b(G369), .O(G435) );
nand2 gate109( .a(G370), .b(G371), .O(G438) );

  xor2  gate743(.a(G373), .b(G372), .O(gate110inter0));
  nand2 gate744(.a(gate110inter0), .b(s_28), .O(gate110inter1));
  and2  gate745(.a(G373), .b(G372), .O(gate110inter2));
  inv1  gate746(.a(s_28), .O(gate110inter3));
  inv1  gate747(.a(s_29), .O(gate110inter4));
  nand2 gate748(.a(gate110inter4), .b(gate110inter3), .O(gate110inter5));
  nor2  gate749(.a(gate110inter5), .b(gate110inter2), .O(gate110inter6));
  inv1  gate750(.a(G372), .O(gate110inter7));
  inv1  gate751(.a(G373), .O(gate110inter8));
  nand2 gate752(.a(gate110inter8), .b(gate110inter7), .O(gate110inter9));
  nand2 gate753(.a(s_29), .b(gate110inter3), .O(gate110inter10));
  nor2  gate754(.a(gate110inter10), .b(gate110inter9), .O(gate110inter11));
  nor2  gate755(.a(gate110inter11), .b(gate110inter6), .O(gate110inter12));
  nand2 gate756(.a(gate110inter12), .b(gate110inter1), .O(G441));

  xor2  gate827(.a(G375), .b(G374), .O(gate111inter0));
  nand2 gate828(.a(gate111inter0), .b(s_40), .O(gate111inter1));
  and2  gate829(.a(G375), .b(G374), .O(gate111inter2));
  inv1  gate830(.a(s_40), .O(gate111inter3));
  inv1  gate831(.a(s_41), .O(gate111inter4));
  nand2 gate832(.a(gate111inter4), .b(gate111inter3), .O(gate111inter5));
  nor2  gate833(.a(gate111inter5), .b(gate111inter2), .O(gate111inter6));
  inv1  gate834(.a(G374), .O(gate111inter7));
  inv1  gate835(.a(G375), .O(gate111inter8));
  nand2 gate836(.a(gate111inter8), .b(gate111inter7), .O(gate111inter9));
  nand2 gate837(.a(s_41), .b(gate111inter3), .O(gate111inter10));
  nor2  gate838(.a(gate111inter10), .b(gate111inter9), .O(gate111inter11));
  nor2  gate839(.a(gate111inter11), .b(gate111inter6), .O(gate111inter12));
  nand2 gate840(.a(gate111inter12), .b(gate111inter1), .O(G444));
nand2 gate112( .a(G376), .b(G377), .O(G447) );
nand2 gate113( .a(G378), .b(G379), .O(G450) );
nand2 gate114( .a(G380), .b(G381), .O(G453) );

  xor2  gate603(.a(G383), .b(G382), .O(gate115inter0));
  nand2 gate604(.a(gate115inter0), .b(s_8), .O(gate115inter1));
  and2  gate605(.a(G383), .b(G382), .O(gate115inter2));
  inv1  gate606(.a(s_8), .O(gate115inter3));
  inv1  gate607(.a(s_9), .O(gate115inter4));
  nand2 gate608(.a(gate115inter4), .b(gate115inter3), .O(gate115inter5));
  nor2  gate609(.a(gate115inter5), .b(gate115inter2), .O(gate115inter6));
  inv1  gate610(.a(G382), .O(gate115inter7));
  inv1  gate611(.a(G383), .O(gate115inter8));
  nand2 gate612(.a(gate115inter8), .b(gate115inter7), .O(gate115inter9));
  nand2 gate613(.a(s_9), .b(gate115inter3), .O(gate115inter10));
  nor2  gate614(.a(gate115inter10), .b(gate115inter9), .O(gate115inter11));
  nor2  gate615(.a(gate115inter11), .b(gate115inter6), .O(gate115inter12));
  nand2 gate616(.a(gate115inter12), .b(gate115inter1), .O(G456));
nand2 gate116( .a(G384), .b(G385), .O(G459) );
nand2 gate117( .a(G386), .b(G387), .O(G462) );
nand2 gate118( .a(G388), .b(G389), .O(G465) );
nand2 gate119( .a(G390), .b(G391), .O(G468) );
nand2 gate120( .a(G392), .b(G393), .O(G471) );
nand2 gate121( .a(G394), .b(G395), .O(G474) );
nand2 gate122( .a(G396), .b(G397), .O(G477) );
nand2 gate123( .a(G398), .b(G399), .O(G480) );
nand2 gate124( .a(G400), .b(G401), .O(G483) );
nand2 gate125( .a(G402), .b(G403), .O(G486) );
nand2 gate126( .a(G404), .b(G405), .O(G489) );
nand2 gate127( .a(G406), .b(G407), .O(G492) );
nand2 gate128( .a(G408), .b(G409), .O(G495) );
nand2 gate129( .a(G410), .b(G411), .O(G498) );
nand2 gate130( .a(G412), .b(G413), .O(G501) );

  xor2  gate799(.a(G415), .b(G414), .O(gate131inter0));
  nand2 gate800(.a(gate131inter0), .b(s_36), .O(gate131inter1));
  and2  gate801(.a(G415), .b(G414), .O(gate131inter2));
  inv1  gate802(.a(s_36), .O(gate131inter3));
  inv1  gate803(.a(s_37), .O(gate131inter4));
  nand2 gate804(.a(gate131inter4), .b(gate131inter3), .O(gate131inter5));
  nor2  gate805(.a(gate131inter5), .b(gate131inter2), .O(gate131inter6));
  inv1  gate806(.a(G414), .O(gate131inter7));
  inv1  gate807(.a(G415), .O(gate131inter8));
  nand2 gate808(.a(gate131inter8), .b(gate131inter7), .O(gate131inter9));
  nand2 gate809(.a(s_37), .b(gate131inter3), .O(gate131inter10));
  nor2  gate810(.a(gate131inter10), .b(gate131inter9), .O(gate131inter11));
  nor2  gate811(.a(gate131inter11), .b(gate131inter6), .O(gate131inter12));
  nand2 gate812(.a(gate131inter12), .b(gate131inter1), .O(G504));

  xor2  gate1065(.a(G417), .b(G416), .O(gate132inter0));
  nand2 gate1066(.a(gate132inter0), .b(s_74), .O(gate132inter1));
  and2  gate1067(.a(G417), .b(G416), .O(gate132inter2));
  inv1  gate1068(.a(s_74), .O(gate132inter3));
  inv1  gate1069(.a(s_75), .O(gate132inter4));
  nand2 gate1070(.a(gate132inter4), .b(gate132inter3), .O(gate132inter5));
  nor2  gate1071(.a(gate132inter5), .b(gate132inter2), .O(gate132inter6));
  inv1  gate1072(.a(G416), .O(gate132inter7));
  inv1  gate1073(.a(G417), .O(gate132inter8));
  nand2 gate1074(.a(gate132inter8), .b(gate132inter7), .O(gate132inter9));
  nand2 gate1075(.a(s_75), .b(gate132inter3), .O(gate132inter10));
  nor2  gate1076(.a(gate132inter10), .b(gate132inter9), .O(gate132inter11));
  nor2  gate1077(.a(gate132inter11), .b(gate132inter6), .O(gate132inter12));
  nand2 gate1078(.a(gate132inter12), .b(gate132inter1), .O(G507));

  xor2  gate1457(.a(G419), .b(G418), .O(gate133inter0));
  nand2 gate1458(.a(gate133inter0), .b(s_130), .O(gate133inter1));
  and2  gate1459(.a(G419), .b(G418), .O(gate133inter2));
  inv1  gate1460(.a(s_130), .O(gate133inter3));
  inv1  gate1461(.a(s_131), .O(gate133inter4));
  nand2 gate1462(.a(gate133inter4), .b(gate133inter3), .O(gate133inter5));
  nor2  gate1463(.a(gate133inter5), .b(gate133inter2), .O(gate133inter6));
  inv1  gate1464(.a(G418), .O(gate133inter7));
  inv1  gate1465(.a(G419), .O(gate133inter8));
  nand2 gate1466(.a(gate133inter8), .b(gate133inter7), .O(gate133inter9));
  nand2 gate1467(.a(s_131), .b(gate133inter3), .O(gate133inter10));
  nor2  gate1468(.a(gate133inter10), .b(gate133inter9), .O(gate133inter11));
  nor2  gate1469(.a(gate133inter11), .b(gate133inter6), .O(gate133inter12));
  nand2 gate1470(.a(gate133inter12), .b(gate133inter1), .O(G510));
nand2 gate134( .a(G420), .b(G421), .O(G513) );
nand2 gate135( .a(G422), .b(G423), .O(G516) );
nand2 gate136( .a(G424), .b(G425), .O(G519) );
nand2 gate137( .a(G426), .b(G429), .O(G522) );
nand2 gate138( .a(G432), .b(G435), .O(G525) );

  xor2  gate1373(.a(G441), .b(G438), .O(gate139inter0));
  nand2 gate1374(.a(gate139inter0), .b(s_118), .O(gate139inter1));
  and2  gate1375(.a(G441), .b(G438), .O(gate139inter2));
  inv1  gate1376(.a(s_118), .O(gate139inter3));
  inv1  gate1377(.a(s_119), .O(gate139inter4));
  nand2 gate1378(.a(gate139inter4), .b(gate139inter3), .O(gate139inter5));
  nor2  gate1379(.a(gate139inter5), .b(gate139inter2), .O(gate139inter6));
  inv1  gate1380(.a(G438), .O(gate139inter7));
  inv1  gate1381(.a(G441), .O(gate139inter8));
  nand2 gate1382(.a(gate139inter8), .b(gate139inter7), .O(gate139inter9));
  nand2 gate1383(.a(s_119), .b(gate139inter3), .O(gate139inter10));
  nor2  gate1384(.a(gate139inter10), .b(gate139inter9), .O(gate139inter11));
  nor2  gate1385(.a(gate139inter11), .b(gate139inter6), .O(gate139inter12));
  nand2 gate1386(.a(gate139inter12), .b(gate139inter1), .O(G528));
nand2 gate140( .a(G444), .b(G447), .O(G531) );

  xor2  gate687(.a(G453), .b(G450), .O(gate141inter0));
  nand2 gate688(.a(gate141inter0), .b(s_20), .O(gate141inter1));
  and2  gate689(.a(G453), .b(G450), .O(gate141inter2));
  inv1  gate690(.a(s_20), .O(gate141inter3));
  inv1  gate691(.a(s_21), .O(gate141inter4));
  nand2 gate692(.a(gate141inter4), .b(gate141inter3), .O(gate141inter5));
  nor2  gate693(.a(gate141inter5), .b(gate141inter2), .O(gate141inter6));
  inv1  gate694(.a(G450), .O(gate141inter7));
  inv1  gate695(.a(G453), .O(gate141inter8));
  nand2 gate696(.a(gate141inter8), .b(gate141inter7), .O(gate141inter9));
  nand2 gate697(.a(s_21), .b(gate141inter3), .O(gate141inter10));
  nor2  gate698(.a(gate141inter10), .b(gate141inter9), .O(gate141inter11));
  nor2  gate699(.a(gate141inter11), .b(gate141inter6), .O(gate141inter12));
  nand2 gate700(.a(gate141inter12), .b(gate141inter1), .O(G534));
nand2 gate142( .a(G456), .b(G459), .O(G537) );
nand2 gate143( .a(G462), .b(G465), .O(G540) );
nand2 gate144( .a(G468), .b(G471), .O(G543) );
nand2 gate145( .a(G474), .b(G477), .O(G546) );
nand2 gate146( .a(G480), .b(G483), .O(G549) );
nand2 gate147( .a(G486), .b(G489), .O(G552) );
nand2 gate148( .a(G492), .b(G495), .O(G555) );
nand2 gate149( .a(G498), .b(G501), .O(G558) );
nand2 gate150( .a(G504), .b(G507), .O(G561) );
nand2 gate151( .a(G510), .b(G513), .O(G564) );
nand2 gate152( .a(G516), .b(G519), .O(G567) );
nand2 gate153( .a(G426), .b(G522), .O(G570) );

  xor2  gate869(.a(G522), .b(G429), .O(gate154inter0));
  nand2 gate870(.a(gate154inter0), .b(s_46), .O(gate154inter1));
  and2  gate871(.a(G522), .b(G429), .O(gate154inter2));
  inv1  gate872(.a(s_46), .O(gate154inter3));
  inv1  gate873(.a(s_47), .O(gate154inter4));
  nand2 gate874(.a(gate154inter4), .b(gate154inter3), .O(gate154inter5));
  nor2  gate875(.a(gate154inter5), .b(gate154inter2), .O(gate154inter6));
  inv1  gate876(.a(G429), .O(gate154inter7));
  inv1  gate877(.a(G522), .O(gate154inter8));
  nand2 gate878(.a(gate154inter8), .b(gate154inter7), .O(gate154inter9));
  nand2 gate879(.a(s_47), .b(gate154inter3), .O(gate154inter10));
  nor2  gate880(.a(gate154inter10), .b(gate154inter9), .O(gate154inter11));
  nor2  gate881(.a(gate154inter11), .b(gate154inter6), .O(gate154inter12));
  nand2 gate882(.a(gate154inter12), .b(gate154inter1), .O(G571));
nand2 gate155( .a(G432), .b(G525), .O(G572) );
nand2 gate156( .a(G435), .b(G525), .O(G573) );
nand2 gate157( .a(G438), .b(G528), .O(G574) );
nand2 gate158( .a(G441), .b(G528), .O(G575) );
nand2 gate159( .a(G444), .b(G531), .O(G576) );
nand2 gate160( .a(G447), .b(G531), .O(G577) );
nand2 gate161( .a(G450), .b(G534), .O(G578) );
nand2 gate162( .a(G453), .b(G534), .O(G579) );
nand2 gate163( .a(G456), .b(G537), .O(G580) );
nand2 gate164( .a(G459), .b(G537), .O(G581) );
nand2 gate165( .a(G462), .b(G540), .O(G582) );
nand2 gate166( .a(G465), .b(G540), .O(G583) );
nand2 gate167( .a(G468), .b(G543), .O(G584) );
nand2 gate168( .a(G471), .b(G543), .O(G585) );
nand2 gate169( .a(G474), .b(G546), .O(G586) );

  xor2  gate1135(.a(G546), .b(G477), .O(gate170inter0));
  nand2 gate1136(.a(gate170inter0), .b(s_84), .O(gate170inter1));
  and2  gate1137(.a(G546), .b(G477), .O(gate170inter2));
  inv1  gate1138(.a(s_84), .O(gate170inter3));
  inv1  gate1139(.a(s_85), .O(gate170inter4));
  nand2 gate1140(.a(gate170inter4), .b(gate170inter3), .O(gate170inter5));
  nor2  gate1141(.a(gate170inter5), .b(gate170inter2), .O(gate170inter6));
  inv1  gate1142(.a(G477), .O(gate170inter7));
  inv1  gate1143(.a(G546), .O(gate170inter8));
  nand2 gate1144(.a(gate170inter8), .b(gate170inter7), .O(gate170inter9));
  nand2 gate1145(.a(s_85), .b(gate170inter3), .O(gate170inter10));
  nor2  gate1146(.a(gate170inter10), .b(gate170inter9), .O(gate170inter11));
  nor2  gate1147(.a(gate170inter11), .b(gate170inter6), .O(gate170inter12));
  nand2 gate1148(.a(gate170inter12), .b(gate170inter1), .O(G587));
nand2 gate171( .a(G480), .b(G549), .O(G588) );
nand2 gate172( .a(G483), .b(G549), .O(G589) );
nand2 gate173( .a(G486), .b(G552), .O(G590) );
nand2 gate174( .a(G489), .b(G552), .O(G591) );

  xor2  gate1429(.a(G555), .b(G492), .O(gate175inter0));
  nand2 gate1430(.a(gate175inter0), .b(s_126), .O(gate175inter1));
  and2  gate1431(.a(G555), .b(G492), .O(gate175inter2));
  inv1  gate1432(.a(s_126), .O(gate175inter3));
  inv1  gate1433(.a(s_127), .O(gate175inter4));
  nand2 gate1434(.a(gate175inter4), .b(gate175inter3), .O(gate175inter5));
  nor2  gate1435(.a(gate175inter5), .b(gate175inter2), .O(gate175inter6));
  inv1  gate1436(.a(G492), .O(gate175inter7));
  inv1  gate1437(.a(G555), .O(gate175inter8));
  nand2 gate1438(.a(gate175inter8), .b(gate175inter7), .O(gate175inter9));
  nand2 gate1439(.a(s_127), .b(gate175inter3), .O(gate175inter10));
  nor2  gate1440(.a(gate175inter10), .b(gate175inter9), .O(gate175inter11));
  nor2  gate1441(.a(gate175inter11), .b(gate175inter6), .O(gate175inter12));
  nand2 gate1442(.a(gate175inter12), .b(gate175inter1), .O(G592));
nand2 gate176( .a(G495), .b(G555), .O(G593) );

  xor2  gate1289(.a(G558), .b(G498), .O(gate177inter0));
  nand2 gate1290(.a(gate177inter0), .b(s_106), .O(gate177inter1));
  and2  gate1291(.a(G558), .b(G498), .O(gate177inter2));
  inv1  gate1292(.a(s_106), .O(gate177inter3));
  inv1  gate1293(.a(s_107), .O(gate177inter4));
  nand2 gate1294(.a(gate177inter4), .b(gate177inter3), .O(gate177inter5));
  nor2  gate1295(.a(gate177inter5), .b(gate177inter2), .O(gate177inter6));
  inv1  gate1296(.a(G498), .O(gate177inter7));
  inv1  gate1297(.a(G558), .O(gate177inter8));
  nand2 gate1298(.a(gate177inter8), .b(gate177inter7), .O(gate177inter9));
  nand2 gate1299(.a(s_107), .b(gate177inter3), .O(gate177inter10));
  nor2  gate1300(.a(gate177inter10), .b(gate177inter9), .O(gate177inter11));
  nor2  gate1301(.a(gate177inter11), .b(gate177inter6), .O(gate177inter12));
  nand2 gate1302(.a(gate177inter12), .b(gate177inter1), .O(G594));
nand2 gate178( .a(G501), .b(G558), .O(G595) );
nand2 gate179( .a(G504), .b(G561), .O(G596) );

  xor2  gate1107(.a(G561), .b(G507), .O(gate180inter0));
  nand2 gate1108(.a(gate180inter0), .b(s_80), .O(gate180inter1));
  and2  gate1109(.a(G561), .b(G507), .O(gate180inter2));
  inv1  gate1110(.a(s_80), .O(gate180inter3));
  inv1  gate1111(.a(s_81), .O(gate180inter4));
  nand2 gate1112(.a(gate180inter4), .b(gate180inter3), .O(gate180inter5));
  nor2  gate1113(.a(gate180inter5), .b(gate180inter2), .O(gate180inter6));
  inv1  gate1114(.a(G507), .O(gate180inter7));
  inv1  gate1115(.a(G561), .O(gate180inter8));
  nand2 gate1116(.a(gate180inter8), .b(gate180inter7), .O(gate180inter9));
  nand2 gate1117(.a(s_81), .b(gate180inter3), .O(gate180inter10));
  nor2  gate1118(.a(gate180inter10), .b(gate180inter9), .O(gate180inter11));
  nor2  gate1119(.a(gate180inter11), .b(gate180inter6), .O(gate180inter12));
  nand2 gate1120(.a(gate180inter12), .b(gate180inter1), .O(G597));
nand2 gate181( .a(G510), .b(G564), .O(G598) );
nand2 gate182( .a(G513), .b(G564), .O(G599) );

  xor2  gate1443(.a(G567), .b(G516), .O(gate183inter0));
  nand2 gate1444(.a(gate183inter0), .b(s_128), .O(gate183inter1));
  and2  gate1445(.a(G567), .b(G516), .O(gate183inter2));
  inv1  gate1446(.a(s_128), .O(gate183inter3));
  inv1  gate1447(.a(s_129), .O(gate183inter4));
  nand2 gate1448(.a(gate183inter4), .b(gate183inter3), .O(gate183inter5));
  nor2  gate1449(.a(gate183inter5), .b(gate183inter2), .O(gate183inter6));
  inv1  gate1450(.a(G516), .O(gate183inter7));
  inv1  gate1451(.a(G567), .O(gate183inter8));
  nand2 gate1452(.a(gate183inter8), .b(gate183inter7), .O(gate183inter9));
  nand2 gate1453(.a(s_129), .b(gate183inter3), .O(gate183inter10));
  nor2  gate1454(.a(gate183inter10), .b(gate183inter9), .O(gate183inter11));
  nor2  gate1455(.a(gate183inter11), .b(gate183inter6), .O(gate183inter12));
  nand2 gate1456(.a(gate183inter12), .b(gate183inter1), .O(G600));
nand2 gate184( .a(G519), .b(G567), .O(G601) );
nand2 gate185( .a(G570), .b(G571), .O(G602) );
nand2 gate186( .a(G572), .b(G573), .O(G607) );

  xor2  gate855(.a(G575), .b(G574), .O(gate187inter0));
  nand2 gate856(.a(gate187inter0), .b(s_44), .O(gate187inter1));
  and2  gate857(.a(G575), .b(G574), .O(gate187inter2));
  inv1  gate858(.a(s_44), .O(gate187inter3));
  inv1  gate859(.a(s_45), .O(gate187inter4));
  nand2 gate860(.a(gate187inter4), .b(gate187inter3), .O(gate187inter5));
  nor2  gate861(.a(gate187inter5), .b(gate187inter2), .O(gate187inter6));
  inv1  gate862(.a(G574), .O(gate187inter7));
  inv1  gate863(.a(G575), .O(gate187inter8));
  nand2 gate864(.a(gate187inter8), .b(gate187inter7), .O(gate187inter9));
  nand2 gate865(.a(s_45), .b(gate187inter3), .O(gate187inter10));
  nor2  gate866(.a(gate187inter10), .b(gate187inter9), .O(gate187inter11));
  nor2  gate867(.a(gate187inter11), .b(gate187inter6), .O(gate187inter12));
  nand2 gate868(.a(gate187inter12), .b(gate187inter1), .O(G612));
nand2 gate188( .a(G576), .b(G577), .O(G617) );

  xor2  gate1121(.a(G579), .b(G578), .O(gate189inter0));
  nand2 gate1122(.a(gate189inter0), .b(s_82), .O(gate189inter1));
  and2  gate1123(.a(G579), .b(G578), .O(gate189inter2));
  inv1  gate1124(.a(s_82), .O(gate189inter3));
  inv1  gate1125(.a(s_83), .O(gate189inter4));
  nand2 gate1126(.a(gate189inter4), .b(gate189inter3), .O(gate189inter5));
  nor2  gate1127(.a(gate189inter5), .b(gate189inter2), .O(gate189inter6));
  inv1  gate1128(.a(G578), .O(gate189inter7));
  inv1  gate1129(.a(G579), .O(gate189inter8));
  nand2 gate1130(.a(gate189inter8), .b(gate189inter7), .O(gate189inter9));
  nand2 gate1131(.a(s_83), .b(gate189inter3), .O(gate189inter10));
  nor2  gate1132(.a(gate189inter10), .b(gate189inter9), .O(gate189inter11));
  nor2  gate1133(.a(gate189inter11), .b(gate189inter6), .O(gate189inter12));
  nand2 gate1134(.a(gate189inter12), .b(gate189inter1), .O(G622));
nand2 gate190( .a(G580), .b(G581), .O(G627) );
nand2 gate191( .a(G582), .b(G583), .O(G632) );
nand2 gate192( .a(G584), .b(G585), .O(G637) );
nand2 gate193( .a(G586), .b(G587), .O(G642) );
nand2 gate194( .a(G588), .b(G589), .O(G645) );
nand2 gate195( .a(G590), .b(G591), .O(G648) );
nand2 gate196( .a(G592), .b(G593), .O(G651) );

  xor2  gate673(.a(G595), .b(G594), .O(gate197inter0));
  nand2 gate674(.a(gate197inter0), .b(s_18), .O(gate197inter1));
  and2  gate675(.a(G595), .b(G594), .O(gate197inter2));
  inv1  gate676(.a(s_18), .O(gate197inter3));
  inv1  gate677(.a(s_19), .O(gate197inter4));
  nand2 gate678(.a(gate197inter4), .b(gate197inter3), .O(gate197inter5));
  nor2  gate679(.a(gate197inter5), .b(gate197inter2), .O(gate197inter6));
  inv1  gate680(.a(G594), .O(gate197inter7));
  inv1  gate681(.a(G595), .O(gate197inter8));
  nand2 gate682(.a(gate197inter8), .b(gate197inter7), .O(gate197inter9));
  nand2 gate683(.a(s_19), .b(gate197inter3), .O(gate197inter10));
  nor2  gate684(.a(gate197inter10), .b(gate197inter9), .O(gate197inter11));
  nor2  gate685(.a(gate197inter11), .b(gate197inter6), .O(gate197inter12));
  nand2 gate686(.a(gate197inter12), .b(gate197inter1), .O(G654));
nand2 gate198( .a(G596), .b(G597), .O(G657) );
nand2 gate199( .a(G598), .b(G599), .O(G660) );
nand2 gate200( .a(G600), .b(G601), .O(G663) );
nand2 gate201( .a(G602), .b(G607), .O(G666) );
nand2 gate202( .a(G612), .b(G617), .O(G669) );
nand2 gate203( .a(G602), .b(G612), .O(G672) );
nand2 gate204( .a(G607), .b(G617), .O(G675) );
nand2 gate205( .a(G622), .b(G627), .O(G678) );

  xor2  gate547(.a(G637), .b(G632), .O(gate206inter0));
  nand2 gate548(.a(gate206inter0), .b(s_0), .O(gate206inter1));
  and2  gate549(.a(G637), .b(G632), .O(gate206inter2));
  inv1  gate550(.a(s_0), .O(gate206inter3));
  inv1  gate551(.a(s_1), .O(gate206inter4));
  nand2 gate552(.a(gate206inter4), .b(gate206inter3), .O(gate206inter5));
  nor2  gate553(.a(gate206inter5), .b(gate206inter2), .O(gate206inter6));
  inv1  gate554(.a(G632), .O(gate206inter7));
  inv1  gate555(.a(G637), .O(gate206inter8));
  nand2 gate556(.a(gate206inter8), .b(gate206inter7), .O(gate206inter9));
  nand2 gate557(.a(s_1), .b(gate206inter3), .O(gate206inter10));
  nor2  gate558(.a(gate206inter10), .b(gate206inter9), .O(gate206inter11));
  nor2  gate559(.a(gate206inter11), .b(gate206inter6), .O(gate206inter12));
  nand2 gate560(.a(gate206inter12), .b(gate206inter1), .O(G681));
nand2 gate207( .a(G622), .b(G632), .O(G684) );
nand2 gate208( .a(G627), .b(G637), .O(G687) );
nand2 gate209( .a(G602), .b(G666), .O(G690) );
nand2 gate210( .a(G607), .b(G666), .O(G691) );
nand2 gate211( .a(G612), .b(G669), .O(G692) );
nand2 gate212( .a(G617), .b(G669), .O(G693) );
nand2 gate213( .a(G602), .b(G672), .O(G694) );
nand2 gate214( .a(G612), .b(G672), .O(G695) );
nand2 gate215( .a(G607), .b(G675), .O(G696) );
nand2 gate216( .a(G617), .b(G675), .O(G697) );
nand2 gate217( .a(G622), .b(G678), .O(G698) );

  xor2  gate883(.a(G678), .b(G627), .O(gate218inter0));
  nand2 gate884(.a(gate218inter0), .b(s_48), .O(gate218inter1));
  and2  gate885(.a(G678), .b(G627), .O(gate218inter2));
  inv1  gate886(.a(s_48), .O(gate218inter3));
  inv1  gate887(.a(s_49), .O(gate218inter4));
  nand2 gate888(.a(gate218inter4), .b(gate218inter3), .O(gate218inter5));
  nor2  gate889(.a(gate218inter5), .b(gate218inter2), .O(gate218inter6));
  inv1  gate890(.a(G627), .O(gate218inter7));
  inv1  gate891(.a(G678), .O(gate218inter8));
  nand2 gate892(.a(gate218inter8), .b(gate218inter7), .O(gate218inter9));
  nand2 gate893(.a(s_49), .b(gate218inter3), .O(gate218inter10));
  nor2  gate894(.a(gate218inter10), .b(gate218inter9), .O(gate218inter11));
  nor2  gate895(.a(gate218inter11), .b(gate218inter6), .O(gate218inter12));
  nand2 gate896(.a(gate218inter12), .b(gate218inter1), .O(G699));
nand2 gate219( .a(G632), .b(G681), .O(G700) );
nand2 gate220( .a(G637), .b(G681), .O(G701) );
nand2 gate221( .a(G622), .b(G684), .O(G702) );
nand2 gate222( .a(G632), .b(G684), .O(G703) );
nand2 gate223( .a(G627), .b(G687), .O(G704) );
nand2 gate224( .a(G637), .b(G687), .O(G705) );
nand2 gate225( .a(G690), .b(G691), .O(G706) );
nand2 gate226( .a(G692), .b(G693), .O(G709) );
nand2 gate227( .a(G694), .b(G695), .O(G712) );
nand2 gate228( .a(G696), .b(G697), .O(G715) );
nand2 gate229( .a(G698), .b(G699), .O(G718) );
nand2 gate230( .a(G700), .b(G701), .O(G721) );

  xor2  gate1009(.a(G703), .b(G702), .O(gate231inter0));
  nand2 gate1010(.a(gate231inter0), .b(s_66), .O(gate231inter1));
  and2  gate1011(.a(G703), .b(G702), .O(gate231inter2));
  inv1  gate1012(.a(s_66), .O(gate231inter3));
  inv1  gate1013(.a(s_67), .O(gate231inter4));
  nand2 gate1014(.a(gate231inter4), .b(gate231inter3), .O(gate231inter5));
  nor2  gate1015(.a(gate231inter5), .b(gate231inter2), .O(gate231inter6));
  inv1  gate1016(.a(G702), .O(gate231inter7));
  inv1  gate1017(.a(G703), .O(gate231inter8));
  nand2 gate1018(.a(gate231inter8), .b(gate231inter7), .O(gate231inter9));
  nand2 gate1019(.a(s_67), .b(gate231inter3), .O(gate231inter10));
  nor2  gate1020(.a(gate231inter10), .b(gate231inter9), .O(gate231inter11));
  nor2  gate1021(.a(gate231inter11), .b(gate231inter6), .O(gate231inter12));
  nand2 gate1022(.a(gate231inter12), .b(gate231inter1), .O(G724));

  xor2  gate1317(.a(G705), .b(G704), .O(gate232inter0));
  nand2 gate1318(.a(gate232inter0), .b(s_110), .O(gate232inter1));
  and2  gate1319(.a(G705), .b(G704), .O(gate232inter2));
  inv1  gate1320(.a(s_110), .O(gate232inter3));
  inv1  gate1321(.a(s_111), .O(gate232inter4));
  nand2 gate1322(.a(gate232inter4), .b(gate232inter3), .O(gate232inter5));
  nor2  gate1323(.a(gate232inter5), .b(gate232inter2), .O(gate232inter6));
  inv1  gate1324(.a(G704), .O(gate232inter7));
  inv1  gate1325(.a(G705), .O(gate232inter8));
  nand2 gate1326(.a(gate232inter8), .b(gate232inter7), .O(gate232inter9));
  nand2 gate1327(.a(s_111), .b(gate232inter3), .O(gate232inter10));
  nor2  gate1328(.a(gate232inter10), .b(gate232inter9), .O(gate232inter11));
  nor2  gate1329(.a(gate232inter11), .b(gate232inter6), .O(gate232inter12));
  nand2 gate1330(.a(gate232inter12), .b(gate232inter1), .O(G727));
nand2 gate233( .a(G242), .b(G718), .O(G730) );

  xor2  gate1345(.a(G721), .b(G245), .O(gate234inter0));
  nand2 gate1346(.a(gate234inter0), .b(s_114), .O(gate234inter1));
  and2  gate1347(.a(G721), .b(G245), .O(gate234inter2));
  inv1  gate1348(.a(s_114), .O(gate234inter3));
  inv1  gate1349(.a(s_115), .O(gate234inter4));
  nand2 gate1350(.a(gate234inter4), .b(gate234inter3), .O(gate234inter5));
  nor2  gate1351(.a(gate234inter5), .b(gate234inter2), .O(gate234inter6));
  inv1  gate1352(.a(G245), .O(gate234inter7));
  inv1  gate1353(.a(G721), .O(gate234inter8));
  nand2 gate1354(.a(gate234inter8), .b(gate234inter7), .O(gate234inter9));
  nand2 gate1355(.a(s_115), .b(gate234inter3), .O(gate234inter10));
  nor2  gate1356(.a(gate234inter10), .b(gate234inter9), .O(gate234inter11));
  nor2  gate1357(.a(gate234inter11), .b(gate234inter6), .O(gate234inter12));
  nand2 gate1358(.a(gate234inter12), .b(gate234inter1), .O(G733));

  xor2  gate1331(.a(G724), .b(G248), .O(gate235inter0));
  nand2 gate1332(.a(gate235inter0), .b(s_112), .O(gate235inter1));
  and2  gate1333(.a(G724), .b(G248), .O(gate235inter2));
  inv1  gate1334(.a(s_112), .O(gate235inter3));
  inv1  gate1335(.a(s_113), .O(gate235inter4));
  nand2 gate1336(.a(gate235inter4), .b(gate235inter3), .O(gate235inter5));
  nor2  gate1337(.a(gate235inter5), .b(gate235inter2), .O(gate235inter6));
  inv1  gate1338(.a(G248), .O(gate235inter7));
  inv1  gate1339(.a(G724), .O(gate235inter8));
  nand2 gate1340(.a(gate235inter8), .b(gate235inter7), .O(gate235inter9));
  nand2 gate1341(.a(s_113), .b(gate235inter3), .O(gate235inter10));
  nor2  gate1342(.a(gate235inter10), .b(gate235inter9), .O(gate235inter11));
  nor2  gate1343(.a(gate235inter11), .b(gate235inter6), .O(gate235inter12));
  nand2 gate1344(.a(gate235inter12), .b(gate235inter1), .O(G736));
nand2 gate236( .a(G251), .b(G727), .O(G739) );

  xor2  gate1023(.a(G706), .b(G254), .O(gate237inter0));
  nand2 gate1024(.a(gate237inter0), .b(s_68), .O(gate237inter1));
  and2  gate1025(.a(G706), .b(G254), .O(gate237inter2));
  inv1  gate1026(.a(s_68), .O(gate237inter3));
  inv1  gate1027(.a(s_69), .O(gate237inter4));
  nand2 gate1028(.a(gate237inter4), .b(gate237inter3), .O(gate237inter5));
  nor2  gate1029(.a(gate237inter5), .b(gate237inter2), .O(gate237inter6));
  inv1  gate1030(.a(G254), .O(gate237inter7));
  inv1  gate1031(.a(G706), .O(gate237inter8));
  nand2 gate1032(.a(gate237inter8), .b(gate237inter7), .O(gate237inter9));
  nand2 gate1033(.a(s_69), .b(gate237inter3), .O(gate237inter10));
  nor2  gate1034(.a(gate237inter10), .b(gate237inter9), .O(gate237inter11));
  nor2  gate1035(.a(gate237inter11), .b(gate237inter6), .O(gate237inter12));
  nand2 gate1036(.a(gate237inter12), .b(gate237inter1), .O(G742));
nand2 gate238( .a(G257), .b(G709), .O(G745) );
nand2 gate239( .a(G260), .b(G712), .O(G748) );
nand2 gate240( .a(G263), .b(G715), .O(G751) );
nand2 gate241( .a(G242), .b(G730), .O(G754) );

  xor2  gate1387(.a(G730), .b(G718), .O(gate242inter0));
  nand2 gate1388(.a(gate242inter0), .b(s_120), .O(gate242inter1));
  and2  gate1389(.a(G730), .b(G718), .O(gate242inter2));
  inv1  gate1390(.a(s_120), .O(gate242inter3));
  inv1  gate1391(.a(s_121), .O(gate242inter4));
  nand2 gate1392(.a(gate242inter4), .b(gate242inter3), .O(gate242inter5));
  nor2  gate1393(.a(gate242inter5), .b(gate242inter2), .O(gate242inter6));
  inv1  gate1394(.a(G718), .O(gate242inter7));
  inv1  gate1395(.a(G730), .O(gate242inter8));
  nand2 gate1396(.a(gate242inter8), .b(gate242inter7), .O(gate242inter9));
  nand2 gate1397(.a(s_121), .b(gate242inter3), .O(gate242inter10));
  nor2  gate1398(.a(gate242inter10), .b(gate242inter9), .O(gate242inter11));
  nor2  gate1399(.a(gate242inter11), .b(gate242inter6), .O(gate242inter12));
  nand2 gate1400(.a(gate242inter12), .b(gate242inter1), .O(G755));
nand2 gate243( .a(G245), .b(G733), .O(G756) );
nand2 gate244( .a(G721), .b(G733), .O(G757) );
nand2 gate245( .a(G248), .b(G736), .O(G758) );
nand2 gate246( .a(G724), .b(G736), .O(G759) );
nand2 gate247( .a(G251), .b(G739), .O(G760) );
nand2 gate248( .a(G727), .b(G739), .O(G761) );
nand2 gate249( .a(G254), .b(G742), .O(G762) );
nand2 gate250( .a(G706), .b(G742), .O(G763) );
nand2 gate251( .a(G257), .b(G745), .O(G764) );
nand2 gate252( .a(G709), .b(G745), .O(G765) );
nand2 gate253( .a(G260), .b(G748), .O(G766) );
nand2 gate254( .a(G712), .b(G748), .O(G767) );

  xor2  gate1191(.a(G751), .b(G263), .O(gate255inter0));
  nand2 gate1192(.a(gate255inter0), .b(s_92), .O(gate255inter1));
  and2  gate1193(.a(G751), .b(G263), .O(gate255inter2));
  inv1  gate1194(.a(s_92), .O(gate255inter3));
  inv1  gate1195(.a(s_93), .O(gate255inter4));
  nand2 gate1196(.a(gate255inter4), .b(gate255inter3), .O(gate255inter5));
  nor2  gate1197(.a(gate255inter5), .b(gate255inter2), .O(gate255inter6));
  inv1  gate1198(.a(G263), .O(gate255inter7));
  inv1  gate1199(.a(G751), .O(gate255inter8));
  nand2 gate1200(.a(gate255inter8), .b(gate255inter7), .O(gate255inter9));
  nand2 gate1201(.a(s_93), .b(gate255inter3), .O(gate255inter10));
  nor2  gate1202(.a(gate255inter10), .b(gate255inter9), .O(gate255inter11));
  nor2  gate1203(.a(gate255inter11), .b(gate255inter6), .O(gate255inter12));
  nand2 gate1204(.a(gate255inter12), .b(gate255inter1), .O(G768));
nand2 gate256( .a(G715), .b(G751), .O(G769) );
nand2 gate257( .a(G754), .b(G755), .O(G770) );
nand2 gate258( .a(G756), .b(G757), .O(G773) );
nand2 gate259( .a(G758), .b(G759), .O(G776) );
nand2 gate260( .a(G760), .b(G761), .O(G779) );
nand2 gate261( .a(G762), .b(G763), .O(G782) );
nand2 gate262( .a(G764), .b(G765), .O(G785) );
nand2 gate263( .a(G766), .b(G767), .O(G788) );

  xor2  gate617(.a(G769), .b(G768), .O(gate264inter0));
  nand2 gate618(.a(gate264inter0), .b(s_10), .O(gate264inter1));
  and2  gate619(.a(G769), .b(G768), .O(gate264inter2));
  inv1  gate620(.a(s_10), .O(gate264inter3));
  inv1  gate621(.a(s_11), .O(gate264inter4));
  nand2 gate622(.a(gate264inter4), .b(gate264inter3), .O(gate264inter5));
  nor2  gate623(.a(gate264inter5), .b(gate264inter2), .O(gate264inter6));
  inv1  gate624(.a(G768), .O(gate264inter7));
  inv1  gate625(.a(G769), .O(gate264inter8));
  nand2 gate626(.a(gate264inter8), .b(gate264inter7), .O(gate264inter9));
  nand2 gate627(.a(s_11), .b(gate264inter3), .O(gate264inter10));
  nor2  gate628(.a(gate264inter10), .b(gate264inter9), .O(gate264inter11));
  nor2  gate629(.a(gate264inter11), .b(gate264inter6), .O(gate264inter12));
  nand2 gate630(.a(gate264inter12), .b(gate264inter1), .O(G791));
nand2 gate265( .a(G642), .b(G770), .O(G794) );
nand2 gate266( .a(G645), .b(G773), .O(G797) );
nand2 gate267( .a(G648), .b(G776), .O(G800) );

  xor2  gate1401(.a(G779), .b(G651), .O(gate268inter0));
  nand2 gate1402(.a(gate268inter0), .b(s_122), .O(gate268inter1));
  and2  gate1403(.a(G779), .b(G651), .O(gate268inter2));
  inv1  gate1404(.a(s_122), .O(gate268inter3));
  inv1  gate1405(.a(s_123), .O(gate268inter4));
  nand2 gate1406(.a(gate268inter4), .b(gate268inter3), .O(gate268inter5));
  nor2  gate1407(.a(gate268inter5), .b(gate268inter2), .O(gate268inter6));
  inv1  gate1408(.a(G651), .O(gate268inter7));
  inv1  gate1409(.a(G779), .O(gate268inter8));
  nand2 gate1410(.a(gate268inter8), .b(gate268inter7), .O(gate268inter9));
  nand2 gate1411(.a(s_123), .b(gate268inter3), .O(gate268inter10));
  nor2  gate1412(.a(gate268inter10), .b(gate268inter9), .O(gate268inter11));
  nor2  gate1413(.a(gate268inter11), .b(gate268inter6), .O(gate268inter12));
  nand2 gate1414(.a(gate268inter12), .b(gate268inter1), .O(G803));
nand2 gate269( .a(G654), .b(G782), .O(G806) );
nand2 gate270( .a(G657), .b(G785), .O(G809) );
nand2 gate271( .a(G660), .b(G788), .O(G812) );
nand2 gate272( .a(G663), .b(G791), .O(G815) );
nand2 gate273( .a(G642), .b(G794), .O(G818) );
nand2 gate274( .a(G770), .b(G794), .O(G819) );
nand2 gate275( .a(G645), .b(G797), .O(G820) );
nand2 gate276( .a(G773), .b(G797), .O(G821) );
nand2 gate277( .a(G648), .b(G800), .O(G822) );

  xor2  gate729(.a(G800), .b(G776), .O(gate278inter0));
  nand2 gate730(.a(gate278inter0), .b(s_26), .O(gate278inter1));
  and2  gate731(.a(G800), .b(G776), .O(gate278inter2));
  inv1  gate732(.a(s_26), .O(gate278inter3));
  inv1  gate733(.a(s_27), .O(gate278inter4));
  nand2 gate734(.a(gate278inter4), .b(gate278inter3), .O(gate278inter5));
  nor2  gate735(.a(gate278inter5), .b(gate278inter2), .O(gate278inter6));
  inv1  gate736(.a(G776), .O(gate278inter7));
  inv1  gate737(.a(G800), .O(gate278inter8));
  nand2 gate738(.a(gate278inter8), .b(gate278inter7), .O(gate278inter9));
  nand2 gate739(.a(s_27), .b(gate278inter3), .O(gate278inter10));
  nor2  gate740(.a(gate278inter10), .b(gate278inter9), .O(gate278inter11));
  nor2  gate741(.a(gate278inter11), .b(gate278inter6), .O(gate278inter12));
  nand2 gate742(.a(gate278inter12), .b(gate278inter1), .O(G823));
nand2 gate279( .a(G651), .b(G803), .O(G824) );
nand2 gate280( .a(G779), .b(G803), .O(G825) );
nand2 gate281( .a(G654), .b(G806), .O(G826) );
nand2 gate282( .a(G782), .b(G806), .O(G827) );
nand2 gate283( .a(G657), .b(G809), .O(G828) );
nand2 gate284( .a(G785), .b(G809), .O(G829) );
nand2 gate285( .a(G660), .b(G812), .O(G830) );
nand2 gate286( .a(G788), .b(G812), .O(G831) );
nand2 gate287( .a(G663), .b(G815), .O(G832) );
nand2 gate288( .a(G791), .b(G815), .O(G833) );
nand2 gate289( .a(G818), .b(G819), .O(G834) );
nand2 gate290( .a(G820), .b(G821), .O(G847) );

  xor2  gate939(.a(G823), .b(G822), .O(gate291inter0));
  nand2 gate940(.a(gate291inter0), .b(s_56), .O(gate291inter1));
  and2  gate941(.a(G823), .b(G822), .O(gate291inter2));
  inv1  gate942(.a(s_56), .O(gate291inter3));
  inv1  gate943(.a(s_57), .O(gate291inter4));
  nand2 gate944(.a(gate291inter4), .b(gate291inter3), .O(gate291inter5));
  nor2  gate945(.a(gate291inter5), .b(gate291inter2), .O(gate291inter6));
  inv1  gate946(.a(G822), .O(gate291inter7));
  inv1  gate947(.a(G823), .O(gate291inter8));
  nand2 gate948(.a(gate291inter8), .b(gate291inter7), .O(gate291inter9));
  nand2 gate949(.a(s_57), .b(gate291inter3), .O(gate291inter10));
  nor2  gate950(.a(gate291inter10), .b(gate291inter9), .O(gate291inter11));
  nor2  gate951(.a(gate291inter11), .b(gate291inter6), .O(gate291inter12));
  nand2 gate952(.a(gate291inter12), .b(gate291inter1), .O(G860));
nand2 gate292( .a(G824), .b(G825), .O(G873) );
nand2 gate293( .a(G828), .b(G829), .O(G886) );
nand2 gate294( .a(G832), .b(G833), .O(G899) );
nand2 gate295( .a(G830), .b(G831), .O(G912) );

  xor2  gate561(.a(G827), .b(G826), .O(gate296inter0));
  nand2 gate562(.a(gate296inter0), .b(s_2), .O(gate296inter1));
  and2  gate563(.a(G827), .b(G826), .O(gate296inter2));
  inv1  gate564(.a(s_2), .O(gate296inter3));
  inv1  gate565(.a(s_3), .O(gate296inter4));
  nand2 gate566(.a(gate296inter4), .b(gate296inter3), .O(gate296inter5));
  nor2  gate567(.a(gate296inter5), .b(gate296inter2), .O(gate296inter6));
  inv1  gate568(.a(G826), .O(gate296inter7));
  inv1  gate569(.a(G827), .O(gate296inter8));
  nand2 gate570(.a(gate296inter8), .b(gate296inter7), .O(gate296inter9));
  nand2 gate571(.a(s_3), .b(gate296inter3), .O(gate296inter10));
  nor2  gate572(.a(gate296inter10), .b(gate296inter9), .O(gate296inter11));
  nor2  gate573(.a(gate296inter11), .b(gate296inter6), .O(gate296inter12));
  nand2 gate574(.a(gate296inter12), .b(gate296inter1), .O(G925));
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );
nand2 gate387( .a(G1), .b(G1036), .O(G1132) );
nand2 gate388( .a(G2), .b(G1039), .O(G1135) );
nand2 gate389( .a(G3), .b(G1042), .O(G1138) );
nand2 gate390( .a(G4), .b(G1045), .O(G1141) );
nand2 gate391( .a(G5), .b(G1048), .O(G1144) );
nand2 gate392( .a(G6), .b(G1051), .O(G1147) );
nand2 gate393( .a(G7), .b(G1054), .O(G1150) );
nand2 gate394( .a(G8), .b(G1057), .O(G1153) );
nand2 gate395( .a(G9), .b(G1060), .O(G1156) );
nand2 gate396( .a(G10), .b(G1063), .O(G1159) );
nand2 gate397( .a(G11), .b(G1066), .O(G1162) );

  xor2  gate631(.a(G1069), .b(G12), .O(gate398inter0));
  nand2 gate632(.a(gate398inter0), .b(s_12), .O(gate398inter1));
  and2  gate633(.a(G1069), .b(G12), .O(gate398inter2));
  inv1  gate634(.a(s_12), .O(gate398inter3));
  inv1  gate635(.a(s_13), .O(gate398inter4));
  nand2 gate636(.a(gate398inter4), .b(gate398inter3), .O(gate398inter5));
  nor2  gate637(.a(gate398inter5), .b(gate398inter2), .O(gate398inter6));
  inv1  gate638(.a(G12), .O(gate398inter7));
  inv1  gate639(.a(G1069), .O(gate398inter8));
  nand2 gate640(.a(gate398inter8), .b(gate398inter7), .O(gate398inter9));
  nand2 gate641(.a(s_13), .b(gate398inter3), .O(gate398inter10));
  nor2  gate642(.a(gate398inter10), .b(gate398inter9), .O(gate398inter11));
  nor2  gate643(.a(gate398inter11), .b(gate398inter6), .O(gate398inter12));
  nand2 gate644(.a(gate398inter12), .b(gate398inter1), .O(G1165));
nand2 gate399( .a(G13), .b(G1072), .O(G1168) );
nand2 gate400( .a(G14), .b(G1075), .O(G1171) );
nand2 gate401( .a(G15), .b(G1078), .O(G1174) );
nand2 gate402( .a(G16), .b(G1081), .O(G1177) );

  xor2  gate813(.a(G1084), .b(G17), .O(gate403inter0));
  nand2 gate814(.a(gate403inter0), .b(s_38), .O(gate403inter1));
  and2  gate815(.a(G1084), .b(G17), .O(gate403inter2));
  inv1  gate816(.a(s_38), .O(gate403inter3));
  inv1  gate817(.a(s_39), .O(gate403inter4));
  nand2 gate818(.a(gate403inter4), .b(gate403inter3), .O(gate403inter5));
  nor2  gate819(.a(gate403inter5), .b(gate403inter2), .O(gate403inter6));
  inv1  gate820(.a(G17), .O(gate403inter7));
  inv1  gate821(.a(G1084), .O(gate403inter8));
  nand2 gate822(.a(gate403inter8), .b(gate403inter7), .O(gate403inter9));
  nand2 gate823(.a(s_39), .b(gate403inter3), .O(gate403inter10));
  nor2  gate824(.a(gate403inter10), .b(gate403inter9), .O(gate403inter11));
  nor2  gate825(.a(gate403inter11), .b(gate403inter6), .O(gate403inter12));
  nand2 gate826(.a(gate403inter12), .b(gate403inter1), .O(G1180));
nand2 gate404( .a(G18), .b(G1087), .O(G1183) );
nand2 gate405( .a(G19), .b(G1090), .O(G1186) );
nand2 gate406( .a(G20), .b(G1093), .O(G1189) );
nand2 gate407( .a(G21), .b(G1096), .O(G1192) );
nand2 gate408( .a(G22), .b(G1099), .O(G1195) );
nand2 gate409( .a(G23), .b(G1102), .O(G1198) );

  xor2  gate715(.a(G1105), .b(G24), .O(gate410inter0));
  nand2 gate716(.a(gate410inter0), .b(s_24), .O(gate410inter1));
  and2  gate717(.a(G1105), .b(G24), .O(gate410inter2));
  inv1  gate718(.a(s_24), .O(gate410inter3));
  inv1  gate719(.a(s_25), .O(gate410inter4));
  nand2 gate720(.a(gate410inter4), .b(gate410inter3), .O(gate410inter5));
  nor2  gate721(.a(gate410inter5), .b(gate410inter2), .O(gate410inter6));
  inv1  gate722(.a(G24), .O(gate410inter7));
  inv1  gate723(.a(G1105), .O(gate410inter8));
  nand2 gate724(.a(gate410inter8), .b(gate410inter7), .O(gate410inter9));
  nand2 gate725(.a(s_25), .b(gate410inter3), .O(gate410inter10));
  nor2  gate726(.a(gate410inter10), .b(gate410inter9), .O(gate410inter11));
  nor2  gate727(.a(gate410inter11), .b(gate410inter6), .O(gate410inter12));
  nand2 gate728(.a(gate410inter12), .b(gate410inter1), .O(G1201));
nand2 gate411( .a(G25), .b(G1108), .O(G1204) );

  xor2  gate589(.a(G1111), .b(G26), .O(gate412inter0));
  nand2 gate590(.a(gate412inter0), .b(s_6), .O(gate412inter1));
  and2  gate591(.a(G1111), .b(G26), .O(gate412inter2));
  inv1  gate592(.a(s_6), .O(gate412inter3));
  inv1  gate593(.a(s_7), .O(gate412inter4));
  nand2 gate594(.a(gate412inter4), .b(gate412inter3), .O(gate412inter5));
  nor2  gate595(.a(gate412inter5), .b(gate412inter2), .O(gate412inter6));
  inv1  gate596(.a(G26), .O(gate412inter7));
  inv1  gate597(.a(G1111), .O(gate412inter8));
  nand2 gate598(.a(gate412inter8), .b(gate412inter7), .O(gate412inter9));
  nand2 gate599(.a(s_7), .b(gate412inter3), .O(gate412inter10));
  nor2  gate600(.a(gate412inter10), .b(gate412inter9), .O(gate412inter11));
  nor2  gate601(.a(gate412inter11), .b(gate412inter6), .O(gate412inter12));
  nand2 gate602(.a(gate412inter12), .b(gate412inter1), .O(G1207));

  xor2  gate1051(.a(G1114), .b(G27), .O(gate413inter0));
  nand2 gate1052(.a(gate413inter0), .b(s_72), .O(gate413inter1));
  and2  gate1053(.a(G1114), .b(G27), .O(gate413inter2));
  inv1  gate1054(.a(s_72), .O(gate413inter3));
  inv1  gate1055(.a(s_73), .O(gate413inter4));
  nand2 gate1056(.a(gate413inter4), .b(gate413inter3), .O(gate413inter5));
  nor2  gate1057(.a(gate413inter5), .b(gate413inter2), .O(gate413inter6));
  inv1  gate1058(.a(G27), .O(gate413inter7));
  inv1  gate1059(.a(G1114), .O(gate413inter8));
  nand2 gate1060(.a(gate413inter8), .b(gate413inter7), .O(gate413inter9));
  nand2 gate1061(.a(s_73), .b(gate413inter3), .O(gate413inter10));
  nor2  gate1062(.a(gate413inter10), .b(gate413inter9), .O(gate413inter11));
  nor2  gate1063(.a(gate413inter11), .b(gate413inter6), .O(gate413inter12));
  nand2 gate1064(.a(gate413inter12), .b(gate413inter1), .O(G1210));
nand2 gate414( .a(G28), .b(G1117), .O(G1213) );
nand2 gate415( .a(G29), .b(G1120), .O(G1216) );
nand2 gate416( .a(G30), .b(G1123), .O(G1219) );

  xor2  gate771(.a(G1126), .b(G31), .O(gate417inter0));
  nand2 gate772(.a(gate417inter0), .b(s_32), .O(gate417inter1));
  and2  gate773(.a(G1126), .b(G31), .O(gate417inter2));
  inv1  gate774(.a(s_32), .O(gate417inter3));
  inv1  gate775(.a(s_33), .O(gate417inter4));
  nand2 gate776(.a(gate417inter4), .b(gate417inter3), .O(gate417inter5));
  nor2  gate777(.a(gate417inter5), .b(gate417inter2), .O(gate417inter6));
  inv1  gate778(.a(G31), .O(gate417inter7));
  inv1  gate779(.a(G1126), .O(gate417inter8));
  nand2 gate780(.a(gate417inter8), .b(gate417inter7), .O(gate417inter9));
  nand2 gate781(.a(s_33), .b(gate417inter3), .O(gate417inter10));
  nor2  gate782(.a(gate417inter10), .b(gate417inter9), .O(gate417inter11));
  nor2  gate783(.a(gate417inter11), .b(gate417inter6), .O(gate417inter12));
  nand2 gate784(.a(gate417inter12), .b(gate417inter1), .O(G1222));
nand2 gate418( .a(G32), .b(G1129), .O(G1225) );
nand2 gate419( .a(G1), .b(G1132), .O(G1228) );
nand2 gate420( .a(G1036), .b(G1132), .O(G1229) );
nand2 gate421( .a(G2), .b(G1135), .O(G1230) );
nand2 gate422( .a(G1039), .b(G1135), .O(G1231) );
nand2 gate423( .a(G3), .b(G1138), .O(G1232) );
nand2 gate424( .a(G1042), .b(G1138), .O(G1233) );
nand2 gate425( .a(G4), .b(G1141), .O(G1234) );
nand2 gate426( .a(G1045), .b(G1141), .O(G1235) );
nand2 gate427( .a(G5), .b(G1144), .O(G1236) );
nand2 gate428( .a(G1048), .b(G1144), .O(G1237) );
nand2 gate429( .a(G6), .b(G1147), .O(G1238) );
nand2 gate430( .a(G1051), .b(G1147), .O(G1239) );
nand2 gate431( .a(G7), .b(G1150), .O(G1240) );

  xor2  gate925(.a(G1150), .b(G1054), .O(gate432inter0));
  nand2 gate926(.a(gate432inter0), .b(s_54), .O(gate432inter1));
  and2  gate927(.a(G1150), .b(G1054), .O(gate432inter2));
  inv1  gate928(.a(s_54), .O(gate432inter3));
  inv1  gate929(.a(s_55), .O(gate432inter4));
  nand2 gate930(.a(gate432inter4), .b(gate432inter3), .O(gate432inter5));
  nor2  gate931(.a(gate432inter5), .b(gate432inter2), .O(gate432inter6));
  inv1  gate932(.a(G1054), .O(gate432inter7));
  inv1  gate933(.a(G1150), .O(gate432inter8));
  nand2 gate934(.a(gate432inter8), .b(gate432inter7), .O(gate432inter9));
  nand2 gate935(.a(s_55), .b(gate432inter3), .O(gate432inter10));
  nor2  gate936(.a(gate432inter10), .b(gate432inter9), .O(gate432inter11));
  nor2  gate937(.a(gate432inter11), .b(gate432inter6), .O(gate432inter12));
  nand2 gate938(.a(gate432inter12), .b(gate432inter1), .O(G1241));
nand2 gate433( .a(G8), .b(G1153), .O(G1242) );
nand2 gate434( .a(G1057), .b(G1153), .O(G1243) );

  xor2  gate1233(.a(G1156), .b(G9), .O(gate435inter0));
  nand2 gate1234(.a(gate435inter0), .b(s_98), .O(gate435inter1));
  and2  gate1235(.a(G1156), .b(G9), .O(gate435inter2));
  inv1  gate1236(.a(s_98), .O(gate435inter3));
  inv1  gate1237(.a(s_99), .O(gate435inter4));
  nand2 gate1238(.a(gate435inter4), .b(gate435inter3), .O(gate435inter5));
  nor2  gate1239(.a(gate435inter5), .b(gate435inter2), .O(gate435inter6));
  inv1  gate1240(.a(G9), .O(gate435inter7));
  inv1  gate1241(.a(G1156), .O(gate435inter8));
  nand2 gate1242(.a(gate435inter8), .b(gate435inter7), .O(gate435inter9));
  nand2 gate1243(.a(s_99), .b(gate435inter3), .O(gate435inter10));
  nor2  gate1244(.a(gate435inter10), .b(gate435inter9), .O(gate435inter11));
  nor2  gate1245(.a(gate435inter11), .b(gate435inter6), .O(gate435inter12));
  nand2 gate1246(.a(gate435inter12), .b(gate435inter1), .O(G1244));
nand2 gate436( .a(G1060), .b(G1156), .O(G1245) );
nand2 gate437( .a(G10), .b(G1159), .O(G1246) );
nand2 gate438( .a(G1063), .b(G1159), .O(G1247) );
nand2 gate439( .a(G11), .b(G1162), .O(G1248) );
nand2 gate440( .a(G1066), .b(G1162), .O(G1249) );
nand2 gate441( .a(G12), .b(G1165), .O(G1250) );
nand2 gate442( .a(G1069), .b(G1165), .O(G1251) );
nand2 gate443( .a(G13), .b(G1168), .O(G1252) );
nand2 gate444( .a(G1072), .b(G1168), .O(G1253) );
nand2 gate445( .a(G14), .b(G1171), .O(G1254) );
nand2 gate446( .a(G1075), .b(G1171), .O(G1255) );
nand2 gate447( .a(G15), .b(G1174), .O(G1256) );
nand2 gate448( .a(G1078), .b(G1174), .O(G1257) );
nand2 gate449( .a(G16), .b(G1177), .O(G1258) );
nand2 gate450( .a(G1081), .b(G1177), .O(G1259) );
nand2 gate451( .a(G17), .b(G1180), .O(G1260) );
nand2 gate452( .a(G1084), .b(G1180), .O(G1261) );
nand2 gate453( .a(G18), .b(G1183), .O(G1262) );
nand2 gate454( .a(G1087), .b(G1183), .O(G1263) );
nand2 gate455( .a(G19), .b(G1186), .O(G1264) );
nand2 gate456( .a(G1090), .b(G1186), .O(G1265) );
nand2 gate457( .a(G20), .b(G1189), .O(G1266) );
nand2 gate458( .a(G1093), .b(G1189), .O(G1267) );
nand2 gate459( .a(G21), .b(G1192), .O(G1268) );

  xor2  gate659(.a(G1192), .b(G1096), .O(gate460inter0));
  nand2 gate660(.a(gate460inter0), .b(s_16), .O(gate460inter1));
  and2  gate661(.a(G1192), .b(G1096), .O(gate460inter2));
  inv1  gate662(.a(s_16), .O(gate460inter3));
  inv1  gate663(.a(s_17), .O(gate460inter4));
  nand2 gate664(.a(gate460inter4), .b(gate460inter3), .O(gate460inter5));
  nor2  gate665(.a(gate460inter5), .b(gate460inter2), .O(gate460inter6));
  inv1  gate666(.a(G1096), .O(gate460inter7));
  inv1  gate667(.a(G1192), .O(gate460inter8));
  nand2 gate668(.a(gate460inter8), .b(gate460inter7), .O(gate460inter9));
  nand2 gate669(.a(s_17), .b(gate460inter3), .O(gate460inter10));
  nor2  gate670(.a(gate460inter10), .b(gate460inter9), .O(gate460inter11));
  nor2  gate671(.a(gate460inter11), .b(gate460inter6), .O(gate460inter12));
  nand2 gate672(.a(gate460inter12), .b(gate460inter1), .O(G1269));
nand2 gate461( .a(G22), .b(G1195), .O(G1270) );
nand2 gate462( .a(G1099), .b(G1195), .O(G1271) );
nand2 gate463( .a(G23), .b(G1198), .O(G1272) );

  xor2  gate757(.a(G1198), .b(G1102), .O(gate464inter0));
  nand2 gate758(.a(gate464inter0), .b(s_30), .O(gate464inter1));
  and2  gate759(.a(G1198), .b(G1102), .O(gate464inter2));
  inv1  gate760(.a(s_30), .O(gate464inter3));
  inv1  gate761(.a(s_31), .O(gate464inter4));
  nand2 gate762(.a(gate464inter4), .b(gate464inter3), .O(gate464inter5));
  nor2  gate763(.a(gate464inter5), .b(gate464inter2), .O(gate464inter6));
  inv1  gate764(.a(G1102), .O(gate464inter7));
  inv1  gate765(.a(G1198), .O(gate464inter8));
  nand2 gate766(.a(gate464inter8), .b(gate464inter7), .O(gate464inter9));
  nand2 gate767(.a(s_31), .b(gate464inter3), .O(gate464inter10));
  nor2  gate768(.a(gate464inter10), .b(gate464inter9), .O(gate464inter11));
  nor2  gate769(.a(gate464inter11), .b(gate464inter6), .O(gate464inter12));
  nand2 gate770(.a(gate464inter12), .b(gate464inter1), .O(G1273));
nand2 gate465( .a(G24), .b(G1201), .O(G1274) );
nand2 gate466( .a(G1105), .b(G1201), .O(G1275) );
nand2 gate467( .a(G25), .b(G1204), .O(G1276) );

  xor2  gate1247(.a(G1204), .b(G1108), .O(gate468inter0));
  nand2 gate1248(.a(gate468inter0), .b(s_100), .O(gate468inter1));
  and2  gate1249(.a(G1204), .b(G1108), .O(gate468inter2));
  inv1  gate1250(.a(s_100), .O(gate468inter3));
  inv1  gate1251(.a(s_101), .O(gate468inter4));
  nand2 gate1252(.a(gate468inter4), .b(gate468inter3), .O(gate468inter5));
  nor2  gate1253(.a(gate468inter5), .b(gate468inter2), .O(gate468inter6));
  inv1  gate1254(.a(G1108), .O(gate468inter7));
  inv1  gate1255(.a(G1204), .O(gate468inter8));
  nand2 gate1256(.a(gate468inter8), .b(gate468inter7), .O(gate468inter9));
  nand2 gate1257(.a(s_101), .b(gate468inter3), .O(gate468inter10));
  nor2  gate1258(.a(gate468inter10), .b(gate468inter9), .O(gate468inter11));
  nor2  gate1259(.a(gate468inter11), .b(gate468inter6), .O(gate468inter12));
  nand2 gate1260(.a(gate468inter12), .b(gate468inter1), .O(G1277));
nand2 gate469( .a(G26), .b(G1207), .O(G1278) );
nand2 gate470( .a(G1111), .b(G1207), .O(G1279) );

  xor2  gate785(.a(G1210), .b(G27), .O(gate471inter0));
  nand2 gate786(.a(gate471inter0), .b(s_34), .O(gate471inter1));
  and2  gate787(.a(G1210), .b(G27), .O(gate471inter2));
  inv1  gate788(.a(s_34), .O(gate471inter3));
  inv1  gate789(.a(s_35), .O(gate471inter4));
  nand2 gate790(.a(gate471inter4), .b(gate471inter3), .O(gate471inter5));
  nor2  gate791(.a(gate471inter5), .b(gate471inter2), .O(gate471inter6));
  inv1  gate792(.a(G27), .O(gate471inter7));
  inv1  gate793(.a(G1210), .O(gate471inter8));
  nand2 gate794(.a(gate471inter8), .b(gate471inter7), .O(gate471inter9));
  nand2 gate795(.a(s_35), .b(gate471inter3), .O(gate471inter10));
  nor2  gate796(.a(gate471inter10), .b(gate471inter9), .O(gate471inter11));
  nor2  gate797(.a(gate471inter11), .b(gate471inter6), .O(gate471inter12));
  nand2 gate798(.a(gate471inter12), .b(gate471inter1), .O(G1280));
nand2 gate472( .a(G1114), .b(G1210), .O(G1281) );
nand2 gate473( .a(G28), .b(G1213), .O(G1282) );
nand2 gate474( .a(G1117), .b(G1213), .O(G1283) );
nand2 gate475( .a(G29), .b(G1216), .O(G1284) );
nand2 gate476( .a(G1120), .b(G1216), .O(G1285) );
nand2 gate477( .a(G30), .b(G1219), .O(G1286) );
nand2 gate478( .a(G1123), .b(G1219), .O(G1287) );
nand2 gate479( .a(G31), .b(G1222), .O(G1288) );
nand2 gate480( .a(G1126), .b(G1222), .O(G1289) );
nand2 gate481( .a(G32), .b(G1225), .O(G1290) );
nand2 gate482( .a(G1129), .b(G1225), .O(G1291) );
nand2 gate483( .a(G1228), .b(G1229), .O(G1292) );

  xor2  gate953(.a(G1231), .b(G1230), .O(gate484inter0));
  nand2 gate954(.a(gate484inter0), .b(s_58), .O(gate484inter1));
  and2  gate955(.a(G1231), .b(G1230), .O(gate484inter2));
  inv1  gate956(.a(s_58), .O(gate484inter3));
  inv1  gate957(.a(s_59), .O(gate484inter4));
  nand2 gate958(.a(gate484inter4), .b(gate484inter3), .O(gate484inter5));
  nor2  gate959(.a(gate484inter5), .b(gate484inter2), .O(gate484inter6));
  inv1  gate960(.a(G1230), .O(gate484inter7));
  inv1  gate961(.a(G1231), .O(gate484inter8));
  nand2 gate962(.a(gate484inter8), .b(gate484inter7), .O(gate484inter9));
  nand2 gate963(.a(s_59), .b(gate484inter3), .O(gate484inter10));
  nor2  gate964(.a(gate484inter10), .b(gate484inter9), .O(gate484inter11));
  nor2  gate965(.a(gate484inter11), .b(gate484inter6), .O(gate484inter12));
  nand2 gate966(.a(gate484inter12), .b(gate484inter1), .O(G1293));
nand2 gate485( .a(G1232), .b(G1233), .O(G1294) );
nand2 gate486( .a(G1234), .b(G1235), .O(G1295) );
nand2 gate487( .a(G1236), .b(G1237), .O(G1296) );

  xor2  gate1303(.a(G1239), .b(G1238), .O(gate488inter0));
  nand2 gate1304(.a(gate488inter0), .b(s_108), .O(gate488inter1));
  and2  gate1305(.a(G1239), .b(G1238), .O(gate488inter2));
  inv1  gate1306(.a(s_108), .O(gate488inter3));
  inv1  gate1307(.a(s_109), .O(gate488inter4));
  nand2 gate1308(.a(gate488inter4), .b(gate488inter3), .O(gate488inter5));
  nor2  gate1309(.a(gate488inter5), .b(gate488inter2), .O(gate488inter6));
  inv1  gate1310(.a(G1238), .O(gate488inter7));
  inv1  gate1311(.a(G1239), .O(gate488inter8));
  nand2 gate1312(.a(gate488inter8), .b(gate488inter7), .O(gate488inter9));
  nand2 gate1313(.a(s_109), .b(gate488inter3), .O(gate488inter10));
  nor2  gate1314(.a(gate488inter10), .b(gate488inter9), .O(gate488inter11));
  nor2  gate1315(.a(gate488inter11), .b(gate488inter6), .O(gate488inter12));
  nand2 gate1316(.a(gate488inter12), .b(gate488inter1), .O(G1297));

  xor2  gate911(.a(G1241), .b(G1240), .O(gate489inter0));
  nand2 gate912(.a(gate489inter0), .b(s_52), .O(gate489inter1));
  and2  gate913(.a(G1241), .b(G1240), .O(gate489inter2));
  inv1  gate914(.a(s_52), .O(gate489inter3));
  inv1  gate915(.a(s_53), .O(gate489inter4));
  nand2 gate916(.a(gate489inter4), .b(gate489inter3), .O(gate489inter5));
  nor2  gate917(.a(gate489inter5), .b(gate489inter2), .O(gate489inter6));
  inv1  gate918(.a(G1240), .O(gate489inter7));
  inv1  gate919(.a(G1241), .O(gate489inter8));
  nand2 gate920(.a(gate489inter8), .b(gate489inter7), .O(gate489inter9));
  nand2 gate921(.a(s_53), .b(gate489inter3), .O(gate489inter10));
  nor2  gate922(.a(gate489inter10), .b(gate489inter9), .O(gate489inter11));
  nor2  gate923(.a(gate489inter11), .b(gate489inter6), .O(gate489inter12));
  nand2 gate924(.a(gate489inter12), .b(gate489inter1), .O(G1298));
nand2 gate490( .a(G1242), .b(G1243), .O(G1299) );

  xor2  gate701(.a(G1245), .b(G1244), .O(gate491inter0));
  nand2 gate702(.a(gate491inter0), .b(s_22), .O(gate491inter1));
  and2  gate703(.a(G1245), .b(G1244), .O(gate491inter2));
  inv1  gate704(.a(s_22), .O(gate491inter3));
  inv1  gate705(.a(s_23), .O(gate491inter4));
  nand2 gate706(.a(gate491inter4), .b(gate491inter3), .O(gate491inter5));
  nor2  gate707(.a(gate491inter5), .b(gate491inter2), .O(gate491inter6));
  inv1  gate708(.a(G1244), .O(gate491inter7));
  inv1  gate709(.a(G1245), .O(gate491inter8));
  nand2 gate710(.a(gate491inter8), .b(gate491inter7), .O(gate491inter9));
  nand2 gate711(.a(s_23), .b(gate491inter3), .O(gate491inter10));
  nor2  gate712(.a(gate491inter10), .b(gate491inter9), .O(gate491inter11));
  nor2  gate713(.a(gate491inter11), .b(gate491inter6), .O(gate491inter12));
  nand2 gate714(.a(gate491inter12), .b(gate491inter1), .O(G1300));
nand2 gate492( .a(G1246), .b(G1247), .O(G1301) );
nand2 gate493( .a(G1248), .b(G1249), .O(G1302) );
nand2 gate494( .a(G1250), .b(G1251), .O(G1303) );
nand2 gate495( .a(G1252), .b(G1253), .O(G1304) );
nand2 gate496( .a(G1254), .b(G1255), .O(G1305) );
nand2 gate497( .a(G1256), .b(G1257), .O(G1306) );
nand2 gate498( .a(G1258), .b(G1259), .O(G1307) );
nand2 gate499( .a(G1260), .b(G1261), .O(G1308) );
nand2 gate500( .a(G1262), .b(G1263), .O(G1309) );

  xor2  gate1359(.a(G1265), .b(G1264), .O(gate501inter0));
  nand2 gate1360(.a(gate501inter0), .b(s_116), .O(gate501inter1));
  and2  gate1361(.a(G1265), .b(G1264), .O(gate501inter2));
  inv1  gate1362(.a(s_116), .O(gate501inter3));
  inv1  gate1363(.a(s_117), .O(gate501inter4));
  nand2 gate1364(.a(gate501inter4), .b(gate501inter3), .O(gate501inter5));
  nor2  gate1365(.a(gate501inter5), .b(gate501inter2), .O(gate501inter6));
  inv1  gate1366(.a(G1264), .O(gate501inter7));
  inv1  gate1367(.a(G1265), .O(gate501inter8));
  nand2 gate1368(.a(gate501inter8), .b(gate501inter7), .O(gate501inter9));
  nand2 gate1369(.a(s_117), .b(gate501inter3), .O(gate501inter10));
  nor2  gate1370(.a(gate501inter10), .b(gate501inter9), .O(gate501inter11));
  nor2  gate1371(.a(gate501inter11), .b(gate501inter6), .O(gate501inter12));
  nand2 gate1372(.a(gate501inter12), .b(gate501inter1), .O(G1310));
nand2 gate502( .a(G1266), .b(G1267), .O(G1311) );
nand2 gate503( .a(G1268), .b(G1269), .O(G1312) );
nand2 gate504( .a(G1270), .b(G1271), .O(G1313) );
nand2 gate505( .a(G1272), .b(G1273), .O(G1314) );
nand2 gate506( .a(G1274), .b(G1275), .O(G1315) );
nand2 gate507( .a(G1276), .b(G1277), .O(G1316) );
nand2 gate508( .a(G1278), .b(G1279), .O(G1317) );
nand2 gate509( .a(G1280), .b(G1281), .O(G1318) );
nand2 gate510( .a(G1282), .b(G1283), .O(G1319) );
nand2 gate511( .a(G1284), .b(G1285), .O(G1320) );
nand2 gate512( .a(G1286), .b(G1287), .O(G1321) );
nand2 gate513( .a(G1288), .b(G1289), .O(G1322) );
nand2 gate514( .a(G1290), .b(G1291), .O(G1323) );
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule