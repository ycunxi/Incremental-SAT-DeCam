module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);

input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;//RE__PI;

input s_0,s_1;//RE__ALLOW(00,01,10,11);
input s_2,s_3;//RE__ALLOW(00,01,10,11);
input s_4,s_5;//RE__ALLOW(00,01,10,11);
input s_6,s_7;//RE__ALLOW(00,01,10,11);
input s_8,s_9;//RE__ALLOW(00,01,10,11);
input s_10,s_11;//RE__ALLOW(00,01,10,11);
input s_12,s_13;//RE__ALLOW(00,01,10,11);
input s_14,s_15;//RE__ALLOW(00,01,10,11);
input s_16,s_17;//RE__ALLOW(00,01,10,11);
input s_18,s_19;//RE__ALLOW(00,01,10,11);
input s_20,s_21;//RE__ALLOW(00,01,10,11);
input s_22,s_23;//RE__ALLOW(00,01,10,11);
input s_24,s_25;//RE__ALLOW(00,01,10,11);
input s_26,s_27;//RE__ALLOW(00,01,10,11);
input s_28,s_29;//RE__ALLOW(00,01,10,11);
input s_30,s_31;//RE__ALLOW(00,01,10,11);
input s_32,s_33;//RE__ALLOW(00,01,10,11);
input s_34,s_35;//RE__ALLOW(00,01,10,11);
input s_36,s_37;//RE__ALLOW(00,01,10,11);
input s_38,s_39;//RE__ALLOW(00,01,10,11);
input s_40,s_41;//RE__ALLOW(00,01,10,11);
input s_42,s_43;//RE__ALLOW(00,01,10,11);
input s_44,s_45;//RE__ALLOW(00,01,10,11);
input s_46,s_47;//RE__ALLOW(00,01,10,11);
input s_48,s_49;//RE__ALLOW(00,01,10,11);
input s_50,s_51;//RE__ALLOW(00,01,10,11);
input s_52,s_53;//RE__ALLOW(00,01,10,11);
input s_54,s_55;//RE__ALLOW(00,01,10,11);
input s_56,s_57;//RE__ALLOW(00,01,10,11);
input s_58,s_59;//RE__ALLOW(00,01,10,11);
input s_60,s_61;//RE__ALLOW(00,01,10,11);
input s_62,s_63;//RE__ALLOW(00,01,10,11);
input s_64,s_65;//RE__ALLOW(00,01,10,11);
input s_66,s_67;//RE__ALLOW(00,01,10,11);
input s_68,s_69;//RE__ALLOW(00,01,10,11);
input s_70,s_71;//RE__ALLOW(00,01,10,11);
input s_72,s_73;//RE__ALLOW(00,01,10,11);
input s_74,s_75;//RE__ALLOW(00,01,10,11);
input s_76,s_77;//RE__ALLOW(00,01,10,11);
input s_78,s_79;//RE__ALLOW(00,01,10,11);
input s_80,s_81;//RE__ALLOW(00,01,10,11);
input s_82,s_83;//RE__ALLOW(00,01,10,11);
input s_84,s_85;//RE__ALLOW(00,01,10,11);
input s_86,s_87;//RE__ALLOW(00,01,10,11);
input s_88,s_89;//RE__ALLOW(00,01,10,11);
input s_90,s_91;//RE__ALLOW(00,01,10,11);
input s_92,s_93;//RE__ALLOW(00,01,10,11);
input s_94,s_95;//RE__ALLOW(00,01,10,11);
input s_96,s_97;//RE__ALLOW(00,01,10,11);
input s_98,s_99;//RE__ALLOW(00,01,10,11);
input s_100,s_101;//RE__ALLOW(00,01,10,11);
input s_102,s_103;//RE__ALLOW(00,01,10,11);
input s_104,s_105;//RE__ALLOW(00,01,10,11);
input s_106,s_107;//RE__ALLOW(00,01,10,11);
input s_108,s_109;//RE__ALLOW(00,01,10,11);
input s_110,s_111;//RE__ALLOW(00,01,10,11);
input s_112,s_113;//RE__ALLOW(00,01,10,11);
input s_114,s_115;//RE__ALLOW(00,01,10,11);
input s_116,s_117;//RE__ALLOW(00,01,10,11);
input s_118,s_119;//RE__ALLOW(00,01,10,11);
input s_120,s_121;//RE__ALLOW(00,01,10,11);
input s_122,s_123;//RE__ALLOW(00,01,10,11);
input s_124,s_125;//RE__ALLOW(00,01,10,11);
input s_126,s_127;//RE__ALLOW(00,01,10,11);
input s_128,s_129;//RE__ALLOW(00,01,10,11);
input s_130,s_131;//RE__ALLOW(00,01,10,11);
input s_132,s_133;//RE__ALLOW(00,01,10,11);
input s_134,s_135;//RE__ALLOW(00,01,10,11);
input s_136,s_137;//RE__ALLOW(00,01,10,11);
input s_138,s_139;//RE__ALLOW(00,01,10,11);
input s_140,s_141;//RE__ALLOW(00,01,10,11);
input s_142,s_143;//RE__ALLOW(00,01,10,11);
input s_144,s_145;//RE__ALLOW(00,01,10,11);
input s_146,s_147;//RE__ALLOW(00,01,10,11);
input s_148,s_149;//RE__ALLOW(00,01,10,11);
input s_150,s_151;//RE__ALLOW(00,01,10,11);
input s_152,s_153;//RE__ALLOW(00,01,10,11);
input s_154,s_155;//RE__ALLOW(00,01,10,11);
input s_156,s_157;//RE__ALLOW(00,01,10,11);
input s_158,s_159;//RE__ALLOW(00,01,10,11);
input s_160,s_161;//RE__ALLOW(00,01,10,11);
input s_162,s_163;//RE__ALLOW(00,01,10,11);
input s_164,s_165;//RE__ALLOW(00,01,10,11);
input s_166,s_167;//RE__ALLOW(00,01,10,11);
input s_168,s_169;//RE__ALLOW(00,01,10,11);
input s_170,s_171;//RE__ALLOW(00,01,10,11);
input s_172,s_173;//RE__ALLOW(00,01,10,11);
input s_174,s_175;//RE__ALLOW(00,01,10,11);
input s_176,s_177;//RE__ALLOW(00,01,10,11);
input s_178,s_179;//RE__ALLOW(00,01,10,11);
input s_180,s_181;//RE__ALLOW(00,01,10,11);
input s_182,s_183;//RE__ALLOW(00,01,10,11);
input s_184,s_185;//RE__ALLOW(00,01,10,11);
input s_186,s_187;//RE__ALLOW(00,01,10,11);
input s_188,s_189;//RE__ALLOW(00,01,10,11);
input s_190,s_191;//RE__ALLOW(00,01,10,11);
input s_192,s_193;//RE__ALLOW(00,01,10,11);
input s_194,s_195;//RE__ALLOW(00,01,10,11);
input s_196,s_197;//RE__ALLOW(00,01,10,11);
input s_198,s_199;//RE__ALLOW(00,01,10,11);
input s_200,s_201;//RE__ALLOW(00,01,10,11);
input s_202,s_203;//RE__ALLOW(00,01,10,11);
input s_204,s_205;//RE__ALLOW(00,01,10,11);
input s_206,s_207;//RE__ALLOW(00,01,10,11);
input s_208,s_209;//RE__ALLOW(00,01,10,11);
input s_210,s_211;//RE__ALLOW(00,01,10,11);
input s_212,s_213;//RE__ALLOW(00,01,10,11);
input s_214,s_215;//RE__ALLOW(00,01,10,11);
input s_216,s_217;//RE__ALLOW(00,01,10,11);
input s_218,s_219;//RE__ALLOW(00,01,10,11);
input s_220,s_221;//RE__ALLOW(00,01,10,11);
input s_222,s_223;//RE__ALLOW(00,01,10,11);
input s_224,s_225;//RE__ALLOW(00,01,10,11);
input s_226,s_227;//RE__ALLOW(00,01,10,11);
input s_228,s_229;//RE__ALLOW(00,01,10,11);
input s_230,s_231;//RE__ALLOW(00,01,10,11);
input s_232,s_233;//RE__ALLOW(00,01,10,11);
input s_234,s_235;//RE__ALLOW(00,01,10,11);
input s_236,s_237;//RE__ALLOW(00,01,10,11);
input s_238,s_239;//RE__ALLOW(00,01,10,11);
input s_240,s_241;//RE__ALLOW(00,01,10,11);
input s_242,s_243;//RE__ALLOW(00,01,10,11);
input s_244,s_245;//RE__ALLOW(00,01,10,11);
input s_246,s_247;//RE__ALLOW(00,01,10,11);
input s_248,s_249;//RE__ALLOW(00,01,10,11);
input s_250,s_251;//RE__ALLOW(00,01,10,11);
input s_252,s_253;//RE__ALLOW(00,01,10,11);
input s_254,s_255;//RE__ALLOW(00,01,10,11);
input s_256,s_257;//RE__ALLOW(00,01,10,11);
input s_258,s_259;//RE__ALLOW(00,01,10,11);
input s_260,s_261;//RE__ALLOW(00,01,10,11);
input s_262,s_263;//RE__ALLOW(00,01,10,11);
input s_264,s_265;//RE__ALLOW(00,01,10,11);
input s_266,s_267;//RE__ALLOW(00,01,10,11);
input s_268,s_269;//RE__ALLOW(00,01,10,11);
input s_270,s_271;//RE__ALLOW(00,01,10,11);
input s_272,s_273;//RE__ALLOW(00,01,10,11);
input s_274,s_275;//RE__ALLOW(00,01,10,11);
input s_276,s_277;//RE__ALLOW(00,01,10,11);
input s_278,s_279;//RE__ALLOW(00,01,10,11);
input s_280,s_281;//RE__ALLOW(00,01,10,11);
input s_282,s_283;//RE__ALLOW(00,01,10,11);
input s_284,s_285;//RE__ALLOW(00,01,10,11);
input s_286,s_287;//RE__ALLOW(00,01,10,11);
input s_288,s_289;//RE__ALLOW(00,01,10,11);
input s_290,s_291;//RE__ALLOW(00,01,10,11);
input s_292,s_293;//RE__ALLOW(00,01,10,11);
input s_294,s_295;//RE__ALLOW(00,01,10,11);
input s_296,s_297;//RE__ALLOW(00,01,10,11);
input s_298,s_299;//RE__ALLOW(00,01,10,11);
input s_300,s_301;//RE__ALLOW(00,01,10,11);
input s_302,s_303;//RE__ALLOW(00,01,10,11);
input s_304,s_305;//RE__ALLOW(00,01,10,11);
input s_306,s_307;//RE__ALLOW(00,01,10,11);
input s_308,s_309;//RE__ALLOW(00,01,10,11);
input s_310,s_311;//RE__ALLOW(00,01,10,11);
input s_312,s_313;//RE__ALLOW(00,01,10,11);
input s_314,s_315;//RE__ALLOW(00,01,10,11);
input s_316,s_317;//RE__ALLOW(00,01,10,11);
input s_318,s_319;//RE__ALLOW(00,01,10,11);
input s_320,s_321;//RE__ALLOW(00,01,10,11);
input s_322,s_323;//RE__ALLOW(00,01,10,11);
input s_324,s_325;//RE__ALLOW(00,01,10,11);
input s_326,s_327;//RE__ALLOW(00,01,10,11);
input s_328,s_329;//RE__ALLOW(00,01,10,11);
input s_330,s_331;//RE__ALLOW(00,01,10,11);
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;

  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate157inter0, gate157inter1, gate157inter2, gate157inter3, gate157inter4, gate157inter5, gate157inter6, gate157inter7, gate157inter8, gate157inter9, gate157inter10, gate157inter11, gate157inter12, gate250inter0, gate250inter1, gate250inter2, gate250inter3, gate250inter4, gate250inter5, gate250inter6, gate250inter7, gate250inter8, gate250inter9, gate250inter10, gate250inter11, gate250inter12, gate253inter0, gate253inter1, gate253inter2, gate253inter3, gate253inter4, gate253inter5, gate253inter6, gate253inter7, gate253inter8, gate253inter9, gate253inter10, gate253inter11, gate253inter12, gate251inter0, gate251inter1, gate251inter2, gate251inter3, gate251inter4, gate251inter5, gate251inter6, gate251inter7, gate251inter8, gate251inter9, gate251inter10, gate251inter11, gate251inter12, gate52inter0, gate52inter1, gate52inter2, gate52inter3, gate52inter4, gate52inter5, gate52inter6, gate52inter7, gate52inter8, gate52inter9, gate52inter10, gate52inter11, gate52inter12, gate509inter0, gate509inter1, gate509inter2, gate509inter3, gate509inter4, gate509inter5, gate509inter6, gate509inter7, gate509inter8, gate509inter9, gate509inter10, gate509inter11, gate509inter12, gate274inter0, gate274inter1, gate274inter2, gate274inter3, gate274inter4, gate274inter5, gate274inter6, gate274inter7, gate274inter8, gate274inter9, gate274inter10, gate274inter11, gate274inter12, gate56inter0, gate56inter1, gate56inter2, gate56inter3, gate56inter4, gate56inter5, gate56inter6, gate56inter7, gate56inter8, gate56inter9, gate56inter10, gate56inter11, gate56inter12, gate139inter0, gate139inter1, gate139inter2, gate139inter3, gate139inter4, gate139inter5, gate139inter6, gate139inter7, gate139inter8, gate139inter9, gate139inter10, gate139inter11, gate139inter12, gate208inter0, gate208inter1, gate208inter2, gate208inter3, gate208inter4, gate208inter5, gate208inter6, gate208inter7, gate208inter8, gate208inter9, gate208inter10, gate208inter11, gate208inter12, gate158inter0, gate158inter1, gate158inter2, gate158inter3, gate158inter4, gate158inter5, gate158inter6, gate158inter7, gate158inter8, gate158inter9, gate158inter10, gate158inter11, gate158inter12, gate287inter0, gate287inter1, gate287inter2, gate287inter3, gate287inter4, gate287inter5, gate287inter6, gate287inter7, gate287inter8, gate287inter9, gate287inter10, gate287inter11, gate287inter12, gate437inter0, gate437inter1, gate437inter2, gate437inter3, gate437inter4, gate437inter5, gate437inter6, gate437inter7, gate437inter8, gate437inter9, gate437inter10, gate437inter11, gate437inter12, gate74inter0, gate74inter1, gate74inter2, gate74inter3, gate74inter4, gate74inter5, gate74inter6, gate74inter7, gate74inter8, gate74inter9, gate74inter10, gate74inter11, gate74inter12, gate249inter0, gate249inter1, gate249inter2, gate249inter3, gate249inter4, gate249inter5, gate249inter6, gate249inter7, gate249inter8, gate249inter9, gate249inter10, gate249inter11, gate249inter12, gate43inter0, gate43inter1, gate43inter2, gate43inter3, gate43inter4, gate43inter5, gate43inter6, gate43inter7, gate43inter8, gate43inter9, gate43inter10, gate43inter11, gate43inter12, gate278inter0, gate278inter1, gate278inter2, gate278inter3, gate278inter4, gate278inter5, gate278inter6, gate278inter7, gate278inter8, gate278inter9, gate278inter10, gate278inter11, gate278inter12, gate484inter0, gate484inter1, gate484inter2, gate484inter3, gate484inter4, gate484inter5, gate484inter6, gate484inter7, gate484inter8, gate484inter9, gate484inter10, gate484inter11, gate484inter12, gate210inter0, gate210inter1, gate210inter2, gate210inter3, gate210inter4, gate210inter5, gate210inter6, gate210inter7, gate210inter8, gate210inter9, gate210inter10, gate210inter11, gate210inter12, gate54inter0, gate54inter1, gate54inter2, gate54inter3, gate54inter4, gate54inter5, gate54inter6, gate54inter7, gate54inter8, gate54inter9, gate54inter10, gate54inter11, gate54inter12, gate99inter0, gate99inter1, gate99inter2, gate99inter3, gate99inter4, gate99inter5, gate99inter6, gate99inter7, gate99inter8, gate99inter9, gate99inter10, gate99inter11, gate99inter12, gate115inter0, gate115inter1, gate115inter2, gate115inter3, gate115inter4, gate115inter5, gate115inter6, gate115inter7, gate115inter8, gate115inter9, gate115inter10, gate115inter11, gate115inter12, gate15inter0, gate15inter1, gate15inter2, gate15inter3, gate15inter4, gate15inter5, gate15inter6, gate15inter7, gate15inter8, gate15inter9, gate15inter10, gate15inter11, gate15inter12, gate235inter0, gate235inter1, gate235inter2, gate235inter3, gate235inter4, gate235inter5, gate235inter6, gate235inter7, gate235inter8, gate235inter9, gate235inter10, gate235inter11, gate235inter12, gate282inter0, gate282inter1, gate282inter2, gate282inter3, gate282inter4, gate282inter5, gate282inter6, gate282inter7, gate282inter8, gate282inter9, gate282inter10, gate282inter11, gate282inter12, gate173inter0, gate173inter1, gate173inter2, gate173inter3, gate173inter4, gate173inter5, gate173inter6, gate173inter7, gate173inter8, gate173inter9, gate173inter10, gate173inter11, gate173inter12, gate244inter0, gate244inter1, gate244inter2, gate244inter3, gate244inter4, gate244inter5, gate244inter6, gate244inter7, gate244inter8, gate244inter9, gate244inter10, gate244inter11, gate244inter12, gate119inter0, gate119inter1, gate119inter2, gate119inter3, gate119inter4, gate119inter5, gate119inter6, gate119inter7, gate119inter8, gate119inter9, gate119inter10, gate119inter11, gate119inter12, gate438inter0, gate438inter1, gate438inter2, gate438inter3, gate438inter4, gate438inter5, gate438inter6, gate438inter7, gate438inter8, gate438inter9, gate438inter10, gate438inter11, gate438inter12, gate492inter0, gate492inter1, gate492inter2, gate492inter3, gate492inter4, gate492inter5, gate492inter6, gate492inter7, gate492inter8, gate492inter9, gate492inter10, gate492inter11, gate492inter12, gate36inter0, gate36inter1, gate36inter2, gate36inter3, gate36inter4, gate36inter5, gate36inter6, gate36inter7, gate36inter8, gate36inter9, gate36inter10, gate36inter11, gate36inter12, gate432inter0, gate432inter1, gate432inter2, gate432inter3, gate432inter4, gate432inter5, gate432inter6, gate432inter7, gate432inter8, gate432inter9, gate432inter10, gate432inter11, gate432inter12, gate156inter0, gate156inter1, gate156inter2, gate156inter3, gate156inter4, gate156inter5, gate156inter6, gate156inter7, gate156inter8, gate156inter9, gate156inter10, gate156inter11, gate156inter12, gate186inter0, gate186inter1, gate186inter2, gate186inter3, gate186inter4, gate186inter5, gate186inter6, gate186inter7, gate186inter8, gate186inter9, gate186inter10, gate186inter11, gate186inter12, gate399inter0, gate399inter1, gate399inter2, gate399inter3, gate399inter4, gate399inter5, gate399inter6, gate399inter7, gate399inter8, gate399inter9, gate399inter10, gate399inter11, gate399inter12, gate290inter0, gate290inter1, gate290inter2, gate290inter3, gate290inter4, gate290inter5, gate290inter6, gate290inter7, gate290inter8, gate290inter9, gate290inter10, gate290inter11, gate290inter12, gate394inter0, gate394inter1, gate394inter2, gate394inter3, gate394inter4, gate394inter5, gate394inter6, gate394inter7, gate394inter8, gate394inter9, gate394inter10, gate394inter11, gate394inter12, gate264inter0, gate264inter1, gate264inter2, gate264inter3, gate264inter4, gate264inter5, gate264inter6, gate264inter7, gate264inter8, gate264inter9, gate264inter10, gate264inter11, gate264inter12, gate184inter0, gate184inter1, gate184inter2, gate184inter3, gate184inter4, gate184inter5, gate184inter6, gate184inter7, gate184inter8, gate184inter9, gate184inter10, gate184inter11, gate184inter12, gate198inter0, gate198inter1, gate198inter2, gate198inter3, gate198inter4, gate198inter5, gate198inter6, gate198inter7, gate198inter8, gate198inter9, gate198inter10, gate198inter11, gate198inter12, gate197inter0, gate197inter1, gate197inter2, gate197inter3, gate197inter4, gate197inter5, gate197inter6, gate197inter7, gate197inter8, gate197inter9, gate197inter10, gate197inter11, gate197inter12, gate387inter0, gate387inter1, gate387inter2, gate387inter3, gate387inter4, gate387inter5, gate387inter6, gate387inter7, gate387inter8, gate387inter9, gate387inter10, gate387inter11, gate387inter12, gate150inter0, gate150inter1, gate150inter2, gate150inter3, gate150inter4, gate150inter5, gate150inter6, gate150inter7, gate150inter8, gate150inter9, gate150inter10, gate150inter11, gate150inter12, gate68inter0, gate68inter1, gate68inter2, gate68inter3, gate68inter4, gate68inter5, gate68inter6, gate68inter7, gate68inter8, gate68inter9, gate68inter10, gate68inter11, gate68inter12, gate147inter0, gate147inter1, gate147inter2, gate147inter3, gate147inter4, gate147inter5, gate147inter6, gate147inter7, gate147inter8, gate147inter9, gate147inter10, gate147inter11, gate147inter12, gate86inter0, gate86inter1, gate86inter2, gate86inter3, gate86inter4, gate86inter5, gate86inter6, gate86inter7, gate86inter8, gate86inter9, gate86inter10, gate86inter11, gate86inter12, gate407inter0, gate407inter1, gate407inter2, gate407inter3, gate407inter4, gate407inter5, gate407inter6, gate407inter7, gate407inter8, gate407inter9, gate407inter10, gate407inter11, gate407inter12, gate151inter0, gate151inter1, gate151inter2, gate151inter3, gate151inter4, gate151inter5, gate151inter6, gate151inter7, gate151inter8, gate151inter9, gate151inter10, gate151inter11, gate151inter12, gate72inter0, gate72inter1, gate72inter2, gate72inter3, gate72inter4, gate72inter5, gate72inter6, gate72inter7, gate72inter8, gate72inter9, gate72inter10, gate72inter11, gate72inter12, gate227inter0, gate227inter1, gate227inter2, gate227inter3, gate227inter4, gate227inter5, gate227inter6, gate227inter7, gate227inter8, gate227inter9, gate227inter10, gate227inter11, gate227inter12, gate502inter0, gate502inter1, gate502inter2, gate502inter3, gate502inter4, gate502inter5, gate502inter6, gate502inter7, gate502inter8, gate502inter9, gate502inter10, gate502inter11, gate502inter12, gate160inter0, gate160inter1, gate160inter2, gate160inter3, gate160inter4, gate160inter5, gate160inter6, gate160inter7, gate160inter8, gate160inter9, gate160inter10, gate160inter11, gate160inter12, gate16inter0, gate16inter1, gate16inter2, gate16inter3, gate16inter4, gate16inter5, gate16inter6, gate16inter7, gate16inter8, gate16inter9, gate16inter10, gate16inter11, gate16inter12, gate391inter0, gate391inter1, gate391inter2, gate391inter3, gate391inter4, gate391inter5, gate391inter6, gate391inter7, gate391inter8, gate391inter9, gate391inter10, gate391inter11, gate391inter12, gate196inter0, gate196inter1, gate196inter2, gate196inter3, gate196inter4, gate196inter5, gate196inter6, gate196inter7, gate196inter8, gate196inter9, gate196inter10, gate196inter11, gate196inter12, gate225inter0, gate225inter1, gate225inter2, gate225inter3, gate225inter4, gate225inter5, gate225inter6, gate225inter7, gate225inter8, gate225inter9, gate225inter10, gate225inter11, gate225inter12, gate109inter0, gate109inter1, gate109inter2, gate109inter3, gate109inter4, gate109inter5, gate109inter6, gate109inter7, gate109inter8, gate109inter9, gate109inter10, gate109inter11, gate109inter12, gate285inter0, gate285inter1, gate285inter2, gate285inter3, gate285inter4, gate285inter5, gate285inter6, gate285inter7, gate285inter8, gate285inter9, gate285inter10, gate285inter11, gate285inter12, gate258inter0, gate258inter1, gate258inter2, gate258inter3, gate258inter4, gate258inter5, gate258inter6, gate258inter7, gate258inter8, gate258inter9, gate258inter10, gate258inter11, gate258inter12, gate118inter0, gate118inter1, gate118inter2, gate118inter3, gate118inter4, gate118inter5, gate118inter6, gate118inter7, gate118inter8, gate118inter9, gate118inter10, gate118inter11, gate118inter12, gate286inter0, gate286inter1, gate286inter2, gate286inter3, gate286inter4, gate286inter5, gate286inter6, gate286inter7, gate286inter8, gate286inter9, gate286inter10, gate286inter11, gate286inter12, gate94inter0, gate94inter1, gate94inter2, gate94inter3, gate94inter4, gate94inter5, gate94inter6, gate94inter7, gate94inter8, gate94inter9, gate94inter10, gate94inter11, gate94inter12, gate76inter0, gate76inter1, gate76inter2, gate76inter3, gate76inter4, gate76inter5, gate76inter6, gate76inter7, gate76inter8, gate76inter9, gate76inter10, gate76inter11, gate76inter12, gate257inter0, gate257inter1, gate257inter2, gate257inter3, gate257inter4, gate257inter5, gate257inter6, gate257inter7, gate257inter8, gate257inter9, gate257inter10, gate257inter11, gate257inter12, gate134inter0, gate134inter1, gate134inter2, gate134inter3, gate134inter4, gate134inter5, gate134inter6, gate134inter7, gate134inter8, gate134inter9, gate134inter10, gate134inter11, gate134inter12, gate429inter0, gate429inter1, gate429inter2, gate429inter3, gate429inter4, gate429inter5, gate429inter6, gate429inter7, gate429inter8, gate429inter9, gate429inter10, gate429inter11, gate429inter12, gate460inter0, gate460inter1, gate460inter2, gate460inter3, gate460inter4, gate460inter5, gate460inter6, gate460inter7, gate460inter8, gate460inter9, gate460inter10, gate460inter11, gate460inter12, gate451inter0, gate451inter1, gate451inter2, gate451inter3, gate451inter4, gate451inter5, gate451inter6, gate451inter7, gate451inter8, gate451inter9, gate451inter10, gate451inter11, gate451inter12, gate265inter0, gate265inter1, gate265inter2, gate265inter3, gate265inter4, gate265inter5, gate265inter6, gate265inter7, gate265inter8, gate265inter9, gate265inter10, gate265inter11, gate265inter12, gate155inter0, gate155inter1, gate155inter2, gate155inter3, gate155inter4, gate155inter5, gate155inter6, gate155inter7, gate155inter8, gate155inter9, gate155inter10, gate155inter11, gate155inter12, gate229inter0, gate229inter1, gate229inter2, gate229inter3, gate229inter4, gate229inter5, gate229inter6, gate229inter7, gate229inter8, gate229inter9, gate229inter10, gate229inter11, gate229inter12, gate398inter0, gate398inter1, gate398inter2, gate398inter3, gate398inter4, gate398inter5, gate398inter6, gate398inter7, gate398inter8, gate398inter9, gate398inter10, gate398inter11, gate398inter12, gate14inter0, gate14inter1, gate14inter2, gate14inter3, gate14inter4, gate14inter5, gate14inter6, gate14inter7, gate14inter8, gate14inter9, gate14inter10, gate14inter11, gate14inter12, gate462inter0, gate462inter1, gate462inter2, gate462inter3, gate462inter4, gate462inter5, gate462inter6, gate462inter7, gate462inter8, gate462inter9, gate462inter10, gate462inter11, gate462inter12, gate110inter0, gate110inter1, gate110inter2, gate110inter3, gate110inter4, gate110inter5, gate110inter6, gate110inter7, gate110inter8, gate110inter9, gate110inter10, gate110inter11, gate110inter12, gate167inter0, gate167inter1, gate167inter2, gate167inter3, gate167inter4, gate167inter5, gate167inter6, gate167inter7, gate167inter8, gate167inter9, gate167inter10, gate167inter11, gate167inter12, gate203inter0, gate203inter1, gate203inter2, gate203inter3, gate203inter4, gate203inter5, gate203inter6, gate203inter7, gate203inter8, gate203inter9, gate203inter10, gate203inter11, gate203inter12, gate488inter0, gate488inter1, gate488inter2, gate488inter3, gate488inter4, gate488inter5, gate488inter6, gate488inter7, gate488inter8, gate488inter9, gate488inter10, gate488inter11, gate488inter12, gate269inter0, gate269inter1, gate269inter2, gate269inter3, gate269inter4, gate269inter5, gate269inter6, gate269inter7, gate269inter8, gate269inter9, gate269inter10, gate269inter11, gate269inter12, gate165inter0, gate165inter1, gate165inter2, gate165inter3, gate165inter4, gate165inter5, gate165inter6, gate165inter7, gate165inter8, gate165inter9, gate165inter10, gate165inter11, gate165inter12, gate279inter0, gate279inter1, gate279inter2, gate279inter3, gate279inter4, gate279inter5, gate279inter6, gate279inter7, gate279inter8, gate279inter9, gate279inter10, gate279inter11, gate279inter12, gate93inter0, gate93inter1, gate93inter2, gate93inter3, gate93inter4, gate93inter5, gate93inter6, gate93inter7, gate93inter8, gate93inter9, gate93inter10, gate93inter11, gate93inter12, gate58inter0, gate58inter1, gate58inter2, gate58inter3, gate58inter4, gate58inter5, gate58inter6, gate58inter7, gate58inter8, gate58inter9, gate58inter10, gate58inter11, gate58inter12, gate388inter0, gate388inter1, gate388inter2, gate388inter3, gate388inter4, gate388inter5, gate388inter6, gate388inter7, gate388inter8, gate388inter9, gate388inter10, gate388inter11, gate388inter12, gate159inter0, gate159inter1, gate159inter2, gate159inter3, gate159inter4, gate159inter5, gate159inter6, gate159inter7, gate159inter8, gate159inter9, gate159inter10, gate159inter11, gate159inter12, gate446inter0, gate446inter1, gate446inter2, gate446inter3, gate446inter4, gate446inter5, gate446inter6, gate446inter7, gate446inter8, gate446inter9, gate446inter10, gate446inter11, gate446inter12, gate105inter0, gate105inter1, gate105inter2, gate105inter3, gate105inter4, gate105inter5, gate105inter6, gate105inter7, gate105inter8, gate105inter9, gate105inter10, gate105inter11, gate105inter12, gate500inter0, gate500inter1, gate500inter2, gate500inter3, gate500inter4, gate500inter5, gate500inter6, gate500inter7, gate500inter8, gate500inter9, gate500inter10, gate500inter11, gate500inter12, gate396inter0, gate396inter1, gate396inter2, gate396inter3, gate396inter4, gate396inter5, gate396inter6, gate396inter7, gate396inter8, gate396inter9, gate396inter10, gate396inter11, gate396inter12, gate27inter0, gate27inter1, gate27inter2, gate27inter3, gate27inter4, gate27inter5, gate27inter6, gate27inter7, gate27inter8, gate27inter9, gate27inter10, gate27inter11, gate27inter12, gate271inter0, gate271inter1, gate271inter2, gate271inter3, gate271inter4, gate271inter5, gate271inter6, gate271inter7, gate271inter8, gate271inter9, gate271inter10, gate271inter11, gate271inter12, gate392inter0, gate392inter1, gate392inter2, gate392inter3, gate392inter4, gate392inter5, gate392inter6, gate392inter7, gate392inter8, gate392inter9, gate392inter10, gate392inter11, gate392inter12, gate277inter0, gate277inter1, gate277inter2, gate277inter3, gate277inter4, gate277inter5, gate277inter6, gate277inter7, gate277inter8, gate277inter9, gate277inter10, gate277inter11, gate277inter12, gate205inter0, gate205inter1, gate205inter2, gate205inter3, gate205inter4, gate205inter5, gate205inter6, gate205inter7, gate205inter8, gate205inter9, gate205inter10, gate205inter11, gate205inter12, gate226inter0, gate226inter1, gate226inter2, gate226inter3, gate226inter4, gate226inter5, gate226inter6, gate226inter7, gate226inter8, gate226inter9, gate226inter10, gate226inter11, gate226inter12, gate132inter0, gate132inter1, gate132inter2, gate132inter3, gate132inter4, gate132inter5, gate132inter6, gate132inter7, gate132inter8, gate132inter9, gate132inter10, gate132inter11, gate132inter12, gate19inter0, gate19inter1, gate19inter2, gate19inter3, gate19inter4, gate19inter5, gate19inter6, gate19inter7, gate19inter8, gate19inter9, gate19inter10, gate19inter11, gate19inter12, gate493inter0, gate493inter1, gate493inter2, gate493inter3, gate493inter4, gate493inter5, gate493inter6, gate493inter7, gate493inter8, gate493inter9, gate493inter10, gate493inter11, gate493inter12, gate34inter0, gate34inter1, gate34inter2, gate34inter3, gate34inter4, gate34inter5, gate34inter6, gate34inter7, gate34inter8, gate34inter9, gate34inter10, gate34inter11, gate34inter12, gate237inter0, gate237inter1, gate237inter2, gate237inter3, gate237inter4, gate237inter5, gate237inter6, gate237inter7, gate237inter8, gate237inter9, gate237inter10, gate237inter11, gate237inter12, gate107inter0, gate107inter1, gate107inter2, gate107inter3, gate107inter4, gate107inter5, gate107inter6, gate107inter7, gate107inter8, gate107inter9, gate107inter10, gate107inter11, gate107inter12, gate45inter0, gate45inter1, gate45inter2, gate45inter3, gate45inter4, gate45inter5, gate45inter6, gate45inter7, gate45inter8, gate45inter9, gate45inter10, gate45inter11, gate45inter12, gate22inter0, gate22inter1, gate22inter2, gate22inter3, gate22inter4, gate22inter5, gate22inter6, gate22inter7, gate22inter8, gate22inter9, gate22inter10, gate22inter11, gate22inter12, gate48inter0, gate48inter1, gate48inter2, gate48inter3, gate48inter4, gate48inter5, gate48inter6, gate48inter7, gate48inter8, gate48inter9, gate48inter10, gate48inter11, gate48inter12, gate31inter0, gate31inter1, gate31inter2, gate31inter3, gate31inter4, gate31inter5, gate31inter6, gate31inter7, gate31inter8, gate31inter9, gate31inter10, gate31inter11, gate31inter12, gate267inter0, gate267inter1, gate267inter2, gate267inter3, gate267inter4, gate267inter5, gate267inter6, gate267inter7, gate267inter8, gate267inter9, gate267inter10, gate267inter11, gate267inter12, gate473inter0, gate473inter1, gate473inter2, gate473inter3, gate473inter4, gate473inter5, gate473inter6, gate473inter7, gate473inter8, gate473inter9, gate473inter10, gate473inter11, gate473inter12, gate106inter0, gate106inter1, gate106inter2, gate106inter3, gate106inter4, gate106inter5, gate106inter6, gate106inter7, gate106inter8, gate106inter9, gate106inter10, gate106inter11, gate106inter12, gate474inter0, gate474inter1, gate474inter2, gate474inter3, gate474inter4, gate474inter5, gate474inter6, gate474inter7, gate474inter8, gate474inter9, gate474inter10, gate474inter11, gate474inter12, gate292inter0, gate292inter1, gate292inter2, gate292inter3, gate292inter4, gate292inter5, gate292inter6, gate292inter7, gate292inter8, gate292inter9, gate292inter10, gate292inter11, gate292inter12, gate255inter0, gate255inter1, gate255inter2, gate255inter3, gate255inter4, gate255inter5, gate255inter6, gate255inter7, gate255inter8, gate255inter9, gate255inter10, gate255inter11, gate255inter12, gate87inter0, gate87inter1, gate87inter2, gate87inter3, gate87inter4, gate87inter5, gate87inter6, gate87inter7, gate87inter8, gate87inter9, gate87inter10, gate87inter11, gate87inter12, gate472inter0, gate472inter1, gate472inter2, gate472inter3, gate472inter4, gate472inter5, gate472inter6, gate472inter7, gate472inter8, gate472inter9, gate472inter10, gate472inter11, gate472inter12, gate92inter0, gate92inter1, gate92inter2, gate92inter3, gate92inter4, gate92inter5, gate92inter6, gate92inter7, gate92inter8, gate92inter9, gate92inter10, gate92inter11, gate92inter12, gate400inter0, gate400inter1, gate400inter2, gate400inter3, gate400inter4, gate400inter5, gate400inter6, gate400inter7, gate400inter8, gate400inter9, gate400inter10, gate400inter11, gate400inter12, gate57inter0, gate57inter1, gate57inter2, gate57inter3, gate57inter4, gate57inter5, gate57inter6, gate57inter7, gate57inter8, gate57inter9, gate57inter10, gate57inter11, gate57inter12, gate448inter0, gate448inter1, gate448inter2, gate448inter3, gate448inter4, gate448inter5, gate448inter6, gate448inter7, gate448inter8, gate448inter9, gate448inter10, gate448inter11, gate448inter12, gate195inter0, gate195inter1, gate195inter2, gate195inter3, gate195inter4, gate195inter5, gate195inter6, gate195inter7, gate195inter8, gate195inter9, gate195inter10, gate195inter11, gate195inter12, gate138inter0, gate138inter1, gate138inter2, gate138inter3, gate138inter4, gate138inter5, gate138inter6, gate138inter7, gate138inter8, gate138inter9, gate138inter10, gate138inter11, gate138inter12, gate133inter0, gate133inter1, gate133inter2, gate133inter3, gate133inter4, gate133inter5, gate133inter6, gate133inter7, gate133inter8, gate133inter9, gate133inter10, gate133inter11, gate133inter12, gate44inter0, gate44inter1, gate44inter2, gate44inter3, gate44inter4, gate44inter5, gate44inter6, gate44inter7, gate44inter8, gate44inter9, gate44inter10, gate44inter11, gate44inter12, gate79inter0, gate79inter1, gate79inter2, gate79inter3, gate79inter4, gate79inter5, gate79inter6, gate79inter7, gate79inter8, gate79inter9, gate79inter10, gate79inter11, gate79inter12, gate137inter0, gate137inter1, gate137inter2, gate137inter3, gate137inter4, gate137inter5, gate137inter6, gate137inter7, gate137inter8, gate137inter9, gate137inter10, gate137inter11, gate137inter12, gate256inter0, gate256inter1, gate256inter2, gate256inter3, gate256inter4, gate256inter5, gate256inter6, gate256inter7, gate256inter8, gate256inter9, gate256inter10, gate256inter11, gate256inter12, gate180inter0, gate180inter1, gate180inter2, gate180inter3, gate180inter4, gate180inter5, gate180inter6, gate180inter7, gate180inter8, gate180inter9, gate180inter10, gate180inter11, gate180inter12, gate475inter0, gate475inter1, gate475inter2, gate475inter3, gate475inter4, gate475inter5, gate475inter6, gate475inter7, gate475inter8, gate475inter9, gate475inter10, gate475inter11, gate475inter12, gate491inter0, gate491inter1, gate491inter2, gate491inter3, gate491inter4, gate491inter5, gate491inter6, gate491inter7, gate491inter8, gate491inter9, gate491inter10, gate491inter11, gate491inter12, gate506inter0, gate506inter1, gate506inter2, gate506inter3, gate506inter4, gate506inter5, gate506inter6, gate506inter7, gate506inter8, gate506inter9, gate506inter10, gate506inter11, gate506inter12, gate427inter0, gate427inter1, gate427inter2, gate427inter3, gate427inter4, gate427inter5, gate427inter6, gate427inter7, gate427inter8, gate427inter9, gate427inter10, gate427inter11, gate427inter12, gate463inter0, gate463inter1, gate463inter2, gate463inter3, gate463inter4, gate463inter5, gate463inter6, gate463inter7, gate463inter8, gate463inter9, gate463inter10, gate463inter11, gate463inter12, gate422inter0, gate422inter1, gate422inter2, gate422inter3, gate422inter4, gate422inter5, gate422inter6, gate422inter7, gate422inter8, gate422inter9, gate422inter10, gate422inter11, gate422inter12, gate454inter0, gate454inter1, gate454inter2, gate454inter3, gate454inter4, gate454inter5, gate454inter6, gate454inter7, gate454inter8, gate454inter9, gate454inter10, gate454inter11, gate454inter12, gate91inter0, gate91inter1, gate91inter2, gate91inter3, gate91inter4, gate91inter5, gate91inter6, gate91inter7, gate91inter8, gate91inter9, gate91inter10, gate91inter11, gate91inter12, gate490inter0, gate490inter1, gate490inter2, gate490inter3, gate490inter4, gate490inter5, gate490inter6, gate490inter7, gate490inter8, gate490inter9, gate490inter10, gate490inter11, gate490inter12, gate202inter0, gate202inter1, gate202inter2, gate202inter3, gate202inter4, gate202inter5, gate202inter6, gate202inter7, gate202inter8, gate202inter9, gate202inter10, gate202inter11, gate202inter12, gate104inter0, gate104inter1, gate104inter2, gate104inter3, gate104inter4, gate104inter5, gate104inter6, gate104inter7, gate104inter8, gate104inter9, gate104inter10, gate104inter11, gate104inter12, gate55inter0, gate55inter1, gate55inter2, gate55inter3, gate55inter4, gate55inter5, gate55inter6, gate55inter7, gate55inter8, gate55inter9, gate55inter10, gate55inter11, gate55inter12, gate445inter0, gate445inter1, gate445inter2, gate445inter3, gate445inter4, gate445inter5, gate445inter6, gate445inter7, gate445inter8, gate445inter9, gate445inter10, gate445inter11, gate445inter12, gate224inter0, gate224inter1, gate224inter2, gate224inter3, gate224inter4, gate224inter5, gate224inter6, gate224inter7, gate224inter8, gate224inter9, gate224inter10, gate224inter11, gate224inter12, gate485inter0, gate485inter1, gate485inter2, gate485inter3, gate485inter4, gate485inter5, gate485inter6, gate485inter7, gate485inter8, gate485inter9, gate485inter10, gate485inter11, gate485inter12, gate442inter0, gate442inter1, gate442inter2, gate442inter3, gate442inter4, gate442inter5, gate442inter6, gate442inter7, gate442inter8, gate442inter9, gate442inter10, gate442inter11, gate442inter12, gate245inter0, gate245inter1, gate245inter2, gate245inter3, gate245inter4, gate245inter5, gate245inter6, gate245inter7, gate245inter8, gate245inter9, gate245inter10, gate245inter11, gate245inter12, gate281inter0, gate281inter1, gate281inter2, gate281inter3, gate281inter4, gate281inter5, gate281inter6, gate281inter7, gate281inter8, gate281inter9, gate281inter10, gate281inter11, gate281inter12, gate414inter0, gate414inter1, gate414inter2, gate414inter3, gate414inter4, gate414inter5, gate414inter6, gate414inter7, gate414inter8, gate414inter9, gate414inter10, gate414inter11, gate414inter12, gate97inter0, gate97inter1, gate97inter2, gate97inter3, gate97inter4, gate97inter5, gate97inter6, gate97inter7, gate97inter8, gate97inter9, gate97inter10, gate97inter11, gate97inter12, gate468inter0, gate468inter1, gate468inter2, gate468inter3, gate468inter4, gate468inter5, gate468inter6, gate468inter7, gate468inter8, gate468inter9, gate468inter10, gate468inter11, gate468inter12, gate144inter0, gate144inter1, gate144inter2, gate144inter3, gate144inter4, gate144inter5, gate144inter6, gate144inter7, gate144inter8, gate144inter9, gate144inter10, gate144inter11, gate144inter12, gate199inter0, gate199inter1, gate199inter2, gate199inter3, gate199inter4, gate199inter5, gate199inter6, gate199inter7, gate199inter8, gate199inter9, gate199inter10, gate199inter11, gate199inter12, gate32inter0, gate32inter1, gate32inter2, gate32inter3, gate32inter4, gate32inter5, gate32inter6, gate32inter7, gate32inter8, gate32inter9, gate32inter10, gate32inter11, gate32inter12, gate166inter0, gate166inter1, gate166inter2, gate166inter3, gate166inter4, gate166inter5, gate166inter6, gate166inter7, gate166inter8, gate166inter9, gate166inter10, gate166inter11, gate166inter12, gate209inter0, gate209inter1, gate209inter2, gate209inter3, gate209inter4, gate209inter5, gate209inter6, gate209inter7, gate209inter8, gate209inter9, gate209inter10, gate209inter11, gate209inter12, gate9inter0, gate9inter1, gate9inter2, gate9inter3, gate9inter4, gate9inter5, gate9inter6, gate9inter7, gate9inter8, gate9inter9, gate9inter10, gate9inter11, gate9inter12, gate486inter0, gate486inter1, gate486inter2, gate486inter3, gate486inter4, gate486inter5, gate486inter6, gate486inter7, gate486inter8, gate486inter9, gate486inter10, gate486inter11, gate486inter12, gate452inter0, gate452inter1, gate452inter2, gate452inter3, gate452inter4, gate452inter5, gate452inter6, gate452inter7, gate452inter8, gate452inter9, gate452inter10, gate452inter11, gate452inter12, gate495inter0, gate495inter1, gate495inter2, gate495inter3, gate495inter4, gate495inter5, gate495inter6, gate495inter7, gate495inter8, gate495inter9, gate495inter10, gate495inter11, gate495inter12, gate487inter0, gate487inter1, gate487inter2, gate487inter3, gate487inter4, gate487inter5, gate487inter6, gate487inter7, gate487inter8, gate487inter9, gate487inter10, gate487inter11, gate487inter12, gate449inter0, gate449inter1, gate449inter2, gate449inter3, gate449inter4, gate449inter5, gate449inter6, gate449inter7, gate449inter8, gate449inter9, gate449inter10, gate449inter11, gate449inter12, gate85inter0, gate85inter1, gate85inter2, gate85inter3, gate85inter4, gate85inter5, gate85inter6, gate85inter7, gate85inter8, gate85inter9, gate85inter10, gate85inter11, gate85inter12, gate236inter0, gate236inter1, gate236inter2, gate236inter3, gate236inter4, gate236inter5, gate236inter6, gate236inter7, gate236inter8, gate236inter9, gate236inter10, gate236inter11, gate236inter12, gate252inter0, gate252inter1, gate252inter2, gate252inter3, gate252inter4, gate252inter5, gate252inter6, gate252inter7, gate252inter8, gate252inter9, gate252inter10, gate252inter11, gate252inter12, gate135inter0, gate135inter1, gate135inter2, gate135inter3, gate135inter4, gate135inter5, gate135inter6, gate135inter7, gate135inter8, gate135inter9, gate135inter10, gate135inter11, gate135inter12, gate70inter0, gate70inter1, gate70inter2, gate70inter3, gate70inter4, gate70inter5, gate70inter6, gate70inter7, gate70inter8, gate70inter9, gate70inter10, gate70inter11, gate70inter12, gate512inter0, gate512inter1, gate512inter2, gate512inter3, gate512inter4, gate512inter5, gate512inter6, gate512inter7, gate512inter8, gate512inter9, gate512inter10, gate512inter11, gate512inter12, gate247inter0, gate247inter1, gate247inter2, gate247inter3, gate247inter4, gate247inter5, gate247inter6, gate247inter7, gate247inter8, gate247inter9, gate247inter10, gate247inter11, gate247inter12, gate141inter0, gate141inter1, gate141inter2, gate141inter3, gate141inter4, gate141inter5, gate141inter6, gate141inter7, gate141inter8, gate141inter9, gate141inter10, gate141inter11, gate141inter12, gate213inter0, gate213inter1, gate213inter2, gate213inter3, gate213inter4, gate213inter5, gate213inter6, gate213inter7, gate213inter8, gate213inter9, gate213inter10, gate213inter11, gate213inter12;



and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );

  xor2  gate2661(.a(G2), .b(G1), .O(gate9inter0));
  nand2 gate2662(.a(gate9inter0), .b(s_302), .O(gate9inter1));
  and2  gate2663(.a(G2), .b(G1), .O(gate9inter2));
  inv1  gate2664(.a(s_302), .O(gate9inter3));
  inv1  gate2665(.a(s_303), .O(gate9inter4));
  nand2 gate2666(.a(gate9inter4), .b(gate9inter3), .O(gate9inter5));
  nor2  gate2667(.a(gate9inter5), .b(gate9inter2), .O(gate9inter6));
  inv1  gate2668(.a(G1), .O(gate9inter7));
  inv1  gate2669(.a(G2), .O(gate9inter8));
  nand2 gate2670(.a(gate9inter8), .b(gate9inter7), .O(gate9inter9));
  nand2 gate2671(.a(s_303), .b(gate9inter3), .O(gate9inter10));
  nor2  gate2672(.a(gate9inter10), .b(gate9inter9), .O(gate9inter11));
  nor2  gate2673(.a(gate9inter11), .b(gate9inter6), .O(gate9inter12));
  nand2 gate2674(.a(gate9inter12), .b(gate9inter1), .O(G266));
nand2 gate10( .a(G3), .b(G4), .O(G269) );
nand2 gate11( .a(G5), .b(G6), .O(G272) );
nand2 gate12( .a(G7), .b(G8), .O(G275) );
nand2 gate13( .a(G9), .b(G10), .O(G278) );

  xor2  gate1555(.a(G12), .b(G11), .O(gate14inter0));
  nand2 gate1556(.a(gate14inter0), .b(s_144), .O(gate14inter1));
  and2  gate1557(.a(G12), .b(G11), .O(gate14inter2));
  inv1  gate1558(.a(s_144), .O(gate14inter3));
  inv1  gate1559(.a(s_145), .O(gate14inter4));
  nand2 gate1560(.a(gate14inter4), .b(gate14inter3), .O(gate14inter5));
  nor2  gate1561(.a(gate14inter5), .b(gate14inter2), .O(gate14inter6));
  inv1  gate1562(.a(G11), .O(gate14inter7));
  inv1  gate1563(.a(G12), .O(gate14inter8));
  nand2 gate1564(.a(gate14inter8), .b(gate14inter7), .O(gate14inter9));
  nand2 gate1565(.a(s_145), .b(gate14inter3), .O(gate14inter10));
  nor2  gate1566(.a(gate14inter10), .b(gate14inter9), .O(gate14inter11));
  nor2  gate1567(.a(gate14inter11), .b(gate14inter6), .O(gate14inter12));
  nand2 gate1568(.a(gate14inter12), .b(gate14inter1), .O(G281));

  xor2  gate855(.a(G14), .b(G13), .O(gate15inter0));
  nand2 gate856(.a(gate15inter0), .b(s_44), .O(gate15inter1));
  and2  gate857(.a(G14), .b(G13), .O(gate15inter2));
  inv1  gate858(.a(s_44), .O(gate15inter3));
  inv1  gate859(.a(s_45), .O(gate15inter4));
  nand2 gate860(.a(gate15inter4), .b(gate15inter3), .O(gate15inter5));
  nor2  gate861(.a(gate15inter5), .b(gate15inter2), .O(gate15inter6));
  inv1  gate862(.a(G13), .O(gate15inter7));
  inv1  gate863(.a(G14), .O(gate15inter8));
  nand2 gate864(.a(gate15inter8), .b(gate15inter7), .O(gate15inter9));
  nand2 gate865(.a(s_45), .b(gate15inter3), .O(gate15inter10));
  nor2  gate866(.a(gate15inter10), .b(gate15inter9), .O(gate15inter11));
  nor2  gate867(.a(gate15inter11), .b(gate15inter6), .O(gate15inter12));
  nand2 gate868(.a(gate15inter12), .b(gate15inter1), .O(G284));

  xor2  gate1275(.a(G16), .b(G15), .O(gate16inter0));
  nand2 gate1276(.a(gate16inter0), .b(s_104), .O(gate16inter1));
  and2  gate1277(.a(G16), .b(G15), .O(gate16inter2));
  inv1  gate1278(.a(s_104), .O(gate16inter3));
  inv1  gate1279(.a(s_105), .O(gate16inter4));
  nand2 gate1280(.a(gate16inter4), .b(gate16inter3), .O(gate16inter5));
  nor2  gate1281(.a(gate16inter5), .b(gate16inter2), .O(gate16inter6));
  inv1  gate1282(.a(G15), .O(gate16inter7));
  inv1  gate1283(.a(G16), .O(gate16inter8));
  nand2 gate1284(.a(gate16inter8), .b(gate16inter7), .O(gate16inter9));
  nand2 gate1285(.a(s_105), .b(gate16inter3), .O(gate16inter10));
  nor2  gate1286(.a(gate16inter10), .b(gate16inter9), .O(gate16inter11));
  nor2  gate1287(.a(gate16inter11), .b(gate16inter6), .O(gate16inter12));
  nand2 gate1288(.a(gate16inter12), .b(gate16inter1), .O(G287));
nand2 gate17( .a(G17), .b(G18), .O(G290) );
nand2 gate18( .a(G19), .b(G20), .O(G293) );

  xor2  gate1891(.a(G22), .b(G21), .O(gate19inter0));
  nand2 gate1892(.a(gate19inter0), .b(s_192), .O(gate19inter1));
  and2  gate1893(.a(G22), .b(G21), .O(gate19inter2));
  inv1  gate1894(.a(s_192), .O(gate19inter3));
  inv1  gate1895(.a(s_193), .O(gate19inter4));
  nand2 gate1896(.a(gate19inter4), .b(gate19inter3), .O(gate19inter5));
  nor2  gate1897(.a(gate19inter5), .b(gate19inter2), .O(gate19inter6));
  inv1  gate1898(.a(G21), .O(gate19inter7));
  inv1  gate1899(.a(G22), .O(gate19inter8));
  nand2 gate1900(.a(gate19inter8), .b(gate19inter7), .O(gate19inter9));
  nand2 gate1901(.a(s_193), .b(gate19inter3), .O(gate19inter10));
  nor2  gate1902(.a(gate19inter10), .b(gate19inter9), .O(gate19inter11));
  nor2  gate1903(.a(gate19inter11), .b(gate19inter6), .O(gate19inter12));
  nand2 gate1904(.a(gate19inter12), .b(gate19inter1), .O(G296));
nand2 gate20( .a(G23), .b(G24), .O(G299) );
nand2 gate21( .a(G25), .b(G26), .O(G302) );

  xor2  gate1975(.a(G28), .b(G27), .O(gate22inter0));
  nand2 gate1976(.a(gate22inter0), .b(s_204), .O(gate22inter1));
  and2  gate1977(.a(G28), .b(G27), .O(gate22inter2));
  inv1  gate1978(.a(s_204), .O(gate22inter3));
  inv1  gate1979(.a(s_205), .O(gate22inter4));
  nand2 gate1980(.a(gate22inter4), .b(gate22inter3), .O(gate22inter5));
  nor2  gate1981(.a(gate22inter5), .b(gate22inter2), .O(gate22inter6));
  inv1  gate1982(.a(G27), .O(gate22inter7));
  inv1  gate1983(.a(G28), .O(gate22inter8));
  nand2 gate1984(.a(gate22inter8), .b(gate22inter7), .O(gate22inter9));
  nand2 gate1985(.a(s_205), .b(gate22inter3), .O(gate22inter10));
  nor2  gate1986(.a(gate22inter10), .b(gate22inter9), .O(gate22inter11));
  nor2  gate1987(.a(gate22inter11), .b(gate22inter6), .O(gate22inter12));
  nand2 gate1988(.a(gate22inter12), .b(gate22inter1), .O(G305));
nand2 gate23( .a(G29), .b(G30), .O(G308) );
nand2 gate24( .a(G31), .b(G32), .O(G311) );
nand2 gate25( .a(G1), .b(G5), .O(G314) );
nand2 gate26( .a(G9), .b(G13), .O(G317) );

  xor2  gate1793(.a(G6), .b(G2), .O(gate27inter0));
  nand2 gate1794(.a(gate27inter0), .b(s_178), .O(gate27inter1));
  and2  gate1795(.a(G6), .b(G2), .O(gate27inter2));
  inv1  gate1796(.a(s_178), .O(gate27inter3));
  inv1  gate1797(.a(s_179), .O(gate27inter4));
  nand2 gate1798(.a(gate27inter4), .b(gate27inter3), .O(gate27inter5));
  nor2  gate1799(.a(gate27inter5), .b(gate27inter2), .O(gate27inter6));
  inv1  gate1800(.a(G2), .O(gate27inter7));
  inv1  gate1801(.a(G6), .O(gate27inter8));
  nand2 gate1802(.a(gate27inter8), .b(gate27inter7), .O(gate27inter9));
  nand2 gate1803(.a(s_179), .b(gate27inter3), .O(gate27inter10));
  nor2  gate1804(.a(gate27inter10), .b(gate27inter9), .O(gate27inter11));
  nor2  gate1805(.a(gate27inter11), .b(gate27inter6), .O(gate27inter12));
  nand2 gate1806(.a(gate27inter12), .b(gate27inter1), .O(G320));
nand2 gate28( .a(G10), .b(G14), .O(G323) );
nand2 gate29( .a(G3), .b(G7), .O(G326) );
nand2 gate30( .a(G11), .b(G15), .O(G329) );

  xor2  gate2003(.a(G8), .b(G4), .O(gate31inter0));
  nand2 gate2004(.a(gate31inter0), .b(s_208), .O(gate31inter1));
  and2  gate2005(.a(G8), .b(G4), .O(gate31inter2));
  inv1  gate2006(.a(s_208), .O(gate31inter3));
  inv1  gate2007(.a(s_209), .O(gate31inter4));
  nand2 gate2008(.a(gate31inter4), .b(gate31inter3), .O(gate31inter5));
  nor2  gate2009(.a(gate31inter5), .b(gate31inter2), .O(gate31inter6));
  inv1  gate2010(.a(G4), .O(gate31inter7));
  inv1  gate2011(.a(G8), .O(gate31inter8));
  nand2 gate2012(.a(gate31inter8), .b(gate31inter7), .O(gate31inter9));
  nand2 gate2013(.a(s_209), .b(gate31inter3), .O(gate31inter10));
  nor2  gate2014(.a(gate31inter10), .b(gate31inter9), .O(gate31inter11));
  nor2  gate2015(.a(gate31inter11), .b(gate31inter6), .O(gate31inter12));
  nand2 gate2016(.a(gate31inter12), .b(gate31inter1), .O(G332));

  xor2  gate2619(.a(G16), .b(G12), .O(gate32inter0));
  nand2 gate2620(.a(gate32inter0), .b(s_296), .O(gate32inter1));
  and2  gate2621(.a(G16), .b(G12), .O(gate32inter2));
  inv1  gate2622(.a(s_296), .O(gate32inter3));
  inv1  gate2623(.a(s_297), .O(gate32inter4));
  nand2 gate2624(.a(gate32inter4), .b(gate32inter3), .O(gate32inter5));
  nor2  gate2625(.a(gate32inter5), .b(gate32inter2), .O(gate32inter6));
  inv1  gate2626(.a(G12), .O(gate32inter7));
  inv1  gate2627(.a(G16), .O(gate32inter8));
  nand2 gate2628(.a(gate32inter8), .b(gate32inter7), .O(gate32inter9));
  nand2 gate2629(.a(s_297), .b(gate32inter3), .O(gate32inter10));
  nor2  gate2630(.a(gate32inter10), .b(gate32inter9), .O(gate32inter11));
  nor2  gate2631(.a(gate32inter11), .b(gate32inter6), .O(gate32inter12));
  nand2 gate2632(.a(gate32inter12), .b(gate32inter1), .O(G335));
nand2 gate33( .a(G17), .b(G21), .O(G338) );

  xor2  gate1919(.a(G29), .b(G25), .O(gate34inter0));
  nand2 gate1920(.a(gate34inter0), .b(s_196), .O(gate34inter1));
  and2  gate1921(.a(G29), .b(G25), .O(gate34inter2));
  inv1  gate1922(.a(s_196), .O(gate34inter3));
  inv1  gate1923(.a(s_197), .O(gate34inter4));
  nand2 gate1924(.a(gate34inter4), .b(gate34inter3), .O(gate34inter5));
  nor2  gate1925(.a(gate34inter5), .b(gate34inter2), .O(gate34inter6));
  inv1  gate1926(.a(G25), .O(gate34inter7));
  inv1  gate1927(.a(G29), .O(gate34inter8));
  nand2 gate1928(.a(gate34inter8), .b(gate34inter7), .O(gate34inter9));
  nand2 gate1929(.a(s_197), .b(gate34inter3), .O(gate34inter10));
  nor2  gate1930(.a(gate34inter10), .b(gate34inter9), .O(gate34inter11));
  nor2  gate1931(.a(gate34inter11), .b(gate34inter6), .O(gate34inter12));
  nand2 gate1932(.a(gate34inter12), .b(gate34inter1), .O(G341));
nand2 gate35( .a(G18), .b(G22), .O(G344) );

  xor2  gate967(.a(G30), .b(G26), .O(gate36inter0));
  nand2 gate968(.a(gate36inter0), .b(s_60), .O(gate36inter1));
  and2  gate969(.a(G30), .b(G26), .O(gate36inter2));
  inv1  gate970(.a(s_60), .O(gate36inter3));
  inv1  gate971(.a(s_61), .O(gate36inter4));
  nand2 gate972(.a(gate36inter4), .b(gate36inter3), .O(gate36inter5));
  nor2  gate973(.a(gate36inter5), .b(gate36inter2), .O(gate36inter6));
  inv1  gate974(.a(G26), .O(gate36inter7));
  inv1  gate975(.a(G30), .O(gate36inter8));
  nand2 gate976(.a(gate36inter8), .b(gate36inter7), .O(gate36inter9));
  nand2 gate977(.a(s_61), .b(gate36inter3), .O(gate36inter10));
  nor2  gate978(.a(gate36inter10), .b(gate36inter9), .O(gate36inter11));
  nor2  gate979(.a(gate36inter11), .b(gate36inter6), .O(gate36inter12));
  nand2 gate980(.a(gate36inter12), .b(gate36inter1), .O(G347));
nand2 gate37( .a(G19), .b(G23), .O(G350) );
nand2 gate38( .a(G27), .b(G31), .O(G353) );
nand2 gate39( .a(G20), .b(G24), .O(G356) );
nand2 gate40( .a(G28), .b(G32), .O(G359) );
nand2 gate41( .a(G1), .b(G266), .O(G362) );
nand2 gate42( .a(G2), .b(G266), .O(G363) );

  xor2  gate757(.a(G269), .b(G3), .O(gate43inter0));
  nand2 gate758(.a(gate43inter0), .b(s_30), .O(gate43inter1));
  and2  gate759(.a(G269), .b(G3), .O(gate43inter2));
  inv1  gate760(.a(s_30), .O(gate43inter3));
  inv1  gate761(.a(s_31), .O(gate43inter4));
  nand2 gate762(.a(gate43inter4), .b(gate43inter3), .O(gate43inter5));
  nor2  gate763(.a(gate43inter5), .b(gate43inter2), .O(gate43inter6));
  inv1  gate764(.a(G3), .O(gate43inter7));
  inv1  gate765(.a(G269), .O(gate43inter8));
  nand2 gate766(.a(gate43inter8), .b(gate43inter7), .O(gate43inter9));
  nand2 gate767(.a(s_31), .b(gate43inter3), .O(gate43inter10));
  nor2  gate768(.a(gate43inter10), .b(gate43inter9), .O(gate43inter11));
  nor2  gate769(.a(gate43inter11), .b(gate43inter6), .O(gate43inter12));
  nand2 gate770(.a(gate43inter12), .b(gate43inter1), .O(G364));

  xor2  gate2227(.a(G269), .b(G4), .O(gate44inter0));
  nand2 gate2228(.a(gate44inter0), .b(s_240), .O(gate44inter1));
  and2  gate2229(.a(G269), .b(G4), .O(gate44inter2));
  inv1  gate2230(.a(s_240), .O(gate44inter3));
  inv1  gate2231(.a(s_241), .O(gate44inter4));
  nand2 gate2232(.a(gate44inter4), .b(gate44inter3), .O(gate44inter5));
  nor2  gate2233(.a(gate44inter5), .b(gate44inter2), .O(gate44inter6));
  inv1  gate2234(.a(G4), .O(gate44inter7));
  inv1  gate2235(.a(G269), .O(gate44inter8));
  nand2 gate2236(.a(gate44inter8), .b(gate44inter7), .O(gate44inter9));
  nand2 gate2237(.a(s_241), .b(gate44inter3), .O(gate44inter10));
  nor2  gate2238(.a(gate44inter10), .b(gate44inter9), .O(gate44inter11));
  nor2  gate2239(.a(gate44inter11), .b(gate44inter6), .O(gate44inter12));
  nand2 gate2240(.a(gate44inter12), .b(gate44inter1), .O(G365));

  xor2  gate1961(.a(G272), .b(G5), .O(gate45inter0));
  nand2 gate1962(.a(gate45inter0), .b(s_202), .O(gate45inter1));
  and2  gate1963(.a(G272), .b(G5), .O(gate45inter2));
  inv1  gate1964(.a(s_202), .O(gate45inter3));
  inv1  gate1965(.a(s_203), .O(gate45inter4));
  nand2 gate1966(.a(gate45inter4), .b(gate45inter3), .O(gate45inter5));
  nor2  gate1967(.a(gate45inter5), .b(gate45inter2), .O(gate45inter6));
  inv1  gate1968(.a(G5), .O(gate45inter7));
  inv1  gate1969(.a(G272), .O(gate45inter8));
  nand2 gate1970(.a(gate45inter8), .b(gate45inter7), .O(gate45inter9));
  nand2 gate1971(.a(s_203), .b(gate45inter3), .O(gate45inter10));
  nor2  gate1972(.a(gate45inter10), .b(gate45inter9), .O(gate45inter11));
  nor2  gate1973(.a(gate45inter11), .b(gate45inter6), .O(gate45inter12));
  nand2 gate1974(.a(gate45inter12), .b(gate45inter1), .O(G366));
nand2 gate46( .a(G6), .b(G272), .O(G367) );
nand2 gate47( .a(G7), .b(G275), .O(G368) );

  xor2  gate1989(.a(G275), .b(G8), .O(gate48inter0));
  nand2 gate1990(.a(gate48inter0), .b(s_206), .O(gate48inter1));
  and2  gate1991(.a(G275), .b(G8), .O(gate48inter2));
  inv1  gate1992(.a(s_206), .O(gate48inter3));
  inv1  gate1993(.a(s_207), .O(gate48inter4));
  nand2 gate1994(.a(gate48inter4), .b(gate48inter3), .O(gate48inter5));
  nor2  gate1995(.a(gate48inter5), .b(gate48inter2), .O(gate48inter6));
  inv1  gate1996(.a(G8), .O(gate48inter7));
  inv1  gate1997(.a(G275), .O(gate48inter8));
  nand2 gate1998(.a(gate48inter8), .b(gate48inter7), .O(gate48inter9));
  nand2 gate1999(.a(s_207), .b(gate48inter3), .O(gate48inter10));
  nor2  gate2000(.a(gate48inter10), .b(gate48inter9), .O(gate48inter11));
  nor2  gate2001(.a(gate48inter11), .b(gate48inter6), .O(gate48inter12));
  nand2 gate2002(.a(gate48inter12), .b(gate48inter1), .O(G369));
nand2 gate49( .a(G9), .b(G278), .O(G370) );
nand2 gate50( .a(G10), .b(G278), .O(G371) );
nand2 gate51( .a(G11), .b(G281), .O(G372) );

  xor2  gate603(.a(G281), .b(G12), .O(gate52inter0));
  nand2 gate604(.a(gate52inter0), .b(s_8), .O(gate52inter1));
  and2  gate605(.a(G281), .b(G12), .O(gate52inter2));
  inv1  gate606(.a(s_8), .O(gate52inter3));
  inv1  gate607(.a(s_9), .O(gate52inter4));
  nand2 gate608(.a(gate52inter4), .b(gate52inter3), .O(gate52inter5));
  nor2  gate609(.a(gate52inter5), .b(gate52inter2), .O(gate52inter6));
  inv1  gate610(.a(G12), .O(gate52inter7));
  inv1  gate611(.a(G281), .O(gate52inter8));
  nand2 gate612(.a(gate52inter8), .b(gate52inter7), .O(gate52inter9));
  nand2 gate613(.a(s_9), .b(gate52inter3), .O(gate52inter10));
  nor2  gate614(.a(gate52inter10), .b(gate52inter9), .O(gate52inter11));
  nor2  gate615(.a(gate52inter11), .b(gate52inter6), .O(gate52inter12));
  nand2 gate616(.a(gate52inter12), .b(gate52inter1), .O(G373));
nand2 gate53( .a(G13), .b(G284), .O(G374) );

  xor2  gate813(.a(G284), .b(G14), .O(gate54inter0));
  nand2 gate814(.a(gate54inter0), .b(s_38), .O(gate54inter1));
  and2  gate815(.a(G284), .b(G14), .O(gate54inter2));
  inv1  gate816(.a(s_38), .O(gate54inter3));
  inv1  gate817(.a(s_39), .O(gate54inter4));
  nand2 gate818(.a(gate54inter4), .b(gate54inter3), .O(gate54inter5));
  nor2  gate819(.a(gate54inter5), .b(gate54inter2), .O(gate54inter6));
  inv1  gate820(.a(G14), .O(gate54inter7));
  inv1  gate821(.a(G284), .O(gate54inter8));
  nand2 gate822(.a(gate54inter8), .b(gate54inter7), .O(gate54inter9));
  nand2 gate823(.a(s_39), .b(gate54inter3), .O(gate54inter10));
  nor2  gate824(.a(gate54inter10), .b(gate54inter9), .O(gate54inter11));
  nor2  gate825(.a(gate54inter11), .b(gate54inter6), .O(gate54inter12));
  nand2 gate826(.a(gate54inter12), .b(gate54inter1), .O(G375));

  xor2  gate2451(.a(G287), .b(G15), .O(gate55inter0));
  nand2 gate2452(.a(gate55inter0), .b(s_272), .O(gate55inter1));
  and2  gate2453(.a(G287), .b(G15), .O(gate55inter2));
  inv1  gate2454(.a(s_272), .O(gate55inter3));
  inv1  gate2455(.a(s_273), .O(gate55inter4));
  nand2 gate2456(.a(gate55inter4), .b(gate55inter3), .O(gate55inter5));
  nor2  gate2457(.a(gate55inter5), .b(gate55inter2), .O(gate55inter6));
  inv1  gate2458(.a(G15), .O(gate55inter7));
  inv1  gate2459(.a(G287), .O(gate55inter8));
  nand2 gate2460(.a(gate55inter8), .b(gate55inter7), .O(gate55inter9));
  nand2 gate2461(.a(s_273), .b(gate55inter3), .O(gate55inter10));
  nor2  gate2462(.a(gate55inter10), .b(gate55inter9), .O(gate55inter11));
  nor2  gate2463(.a(gate55inter11), .b(gate55inter6), .O(gate55inter12));
  nand2 gate2464(.a(gate55inter12), .b(gate55inter1), .O(G376));

  xor2  gate645(.a(G287), .b(G16), .O(gate56inter0));
  nand2 gate646(.a(gate56inter0), .b(s_14), .O(gate56inter1));
  and2  gate647(.a(G287), .b(G16), .O(gate56inter2));
  inv1  gate648(.a(s_14), .O(gate56inter3));
  inv1  gate649(.a(s_15), .O(gate56inter4));
  nand2 gate650(.a(gate56inter4), .b(gate56inter3), .O(gate56inter5));
  nor2  gate651(.a(gate56inter5), .b(gate56inter2), .O(gate56inter6));
  inv1  gate652(.a(G16), .O(gate56inter7));
  inv1  gate653(.a(G287), .O(gate56inter8));
  nand2 gate654(.a(gate56inter8), .b(gate56inter7), .O(gate56inter9));
  nand2 gate655(.a(s_15), .b(gate56inter3), .O(gate56inter10));
  nor2  gate656(.a(gate56inter10), .b(gate56inter9), .O(gate56inter11));
  nor2  gate657(.a(gate56inter11), .b(gate56inter6), .O(gate56inter12));
  nand2 gate658(.a(gate56inter12), .b(gate56inter1), .O(G377));

  xor2  gate2157(.a(G290), .b(G17), .O(gate57inter0));
  nand2 gate2158(.a(gate57inter0), .b(s_230), .O(gate57inter1));
  and2  gate2159(.a(G290), .b(G17), .O(gate57inter2));
  inv1  gate2160(.a(s_230), .O(gate57inter3));
  inv1  gate2161(.a(s_231), .O(gate57inter4));
  nand2 gate2162(.a(gate57inter4), .b(gate57inter3), .O(gate57inter5));
  nor2  gate2163(.a(gate57inter5), .b(gate57inter2), .O(gate57inter6));
  inv1  gate2164(.a(G17), .O(gate57inter7));
  inv1  gate2165(.a(G290), .O(gate57inter8));
  nand2 gate2166(.a(gate57inter8), .b(gate57inter7), .O(gate57inter9));
  nand2 gate2167(.a(s_231), .b(gate57inter3), .O(gate57inter10));
  nor2  gate2168(.a(gate57inter10), .b(gate57inter9), .O(gate57inter11));
  nor2  gate2169(.a(gate57inter11), .b(gate57inter6), .O(gate57inter12));
  nand2 gate2170(.a(gate57inter12), .b(gate57inter1), .O(G378));

  xor2  gate1695(.a(G290), .b(G18), .O(gate58inter0));
  nand2 gate1696(.a(gate58inter0), .b(s_164), .O(gate58inter1));
  and2  gate1697(.a(G290), .b(G18), .O(gate58inter2));
  inv1  gate1698(.a(s_164), .O(gate58inter3));
  inv1  gate1699(.a(s_165), .O(gate58inter4));
  nand2 gate1700(.a(gate58inter4), .b(gate58inter3), .O(gate58inter5));
  nor2  gate1701(.a(gate58inter5), .b(gate58inter2), .O(gate58inter6));
  inv1  gate1702(.a(G18), .O(gate58inter7));
  inv1  gate1703(.a(G290), .O(gate58inter8));
  nand2 gate1704(.a(gate58inter8), .b(gate58inter7), .O(gate58inter9));
  nand2 gate1705(.a(s_165), .b(gate58inter3), .O(gate58inter10));
  nor2  gate1706(.a(gate58inter10), .b(gate58inter9), .O(gate58inter11));
  nor2  gate1707(.a(gate58inter11), .b(gate58inter6), .O(gate58inter12));
  nand2 gate1708(.a(gate58inter12), .b(gate58inter1), .O(G379));
nand2 gate59( .a(G19), .b(G293), .O(G380) );
nand2 gate60( .a(G20), .b(G293), .O(G381) );
nand2 gate61( .a(G21), .b(G296), .O(G382) );
nand2 gate62( .a(G22), .b(G296), .O(G383) );
nand2 gate63( .a(G23), .b(G299), .O(G384) );
nand2 gate64( .a(G24), .b(G299), .O(G385) );
nand2 gate65( .a(G25), .b(G302), .O(G386) );
nand2 gate66( .a(G26), .b(G302), .O(G387) );
nand2 gate67( .a(G27), .b(G305), .O(G388) );

  xor2  gate1149(.a(G305), .b(G28), .O(gate68inter0));
  nand2 gate1150(.a(gate68inter0), .b(s_86), .O(gate68inter1));
  and2  gate1151(.a(G305), .b(G28), .O(gate68inter2));
  inv1  gate1152(.a(s_86), .O(gate68inter3));
  inv1  gate1153(.a(s_87), .O(gate68inter4));
  nand2 gate1154(.a(gate68inter4), .b(gate68inter3), .O(gate68inter5));
  nor2  gate1155(.a(gate68inter5), .b(gate68inter2), .O(gate68inter6));
  inv1  gate1156(.a(G28), .O(gate68inter7));
  inv1  gate1157(.a(G305), .O(gate68inter8));
  nand2 gate1158(.a(gate68inter8), .b(gate68inter7), .O(gate68inter9));
  nand2 gate1159(.a(s_87), .b(gate68inter3), .O(gate68inter10));
  nor2  gate1160(.a(gate68inter10), .b(gate68inter9), .O(gate68inter11));
  nor2  gate1161(.a(gate68inter11), .b(gate68inter6), .O(gate68inter12));
  nand2 gate1162(.a(gate68inter12), .b(gate68inter1), .O(G389));
nand2 gate69( .a(G29), .b(G308), .O(G390) );

  xor2  gate2801(.a(G308), .b(G30), .O(gate70inter0));
  nand2 gate2802(.a(gate70inter0), .b(s_322), .O(gate70inter1));
  and2  gate2803(.a(G308), .b(G30), .O(gate70inter2));
  inv1  gate2804(.a(s_322), .O(gate70inter3));
  inv1  gate2805(.a(s_323), .O(gate70inter4));
  nand2 gate2806(.a(gate70inter4), .b(gate70inter3), .O(gate70inter5));
  nor2  gate2807(.a(gate70inter5), .b(gate70inter2), .O(gate70inter6));
  inv1  gate2808(.a(G30), .O(gate70inter7));
  inv1  gate2809(.a(G308), .O(gate70inter8));
  nand2 gate2810(.a(gate70inter8), .b(gate70inter7), .O(gate70inter9));
  nand2 gate2811(.a(s_323), .b(gate70inter3), .O(gate70inter10));
  nor2  gate2812(.a(gate70inter10), .b(gate70inter9), .O(gate70inter11));
  nor2  gate2813(.a(gate70inter11), .b(gate70inter6), .O(gate70inter12));
  nand2 gate2814(.a(gate70inter12), .b(gate70inter1), .O(G391));
nand2 gate71( .a(G31), .b(G311), .O(G392) );

  xor2  gate1219(.a(G311), .b(G32), .O(gate72inter0));
  nand2 gate1220(.a(gate72inter0), .b(s_96), .O(gate72inter1));
  and2  gate1221(.a(G311), .b(G32), .O(gate72inter2));
  inv1  gate1222(.a(s_96), .O(gate72inter3));
  inv1  gate1223(.a(s_97), .O(gate72inter4));
  nand2 gate1224(.a(gate72inter4), .b(gate72inter3), .O(gate72inter5));
  nor2  gate1225(.a(gate72inter5), .b(gate72inter2), .O(gate72inter6));
  inv1  gate1226(.a(G32), .O(gate72inter7));
  inv1  gate1227(.a(G311), .O(gate72inter8));
  nand2 gate1228(.a(gate72inter8), .b(gate72inter7), .O(gate72inter9));
  nand2 gate1229(.a(s_97), .b(gate72inter3), .O(gate72inter10));
  nor2  gate1230(.a(gate72inter10), .b(gate72inter9), .O(gate72inter11));
  nor2  gate1231(.a(gate72inter11), .b(gate72inter6), .O(gate72inter12));
  nand2 gate1232(.a(gate72inter12), .b(gate72inter1), .O(G393));
nand2 gate73( .a(G1), .b(G314), .O(G394) );

  xor2  gate729(.a(G314), .b(G5), .O(gate74inter0));
  nand2 gate730(.a(gate74inter0), .b(s_26), .O(gate74inter1));
  and2  gate731(.a(G314), .b(G5), .O(gate74inter2));
  inv1  gate732(.a(s_26), .O(gate74inter3));
  inv1  gate733(.a(s_27), .O(gate74inter4));
  nand2 gate734(.a(gate74inter4), .b(gate74inter3), .O(gate74inter5));
  nor2  gate735(.a(gate74inter5), .b(gate74inter2), .O(gate74inter6));
  inv1  gate736(.a(G5), .O(gate74inter7));
  inv1  gate737(.a(G314), .O(gate74inter8));
  nand2 gate738(.a(gate74inter8), .b(gate74inter7), .O(gate74inter9));
  nand2 gate739(.a(s_27), .b(gate74inter3), .O(gate74inter10));
  nor2  gate740(.a(gate74inter10), .b(gate74inter9), .O(gate74inter11));
  nor2  gate741(.a(gate74inter11), .b(gate74inter6), .O(gate74inter12));
  nand2 gate742(.a(gate74inter12), .b(gate74inter1), .O(G395));
nand2 gate75( .a(G9), .b(G317), .O(G396) );

  xor2  gate1415(.a(G317), .b(G13), .O(gate76inter0));
  nand2 gate1416(.a(gate76inter0), .b(s_124), .O(gate76inter1));
  and2  gate1417(.a(G317), .b(G13), .O(gate76inter2));
  inv1  gate1418(.a(s_124), .O(gate76inter3));
  inv1  gate1419(.a(s_125), .O(gate76inter4));
  nand2 gate1420(.a(gate76inter4), .b(gate76inter3), .O(gate76inter5));
  nor2  gate1421(.a(gate76inter5), .b(gate76inter2), .O(gate76inter6));
  inv1  gate1422(.a(G13), .O(gate76inter7));
  inv1  gate1423(.a(G317), .O(gate76inter8));
  nand2 gate1424(.a(gate76inter8), .b(gate76inter7), .O(gate76inter9));
  nand2 gate1425(.a(s_125), .b(gate76inter3), .O(gate76inter10));
  nor2  gate1426(.a(gate76inter10), .b(gate76inter9), .O(gate76inter11));
  nor2  gate1427(.a(gate76inter11), .b(gate76inter6), .O(gate76inter12));
  nand2 gate1428(.a(gate76inter12), .b(gate76inter1), .O(G397));
nand2 gate77( .a(G2), .b(G320), .O(G398) );
nand2 gate78( .a(G6), .b(G320), .O(G399) );

  xor2  gate2241(.a(G323), .b(G10), .O(gate79inter0));
  nand2 gate2242(.a(gate79inter0), .b(s_242), .O(gate79inter1));
  and2  gate2243(.a(G323), .b(G10), .O(gate79inter2));
  inv1  gate2244(.a(s_242), .O(gate79inter3));
  inv1  gate2245(.a(s_243), .O(gate79inter4));
  nand2 gate2246(.a(gate79inter4), .b(gate79inter3), .O(gate79inter5));
  nor2  gate2247(.a(gate79inter5), .b(gate79inter2), .O(gate79inter6));
  inv1  gate2248(.a(G10), .O(gate79inter7));
  inv1  gate2249(.a(G323), .O(gate79inter8));
  nand2 gate2250(.a(gate79inter8), .b(gate79inter7), .O(gate79inter9));
  nand2 gate2251(.a(s_243), .b(gate79inter3), .O(gate79inter10));
  nor2  gate2252(.a(gate79inter10), .b(gate79inter9), .O(gate79inter11));
  nor2  gate2253(.a(gate79inter11), .b(gate79inter6), .O(gate79inter12));
  nand2 gate2254(.a(gate79inter12), .b(gate79inter1), .O(G400));
nand2 gate80( .a(G14), .b(G323), .O(G401) );
nand2 gate81( .a(G3), .b(G326), .O(G402) );
nand2 gate82( .a(G7), .b(G326), .O(G403) );
nand2 gate83( .a(G11), .b(G329), .O(G404) );
nand2 gate84( .a(G15), .b(G329), .O(G405) );

  xor2  gate2745(.a(G332), .b(G4), .O(gate85inter0));
  nand2 gate2746(.a(gate85inter0), .b(s_314), .O(gate85inter1));
  and2  gate2747(.a(G332), .b(G4), .O(gate85inter2));
  inv1  gate2748(.a(s_314), .O(gate85inter3));
  inv1  gate2749(.a(s_315), .O(gate85inter4));
  nand2 gate2750(.a(gate85inter4), .b(gate85inter3), .O(gate85inter5));
  nor2  gate2751(.a(gate85inter5), .b(gate85inter2), .O(gate85inter6));
  inv1  gate2752(.a(G4), .O(gate85inter7));
  inv1  gate2753(.a(G332), .O(gate85inter8));
  nand2 gate2754(.a(gate85inter8), .b(gate85inter7), .O(gate85inter9));
  nand2 gate2755(.a(s_315), .b(gate85inter3), .O(gate85inter10));
  nor2  gate2756(.a(gate85inter10), .b(gate85inter9), .O(gate85inter11));
  nor2  gate2757(.a(gate85inter11), .b(gate85inter6), .O(gate85inter12));
  nand2 gate2758(.a(gate85inter12), .b(gate85inter1), .O(G406));

  xor2  gate1177(.a(G332), .b(G8), .O(gate86inter0));
  nand2 gate1178(.a(gate86inter0), .b(s_90), .O(gate86inter1));
  and2  gate1179(.a(G332), .b(G8), .O(gate86inter2));
  inv1  gate1180(.a(s_90), .O(gate86inter3));
  inv1  gate1181(.a(s_91), .O(gate86inter4));
  nand2 gate1182(.a(gate86inter4), .b(gate86inter3), .O(gate86inter5));
  nor2  gate1183(.a(gate86inter5), .b(gate86inter2), .O(gate86inter6));
  inv1  gate1184(.a(G8), .O(gate86inter7));
  inv1  gate1185(.a(G332), .O(gate86inter8));
  nand2 gate1186(.a(gate86inter8), .b(gate86inter7), .O(gate86inter9));
  nand2 gate1187(.a(s_91), .b(gate86inter3), .O(gate86inter10));
  nor2  gate1188(.a(gate86inter10), .b(gate86inter9), .O(gate86inter11));
  nor2  gate1189(.a(gate86inter11), .b(gate86inter6), .O(gate86inter12));
  nand2 gate1190(.a(gate86inter12), .b(gate86inter1), .O(G407));

  xor2  gate2101(.a(G335), .b(G12), .O(gate87inter0));
  nand2 gate2102(.a(gate87inter0), .b(s_222), .O(gate87inter1));
  and2  gate2103(.a(G335), .b(G12), .O(gate87inter2));
  inv1  gate2104(.a(s_222), .O(gate87inter3));
  inv1  gate2105(.a(s_223), .O(gate87inter4));
  nand2 gate2106(.a(gate87inter4), .b(gate87inter3), .O(gate87inter5));
  nor2  gate2107(.a(gate87inter5), .b(gate87inter2), .O(gate87inter6));
  inv1  gate2108(.a(G12), .O(gate87inter7));
  inv1  gate2109(.a(G335), .O(gate87inter8));
  nand2 gate2110(.a(gate87inter8), .b(gate87inter7), .O(gate87inter9));
  nand2 gate2111(.a(s_223), .b(gate87inter3), .O(gate87inter10));
  nor2  gate2112(.a(gate87inter10), .b(gate87inter9), .O(gate87inter11));
  nor2  gate2113(.a(gate87inter11), .b(gate87inter6), .O(gate87inter12));
  nand2 gate2114(.a(gate87inter12), .b(gate87inter1), .O(G408));
nand2 gate88( .a(G16), .b(G335), .O(G409) );
nand2 gate89( .a(G17), .b(G338), .O(G410) );
nand2 gate90( .a(G21), .b(G338), .O(G411) );

  xor2  gate2395(.a(G341), .b(G25), .O(gate91inter0));
  nand2 gate2396(.a(gate91inter0), .b(s_264), .O(gate91inter1));
  and2  gate2397(.a(G341), .b(G25), .O(gate91inter2));
  inv1  gate2398(.a(s_264), .O(gate91inter3));
  inv1  gate2399(.a(s_265), .O(gate91inter4));
  nand2 gate2400(.a(gate91inter4), .b(gate91inter3), .O(gate91inter5));
  nor2  gate2401(.a(gate91inter5), .b(gate91inter2), .O(gate91inter6));
  inv1  gate2402(.a(G25), .O(gate91inter7));
  inv1  gate2403(.a(G341), .O(gate91inter8));
  nand2 gate2404(.a(gate91inter8), .b(gate91inter7), .O(gate91inter9));
  nand2 gate2405(.a(s_265), .b(gate91inter3), .O(gate91inter10));
  nor2  gate2406(.a(gate91inter10), .b(gate91inter9), .O(gate91inter11));
  nor2  gate2407(.a(gate91inter11), .b(gate91inter6), .O(gate91inter12));
  nand2 gate2408(.a(gate91inter12), .b(gate91inter1), .O(G412));

  xor2  gate2129(.a(G341), .b(G29), .O(gate92inter0));
  nand2 gate2130(.a(gate92inter0), .b(s_226), .O(gate92inter1));
  and2  gate2131(.a(G341), .b(G29), .O(gate92inter2));
  inv1  gate2132(.a(s_226), .O(gate92inter3));
  inv1  gate2133(.a(s_227), .O(gate92inter4));
  nand2 gate2134(.a(gate92inter4), .b(gate92inter3), .O(gate92inter5));
  nor2  gate2135(.a(gate92inter5), .b(gate92inter2), .O(gate92inter6));
  inv1  gate2136(.a(G29), .O(gate92inter7));
  inv1  gate2137(.a(G341), .O(gate92inter8));
  nand2 gate2138(.a(gate92inter8), .b(gate92inter7), .O(gate92inter9));
  nand2 gate2139(.a(s_227), .b(gate92inter3), .O(gate92inter10));
  nor2  gate2140(.a(gate92inter10), .b(gate92inter9), .O(gate92inter11));
  nor2  gate2141(.a(gate92inter11), .b(gate92inter6), .O(gate92inter12));
  nand2 gate2142(.a(gate92inter12), .b(gate92inter1), .O(G413));

  xor2  gate1681(.a(G344), .b(G18), .O(gate93inter0));
  nand2 gate1682(.a(gate93inter0), .b(s_162), .O(gate93inter1));
  and2  gate1683(.a(G344), .b(G18), .O(gate93inter2));
  inv1  gate1684(.a(s_162), .O(gate93inter3));
  inv1  gate1685(.a(s_163), .O(gate93inter4));
  nand2 gate1686(.a(gate93inter4), .b(gate93inter3), .O(gate93inter5));
  nor2  gate1687(.a(gate93inter5), .b(gate93inter2), .O(gate93inter6));
  inv1  gate1688(.a(G18), .O(gate93inter7));
  inv1  gate1689(.a(G344), .O(gate93inter8));
  nand2 gate1690(.a(gate93inter8), .b(gate93inter7), .O(gate93inter9));
  nand2 gate1691(.a(s_163), .b(gate93inter3), .O(gate93inter10));
  nor2  gate1692(.a(gate93inter10), .b(gate93inter9), .O(gate93inter11));
  nor2  gate1693(.a(gate93inter11), .b(gate93inter6), .O(gate93inter12));
  nand2 gate1694(.a(gate93inter12), .b(gate93inter1), .O(G414));

  xor2  gate1401(.a(G344), .b(G22), .O(gate94inter0));
  nand2 gate1402(.a(gate94inter0), .b(s_122), .O(gate94inter1));
  and2  gate1403(.a(G344), .b(G22), .O(gate94inter2));
  inv1  gate1404(.a(s_122), .O(gate94inter3));
  inv1  gate1405(.a(s_123), .O(gate94inter4));
  nand2 gate1406(.a(gate94inter4), .b(gate94inter3), .O(gate94inter5));
  nor2  gate1407(.a(gate94inter5), .b(gate94inter2), .O(gate94inter6));
  inv1  gate1408(.a(G22), .O(gate94inter7));
  inv1  gate1409(.a(G344), .O(gate94inter8));
  nand2 gate1410(.a(gate94inter8), .b(gate94inter7), .O(gate94inter9));
  nand2 gate1411(.a(s_123), .b(gate94inter3), .O(gate94inter10));
  nor2  gate1412(.a(gate94inter10), .b(gate94inter9), .O(gate94inter11));
  nor2  gate1413(.a(gate94inter11), .b(gate94inter6), .O(gate94inter12));
  nand2 gate1414(.a(gate94inter12), .b(gate94inter1), .O(G415));
nand2 gate95( .a(G26), .b(G347), .O(G416) );
nand2 gate96( .a(G30), .b(G347), .O(G417) );

  xor2  gate2563(.a(G350), .b(G19), .O(gate97inter0));
  nand2 gate2564(.a(gate97inter0), .b(s_288), .O(gate97inter1));
  and2  gate2565(.a(G350), .b(G19), .O(gate97inter2));
  inv1  gate2566(.a(s_288), .O(gate97inter3));
  inv1  gate2567(.a(s_289), .O(gate97inter4));
  nand2 gate2568(.a(gate97inter4), .b(gate97inter3), .O(gate97inter5));
  nor2  gate2569(.a(gate97inter5), .b(gate97inter2), .O(gate97inter6));
  inv1  gate2570(.a(G19), .O(gate97inter7));
  inv1  gate2571(.a(G350), .O(gate97inter8));
  nand2 gate2572(.a(gate97inter8), .b(gate97inter7), .O(gate97inter9));
  nand2 gate2573(.a(s_289), .b(gate97inter3), .O(gate97inter10));
  nor2  gate2574(.a(gate97inter10), .b(gate97inter9), .O(gate97inter11));
  nor2  gate2575(.a(gate97inter11), .b(gate97inter6), .O(gate97inter12));
  nand2 gate2576(.a(gate97inter12), .b(gate97inter1), .O(G418));
nand2 gate98( .a(G23), .b(G350), .O(G419) );

  xor2  gate827(.a(G353), .b(G27), .O(gate99inter0));
  nand2 gate828(.a(gate99inter0), .b(s_40), .O(gate99inter1));
  and2  gate829(.a(G353), .b(G27), .O(gate99inter2));
  inv1  gate830(.a(s_40), .O(gate99inter3));
  inv1  gate831(.a(s_41), .O(gate99inter4));
  nand2 gate832(.a(gate99inter4), .b(gate99inter3), .O(gate99inter5));
  nor2  gate833(.a(gate99inter5), .b(gate99inter2), .O(gate99inter6));
  inv1  gate834(.a(G27), .O(gate99inter7));
  inv1  gate835(.a(G353), .O(gate99inter8));
  nand2 gate836(.a(gate99inter8), .b(gate99inter7), .O(gate99inter9));
  nand2 gate837(.a(s_41), .b(gate99inter3), .O(gate99inter10));
  nor2  gate838(.a(gate99inter10), .b(gate99inter9), .O(gate99inter11));
  nor2  gate839(.a(gate99inter11), .b(gate99inter6), .O(gate99inter12));
  nand2 gate840(.a(gate99inter12), .b(gate99inter1), .O(G420));
nand2 gate100( .a(G31), .b(G353), .O(G421) );
nand2 gate101( .a(G20), .b(G356), .O(G422) );
nand2 gate102( .a(G24), .b(G356), .O(G423) );
nand2 gate103( .a(G28), .b(G359), .O(G424) );

  xor2  gate2437(.a(G359), .b(G32), .O(gate104inter0));
  nand2 gate2438(.a(gate104inter0), .b(s_270), .O(gate104inter1));
  and2  gate2439(.a(G359), .b(G32), .O(gate104inter2));
  inv1  gate2440(.a(s_270), .O(gate104inter3));
  inv1  gate2441(.a(s_271), .O(gate104inter4));
  nand2 gate2442(.a(gate104inter4), .b(gate104inter3), .O(gate104inter5));
  nor2  gate2443(.a(gate104inter5), .b(gate104inter2), .O(gate104inter6));
  inv1  gate2444(.a(G32), .O(gate104inter7));
  inv1  gate2445(.a(G359), .O(gate104inter8));
  nand2 gate2446(.a(gate104inter8), .b(gate104inter7), .O(gate104inter9));
  nand2 gate2447(.a(s_271), .b(gate104inter3), .O(gate104inter10));
  nor2  gate2448(.a(gate104inter10), .b(gate104inter9), .O(gate104inter11));
  nor2  gate2449(.a(gate104inter11), .b(gate104inter6), .O(gate104inter12));
  nand2 gate2450(.a(gate104inter12), .b(gate104inter1), .O(G425));

  xor2  gate1751(.a(G363), .b(G362), .O(gate105inter0));
  nand2 gate1752(.a(gate105inter0), .b(s_172), .O(gate105inter1));
  and2  gate1753(.a(G363), .b(G362), .O(gate105inter2));
  inv1  gate1754(.a(s_172), .O(gate105inter3));
  inv1  gate1755(.a(s_173), .O(gate105inter4));
  nand2 gate1756(.a(gate105inter4), .b(gate105inter3), .O(gate105inter5));
  nor2  gate1757(.a(gate105inter5), .b(gate105inter2), .O(gate105inter6));
  inv1  gate1758(.a(G362), .O(gate105inter7));
  inv1  gate1759(.a(G363), .O(gate105inter8));
  nand2 gate1760(.a(gate105inter8), .b(gate105inter7), .O(gate105inter9));
  nand2 gate1761(.a(s_173), .b(gate105inter3), .O(gate105inter10));
  nor2  gate1762(.a(gate105inter10), .b(gate105inter9), .O(gate105inter11));
  nor2  gate1763(.a(gate105inter11), .b(gate105inter6), .O(gate105inter12));
  nand2 gate1764(.a(gate105inter12), .b(gate105inter1), .O(G426));

  xor2  gate2045(.a(G365), .b(G364), .O(gate106inter0));
  nand2 gate2046(.a(gate106inter0), .b(s_214), .O(gate106inter1));
  and2  gate2047(.a(G365), .b(G364), .O(gate106inter2));
  inv1  gate2048(.a(s_214), .O(gate106inter3));
  inv1  gate2049(.a(s_215), .O(gate106inter4));
  nand2 gate2050(.a(gate106inter4), .b(gate106inter3), .O(gate106inter5));
  nor2  gate2051(.a(gate106inter5), .b(gate106inter2), .O(gate106inter6));
  inv1  gate2052(.a(G364), .O(gate106inter7));
  inv1  gate2053(.a(G365), .O(gate106inter8));
  nand2 gate2054(.a(gate106inter8), .b(gate106inter7), .O(gate106inter9));
  nand2 gate2055(.a(s_215), .b(gate106inter3), .O(gate106inter10));
  nor2  gate2056(.a(gate106inter10), .b(gate106inter9), .O(gate106inter11));
  nor2  gate2057(.a(gate106inter11), .b(gate106inter6), .O(gate106inter12));
  nand2 gate2058(.a(gate106inter12), .b(gate106inter1), .O(G429));

  xor2  gate1947(.a(G367), .b(G366), .O(gate107inter0));
  nand2 gate1948(.a(gate107inter0), .b(s_200), .O(gate107inter1));
  and2  gate1949(.a(G367), .b(G366), .O(gate107inter2));
  inv1  gate1950(.a(s_200), .O(gate107inter3));
  inv1  gate1951(.a(s_201), .O(gate107inter4));
  nand2 gate1952(.a(gate107inter4), .b(gate107inter3), .O(gate107inter5));
  nor2  gate1953(.a(gate107inter5), .b(gate107inter2), .O(gate107inter6));
  inv1  gate1954(.a(G366), .O(gate107inter7));
  inv1  gate1955(.a(G367), .O(gate107inter8));
  nand2 gate1956(.a(gate107inter8), .b(gate107inter7), .O(gate107inter9));
  nand2 gate1957(.a(s_201), .b(gate107inter3), .O(gate107inter10));
  nor2  gate1958(.a(gate107inter10), .b(gate107inter9), .O(gate107inter11));
  nor2  gate1959(.a(gate107inter11), .b(gate107inter6), .O(gate107inter12));
  nand2 gate1960(.a(gate107inter12), .b(gate107inter1), .O(G432));
nand2 gate108( .a(G368), .b(G369), .O(G435) );

  xor2  gate1331(.a(G371), .b(G370), .O(gate109inter0));
  nand2 gate1332(.a(gate109inter0), .b(s_112), .O(gate109inter1));
  and2  gate1333(.a(G371), .b(G370), .O(gate109inter2));
  inv1  gate1334(.a(s_112), .O(gate109inter3));
  inv1  gate1335(.a(s_113), .O(gate109inter4));
  nand2 gate1336(.a(gate109inter4), .b(gate109inter3), .O(gate109inter5));
  nor2  gate1337(.a(gate109inter5), .b(gate109inter2), .O(gate109inter6));
  inv1  gate1338(.a(G370), .O(gate109inter7));
  inv1  gate1339(.a(G371), .O(gate109inter8));
  nand2 gate1340(.a(gate109inter8), .b(gate109inter7), .O(gate109inter9));
  nand2 gate1341(.a(s_113), .b(gate109inter3), .O(gate109inter10));
  nor2  gate1342(.a(gate109inter10), .b(gate109inter9), .O(gate109inter11));
  nor2  gate1343(.a(gate109inter11), .b(gate109inter6), .O(gate109inter12));
  nand2 gate1344(.a(gate109inter12), .b(gate109inter1), .O(G438));

  xor2  gate1583(.a(G373), .b(G372), .O(gate110inter0));
  nand2 gate1584(.a(gate110inter0), .b(s_148), .O(gate110inter1));
  and2  gate1585(.a(G373), .b(G372), .O(gate110inter2));
  inv1  gate1586(.a(s_148), .O(gate110inter3));
  inv1  gate1587(.a(s_149), .O(gate110inter4));
  nand2 gate1588(.a(gate110inter4), .b(gate110inter3), .O(gate110inter5));
  nor2  gate1589(.a(gate110inter5), .b(gate110inter2), .O(gate110inter6));
  inv1  gate1590(.a(G372), .O(gate110inter7));
  inv1  gate1591(.a(G373), .O(gate110inter8));
  nand2 gate1592(.a(gate110inter8), .b(gate110inter7), .O(gate110inter9));
  nand2 gate1593(.a(s_149), .b(gate110inter3), .O(gate110inter10));
  nor2  gate1594(.a(gate110inter10), .b(gate110inter9), .O(gate110inter11));
  nor2  gate1595(.a(gate110inter11), .b(gate110inter6), .O(gate110inter12));
  nand2 gate1596(.a(gate110inter12), .b(gate110inter1), .O(G441));
nand2 gate111( .a(G374), .b(G375), .O(G444) );
nand2 gate112( .a(G376), .b(G377), .O(G447) );
nand2 gate113( .a(G378), .b(G379), .O(G450) );
nand2 gate114( .a(G380), .b(G381), .O(G453) );

  xor2  gate841(.a(G383), .b(G382), .O(gate115inter0));
  nand2 gate842(.a(gate115inter0), .b(s_42), .O(gate115inter1));
  and2  gate843(.a(G383), .b(G382), .O(gate115inter2));
  inv1  gate844(.a(s_42), .O(gate115inter3));
  inv1  gate845(.a(s_43), .O(gate115inter4));
  nand2 gate846(.a(gate115inter4), .b(gate115inter3), .O(gate115inter5));
  nor2  gate847(.a(gate115inter5), .b(gate115inter2), .O(gate115inter6));
  inv1  gate848(.a(G382), .O(gate115inter7));
  inv1  gate849(.a(G383), .O(gate115inter8));
  nand2 gate850(.a(gate115inter8), .b(gate115inter7), .O(gate115inter9));
  nand2 gate851(.a(s_43), .b(gate115inter3), .O(gate115inter10));
  nor2  gate852(.a(gate115inter10), .b(gate115inter9), .O(gate115inter11));
  nor2  gate853(.a(gate115inter11), .b(gate115inter6), .O(gate115inter12));
  nand2 gate854(.a(gate115inter12), .b(gate115inter1), .O(G456));
nand2 gate116( .a(G384), .b(G385), .O(G459) );
nand2 gate117( .a(G386), .b(G387), .O(G462) );

  xor2  gate1373(.a(G389), .b(G388), .O(gate118inter0));
  nand2 gate1374(.a(gate118inter0), .b(s_118), .O(gate118inter1));
  and2  gate1375(.a(G389), .b(G388), .O(gate118inter2));
  inv1  gate1376(.a(s_118), .O(gate118inter3));
  inv1  gate1377(.a(s_119), .O(gate118inter4));
  nand2 gate1378(.a(gate118inter4), .b(gate118inter3), .O(gate118inter5));
  nor2  gate1379(.a(gate118inter5), .b(gate118inter2), .O(gate118inter6));
  inv1  gate1380(.a(G388), .O(gate118inter7));
  inv1  gate1381(.a(G389), .O(gate118inter8));
  nand2 gate1382(.a(gate118inter8), .b(gate118inter7), .O(gate118inter9));
  nand2 gate1383(.a(s_119), .b(gate118inter3), .O(gate118inter10));
  nor2  gate1384(.a(gate118inter10), .b(gate118inter9), .O(gate118inter11));
  nor2  gate1385(.a(gate118inter11), .b(gate118inter6), .O(gate118inter12));
  nand2 gate1386(.a(gate118inter12), .b(gate118inter1), .O(G465));

  xor2  gate925(.a(G391), .b(G390), .O(gate119inter0));
  nand2 gate926(.a(gate119inter0), .b(s_54), .O(gate119inter1));
  and2  gate927(.a(G391), .b(G390), .O(gate119inter2));
  inv1  gate928(.a(s_54), .O(gate119inter3));
  inv1  gate929(.a(s_55), .O(gate119inter4));
  nand2 gate930(.a(gate119inter4), .b(gate119inter3), .O(gate119inter5));
  nor2  gate931(.a(gate119inter5), .b(gate119inter2), .O(gate119inter6));
  inv1  gate932(.a(G390), .O(gate119inter7));
  inv1  gate933(.a(G391), .O(gate119inter8));
  nand2 gate934(.a(gate119inter8), .b(gate119inter7), .O(gate119inter9));
  nand2 gate935(.a(s_55), .b(gate119inter3), .O(gate119inter10));
  nor2  gate936(.a(gate119inter10), .b(gate119inter9), .O(gate119inter11));
  nor2  gate937(.a(gate119inter11), .b(gate119inter6), .O(gate119inter12));
  nand2 gate938(.a(gate119inter12), .b(gate119inter1), .O(G468));
nand2 gate120( .a(G392), .b(G393), .O(G471) );
nand2 gate121( .a(G394), .b(G395), .O(G474) );
nand2 gate122( .a(G396), .b(G397), .O(G477) );
nand2 gate123( .a(G398), .b(G399), .O(G480) );
nand2 gate124( .a(G400), .b(G401), .O(G483) );
nand2 gate125( .a(G402), .b(G403), .O(G486) );
nand2 gate126( .a(G404), .b(G405), .O(G489) );
nand2 gate127( .a(G406), .b(G407), .O(G492) );
nand2 gate128( .a(G408), .b(G409), .O(G495) );
nand2 gate129( .a(G410), .b(G411), .O(G498) );
nand2 gate130( .a(G412), .b(G413), .O(G501) );
nand2 gate131( .a(G414), .b(G415), .O(G504) );

  xor2  gate1877(.a(G417), .b(G416), .O(gate132inter0));
  nand2 gate1878(.a(gate132inter0), .b(s_190), .O(gate132inter1));
  and2  gate1879(.a(G417), .b(G416), .O(gate132inter2));
  inv1  gate1880(.a(s_190), .O(gate132inter3));
  inv1  gate1881(.a(s_191), .O(gate132inter4));
  nand2 gate1882(.a(gate132inter4), .b(gate132inter3), .O(gate132inter5));
  nor2  gate1883(.a(gate132inter5), .b(gate132inter2), .O(gate132inter6));
  inv1  gate1884(.a(G416), .O(gate132inter7));
  inv1  gate1885(.a(G417), .O(gate132inter8));
  nand2 gate1886(.a(gate132inter8), .b(gate132inter7), .O(gate132inter9));
  nand2 gate1887(.a(s_191), .b(gate132inter3), .O(gate132inter10));
  nor2  gate1888(.a(gate132inter10), .b(gate132inter9), .O(gate132inter11));
  nor2  gate1889(.a(gate132inter11), .b(gate132inter6), .O(gate132inter12));
  nand2 gate1890(.a(gate132inter12), .b(gate132inter1), .O(G507));

  xor2  gate2213(.a(G419), .b(G418), .O(gate133inter0));
  nand2 gate2214(.a(gate133inter0), .b(s_238), .O(gate133inter1));
  and2  gate2215(.a(G419), .b(G418), .O(gate133inter2));
  inv1  gate2216(.a(s_238), .O(gate133inter3));
  inv1  gate2217(.a(s_239), .O(gate133inter4));
  nand2 gate2218(.a(gate133inter4), .b(gate133inter3), .O(gate133inter5));
  nor2  gate2219(.a(gate133inter5), .b(gate133inter2), .O(gate133inter6));
  inv1  gate2220(.a(G418), .O(gate133inter7));
  inv1  gate2221(.a(G419), .O(gate133inter8));
  nand2 gate2222(.a(gate133inter8), .b(gate133inter7), .O(gate133inter9));
  nand2 gate2223(.a(s_239), .b(gate133inter3), .O(gate133inter10));
  nor2  gate2224(.a(gate133inter10), .b(gate133inter9), .O(gate133inter11));
  nor2  gate2225(.a(gate133inter11), .b(gate133inter6), .O(gate133inter12));
  nand2 gate2226(.a(gate133inter12), .b(gate133inter1), .O(G510));

  xor2  gate1443(.a(G421), .b(G420), .O(gate134inter0));
  nand2 gate1444(.a(gate134inter0), .b(s_128), .O(gate134inter1));
  and2  gate1445(.a(G421), .b(G420), .O(gate134inter2));
  inv1  gate1446(.a(s_128), .O(gate134inter3));
  inv1  gate1447(.a(s_129), .O(gate134inter4));
  nand2 gate1448(.a(gate134inter4), .b(gate134inter3), .O(gate134inter5));
  nor2  gate1449(.a(gate134inter5), .b(gate134inter2), .O(gate134inter6));
  inv1  gate1450(.a(G420), .O(gate134inter7));
  inv1  gate1451(.a(G421), .O(gate134inter8));
  nand2 gate1452(.a(gate134inter8), .b(gate134inter7), .O(gate134inter9));
  nand2 gate1453(.a(s_129), .b(gate134inter3), .O(gate134inter10));
  nor2  gate1454(.a(gate134inter10), .b(gate134inter9), .O(gate134inter11));
  nor2  gate1455(.a(gate134inter11), .b(gate134inter6), .O(gate134inter12));
  nand2 gate1456(.a(gate134inter12), .b(gate134inter1), .O(G513));

  xor2  gate2787(.a(G423), .b(G422), .O(gate135inter0));
  nand2 gate2788(.a(gate135inter0), .b(s_320), .O(gate135inter1));
  and2  gate2789(.a(G423), .b(G422), .O(gate135inter2));
  inv1  gate2790(.a(s_320), .O(gate135inter3));
  inv1  gate2791(.a(s_321), .O(gate135inter4));
  nand2 gate2792(.a(gate135inter4), .b(gate135inter3), .O(gate135inter5));
  nor2  gate2793(.a(gate135inter5), .b(gate135inter2), .O(gate135inter6));
  inv1  gate2794(.a(G422), .O(gate135inter7));
  inv1  gate2795(.a(G423), .O(gate135inter8));
  nand2 gate2796(.a(gate135inter8), .b(gate135inter7), .O(gate135inter9));
  nand2 gate2797(.a(s_321), .b(gate135inter3), .O(gate135inter10));
  nor2  gate2798(.a(gate135inter10), .b(gate135inter9), .O(gate135inter11));
  nor2  gate2799(.a(gate135inter11), .b(gate135inter6), .O(gate135inter12));
  nand2 gate2800(.a(gate135inter12), .b(gate135inter1), .O(G516));
nand2 gate136( .a(G424), .b(G425), .O(G519) );

  xor2  gate2255(.a(G429), .b(G426), .O(gate137inter0));
  nand2 gate2256(.a(gate137inter0), .b(s_244), .O(gate137inter1));
  and2  gate2257(.a(G429), .b(G426), .O(gate137inter2));
  inv1  gate2258(.a(s_244), .O(gate137inter3));
  inv1  gate2259(.a(s_245), .O(gate137inter4));
  nand2 gate2260(.a(gate137inter4), .b(gate137inter3), .O(gate137inter5));
  nor2  gate2261(.a(gate137inter5), .b(gate137inter2), .O(gate137inter6));
  inv1  gate2262(.a(G426), .O(gate137inter7));
  inv1  gate2263(.a(G429), .O(gate137inter8));
  nand2 gate2264(.a(gate137inter8), .b(gate137inter7), .O(gate137inter9));
  nand2 gate2265(.a(s_245), .b(gate137inter3), .O(gate137inter10));
  nor2  gate2266(.a(gate137inter10), .b(gate137inter9), .O(gate137inter11));
  nor2  gate2267(.a(gate137inter11), .b(gate137inter6), .O(gate137inter12));
  nand2 gate2268(.a(gate137inter12), .b(gate137inter1), .O(G522));

  xor2  gate2199(.a(G435), .b(G432), .O(gate138inter0));
  nand2 gate2200(.a(gate138inter0), .b(s_236), .O(gate138inter1));
  and2  gate2201(.a(G435), .b(G432), .O(gate138inter2));
  inv1  gate2202(.a(s_236), .O(gate138inter3));
  inv1  gate2203(.a(s_237), .O(gate138inter4));
  nand2 gate2204(.a(gate138inter4), .b(gate138inter3), .O(gate138inter5));
  nor2  gate2205(.a(gate138inter5), .b(gate138inter2), .O(gate138inter6));
  inv1  gate2206(.a(G432), .O(gate138inter7));
  inv1  gate2207(.a(G435), .O(gate138inter8));
  nand2 gate2208(.a(gate138inter8), .b(gate138inter7), .O(gate138inter9));
  nand2 gate2209(.a(s_237), .b(gate138inter3), .O(gate138inter10));
  nor2  gate2210(.a(gate138inter10), .b(gate138inter9), .O(gate138inter11));
  nor2  gate2211(.a(gate138inter11), .b(gate138inter6), .O(gate138inter12));
  nand2 gate2212(.a(gate138inter12), .b(gate138inter1), .O(G525));

  xor2  gate659(.a(G441), .b(G438), .O(gate139inter0));
  nand2 gate660(.a(gate139inter0), .b(s_16), .O(gate139inter1));
  and2  gate661(.a(G441), .b(G438), .O(gate139inter2));
  inv1  gate662(.a(s_16), .O(gate139inter3));
  inv1  gate663(.a(s_17), .O(gate139inter4));
  nand2 gate664(.a(gate139inter4), .b(gate139inter3), .O(gate139inter5));
  nor2  gate665(.a(gate139inter5), .b(gate139inter2), .O(gate139inter6));
  inv1  gate666(.a(G438), .O(gate139inter7));
  inv1  gate667(.a(G441), .O(gate139inter8));
  nand2 gate668(.a(gate139inter8), .b(gate139inter7), .O(gate139inter9));
  nand2 gate669(.a(s_17), .b(gate139inter3), .O(gate139inter10));
  nor2  gate670(.a(gate139inter10), .b(gate139inter9), .O(gate139inter11));
  nor2  gate671(.a(gate139inter11), .b(gate139inter6), .O(gate139inter12));
  nand2 gate672(.a(gate139inter12), .b(gate139inter1), .O(G528));
nand2 gate140( .a(G444), .b(G447), .O(G531) );

  xor2  gate2843(.a(G453), .b(G450), .O(gate141inter0));
  nand2 gate2844(.a(gate141inter0), .b(s_328), .O(gate141inter1));
  and2  gate2845(.a(G453), .b(G450), .O(gate141inter2));
  inv1  gate2846(.a(s_328), .O(gate141inter3));
  inv1  gate2847(.a(s_329), .O(gate141inter4));
  nand2 gate2848(.a(gate141inter4), .b(gate141inter3), .O(gate141inter5));
  nor2  gate2849(.a(gate141inter5), .b(gate141inter2), .O(gate141inter6));
  inv1  gate2850(.a(G450), .O(gate141inter7));
  inv1  gate2851(.a(G453), .O(gate141inter8));
  nand2 gate2852(.a(gate141inter8), .b(gate141inter7), .O(gate141inter9));
  nand2 gate2853(.a(s_329), .b(gate141inter3), .O(gate141inter10));
  nor2  gate2854(.a(gate141inter10), .b(gate141inter9), .O(gate141inter11));
  nor2  gate2855(.a(gate141inter11), .b(gate141inter6), .O(gate141inter12));
  nand2 gate2856(.a(gate141inter12), .b(gate141inter1), .O(G534));
nand2 gate142( .a(G456), .b(G459), .O(G537) );
nand2 gate143( .a(G462), .b(G465), .O(G540) );

  xor2  gate2591(.a(G471), .b(G468), .O(gate144inter0));
  nand2 gate2592(.a(gate144inter0), .b(s_292), .O(gate144inter1));
  and2  gate2593(.a(G471), .b(G468), .O(gate144inter2));
  inv1  gate2594(.a(s_292), .O(gate144inter3));
  inv1  gate2595(.a(s_293), .O(gate144inter4));
  nand2 gate2596(.a(gate144inter4), .b(gate144inter3), .O(gate144inter5));
  nor2  gate2597(.a(gate144inter5), .b(gate144inter2), .O(gate144inter6));
  inv1  gate2598(.a(G468), .O(gate144inter7));
  inv1  gate2599(.a(G471), .O(gate144inter8));
  nand2 gate2600(.a(gate144inter8), .b(gate144inter7), .O(gate144inter9));
  nand2 gate2601(.a(s_293), .b(gate144inter3), .O(gate144inter10));
  nor2  gate2602(.a(gate144inter10), .b(gate144inter9), .O(gate144inter11));
  nor2  gate2603(.a(gate144inter11), .b(gate144inter6), .O(gate144inter12));
  nand2 gate2604(.a(gate144inter12), .b(gate144inter1), .O(G543));
nand2 gate145( .a(G474), .b(G477), .O(G546) );
nand2 gate146( .a(G480), .b(G483), .O(G549) );

  xor2  gate1163(.a(G489), .b(G486), .O(gate147inter0));
  nand2 gate1164(.a(gate147inter0), .b(s_88), .O(gate147inter1));
  and2  gate1165(.a(G489), .b(G486), .O(gate147inter2));
  inv1  gate1166(.a(s_88), .O(gate147inter3));
  inv1  gate1167(.a(s_89), .O(gate147inter4));
  nand2 gate1168(.a(gate147inter4), .b(gate147inter3), .O(gate147inter5));
  nor2  gate1169(.a(gate147inter5), .b(gate147inter2), .O(gate147inter6));
  inv1  gate1170(.a(G486), .O(gate147inter7));
  inv1  gate1171(.a(G489), .O(gate147inter8));
  nand2 gate1172(.a(gate147inter8), .b(gate147inter7), .O(gate147inter9));
  nand2 gate1173(.a(s_89), .b(gate147inter3), .O(gate147inter10));
  nor2  gate1174(.a(gate147inter10), .b(gate147inter9), .O(gate147inter11));
  nor2  gate1175(.a(gate147inter11), .b(gate147inter6), .O(gate147inter12));
  nand2 gate1176(.a(gate147inter12), .b(gate147inter1), .O(G552));
nand2 gate148( .a(G492), .b(G495), .O(G555) );
nand2 gate149( .a(G498), .b(G501), .O(G558) );

  xor2  gate1135(.a(G507), .b(G504), .O(gate150inter0));
  nand2 gate1136(.a(gate150inter0), .b(s_84), .O(gate150inter1));
  and2  gate1137(.a(G507), .b(G504), .O(gate150inter2));
  inv1  gate1138(.a(s_84), .O(gate150inter3));
  inv1  gate1139(.a(s_85), .O(gate150inter4));
  nand2 gate1140(.a(gate150inter4), .b(gate150inter3), .O(gate150inter5));
  nor2  gate1141(.a(gate150inter5), .b(gate150inter2), .O(gate150inter6));
  inv1  gate1142(.a(G504), .O(gate150inter7));
  inv1  gate1143(.a(G507), .O(gate150inter8));
  nand2 gate1144(.a(gate150inter8), .b(gate150inter7), .O(gate150inter9));
  nand2 gate1145(.a(s_85), .b(gate150inter3), .O(gate150inter10));
  nor2  gate1146(.a(gate150inter10), .b(gate150inter9), .O(gate150inter11));
  nor2  gate1147(.a(gate150inter11), .b(gate150inter6), .O(gate150inter12));
  nand2 gate1148(.a(gate150inter12), .b(gate150inter1), .O(G561));

  xor2  gate1205(.a(G513), .b(G510), .O(gate151inter0));
  nand2 gate1206(.a(gate151inter0), .b(s_94), .O(gate151inter1));
  and2  gate1207(.a(G513), .b(G510), .O(gate151inter2));
  inv1  gate1208(.a(s_94), .O(gate151inter3));
  inv1  gate1209(.a(s_95), .O(gate151inter4));
  nand2 gate1210(.a(gate151inter4), .b(gate151inter3), .O(gate151inter5));
  nor2  gate1211(.a(gate151inter5), .b(gate151inter2), .O(gate151inter6));
  inv1  gate1212(.a(G510), .O(gate151inter7));
  inv1  gate1213(.a(G513), .O(gate151inter8));
  nand2 gate1214(.a(gate151inter8), .b(gate151inter7), .O(gate151inter9));
  nand2 gate1215(.a(s_95), .b(gate151inter3), .O(gate151inter10));
  nor2  gate1216(.a(gate151inter10), .b(gate151inter9), .O(gate151inter11));
  nor2  gate1217(.a(gate151inter11), .b(gate151inter6), .O(gate151inter12));
  nand2 gate1218(.a(gate151inter12), .b(gate151inter1), .O(G564));
nand2 gate152( .a(G516), .b(G519), .O(G567) );
nand2 gate153( .a(G426), .b(G522), .O(G570) );
nand2 gate154( .a(G429), .b(G522), .O(G571) );

  xor2  gate1513(.a(G525), .b(G432), .O(gate155inter0));
  nand2 gate1514(.a(gate155inter0), .b(s_138), .O(gate155inter1));
  and2  gate1515(.a(G525), .b(G432), .O(gate155inter2));
  inv1  gate1516(.a(s_138), .O(gate155inter3));
  inv1  gate1517(.a(s_139), .O(gate155inter4));
  nand2 gate1518(.a(gate155inter4), .b(gate155inter3), .O(gate155inter5));
  nor2  gate1519(.a(gate155inter5), .b(gate155inter2), .O(gate155inter6));
  inv1  gate1520(.a(G432), .O(gate155inter7));
  inv1  gate1521(.a(G525), .O(gate155inter8));
  nand2 gate1522(.a(gate155inter8), .b(gate155inter7), .O(gate155inter9));
  nand2 gate1523(.a(s_139), .b(gate155inter3), .O(gate155inter10));
  nor2  gate1524(.a(gate155inter10), .b(gate155inter9), .O(gate155inter11));
  nor2  gate1525(.a(gate155inter11), .b(gate155inter6), .O(gate155inter12));
  nand2 gate1526(.a(gate155inter12), .b(gate155inter1), .O(G572));

  xor2  gate995(.a(G525), .b(G435), .O(gate156inter0));
  nand2 gate996(.a(gate156inter0), .b(s_64), .O(gate156inter1));
  and2  gate997(.a(G525), .b(G435), .O(gate156inter2));
  inv1  gate998(.a(s_64), .O(gate156inter3));
  inv1  gate999(.a(s_65), .O(gate156inter4));
  nand2 gate1000(.a(gate156inter4), .b(gate156inter3), .O(gate156inter5));
  nor2  gate1001(.a(gate156inter5), .b(gate156inter2), .O(gate156inter6));
  inv1  gate1002(.a(G435), .O(gate156inter7));
  inv1  gate1003(.a(G525), .O(gate156inter8));
  nand2 gate1004(.a(gate156inter8), .b(gate156inter7), .O(gate156inter9));
  nand2 gate1005(.a(s_65), .b(gate156inter3), .O(gate156inter10));
  nor2  gate1006(.a(gate156inter10), .b(gate156inter9), .O(gate156inter11));
  nor2  gate1007(.a(gate156inter11), .b(gate156inter6), .O(gate156inter12));
  nand2 gate1008(.a(gate156inter12), .b(gate156inter1), .O(G573));

  xor2  gate547(.a(G528), .b(G438), .O(gate157inter0));
  nand2 gate548(.a(gate157inter0), .b(s_0), .O(gate157inter1));
  and2  gate549(.a(G528), .b(G438), .O(gate157inter2));
  inv1  gate550(.a(s_0), .O(gate157inter3));
  inv1  gate551(.a(s_1), .O(gate157inter4));
  nand2 gate552(.a(gate157inter4), .b(gate157inter3), .O(gate157inter5));
  nor2  gate553(.a(gate157inter5), .b(gate157inter2), .O(gate157inter6));
  inv1  gate554(.a(G438), .O(gate157inter7));
  inv1  gate555(.a(G528), .O(gate157inter8));
  nand2 gate556(.a(gate157inter8), .b(gate157inter7), .O(gate157inter9));
  nand2 gate557(.a(s_1), .b(gate157inter3), .O(gate157inter10));
  nor2  gate558(.a(gate157inter10), .b(gate157inter9), .O(gate157inter11));
  nor2  gate559(.a(gate157inter11), .b(gate157inter6), .O(gate157inter12));
  nand2 gate560(.a(gate157inter12), .b(gate157inter1), .O(G574));

  xor2  gate687(.a(G528), .b(G441), .O(gate158inter0));
  nand2 gate688(.a(gate158inter0), .b(s_20), .O(gate158inter1));
  and2  gate689(.a(G528), .b(G441), .O(gate158inter2));
  inv1  gate690(.a(s_20), .O(gate158inter3));
  inv1  gate691(.a(s_21), .O(gate158inter4));
  nand2 gate692(.a(gate158inter4), .b(gate158inter3), .O(gate158inter5));
  nor2  gate693(.a(gate158inter5), .b(gate158inter2), .O(gate158inter6));
  inv1  gate694(.a(G441), .O(gate158inter7));
  inv1  gate695(.a(G528), .O(gate158inter8));
  nand2 gate696(.a(gate158inter8), .b(gate158inter7), .O(gate158inter9));
  nand2 gate697(.a(s_21), .b(gate158inter3), .O(gate158inter10));
  nor2  gate698(.a(gate158inter10), .b(gate158inter9), .O(gate158inter11));
  nor2  gate699(.a(gate158inter11), .b(gate158inter6), .O(gate158inter12));
  nand2 gate700(.a(gate158inter12), .b(gate158inter1), .O(G575));

  xor2  gate1723(.a(G531), .b(G444), .O(gate159inter0));
  nand2 gate1724(.a(gate159inter0), .b(s_168), .O(gate159inter1));
  and2  gate1725(.a(G531), .b(G444), .O(gate159inter2));
  inv1  gate1726(.a(s_168), .O(gate159inter3));
  inv1  gate1727(.a(s_169), .O(gate159inter4));
  nand2 gate1728(.a(gate159inter4), .b(gate159inter3), .O(gate159inter5));
  nor2  gate1729(.a(gate159inter5), .b(gate159inter2), .O(gate159inter6));
  inv1  gate1730(.a(G444), .O(gate159inter7));
  inv1  gate1731(.a(G531), .O(gate159inter8));
  nand2 gate1732(.a(gate159inter8), .b(gate159inter7), .O(gate159inter9));
  nand2 gate1733(.a(s_169), .b(gate159inter3), .O(gate159inter10));
  nor2  gate1734(.a(gate159inter10), .b(gate159inter9), .O(gate159inter11));
  nor2  gate1735(.a(gate159inter11), .b(gate159inter6), .O(gate159inter12));
  nand2 gate1736(.a(gate159inter12), .b(gate159inter1), .O(G576));

  xor2  gate1261(.a(G531), .b(G447), .O(gate160inter0));
  nand2 gate1262(.a(gate160inter0), .b(s_102), .O(gate160inter1));
  and2  gate1263(.a(G531), .b(G447), .O(gate160inter2));
  inv1  gate1264(.a(s_102), .O(gate160inter3));
  inv1  gate1265(.a(s_103), .O(gate160inter4));
  nand2 gate1266(.a(gate160inter4), .b(gate160inter3), .O(gate160inter5));
  nor2  gate1267(.a(gate160inter5), .b(gate160inter2), .O(gate160inter6));
  inv1  gate1268(.a(G447), .O(gate160inter7));
  inv1  gate1269(.a(G531), .O(gate160inter8));
  nand2 gate1270(.a(gate160inter8), .b(gate160inter7), .O(gate160inter9));
  nand2 gate1271(.a(s_103), .b(gate160inter3), .O(gate160inter10));
  nor2  gate1272(.a(gate160inter10), .b(gate160inter9), .O(gate160inter11));
  nor2  gate1273(.a(gate160inter11), .b(gate160inter6), .O(gate160inter12));
  nand2 gate1274(.a(gate160inter12), .b(gate160inter1), .O(G577));
nand2 gate161( .a(G450), .b(G534), .O(G578) );
nand2 gate162( .a(G453), .b(G534), .O(G579) );
nand2 gate163( .a(G456), .b(G537), .O(G580) );
nand2 gate164( .a(G459), .b(G537), .O(G581) );

  xor2  gate1653(.a(G540), .b(G462), .O(gate165inter0));
  nand2 gate1654(.a(gate165inter0), .b(s_158), .O(gate165inter1));
  and2  gate1655(.a(G540), .b(G462), .O(gate165inter2));
  inv1  gate1656(.a(s_158), .O(gate165inter3));
  inv1  gate1657(.a(s_159), .O(gate165inter4));
  nand2 gate1658(.a(gate165inter4), .b(gate165inter3), .O(gate165inter5));
  nor2  gate1659(.a(gate165inter5), .b(gate165inter2), .O(gate165inter6));
  inv1  gate1660(.a(G462), .O(gate165inter7));
  inv1  gate1661(.a(G540), .O(gate165inter8));
  nand2 gate1662(.a(gate165inter8), .b(gate165inter7), .O(gate165inter9));
  nand2 gate1663(.a(s_159), .b(gate165inter3), .O(gate165inter10));
  nor2  gate1664(.a(gate165inter10), .b(gate165inter9), .O(gate165inter11));
  nor2  gate1665(.a(gate165inter11), .b(gate165inter6), .O(gate165inter12));
  nand2 gate1666(.a(gate165inter12), .b(gate165inter1), .O(G582));

  xor2  gate2633(.a(G540), .b(G465), .O(gate166inter0));
  nand2 gate2634(.a(gate166inter0), .b(s_298), .O(gate166inter1));
  and2  gate2635(.a(G540), .b(G465), .O(gate166inter2));
  inv1  gate2636(.a(s_298), .O(gate166inter3));
  inv1  gate2637(.a(s_299), .O(gate166inter4));
  nand2 gate2638(.a(gate166inter4), .b(gate166inter3), .O(gate166inter5));
  nor2  gate2639(.a(gate166inter5), .b(gate166inter2), .O(gate166inter6));
  inv1  gate2640(.a(G465), .O(gate166inter7));
  inv1  gate2641(.a(G540), .O(gate166inter8));
  nand2 gate2642(.a(gate166inter8), .b(gate166inter7), .O(gate166inter9));
  nand2 gate2643(.a(s_299), .b(gate166inter3), .O(gate166inter10));
  nor2  gate2644(.a(gate166inter10), .b(gate166inter9), .O(gate166inter11));
  nor2  gate2645(.a(gate166inter11), .b(gate166inter6), .O(gate166inter12));
  nand2 gate2646(.a(gate166inter12), .b(gate166inter1), .O(G583));

  xor2  gate1597(.a(G543), .b(G468), .O(gate167inter0));
  nand2 gate1598(.a(gate167inter0), .b(s_150), .O(gate167inter1));
  and2  gate1599(.a(G543), .b(G468), .O(gate167inter2));
  inv1  gate1600(.a(s_150), .O(gate167inter3));
  inv1  gate1601(.a(s_151), .O(gate167inter4));
  nand2 gate1602(.a(gate167inter4), .b(gate167inter3), .O(gate167inter5));
  nor2  gate1603(.a(gate167inter5), .b(gate167inter2), .O(gate167inter6));
  inv1  gate1604(.a(G468), .O(gate167inter7));
  inv1  gate1605(.a(G543), .O(gate167inter8));
  nand2 gate1606(.a(gate167inter8), .b(gate167inter7), .O(gate167inter9));
  nand2 gate1607(.a(s_151), .b(gate167inter3), .O(gate167inter10));
  nor2  gate1608(.a(gate167inter10), .b(gate167inter9), .O(gate167inter11));
  nor2  gate1609(.a(gate167inter11), .b(gate167inter6), .O(gate167inter12));
  nand2 gate1610(.a(gate167inter12), .b(gate167inter1), .O(G584));
nand2 gate168( .a(G471), .b(G543), .O(G585) );
nand2 gate169( .a(G474), .b(G546), .O(G586) );
nand2 gate170( .a(G477), .b(G546), .O(G587) );
nand2 gate171( .a(G480), .b(G549), .O(G588) );
nand2 gate172( .a(G483), .b(G549), .O(G589) );

  xor2  gate897(.a(G552), .b(G486), .O(gate173inter0));
  nand2 gate898(.a(gate173inter0), .b(s_50), .O(gate173inter1));
  and2  gate899(.a(G552), .b(G486), .O(gate173inter2));
  inv1  gate900(.a(s_50), .O(gate173inter3));
  inv1  gate901(.a(s_51), .O(gate173inter4));
  nand2 gate902(.a(gate173inter4), .b(gate173inter3), .O(gate173inter5));
  nor2  gate903(.a(gate173inter5), .b(gate173inter2), .O(gate173inter6));
  inv1  gate904(.a(G486), .O(gate173inter7));
  inv1  gate905(.a(G552), .O(gate173inter8));
  nand2 gate906(.a(gate173inter8), .b(gate173inter7), .O(gate173inter9));
  nand2 gate907(.a(s_51), .b(gate173inter3), .O(gate173inter10));
  nor2  gate908(.a(gate173inter10), .b(gate173inter9), .O(gate173inter11));
  nor2  gate909(.a(gate173inter11), .b(gate173inter6), .O(gate173inter12));
  nand2 gate910(.a(gate173inter12), .b(gate173inter1), .O(G590));
nand2 gate174( .a(G489), .b(G552), .O(G591) );
nand2 gate175( .a(G492), .b(G555), .O(G592) );
nand2 gate176( .a(G495), .b(G555), .O(G593) );
nand2 gate177( .a(G498), .b(G558), .O(G594) );
nand2 gate178( .a(G501), .b(G558), .O(G595) );
nand2 gate179( .a(G504), .b(G561), .O(G596) );

  xor2  gate2283(.a(G561), .b(G507), .O(gate180inter0));
  nand2 gate2284(.a(gate180inter0), .b(s_248), .O(gate180inter1));
  and2  gate2285(.a(G561), .b(G507), .O(gate180inter2));
  inv1  gate2286(.a(s_248), .O(gate180inter3));
  inv1  gate2287(.a(s_249), .O(gate180inter4));
  nand2 gate2288(.a(gate180inter4), .b(gate180inter3), .O(gate180inter5));
  nor2  gate2289(.a(gate180inter5), .b(gate180inter2), .O(gate180inter6));
  inv1  gate2290(.a(G507), .O(gate180inter7));
  inv1  gate2291(.a(G561), .O(gate180inter8));
  nand2 gate2292(.a(gate180inter8), .b(gate180inter7), .O(gate180inter9));
  nand2 gate2293(.a(s_249), .b(gate180inter3), .O(gate180inter10));
  nor2  gate2294(.a(gate180inter10), .b(gate180inter9), .O(gate180inter11));
  nor2  gate2295(.a(gate180inter11), .b(gate180inter6), .O(gate180inter12));
  nand2 gate2296(.a(gate180inter12), .b(gate180inter1), .O(G597));
nand2 gate181( .a(G510), .b(G564), .O(G598) );
nand2 gate182( .a(G513), .b(G564), .O(G599) );
nand2 gate183( .a(G516), .b(G567), .O(G600) );

  xor2  gate1079(.a(G567), .b(G519), .O(gate184inter0));
  nand2 gate1080(.a(gate184inter0), .b(s_76), .O(gate184inter1));
  and2  gate1081(.a(G567), .b(G519), .O(gate184inter2));
  inv1  gate1082(.a(s_76), .O(gate184inter3));
  inv1  gate1083(.a(s_77), .O(gate184inter4));
  nand2 gate1084(.a(gate184inter4), .b(gate184inter3), .O(gate184inter5));
  nor2  gate1085(.a(gate184inter5), .b(gate184inter2), .O(gate184inter6));
  inv1  gate1086(.a(G519), .O(gate184inter7));
  inv1  gate1087(.a(G567), .O(gate184inter8));
  nand2 gate1088(.a(gate184inter8), .b(gate184inter7), .O(gate184inter9));
  nand2 gate1089(.a(s_77), .b(gate184inter3), .O(gate184inter10));
  nor2  gate1090(.a(gate184inter10), .b(gate184inter9), .O(gate184inter11));
  nor2  gate1091(.a(gate184inter11), .b(gate184inter6), .O(gate184inter12));
  nand2 gate1092(.a(gate184inter12), .b(gate184inter1), .O(G601));
nand2 gate185( .a(G570), .b(G571), .O(G602) );

  xor2  gate1009(.a(G573), .b(G572), .O(gate186inter0));
  nand2 gate1010(.a(gate186inter0), .b(s_66), .O(gate186inter1));
  and2  gate1011(.a(G573), .b(G572), .O(gate186inter2));
  inv1  gate1012(.a(s_66), .O(gate186inter3));
  inv1  gate1013(.a(s_67), .O(gate186inter4));
  nand2 gate1014(.a(gate186inter4), .b(gate186inter3), .O(gate186inter5));
  nor2  gate1015(.a(gate186inter5), .b(gate186inter2), .O(gate186inter6));
  inv1  gate1016(.a(G572), .O(gate186inter7));
  inv1  gate1017(.a(G573), .O(gate186inter8));
  nand2 gate1018(.a(gate186inter8), .b(gate186inter7), .O(gate186inter9));
  nand2 gate1019(.a(s_67), .b(gate186inter3), .O(gate186inter10));
  nor2  gate1020(.a(gate186inter10), .b(gate186inter9), .O(gate186inter11));
  nor2  gate1021(.a(gate186inter11), .b(gate186inter6), .O(gate186inter12));
  nand2 gate1022(.a(gate186inter12), .b(gate186inter1), .O(G607));
nand2 gate187( .a(G574), .b(G575), .O(G612) );
nand2 gate188( .a(G576), .b(G577), .O(G617) );
nand2 gate189( .a(G578), .b(G579), .O(G622) );
nand2 gate190( .a(G580), .b(G581), .O(G627) );
nand2 gate191( .a(G582), .b(G583), .O(G632) );
nand2 gate192( .a(G584), .b(G585), .O(G637) );
nand2 gate193( .a(G586), .b(G587), .O(G642) );
nand2 gate194( .a(G588), .b(G589), .O(G645) );

  xor2  gate2185(.a(G591), .b(G590), .O(gate195inter0));
  nand2 gate2186(.a(gate195inter0), .b(s_234), .O(gate195inter1));
  and2  gate2187(.a(G591), .b(G590), .O(gate195inter2));
  inv1  gate2188(.a(s_234), .O(gate195inter3));
  inv1  gate2189(.a(s_235), .O(gate195inter4));
  nand2 gate2190(.a(gate195inter4), .b(gate195inter3), .O(gate195inter5));
  nor2  gate2191(.a(gate195inter5), .b(gate195inter2), .O(gate195inter6));
  inv1  gate2192(.a(G590), .O(gate195inter7));
  inv1  gate2193(.a(G591), .O(gate195inter8));
  nand2 gate2194(.a(gate195inter8), .b(gate195inter7), .O(gate195inter9));
  nand2 gate2195(.a(s_235), .b(gate195inter3), .O(gate195inter10));
  nor2  gate2196(.a(gate195inter10), .b(gate195inter9), .O(gate195inter11));
  nor2  gate2197(.a(gate195inter11), .b(gate195inter6), .O(gate195inter12));
  nand2 gate2198(.a(gate195inter12), .b(gate195inter1), .O(G648));

  xor2  gate1303(.a(G593), .b(G592), .O(gate196inter0));
  nand2 gate1304(.a(gate196inter0), .b(s_108), .O(gate196inter1));
  and2  gate1305(.a(G593), .b(G592), .O(gate196inter2));
  inv1  gate1306(.a(s_108), .O(gate196inter3));
  inv1  gate1307(.a(s_109), .O(gate196inter4));
  nand2 gate1308(.a(gate196inter4), .b(gate196inter3), .O(gate196inter5));
  nor2  gate1309(.a(gate196inter5), .b(gate196inter2), .O(gate196inter6));
  inv1  gate1310(.a(G592), .O(gate196inter7));
  inv1  gate1311(.a(G593), .O(gate196inter8));
  nand2 gate1312(.a(gate196inter8), .b(gate196inter7), .O(gate196inter9));
  nand2 gate1313(.a(s_109), .b(gate196inter3), .O(gate196inter10));
  nor2  gate1314(.a(gate196inter10), .b(gate196inter9), .O(gate196inter11));
  nor2  gate1315(.a(gate196inter11), .b(gate196inter6), .O(gate196inter12));
  nand2 gate1316(.a(gate196inter12), .b(gate196inter1), .O(G651));

  xor2  gate1107(.a(G595), .b(G594), .O(gate197inter0));
  nand2 gate1108(.a(gate197inter0), .b(s_80), .O(gate197inter1));
  and2  gate1109(.a(G595), .b(G594), .O(gate197inter2));
  inv1  gate1110(.a(s_80), .O(gate197inter3));
  inv1  gate1111(.a(s_81), .O(gate197inter4));
  nand2 gate1112(.a(gate197inter4), .b(gate197inter3), .O(gate197inter5));
  nor2  gate1113(.a(gate197inter5), .b(gate197inter2), .O(gate197inter6));
  inv1  gate1114(.a(G594), .O(gate197inter7));
  inv1  gate1115(.a(G595), .O(gate197inter8));
  nand2 gate1116(.a(gate197inter8), .b(gate197inter7), .O(gate197inter9));
  nand2 gate1117(.a(s_81), .b(gate197inter3), .O(gate197inter10));
  nor2  gate1118(.a(gate197inter10), .b(gate197inter9), .O(gate197inter11));
  nor2  gate1119(.a(gate197inter11), .b(gate197inter6), .O(gate197inter12));
  nand2 gate1120(.a(gate197inter12), .b(gate197inter1), .O(G654));

  xor2  gate1093(.a(G597), .b(G596), .O(gate198inter0));
  nand2 gate1094(.a(gate198inter0), .b(s_78), .O(gate198inter1));
  and2  gate1095(.a(G597), .b(G596), .O(gate198inter2));
  inv1  gate1096(.a(s_78), .O(gate198inter3));
  inv1  gate1097(.a(s_79), .O(gate198inter4));
  nand2 gate1098(.a(gate198inter4), .b(gate198inter3), .O(gate198inter5));
  nor2  gate1099(.a(gate198inter5), .b(gate198inter2), .O(gate198inter6));
  inv1  gate1100(.a(G596), .O(gate198inter7));
  inv1  gate1101(.a(G597), .O(gate198inter8));
  nand2 gate1102(.a(gate198inter8), .b(gate198inter7), .O(gate198inter9));
  nand2 gate1103(.a(s_79), .b(gate198inter3), .O(gate198inter10));
  nor2  gate1104(.a(gate198inter10), .b(gate198inter9), .O(gate198inter11));
  nor2  gate1105(.a(gate198inter11), .b(gate198inter6), .O(gate198inter12));
  nand2 gate1106(.a(gate198inter12), .b(gate198inter1), .O(G657));

  xor2  gate2605(.a(G599), .b(G598), .O(gate199inter0));
  nand2 gate2606(.a(gate199inter0), .b(s_294), .O(gate199inter1));
  and2  gate2607(.a(G599), .b(G598), .O(gate199inter2));
  inv1  gate2608(.a(s_294), .O(gate199inter3));
  inv1  gate2609(.a(s_295), .O(gate199inter4));
  nand2 gate2610(.a(gate199inter4), .b(gate199inter3), .O(gate199inter5));
  nor2  gate2611(.a(gate199inter5), .b(gate199inter2), .O(gate199inter6));
  inv1  gate2612(.a(G598), .O(gate199inter7));
  inv1  gate2613(.a(G599), .O(gate199inter8));
  nand2 gate2614(.a(gate199inter8), .b(gate199inter7), .O(gate199inter9));
  nand2 gate2615(.a(s_295), .b(gate199inter3), .O(gate199inter10));
  nor2  gate2616(.a(gate199inter10), .b(gate199inter9), .O(gate199inter11));
  nor2  gate2617(.a(gate199inter11), .b(gate199inter6), .O(gate199inter12));
  nand2 gate2618(.a(gate199inter12), .b(gate199inter1), .O(G660));
nand2 gate200( .a(G600), .b(G601), .O(G663) );
nand2 gate201( .a(G602), .b(G607), .O(G666) );

  xor2  gate2423(.a(G617), .b(G612), .O(gate202inter0));
  nand2 gate2424(.a(gate202inter0), .b(s_268), .O(gate202inter1));
  and2  gate2425(.a(G617), .b(G612), .O(gate202inter2));
  inv1  gate2426(.a(s_268), .O(gate202inter3));
  inv1  gate2427(.a(s_269), .O(gate202inter4));
  nand2 gate2428(.a(gate202inter4), .b(gate202inter3), .O(gate202inter5));
  nor2  gate2429(.a(gate202inter5), .b(gate202inter2), .O(gate202inter6));
  inv1  gate2430(.a(G612), .O(gate202inter7));
  inv1  gate2431(.a(G617), .O(gate202inter8));
  nand2 gate2432(.a(gate202inter8), .b(gate202inter7), .O(gate202inter9));
  nand2 gate2433(.a(s_269), .b(gate202inter3), .O(gate202inter10));
  nor2  gate2434(.a(gate202inter10), .b(gate202inter9), .O(gate202inter11));
  nor2  gate2435(.a(gate202inter11), .b(gate202inter6), .O(gate202inter12));
  nand2 gate2436(.a(gate202inter12), .b(gate202inter1), .O(G669));

  xor2  gate1611(.a(G612), .b(G602), .O(gate203inter0));
  nand2 gate1612(.a(gate203inter0), .b(s_152), .O(gate203inter1));
  and2  gate1613(.a(G612), .b(G602), .O(gate203inter2));
  inv1  gate1614(.a(s_152), .O(gate203inter3));
  inv1  gate1615(.a(s_153), .O(gate203inter4));
  nand2 gate1616(.a(gate203inter4), .b(gate203inter3), .O(gate203inter5));
  nor2  gate1617(.a(gate203inter5), .b(gate203inter2), .O(gate203inter6));
  inv1  gate1618(.a(G602), .O(gate203inter7));
  inv1  gate1619(.a(G612), .O(gate203inter8));
  nand2 gate1620(.a(gate203inter8), .b(gate203inter7), .O(gate203inter9));
  nand2 gate1621(.a(s_153), .b(gate203inter3), .O(gate203inter10));
  nor2  gate1622(.a(gate203inter10), .b(gate203inter9), .O(gate203inter11));
  nor2  gate1623(.a(gate203inter11), .b(gate203inter6), .O(gate203inter12));
  nand2 gate1624(.a(gate203inter12), .b(gate203inter1), .O(G672));
nand2 gate204( .a(G607), .b(G617), .O(G675) );

  xor2  gate1849(.a(G627), .b(G622), .O(gate205inter0));
  nand2 gate1850(.a(gate205inter0), .b(s_186), .O(gate205inter1));
  and2  gate1851(.a(G627), .b(G622), .O(gate205inter2));
  inv1  gate1852(.a(s_186), .O(gate205inter3));
  inv1  gate1853(.a(s_187), .O(gate205inter4));
  nand2 gate1854(.a(gate205inter4), .b(gate205inter3), .O(gate205inter5));
  nor2  gate1855(.a(gate205inter5), .b(gate205inter2), .O(gate205inter6));
  inv1  gate1856(.a(G622), .O(gate205inter7));
  inv1  gate1857(.a(G627), .O(gate205inter8));
  nand2 gate1858(.a(gate205inter8), .b(gate205inter7), .O(gate205inter9));
  nand2 gate1859(.a(s_187), .b(gate205inter3), .O(gate205inter10));
  nor2  gate1860(.a(gate205inter10), .b(gate205inter9), .O(gate205inter11));
  nor2  gate1861(.a(gate205inter11), .b(gate205inter6), .O(gate205inter12));
  nand2 gate1862(.a(gate205inter12), .b(gate205inter1), .O(G678));
nand2 gate206( .a(G632), .b(G637), .O(G681) );
nand2 gate207( .a(G622), .b(G632), .O(G684) );

  xor2  gate673(.a(G637), .b(G627), .O(gate208inter0));
  nand2 gate674(.a(gate208inter0), .b(s_18), .O(gate208inter1));
  and2  gate675(.a(G637), .b(G627), .O(gate208inter2));
  inv1  gate676(.a(s_18), .O(gate208inter3));
  inv1  gate677(.a(s_19), .O(gate208inter4));
  nand2 gate678(.a(gate208inter4), .b(gate208inter3), .O(gate208inter5));
  nor2  gate679(.a(gate208inter5), .b(gate208inter2), .O(gate208inter6));
  inv1  gate680(.a(G627), .O(gate208inter7));
  inv1  gate681(.a(G637), .O(gate208inter8));
  nand2 gate682(.a(gate208inter8), .b(gate208inter7), .O(gate208inter9));
  nand2 gate683(.a(s_19), .b(gate208inter3), .O(gate208inter10));
  nor2  gate684(.a(gate208inter10), .b(gate208inter9), .O(gate208inter11));
  nor2  gate685(.a(gate208inter11), .b(gate208inter6), .O(gate208inter12));
  nand2 gate686(.a(gate208inter12), .b(gate208inter1), .O(G687));

  xor2  gate2647(.a(G666), .b(G602), .O(gate209inter0));
  nand2 gate2648(.a(gate209inter0), .b(s_300), .O(gate209inter1));
  and2  gate2649(.a(G666), .b(G602), .O(gate209inter2));
  inv1  gate2650(.a(s_300), .O(gate209inter3));
  inv1  gate2651(.a(s_301), .O(gate209inter4));
  nand2 gate2652(.a(gate209inter4), .b(gate209inter3), .O(gate209inter5));
  nor2  gate2653(.a(gate209inter5), .b(gate209inter2), .O(gate209inter6));
  inv1  gate2654(.a(G602), .O(gate209inter7));
  inv1  gate2655(.a(G666), .O(gate209inter8));
  nand2 gate2656(.a(gate209inter8), .b(gate209inter7), .O(gate209inter9));
  nand2 gate2657(.a(s_301), .b(gate209inter3), .O(gate209inter10));
  nor2  gate2658(.a(gate209inter10), .b(gate209inter9), .O(gate209inter11));
  nor2  gate2659(.a(gate209inter11), .b(gate209inter6), .O(gate209inter12));
  nand2 gate2660(.a(gate209inter12), .b(gate209inter1), .O(G690));

  xor2  gate799(.a(G666), .b(G607), .O(gate210inter0));
  nand2 gate800(.a(gate210inter0), .b(s_36), .O(gate210inter1));
  and2  gate801(.a(G666), .b(G607), .O(gate210inter2));
  inv1  gate802(.a(s_36), .O(gate210inter3));
  inv1  gate803(.a(s_37), .O(gate210inter4));
  nand2 gate804(.a(gate210inter4), .b(gate210inter3), .O(gate210inter5));
  nor2  gate805(.a(gate210inter5), .b(gate210inter2), .O(gate210inter6));
  inv1  gate806(.a(G607), .O(gate210inter7));
  inv1  gate807(.a(G666), .O(gate210inter8));
  nand2 gate808(.a(gate210inter8), .b(gate210inter7), .O(gate210inter9));
  nand2 gate809(.a(s_37), .b(gate210inter3), .O(gate210inter10));
  nor2  gate810(.a(gate210inter10), .b(gate210inter9), .O(gate210inter11));
  nor2  gate811(.a(gate210inter11), .b(gate210inter6), .O(gate210inter12));
  nand2 gate812(.a(gate210inter12), .b(gate210inter1), .O(G691));
nand2 gate211( .a(G612), .b(G669), .O(G692) );
nand2 gate212( .a(G617), .b(G669), .O(G693) );

  xor2  gate2857(.a(G672), .b(G602), .O(gate213inter0));
  nand2 gate2858(.a(gate213inter0), .b(s_330), .O(gate213inter1));
  and2  gate2859(.a(G672), .b(G602), .O(gate213inter2));
  inv1  gate2860(.a(s_330), .O(gate213inter3));
  inv1  gate2861(.a(s_331), .O(gate213inter4));
  nand2 gate2862(.a(gate213inter4), .b(gate213inter3), .O(gate213inter5));
  nor2  gate2863(.a(gate213inter5), .b(gate213inter2), .O(gate213inter6));
  inv1  gate2864(.a(G602), .O(gate213inter7));
  inv1  gate2865(.a(G672), .O(gate213inter8));
  nand2 gate2866(.a(gate213inter8), .b(gate213inter7), .O(gate213inter9));
  nand2 gate2867(.a(s_331), .b(gate213inter3), .O(gate213inter10));
  nor2  gate2868(.a(gate213inter10), .b(gate213inter9), .O(gate213inter11));
  nor2  gate2869(.a(gate213inter11), .b(gate213inter6), .O(gate213inter12));
  nand2 gate2870(.a(gate213inter12), .b(gate213inter1), .O(G694));
nand2 gate214( .a(G612), .b(G672), .O(G695) );
nand2 gate215( .a(G607), .b(G675), .O(G696) );
nand2 gate216( .a(G617), .b(G675), .O(G697) );
nand2 gate217( .a(G622), .b(G678), .O(G698) );
nand2 gate218( .a(G627), .b(G678), .O(G699) );
nand2 gate219( .a(G632), .b(G681), .O(G700) );
nand2 gate220( .a(G637), .b(G681), .O(G701) );
nand2 gate221( .a(G622), .b(G684), .O(G702) );
nand2 gate222( .a(G632), .b(G684), .O(G703) );
nand2 gate223( .a(G627), .b(G687), .O(G704) );

  xor2  gate2479(.a(G687), .b(G637), .O(gate224inter0));
  nand2 gate2480(.a(gate224inter0), .b(s_276), .O(gate224inter1));
  and2  gate2481(.a(G687), .b(G637), .O(gate224inter2));
  inv1  gate2482(.a(s_276), .O(gate224inter3));
  inv1  gate2483(.a(s_277), .O(gate224inter4));
  nand2 gate2484(.a(gate224inter4), .b(gate224inter3), .O(gate224inter5));
  nor2  gate2485(.a(gate224inter5), .b(gate224inter2), .O(gate224inter6));
  inv1  gate2486(.a(G637), .O(gate224inter7));
  inv1  gate2487(.a(G687), .O(gate224inter8));
  nand2 gate2488(.a(gate224inter8), .b(gate224inter7), .O(gate224inter9));
  nand2 gate2489(.a(s_277), .b(gate224inter3), .O(gate224inter10));
  nor2  gate2490(.a(gate224inter10), .b(gate224inter9), .O(gate224inter11));
  nor2  gate2491(.a(gate224inter11), .b(gate224inter6), .O(gate224inter12));
  nand2 gate2492(.a(gate224inter12), .b(gate224inter1), .O(G705));

  xor2  gate1317(.a(G691), .b(G690), .O(gate225inter0));
  nand2 gate1318(.a(gate225inter0), .b(s_110), .O(gate225inter1));
  and2  gate1319(.a(G691), .b(G690), .O(gate225inter2));
  inv1  gate1320(.a(s_110), .O(gate225inter3));
  inv1  gate1321(.a(s_111), .O(gate225inter4));
  nand2 gate1322(.a(gate225inter4), .b(gate225inter3), .O(gate225inter5));
  nor2  gate1323(.a(gate225inter5), .b(gate225inter2), .O(gate225inter6));
  inv1  gate1324(.a(G690), .O(gate225inter7));
  inv1  gate1325(.a(G691), .O(gate225inter8));
  nand2 gate1326(.a(gate225inter8), .b(gate225inter7), .O(gate225inter9));
  nand2 gate1327(.a(s_111), .b(gate225inter3), .O(gate225inter10));
  nor2  gate1328(.a(gate225inter10), .b(gate225inter9), .O(gate225inter11));
  nor2  gate1329(.a(gate225inter11), .b(gate225inter6), .O(gate225inter12));
  nand2 gate1330(.a(gate225inter12), .b(gate225inter1), .O(G706));

  xor2  gate1863(.a(G693), .b(G692), .O(gate226inter0));
  nand2 gate1864(.a(gate226inter0), .b(s_188), .O(gate226inter1));
  and2  gate1865(.a(G693), .b(G692), .O(gate226inter2));
  inv1  gate1866(.a(s_188), .O(gate226inter3));
  inv1  gate1867(.a(s_189), .O(gate226inter4));
  nand2 gate1868(.a(gate226inter4), .b(gate226inter3), .O(gate226inter5));
  nor2  gate1869(.a(gate226inter5), .b(gate226inter2), .O(gate226inter6));
  inv1  gate1870(.a(G692), .O(gate226inter7));
  inv1  gate1871(.a(G693), .O(gate226inter8));
  nand2 gate1872(.a(gate226inter8), .b(gate226inter7), .O(gate226inter9));
  nand2 gate1873(.a(s_189), .b(gate226inter3), .O(gate226inter10));
  nor2  gate1874(.a(gate226inter10), .b(gate226inter9), .O(gate226inter11));
  nor2  gate1875(.a(gate226inter11), .b(gate226inter6), .O(gate226inter12));
  nand2 gate1876(.a(gate226inter12), .b(gate226inter1), .O(G709));

  xor2  gate1233(.a(G695), .b(G694), .O(gate227inter0));
  nand2 gate1234(.a(gate227inter0), .b(s_98), .O(gate227inter1));
  and2  gate1235(.a(G695), .b(G694), .O(gate227inter2));
  inv1  gate1236(.a(s_98), .O(gate227inter3));
  inv1  gate1237(.a(s_99), .O(gate227inter4));
  nand2 gate1238(.a(gate227inter4), .b(gate227inter3), .O(gate227inter5));
  nor2  gate1239(.a(gate227inter5), .b(gate227inter2), .O(gate227inter6));
  inv1  gate1240(.a(G694), .O(gate227inter7));
  inv1  gate1241(.a(G695), .O(gate227inter8));
  nand2 gate1242(.a(gate227inter8), .b(gate227inter7), .O(gate227inter9));
  nand2 gate1243(.a(s_99), .b(gate227inter3), .O(gate227inter10));
  nor2  gate1244(.a(gate227inter10), .b(gate227inter9), .O(gate227inter11));
  nor2  gate1245(.a(gate227inter11), .b(gate227inter6), .O(gate227inter12));
  nand2 gate1246(.a(gate227inter12), .b(gate227inter1), .O(G712));
nand2 gate228( .a(G696), .b(G697), .O(G715) );

  xor2  gate1527(.a(G699), .b(G698), .O(gate229inter0));
  nand2 gate1528(.a(gate229inter0), .b(s_140), .O(gate229inter1));
  and2  gate1529(.a(G699), .b(G698), .O(gate229inter2));
  inv1  gate1530(.a(s_140), .O(gate229inter3));
  inv1  gate1531(.a(s_141), .O(gate229inter4));
  nand2 gate1532(.a(gate229inter4), .b(gate229inter3), .O(gate229inter5));
  nor2  gate1533(.a(gate229inter5), .b(gate229inter2), .O(gate229inter6));
  inv1  gate1534(.a(G698), .O(gate229inter7));
  inv1  gate1535(.a(G699), .O(gate229inter8));
  nand2 gate1536(.a(gate229inter8), .b(gate229inter7), .O(gate229inter9));
  nand2 gate1537(.a(s_141), .b(gate229inter3), .O(gate229inter10));
  nor2  gate1538(.a(gate229inter10), .b(gate229inter9), .O(gate229inter11));
  nor2  gate1539(.a(gate229inter11), .b(gate229inter6), .O(gate229inter12));
  nand2 gate1540(.a(gate229inter12), .b(gate229inter1), .O(G718));
nand2 gate230( .a(G700), .b(G701), .O(G721) );
nand2 gate231( .a(G702), .b(G703), .O(G724) );
nand2 gate232( .a(G704), .b(G705), .O(G727) );
nand2 gate233( .a(G242), .b(G718), .O(G730) );
nand2 gate234( .a(G245), .b(G721), .O(G733) );

  xor2  gate869(.a(G724), .b(G248), .O(gate235inter0));
  nand2 gate870(.a(gate235inter0), .b(s_46), .O(gate235inter1));
  and2  gate871(.a(G724), .b(G248), .O(gate235inter2));
  inv1  gate872(.a(s_46), .O(gate235inter3));
  inv1  gate873(.a(s_47), .O(gate235inter4));
  nand2 gate874(.a(gate235inter4), .b(gate235inter3), .O(gate235inter5));
  nor2  gate875(.a(gate235inter5), .b(gate235inter2), .O(gate235inter6));
  inv1  gate876(.a(G248), .O(gate235inter7));
  inv1  gate877(.a(G724), .O(gate235inter8));
  nand2 gate878(.a(gate235inter8), .b(gate235inter7), .O(gate235inter9));
  nand2 gate879(.a(s_47), .b(gate235inter3), .O(gate235inter10));
  nor2  gate880(.a(gate235inter10), .b(gate235inter9), .O(gate235inter11));
  nor2  gate881(.a(gate235inter11), .b(gate235inter6), .O(gate235inter12));
  nand2 gate882(.a(gate235inter12), .b(gate235inter1), .O(G736));

  xor2  gate2759(.a(G727), .b(G251), .O(gate236inter0));
  nand2 gate2760(.a(gate236inter0), .b(s_316), .O(gate236inter1));
  and2  gate2761(.a(G727), .b(G251), .O(gate236inter2));
  inv1  gate2762(.a(s_316), .O(gate236inter3));
  inv1  gate2763(.a(s_317), .O(gate236inter4));
  nand2 gate2764(.a(gate236inter4), .b(gate236inter3), .O(gate236inter5));
  nor2  gate2765(.a(gate236inter5), .b(gate236inter2), .O(gate236inter6));
  inv1  gate2766(.a(G251), .O(gate236inter7));
  inv1  gate2767(.a(G727), .O(gate236inter8));
  nand2 gate2768(.a(gate236inter8), .b(gate236inter7), .O(gate236inter9));
  nand2 gate2769(.a(s_317), .b(gate236inter3), .O(gate236inter10));
  nor2  gate2770(.a(gate236inter10), .b(gate236inter9), .O(gate236inter11));
  nor2  gate2771(.a(gate236inter11), .b(gate236inter6), .O(gate236inter12));
  nand2 gate2772(.a(gate236inter12), .b(gate236inter1), .O(G739));

  xor2  gate1933(.a(G706), .b(G254), .O(gate237inter0));
  nand2 gate1934(.a(gate237inter0), .b(s_198), .O(gate237inter1));
  and2  gate1935(.a(G706), .b(G254), .O(gate237inter2));
  inv1  gate1936(.a(s_198), .O(gate237inter3));
  inv1  gate1937(.a(s_199), .O(gate237inter4));
  nand2 gate1938(.a(gate237inter4), .b(gate237inter3), .O(gate237inter5));
  nor2  gate1939(.a(gate237inter5), .b(gate237inter2), .O(gate237inter6));
  inv1  gate1940(.a(G254), .O(gate237inter7));
  inv1  gate1941(.a(G706), .O(gate237inter8));
  nand2 gate1942(.a(gate237inter8), .b(gate237inter7), .O(gate237inter9));
  nand2 gate1943(.a(s_199), .b(gate237inter3), .O(gate237inter10));
  nor2  gate1944(.a(gate237inter10), .b(gate237inter9), .O(gate237inter11));
  nor2  gate1945(.a(gate237inter11), .b(gate237inter6), .O(gate237inter12));
  nand2 gate1946(.a(gate237inter12), .b(gate237inter1), .O(G742));
nand2 gate238( .a(G257), .b(G709), .O(G745) );
nand2 gate239( .a(G260), .b(G712), .O(G748) );
nand2 gate240( .a(G263), .b(G715), .O(G751) );
nand2 gate241( .a(G242), .b(G730), .O(G754) );
nand2 gate242( .a(G718), .b(G730), .O(G755) );
nand2 gate243( .a(G245), .b(G733), .O(G756) );

  xor2  gate911(.a(G733), .b(G721), .O(gate244inter0));
  nand2 gate912(.a(gate244inter0), .b(s_52), .O(gate244inter1));
  and2  gate913(.a(G733), .b(G721), .O(gate244inter2));
  inv1  gate914(.a(s_52), .O(gate244inter3));
  inv1  gate915(.a(s_53), .O(gate244inter4));
  nand2 gate916(.a(gate244inter4), .b(gate244inter3), .O(gate244inter5));
  nor2  gate917(.a(gate244inter5), .b(gate244inter2), .O(gate244inter6));
  inv1  gate918(.a(G721), .O(gate244inter7));
  inv1  gate919(.a(G733), .O(gate244inter8));
  nand2 gate920(.a(gate244inter8), .b(gate244inter7), .O(gate244inter9));
  nand2 gate921(.a(s_53), .b(gate244inter3), .O(gate244inter10));
  nor2  gate922(.a(gate244inter10), .b(gate244inter9), .O(gate244inter11));
  nor2  gate923(.a(gate244inter11), .b(gate244inter6), .O(gate244inter12));
  nand2 gate924(.a(gate244inter12), .b(gate244inter1), .O(G757));

  xor2  gate2521(.a(G736), .b(G248), .O(gate245inter0));
  nand2 gate2522(.a(gate245inter0), .b(s_282), .O(gate245inter1));
  and2  gate2523(.a(G736), .b(G248), .O(gate245inter2));
  inv1  gate2524(.a(s_282), .O(gate245inter3));
  inv1  gate2525(.a(s_283), .O(gate245inter4));
  nand2 gate2526(.a(gate245inter4), .b(gate245inter3), .O(gate245inter5));
  nor2  gate2527(.a(gate245inter5), .b(gate245inter2), .O(gate245inter6));
  inv1  gate2528(.a(G248), .O(gate245inter7));
  inv1  gate2529(.a(G736), .O(gate245inter8));
  nand2 gate2530(.a(gate245inter8), .b(gate245inter7), .O(gate245inter9));
  nand2 gate2531(.a(s_283), .b(gate245inter3), .O(gate245inter10));
  nor2  gate2532(.a(gate245inter10), .b(gate245inter9), .O(gate245inter11));
  nor2  gate2533(.a(gate245inter11), .b(gate245inter6), .O(gate245inter12));
  nand2 gate2534(.a(gate245inter12), .b(gate245inter1), .O(G758));
nand2 gate246( .a(G724), .b(G736), .O(G759) );

  xor2  gate2829(.a(G739), .b(G251), .O(gate247inter0));
  nand2 gate2830(.a(gate247inter0), .b(s_326), .O(gate247inter1));
  and2  gate2831(.a(G739), .b(G251), .O(gate247inter2));
  inv1  gate2832(.a(s_326), .O(gate247inter3));
  inv1  gate2833(.a(s_327), .O(gate247inter4));
  nand2 gate2834(.a(gate247inter4), .b(gate247inter3), .O(gate247inter5));
  nor2  gate2835(.a(gate247inter5), .b(gate247inter2), .O(gate247inter6));
  inv1  gate2836(.a(G251), .O(gate247inter7));
  inv1  gate2837(.a(G739), .O(gate247inter8));
  nand2 gate2838(.a(gate247inter8), .b(gate247inter7), .O(gate247inter9));
  nand2 gate2839(.a(s_327), .b(gate247inter3), .O(gate247inter10));
  nor2  gate2840(.a(gate247inter10), .b(gate247inter9), .O(gate247inter11));
  nor2  gate2841(.a(gate247inter11), .b(gate247inter6), .O(gate247inter12));
  nand2 gate2842(.a(gate247inter12), .b(gate247inter1), .O(G760));
nand2 gate248( .a(G727), .b(G739), .O(G761) );

  xor2  gate743(.a(G742), .b(G254), .O(gate249inter0));
  nand2 gate744(.a(gate249inter0), .b(s_28), .O(gate249inter1));
  and2  gate745(.a(G742), .b(G254), .O(gate249inter2));
  inv1  gate746(.a(s_28), .O(gate249inter3));
  inv1  gate747(.a(s_29), .O(gate249inter4));
  nand2 gate748(.a(gate249inter4), .b(gate249inter3), .O(gate249inter5));
  nor2  gate749(.a(gate249inter5), .b(gate249inter2), .O(gate249inter6));
  inv1  gate750(.a(G254), .O(gate249inter7));
  inv1  gate751(.a(G742), .O(gate249inter8));
  nand2 gate752(.a(gate249inter8), .b(gate249inter7), .O(gate249inter9));
  nand2 gate753(.a(s_29), .b(gate249inter3), .O(gate249inter10));
  nor2  gate754(.a(gate249inter10), .b(gate249inter9), .O(gate249inter11));
  nor2  gate755(.a(gate249inter11), .b(gate249inter6), .O(gate249inter12));
  nand2 gate756(.a(gate249inter12), .b(gate249inter1), .O(G762));

  xor2  gate561(.a(G742), .b(G706), .O(gate250inter0));
  nand2 gate562(.a(gate250inter0), .b(s_2), .O(gate250inter1));
  and2  gate563(.a(G742), .b(G706), .O(gate250inter2));
  inv1  gate564(.a(s_2), .O(gate250inter3));
  inv1  gate565(.a(s_3), .O(gate250inter4));
  nand2 gate566(.a(gate250inter4), .b(gate250inter3), .O(gate250inter5));
  nor2  gate567(.a(gate250inter5), .b(gate250inter2), .O(gate250inter6));
  inv1  gate568(.a(G706), .O(gate250inter7));
  inv1  gate569(.a(G742), .O(gate250inter8));
  nand2 gate570(.a(gate250inter8), .b(gate250inter7), .O(gate250inter9));
  nand2 gate571(.a(s_3), .b(gate250inter3), .O(gate250inter10));
  nor2  gate572(.a(gate250inter10), .b(gate250inter9), .O(gate250inter11));
  nor2  gate573(.a(gate250inter11), .b(gate250inter6), .O(gate250inter12));
  nand2 gate574(.a(gate250inter12), .b(gate250inter1), .O(G763));

  xor2  gate589(.a(G745), .b(G257), .O(gate251inter0));
  nand2 gate590(.a(gate251inter0), .b(s_6), .O(gate251inter1));
  and2  gate591(.a(G745), .b(G257), .O(gate251inter2));
  inv1  gate592(.a(s_6), .O(gate251inter3));
  inv1  gate593(.a(s_7), .O(gate251inter4));
  nand2 gate594(.a(gate251inter4), .b(gate251inter3), .O(gate251inter5));
  nor2  gate595(.a(gate251inter5), .b(gate251inter2), .O(gate251inter6));
  inv1  gate596(.a(G257), .O(gate251inter7));
  inv1  gate597(.a(G745), .O(gate251inter8));
  nand2 gate598(.a(gate251inter8), .b(gate251inter7), .O(gate251inter9));
  nand2 gate599(.a(s_7), .b(gate251inter3), .O(gate251inter10));
  nor2  gate600(.a(gate251inter10), .b(gate251inter9), .O(gate251inter11));
  nor2  gate601(.a(gate251inter11), .b(gate251inter6), .O(gate251inter12));
  nand2 gate602(.a(gate251inter12), .b(gate251inter1), .O(G764));

  xor2  gate2773(.a(G745), .b(G709), .O(gate252inter0));
  nand2 gate2774(.a(gate252inter0), .b(s_318), .O(gate252inter1));
  and2  gate2775(.a(G745), .b(G709), .O(gate252inter2));
  inv1  gate2776(.a(s_318), .O(gate252inter3));
  inv1  gate2777(.a(s_319), .O(gate252inter4));
  nand2 gate2778(.a(gate252inter4), .b(gate252inter3), .O(gate252inter5));
  nor2  gate2779(.a(gate252inter5), .b(gate252inter2), .O(gate252inter6));
  inv1  gate2780(.a(G709), .O(gate252inter7));
  inv1  gate2781(.a(G745), .O(gate252inter8));
  nand2 gate2782(.a(gate252inter8), .b(gate252inter7), .O(gate252inter9));
  nand2 gate2783(.a(s_319), .b(gate252inter3), .O(gate252inter10));
  nor2  gate2784(.a(gate252inter10), .b(gate252inter9), .O(gate252inter11));
  nor2  gate2785(.a(gate252inter11), .b(gate252inter6), .O(gate252inter12));
  nand2 gate2786(.a(gate252inter12), .b(gate252inter1), .O(G765));

  xor2  gate575(.a(G748), .b(G260), .O(gate253inter0));
  nand2 gate576(.a(gate253inter0), .b(s_4), .O(gate253inter1));
  and2  gate577(.a(G748), .b(G260), .O(gate253inter2));
  inv1  gate578(.a(s_4), .O(gate253inter3));
  inv1  gate579(.a(s_5), .O(gate253inter4));
  nand2 gate580(.a(gate253inter4), .b(gate253inter3), .O(gate253inter5));
  nor2  gate581(.a(gate253inter5), .b(gate253inter2), .O(gate253inter6));
  inv1  gate582(.a(G260), .O(gate253inter7));
  inv1  gate583(.a(G748), .O(gate253inter8));
  nand2 gate584(.a(gate253inter8), .b(gate253inter7), .O(gate253inter9));
  nand2 gate585(.a(s_5), .b(gate253inter3), .O(gate253inter10));
  nor2  gate586(.a(gate253inter10), .b(gate253inter9), .O(gate253inter11));
  nor2  gate587(.a(gate253inter11), .b(gate253inter6), .O(gate253inter12));
  nand2 gate588(.a(gate253inter12), .b(gate253inter1), .O(G766));
nand2 gate254( .a(G712), .b(G748), .O(G767) );

  xor2  gate2087(.a(G751), .b(G263), .O(gate255inter0));
  nand2 gate2088(.a(gate255inter0), .b(s_220), .O(gate255inter1));
  and2  gate2089(.a(G751), .b(G263), .O(gate255inter2));
  inv1  gate2090(.a(s_220), .O(gate255inter3));
  inv1  gate2091(.a(s_221), .O(gate255inter4));
  nand2 gate2092(.a(gate255inter4), .b(gate255inter3), .O(gate255inter5));
  nor2  gate2093(.a(gate255inter5), .b(gate255inter2), .O(gate255inter6));
  inv1  gate2094(.a(G263), .O(gate255inter7));
  inv1  gate2095(.a(G751), .O(gate255inter8));
  nand2 gate2096(.a(gate255inter8), .b(gate255inter7), .O(gate255inter9));
  nand2 gate2097(.a(s_221), .b(gate255inter3), .O(gate255inter10));
  nor2  gate2098(.a(gate255inter10), .b(gate255inter9), .O(gate255inter11));
  nor2  gate2099(.a(gate255inter11), .b(gate255inter6), .O(gate255inter12));
  nand2 gate2100(.a(gate255inter12), .b(gate255inter1), .O(G768));

  xor2  gate2269(.a(G751), .b(G715), .O(gate256inter0));
  nand2 gate2270(.a(gate256inter0), .b(s_246), .O(gate256inter1));
  and2  gate2271(.a(G751), .b(G715), .O(gate256inter2));
  inv1  gate2272(.a(s_246), .O(gate256inter3));
  inv1  gate2273(.a(s_247), .O(gate256inter4));
  nand2 gate2274(.a(gate256inter4), .b(gate256inter3), .O(gate256inter5));
  nor2  gate2275(.a(gate256inter5), .b(gate256inter2), .O(gate256inter6));
  inv1  gate2276(.a(G715), .O(gate256inter7));
  inv1  gate2277(.a(G751), .O(gate256inter8));
  nand2 gate2278(.a(gate256inter8), .b(gate256inter7), .O(gate256inter9));
  nand2 gate2279(.a(s_247), .b(gate256inter3), .O(gate256inter10));
  nor2  gate2280(.a(gate256inter10), .b(gate256inter9), .O(gate256inter11));
  nor2  gate2281(.a(gate256inter11), .b(gate256inter6), .O(gate256inter12));
  nand2 gate2282(.a(gate256inter12), .b(gate256inter1), .O(G769));

  xor2  gate1429(.a(G755), .b(G754), .O(gate257inter0));
  nand2 gate1430(.a(gate257inter0), .b(s_126), .O(gate257inter1));
  and2  gate1431(.a(G755), .b(G754), .O(gate257inter2));
  inv1  gate1432(.a(s_126), .O(gate257inter3));
  inv1  gate1433(.a(s_127), .O(gate257inter4));
  nand2 gate1434(.a(gate257inter4), .b(gate257inter3), .O(gate257inter5));
  nor2  gate1435(.a(gate257inter5), .b(gate257inter2), .O(gate257inter6));
  inv1  gate1436(.a(G754), .O(gate257inter7));
  inv1  gate1437(.a(G755), .O(gate257inter8));
  nand2 gate1438(.a(gate257inter8), .b(gate257inter7), .O(gate257inter9));
  nand2 gate1439(.a(s_127), .b(gate257inter3), .O(gate257inter10));
  nor2  gate1440(.a(gate257inter10), .b(gate257inter9), .O(gate257inter11));
  nor2  gate1441(.a(gate257inter11), .b(gate257inter6), .O(gate257inter12));
  nand2 gate1442(.a(gate257inter12), .b(gate257inter1), .O(G770));

  xor2  gate1359(.a(G757), .b(G756), .O(gate258inter0));
  nand2 gate1360(.a(gate258inter0), .b(s_116), .O(gate258inter1));
  and2  gate1361(.a(G757), .b(G756), .O(gate258inter2));
  inv1  gate1362(.a(s_116), .O(gate258inter3));
  inv1  gate1363(.a(s_117), .O(gate258inter4));
  nand2 gate1364(.a(gate258inter4), .b(gate258inter3), .O(gate258inter5));
  nor2  gate1365(.a(gate258inter5), .b(gate258inter2), .O(gate258inter6));
  inv1  gate1366(.a(G756), .O(gate258inter7));
  inv1  gate1367(.a(G757), .O(gate258inter8));
  nand2 gate1368(.a(gate258inter8), .b(gate258inter7), .O(gate258inter9));
  nand2 gate1369(.a(s_117), .b(gate258inter3), .O(gate258inter10));
  nor2  gate1370(.a(gate258inter10), .b(gate258inter9), .O(gate258inter11));
  nor2  gate1371(.a(gate258inter11), .b(gate258inter6), .O(gate258inter12));
  nand2 gate1372(.a(gate258inter12), .b(gate258inter1), .O(G773));
nand2 gate259( .a(G758), .b(G759), .O(G776) );
nand2 gate260( .a(G760), .b(G761), .O(G779) );
nand2 gate261( .a(G762), .b(G763), .O(G782) );
nand2 gate262( .a(G764), .b(G765), .O(G785) );
nand2 gate263( .a(G766), .b(G767), .O(G788) );

  xor2  gate1065(.a(G769), .b(G768), .O(gate264inter0));
  nand2 gate1066(.a(gate264inter0), .b(s_74), .O(gate264inter1));
  and2  gate1067(.a(G769), .b(G768), .O(gate264inter2));
  inv1  gate1068(.a(s_74), .O(gate264inter3));
  inv1  gate1069(.a(s_75), .O(gate264inter4));
  nand2 gate1070(.a(gate264inter4), .b(gate264inter3), .O(gate264inter5));
  nor2  gate1071(.a(gate264inter5), .b(gate264inter2), .O(gate264inter6));
  inv1  gate1072(.a(G768), .O(gate264inter7));
  inv1  gate1073(.a(G769), .O(gate264inter8));
  nand2 gate1074(.a(gate264inter8), .b(gate264inter7), .O(gate264inter9));
  nand2 gate1075(.a(s_75), .b(gate264inter3), .O(gate264inter10));
  nor2  gate1076(.a(gate264inter10), .b(gate264inter9), .O(gate264inter11));
  nor2  gate1077(.a(gate264inter11), .b(gate264inter6), .O(gate264inter12));
  nand2 gate1078(.a(gate264inter12), .b(gate264inter1), .O(G791));

  xor2  gate1499(.a(G770), .b(G642), .O(gate265inter0));
  nand2 gate1500(.a(gate265inter0), .b(s_136), .O(gate265inter1));
  and2  gate1501(.a(G770), .b(G642), .O(gate265inter2));
  inv1  gate1502(.a(s_136), .O(gate265inter3));
  inv1  gate1503(.a(s_137), .O(gate265inter4));
  nand2 gate1504(.a(gate265inter4), .b(gate265inter3), .O(gate265inter5));
  nor2  gate1505(.a(gate265inter5), .b(gate265inter2), .O(gate265inter6));
  inv1  gate1506(.a(G642), .O(gate265inter7));
  inv1  gate1507(.a(G770), .O(gate265inter8));
  nand2 gate1508(.a(gate265inter8), .b(gate265inter7), .O(gate265inter9));
  nand2 gate1509(.a(s_137), .b(gate265inter3), .O(gate265inter10));
  nor2  gate1510(.a(gate265inter10), .b(gate265inter9), .O(gate265inter11));
  nor2  gate1511(.a(gate265inter11), .b(gate265inter6), .O(gate265inter12));
  nand2 gate1512(.a(gate265inter12), .b(gate265inter1), .O(G794));
nand2 gate266( .a(G645), .b(G773), .O(G797) );

  xor2  gate2017(.a(G776), .b(G648), .O(gate267inter0));
  nand2 gate2018(.a(gate267inter0), .b(s_210), .O(gate267inter1));
  and2  gate2019(.a(G776), .b(G648), .O(gate267inter2));
  inv1  gate2020(.a(s_210), .O(gate267inter3));
  inv1  gate2021(.a(s_211), .O(gate267inter4));
  nand2 gate2022(.a(gate267inter4), .b(gate267inter3), .O(gate267inter5));
  nor2  gate2023(.a(gate267inter5), .b(gate267inter2), .O(gate267inter6));
  inv1  gate2024(.a(G648), .O(gate267inter7));
  inv1  gate2025(.a(G776), .O(gate267inter8));
  nand2 gate2026(.a(gate267inter8), .b(gate267inter7), .O(gate267inter9));
  nand2 gate2027(.a(s_211), .b(gate267inter3), .O(gate267inter10));
  nor2  gate2028(.a(gate267inter10), .b(gate267inter9), .O(gate267inter11));
  nor2  gate2029(.a(gate267inter11), .b(gate267inter6), .O(gate267inter12));
  nand2 gate2030(.a(gate267inter12), .b(gate267inter1), .O(G800));
nand2 gate268( .a(G651), .b(G779), .O(G803) );

  xor2  gate1639(.a(G782), .b(G654), .O(gate269inter0));
  nand2 gate1640(.a(gate269inter0), .b(s_156), .O(gate269inter1));
  and2  gate1641(.a(G782), .b(G654), .O(gate269inter2));
  inv1  gate1642(.a(s_156), .O(gate269inter3));
  inv1  gate1643(.a(s_157), .O(gate269inter4));
  nand2 gate1644(.a(gate269inter4), .b(gate269inter3), .O(gate269inter5));
  nor2  gate1645(.a(gate269inter5), .b(gate269inter2), .O(gate269inter6));
  inv1  gate1646(.a(G654), .O(gate269inter7));
  inv1  gate1647(.a(G782), .O(gate269inter8));
  nand2 gate1648(.a(gate269inter8), .b(gate269inter7), .O(gate269inter9));
  nand2 gate1649(.a(s_157), .b(gate269inter3), .O(gate269inter10));
  nor2  gate1650(.a(gate269inter10), .b(gate269inter9), .O(gate269inter11));
  nor2  gate1651(.a(gate269inter11), .b(gate269inter6), .O(gate269inter12));
  nand2 gate1652(.a(gate269inter12), .b(gate269inter1), .O(G806));
nand2 gate270( .a(G657), .b(G785), .O(G809) );

  xor2  gate1807(.a(G788), .b(G660), .O(gate271inter0));
  nand2 gate1808(.a(gate271inter0), .b(s_180), .O(gate271inter1));
  and2  gate1809(.a(G788), .b(G660), .O(gate271inter2));
  inv1  gate1810(.a(s_180), .O(gate271inter3));
  inv1  gate1811(.a(s_181), .O(gate271inter4));
  nand2 gate1812(.a(gate271inter4), .b(gate271inter3), .O(gate271inter5));
  nor2  gate1813(.a(gate271inter5), .b(gate271inter2), .O(gate271inter6));
  inv1  gate1814(.a(G660), .O(gate271inter7));
  inv1  gate1815(.a(G788), .O(gate271inter8));
  nand2 gate1816(.a(gate271inter8), .b(gate271inter7), .O(gate271inter9));
  nand2 gate1817(.a(s_181), .b(gate271inter3), .O(gate271inter10));
  nor2  gate1818(.a(gate271inter10), .b(gate271inter9), .O(gate271inter11));
  nor2  gate1819(.a(gate271inter11), .b(gate271inter6), .O(gate271inter12));
  nand2 gate1820(.a(gate271inter12), .b(gate271inter1), .O(G812));
nand2 gate272( .a(G663), .b(G791), .O(G815) );
nand2 gate273( .a(G642), .b(G794), .O(G818) );

  xor2  gate631(.a(G794), .b(G770), .O(gate274inter0));
  nand2 gate632(.a(gate274inter0), .b(s_12), .O(gate274inter1));
  and2  gate633(.a(G794), .b(G770), .O(gate274inter2));
  inv1  gate634(.a(s_12), .O(gate274inter3));
  inv1  gate635(.a(s_13), .O(gate274inter4));
  nand2 gate636(.a(gate274inter4), .b(gate274inter3), .O(gate274inter5));
  nor2  gate637(.a(gate274inter5), .b(gate274inter2), .O(gate274inter6));
  inv1  gate638(.a(G770), .O(gate274inter7));
  inv1  gate639(.a(G794), .O(gate274inter8));
  nand2 gate640(.a(gate274inter8), .b(gate274inter7), .O(gate274inter9));
  nand2 gate641(.a(s_13), .b(gate274inter3), .O(gate274inter10));
  nor2  gate642(.a(gate274inter10), .b(gate274inter9), .O(gate274inter11));
  nor2  gate643(.a(gate274inter11), .b(gate274inter6), .O(gate274inter12));
  nand2 gate644(.a(gate274inter12), .b(gate274inter1), .O(G819));
nand2 gate275( .a(G645), .b(G797), .O(G820) );
nand2 gate276( .a(G773), .b(G797), .O(G821) );

  xor2  gate1835(.a(G800), .b(G648), .O(gate277inter0));
  nand2 gate1836(.a(gate277inter0), .b(s_184), .O(gate277inter1));
  and2  gate1837(.a(G800), .b(G648), .O(gate277inter2));
  inv1  gate1838(.a(s_184), .O(gate277inter3));
  inv1  gate1839(.a(s_185), .O(gate277inter4));
  nand2 gate1840(.a(gate277inter4), .b(gate277inter3), .O(gate277inter5));
  nor2  gate1841(.a(gate277inter5), .b(gate277inter2), .O(gate277inter6));
  inv1  gate1842(.a(G648), .O(gate277inter7));
  inv1  gate1843(.a(G800), .O(gate277inter8));
  nand2 gate1844(.a(gate277inter8), .b(gate277inter7), .O(gate277inter9));
  nand2 gate1845(.a(s_185), .b(gate277inter3), .O(gate277inter10));
  nor2  gate1846(.a(gate277inter10), .b(gate277inter9), .O(gate277inter11));
  nor2  gate1847(.a(gate277inter11), .b(gate277inter6), .O(gate277inter12));
  nand2 gate1848(.a(gate277inter12), .b(gate277inter1), .O(G822));

  xor2  gate771(.a(G800), .b(G776), .O(gate278inter0));
  nand2 gate772(.a(gate278inter0), .b(s_32), .O(gate278inter1));
  and2  gate773(.a(G800), .b(G776), .O(gate278inter2));
  inv1  gate774(.a(s_32), .O(gate278inter3));
  inv1  gate775(.a(s_33), .O(gate278inter4));
  nand2 gate776(.a(gate278inter4), .b(gate278inter3), .O(gate278inter5));
  nor2  gate777(.a(gate278inter5), .b(gate278inter2), .O(gate278inter6));
  inv1  gate778(.a(G776), .O(gate278inter7));
  inv1  gate779(.a(G800), .O(gate278inter8));
  nand2 gate780(.a(gate278inter8), .b(gate278inter7), .O(gate278inter9));
  nand2 gate781(.a(s_33), .b(gate278inter3), .O(gate278inter10));
  nor2  gate782(.a(gate278inter10), .b(gate278inter9), .O(gate278inter11));
  nor2  gate783(.a(gate278inter11), .b(gate278inter6), .O(gate278inter12));
  nand2 gate784(.a(gate278inter12), .b(gate278inter1), .O(G823));

  xor2  gate1667(.a(G803), .b(G651), .O(gate279inter0));
  nand2 gate1668(.a(gate279inter0), .b(s_160), .O(gate279inter1));
  and2  gate1669(.a(G803), .b(G651), .O(gate279inter2));
  inv1  gate1670(.a(s_160), .O(gate279inter3));
  inv1  gate1671(.a(s_161), .O(gate279inter4));
  nand2 gate1672(.a(gate279inter4), .b(gate279inter3), .O(gate279inter5));
  nor2  gate1673(.a(gate279inter5), .b(gate279inter2), .O(gate279inter6));
  inv1  gate1674(.a(G651), .O(gate279inter7));
  inv1  gate1675(.a(G803), .O(gate279inter8));
  nand2 gate1676(.a(gate279inter8), .b(gate279inter7), .O(gate279inter9));
  nand2 gate1677(.a(s_161), .b(gate279inter3), .O(gate279inter10));
  nor2  gate1678(.a(gate279inter10), .b(gate279inter9), .O(gate279inter11));
  nor2  gate1679(.a(gate279inter11), .b(gate279inter6), .O(gate279inter12));
  nand2 gate1680(.a(gate279inter12), .b(gate279inter1), .O(G824));
nand2 gate280( .a(G779), .b(G803), .O(G825) );

  xor2  gate2535(.a(G806), .b(G654), .O(gate281inter0));
  nand2 gate2536(.a(gate281inter0), .b(s_284), .O(gate281inter1));
  and2  gate2537(.a(G806), .b(G654), .O(gate281inter2));
  inv1  gate2538(.a(s_284), .O(gate281inter3));
  inv1  gate2539(.a(s_285), .O(gate281inter4));
  nand2 gate2540(.a(gate281inter4), .b(gate281inter3), .O(gate281inter5));
  nor2  gate2541(.a(gate281inter5), .b(gate281inter2), .O(gate281inter6));
  inv1  gate2542(.a(G654), .O(gate281inter7));
  inv1  gate2543(.a(G806), .O(gate281inter8));
  nand2 gate2544(.a(gate281inter8), .b(gate281inter7), .O(gate281inter9));
  nand2 gate2545(.a(s_285), .b(gate281inter3), .O(gate281inter10));
  nor2  gate2546(.a(gate281inter10), .b(gate281inter9), .O(gate281inter11));
  nor2  gate2547(.a(gate281inter11), .b(gate281inter6), .O(gate281inter12));
  nand2 gate2548(.a(gate281inter12), .b(gate281inter1), .O(G826));

  xor2  gate883(.a(G806), .b(G782), .O(gate282inter0));
  nand2 gate884(.a(gate282inter0), .b(s_48), .O(gate282inter1));
  and2  gate885(.a(G806), .b(G782), .O(gate282inter2));
  inv1  gate886(.a(s_48), .O(gate282inter3));
  inv1  gate887(.a(s_49), .O(gate282inter4));
  nand2 gate888(.a(gate282inter4), .b(gate282inter3), .O(gate282inter5));
  nor2  gate889(.a(gate282inter5), .b(gate282inter2), .O(gate282inter6));
  inv1  gate890(.a(G782), .O(gate282inter7));
  inv1  gate891(.a(G806), .O(gate282inter8));
  nand2 gate892(.a(gate282inter8), .b(gate282inter7), .O(gate282inter9));
  nand2 gate893(.a(s_49), .b(gate282inter3), .O(gate282inter10));
  nor2  gate894(.a(gate282inter10), .b(gate282inter9), .O(gate282inter11));
  nor2  gate895(.a(gate282inter11), .b(gate282inter6), .O(gate282inter12));
  nand2 gate896(.a(gate282inter12), .b(gate282inter1), .O(G827));
nand2 gate283( .a(G657), .b(G809), .O(G828) );
nand2 gate284( .a(G785), .b(G809), .O(G829) );

  xor2  gate1345(.a(G812), .b(G660), .O(gate285inter0));
  nand2 gate1346(.a(gate285inter0), .b(s_114), .O(gate285inter1));
  and2  gate1347(.a(G812), .b(G660), .O(gate285inter2));
  inv1  gate1348(.a(s_114), .O(gate285inter3));
  inv1  gate1349(.a(s_115), .O(gate285inter4));
  nand2 gate1350(.a(gate285inter4), .b(gate285inter3), .O(gate285inter5));
  nor2  gate1351(.a(gate285inter5), .b(gate285inter2), .O(gate285inter6));
  inv1  gate1352(.a(G660), .O(gate285inter7));
  inv1  gate1353(.a(G812), .O(gate285inter8));
  nand2 gate1354(.a(gate285inter8), .b(gate285inter7), .O(gate285inter9));
  nand2 gate1355(.a(s_115), .b(gate285inter3), .O(gate285inter10));
  nor2  gate1356(.a(gate285inter10), .b(gate285inter9), .O(gate285inter11));
  nor2  gate1357(.a(gate285inter11), .b(gate285inter6), .O(gate285inter12));
  nand2 gate1358(.a(gate285inter12), .b(gate285inter1), .O(G830));

  xor2  gate1387(.a(G812), .b(G788), .O(gate286inter0));
  nand2 gate1388(.a(gate286inter0), .b(s_120), .O(gate286inter1));
  and2  gate1389(.a(G812), .b(G788), .O(gate286inter2));
  inv1  gate1390(.a(s_120), .O(gate286inter3));
  inv1  gate1391(.a(s_121), .O(gate286inter4));
  nand2 gate1392(.a(gate286inter4), .b(gate286inter3), .O(gate286inter5));
  nor2  gate1393(.a(gate286inter5), .b(gate286inter2), .O(gate286inter6));
  inv1  gate1394(.a(G788), .O(gate286inter7));
  inv1  gate1395(.a(G812), .O(gate286inter8));
  nand2 gate1396(.a(gate286inter8), .b(gate286inter7), .O(gate286inter9));
  nand2 gate1397(.a(s_121), .b(gate286inter3), .O(gate286inter10));
  nor2  gate1398(.a(gate286inter10), .b(gate286inter9), .O(gate286inter11));
  nor2  gate1399(.a(gate286inter11), .b(gate286inter6), .O(gate286inter12));
  nand2 gate1400(.a(gate286inter12), .b(gate286inter1), .O(G831));

  xor2  gate701(.a(G815), .b(G663), .O(gate287inter0));
  nand2 gate702(.a(gate287inter0), .b(s_22), .O(gate287inter1));
  and2  gate703(.a(G815), .b(G663), .O(gate287inter2));
  inv1  gate704(.a(s_22), .O(gate287inter3));
  inv1  gate705(.a(s_23), .O(gate287inter4));
  nand2 gate706(.a(gate287inter4), .b(gate287inter3), .O(gate287inter5));
  nor2  gate707(.a(gate287inter5), .b(gate287inter2), .O(gate287inter6));
  inv1  gate708(.a(G663), .O(gate287inter7));
  inv1  gate709(.a(G815), .O(gate287inter8));
  nand2 gate710(.a(gate287inter8), .b(gate287inter7), .O(gate287inter9));
  nand2 gate711(.a(s_23), .b(gate287inter3), .O(gate287inter10));
  nor2  gate712(.a(gate287inter10), .b(gate287inter9), .O(gate287inter11));
  nor2  gate713(.a(gate287inter11), .b(gate287inter6), .O(gate287inter12));
  nand2 gate714(.a(gate287inter12), .b(gate287inter1), .O(G832));
nand2 gate288( .a(G791), .b(G815), .O(G833) );
nand2 gate289( .a(G818), .b(G819), .O(G834) );

  xor2  gate1037(.a(G821), .b(G820), .O(gate290inter0));
  nand2 gate1038(.a(gate290inter0), .b(s_70), .O(gate290inter1));
  and2  gate1039(.a(G821), .b(G820), .O(gate290inter2));
  inv1  gate1040(.a(s_70), .O(gate290inter3));
  inv1  gate1041(.a(s_71), .O(gate290inter4));
  nand2 gate1042(.a(gate290inter4), .b(gate290inter3), .O(gate290inter5));
  nor2  gate1043(.a(gate290inter5), .b(gate290inter2), .O(gate290inter6));
  inv1  gate1044(.a(G820), .O(gate290inter7));
  inv1  gate1045(.a(G821), .O(gate290inter8));
  nand2 gate1046(.a(gate290inter8), .b(gate290inter7), .O(gate290inter9));
  nand2 gate1047(.a(s_71), .b(gate290inter3), .O(gate290inter10));
  nor2  gate1048(.a(gate290inter10), .b(gate290inter9), .O(gate290inter11));
  nor2  gate1049(.a(gate290inter11), .b(gate290inter6), .O(gate290inter12));
  nand2 gate1050(.a(gate290inter12), .b(gate290inter1), .O(G847));
nand2 gate291( .a(G822), .b(G823), .O(G860) );

  xor2  gate2073(.a(G825), .b(G824), .O(gate292inter0));
  nand2 gate2074(.a(gate292inter0), .b(s_218), .O(gate292inter1));
  and2  gate2075(.a(G825), .b(G824), .O(gate292inter2));
  inv1  gate2076(.a(s_218), .O(gate292inter3));
  inv1  gate2077(.a(s_219), .O(gate292inter4));
  nand2 gate2078(.a(gate292inter4), .b(gate292inter3), .O(gate292inter5));
  nor2  gate2079(.a(gate292inter5), .b(gate292inter2), .O(gate292inter6));
  inv1  gate2080(.a(G824), .O(gate292inter7));
  inv1  gate2081(.a(G825), .O(gate292inter8));
  nand2 gate2082(.a(gate292inter8), .b(gate292inter7), .O(gate292inter9));
  nand2 gate2083(.a(s_219), .b(gate292inter3), .O(gate292inter10));
  nor2  gate2084(.a(gate292inter10), .b(gate292inter9), .O(gate292inter11));
  nor2  gate2085(.a(gate292inter11), .b(gate292inter6), .O(gate292inter12));
  nand2 gate2086(.a(gate292inter12), .b(gate292inter1), .O(G873));
nand2 gate293( .a(G828), .b(G829), .O(G886) );
nand2 gate294( .a(G832), .b(G833), .O(G899) );
nand2 gate295( .a(G830), .b(G831), .O(G912) );
nand2 gate296( .a(G826), .b(G827), .O(G925) );
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );

  xor2  gate1121(.a(G1036), .b(G1), .O(gate387inter0));
  nand2 gate1122(.a(gate387inter0), .b(s_82), .O(gate387inter1));
  and2  gate1123(.a(G1036), .b(G1), .O(gate387inter2));
  inv1  gate1124(.a(s_82), .O(gate387inter3));
  inv1  gate1125(.a(s_83), .O(gate387inter4));
  nand2 gate1126(.a(gate387inter4), .b(gate387inter3), .O(gate387inter5));
  nor2  gate1127(.a(gate387inter5), .b(gate387inter2), .O(gate387inter6));
  inv1  gate1128(.a(G1), .O(gate387inter7));
  inv1  gate1129(.a(G1036), .O(gate387inter8));
  nand2 gate1130(.a(gate387inter8), .b(gate387inter7), .O(gate387inter9));
  nand2 gate1131(.a(s_83), .b(gate387inter3), .O(gate387inter10));
  nor2  gate1132(.a(gate387inter10), .b(gate387inter9), .O(gate387inter11));
  nor2  gate1133(.a(gate387inter11), .b(gate387inter6), .O(gate387inter12));
  nand2 gate1134(.a(gate387inter12), .b(gate387inter1), .O(G1132));

  xor2  gate1709(.a(G1039), .b(G2), .O(gate388inter0));
  nand2 gate1710(.a(gate388inter0), .b(s_166), .O(gate388inter1));
  and2  gate1711(.a(G1039), .b(G2), .O(gate388inter2));
  inv1  gate1712(.a(s_166), .O(gate388inter3));
  inv1  gate1713(.a(s_167), .O(gate388inter4));
  nand2 gate1714(.a(gate388inter4), .b(gate388inter3), .O(gate388inter5));
  nor2  gate1715(.a(gate388inter5), .b(gate388inter2), .O(gate388inter6));
  inv1  gate1716(.a(G2), .O(gate388inter7));
  inv1  gate1717(.a(G1039), .O(gate388inter8));
  nand2 gate1718(.a(gate388inter8), .b(gate388inter7), .O(gate388inter9));
  nand2 gate1719(.a(s_167), .b(gate388inter3), .O(gate388inter10));
  nor2  gate1720(.a(gate388inter10), .b(gate388inter9), .O(gate388inter11));
  nor2  gate1721(.a(gate388inter11), .b(gate388inter6), .O(gate388inter12));
  nand2 gate1722(.a(gate388inter12), .b(gate388inter1), .O(G1135));
nand2 gate389( .a(G3), .b(G1042), .O(G1138) );
nand2 gate390( .a(G4), .b(G1045), .O(G1141) );

  xor2  gate1289(.a(G1048), .b(G5), .O(gate391inter0));
  nand2 gate1290(.a(gate391inter0), .b(s_106), .O(gate391inter1));
  and2  gate1291(.a(G1048), .b(G5), .O(gate391inter2));
  inv1  gate1292(.a(s_106), .O(gate391inter3));
  inv1  gate1293(.a(s_107), .O(gate391inter4));
  nand2 gate1294(.a(gate391inter4), .b(gate391inter3), .O(gate391inter5));
  nor2  gate1295(.a(gate391inter5), .b(gate391inter2), .O(gate391inter6));
  inv1  gate1296(.a(G5), .O(gate391inter7));
  inv1  gate1297(.a(G1048), .O(gate391inter8));
  nand2 gate1298(.a(gate391inter8), .b(gate391inter7), .O(gate391inter9));
  nand2 gate1299(.a(s_107), .b(gate391inter3), .O(gate391inter10));
  nor2  gate1300(.a(gate391inter10), .b(gate391inter9), .O(gate391inter11));
  nor2  gate1301(.a(gate391inter11), .b(gate391inter6), .O(gate391inter12));
  nand2 gate1302(.a(gate391inter12), .b(gate391inter1), .O(G1144));

  xor2  gate1821(.a(G1051), .b(G6), .O(gate392inter0));
  nand2 gate1822(.a(gate392inter0), .b(s_182), .O(gate392inter1));
  and2  gate1823(.a(G1051), .b(G6), .O(gate392inter2));
  inv1  gate1824(.a(s_182), .O(gate392inter3));
  inv1  gate1825(.a(s_183), .O(gate392inter4));
  nand2 gate1826(.a(gate392inter4), .b(gate392inter3), .O(gate392inter5));
  nor2  gate1827(.a(gate392inter5), .b(gate392inter2), .O(gate392inter6));
  inv1  gate1828(.a(G6), .O(gate392inter7));
  inv1  gate1829(.a(G1051), .O(gate392inter8));
  nand2 gate1830(.a(gate392inter8), .b(gate392inter7), .O(gate392inter9));
  nand2 gate1831(.a(s_183), .b(gate392inter3), .O(gate392inter10));
  nor2  gate1832(.a(gate392inter10), .b(gate392inter9), .O(gate392inter11));
  nor2  gate1833(.a(gate392inter11), .b(gate392inter6), .O(gate392inter12));
  nand2 gate1834(.a(gate392inter12), .b(gate392inter1), .O(G1147));
nand2 gate393( .a(G7), .b(G1054), .O(G1150) );

  xor2  gate1051(.a(G1057), .b(G8), .O(gate394inter0));
  nand2 gate1052(.a(gate394inter0), .b(s_72), .O(gate394inter1));
  and2  gate1053(.a(G1057), .b(G8), .O(gate394inter2));
  inv1  gate1054(.a(s_72), .O(gate394inter3));
  inv1  gate1055(.a(s_73), .O(gate394inter4));
  nand2 gate1056(.a(gate394inter4), .b(gate394inter3), .O(gate394inter5));
  nor2  gate1057(.a(gate394inter5), .b(gate394inter2), .O(gate394inter6));
  inv1  gate1058(.a(G8), .O(gate394inter7));
  inv1  gate1059(.a(G1057), .O(gate394inter8));
  nand2 gate1060(.a(gate394inter8), .b(gate394inter7), .O(gate394inter9));
  nand2 gate1061(.a(s_73), .b(gate394inter3), .O(gate394inter10));
  nor2  gate1062(.a(gate394inter10), .b(gate394inter9), .O(gate394inter11));
  nor2  gate1063(.a(gate394inter11), .b(gate394inter6), .O(gate394inter12));
  nand2 gate1064(.a(gate394inter12), .b(gate394inter1), .O(G1153));
nand2 gate395( .a(G9), .b(G1060), .O(G1156) );

  xor2  gate1779(.a(G1063), .b(G10), .O(gate396inter0));
  nand2 gate1780(.a(gate396inter0), .b(s_176), .O(gate396inter1));
  and2  gate1781(.a(G1063), .b(G10), .O(gate396inter2));
  inv1  gate1782(.a(s_176), .O(gate396inter3));
  inv1  gate1783(.a(s_177), .O(gate396inter4));
  nand2 gate1784(.a(gate396inter4), .b(gate396inter3), .O(gate396inter5));
  nor2  gate1785(.a(gate396inter5), .b(gate396inter2), .O(gate396inter6));
  inv1  gate1786(.a(G10), .O(gate396inter7));
  inv1  gate1787(.a(G1063), .O(gate396inter8));
  nand2 gate1788(.a(gate396inter8), .b(gate396inter7), .O(gate396inter9));
  nand2 gate1789(.a(s_177), .b(gate396inter3), .O(gate396inter10));
  nor2  gate1790(.a(gate396inter10), .b(gate396inter9), .O(gate396inter11));
  nor2  gate1791(.a(gate396inter11), .b(gate396inter6), .O(gate396inter12));
  nand2 gate1792(.a(gate396inter12), .b(gate396inter1), .O(G1159));
nand2 gate397( .a(G11), .b(G1066), .O(G1162) );

  xor2  gate1541(.a(G1069), .b(G12), .O(gate398inter0));
  nand2 gate1542(.a(gate398inter0), .b(s_142), .O(gate398inter1));
  and2  gate1543(.a(G1069), .b(G12), .O(gate398inter2));
  inv1  gate1544(.a(s_142), .O(gate398inter3));
  inv1  gate1545(.a(s_143), .O(gate398inter4));
  nand2 gate1546(.a(gate398inter4), .b(gate398inter3), .O(gate398inter5));
  nor2  gate1547(.a(gate398inter5), .b(gate398inter2), .O(gate398inter6));
  inv1  gate1548(.a(G12), .O(gate398inter7));
  inv1  gate1549(.a(G1069), .O(gate398inter8));
  nand2 gate1550(.a(gate398inter8), .b(gate398inter7), .O(gate398inter9));
  nand2 gate1551(.a(s_143), .b(gate398inter3), .O(gate398inter10));
  nor2  gate1552(.a(gate398inter10), .b(gate398inter9), .O(gate398inter11));
  nor2  gate1553(.a(gate398inter11), .b(gate398inter6), .O(gate398inter12));
  nand2 gate1554(.a(gate398inter12), .b(gate398inter1), .O(G1165));

  xor2  gate1023(.a(G1072), .b(G13), .O(gate399inter0));
  nand2 gate1024(.a(gate399inter0), .b(s_68), .O(gate399inter1));
  and2  gate1025(.a(G1072), .b(G13), .O(gate399inter2));
  inv1  gate1026(.a(s_68), .O(gate399inter3));
  inv1  gate1027(.a(s_69), .O(gate399inter4));
  nand2 gate1028(.a(gate399inter4), .b(gate399inter3), .O(gate399inter5));
  nor2  gate1029(.a(gate399inter5), .b(gate399inter2), .O(gate399inter6));
  inv1  gate1030(.a(G13), .O(gate399inter7));
  inv1  gate1031(.a(G1072), .O(gate399inter8));
  nand2 gate1032(.a(gate399inter8), .b(gate399inter7), .O(gate399inter9));
  nand2 gate1033(.a(s_69), .b(gate399inter3), .O(gate399inter10));
  nor2  gate1034(.a(gate399inter10), .b(gate399inter9), .O(gate399inter11));
  nor2  gate1035(.a(gate399inter11), .b(gate399inter6), .O(gate399inter12));
  nand2 gate1036(.a(gate399inter12), .b(gate399inter1), .O(G1168));

  xor2  gate2143(.a(G1075), .b(G14), .O(gate400inter0));
  nand2 gate2144(.a(gate400inter0), .b(s_228), .O(gate400inter1));
  and2  gate2145(.a(G1075), .b(G14), .O(gate400inter2));
  inv1  gate2146(.a(s_228), .O(gate400inter3));
  inv1  gate2147(.a(s_229), .O(gate400inter4));
  nand2 gate2148(.a(gate400inter4), .b(gate400inter3), .O(gate400inter5));
  nor2  gate2149(.a(gate400inter5), .b(gate400inter2), .O(gate400inter6));
  inv1  gate2150(.a(G14), .O(gate400inter7));
  inv1  gate2151(.a(G1075), .O(gate400inter8));
  nand2 gate2152(.a(gate400inter8), .b(gate400inter7), .O(gate400inter9));
  nand2 gate2153(.a(s_229), .b(gate400inter3), .O(gate400inter10));
  nor2  gate2154(.a(gate400inter10), .b(gate400inter9), .O(gate400inter11));
  nor2  gate2155(.a(gate400inter11), .b(gate400inter6), .O(gate400inter12));
  nand2 gate2156(.a(gate400inter12), .b(gate400inter1), .O(G1171));
nand2 gate401( .a(G15), .b(G1078), .O(G1174) );
nand2 gate402( .a(G16), .b(G1081), .O(G1177) );
nand2 gate403( .a(G17), .b(G1084), .O(G1180) );
nand2 gate404( .a(G18), .b(G1087), .O(G1183) );
nand2 gate405( .a(G19), .b(G1090), .O(G1186) );
nand2 gate406( .a(G20), .b(G1093), .O(G1189) );

  xor2  gate1191(.a(G1096), .b(G21), .O(gate407inter0));
  nand2 gate1192(.a(gate407inter0), .b(s_92), .O(gate407inter1));
  and2  gate1193(.a(G1096), .b(G21), .O(gate407inter2));
  inv1  gate1194(.a(s_92), .O(gate407inter3));
  inv1  gate1195(.a(s_93), .O(gate407inter4));
  nand2 gate1196(.a(gate407inter4), .b(gate407inter3), .O(gate407inter5));
  nor2  gate1197(.a(gate407inter5), .b(gate407inter2), .O(gate407inter6));
  inv1  gate1198(.a(G21), .O(gate407inter7));
  inv1  gate1199(.a(G1096), .O(gate407inter8));
  nand2 gate1200(.a(gate407inter8), .b(gate407inter7), .O(gate407inter9));
  nand2 gate1201(.a(s_93), .b(gate407inter3), .O(gate407inter10));
  nor2  gate1202(.a(gate407inter10), .b(gate407inter9), .O(gate407inter11));
  nor2  gate1203(.a(gate407inter11), .b(gate407inter6), .O(gate407inter12));
  nand2 gate1204(.a(gate407inter12), .b(gate407inter1), .O(G1192));
nand2 gate408( .a(G22), .b(G1099), .O(G1195) );
nand2 gate409( .a(G23), .b(G1102), .O(G1198) );
nand2 gate410( .a(G24), .b(G1105), .O(G1201) );
nand2 gate411( .a(G25), .b(G1108), .O(G1204) );
nand2 gate412( .a(G26), .b(G1111), .O(G1207) );
nand2 gate413( .a(G27), .b(G1114), .O(G1210) );

  xor2  gate2549(.a(G1117), .b(G28), .O(gate414inter0));
  nand2 gate2550(.a(gate414inter0), .b(s_286), .O(gate414inter1));
  and2  gate2551(.a(G1117), .b(G28), .O(gate414inter2));
  inv1  gate2552(.a(s_286), .O(gate414inter3));
  inv1  gate2553(.a(s_287), .O(gate414inter4));
  nand2 gate2554(.a(gate414inter4), .b(gate414inter3), .O(gate414inter5));
  nor2  gate2555(.a(gate414inter5), .b(gate414inter2), .O(gate414inter6));
  inv1  gate2556(.a(G28), .O(gate414inter7));
  inv1  gate2557(.a(G1117), .O(gate414inter8));
  nand2 gate2558(.a(gate414inter8), .b(gate414inter7), .O(gate414inter9));
  nand2 gate2559(.a(s_287), .b(gate414inter3), .O(gate414inter10));
  nor2  gate2560(.a(gate414inter10), .b(gate414inter9), .O(gate414inter11));
  nor2  gate2561(.a(gate414inter11), .b(gate414inter6), .O(gate414inter12));
  nand2 gate2562(.a(gate414inter12), .b(gate414inter1), .O(G1213));
nand2 gate415( .a(G29), .b(G1120), .O(G1216) );
nand2 gate416( .a(G30), .b(G1123), .O(G1219) );
nand2 gate417( .a(G31), .b(G1126), .O(G1222) );
nand2 gate418( .a(G32), .b(G1129), .O(G1225) );
nand2 gate419( .a(G1), .b(G1132), .O(G1228) );
nand2 gate420( .a(G1036), .b(G1132), .O(G1229) );
nand2 gate421( .a(G2), .b(G1135), .O(G1230) );

  xor2  gate2367(.a(G1135), .b(G1039), .O(gate422inter0));
  nand2 gate2368(.a(gate422inter0), .b(s_260), .O(gate422inter1));
  and2  gate2369(.a(G1135), .b(G1039), .O(gate422inter2));
  inv1  gate2370(.a(s_260), .O(gate422inter3));
  inv1  gate2371(.a(s_261), .O(gate422inter4));
  nand2 gate2372(.a(gate422inter4), .b(gate422inter3), .O(gate422inter5));
  nor2  gate2373(.a(gate422inter5), .b(gate422inter2), .O(gate422inter6));
  inv1  gate2374(.a(G1039), .O(gate422inter7));
  inv1  gate2375(.a(G1135), .O(gate422inter8));
  nand2 gate2376(.a(gate422inter8), .b(gate422inter7), .O(gate422inter9));
  nand2 gate2377(.a(s_261), .b(gate422inter3), .O(gate422inter10));
  nor2  gate2378(.a(gate422inter10), .b(gate422inter9), .O(gate422inter11));
  nor2  gate2379(.a(gate422inter11), .b(gate422inter6), .O(gate422inter12));
  nand2 gate2380(.a(gate422inter12), .b(gate422inter1), .O(G1231));
nand2 gate423( .a(G3), .b(G1138), .O(G1232) );
nand2 gate424( .a(G1042), .b(G1138), .O(G1233) );
nand2 gate425( .a(G4), .b(G1141), .O(G1234) );
nand2 gate426( .a(G1045), .b(G1141), .O(G1235) );

  xor2  gate2339(.a(G1144), .b(G5), .O(gate427inter0));
  nand2 gate2340(.a(gate427inter0), .b(s_256), .O(gate427inter1));
  and2  gate2341(.a(G1144), .b(G5), .O(gate427inter2));
  inv1  gate2342(.a(s_256), .O(gate427inter3));
  inv1  gate2343(.a(s_257), .O(gate427inter4));
  nand2 gate2344(.a(gate427inter4), .b(gate427inter3), .O(gate427inter5));
  nor2  gate2345(.a(gate427inter5), .b(gate427inter2), .O(gate427inter6));
  inv1  gate2346(.a(G5), .O(gate427inter7));
  inv1  gate2347(.a(G1144), .O(gate427inter8));
  nand2 gate2348(.a(gate427inter8), .b(gate427inter7), .O(gate427inter9));
  nand2 gate2349(.a(s_257), .b(gate427inter3), .O(gate427inter10));
  nor2  gate2350(.a(gate427inter10), .b(gate427inter9), .O(gate427inter11));
  nor2  gate2351(.a(gate427inter11), .b(gate427inter6), .O(gate427inter12));
  nand2 gate2352(.a(gate427inter12), .b(gate427inter1), .O(G1236));
nand2 gate428( .a(G1048), .b(G1144), .O(G1237) );

  xor2  gate1457(.a(G1147), .b(G6), .O(gate429inter0));
  nand2 gate1458(.a(gate429inter0), .b(s_130), .O(gate429inter1));
  and2  gate1459(.a(G1147), .b(G6), .O(gate429inter2));
  inv1  gate1460(.a(s_130), .O(gate429inter3));
  inv1  gate1461(.a(s_131), .O(gate429inter4));
  nand2 gate1462(.a(gate429inter4), .b(gate429inter3), .O(gate429inter5));
  nor2  gate1463(.a(gate429inter5), .b(gate429inter2), .O(gate429inter6));
  inv1  gate1464(.a(G6), .O(gate429inter7));
  inv1  gate1465(.a(G1147), .O(gate429inter8));
  nand2 gate1466(.a(gate429inter8), .b(gate429inter7), .O(gate429inter9));
  nand2 gate1467(.a(s_131), .b(gate429inter3), .O(gate429inter10));
  nor2  gate1468(.a(gate429inter10), .b(gate429inter9), .O(gate429inter11));
  nor2  gate1469(.a(gate429inter11), .b(gate429inter6), .O(gate429inter12));
  nand2 gate1470(.a(gate429inter12), .b(gate429inter1), .O(G1238));
nand2 gate430( .a(G1051), .b(G1147), .O(G1239) );
nand2 gate431( .a(G7), .b(G1150), .O(G1240) );

  xor2  gate981(.a(G1150), .b(G1054), .O(gate432inter0));
  nand2 gate982(.a(gate432inter0), .b(s_62), .O(gate432inter1));
  and2  gate983(.a(G1150), .b(G1054), .O(gate432inter2));
  inv1  gate984(.a(s_62), .O(gate432inter3));
  inv1  gate985(.a(s_63), .O(gate432inter4));
  nand2 gate986(.a(gate432inter4), .b(gate432inter3), .O(gate432inter5));
  nor2  gate987(.a(gate432inter5), .b(gate432inter2), .O(gate432inter6));
  inv1  gate988(.a(G1054), .O(gate432inter7));
  inv1  gate989(.a(G1150), .O(gate432inter8));
  nand2 gate990(.a(gate432inter8), .b(gate432inter7), .O(gate432inter9));
  nand2 gate991(.a(s_63), .b(gate432inter3), .O(gate432inter10));
  nor2  gate992(.a(gate432inter10), .b(gate432inter9), .O(gate432inter11));
  nor2  gate993(.a(gate432inter11), .b(gate432inter6), .O(gate432inter12));
  nand2 gate994(.a(gate432inter12), .b(gate432inter1), .O(G1241));
nand2 gate433( .a(G8), .b(G1153), .O(G1242) );
nand2 gate434( .a(G1057), .b(G1153), .O(G1243) );
nand2 gate435( .a(G9), .b(G1156), .O(G1244) );
nand2 gate436( .a(G1060), .b(G1156), .O(G1245) );

  xor2  gate715(.a(G1159), .b(G10), .O(gate437inter0));
  nand2 gate716(.a(gate437inter0), .b(s_24), .O(gate437inter1));
  and2  gate717(.a(G1159), .b(G10), .O(gate437inter2));
  inv1  gate718(.a(s_24), .O(gate437inter3));
  inv1  gate719(.a(s_25), .O(gate437inter4));
  nand2 gate720(.a(gate437inter4), .b(gate437inter3), .O(gate437inter5));
  nor2  gate721(.a(gate437inter5), .b(gate437inter2), .O(gate437inter6));
  inv1  gate722(.a(G10), .O(gate437inter7));
  inv1  gate723(.a(G1159), .O(gate437inter8));
  nand2 gate724(.a(gate437inter8), .b(gate437inter7), .O(gate437inter9));
  nand2 gate725(.a(s_25), .b(gate437inter3), .O(gate437inter10));
  nor2  gate726(.a(gate437inter10), .b(gate437inter9), .O(gate437inter11));
  nor2  gate727(.a(gate437inter11), .b(gate437inter6), .O(gate437inter12));
  nand2 gate728(.a(gate437inter12), .b(gate437inter1), .O(G1246));

  xor2  gate939(.a(G1159), .b(G1063), .O(gate438inter0));
  nand2 gate940(.a(gate438inter0), .b(s_56), .O(gate438inter1));
  and2  gate941(.a(G1159), .b(G1063), .O(gate438inter2));
  inv1  gate942(.a(s_56), .O(gate438inter3));
  inv1  gate943(.a(s_57), .O(gate438inter4));
  nand2 gate944(.a(gate438inter4), .b(gate438inter3), .O(gate438inter5));
  nor2  gate945(.a(gate438inter5), .b(gate438inter2), .O(gate438inter6));
  inv1  gate946(.a(G1063), .O(gate438inter7));
  inv1  gate947(.a(G1159), .O(gate438inter8));
  nand2 gate948(.a(gate438inter8), .b(gate438inter7), .O(gate438inter9));
  nand2 gate949(.a(s_57), .b(gate438inter3), .O(gate438inter10));
  nor2  gate950(.a(gate438inter10), .b(gate438inter9), .O(gate438inter11));
  nor2  gate951(.a(gate438inter11), .b(gate438inter6), .O(gate438inter12));
  nand2 gate952(.a(gate438inter12), .b(gate438inter1), .O(G1247));
nand2 gate439( .a(G11), .b(G1162), .O(G1248) );
nand2 gate440( .a(G1066), .b(G1162), .O(G1249) );
nand2 gate441( .a(G12), .b(G1165), .O(G1250) );

  xor2  gate2507(.a(G1165), .b(G1069), .O(gate442inter0));
  nand2 gate2508(.a(gate442inter0), .b(s_280), .O(gate442inter1));
  and2  gate2509(.a(G1165), .b(G1069), .O(gate442inter2));
  inv1  gate2510(.a(s_280), .O(gate442inter3));
  inv1  gate2511(.a(s_281), .O(gate442inter4));
  nand2 gate2512(.a(gate442inter4), .b(gate442inter3), .O(gate442inter5));
  nor2  gate2513(.a(gate442inter5), .b(gate442inter2), .O(gate442inter6));
  inv1  gate2514(.a(G1069), .O(gate442inter7));
  inv1  gate2515(.a(G1165), .O(gate442inter8));
  nand2 gate2516(.a(gate442inter8), .b(gate442inter7), .O(gate442inter9));
  nand2 gate2517(.a(s_281), .b(gate442inter3), .O(gate442inter10));
  nor2  gate2518(.a(gate442inter10), .b(gate442inter9), .O(gate442inter11));
  nor2  gate2519(.a(gate442inter11), .b(gate442inter6), .O(gate442inter12));
  nand2 gate2520(.a(gate442inter12), .b(gate442inter1), .O(G1251));
nand2 gate443( .a(G13), .b(G1168), .O(G1252) );
nand2 gate444( .a(G1072), .b(G1168), .O(G1253) );

  xor2  gate2465(.a(G1171), .b(G14), .O(gate445inter0));
  nand2 gate2466(.a(gate445inter0), .b(s_274), .O(gate445inter1));
  and2  gate2467(.a(G1171), .b(G14), .O(gate445inter2));
  inv1  gate2468(.a(s_274), .O(gate445inter3));
  inv1  gate2469(.a(s_275), .O(gate445inter4));
  nand2 gate2470(.a(gate445inter4), .b(gate445inter3), .O(gate445inter5));
  nor2  gate2471(.a(gate445inter5), .b(gate445inter2), .O(gate445inter6));
  inv1  gate2472(.a(G14), .O(gate445inter7));
  inv1  gate2473(.a(G1171), .O(gate445inter8));
  nand2 gate2474(.a(gate445inter8), .b(gate445inter7), .O(gate445inter9));
  nand2 gate2475(.a(s_275), .b(gate445inter3), .O(gate445inter10));
  nor2  gate2476(.a(gate445inter10), .b(gate445inter9), .O(gate445inter11));
  nor2  gate2477(.a(gate445inter11), .b(gate445inter6), .O(gate445inter12));
  nand2 gate2478(.a(gate445inter12), .b(gate445inter1), .O(G1254));

  xor2  gate1737(.a(G1171), .b(G1075), .O(gate446inter0));
  nand2 gate1738(.a(gate446inter0), .b(s_170), .O(gate446inter1));
  and2  gate1739(.a(G1171), .b(G1075), .O(gate446inter2));
  inv1  gate1740(.a(s_170), .O(gate446inter3));
  inv1  gate1741(.a(s_171), .O(gate446inter4));
  nand2 gate1742(.a(gate446inter4), .b(gate446inter3), .O(gate446inter5));
  nor2  gate1743(.a(gate446inter5), .b(gate446inter2), .O(gate446inter6));
  inv1  gate1744(.a(G1075), .O(gate446inter7));
  inv1  gate1745(.a(G1171), .O(gate446inter8));
  nand2 gate1746(.a(gate446inter8), .b(gate446inter7), .O(gate446inter9));
  nand2 gate1747(.a(s_171), .b(gate446inter3), .O(gate446inter10));
  nor2  gate1748(.a(gate446inter10), .b(gate446inter9), .O(gate446inter11));
  nor2  gate1749(.a(gate446inter11), .b(gate446inter6), .O(gate446inter12));
  nand2 gate1750(.a(gate446inter12), .b(gate446inter1), .O(G1255));
nand2 gate447( .a(G15), .b(G1174), .O(G1256) );

  xor2  gate2171(.a(G1174), .b(G1078), .O(gate448inter0));
  nand2 gate2172(.a(gate448inter0), .b(s_232), .O(gate448inter1));
  and2  gate2173(.a(G1174), .b(G1078), .O(gate448inter2));
  inv1  gate2174(.a(s_232), .O(gate448inter3));
  inv1  gate2175(.a(s_233), .O(gate448inter4));
  nand2 gate2176(.a(gate448inter4), .b(gate448inter3), .O(gate448inter5));
  nor2  gate2177(.a(gate448inter5), .b(gate448inter2), .O(gate448inter6));
  inv1  gate2178(.a(G1078), .O(gate448inter7));
  inv1  gate2179(.a(G1174), .O(gate448inter8));
  nand2 gate2180(.a(gate448inter8), .b(gate448inter7), .O(gate448inter9));
  nand2 gate2181(.a(s_233), .b(gate448inter3), .O(gate448inter10));
  nor2  gate2182(.a(gate448inter10), .b(gate448inter9), .O(gate448inter11));
  nor2  gate2183(.a(gate448inter11), .b(gate448inter6), .O(gate448inter12));
  nand2 gate2184(.a(gate448inter12), .b(gate448inter1), .O(G1257));

  xor2  gate2731(.a(G1177), .b(G16), .O(gate449inter0));
  nand2 gate2732(.a(gate449inter0), .b(s_312), .O(gate449inter1));
  and2  gate2733(.a(G1177), .b(G16), .O(gate449inter2));
  inv1  gate2734(.a(s_312), .O(gate449inter3));
  inv1  gate2735(.a(s_313), .O(gate449inter4));
  nand2 gate2736(.a(gate449inter4), .b(gate449inter3), .O(gate449inter5));
  nor2  gate2737(.a(gate449inter5), .b(gate449inter2), .O(gate449inter6));
  inv1  gate2738(.a(G16), .O(gate449inter7));
  inv1  gate2739(.a(G1177), .O(gate449inter8));
  nand2 gate2740(.a(gate449inter8), .b(gate449inter7), .O(gate449inter9));
  nand2 gate2741(.a(s_313), .b(gate449inter3), .O(gate449inter10));
  nor2  gate2742(.a(gate449inter10), .b(gate449inter9), .O(gate449inter11));
  nor2  gate2743(.a(gate449inter11), .b(gate449inter6), .O(gate449inter12));
  nand2 gate2744(.a(gate449inter12), .b(gate449inter1), .O(G1258));
nand2 gate450( .a(G1081), .b(G1177), .O(G1259) );

  xor2  gate1485(.a(G1180), .b(G17), .O(gate451inter0));
  nand2 gate1486(.a(gate451inter0), .b(s_134), .O(gate451inter1));
  and2  gate1487(.a(G1180), .b(G17), .O(gate451inter2));
  inv1  gate1488(.a(s_134), .O(gate451inter3));
  inv1  gate1489(.a(s_135), .O(gate451inter4));
  nand2 gate1490(.a(gate451inter4), .b(gate451inter3), .O(gate451inter5));
  nor2  gate1491(.a(gate451inter5), .b(gate451inter2), .O(gate451inter6));
  inv1  gate1492(.a(G17), .O(gate451inter7));
  inv1  gate1493(.a(G1180), .O(gate451inter8));
  nand2 gate1494(.a(gate451inter8), .b(gate451inter7), .O(gate451inter9));
  nand2 gate1495(.a(s_135), .b(gate451inter3), .O(gate451inter10));
  nor2  gate1496(.a(gate451inter10), .b(gate451inter9), .O(gate451inter11));
  nor2  gate1497(.a(gate451inter11), .b(gate451inter6), .O(gate451inter12));
  nand2 gate1498(.a(gate451inter12), .b(gate451inter1), .O(G1260));

  xor2  gate2689(.a(G1180), .b(G1084), .O(gate452inter0));
  nand2 gate2690(.a(gate452inter0), .b(s_306), .O(gate452inter1));
  and2  gate2691(.a(G1180), .b(G1084), .O(gate452inter2));
  inv1  gate2692(.a(s_306), .O(gate452inter3));
  inv1  gate2693(.a(s_307), .O(gate452inter4));
  nand2 gate2694(.a(gate452inter4), .b(gate452inter3), .O(gate452inter5));
  nor2  gate2695(.a(gate452inter5), .b(gate452inter2), .O(gate452inter6));
  inv1  gate2696(.a(G1084), .O(gate452inter7));
  inv1  gate2697(.a(G1180), .O(gate452inter8));
  nand2 gate2698(.a(gate452inter8), .b(gate452inter7), .O(gate452inter9));
  nand2 gate2699(.a(s_307), .b(gate452inter3), .O(gate452inter10));
  nor2  gate2700(.a(gate452inter10), .b(gate452inter9), .O(gate452inter11));
  nor2  gate2701(.a(gate452inter11), .b(gate452inter6), .O(gate452inter12));
  nand2 gate2702(.a(gate452inter12), .b(gate452inter1), .O(G1261));
nand2 gate453( .a(G18), .b(G1183), .O(G1262) );

  xor2  gate2381(.a(G1183), .b(G1087), .O(gate454inter0));
  nand2 gate2382(.a(gate454inter0), .b(s_262), .O(gate454inter1));
  and2  gate2383(.a(G1183), .b(G1087), .O(gate454inter2));
  inv1  gate2384(.a(s_262), .O(gate454inter3));
  inv1  gate2385(.a(s_263), .O(gate454inter4));
  nand2 gate2386(.a(gate454inter4), .b(gate454inter3), .O(gate454inter5));
  nor2  gate2387(.a(gate454inter5), .b(gate454inter2), .O(gate454inter6));
  inv1  gate2388(.a(G1087), .O(gate454inter7));
  inv1  gate2389(.a(G1183), .O(gate454inter8));
  nand2 gate2390(.a(gate454inter8), .b(gate454inter7), .O(gate454inter9));
  nand2 gate2391(.a(s_263), .b(gate454inter3), .O(gate454inter10));
  nor2  gate2392(.a(gate454inter10), .b(gate454inter9), .O(gate454inter11));
  nor2  gate2393(.a(gate454inter11), .b(gate454inter6), .O(gate454inter12));
  nand2 gate2394(.a(gate454inter12), .b(gate454inter1), .O(G1263));
nand2 gate455( .a(G19), .b(G1186), .O(G1264) );
nand2 gate456( .a(G1090), .b(G1186), .O(G1265) );
nand2 gate457( .a(G20), .b(G1189), .O(G1266) );
nand2 gate458( .a(G1093), .b(G1189), .O(G1267) );
nand2 gate459( .a(G21), .b(G1192), .O(G1268) );

  xor2  gate1471(.a(G1192), .b(G1096), .O(gate460inter0));
  nand2 gate1472(.a(gate460inter0), .b(s_132), .O(gate460inter1));
  and2  gate1473(.a(G1192), .b(G1096), .O(gate460inter2));
  inv1  gate1474(.a(s_132), .O(gate460inter3));
  inv1  gate1475(.a(s_133), .O(gate460inter4));
  nand2 gate1476(.a(gate460inter4), .b(gate460inter3), .O(gate460inter5));
  nor2  gate1477(.a(gate460inter5), .b(gate460inter2), .O(gate460inter6));
  inv1  gate1478(.a(G1096), .O(gate460inter7));
  inv1  gate1479(.a(G1192), .O(gate460inter8));
  nand2 gate1480(.a(gate460inter8), .b(gate460inter7), .O(gate460inter9));
  nand2 gate1481(.a(s_133), .b(gate460inter3), .O(gate460inter10));
  nor2  gate1482(.a(gate460inter10), .b(gate460inter9), .O(gate460inter11));
  nor2  gate1483(.a(gate460inter11), .b(gate460inter6), .O(gate460inter12));
  nand2 gate1484(.a(gate460inter12), .b(gate460inter1), .O(G1269));
nand2 gate461( .a(G22), .b(G1195), .O(G1270) );

  xor2  gate1569(.a(G1195), .b(G1099), .O(gate462inter0));
  nand2 gate1570(.a(gate462inter0), .b(s_146), .O(gate462inter1));
  and2  gate1571(.a(G1195), .b(G1099), .O(gate462inter2));
  inv1  gate1572(.a(s_146), .O(gate462inter3));
  inv1  gate1573(.a(s_147), .O(gate462inter4));
  nand2 gate1574(.a(gate462inter4), .b(gate462inter3), .O(gate462inter5));
  nor2  gate1575(.a(gate462inter5), .b(gate462inter2), .O(gate462inter6));
  inv1  gate1576(.a(G1099), .O(gate462inter7));
  inv1  gate1577(.a(G1195), .O(gate462inter8));
  nand2 gate1578(.a(gate462inter8), .b(gate462inter7), .O(gate462inter9));
  nand2 gate1579(.a(s_147), .b(gate462inter3), .O(gate462inter10));
  nor2  gate1580(.a(gate462inter10), .b(gate462inter9), .O(gate462inter11));
  nor2  gate1581(.a(gate462inter11), .b(gate462inter6), .O(gate462inter12));
  nand2 gate1582(.a(gate462inter12), .b(gate462inter1), .O(G1271));

  xor2  gate2353(.a(G1198), .b(G23), .O(gate463inter0));
  nand2 gate2354(.a(gate463inter0), .b(s_258), .O(gate463inter1));
  and2  gate2355(.a(G1198), .b(G23), .O(gate463inter2));
  inv1  gate2356(.a(s_258), .O(gate463inter3));
  inv1  gate2357(.a(s_259), .O(gate463inter4));
  nand2 gate2358(.a(gate463inter4), .b(gate463inter3), .O(gate463inter5));
  nor2  gate2359(.a(gate463inter5), .b(gate463inter2), .O(gate463inter6));
  inv1  gate2360(.a(G23), .O(gate463inter7));
  inv1  gate2361(.a(G1198), .O(gate463inter8));
  nand2 gate2362(.a(gate463inter8), .b(gate463inter7), .O(gate463inter9));
  nand2 gate2363(.a(s_259), .b(gate463inter3), .O(gate463inter10));
  nor2  gate2364(.a(gate463inter10), .b(gate463inter9), .O(gate463inter11));
  nor2  gate2365(.a(gate463inter11), .b(gate463inter6), .O(gate463inter12));
  nand2 gate2366(.a(gate463inter12), .b(gate463inter1), .O(G1272));
nand2 gate464( .a(G1102), .b(G1198), .O(G1273) );
nand2 gate465( .a(G24), .b(G1201), .O(G1274) );
nand2 gate466( .a(G1105), .b(G1201), .O(G1275) );
nand2 gate467( .a(G25), .b(G1204), .O(G1276) );

  xor2  gate2577(.a(G1204), .b(G1108), .O(gate468inter0));
  nand2 gate2578(.a(gate468inter0), .b(s_290), .O(gate468inter1));
  and2  gate2579(.a(G1204), .b(G1108), .O(gate468inter2));
  inv1  gate2580(.a(s_290), .O(gate468inter3));
  inv1  gate2581(.a(s_291), .O(gate468inter4));
  nand2 gate2582(.a(gate468inter4), .b(gate468inter3), .O(gate468inter5));
  nor2  gate2583(.a(gate468inter5), .b(gate468inter2), .O(gate468inter6));
  inv1  gate2584(.a(G1108), .O(gate468inter7));
  inv1  gate2585(.a(G1204), .O(gate468inter8));
  nand2 gate2586(.a(gate468inter8), .b(gate468inter7), .O(gate468inter9));
  nand2 gate2587(.a(s_291), .b(gate468inter3), .O(gate468inter10));
  nor2  gate2588(.a(gate468inter10), .b(gate468inter9), .O(gate468inter11));
  nor2  gate2589(.a(gate468inter11), .b(gate468inter6), .O(gate468inter12));
  nand2 gate2590(.a(gate468inter12), .b(gate468inter1), .O(G1277));
nand2 gate469( .a(G26), .b(G1207), .O(G1278) );
nand2 gate470( .a(G1111), .b(G1207), .O(G1279) );
nand2 gate471( .a(G27), .b(G1210), .O(G1280) );

  xor2  gate2115(.a(G1210), .b(G1114), .O(gate472inter0));
  nand2 gate2116(.a(gate472inter0), .b(s_224), .O(gate472inter1));
  and2  gate2117(.a(G1210), .b(G1114), .O(gate472inter2));
  inv1  gate2118(.a(s_224), .O(gate472inter3));
  inv1  gate2119(.a(s_225), .O(gate472inter4));
  nand2 gate2120(.a(gate472inter4), .b(gate472inter3), .O(gate472inter5));
  nor2  gate2121(.a(gate472inter5), .b(gate472inter2), .O(gate472inter6));
  inv1  gate2122(.a(G1114), .O(gate472inter7));
  inv1  gate2123(.a(G1210), .O(gate472inter8));
  nand2 gate2124(.a(gate472inter8), .b(gate472inter7), .O(gate472inter9));
  nand2 gate2125(.a(s_225), .b(gate472inter3), .O(gate472inter10));
  nor2  gate2126(.a(gate472inter10), .b(gate472inter9), .O(gate472inter11));
  nor2  gate2127(.a(gate472inter11), .b(gate472inter6), .O(gate472inter12));
  nand2 gate2128(.a(gate472inter12), .b(gate472inter1), .O(G1281));

  xor2  gate2031(.a(G1213), .b(G28), .O(gate473inter0));
  nand2 gate2032(.a(gate473inter0), .b(s_212), .O(gate473inter1));
  and2  gate2033(.a(G1213), .b(G28), .O(gate473inter2));
  inv1  gate2034(.a(s_212), .O(gate473inter3));
  inv1  gate2035(.a(s_213), .O(gate473inter4));
  nand2 gate2036(.a(gate473inter4), .b(gate473inter3), .O(gate473inter5));
  nor2  gate2037(.a(gate473inter5), .b(gate473inter2), .O(gate473inter6));
  inv1  gate2038(.a(G28), .O(gate473inter7));
  inv1  gate2039(.a(G1213), .O(gate473inter8));
  nand2 gate2040(.a(gate473inter8), .b(gate473inter7), .O(gate473inter9));
  nand2 gate2041(.a(s_213), .b(gate473inter3), .O(gate473inter10));
  nor2  gate2042(.a(gate473inter10), .b(gate473inter9), .O(gate473inter11));
  nor2  gate2043(.a(gate473inter11), .b(gate473inter6), .O(gate473inter12));
  nand2 gate2044(.a(gate473inter12), .b(gate473inter1), .O(G1282));

  xor2  gate2059(.a(G1213), .b(G1117), .O(gate474inter0));
  nand2 gate2060(.a(gate474inter0), .b(s_216), .O(gate474inter1));
  and2  gate2061(.a(G1213), .b(G1117), .O(gate474inter2));
  inv1  gate2062(.a(s_216), .O(gate474inter3));
  inv1  gate2063(.a(s_217), .O(gate474inter4));
  nand2 gate2064(.a(gate474inter4), .b(gate474inter3), .O(gate474inter5));
  nor2  gate2065(.a(gate474inter5), .b(gate474inter2), .O(gate474inter6));
  inv1  gate2066(.a(G1117), .O(gate474inter7));
  inv1  gate2067(.a(G1213), .O(gate474inter8));
  nand2 gate2068(.a(gate474inter8), .b(gate474inter7), .O(gate474inter9));
  nand2 gate2069(.a(s_217), .b(gate474inter3), .O(gate474inter10));
  nor2  gate2070(.a(gate474inter10), .b(gate474inter9), .O(gate474inter11));
  nor2  gate2071(.a(gate474inter11), .b(gate474inter6), .O(gate474inter12));
  nand2 gate2072(.a(gate474inter12), .b(gate474inter1), .O(G1283));

  xor2  gate2297(.a(G1216), .b(G29), .O(gate475inter0));
  nand2 gate2298(.a(gate475inter0), .b(s_250), .O(gate475inter1));
  and2  gate2299(.a(G1216), .b(G29), .O(gate475inter2));
  inv1  gate2300(.a(s_250), .O(gate475inter3));
  inv1  gate2301(.a(s_251), .O(gate475inter4));
  nand2 gate2302(.a(gate475inter4), .b(gate475inter3), .O(gate475inter5));
  nor2  gate2303(.a(gate475inter5), .b(gate475inter2), .O(gate475inter6));
  inv1  gate2304(.a(G29), .O(gate475inter7));
  inv1  gate2305(.a(G1216), .O(gate475inter8));
  nand2 gate2306(.a(gate475inter8), .b(gate475inter7), .O(gate475inter9));
  nand2 gate2307(.a(s_251), .b(gate475inter3), .O(gate475inter10));
  nor2  gate2308(.a(gate475inter10), .b(gate475inter9), .O(gate475inter11));
  nor2  gate2309(.a(gate475inter11), .b(gate475inter6), .O(gate475inter12));
  nand2 gate2310(.a(gate475inter12), .b(gate475inter1), .O(G1284));
nand2 gate476( .a(G1120), .b(G1216), .O(G1285) );
nand2 gate477( .a(G30), .b(G1219), .O(G1286) );
nand2 gate478( .a(G1123), .b(G1219), .O(G1287) );
nand2 gate479( .a(G31), .b(G1222), .O(G1288) );
nand2 gate480( .a(G1126), .b(G1222), .O(G1289) );
nand2 gate481( .a(G32), .b(G1225), .O(G1290) );
nand2 gate482( .a(G1129), .b(G1225), .O(G1291) );
nand2 gate483( .a(G1228), .b(G1229), .O(G1292) );

  xor2  gate785(.a(G1231), .b(G1230), .O(gate484inter0));
  nand2 gate786(.a(gate484inter0), .b(s_34), .O(gate484inter1));
  and2  gate787(.a(G1231), .b(G1230), .O(gate484inter2));
  inv1  gate788(.a(s_34), .O(gate484inter3));
  inv1  gate789(.a(s_35), .O(gate484inter4));
  nand2 gate790(.a(gate484inter4), .b(gate484inter3), .O(gate484inter5));
  nor2  gate791(.a(gate484inter5), .b(gate484inter2), .O(gate484inter6));
  inv1  gate792(.a(G1230), .O(gate484inter7));
  inv1  gate793(.a(G1231), .O(gate484inter8));
  nand2 gate794(.a(gate484inter8), .b(gate484inter7), .O(gate484inter9));
  nand2 gate795(.a(s_35), .b(gate484inter3), .O(gate484inter10));
  nor2  gate796(.a(gate484inter10), .b(gate484inter9), .O(gate484inter11));
  nor2  gate797(.a(gate484inter11), .b(gate484inter6), .O(gate484inter12));
  nand2 gate798(.a(gate484inter12), .b(gate484inter1), .O(G1293));

  xor2  gate2493(.a(G1233), .b(G1232), .O(gate485inter0));
  nand2 gate2494(.a(gate485inter0), .b(s_278), .O(gate485inter1));
  and2  gate2495(.a(G1233), .b(G1232), .O(gate485inter2));
  inv1  gate2496(.a(s_278), .O(gate485inter3));
  inv1  gate2497(.a(s_279), .O(gate485inter4));
  nand2 gate2498(.a(gate485inter4), .b(gate485inter3), .O(gate485inter5));
  nor2  gate2499(.a(gate485inter5), .b(gate485inter2), .O(gate485inter6));
  inv1  gate2500(.a(G1232), .O(gate485inter7));
  inv1  gate2501(.a(G1233), .O(gate485inter8));
  nand2 gate2502(.a(gate485inter8), .b(gate485inter7), .O(gate485inter9));
  nand2 gate2503(.a(s_279), .b(gate485inter3), .O(gate485inter10));
  nor2  gate2504(.a(gate485inter10), .b(gate485inter9), .O(gate485inter11));
  nor2  gate2505(.a(gate485inter11), .b(gate485inter6), .O(gate485inter12));
  nand2 gate2506(.a(gate485inter12), .b(gate485inter1), .O(G1294));

  xor2  gate2675(.a(G1235), .b(G1234), .O(gate486inter0));
  nand2 gate2676(.a(gate486inter0), .b(s_304), .O(gate486inter1));
  and2  gate2677(.a(G1235), .b(G1234), .O(gate486inter2));
  inv1  gate2678(.a(s_304), .O(gate486inter3));
  inv1  gate2679(.a(s_305), .O(gate486inter4));
  nand2 gate2680(.a(gate486inter4), .b(gate486inter3), .O(gate486inter5));
  nor2  gate2681(.a(gate486inter5), .b(gate486inter2), .O(gate486inter6));
  inv1  gate2682(.a(G1234), .O(gate486inter7));
  inv1  gate2683(.a(G1235), .O(gate486inter8));
  nand2 gate2684(.a(gate486inter8), .b(gate486inter7), .O(gate486inter9));
  nand2 gate2685(.a(s_305), .b(gate486inter3), .O(gate486inter10));
  nor2  gate2686(.a(gate486inter10), .b(gate486inter9), .O(gate486inter11));
  nor2  gate2687(.a(gate486inter11), .b(gate486inter6), .O(gate486inter12));
  nand2 gate2688(.a(gate486inter12), .b(gate486inter1), .O(G1295));

  xor2  gate2717(.a(G1237), .b(G1236), .O(gate487inter0));
  nand2 gate2718(.a(gate487inter0), .b(s_310), .O(gate487inter1));
  and2  gate2719(.a(G1237), .b(G1236), .O(gate487inter2));
  inv1  gate2720(.a(s_310), .O(gate487inter3));
  inv1  gate2721(.a(s_311), .O(gate487inter4));
  nand2 gate2722(.a(gate487inter4), .b(gate487inter3), .O(gate487inter5));
  nor2  gate2723(.a(gate487inter5), .b(gate487inter2), .O(gate487inter6));
  inv1  gate2724(.a(G1236), .O(gate487inter7));
  inv1  gate2725(.a(G1237), .O(gate487inter8));
  nand2 gate2726(.a(gate487inter8), .b(gate487inter7), .O(gate487inter9));
  nand2 gate2727(.a(s_311), .b(gate487inter3), .O(gate487inter10));
  nor2  gate2728(.a(gate487inter10), .b(gate487inter9), .O(gate487inter11));
  nor2  gate2729(.a(gate487inter11), .b(gate487inter6), .O(gate487inter12));
  nand2 gate2730(.a(gate487inter12), .b(gate487inter1), .O(G1296));

  xor2  gate1625(.a(G1239), .b(G1238), .O(gate488inter0));
  nand2 gate1626(.a(gate488inter0), .b(s_154), .O(gate488inter1));
  and2  gate1627(.a(G1239), .b(G1238), .O(gate488inter2));
  inv1  gate1628(.a(s_154), .O(gate488inter3));
  inv1  gate1629(.a(s_155), .O(gate488inter4));
  nand2 gate1630(.a(gate488inter4), .b(gate488inter3), .O(gate488inter5));
  nor2  gate1631(.a(gate488inter5), .b(gate488inter2), .O(gate488inter6));
  inv1  gate1632(.a(G1238), .O(gate488inter7));
  inv1  gate1633(.a(G1239), .O(gate488inter8));
  nand2 gate1634(.a(gate488inter8), .b(gate488inter7), .O(gate488inter9));
  nand2 gate1635(.a(s_155), .b(gate488inter3), .O(gate488inter10));
  nor2  gate1636(.a(gate488inter10), .b(gate488inter9), .O(gate488inter11));
  nor2  gate1637(.a(gate488inter11), .b(gate488inter6), .O(gate488inter12));
  nand2 gate1638(.a(gate488inter12), .b(gate488inter1), .O(G1297));
nand2 gate489( .a(G1240), .b(G1241), .O(G1298) );

  xor2  gate2409(.a(G1243), .b(G1242), .O(gate490inter0));
  nand2 gate2410(.a(gate490inter0), .b(s_266), .O(gate490inter1));
  and2  gate2411(.a(G1243), .b(G1242), .O(gate490inter2));
  inv1  gate2412(.a(s_266), .O(gate490inter3));
  inv1  gate2413(.a(s_267), .O(gate490inter4));
  nand2 gate2414(.a(gate490inter4), .b(gate490inter3), .O(gate490inter5));
  nor2  gate2415(.a(gate490inter5), .b(gate490inter2), .O(gate490inter6));
  inv1  gate2416(.a(G1242), .O(gate490inter7));
  inv1  gate2417(.a(G1243), .O(gate490inter8));
  nand2 gate2418(.a(gate490inter8), .b(gate490inter7), .O(gate490inter9));
  nand2 gate2419(.a(s_267), .b(gate490inter3), .O(gate490inter10));
  nor2  gate2420(.a(gate490inter10), .b(gate490inter9), .O(gate490inter11));
  nor2  gate2421(.a(gate490inter11), .b(gate490inter6), .O(gate490inter12));
  nand2 gate2422(.a(gate490inter12), .b(gate490inter1), .O(G1299));

  xor2  gate2311(.a(G1245), .b(G1244), .O(gate491inter0));
  nand2 gate2312(.a(gate491inter0), .b(s_252), .O(gate491inter1));
  and2  gate2313(.a(G1245), .b(G1244), .O(gate491inter2));
  inv1  gate2314(.a(s_252), .O(gate491inter3));
  inv1  gate2315(.a(s_253), .O(gate491inter4));
  nand2 gate2316(.a(gate491inter4), .b(gate491inter3), .O(gate491inter5));
  nor2  gate2317(.a(gate491inter5), .b(gate491inter2), .O(gate491inter6));
  inv1  gate2318(.a(G1244), .O(gate491inter7));
  inv1  gate2319(.a(G1245), .O(gate491inter8));
  nand2 gate2320(.a(gate491inter8), .b(gate491inter7), .O(gate491inter9));
  nand2 gate2321(.a(s_253), .b(gate491inter3), .O(gate491inter10));
  nor2  gate2322(.a(gate491inter10), .b(gate491inter9), .O(gate491inter11));
  nor2  gate2323(.a(gate491inter11), .b(gate491inter6), .O(gate491inter12));
  nand2 gate2324(.a(gate491inter12), .b(gate491inter1), .O(G1300));

  xor2  gate953(.a(G1247), .b(G1246), .O(gate492inter0));
  nand2 gate954(.a(gate492inter0), .b(s_58), .O(gate492inter1));
  and2  gate955(.a(G1247), .b(G1246), .O(gate492inter2));
  inv1  gate956(.a(s_58), .O(gate492inter3));
  inv1  gate957(.a(s_59), .O(gate492inter4));
  nand2 gate958(.a(gate492inter4), .b(gate492inter3), .O(gate492inter5));
  nor2  gate959(.a(gate492inter5), .b(gate492inter2), .O(gate492inter6));
  inv1  gate960(.a(G1246), .O(gate492inter7));
  inv1  gate961(.a(G1247), .O(gate492inter8));
  nand2 gate962(.a(gate492inter8), .b(gate492inter7), .O(gate492inter9));
  nand2 gate963(.a(s_59), .b(gate492inter3), .O(gate492inter10));
  nor2  gate964(.a(gate492inter10), .b(gate492inter9), .O(gate492inter11));
  nor2  gate965(.a(gate492inter11), .b(gate492inter6), .O(gate492inter12));
  nand2 gate966(.a(gate492inter12), .b(gate492inter1), .O(G1301));

  xor2  gate1905(.a(G1249), .b(G1248), .O(gate493inter0));
  nand2 gate1906(.a(gate493inter0), .b(s_194), .O(gate493inter1));
  and2  gate1907(.a(G1249), .b(G1248), .O(gate493inter2));
  inv1  gate1908(.a(s_194), .O(gate493inter3));
  inv1  gate1909(.a(s_195), .O(gate493inter4));
  nand2 gate1910(.a(gate493inter4), .b(gate493inter3), .O(gate493inter5));
  nor2  gate1911(.a(gate493inter5), .b(gate493inter2), .O(gate493inter6));
  inv1  gate1912(.a(G1248), .O(gate493inter7));
  inv1  gate1913(.a(G1249), .O(gate493inter8));
  nand2 gate1914(.a(gate493inter8), .b(gate493inter7), .O(gate493inter9));
  nand2 gate1915(.a(s_195), .b(gate493inter3), .O(gate493inter10));
  nor2  gate1916(.a(gate493inter10), .b(gate493inter9), .O(gate493inter11));
  nor2  gate1917(.a(gate493inter11), .b(gate493inter6), .O(gate493inter12));
  nand2 gate1918(.a(gate493inter12), .b(gate493inter1), .O(G1302));
nand2 gate494( .a(G1250), .b(G1251), .O(G1303) );

  xor2  gate2703(.a(G1253), .b(G1252), .O(gate495inter0));
  nand2 gate2704(.a(gate495inter0), .b(s_308), .O(gate495inter1));
  and2  gate2705(.a(G1253), .b(G1252), .O(gate495inter2));
  inv1  gate2706(.a(s_308), .O(gate495inter3));
  inv1  gate2707(.a(s_309), .O(gate495inter4));
  nand2 gate2708(.a(gate495inter4), .b(gate495inter3), .O(gate495inter5));
  nor2  gate2709(.a(gate495inter5), .b(gate495inter2), .O(gate495inter6));
  inv1  gate2710(.a(G1252), .O(gate495inter7));
  inv1  gate2711(.a(G1253), .O(gate495inter8));
  nand2 gate2712(.a(gate495inter8), .b(gate495inter7), .O(gate495inter9));
  nand2 gate2713(.a(s_309), .b(gate495inter3), .O(gate495inter10));
  nor2  gate2714(.a(gate495inter10), .b(gate495inter9), .O(gate495inter11));
  nor2  gate2715(.a(gate495inter11), .b(gate495inter6), .O(gate495inter12));
  nand2 gate2716(.a(gate495inter12), .b(gate495inter1), .O(G1304));
nand2 gate496( .a(G1254), .b(G1255), .O(G1305) );
nand2 gate497( .a(G1256), .b(G1257), .O(G1306) );
nand2 gate498( .a(G1258), .b(G1259), .O(G1307) );
nand2 gate499( .a(G1260), .b(G1261), .O(G1308) );

  xor2  gate1765(.a(G1263), .b(G1262), .O(gate500inter0));
  nand2 gate1766(.a(gate500inter0), .b(s_174), .O(gate500inter1));
  and2  gate1767(.a(G1263), .b(G1262), .O(gate500inter2));
  inv1  gate1768(.a(s_174), .O(gate500inter3));
  inv1  gate1769(.a(s_175), .O(gate500inter4));
  nand2 gate1770(.a(gate500inter4), .b(gate500inter3), .O(gate500inter5));
  nor2  gate1771(.a(gate500inter5), .b(gate500inter2), .O(gate500inter6));
  inv1  gate1772(.a(G1262), .O(gate500inter7));
  inv1  gate1773(.a(G1263), .O(gate500inter8));
  nand2 gate1774(.a(gate500inter8), .b(gate500inter7), .O(gate500inter9));
  nand2 gate1775(.a(s_175), .b(gate500inter3), .O(gate500inter10));
  nor2  gate1776(.a(gate500inter10), .b(gate500inter9), .O(gate500inter11));
  nor2  gate1777(.a(gate500inter11), .b(gate500inter6), .O(gate500inter12));
  nand2 gate1778(.a(gate500inter12), .b(gate500inter1), .O(G1309));
nand2 gate501( .a(G1264), .b(G1265), .O(G1310) );

  xor2  gate1247(.a(G1267), .b(G1266), .O(gate502inter0));
  nand2 gate1248(.a(gate502inter0), .b(s_100), .O(gate502inter1));
  and2  gate1249(.a(G1267), .b(G1266), .O(gate502inter2));
  inv1  gate1250(.a(s_100), .O(gate502inter3));
  inv1  gate1251(.a(s_101), .O(gate502inter4));
  nand2 gate1252(.a(gate502inter4), .b(gate502inter3), .O(gate502inter5));
  nor2  gate1253(.a(gate502inter5), .b(gate502inter2), .O(gate502inter6));
  inv1  gate1254(.a(G1266), .O(gate502inter7));
  inv1  gate1255(.a(G1267), .O(gate502inter8));
  nand2 gate1256(.a(gate502inter8), .b(gate502inter7), .O(gate502inter9));
  nand2 gate1257(.a(s_101), .b(gate502inter3), .O(gate502inter10));
  nor2  gate1258(.a(gate502inter10), .b(gate502inter9), .O(gate502inter11));
  nor2  gate1259(.a(gate502inter11), .b(gate502inter6), .O(gate502inter12));
  nand2 gate1260(.a(gate502inter12), .b(gate502inter1), .O(G1311));
nand2 gate503( .a(G1268), .b(G1269), .O(G1312) );
nand2 gate504( .a(G1270), .b(G1271), .O(G1313) );
nand2 gate505( .a(G1272), .b(G1273), .O(G1314) );

  xor2  gate2325(.a(G1275), .b(G1274), .O(gate506inter0));
  nand2 gate2326(.a(gate506inter0), .b(s_254), .O(gate506inter1));
  and2  gate2327(.a(G1275), .b(G1274), .O(gate506inter2));
  inv1  gate2328(.a(s_254), .O(gate506inter3));
  inv1  gate2329(.a(s_255), .O(gate506inter4));
  nand2 gate2330(.a(gate506inter4), .b(gate506inter3), .O(gate506inter5));
  nor2  gate2331(.a(gate506inter5), .b(gate506inter2), .O(gate506inter6));
  inv1  gate2332(.a(G1274), .O(gate506inter7));
  inv1  gate2333(.a(G1275), .O(gate506inter8));
  nand2 gate2334(.a(gate506inter8), .b(gate506inter7), .O(gate506inter9));
  nand2 gate2335(.a(s_255), .b(gate506inter3), .O(gate506inter10));
  nor2  gate2336(.a(gate506inter10), .b(gate506inter9), .O(gate506inter11));
  nor2  gate2337(.a(gate506inter11), .b(gate506inter6), .O(gate506inter12));
  nand2 gate2338(.a(gate506inter12), .b(gate506inter1), .O(G1315));
nand2 gate507( .a(G1276), .b(G1277), .O(G1316) );
nand2 gate508( .a(G1278), .b(G1279), .O(G1317) );

  xor2  gate617(.a(G1281), .b(G1280), .O(gate509inter0));
  nand2 gate618(.a(gate509inter0), .b(s_10), .O(gate509inter1));
  and2  gate619(.a(G1281), .b(G1280), .O(gate509inter2));
  inv1  gate620(.a(s_10), .O(gate509inter3));
  inv1  gate621(.a(s_11), .O(gate509inter4));
  nand2 gate622(.a(gate509inter4), .b(gate509inter3), .O(gate509inter5));
  nor2  gate623(.a(gate509inter5), .b(gate509inter2), .O(gate509inter6));
  inv1  gate624(.a(G1280), .O(gate509inter7));
  inv1  gate625(.a(G1281), .O(gate509inter8));
  nand2 gate626(.a(gate509inter8), .b(gate509inter7), .O(gate509inter9));
  nand2 gate627(.a(s_11), .b(gate509inter3), .O(gate509inter10));
  nor2  gate628(.a(gate509inter10), .b(gate509inter9), .O(gate509inter11));
  nor2  gate629(.a(gate509inter11), .b(gate509inter6), .O(gate509inter12));
  nand2 gate630(.a(gate509inter12), .b(gate509inter1), .O(G1318));
nand2 gate510( .a(G1282), .b(G1283), .O(G1319) );
nand2 gate511( .a(G1284), .b(G1285), .O(G1320) );

  xor2  gate2815(.a(G1287), .b(G1286), .O(gate512inter0));
  nand2 gate2816(.a(gate512inter0), .b(s_324), .O(gate512inter1));
  and2  gate2817(.a(G1287), .b(G1286), .O(gate512inter2));
  inv1  gate2818(.a(s_324), .O(gate512inter3));
  inv1  gate2819(.a(s_325), .O(gate512inter4));
  nand2 gate2820(.a(gate512inter4), .b(gate512inter3), .O(gate512inter5));
  nor2  gate2821(.a(gate512inter5), .b(gate512inter2), .O(gate512inter6));
  inv1  gate2822(.a(G1286), .O(gate512inter7));
  inv1  gate2823(.a(G1287), .O(gate512inter8));
  nand2 gate2824(.a(gate512inter8), .b(gate512inter7), .O(gate512inter9));
  nand2 gate2825(.a(s_325), .b(gate512inter3), .O(gate512inter10));
  nor2  gate2826(.a(gate512inter10), .b(gate512inter9), .O(gate512inter11));
  nor2  gate2827(.a(gate512inter11), .b(gate512inter6), .O(gate512inter12));
  nand2 gate2828(.a(gate512inter12), .b(gate512inter1), .O(G1321));
nand2 gate513( .a(G1288), .b(G1289), .O(G1322) );
nand2 gate514( .a(G1290), .b(G1291), .O(G1323) );
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule